-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qCqweJcc6zsP8MeHYacR9I5hc0gpY1h5MkISUQ5A+1l6FLVwrP/jJjzp5/0padrAdKx5xFurvETh
UWcMo3+v8r3AHMzsJq3+sfeIvYoqmkoHVSdBIwQTwMV78o9FAumYI0cwLdMG/kl9iyvtLYBCJAnF
bcJTji3+zDV26SDbkREoIGLpBHVeUGqLQHIqSi/SQOyXGJDyPiBwD29FtC2wj60p/1CIfjG4im41
W2vUyZKbD7bntoDpMHK3l62OYGGP9NPHsUdishxSdmBpeu76lIVMtrlHulbvA7RzOWKR15quHEe8
bX0N4+BOXQ2C+jd8DLfndlRnHi8P2fPJIqmzxA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
UQMLVnhWFQM2yzX4xwgjY/68o4qk+V/TaNjcTDzfoiHJBp34seVwV9zWGAN3ycIK9eGz3MlrIYEy
5Cv0hh4Og3HrdZ0BkUfJ6eXlR2BI3NauMfXxTInuyeceLk5oFBd37X3pzwfdgbe8U8VsqqOX8n8F
o5/rKschSxFCY+etZ9w0DKHXX142Iv0dASPv4vF4LtzkaIUDONO+ENKKhFsNFnVbeSvQCWGGsjCf
kd9jCnaTjBVXa2nv2pGV42M0S96dtCUeZN/oM67idOUF7t2Rr3exWfWRlbo/VvJjjUWVo+BUUxFM
jzg0bxKer6UNZ+Rw/pwP7GPLRKtkHVmqi3oT0Ch3h25c9K46dLpgwQmlMZlnlPusBNL7apye5r8M
vuaaNcREl1iXGjyaV99W3WePyVZKLTRgWgR7eI8stH6cAe0ueCUTknDP0u/2KG+QoyfE0UAkyecG
FYvrgOKwJQJk5E0EKfYD5qdIbRyGoaH2ucs31CN4fYZGDzKUXnsDt8HLli8aHqkaIdnETF0njt8M
QrkXBcSYm+YaTJXKa3HZ61V6VPB6yRJVA6mFq1X4o6wik6H7QOZr0iqaqky0TxHarOqkjlNMVSNF
g+GqJcPRTYNS+PK1BpDeLkex504RotZp5iSvYJ8MOvlXv/38Ch6bZMw27opf6/Q9/mGDmMlA9tQH
aE9Fc5z2FOIpimC2Apnirn18Zl7+Uhdnb+qb1xVVj6GGxp/PK4ubufJy4Kfu+/Eb2gsZOUb75EZ9
H/xbk2X5pgp+5e665MV8aO7ZiovdI12P4nbGoxdQ6d6qA/GAWb+3sux6u1NE5ycTCcgpphbcska/
nOnF9eMNxKDUJy3cSGlFxSRA/OB1j35JFQfpg7+3IpgJnCZPMMnZRt5ZV4fP4/j6VT/vBglCqP4E
IR1rXZsKxCt6AWe8ElFSbq3xbmRic7bbOZ0pWOXy6pJD0w7C6CtlY0HibjgKChvWWEv6ItxP3juk
HPJvhOQL5/ihEEYFmBbzaMWbpJStcHtf6sQd3tH3JzBGVLF4xSvUpR5E+AHRruWYUW95laWiaSXs
eOI0XNCDMf5zGKaWkICdla1P87ghTx/L1pG/8a/P6VVK6x6FLRtDN2Tsszvk6Ge1sdxoKNEYeIZU
uB24GQvHHIeUUBZXgJw6xZ27XchxPK6triqa4K0w4u9N2B8UZXKMIylyJxam6oeRkRdDjAmPyoDn
sg410CCsTbuZerfasSqJzDM0xHah351Z6mWmxK5twKmzkJMS9XZcIz+6fTUar1Xvlzq7Rt/xmTMK
oGi/thtzgomTW4b4RPkxzVj9eIhJkNgl9TcRBgo1HL5TtJ0JNCoUWq43zReNnWnQcDx1wxlFWvS5
vYA6WBr9Ss7nC9ItKiXhF7Id6g5d5R1s/1tqROyKZbDsySFmzaoLwv435HR5EnO02v7vrVomN6OB
QFggfeLXFmJxc2zN3OQY+6zAxNOJ9O+XWzZMz3iNAcaqnZkYgFlIcrqoxMZbrQQ655twlDVB6t2W
LAwN0Ew6MT2thD+QAJ6OutRoV2Xx35ijD4PjkehWo28TaNp/Xqzedv90qIxe75kV99i6HbCUj1Wu
labSWjIy7xRzkh1zJb1Ta7VkPIO+sFEHIa+7Bslhc8MfUq5oU1rhby3a7drztlY/QvqkzOun0cy0
fegmx+0EzCQxmzNJMrF8NL3xrKg1qnc/eo2AlXdTkvW2vUMP549PdpLxQ806KIArbV1j5HyYLZQr
4OSm2+g6NJdcD8dUeZpLSVt7lII67WBNjlCnDkPASzXFfTQQi3y0CB4CzKTbiumIJ5QO3a2rYi7p
keesha3CgpN15bvWk8MkHPMKA2r7iMz1nyPnTGw0FbCSGSy11NAd+jUxw4KS9WlVYVBv1p0NyiFQ
MJlvVWLEFGeHmN4FoXiJS3iq2OTBVuukFxL63OZ6ja9Bb3QzsHOehFrgz/MmkmoNvLrDURfWA0nL
h91d5f8/KFKWGwiJd13+R4nrY/LEzMI2zv4IGvIxTORE5bFSA/DP6SJSQ6VKXigyetsX//LuT9tY
5utGdpvQFptDtlP7Fi8uSCMJ0R7uPJrVdLVa1X9GwGZD/CeGjP1lj3touC5sTjkNLMHUg5outhOu
Lr/l1lIcGrPzTQeKbWTICbDSPUNQJ2Ww40Id5dMKmahjGjeVPIa96F8L2JNTf4DCc4qyz462xTJl
UtWfgiY1bTkZDDGMM5Apq63GRzDwnBiXECOTWjXoTJ2DqBH9Ua50XTiMQcJu/JIGABOF7tZieDoo
esKMvfQNU7WXx/SfFrJpYd4DrPIXk3BKUZVETTYwpwJJPCLUFRqkHML3760q2xPxUy2V71xPdENz
NfO6/DcxypVYwkzlibQzf4LuoSbFZOn58V3Gv8ppZixFKQvHPJqfkyqYB1AOD4HrmswC0RjR58NH
13dYIAGNxYLj+f22rUQw23iEwcDmdGxNOov918Y69QFQGgEHBZ45zybCLIAepyd4sugjWOiwhAfq
46cWY6TVGMUadoqaHTJxcabAiiMP6Gqk6rwetB2MVbbYOmUx5EXtEg/KBuJLkxS5OOGIbV4qZgH9
2Xtseb63uP8SyvjW7awDSJv6f943VCQ4pkTV15+gunz4CyIv89Plx9XiSUHO6sqiCDfUfZqjmoDE
81CYJKQU/wtMQ6bT0SzeQs9FfBBeIVr9iGRhXM4Eqo8/I8+15CZyXqZpYNzdYC9U+ofpTZVHSOBU
6S40b/5659DjM6BkPDHI0zQ9l0ZA9Y3eftq34odmefyFzk92iJpkc9+1uH34Da/Z1tAIZTOZU7s7
ycTtGJKXOtjA6XRf2c43K07AbTElGbES7Tj5zldmMONkcNXNQ3/0j4ExPT1Q/s8f9yu+Dw3MZCom
oqGcwBkqSi0CtYp+CIRfTvCSghVhPa6hy/ptTri/AYK5UCBIU6/hz15ZQIYrZki4mAk1+K8j2ZKo
Z1mjrv7Crfg513e95w7pYDWQ+zNoEYokZkicZkcWZtDjZGHqJ/0ouCW8mN8V3cy/VJWaYU8Smz6X
fMRLzGGtAp61v87Aevns0jr3u+NHc2QvocdPwdRRr7zFiSqKItm3yVSi5LUJd+mc+PQqBMIKxgOv
1XkyBNq6rSvSCUQ0/devWOQICXIyvpmNZJKJ9ltEBY5pygaq98nnDdZml5F/Wzapge/592S+ZsuV
wsQ8F4LgqfKuNiZpjCjpY7nemt3F2Wo62pm2NZWbuNOip/j5tXJrog6g5JZxkSOYUC3ITXz1uwxl
BUuvXiw5FQx2clRexjCZuN4gQmsPeLKOHNci/6dDZQw05xjFDeA8jJWOZBYJkOPyEh8SNKUWLqft
jt+bEX+4Bor48Xt399KrSm0o/YPOzwTGVzluLkaEWBIACNG0WfUOBq+E9vr2jBtfqdi2FV5tsh6O
bFY0aGV5RNisMTgdaTAtIGHycL12InmDH6Kh1NOqSd/Yp9hxPWcvwt4kklRpMJUXY4CUmDcBhZq9
5hahwfCkdA/4w6atqu54WKj4nVh+IYwk8sxOv9KYKbvvUv0EInGa1eT81k98bXncVsPOLZmrIBVk
8zj9TIom+q3x8qkyennw16DR9OU164hWNJbRJ8pytTkTElEba9vbYxzJ8sY9WUkq2V0CCDUNVKFJ
HJhj2jb7ga2qhZmypmwFZq32UW9MSCT6jwztdkJ9ljQDHwdjm0hHzPDEEODYAlgnG+IB4gTngTCT
DC/IfnpPl1+FEyybo4FyqkNudSR1CfCw/lTUU9torgXidCWJMAGUnr7eT+386jfyg2TGEhc2wnI4
LjZJImLSdPj12lFCKY74P1t4iYlZrWkSj5ZbPwhEi91TMz97Cbl17QM73/f3RBtRV8J4UbxcspUv
dTgJIbvov7bqxlAxXSQYn7WrAUYaDs+bM1Z3EoM9/K/MVYkrTadMb45Ft8ZJlmCsw6Djv7e85DoP
dT8OgStecwvXcf8wt1z4PLZScQ/tcK0jeCt6bcIC4uGEjoxdJWJ7cl2M/Xgfa9Gz/sw7l47beTZi
nUmiW1QEvyPa0rCwasFQn9YeAiPi/aoUg9YoP0LNknORdPjSg+uGIIpYhFQ6gqn+X15/kfxxyCgZ
a2F0WIP345auklWxKn2ulnSqEvIqJhkoiT+pSWy+Ld9rCYR+FX1pWxPTVC+H6gkBel2B5PEFtpnH
G4vMWddUxzeGz7rJxih2rxiApb2huGJ8s/8lzOcUS9+Nkc6PysOxzpZ/NPzSi9KxLhl+bvcTwigk
2ob0Tuo/cl9mjjEYoqnePiBdjdkx5//AIUQJ9dcrYtqonY7NGuOniXQvmsOYUo4sBruX9PAH2toy
KXAdgeo0VIrYN7zzQK+32Re+kt0/ZS3NW5dZYfOgb8k/4aHqSRAy4BvdAs+uCjvGdYA7fL40P1HL
wYyqnjyJmVWeIdaNmVlqwYPJpBB5cJk/18sAxPGBYHO6xFCP6TLP/IOxEHstt2FsU4zt/dTZgUc7
wQEH1Qh1bRGqBl0kZnr5VxfKXN77e5c9krLNR4JAJkqEcl9dgclrBd4ic8YoaP0UaSjnd0rt/hSc
zH05joDy8lMwpc+83dU96cS4rO9FgaWI3op2hBTXBhS+4Ba4HwSxCtDEu/h5h3TF2kdh7NtES96i
8KYhIeyQZ14DCOylEi0SJb88woKZEzfnHeaQA6RuR5/+1hrRoLF/MqBWQdhT7J0flPXZv0OnRTHv
9OBePG0FHsCAgoNiIClZdyw9e4ed1IN1dB6k+JT2tKcMOriFS0977q+XEea1wAo3BK9XiyIjucQ9
dO6yWUOr1+Z+sKinQCuNjQ4KgAorcCHa1WskuCUHUgSCejxhhz8U/irO0di8y6rR3aDZoAdnArg3
vrPrFm53udwsxnF/zsmMCJJ2sIbaZWR9pT1qvulRmRvNoM7CK/QcL9NZwPJdJljNE8z+cUXjQ/8L
RR+9I+Tvs2tpGCl4/A9UQdWnrzCSd+cEY4BGBpUeM+PiYGGkgp30r6T+GDGqcCVTX90zVcMy1g/8
TgEcJdtw4Ls/AyMvjL8/649Goe0ApfXdEHuv7AjSBckgLItAZV7zesdcIWtBA3vzk4NcYOUXtOmT
q8C+oTiJsN50Sxku6hp3/vmw3pvI0IBo2i40uOU3z+tiK/JOy1aAAp3XZZgYNTOogd1X1HkHs3Gr
u2Ho5ua6OFe0MbNBn2DiXyoeDR/s8H3QJVW/NJrdaUZF5pFgERygefet36TQQSv356qH2UeaSydM
1ZtM1Tds9vwI9aAgLIA5IldSOSaDMvEa1LQIx0tZenNd+dD4XRePtI375AC+lyluQsObc5/B0ZPR
sK4EwyQvc5ebKuPH0r/LZMjIrvrDhLi3odWLdxfS3d4etcJMWVHcs2lw3Z75xCzXV24faG/PsEoD
ygLEGTy9GAtTomUs/iH3V1efHUCmdejjf4BWQKSyRyKqeXcm3GsbdKZ/eJy8FXiahw/tdnH83b1K
F+5a3c4hz1+/s0e4ex42QpbCBUJC+lJmDjdlPSbr4hSTDac++GLCKuhsLOEfG578AFBJ7a6x8dp9
oXRPaX0/sjprnbJlXYzSBawDPzi72NKpbo2X+4rfpOxiLDPrlvtKnYetEg0dznFpTF3+0eoQXyCz
PTJnGKt0gM5slReqoTf2+jeIsJd2B2vYaL0QusQwbRX+kKJUzT8+u2NAPnhe4XLBdDrRlP7C2l5J
0pMN3wv8ViMyzRIHWka8+4qEVFnZ7cOoyizDFYgp+2SHP0ymHZWq9EDpFhwx0B5T+10UfPdiyS1M
Tlpg+cQU5JtipXlM/sdFdUZhYyl5sHifGgS2bXdiIq84NMf8KhNln5v4PGzR2Tum1mzZN4E2oKLT
hD3J4TTspmO9WJqqf0PHkKq2duIcuDKO/Dgq/xClsjDxWAHXIFyj+JCCSubQIUu35ewWEUR1uDJ8
igGZvLD9oufKdMsn2jbeuPqUNgZhQzeBhLrnbtSJixEZKYYee36sczTII6bdcyA+HD8gYxIVxeCP
UHNowq0Azj44HBO/4pva5dH3/eSL3DTpUsCravX3oX8To88kx2nGEZF3BRdPYjmb9HOmrWSo5P4k
bkVHVIhtQ8NN4ZkOETGUj4D6+OG2KkItLvdmMXR+w0u7g1yo6+F5+aSPTaBhQY6P8BvLMd96oRVt
oIbMptiVG26DP57gYBeDZfbSk9/b7Hx70ZbJu/AcbXYxsYWPvVUePJzZSeabuU7bwIYBc6KpP+3Y
fT6rxZZB7RLfGD9ARQabSEUiltBrgFgJoLNtdghDIEQCKtNir90yD/4p84rztq4LonLTS/zH0hsf
IrjTM9uCdbo6ybxkMMwnPzfc76mISqmeXd5GsY8vAXJp13jrNyQkw+PKTm5uXPLJQ7o1glGibP76
eDxWLkrfw8rz5HY21eV4qPnBxdMQVVny9ZzyzbnTVzzUG7BDfkPUvQMv+fygZWjDfnf26OEfm0QT
HAT+uAtkf1L8DrG1FAOzSJ4Q63YyQ9wqedr0YmQ9cwtZVo54qAMm+JuBrVg7dMaa37l9r9+SyLfm
TQ6WCtki76sOPlIAmd+PF49WbT4SF2N2S2+JjMbhMgCMPSGQ8DYbjTgcCPzyYLlb3Mt94/sajfot
P6ZNEmgH/ln/1/+3DW4F1el07+C5Gwbokk6rdp4iQWzL+3l3v+zLHKk+K8JEqW85nCmZ2msHLfTr
EZdHX1Av4Ob/6W462bgPbC4epLVXYuVsYLL8PUmuvVtUDtu7dUfC3RRbvO2ulltcdMMGFy3UwbSa
CyoF8Gty11S7Zk7ujpQr9wrRSjjHP1u51P7wEi/ald8X8k+kYRVy+rdJKKkBf0cXxtVsQ9FKFbZY
fKQRUM4y3PbgArS285EgriLLtG/OxLCRlcGOSPsKYdlDidk/7fWdTbRVLH2kac/Wyoaxo1/kkQ1m
Ea8JRjHuVRl1HfyNGpSbM37iGOSSzdEqGvjwECxHaNysYI2ihBx983ARkOQlU9UWK7ZaErhUiOy8
YGPMe0SuSoYJwjoZ/TRwtFRZm0Q29dUZ/BL+lZKRIdMxuNuuDarpjngpMIiKvfvt/7/X4saPrilY
mFttlucjwKCOZcDQ4e5OyDkxVQ3tPc4+nH6+HGJ/UdtOd4i8R9yoLQ1OO0IRx8kJXSzOrsi8c1tu
ypIoqqfocAkEOUactnrObnKZYFiC4PoXApsMl3iV68R3jYwaH6rGI/8DE3jIpkVaROLyF+xFXscn
VxlBpVj7CVBgCreUryMlI4tC6WgkW5QGLJZRu9tmPGiOcMB3zm9XcYBFiq+N1av4wRzGmhFfdK5y
gJehnVz21UEF+bzcPKO1JZcmxhorKu/wVyKPA7c0zkjzTYEdHxi1XiEpsxmLxi4/Iy+Cn74hozmn
214pTP6zuvuxh7KMJatFMGmmzzjuCMiNPWZcXOpKwubEXT0QoZ816+XtZiWgI+EVozHB1OAm1jOV
FNn7XyxJVHcWlxjIXkiLr5GjoMXMegIm9SGoguqCsL2HUqhxqHsY2YUXEgz9tHaeWF7nVqBQ3lwO
43Ppiu2rUKcp+EFg78e8Kr43UgmfUFp3DkiwIOXql04bImpPyUMa/DbuNNU7pFnQCiMlu0794f98
YrikdUiNBJEIvaz0lhjjgjXc65VtqxBzUCyw6M98tVeYGhwNaq1p6Jkoy10n//z0p+4yqei84O49
lfR1ZeW9KTqFn3m68022NAqb3EUOb/mo8hlDm4/CTaQhPpJMC5brUttfY91v8mjvxIhy8Eymh3rE
XKZgA0569V3uCFj5BzxpvDAXkAvwLlHlt4SfTTrUmejfaJtVNg2sdY46xfkYN6cNPbXjyj9f7Wjb
KlQRdgtEPz2kSt0H/mebq1yUOUwJtALBZIyejCEJ/KvU+dkBFk/vPGI6MmDGcbtKa6M4OL4T7lW3
2hwD0sEmAUFJEumwglpql+Z6YiHI0C/BOyeOGZpTy6n21dXhZuC0UumcBqFQcIqQHTxEHCdyIfvJ
u66d3IgMnD87ZJZLijfyCrpAf1InsDaLwE29WDm3OaE7Vob9eRMD9R2hlmEaS1whvH5j0aqYDQAZ
4jxlaxGWx9MmpYtk/XH3fZXzLPDSKpo16Xh3ojTU0wPR0gFWod6bGierhSgiQSOAPa6r8VwXr0aK
V6h5hsy9tc8q0bTrpuiqLoyLZ/e9CEikE4L9x8uAQ5NIwA894vhycLG7lTLgsFpYWqFD8RwIk4da
KNaXCtG6z/Huy8CI9IxIlrFANf5xrcBKufDifVqGuNTNPUya8g9fYJLmpdf7OqTfDFOass7cHpaT
AZW43rfIfIFwTDhE67VcG87bKjEhT9BGNUOO91G3b7PhtA2wq33VFramOOUywAdVsv/SxQPaOrOW
tb4dLr5plQCnPMraqAPkhzNZ3dykXMOrECeduUNhZxqbqezE44z8m+oF+rHmn/2KAic+Rpsm3M8d
e/qwjKXDvGDvsjyZoQixfxoj/GUGmPki0qOrPoM1mwNZ0tpujuoZGyk6T40vY9LjAwMxjUMKRfeu
mr9GesJN73pCoQq7IMNJaLZXORt76SHCIOAcALRkHBgscqH/Qyg32AsNW1dnkiidsT+OsU4rrSd+
ApXquzlCFthXKSEWxzoW/gJFeMA0E6Jm8MhSIEfepFG35iEhCB4c7M/3Vxrtw47vvot/nk3UDrXW
0pdW6owa49GQyvNw0Wph9m8ZmOsMTWhfLNDdT0m1pjG7asoN/hjm7OgCoLXHlltya/06dA1OsQh+
QySsS/bwf7/uAngXewwDnotpYHZctnJJlf1UpK7rghNElNOQQtyAD+owOyYcJjFAbiqHTYzrk1IG
ESpaX5xgtNwsGcSx9gh2mJbEXIT4vK8rGDi7hnyHWNdV+d2RiaHCFaZC6ZMnkUo88D98VLbkmhUY
iRfDm+5KELe5IdFjGYxiHjdOAGi0Qn0oTRRNxIdvdnfULTKk2p28DuasgiNMYpk0lcRVOzJRNNzS
WndbNh5DShlRPVLxCJDK9wJXRg9WsseoWJwo9XTEfoEyLuyHeAnxN7GJNeB491X4vELZg6ki7F6u
jDNapMPO6hzltGTKZrFKt/zYptkG9uFd/v1TMNWYxbKuazw0y3wvSnOTEb0xiHM6EDVkygDj9tMZ
BXEU8EWLgEFHHB+ieesn1jy8NzsI0z4nYpL65GHDGgUIamgmpRorDGifYwDjDJL7y+pb4F8mxZop
apDUlp9ekj62M/+KUzDq9ORWclHrjD921gvsK2RMKdwee9qc5oE7RdI9HWaNNn5x5R4Q9OwMSgFU
yNoVxgx3om73kxxIZiqinbThiTboRQDmpDrlTSphhVpAuVGo3sIsgyv8i2QBTf/TROHzhetNJUtV
EBAiHMxY6lOs6//7gnThTy9HXag2HCJM57GLf5L0KhD2ol1ldlijCk/4MgdRgKEYjpX54rirl2UY
O2W6VTbnIEcUe4KIs1qlaqrLutKq0Pin6pz6qwTa1yY68/9P7gHjmhLgLSKhHIzmBK+b4S9kL1hY
rccHITlzV0qCc1g0naF1HUFTjeX4jDaLh4AOjbXxRrdwwck0Mj1Xik65v0F8gGb4LaEIexU4xuUh
FK8YEUasTfz+No40/DveahcMT9tRD0THmq7grTJDzSZqYCgXSV9vHs2mSzZMEh+G5M4qZMR9EGJz
1aSSdBpJHlR6HI5IL3xTqtFYQ6f01Y5LqFEGYmIYndmiNIx9/6D5EP9fjnxhYgMH13HtDNRwd/oN
WvKoyhcIxIxBFMdz168OUBP45QPuPtKkqEkJJvkyAJBs9/AZXXOv1TNrqR3QELypZxuBj9tWblFj
7xj2i6VACR2oiPAOr+cfcCVkg/BoF6ZXinkRljWyNwJ8OFsuxKvyl1NhOAbu0uLAQhfdb9jHiA99
6gmhov1Tvi6uX5o6ASNlw0lMFzq0AEX0eS0+EK2qFNCWsaJsR2YwSnmy+jYzFdmULvYvgOnoY/pO
y9nAAaEtE/uvhLa0R9ZBjHC33b5MkPPlZsBOyiI1XzB6YUNzaJO3DdVQwb85JriXW8Tak+am4IMV
uee8FCzaZig8ASVZEXrZQqBT5JVO3aOwGCj283vldlnb6UkOOett2dtXeJO6T0g2FTsZdVrSOhMR
gJLGunLSE5N6Or4atAfKFWIjKqtPgog0F2c0UJOV2yP7vCEfjeITqMXpjPITooa037uHiwujy8cd
qBb+6RveGAbXW+v36LFaRJoENaRqFauK+NcfphQHIJSfOusjFXVyf2kLSEHNaUtb4MhcUi7VgEPz
Yssl3Mn5taWE9kU8MZaTInyvPzUYqUaGDBx1NDToJj+Vm/CjMTMtp9HWYKvdBWbyefFz29Fi+qyK
lflI1bZ5Mp3u91d0Z+K+aSuauOB4Ldi6Pi3J35cfsmrNNzrUzFL4bIoY8a4UToNIj0hFsWpej1XX
4nipuUiCuHP3eBGQN4QoR+QuAxGnauh/gpUQWeYCeMZnPMtQqmSeqU/l4CEKUGJAfdpjHq57lGWI
vAXdg7be2+44OG4NIoygwVOqEI9rS2ZJGZNXteKg3ys0H+UJ4r0Kn1T/beLv3WrIrxnaz9dlT3tJ
v4EgTHbPIczrEoZCHRpVQM3BkFpWFGoAYJ7wD/KwQqv1TSfswt56CLfFDOF7uGff1LSKvQG9IwQE
pumbCEUoDhO1rUN2fvIMFhK5dahqprK3w/xL/y0uR/XP+G4WDbevRJL2yDzji+7paV5YWqPz4oMe
RQS/Fm+k533+/KzAJhc5wYAZsJmTWxweVvhohyhFcf5XsvMbVEHEd0S5VP1dtuvobWwjE1ZWA8RZ
Hri60TKMQo/fLSVX/3RpOSTC2B1aHWci+DbhybjFSjcmaosHI2awLEBbVEcRpYYmez0/e86/iD2C
rZ/d63TJg6fFEGLAWoRLUBI1jNLkxyOAyAJrp0Qp3VhGMbwdeaWEkKJtslVUmZyIY7Y1gukU2rz4
gyfZ4eFXthARO2oZB4dKbT8gL8DRbN002Jsy6kAL4JMM/Mk78QoZdNqhwxIMqiBouxlmNZE/d1zs
XkgVWFtPLmidImXTAxY726LCmnnUahQr4JZiwYqgASjLzhbLO59GYXXzKq4xY5tIsQYkUzw0gmcg
exNbNGV5mu6RGD5pD4o1Gv4v7jkmTWZdmZgf5EzO5mEib30kDwdxTD285S8DD2y2mIQBcu1nynPX
pmyGybBFhRuWGzmqn8WrteVKVCUG9B9C4UGV4YhuHd1NnHEtjLm6CPLZiPb3PlIEVecGHUBeS5Iq
hSu6wlD20WIgBv2TceyS/l7Pgbhqz9CWUScNY3/M3KqlEJ3Gyuq/8sgKEsoNjQpelS+NOsO0iMdC
6r3Ag41eYugmQfs8JZpWwWSoXxfySijYXYIM6iMyZ8p9gVqK1/KwBtSERtunIcBplQKTlh1gdZf/
JWy/6DNHGuiNuLBCAeUaH+x67UA6fPqOs/AON/XN53NN9uztJnCkCBXzS8RYIxS9yA50L6dEQ2Dd
ZVKMG+oGhlTbqtq4QTEQG1ZbFGOkqALPuIwBHiFWMp0BaP2zLxfhbucN2CnN6BV0PwLxUOR9nsVl
BNUGrFvJlWNu4pLO8wsbxdbboYQWceDyHQwf+LgDQy73NaoelFOtLlpmTFNh+a68/KXNj1vOqF8S
8GWVlyp7+g/hnu3/5LryFbyC/82Kz0gn323q0EM3QCOfk1vQRz5Bm2/Crwqiph/xFsf96HlvDOcs
ZN0KHSvGJzRQCNvpJTJ2U4UQYY+sCag3iOoA427Y897B+MpttOWoYmLd4oAdq6hKgHb4ZUjw2qGb
pQfZnDf3CTNaG63N/A==
`protect end_protected
