��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i��͌c�iv����'ό1_��A�����G���H��8���ř��wJ�S��U���A�,�{��k��2�Og�L�@�_=�s�d8�7?:�&�ȁ�꧕��׉�F�d���	\�J	�q/|U��Kt�'���%l)���~��M�	4��ٗ����ɸK���g˟h;&ύd��G�BĕK���	c��*��#sh|���
�@u�\quy�o�mwC�5�9�˖>9��F�~���oI��r?3�:ő�f���Ș��"�}W�w���'�,]�k��ҽp�� �<�;kX��s`���[�ؙ�J�l H1S���|�ooKǷd Iʲ.+���ϤG0J��^V|@i�g/h,
-������*\�2U���(9(2)E�/g�$�g�`7�5����:lֆr6
Y~@�RD�(�A-�ߺ��j�vftr��T8�Ő���vN}� +w2��?�@ů����I�!�K�`�4��ϩ6�R@~3�(���G�j
�Q?���/�Co�_c�Sc�zlT�B^P�Ba�2!f�S�ʷ8
��zM@ �I��ڐ�+���'��7�?���>�`��&(Na�}#N�k2��N��x��3۾�����Ŷ�P�����˻D��:B�D���eQYK�#YANo�{]ᄝ|��;T��_���؈�O�q�2��ߤ���U����ɫJ&S�#�/�
/�7+$���EIȥ�_PSg%
�r@����2��;g�&HO�x��0E�_��F�z�S��~k�/WI��w�7���`~n�M����O�I
����<�䓸��e�1X��RL�߳��;�~��4��O��ŗ��qJ��=���,}�{&ppk&�N�In�	�S��nW��	+�M��Zx��O�~RԶ^˭�_�'h������DA��4s����a2v�ů�W|�}H�S�Z��]X)O6�*ճ��.5	d��FU7M�)�&󮫚u�S����y�-#ʻs�&���'_v�h�Ulwh��֯�Й��6�kxT���!O�q+]M�xo�k�T�!f�N��6uF��/�|�]��O��ž�$t���ttnm��#��+��sAc���&o��^�R˪�PX��0����ć�NEdP&�φ����F㸍��*ǀ�q���:�8�E��6��b��:&��ӷ���o�d�ၿVq�h��w�	o'���x �����1"�@n�Cl������hQ?�ēJ��E���g�Y���}A���$P���$�{׆Mv�+�Σ�{1��b38�\9;J�9֪�*��:#w]:���_N'}Hy������?��Xt��ǀ�d���;�׆ˤ$l�6�K�:у�4	�k������g5�Y��١���0Ο,��Ed3:��� �5��y�q��+��T	- �T?D���b���qv�`�l��k�U�L#4�T�w����ҿ�>騦Q��Ï��2w��5����ϒ�	Q�c-����!�y�u	L����\�LɋS̀U�H���3D���b�Pv"�S��,% �4�~M�Î8�ć=�t�P����B�ZN
��Z�8��X��x�
��8�q�4�'�(%0�#�	��Ui%,�4A$�ٰ}��lj�H�4m����9h�&���JauRi��X̌�2�ρ��	�2"�@�T\�zn:?xQ���e�~����E���\���l�H_qm�9�oO��1�M�a��:jF�^���t��)4��&�H9� �V�E/�˄^�转���R�)V��v�7�v����ʞ}fs��8~D���R��AܮN��&��@LT�h"�/��_�;ac'K;e�:��_�M��KT��� �C��ɾ1�0<�?^	3vD��Ml:>&KE%�_tLjg�n�a��&����F�5��öu|�㑥Emq\������9�d������	�'��?��O2<ʂ]���{̤��::�k��Y��y�o����d�8���
5��H��x2Y�RLR�5��ϐ ���	��}Ҽ*���چ Y�~0~����
Ac�!�_\X1[�z�	Np3���W�E��EFQ�T�����,��M�Qm�U�����Aˤ���	
�u�T�2�Ⱦk^1�R�Z���V��o��p4�**~fo��~&�m�kI�_p����ɵ5ې�ǻe��q���Y �V��D���U��_���2�$F=��U���]�� �=�q�o1�n�B�7����GW�~oP�O(+ �Km����f��Q�]�^�[���a|�$ǥ��A}�gH���cJ�oq�s�ܕ�ܴ{��~�"�L��)��A� �Y�	���ҋ�9�*�0�Ɇc\�����-�kc���~
���$~���O��$� ��Fq,n�-K*�	ɾ�|0b ���_+�e����S�u��R֣��W,��uG:|���c~�k��m�P�S���;�/9��2���M�~�6r��g�*A���R�)�d �,�Į�l��.r0'rv?#�63��>�p!�e{돍GI&H����H���?K�<�/�ܝaゔ�]���ҙ��(�M�X� �z��ocs���fxAТ��I��������;�pJ�/ΕNe�aC�H�t�t'���z����\�y�`Y�Oz�D�#�\���L�4��ʴ3F(�V�V6�p�N�4"�p�p/�b(��lJ�GK{�ng�z�n�~�Ge��o��,�_�X�6���ֹ6hF� ���Kz�����f�fηc2�4���,�tZ����d�ֿ�$8�l��68�Y�V�eu4���L��0(��Zσo(�*��;�E�B}�Z�S��wH�;��f,�=u�
�6��65r���>���).Z�L>�p{��	"�i@|�]���ٍt3Q��'FJUxxap_�S��[�aB5p���ʝ 3bc�A��
��gX#�s�%��ҝu����[L
z�Ms��2¯#��rM�EW� �ȟ��,n�L��'�jpQ<%4�D���Y�"q�s ����6�jJ�G��j�����#`C��E�2�wZ�Ll����j'�n������Yt^
jI_A9i���n���m|���b��h��I�I�B�����\�߁�qܒ�{�?~gIҹ>��uO�V�s�@��p8С���ɽ�o=���(6A![�Sg���Ȍx0�1�♮ذZ��<�#��T�t�Է�5��vl�c'm�;����ۉ�ꂇVrK���'?�w����UYU��j̹<Z�����Ƴ�Lj�_|�Ez�R)'��^��oV��c�'�f�b(å�o0����!��뼭l��)��)��;j1^�Zd�;o�*�+&ٔ���6�?����$M�<)7�̿֟f���岔�6Z�8t�w��@�3Ą<8�u ��<`��%FY��DÎ;�f�(S-$$w��{p8�+��1$��Wq!��G���[޳S& ��[L%`�E��W4 ���1��Jxʉ�u���0����`T��׫��RA0L�an��C�zk�(���i6�C*XK����
����-��8�˝J	!�<jܧ�g�־��Ǖk"�:ʆs�N��z⭤�՟�3 �F�������p��WS�<�F��uhF��W���7w|��7����h�ʩ�S����ł��[�34}$6L�Qɉ�o��F�n�<��6Ha�pt�m�����ʋA;
RG�i���73�Ȱ`�zV�ȱiYP׃]L����л`���7[�S:�L��/���K���$5�[��m>��&�S�xѝ� �mni>s��� ����`��� �c��+K�ɦ�!�V[;�(𞯱	޹��ukqV�$/�#ذw�fħ�*����s�����2}J&�P���B�_�`�)��tI���W��=��=�z�mo�]��hg�j@z�!�3���O����O��=���$��j�h儸ZN��M�@U�FY�Q����I���W�Yd��	�l�M{c3٨|�������*�&`�p��g�辏��F�R��+�-_l�j��۞^��OkWg��G~�69�Y�H*���UR��hb~U�J��MYP���	Y�S��1޿��C���R!j���r0mٝF𐙢Vh�x��	&������:�? rg.�K�O�	�K�ٱ��lf��7�x������'YJ���9����G��W!)�ŹӎA5��ث��%�U��=���\Щ1Yg`cP���I���(+5��DE��X%i����_2eV�-A=�e�Q���ۃ�b\�����-4i����XZ ���kAMg�5�d�沰��캄i-���?:�7�ȟ'=[��vi��!2��n*�87Q ��5FD�ǝG�iRhsH�nĸ�f�t`I�QgM#t�dd~��Ŕ:���η�P���&�YJ�	-|Ǔ�i���!�"�	˾�X�v�:*�91��s�9�zA�V�J�o��q�����������L��o����*Dxz;�!�|��}�`$?U�)ުS�6g���.·)�k����`���~1���E��+k#��)Q�V�5>޸��i�L<��������ta�;}��~�Þ1C6dU9Q~g��[E?���O"	].ʖƢؑ&��� �R��g=G�D�\o>i e��yUݸv��-�,M��f�A�'���ώ
	�9�?.e?\	�a%�������S��f,�+��{HbWiq��2p�z�,Z�y�N���>u	 ew���dwU�X��t��o��>F��L����:�{>�e$��N�7ͱ���R�N�1��@��������Z����a)����k�mq��0�6!Њ���H	E�<��1pi�0��6���&��S�{�(�!��Nι�@�>�?�U�j���2�=]z/��>%��u�!i�D�/u/E�~��rcbWWbخk3��)��U�	6w(K~i��r�Z��F�h�QQ�txE��J�5���'Yx ��m�'6��Lu�\�[`���o+����KTm��S����&��(��� =�lESĜg�܅�:�]�W_Jr�܀O v �����"!��z���7jXZ�� ݇��̝-4@l�`�&�:�����D�������]�?1(����̧��nE<�}E�GP�Ԯ:.tÑ��Hr�{k���m#�س+�&�݋$�3(�h d�'�U�Ýڬ0"~ӂQ��]Nt���vk��V��!��8Ú��Za�Q�p,�w�8-Mֻߚ�u�����֢�x�ǌ"ї5%�:����ǔx�