-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SeYi/kHWCHaBogdXChpTcDKwlQb6icoetEkl4QzwX+orsVtn+xGlHY806Qu0HMYey9E1EOrsX+tk
AlY5ogFYxisqg3eQ3fwj10HnXbtRG+pTP8fBdESj8QqiIXXrpbisEAzvN72d025lfQ41nl/gkPRn
uCKevfvqJxID3oiskXhfiYb+rnQ3Ec4ZsFiYG05aKrcvFwC93k/zCp4T4wAPrgh3ipp5dq6XBmz5
dNjDVpwpo655gPG77f7PHNpVXHpCCmQ/4AbP/PfcoyltRTtgtuGWf6CqKC2vK9cPfMAgSDqrHNkd
YR20T3ZPPX0M8X1cc9tGmZ98XgSAmDRsN1ANsQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30288)
`protect data_block
v7UxEqKLNNo5NYh9rg3iChVpnWaEJtyKCqG6sqXx8Ma3vFNaPgxQWvq8VLZkwEPgjuoOXAC70Koy
V6vxAcsLq1dcj107x3gEfBCcOkqIZoOXeqnOyWRxw4TGckEx3Y5ZdHmQVVxR/V7lmCGfHbnabvWG
WBoHbbooxvu8eqeM4nEJA0vW4rkeItwEIcOzkbuYlZyMxHfXL6FjfDm6SV4PnI7q+1ttGJo/nPLO
ouf1QlmZvtJP+o5f2orvUD1X0DROqUdcKwclYPXxLLrvTrAjXG78Lazj38f6LDXlkX+8vNWz63ux
N9q50kjyO2p+9CQ4TvejxDZkJluOydPorn7al7tiF0VF+u6V8PHN6bpmH05Oc5pkRiWqH7XnR+ja
MB15ABCfycoaLUlsI/UmP82Yw0YjRNl8+pFjxmxrkI7rszZEkbMsYIEgqxHePh3Z7/Ny4mzvGFr+
YRdL0BwOtdzb3nfN5ObwXouCz7YG02zTYgAMiQyGpm4s7emdkngQYlGF7BI3UVBV9rJZCE6hKrT6
U/hVqUKvWu21q7Q+Nscn35mDa7be7VnPRK7HYm9wQUQUQQv6I895FpOHS5Z6vYaB7hbM0aNW36Ox
9VNHATJvf2bNFTdCniYs/jk/SetKXTA7icijpSBexKHWhuWlLdrYlClzSMdvNHHl3zP9iQlf0dF+
96/3E2sX34ocjto3ecbJ24J4U7SogzK4/4sK3lMhFznUhdlH/CCkYy++A+0o3j3/4bnkz9TNt/CC
xF2jPsvTb4vN3NpkARFTemvIl56JQl4Yw10+mTunMRy8V+plMYlbdEK0vLIOSOLrQC5vTnldTQaD
OVLNMzXSelAfYY9/8VJlF2BNzbLejRjpZj35kubIqdUEY9Ajrxt/iyF6YxIzv+44rFm/ufsKbemj
am2W+WKdZ9iTc9hxR5ffy/Gd7t2XvMIze8l5cTkWScdy1aZpI3CBYOYyXxGXkoVNxGzsotOvlQyc
1E/98qNoLn0KGRpsO9MS5psJBuAmg2hPifFTjaJir+G+SjGl82b2j3JcFcr3zU06Y75SJl8raZgp
Swag+69p5axIlOaMWKNWe3HIjpLTOQIv0qWxnxvCVXOFMMhZrAL25ojXz3CkA6wtg9k82wgdveDw
7C7Q844iJV2rNO8Q7RgdubLJQSLcmcZ3Rg5jwViIFgVvXzZVRFNc1rObfb9rj9ys5BCBqxyZhFrx
YPxXaC4j72/G2j9kFV99T+ChXiwIJPXvoHHbsciuQ5DyyJi7ocQne/qvEpkiavvRC3Yse1/GaxGC
D9pANqbDv8eBjsNWyPXztSaTYC+1a+LEhfTmOqxZVbjKzkhW48/hEebBAlgV3oWcRV4A8NFP4ap4
GkJGWlG/nu4DkonIIzDInQOqHHZnT60CYAPVSQ20vcHeLA8LTx/k7nGMgXh9WZ39PFE+UjvE/wYo
23nk85VCDb2zx0xfVV70AVr6/4G6w74MNQiIjAUuNIuYOuwp8bXJ1eWXyV+kvqfy5XJB3VHb56Us
O8FFGVN4psiA/dDpvkqHfhpIAJ1NwPhheafToWEhvsMan7Y7Xv3rF3Cj6t0HJyyClLUHEnk2MQik
K5aNxa5xOW2dAeajHnd/LYqAFLlaIuBkyKG7Szp1wGCQv8cVWlhPqUeQIe4K/yiDT7mEGuBHsx3U
542/HdK6GEd0XFajjhpZjF9Y4YUA+3gFkuQKsq+iM2YEZ6iq8Cs6klE5r2w0Td6KC6V4s8mtp3b4
vFqtUaAeD3CB3X+ktibx0vOVBRS0llUDka1SbJpM0A8klPafCqg41WtTCPcgSiteapiF618CGUuT
b09Ho5zHJR1inJdDOStZ2/DWpAWaoTktU412KzFaJvmEG+zt9dLLfcbfPnIWGcUY6I2A4gKh0CiI
iVEEzjmSx3MzWjKOcP1j3kamm60ZS1Zgg3sUAWr19D2QKlJQDQknDRKnkcR1BxkA1JvAlcmNsSGG
N17lGwYgFNUTmUOZ/VrnLSMQpUcnPXqO/MyWj3fv7cGV0D4P2oPJEnNVNUoVWXqcLnAZBzT+RTSi
5+4387XejLPKJ3jUg/rEefC+drSXlc51sDOBoPAJkDOOcHIuyBva0Nehylhi/a2vkT6uBhqgcqq+
cziaxrwmh1JJOSwhzEQX1xlE13O6Txrthi3QHuLQOYb8Pq2w5xF1oB/pduW0oTzaOiTMixw0xsSZ
knSH7Gim+lHzn/7yQ+9Rsa2WEuTp7L4Nwy8spBml3LwnEdX556oT01ke8dj7lO7NQqDku7lndALd
AncfKUT2O2LqzykJiubkbOX7tYzW0LzQYeKOSjribcPZLodyDg16spbci79oW4C8aXylHBsAWgzu
+y4Z1LBreVa9DhalkjQVbQADFcAUsDy52HAej229JGVEIKUdJH5gUh0PAH3jO3t/fu5BfH3l9mY3
INFIS1RkOerxDp9Hhv6qG0RxkSl5M3v4nAsJGjK3lhZUkhCy/vkmNeDOyKNYs1AehCl+I3ENW5wm
octM4OwCeSOIrxZt/HPa26vVtW6LsYFogEey+p1gnRVvoTakwryIhXg6lx2o5Y0UeA2fY+KnzSeZ
WcJNlI5Y72lQqAGm+MQJ/VMD3zETYcrK+QH5lCSO/RWaxnSWyuKey0iBmuH/dC4Hgh2SBSFs3mRh
oeETE06Zv3gpJGMja1YQd40/3LP8BOGtn1JmRnkfmRoFJwDz+wnZ2P7l6cfhWqAUa7BsGGp7ckXl
OBVk/XQ7owqutNjehUmDbNWP85cRlh8eFX/AT5Pf4Hz7maeqirgIl4Pd1/Sp8wLs/SlbYOvCLTG0
ciuULR2d5tRlkLgklX88ZGmY6ggDcHnAbpf58t17cBOs4zrOAed9MtOVBRbsAEEkjm55IjaJAvDu
vIsYPD3UNe3SvUn4t6rE9IUuQVXQZEA1LKb2T8SlgUbthuW5D5CUWABV+k2R3q+vd5sGAz5k95Hx
r4hTR6bP4WBh1FxNGJxopYjE9zqYGaeTksdFRYkIZmhsdozIAyAmTXROIy8Nkm8MNFO7Z7u/92r9
5Lv76gdqBYVqyO3kWK3RZTmR/U+ZGH2aE319hPz2XAi1+Q9SX3cmSEitONO67M97ipJLTEONrv++
zZLNC3bD9ynHtf+wcQ8CCitUWdJ9WoT762qXa0veQaTjAb3BtWdoAAbqTPp4kzNcRHP+K4KwveLL
xm6GiFW70EfAd7YHlcxEB6LrswE54KPscOf44CcK1IkMMl06W63PW579bSSEGSzf/XwefNC4UrOr
EN/T48UDfqKEUedleNkfoEOndy1T6UAP5Y668VE5maEtvTNgOKNQoOGmoGxyFQMpe2JcxeKJzN+9
/qqrmT0oUV+AiQFC2YJ+/IMyJTts3dD3SGxeTBW8F5O5v4weL1QWX90NfrIUKX/x5NMNq90sSQqX
SlMHjCcI1RoIY5VnSkLaJtwDRi7nXgdUkPHcNJamsCe1F1Q5WEtxq7g7CA6hSTlaRfA+QAPYsiok
7TPFPdR6ZuAyn77TUZxZbVOyuUq2DIuy8KxVvSQ+Nk0KWHkCTQrfVa3P2SkzsgYoFo80TsmGcr8c
pMdl7giRGf/zmzMgWvQENO6T8h074VESPSg5zK4tvJmGBtiFEBMa5qvkePb7511CMUnPqvDOnSjW
X9BJIadcAW6M/9WVXHjaRu6d2VI1oJWbTMHCEiyr2Rl3dJLxyOJMl8muaBOrTmlf8RLqQJF9w3Gm
Ksojl18yc91BZoxVQg8qV6jXtTSsZ+sHjS/ytNQ2/ok2EYsRElXA6B3QKSWEfekt3k7EUxjapiS0
xvTjeSCdFxpEMBCkyxQycpj0gmSL2jtn/Gqk+KKOFHfBl+JbLFIH6UKmD6JRuIxrWOrACok7Vnl1
mpzW8IINeJthR8bgiailInAbpkLIpZrdrlDmH9HGwaMzf6fwZbRH4o/zq3trqgosfBGTOVevo+rg
Y2XhWVD9Z1lxzkXU4ceJKJmbln7YtRqpW9qQAy470FDSMawj7w1a8jtahOlUR5REW1qMhDj3F7u7
v5SfHJ6PmghyCEL5a6NN1BCeiUsRDd+GceFFrpBdOhL0a/CcwYZ5VciGzojSfnCoX+KtKajvJn/G
GbR+Bm5DYp5qTzVz8tHnh4HcubfSSkXBLJvgy9Ukdyf/2+stLdZs/hP9BnHmc+GSg8zcOqsIaP8S
41ND6muZ6RK6A6f/2cFnhXA8P9Oo0aDcuNo4yHkUxf/X3LhM45KtginE+sAdQ6G+1Dmk0watlqYR
gzcm44kx5viSGGpprwX5oTZWmW7vvRMvdQrfo68xMSCQQ6PRnW0A/yRPFxHNU8kRPMUMuTO64UCc
JZ5mXS0vUwvurGh5eM6xA8TuGnqrZys5exE4QeSSZt1VunFA0fpkOlFLjFQYOJ4SnKQBgJMANpyW
+yMghCGAVxXtvDoTmMwyNZ3wf6MH+52+AfyH4O89rVipzdokAqudbMYcTK4ID0lfeDBZsO1cgxYa
/Ph3rpIPP3eeqr0LL/eHdZDKf3yCTRPgUE+d9EDUZmRX+5bvZCKL1ak8/f0Izc9sSxjU4APg9XsJ
+ZPrK5WmocqdDpXVet+YTraxM6MlhIvtn6mFkeWKxbtz6d7IR3yRPCzzLQLNJ9NCsi6BE6pG3n76
ESmvXagTw8vAVGgIg8XUk/WEucJVbSINRoREOFWCpXbBakTselSQ9NHxYu5jAlD4UmZ2Z3VoGtQI
lYvp+H+qMbW3YaZ9LcB6vBZK2O0hdFaCYz3NGaHBhDkm9Co3dLNI6ZeoXzDfQWN6DtfxEnY0vGev
WOcKYpd3MZU7vzRZgf4bj4BlPZBC9x/yH8R8nBGa9o/fB9SwfIj/IaVNwsm/BDsuLE5zGLOj3Uar
Mln772EAZBDX6ihcKiFR9XczwlXoMdAL2SUd4oItus8aAOGWYP4BP2IVf+HQfv/gIUZ87bgGYJkB
szWWjQhcCwEoECnYnkcTswJcuJ/G6mM5S88h3Iyi1ACWK9d9lRTgvVPN1OMxdTG9hQQJQ7zQns7b
IlJfDiPzF0sv6BNna8tDFjeslofjTaHznHZkb4LmrIp1P+Srq7Gn/xMThRgiJmKS7a9CQ+19eHDq
ogMiDd4E93/WVt0iXtt52LOvQxOMX1u4sjtywS+fG/L9s5Uf+IQQ5BmRdpoZGYu5h763Z+RklB83
5RJBK8MSj+ElZNe+uLOyMVd9AvsWoqRgEtYr/uJbkX74cxaXy79DPSn96OlreitvWMzXNPLhcF7F
U8hR7w1SZQlrk9rfuiLAM9zE3RvEUWvzWhyqBdmMPtQmjfD4Jth/Gwo1I/PsH8Tgf74RXWMebc3k
Fw6tLIMEhN/OGlUNkCGgaCEVlDTm+4SShPR72XonQhU4e/DztSNlcdASUIo3sjI/ThpnneywcTVA
X+s5F0ZfdqyR3rOhSwH7J7ow2h5jPW66T6QkI1grtRGZw469Jfww6GpTco5k6WpG+YG/DheS4C/a
C647tE2DYC9AYm9wmUcDiyAwH7zCtictTReACNV2I8kZyL/7I9PM1ldLbKGHYtn8zKYOoxwAU9dq
EBrTrPzvWrmAKAlaXo0+y4u/u/RI/TMmNtXdARIPnN7VaSv3yl342PBTKHDGJaWVuEDsj4fz4Qu+
leseaavnkolCtalP1mmWBvwaYgHmeObrAKkpe4vHEPDBoIOpG+HLmFex49JCS7oWv0tH+pR4b+Y2
mRQdyco7qB0aOi8vjT2TM4MKG3LO8VutWharXAh4szjhCIuSQkd2/Q9QnIIV3tMT7HRx/zuRqAqY
KH2G/GpnRtUdtwRUEBQ88X6J7ZBxxUqzIO0NBeVg6PpflCg7ACVuN31cnxl0jcXgwR7/Qe0ZZMUz
fbCQ8RMFcTx8SXK53g1SfSpQoF5QW0NpCiVYKwUwCFOAZfsrOW7FC5ygnhOk0wD5whHbVtJBcGyN
5w29bXMiYLuE1eqWp6gDgqplDNREqIS7F5bMI7UkMXyuMxylHJh2h1I49dL4ZpRHQmBDnnMLNOlL
oK20IIKHhWSg6CHNaCpWYhdzvxAostDKlBwgMnnIpnXC1JH+Mr87ou0OIre8L7OUbYi4++RUk6W0
e0MT8moVIeXMzieQiFyONc9sH2wTgegoxeyXHpcCAiPSOoRCT/w1jakO3PgvX8yT3mB2Lbnf6YMZ
7gUyORBKWfFKRu6bR4h78s3Umft34hLAeQqOsblN5OUokw8Pz39rZpLvt3wy2s5T0f+8ImcMEKSN
lU2l0hwRfNh9fMtDX3YnpteDeWgPt5FqWhpYn6g745qodXMJ6844I4WVQODFGZttdOXMgYGq9lTd
PBVSeUEkZ8Cn4TX8OEG6DWB1LVQtkUuG4BVp9/3zj2wPKhgsKiqIbICOzp93XWXCMIqAJ5zAsf6Y
SPwcRIpycJH2b9eP1gvh0KjPgkPGHzwVe/YbeCsWS8R+sfksnVpuYYODtKcShJkxaHlUE+4GhI/P
PTjULULUNm4IbNtEgwzAhBlSJwkIo5ndoYHyEVIEPBVAnF8MaGSrZdZV6Myj8udCPVmzriqCzT2c
G3MqDsY9KKLItJkoCIdv6/S32xFIgCvBjDb9Z4vRrIUJbKc0fH6i8632Tov6vfIbJIKl2SWhSai+
CmmqmcL4L3iEWTkkgut/8dRYGJr3Ww7FdsVTuCVqplQjdVgc+vzd7kNmqWYIbBTzmbfKd/YcYb57
0ImcibTzWB20rePROE3wVyNZ/S6UM1ZRr3bPWMgonewKcCzRVCEDZ/bq9xW82bq/6bA8JsAc0iXQ
JChTYPD0/t3wE9zLUTmm9t6ZucZG7qan2MOFmXn7UlRZfrY7unvfvgrysJkT0ABkL0gpoKWJ9RtO
cJYRuQFbCqwrQhJH2+dyWINY5rj21KOcEf1+2uzBVZ4yUAkKSGbg4XEeCHgjdV3cti00XvYRsqan
QFkNjjUbc01PSnYEtSZyoUwwSl4VAt5JPtOYzZeHf4qTlObCWAZmJm2fnhU8d5MPLNMcshaMevy7
UOv/0sdXqifrMbDAS0kWrz7a8wsuSrfgktmOpUzikykRdgVnDJ2ZxfbL7Dh3/smr62QoVdZdZlo7
WuEUwLgbLklZCqi7MyEQr31WAy/hyzmX5KRC7Voro+XjQFWiGAUNkOi4UIUVq4OQrOwUPO2295X0
DV6foyNztMrC5Qi6Cxk9EK4Z21u6TTi7DhOe7hPbBKJQkrwrItrRmAHSnsjo3F1NElBvsBHlRhV9
QS+aHfNNWMIVv4HgQ4DOV6NV7HX4YRDkz1hH9zclxig7GseNcYSbAf7esYOe3yW0NncDUy6Kskx5
h52qokDcMF9jjft4IQDMJOy5x5fl5tz47nKAdEGESi/03xVuMJSw62X6YzvqOPD67kWKY8V8WNGu
5eYNG/+nXR6Xzs0cZ274XefyB836Gf5pW+auJOaObQCU4fkA++/Y0e2fbGBXQHL46aSB/mlDrUa8
MSYmclqyZvXxbaJQK5neXFtezMQHfhObciOBWrsWSb/7x+VjVIV0FcFubROYcdcWEzQGXfeNMcr5
djpkRujDWoQ4HnsJbpmCGZc070e0s01yM1fYLKIGug5c5KhYl9Htgj4NtmMQxYUsly1vaXcWo/95
2zqvqDqQI2SoGRWJoACO4I8QyhhzEP82+ZrF4L0EY5vYr3VntHZWD3QO1WuoKYS+Bf3DwlZrAhF9
UzFy4OZXUCDt/65/k/iONgEyh5Nj1BRr91JSVtaRcAuqFJZPEXFZX9yhVW3DYQzzs0Dg5dMp8sbS
PhjTChVsNJg/yTIf0huXNuDRA0WONtUYHbv6wmUqeE7GlodQP4Ddt2D0wP4NQwbywsLNhBPVwbPo
CzeSXA9+NgitOclMPYGDmA5PGCSITRLMbUqi9BdAVSqrl8Sb/OorUTlkq6vXyp1JwKA7z0zMlrs+
iONyFbhJ6+s6T4h+eOKn0+BQPddSnNlwR2Vkf84ieumtZ/qLNuelWlOc6i0g6RAiR31CRfAcpY8g
oDDpiYevOsRXpsG/dCMPGbS6VNujT60tdolXE0qv0z17q/o6luk8PqlBqA042iSaZO6pmUWaLWix
v8maAwWJnYoVsfKfT+wNfbGF2UFDiKhdBXVcuiBpkCPbpH61k+XU/jdFe2qCVbxzwl3G3kbCA7qs
nHvNsTHf7fQ+d+ClQVIDR3eTVnjDHpwwcKLYZg1gKUWUYsV9lmht+JDudZ3cOw1kCAu4y1aOiOym
I7z7IwLVC1h3AkNxGtxd5dMvzNrp0SQEn/2SJ4bjQnmgFaQKPUtlT7D+6g1HKyvI+EH+uiwi8KXq
aGrzQzf31mzn7TBR9+nnfp1e57cBkNUnVwsxqdZWyvh7b2quFJj98GUm1w70BSFF6ts7Yxobt7S4
FDAYtv2fX6V1BJSInsPsY9nB6rEPjTDLbV/9zA6KK7Wk+P64V1cMU512r7oG0Dh3QwQJcQ9HJWHu
Ck23hMT/46ZKHLNDaNQf5qeYdPZVB4MW6yRD7gs0n+ReuSx2LliKWvSNxon5JX12SD+6Xq033ftw
YCW5H6TQkFFn86r+eZ8QvcsYjT2fEnNTWL06E4/MxiK/vMETQdBj09Ub8vYRcJpTM1tRqHyIU59Q
A41wG3vfdeF4pb88cWJBBU1E4wWjB1PeV3iPYaFJMTZZLDgkMddIchK1/FIUeTwxR1vN/Frg+MFs
DTzZy2speKYpByiyYP9pDOzaDaQAaZ3mHepqj7ENjTFk8Q8qobObIVHghTLuhWrWfq73oK+OeUe5
RZD7WQeQXDz1sqNji8SNPSwp+l6dj3/3GTFBNSqM1RZ5Gf9TW1ykzuDpS5AbD1cp+tPC7nBorI7y
Pd6qXdn85VzI25T7Uyhyf+R/wQcLzNotX16ppC2Gkq3W8CHGi/YURHFQG7b4xgjn4+OSA3MiAfsU
EOD0RiIF+V2KsL6PQx1OX7pEseLejxwtJJoShn1afPH//m61s5jIubcxXXxPOyIVsoKWVZxI8S7t
nF5qaTaz2f8V5n2OhVP8KWAB/NJ1prqPz3rCySCXQKwlkF/b11RT8haBq0RUSQXcUGsMXXJCRr/g
yQR4pE1VaacmtfekWQqHRkoh3WmPRhGCpax8FmZSWwc/W2Qtedkmrf7Bs3VfRSq/rw6k3ccFuMzT
uw5IXytoZgfP4ykq8UzEUwOPMQhhuYWCZ147kY3mdVietmP/BDcxbIGX+ldEVYwOkb0yG7Pa5kCg
/twJ/WEi/MGnjywnxmGehRHZKxdzyd886O+/+62Xx1o8pJbnLgEJTKh2uCwWPr+HTP1wiY9RlAv9
/cEfQ1tYoPXoSsgpqq7pbo8Kv6R/KO/LVY1XjSEhjUhFxphzmS9Wbt4intg8eB1Xtk4igB2UfEVo
Uua9LA/Os7T0c0+0WHlMyH/BOI6nYBKOt7p3MDU+emKAuIbZua6PamcExiqmZUoeGI0NbMEa1/Ov
zRD3CcV85jmgLGJ8AZl9FtR3etMFKPGnnK5Mxocsv5lUCN/xFmKAjG5OKwe3bAlu5XaYmp8Yexc4
FNk+iOUAoxXNQVFcqVKypslH7LDDqPhG8uOVKjvdggD+MSxrrqaRCVAi5wJn4clY5/5pGq9rqliZ
M9QXFpLHkZuy1MQDS/9v7ZaCTWNrYf6i7RtCDReemdNCeCjPIvu/dhNcx+30CwUM0dTyHeEdIgdg
DvcAFK1xcojQFK/AhhZd7r56dJslj7qgAdUz3ZGjpsT6kBzCHbnhYoxJhbDcMhDgk+nn+xwzloae
xLJOqMww5e799dJPmY8avLfYd+DlVZsn+WXvlFBftEq8UXHZMWABrfb7xYZfLiW4ZD752yoemxT8
dnIXficTyEHfLvhgLHsRS/0OPLi2hbL8wRP0gJXnjlshZ647rz/lvsH12XAIXddGpddcnYZMD3Jc
ITW68jlMgcwknpN241IK1PTpfCM9jVLTn7onTbL22tQkkjs5b3BmjDsCAI1TU7z0nDVzGqKCl0+S
TvNHa4oIl44SjlAEFcy/jge+L2puuyrvoeL2VLPPFp0PITrYccTUFpYBMF+B1hR6ilvqh7+AVy7U
JVZZOyxB8D3+oZ7Cfrb14XWCtGK1DGC/mrslWu5Kg7GUzYUQxiF+DcZgaRdO6MG9DkMjtB9lZHGz
P94rlddRiGkJLAX1kgRC+iXkEjWzStbZgK8IGjZLHwvSgb3oe2Qu8508JJBheNv+Q8oWmGn4jNMp
n3Ixaup6Ox6N9uOLU060YvxeacXfbC88SZp9qikZ4+i1P9anhGirq8JyEjWrTm89dC3rJLjYmAZ0
bmqWgadN3CHVbhABjkGUZ06RiECgEh/282AMCGVsBVo3sFanPgFZV0D4OKagsqSc+Yz8/nHht4Zf
kjwYQoI3BmlMt7XiahpYw3V4kXBSsaysz8Dg2s4mRlaPBasq5WErdWyVhMc2k4bsgTLumZjIxsfa
Y3EynaEwMHxaLu35nulJT1l5aMIoc83l+FBTHqWD2aATJk9eY/Zm37D4y2CVVe8Cn/T0f8TUxvG6
3wGtV601ZHcKsZXtXP577c4ix5gKTWkIcRLfDs/pspW97AfQnOj0LZN33BabRZ0eQTd5V1j0NUzd
uGXxpr1hntyK2kZxNxUlPmWbz3M5WrqW3ijKXvaGdvAUWW2/TppmPUMOxnO6JybdCLaCLADVZHUp
bDe0z6D2yIfKNBNwhHgKCyvNzhYnZHQa39q3zUv9eFsd+c9SDorxycTwIAMpGXEQYz4ybV9scrcb
V2rZgwd2dcrjPkKiYLysEqQVeiVVkCrUtxedSP5wZKRHAfPpfaTfopeVvEInlqs2J7n1MXSf+nIV
sF+yI7FqtUIa0bfmYHyINUddn9MwnhXz4O5vl9ZTXHcW6AHFRCIf+4kTK90Bt7yeYO3QvYNKtLOd
JoKOhT9FqM2gfZujBZb+SxOL6cTwFQl+i0hKq51+BbdB6gTd6E3EdT066EeU6qDFZYQHjqWVNov6
waIJP2VxINzjpg7X/yctEeRwh/8NU2o61v88L/8Svc1pCOMT0F7pTNUOQ9LANlPwhnME7l/ZpOVQ
Cq9soNXwEU4c7YelpimUhy/zZhqW4LiFnEKKxYxYRNVyOC8qJzunzGRD/euq5/ezruc21fKhhUbi
m9g36dSo1tLiweNJezROsaDAU/kbHxjaPvSENFxPKfnVht5/DNm9rDKlwMRGWGUSwzjyRHM7Wt8p
4fC4jDOnDrqu3VXMwkUNDk16MHYUg395J5Il0gT9qqGQNxXVObCv9untkus7C6SvlPPlMUsrweF/
iXHUazPd9z4wBiUoPfV9kuBNFkZVKgdDfXfNs/3lW5USMO3MEC0X2jn/v0cCP/OVqLIlU1Uj3fbw
EzbmWBrEyAqtIS5Ueb2LWCimSQjBGjTbUiQ7x2G0Yyv2uJkqM9lb0tZFsDz39jclsHqjl41A94JX
XRGummrF5fssl0Vi6a/y8lE5J3BypYkDNI4ZjjL5uiP/Uq4erZhXAHFQ4tFbnPkDZbq2+r26jYaG
IsrtTRw97+ttaJFaA2NmovH5TtmmwnV0ROLRgI7UWGP/hV6WLJ6+nDQlaDPb+Qp/Pe066laTakOJ
qgNLkLuHX5/CJBRtQsCzLGkwbhK/8nIdYVfhXA9woMDqL2prNHveI/9Vbdt/6um6yMxe48t2080s
rMiRF/IpIgPvKUfQHMuEYx3eUF4FQ8/pmseeooM5SfoctjLTjlYz/M2MNSmg1/FZ7jw8ViJkaEAu
WdmA/2PJ9qdnZCOxSib4ANRxWKZvlNU2MuJKQ8c1GItwG6/zTVh+qi0x0iKrSB/nruNZvtPcMpia
9vffsYGucPU8sBTj/+ky5eAA7M13cIemZBOiN+FZlTt+uSDHhNz0siEtRVo7t9rVVaptLsWV2nN+
bTpVuHd4ht2gzTj72DgaUgkAdrFA6MQZBtU0Xqz8O/4Ev18LwZLVoQLhFe7gB201SVHdHaeL9GOz
NHD1pmLs7/jcwhFXS38zYJEM03HbUZUdC3GbOB2BAt61DqhAcOlTXSzbDdrbzPujVmLFTZkOPoYD
o6jXghFDN73dYihMwZLv9qPZBv1jwi4zWN0woi2SvZ5d678MX47nII/5D5iwz2k3KniBcqEqb1Mm
Ijnk7M52COaiet8RNuRI73N78wC/Qv2QowLYESfWd6Blx/dMQ0AUaLuOcN+TQLXk9uMbPuCV1mXG
XxbyqC7pBAn6JCKFXnCDtjhYi64hk8zHNv6vIjsf6emgAiaKhKJVGY7oj9CaKDHiehrmuovzCrBk
MQlPsYBlxLFAOQrFXLHpf5K7DSASZUNsezwvWnt0Rz2SxQYnXsKtLcSqhQ9O7OWmJL+MX+hgHoLD
FCoSOhQsg0AhWI4yhMFiRYHq62I3Ks1j6KffcLcBDdaH6aLrI3UBhClxNK/TqRAHW39+AJw/V8Ye
JjtfmVr5R9hVJEVlneBqjjUdXENGuvm46y+xbzy/rwJllhTWtErWNCz7UCfgBkqjcIK5vjVP9Hmm
fS2Q7zGiCb0ECKCy4p9fBY0JZUw7Z7ikmk0/jvaAZf0z2vPT5Xispab/eenfk6YzXoot1XQaWyop
xWdZkAR3V8TdIu1bPXIHxLBMBHMbEmXzk6XqMZrYb/IDXTVtf9ogGxRvE/aM5uhM3rEJ/h8HPtli
WuX/0MKJedmD5fnRaS7ukCXNYiHUcLv6HiK018+5L2uIuMC9ndydWj1yX0/EeC5QmFV0qDG6U1ff
V2BK6/+ybu9G1TJRuDDdokv/SGMI2GTfHpafnLWGrbh6S+VQK7LwDjxx41aHsuEzvHimOM+evaKK
NO/vEnQU28ahCfEYhpvRVW0YpTDHNlRy84w0MtFUyRWWKE/87wIbOPr7RgnRWgjHUrox8fwH3Vnc
8ITcEX7QMCKsR0k2UiYLbyfc61TVo/hM6VsPKUPnW1LfF+cJyHFDd/0AHJKRNWsmFnu7bPZpyExS
lyqZgD1IcWKAkhVBsMBreERMd4zpw6mM4EZCDuCdCLDf9RPnHjLhIQ6g5AfnuYVGP/Ixbn++1cpJ
9GD7TDRMtevMvR/lSJGj+r034mLKq2ujbAOUCfonSqhxu/ZEnODyxfDfTUTYbtVYc1+BuEhBECn8
3WyS083MQ1KWKpZG+IUXmz1OyzL8UHoDgqC+GtymL9XEE3SaLY/U4nbmQfayAEGZUvbwFQH6aDR3
/6oFsjxfA3ebzA21t0pPD3AHxdJEJ3uFavUk49+qfLTthAMBqrdB6ahy5lQjRUAQyXt3/0h4cDEi
69YG8UfjETZlBJtlZNJ1jPCPyNdTsLnju+JylnvL3GaqEohIUCKJYTSrLI32FUY+DH09GKbqtt9H
tE2i39f3Hq/l/+hA8tkHpJC1pxOMLOWQM7yFbvY1rd+RC2w4bX2tIKKRnt2p9wYa+wM4hBe6quLb
kbXdnpQo1SJUFW6FlafqI2oOdyGA6Y8fIchFI89Xy7HnH701pJ7PwCInC340y95CE9eq8+8IoZt9
qdz/DrTFKhSme4z5WKIC+Lj59B3qNoYswbsrc3rNnxtoPt7pFzVOSFeE3VxQE73tZP7h7TZ3UqRk
LaVWwPDYFDyQn/QP7J2kRoAoVULnMJw2JBSKpdrKmkeUAaySJIZ1/DUxElimg4Ads94eiXqbV4ix
b0WymZLCA6Bq84eYWpwv7PXIVD5cFrwvD4+HDfANYYfQoEaJb24DUQp+MoVtiZRK3n0wdyP6/kQa
2Lp3qVheZDovQyS4jZOwAzLLsWWjh+ZHAhJ8AB3tnTjVZmGgUjexPIYd6S3ExXh4ky8H8JlnKvzc
rFWckI8UHT2dDFV8qDIWjNlLLuqlZfvaztDCWlp5OPJA8GO3OSEKaFppaK8VR4rT3LA9OFY33Amd
tYCi0hCRrTI1VrM6eCGwwC9nXFoO4YZF5rYfwNjcWxzMPDgjUOpPGKbYzOtP3w7vnEWQKH+m7inF
qyDAg7cpOfwXY+Jia4CzxISYNGmw8LIpsGK7qSWFYM2raE6NtHKUZCuT//12oyl5GTfQJPysHb63
BpRqxc7emhQXJMollnNkKo19tDR1EbODxGLRi0MyNYDdfi5TYCIcn8sE53uTmV82zdU1sEnISN7V
DMcv/XC6rzhWopO49bjYtfhUftzpwjOTPB9+YHbY7aDPIyMOLwqaf14ejpGGLSib463aH2STmMrY
RgdSdMD42RVzbNummk5xcShukdoMV35PWwj5SXcq8HvQfrQNlg7PD5FEzjMJOsgY5GzI5bXjqH7q
euhwZTvjqLmImYFFzJXdQ0h1eBVgwIb40Mn3PhZdiZylYTtNFK/LT+a++7Efm1zIvlvjZIjHVmp9
6XSLW99c23vukx98vjzHBUmoVmFgTZvqKJTJJG8ubDZy04SKP3X9/5+UBa5b5jyfO2cLuSQIFFCR
i3A2vxHrisyZQpK030E6qPmmLs3TxqW5YluPITqO93/s4onIMFeSOYK56zslK+x1v3IvYVf+3WFW
estIrtxUBfLBn+zawjdqvgNMv6+Pn/xCF8Dh55FB1YuzKxVyIesoMK1tAWGrSXcasMErEOAkatxq
3Q1baR3URMVIRQsskRsYRq6ZwRnOdRjfVbZCY3XffRN8itEayx/0azjmu/L6VZGDEiLSAQEpApsa
w6wTZVe2+0v9YmfCVepSANSjR2/FFfLiY6Gfm2lDqC5NSkTaKN6rCacPOKTNcsjFvpkY4F7IcKXO
SBlw7UgUWem9f9AUacNHdTaIgZkSH/EKFxhBf1/wvRaNRBv79JbUUImcNByfmsZUU+3d72iY2V7i
PfeL8lTJ+voEXwwthlUpVJcm5xx0UAnSheTsY0vGWIgn46MXyQeu1YPzXX2bWlAZCCpZqMa2C5T9
yU4yleabDXhYvYpBijLEClHw4SgurDgMjICfapKb03wXOn+RGrFNTnB1X9VbZsuYB5hwZmILwHiS
h9rzzFrQwexgGA7sBEfP9WK46/q/cv2fpfVJ42BvbYmT63nO2k+q2uLeQ9c8Q/Vf+HPcrx9nPFrD
oYGiB6In81YZmXRFhwzJSsio+Kx656WFj4KrkxGFnBKEWaXXceY8G33fLN3ANvAEJE/8nhIG2ZbF
KYAQ7Z03Pk4Jvp3YEzFvZu2ClLM+D2GgsGy4lTXCAjrtFEROUbxu0e+9f+bei6Vz3AT5CyXb9g91
wqZe0OYb4CTHuBd0/ekUxq6rklnYyV1T3gTOC9nUh5/sN8JNEGlxO6h9Pg75bgOf6V3rZYwkHwIj
TaJ/9QQViloa6UuPPLGnv0u4hYmIcgCvDhIVRl9hUsNsQyxUaEzUcaXQaHgkTBg0qZ9uUtyj09OB
qrdyMM825Ec7YtxBjlO0Tb8x3h48C1dwjH/p1J7/3k3rKDvnefAQBDnqxrlZR38LfixU7LhS7bra
720pMEJZH/Xzw7I44zQkl8k/+d28Fnk4qj/E63mVIONl8UuFZPQ2rnk61OEyuov3BNJrXJ3JbaiR
SVAix69odNhS+3fT7cRJLG9sgejGNLP33kjdVu6xyGwiMClU8c1OcpmMXYilJfV4RHvzzPnqrbue
meAsnIQlSCuZio7iGK9E3EXNPX12eNh3lBWrDucytCUflsjExqdDroz8hdM4cS87Sk6Ic/KZoSZg
Ywdh2D5UtrQbodt7mgNreTLrrNTuqQuIUBpF+gNLLmqMtunrbNf8yK42yRA7UKO3+Dwn6h6LKvIN
n7z5ANtRIObGDzRH805qdk/JotSaHBQtlqTbXj1w+amN3WATJ6nIaKxwZDSAG+AifGhI/SRi4S65
ieK4MeEkKXdwb/C0biG/mBSBlIsoLmaOtu8jDOJLp2iSCfIHOLGX7Hx7Y7pCLkH1leZPnPHSqfK0
lQwAusp6bNhD1AWMy5hTN5aEh9X4rrFzZxpNux5ezX9xNjUW4m2ws3d/G1Bvf7Spbqpc+MnKu6qp
W7BNxKtuZWmM9T2gTPM2m1hGCImZa1b2tld97skrASRZhTBM0Q9VXs15VYdZb9hCqJpKzFSl5h5Z
jnmUoz5J0XmMvkIfWVK+6K57NZss2fjdbZC7WVzeCIiLLwN/wDhyC2qdK9x+tcfaLNviDguNyWul
ekAXQkFHT2UXl0EB8BH3so7ECrA+m5NZZd3BxvY25xFM2AzGMK/OC4kzNGTXHp2TWwXHHr/TlEbD
UJCHkyLEv09msKF7PRZexn3ggFq3Zt9pCFn6+6Yk1Xjy7rtWPjuh3Bo43EDe3V0JAJL8mYnUttnm
gUNsPl+BQ9P4U7dXkw8XxKrQPZxpHWk6M2NdYzcx4mnOmsE4YNYEeQohKsoS/Ajzm8fsscS4exL3
fubRtvEyzIZ2LiT3M6nErnY5zYZEWyoBupw0zolE6Pch3wn6JnPQyZgyM3W1Vzbaj0iaHuneLjjV
mZ00K95Mi/IZoTjIYYtHL4Zk8DreRzWw+g3xOJ8FXAT4onF1dnbGujcuGKgq0LWuFW7L6J4pNs+y
vtj+5ixre7vaevUZZYQ1mPKfb28xIu5SlStf8LH8EGGWTOFOJAtR51jnHNXtnCA+3y8A/jDHh+28
ykKYp+Lig++qB+le7InLBjHXCodMfQiAyiL4l/LY7lVncda4ZoIMxnCUFC9UfmxFcnkKOLhgC+Qt
rWszx0JxrTRk456vT4IYKy0aVROaoQpfmksbIe+Fo4uQ/5SNWaS3F/KOETyYczf/lI91MR7+mz0a
s1jGeDyHY0H5D7l59kzn/Jo/U7kIiQTFnmocaaMVX82HWikvU4BsTrk6Xz/2Dt+FZMTlQkEQ1Te9
Mv4n2XZJi6K/JUhNVTdLvKe+tdlHW0OqhSyosY4nxVLV0tDMYzYY3rELOQj9aANfHoinV4L+IngY
rORADFKLKDUajVHuYhB1hs3aooeNRpn+k8YOW/XPICX22ggxqRlqvVOaSmqG3gqfULBO4maVNyaw
L4RYu3wWuEf7TgqvHRHF2/SlaayDF0kWa6WXzq84x39vwwBtNeGeg4JLs/C0UmsurZsjnwdmyLog
JDoAFNAsSIWDxUXK0kHVxm/VxyMiLMDTCt1Hmuq3rIrOH+J2Q143h2ubaTrtRvQr9gAh82CR/IKS
Q1QZBeziU3kh4Ho1jj7ZgkipHTZqtd7HRwZVBfUVNgH3ew7jV5P+IRAiiMp79f4AWjFJMzfCZSmq
tPiJ63UT3EDwLt8ujYOPKO3dGUZ7qFYDqkxCQWXl85d7mcP4Slb7fNf+G8CUsRj5dZLfN+4y/nd1
rmuJOxlKwaAmJf30YcSwXnzUEsLaaA+aHKXDQZZKUoonSi6bud+47/xpDoa2QddrTg2hJYbUmsjF
mOHz7eQ5o0yDTerCei3Ct3bVYaUKEp/yfYxffO6/U9+rQXs8vb/GeVsAArDhQ3Nn1XkJLHcDMIFb
tjwVJF57zcKAHeB4Tf8wm43A+ap9K/AFThrEWqtPrSXJkS6FbxNy5i0dfN3v5Mv8l8DRD2YWnIhd
F2/xOQxPqWdVkIi2rmIrGsnPnknKAAweH+HGLJ/M8uQIVjwlnt4b0vdsjf+hQCAU9JyVI4W+0rwp
sxwUR8p6vmN4R+A80gCc90jF1UC9WwHQBtN8zk2X+CBpqNXOmIXcyUNJcI4gu4Cwd/FSsgzD5jXn
77vIxN5aJ0uahffLywalfmPemXlheDJxLyIeA5VvHggTZ94EctboOJMK4KvpLaXBnpi5FRH1D3Kg
2y33Zn/Vh3YKAuOkwjqnlHjUruDYEs36KMunMuiHy+QSjYBzf8o08CT6EjEbkZkvD9oKyXFl+EG8
K3BwCjWWK4JqyT71Tt32STM6rXklTjI+MycSIHMYyN4oVvgiAZlG3PLmao2wic/Y/Sfs8bw2qYFq
cazYzPNthICxYIrdzpRyYpSPgWAfNHPb/HoLRy0HLsg2ZhrRhlnHDjMgIkeamvFEWirCcdl3pfAg
NjKUlERVuu2p946/olq09aHyUXx0HnR76x34gp4yXFnpvPqVKWuDG03HO83tNHFkz9wPp6PvHtlu
kC8mLUYIqOnyIwE6oixJUtR07hWbzWRTzaMemYZCz5QgWF4+zErQL26bUpQmGLpwD94CWo75URO6
9Z+phAkEieerWP4crq7DtV6bMfCm0u+8l9ZDvfUuFLRg7xx7RUvcX237xLkSyUB9tfXKM+K1UTU2
D6q7js0dgcdgZ7rcQQccgYZJW7T9Fc4Rwx+tQlrg66spxwjn1kdGS5Cl0cP5ZGSz+XSVQhdwCjVw
s+QyylxjTymU43jbPaP9KfwuCMFIceyv0QwNwlDOkvtdM2yHQPxW2JPGPelD2nYQyr7vI0ZngndG
WwhH78fvzGWC+E8/xRaPk4fPXjzvRD/Pr+iR4smqOOaLvg9Xyotw0Yfv4rGydZbPnS6UVFBX2+tP
4nhkxDzPkFY/0dJ9M8ZubUOpEuaPSbHVu2W9LBtqZ7jsh8pqmvZngSC0UPMkwjjM2gKpbmUr0xdB
nphDHOOiXXYe0ZiBHwonutcMStaQAe5GzK+z69b90/wgazY2HeeHYgmkylCwTosZQvXz8L2yoCYF
47gF+YDbWZhS+i8nRa2xBghzlAG24WhZ9f4V0V0xO0EmNwIuwcKdx6LFe7N8TRYjU0lLfqBfgM1d
x09N39/CNi2A4n2b+KTCVD2TXHTRwmUaDiDkdhe/8DLjUZ4bUqWOGyBR89tIoG89p4b0yfHB+NO8
7GQIOb0kwFIdy81WeyXj6ELE547jN1O/rkvu5MFdgG/cPVuzsUFH0+tgHXQ2DFNQofO2mQYQ+6TU
uivHvx0KYsywfE/TfU9jrVzupsVrE9D+zXoXvSVJ3CtFRyJ+EXh74yzRmr5BfZ4hlAHi8LzGy/E+
zNgnmb77Ay8Z+8HbvGJDT+QSXpBzE+yQx0utvc0slTDLVTF2MO/LW8PcQq4m/mtoj+CnHHAb+giH
UMsGXDYF7srGsHX9sVrVrbrNED9MdxecJ+aq6zbDjBOAzxHyZz/iWZtUfHQMehQQHFeLm1GnvtR1
ftSF5topbS5N9/V4gX6uwDrMitH3r3qh54pmHqCJVl3EmO6qppGSFoEhgMBnxy/c5QvJKGYkPSZF
DY5K92Z5LBHNFRt8lkj62IdSW2j4Va4N7Kw6uAgwDC2/gTV1O0zAn7IGINFVkAtFJuuTvzm/1k5u
lGyQn6tLPHz2OPmzU8CddI8rf/3oBMGjFDuzp+uKy0ZgntggmIGZKCxUGyaLShqiztvrtfhi0Hae
kSlf38hG/mO5NtcKtGwtvsSGpX9hUmZJ+E44AYhxqKjK58Urr+yXJ6rTpv3DoKwdPuZbuaEBJi3G
yC/0P8wTeluLzfe8ocFl0eCZ64y9ogPWXu9tuTZYR2e+y0hmk7lv5kf5LZZLKyPzL5x2aTWD5Xos
VCHPAj8+qkH+yQm7nVd+Fd2Ddd3Ygj5h+ZoFg2IOazM/ywX1rtlJvuD6fMpsaIU//a47SfXTTE0t
4A1YFbTTjWdouIv/Rt1urUJN+uXufFqcWTkMAXOKRcaM8X8Z1BJFm7kzNlHe1K8y1ehtUeVlMvvl
T3uYiTWPpV+Ify5vPsQDkX2dufZ+vGclnRrEM0/UWCmkc+WSBxEVqIlKzZR9oj+1udwqCYTtGb44
Iwv1vJaWF+KS/0A2wbb0w0jOUB5OtgyDvgDW1u2fv5kfhSbdWxIV0nJvxCMUyMVFA8uzexgIW80Z
2ayO2PAxwEzsY1soF9s1ZiSwTJniTNDc3i3r8I9nnbhVT+gg+CQ49g4XJQ8KkcZgQufb/z8yoOkB
AaFuwBdxF6WrX4KrGYKPuiTRl7G9LAdeuvHjBihSkV69NiSAaUdzBo8Rq/HDMVKJgZ67zsY9DBhF
l/hzhnTTR5G+D7OH4m/knA0VJSQhZb8Do18baHAkxShLttPYBL469Bp1YHpygS21cNdRVxZpmmH3
1tEnM9+K01mbChic9W7MdWh/1rKILCpNgmfrul9OVXPJPb3DD7+MVN7Lrd71oaPBfwG/mgsWWH7D
Ccw2z8B6NnK5F69PWsjH8BPoe4fYYBOqRkNYSXtH9wodglGalaOJbowkc6axiEirrTQgxcz2YUJn
jrepvaTR5mMctIfrXew/WmZ/CAGny4ScDfcdwjmSp29YsTa/13TJ+3Jix0qsHxV34bQcLFHPQm4E
6qgyn4WXrqea90oQnJqRnUNm3ITb1L/n5B0RI/u1oADDfBKOBLZi1IhlrBHdvZg747PlxVs4K9tw
yNdon13tqZRDyCnEvlsvVRX2ZqqyXolb+cYl9v0f0VfCjcCvBt6ByzCE7Ub4xgbfXkwNdGbKwwnI
gACBOd+iZNe9wMGaUUEUidXrEOvvjdWY7Da4JVRa/MGq0KtBrYjpOhzgVH5ncGHGI+hCjXXtuSxO
00UKGStTto/2/gXSXjMaYylyW4YVZpwG8Vq5Hz8lcFlk+wFsBKJ3IUe5xaBdCxGQSKEVVlzaFCRU
A/eV9j/JEfWzgZggMzR+GTAma74J2xDP3iKHCeJ4Ns2Z6SylcDdAbnoZlBRMllfXdh5+Ae4G+tZk
ThSGDBukr6cHTG6QWe5m08ZbEeW/i8WXkQ0S9EvbSOPKUl6gPe+l1Qt0ojQ2u7k49nKmJYUUYytm
Jj00gM5CEGvBVvfscxdnDSCmVDhLpdf2nks5I8uepBNduSSQ4oy0mE66ojcZP/kfvUsao8xSPjUL
vlPNuEW+LyQZOIe6JUiPRWwWsbTC+gXoE/ClKL64eyx/0mUODd0Y53unhOJKJMJx/SjSaycc65WD
TTTfvzXFGgvlb/MlDCIlJT30YZg+1HggU8FtoEScBa/t3j1bni6PDfWC23kaLuM8ELE4Q2POM2fQ
dki74ODJxXdhrePqALAfQ0uO5UvM/fBNfdWVWXUY/l9S2XhXiT6Eq9KllHCAum9wqUCQYbJPKqos
N4hQhfgjsw4ALBdEco8b9rWbTTwmb9vx7lJK+LJ4CbgmANSEnbykrKujk+E3EydS6yqJno+J1EBK
4IJdj/9rFOVSuhy7VNZmYzreg3YXMeKam+2br4BqGTb2vOR4DlHs1Fc63D0dC1rPG0uwDc7emAGc
uvx7BfWEA6b2/4x3o3pF5Cqn82eOTwBM0sEXFx3Jw3o4NnoYJEA5aDJ5oU/nkiee9PtNQYZffwz1
LOmfuqjyD3NdU2VIwKXjkorWIf4xILrSHFzbllbQPqR9aBUcwiezxdsbLEUfJRILGvlP1LT1/XwY
UGXpwXTThChcBNeNJs5rrxmcfC6sJ3WlfKq3C1sL9dmOzscOSJ7jyIteR1UnPvggIPwGGE5nnQ9t
HrjzhOgBHW5dP/2UebAJVj+nEubHZ4flzXGl936hc6UBMQQO+NaR68AtdH9gW8kVBQhn+BQDf9jY
H3WqU2Ovvutq1fty1lR1Fbwm2vA91EfT+/en77ZdpIR2vIhvEpZ+0taa9oQc06PW/qgMqhZvJ08N
cWXtm8tGPE6SR8bz2dqSFeTX0tF+c0e9B/rCmFiDj2MHkDkijjqYytwWdCUu+mUJYHu+SSJWCyBa
v3gne7DEY2twjVTpY87kKGllmXgg2/ERj0zOqKs/zsORg71s3m6DPwlBcp1BWKu/VhJVuZ+Yis9X
uv+Bm4DXsbCUsJA3MqMX9LeuEJH6Jneuk5Kdq3TdB+V1ZlbwegcX/jKQIR1aaTnGll+kOvuoZ8vI
YadAxdOZhUc7xIn4iRfg0soS6P8VsTGCs958dDExDeg0D0omHCjPL7KUO+Zx0OH+GDA4Jv2Bv2UD
X6bgPNnS4RUi6BBU0SoGY95EJmDPdoopTFd5l01+vKipxnDTJbMLtHan1v6gNbF/3I43kXdopy3R
vNK75aLInQxPKNCHcbSZW2Wb6/WxpQ8vxq1+/mKL6AzynMECEuM+tJW4naJRmgeR0jhrX6aj2Lw+
vIG1FjyIBZsHejkQIQRo1I7jCcPj+1lgOXoPQ4r2OWuvV/ENfdXHRftUzio5ufRMYpFNPxdLmk2I
yQjrJap2i7EItcs9I45gQMfG2MDlpCjV1ePNG6090s7fA3cD7P96/K4IySUWlTpOIy8k609EU04i
7qZ2oGjXor9p0WV1kbdQeQha04fZHnKMZCiM550jX3Yx+9LYIYJ0ev+vE+ZG8NojM/UzQg2B5Mh6
StpVDZfeHflG+wGGJd8jCwCBYw9BqftHosYikY6G20w55sRtqRFKtpE0p0jJjb3Z0Rrfzl1Gyco/
qT41iumzkNjiNVX/M8aeN3CFt8KT0IlgK7xQYzEth78OJJvYebOdGaJY89lPYLsvT9WlbfI3DB4c
UMPihqAMXZHPiH+IZMy76MAGSTFfdRKYRySLiPbQvgu9nIzCY1X6CyzSLFf03BIURwx4/0aGyB5r
DQVS5ol7bVcND7FkvrzfFN4EA7sbM8AGgQyfS/2TMdqyOmKF4N8tbfftleACCCEtu3MaN3GKY47N
pGUcAx2Dg9anDOIgXAHx2yKLtbNboZOGLxsxZar8rVEkqRkoZZql6CsgNxQbeC5SPURSqc411l20
ywy9D/OJUH6Y0W3BWplOs7UwQzdjz+UZBINKUG2SviAGgRPjRfkfeJrcglrPBDerKnL2bOAsshOB
TUaKUaVxafE8kQjKFF3F5sk/38S2vtrlsdDNw/vu6ECCCYDNIUfH4ey+OPYm/5THSl9sAPk8FwYc
XdhAH+rYVS9CPO1mi6EG4RFqnYYQsdwn0J/E4esuJU2yx7tMkbBfymxpMykDjRniKUCk8DeVXN/Y
LPJoPMutArioaJ8xozWpiaNGjdDhOTBJ8vEH0t9Klk3zkvNGASdmTUnjeSYA1SQfNFSuD72HknQb
tkoX4d2wjgGpkcDRi/q0N+FyDv1er+crY2KDSY8O4slR5KRhZRnWEWGwDGOALHN/mGUj3mIAQD5H
qotDxbY7J6DGJlbDyh8186aIQbw8kLH3B7zJjMnVhRHRkwpzt88hwx5/LeJUvTFsfrcnDMQUziOG
zE4TV5RHrxO5OqQhmkIIv2nBe0Hme+FD3kFTNDNbNZoZ3sg112Dv+pbVk+Ij+j/Z0VdOvjLEHCe4
GdXfgMPqAba1wuBIzq8JfEMExhvcMEuj1UG0gOVfj7m+kLwnv31ZWGUlEpxO1sBacKngkann8dZP
Iqr+bvlqrOTwk+ncxqvy+cspDaAN+SFgqatt0/Y8bhq9tN7yHbCNNbDU4d1chhp4XfnOL+Geo2YL
yAm8CTKCj37ZED7CMEXfYjGNukjH5FvEj5mlTFlZ1G7BOpxkO8nelzmnRNIgQ6O7FObld1WPHu50
rLqz/gLaD7wcc6Nbw8NMSdO3wcagF+tS/ZoRYy3Q9t2VWS9aPbRVXHr7bYOLvEuAtA062nlyP785
+uCAg+uvkiPv7KQYu5gWRuI2gkLw3qANMIDlbpTma9SnvHajz0unr4UazsiJQCv6lwCLxy/yj1yU
aJkrsd+lmw3+RQLjsdwnKxHDV+s9EXYdCt1KoHtAlK8jIyR88wxfbefvf7pHKjxiw8Y5LQHk2sF7
4zdKbzWMKrYOA4KTPgVx1keu6nZ+Q4PPYiOXdVrnYaDS5h+vAEwJDCcJ0Ob2S8ndYmE7LOeghUNU
VEN6EwbfHhu5FTINpNgTMwZEd/zNFBGHzLL2Pi6WHEZnEwy5trZIFnIcR9pF3mcGPWTVRWhihWxF
dfs4APIS/rtf4XXXsL8pEweWEcE7OcDGRC0GDO1fX8m/vrAJaruirI8nRLEh1CGClKDy10ogJW4j
0itXFgB2BRoEr8BQadqK2HvK2P1yMr43d9hDyrMQDozHHXilsGn/RmhkkjUfb9tOUXy0C2d//BJK
Wg6TFnKBZHt3JObsYE49P9ZK/uQsWzsK2nHmbtb4rrH1PAZhOYEmzs6irLBuQwRkhyxOZG/Ygn5g
m7Hcvobiicr74OXyLmhA6e57Q4t+6hQ9HIy19sKWEjLAE2YnbJT2myIegGEX7yKLm0ssS+QxJRDr
c2YQO1GIxIYQkVk2T5XWGji6S1HTEmMpqK10yU82B5wuUWmfVuu+IBXBshbeTWX/e641355zUl9/
guG3NDnxmj8RxKlRqV0G6LkTd39QEJq6+ekNUK+2fj6hZvRibuo/VCitrIloQGGzsgqrLDCT3ga8
+5ZGkrjjErBs4I5eqOviRdZnIXcbZJhLS8evBgPQAH/g74MKMD9uRZLa1Y8NNQ5al1FvglVFoi6i
S4ub0bi1TsCy7ZNQQHAtxad5z3h5WQnkWjzRxLi1bxjwAsBXeG4Gq0V0OUIxPysMfDrrQVIVuAOC
igBPihqxU7P5LttnyUggfomFkBysnUZCgDCyQKqnkycQaQuRjngDHEWHzesVkKEmHzj+rqmJ+sGs
1dZlJU68/W3CRbZdIX7RkDzi2bYY9eeanx+kwydwFFHvIPY7adQXP3PMKq0QloIfO+vB95theSAQ
Hlf8JKHQZsRYLIKDZCddoMHJqxaIB9msB7WOZaEschYf5+90zCIASiqgLOMMMZFPkV0ePnfLr9jl
ZI33rvKYPdUiGphLA8ZYVYdd2Csah9EUVpB/Fr1Mql3IUI6/H4sTd1q31MCwMiMQju0TPWZFnoS3
FT+za7NPGevxG8BnnxkUVkowO8UN0+Xy8rb8c//Lr58gjKKJwDRyvpiuLCtwZTEKzrLMQ3TnEvaV
d2L2Yc/KmhZdpQetDFt/vZ56UmBkNlU7EjMC1ZM4rJTBfhFoS2YBoiQG6fKya/DmOZ37L6C8hEuP
AWVfR/RC5x8oJsfihfVDOGQwtXIgjggpCnjpBplOoQa4VP4ohO5B0JBYV9R+tMu7+LHWrHdlN3Wf
m4cGeJI0eNlgwetJCxdmQTrxi4aVNzBaYUU3jMlIEslXimX2TtBoL8pKWmqGQ8QIOAR1QoOy0x/S
h0Dk3N9zCUfB12LhgkVG3K9UV6tT1cZYi4z40worH+FAazVPclrjF/fFwC72Ju/wRrmrAMlpiDyk
PNXq8bFYz5Fop3K6YIj5r3JDqYpPoNYMsgNY+aXeIbfbXLeRkvDJ35kNNkAcgin9sIT/uGZzMefL
TWsZz2dB9obBS/y8mACd48IcnZdb6KdlGe8k7/1F0rGDvbywia8/bC8zuOYTEiSZwaTNQjnoCqU1
KEJdKOoXLdLZD/wghTn9BMxKrdqZiuGPMmJabb677pdFWhu3wf7P2HaqkWQy2+UBiEHeu+y99FaW
EWfSNRss2D9w1F30HyXeI5r4mwOpe81+r0Gmdn1ZC5N540OAtauTs6N6SwijKBEuxrcEgbpVE9xj
UqC7op35A9db/iii0MVo8e65wzwTvGk5eC6UGg/AjBb1B9OE6+vF1SGUVHntW1AhL/obWoh4sPet
ZzPoub0lv30tUGpXYhasTUqY3PJx1ST0M97eTmh6w0CSkFAiJzRiJP+jp5e3P115loJywNkrvyOA
aHXHHzJQ0OMHhJ9tgN/0UhqNvoACaxxBcfVXbgYOWqwCg3Xi2g5Xk2xi1rjwgLfCIp7cY+ENrvYl
39//p0rOXJEFJxH3P8nZj6bcfmQNHb+UGmIK331TXrBB1HH2O8cYRqw1xh2sNrJU2WcGGfBj5w63
fgzHD96GVe7Iqd3iHOUjnwdz9ipb3CDTio8vz/TWeoRDumfiw3GKuU8L9NGdciC034P+z0fm//7P
wsJvBi/bBDo+rEPrvt1GXuLXEdK+/TPeNX9rwgWmGKfn2ZhTfOWrWVtpnv3rLAqXCmZyZmmYdDbp
+uEGa3QiTDKhf7g9ji2NG8mF8GS08kdDeYS8gBZoM25tG3bNzh6KjXztAAPox3H0EvnCJFDn7giO
z2CXuWecbqIoshwOeccwBkyEnN7WXh0isnipOnkjRnXMtf8WUuXPYK0Thku1Ais33vHqRnWI7q7D
pWdjDAsg4Ty5pSJJ0Xve55jcIKNbYYZoWuKDQpg6ztb73/+Rrj/mjeN8tLxWWHt/LwQcgX6wfgKs
Rk9O4XSgqbH8WTAhHcYaqGjL0vJetlESLi+awvFUkhRHonQApbcwbnE1yYCfGEy78D6G5jxaPMCd
p5GO4DbVuNh+jCYgm9xZicUdVQxerOs0n6NUwKegqZy560wbTyEJEOGmTBQ1RYO/8+rm6oGLYuK3
USFnA0NOrGTjid1N6f3ESqmPJZLF8u1FHrcI4/IbkFFJYh8nX/z/RcGVH79SeXm9jgoO9yrXujPO
v4E36+YjpmrNTAhW4+YTK+WsbdvsrtDOV7LrKskY4Xf4abvKRm0vuMHfaeV1AZYKYOhBVhsRrhHa
twWgDvoW4m6VA8SYR2Ipe4S573WRzxiEzLjWjET35JWltOU4+MvwyRyZZHK0woiovTCCy8z9VbES
9jYDRFz7NMUGHBVhcBTQLliUodS26x7u29rfXqtMbVfSGpcgwF+moIZPZ6/wl1yqBISuokAyzCb2
nQr2ejoZokHWeJdNUowHgsDHa6zGuEM16RvXwiFH8YYTs7ukgLTBkho6DC6tyR6gObFzOidfRC1A
KRP0kjT84mWDs6M09/IV+nrN9NMmw+Twcb8RHqHKM1z85JQ/kdO4gbAaoxNh6X5DLLesMMBBJrur
I3VEyfr1AcqP+yOieptWxjAtUfWiiEJ7Mu5AcsN/FcCzKdeQtY8JdseE2j2gguSVybEwtDQoxBsM
8P3r1YfGtAaLcIwMl7fP6J0v6RKhbZj2a69QU4n4Q6IbAoBeRcxu8GDDD3YM/DumW4LXxbZyp5Si
52byK87LIn3LjryL54C4D/sV4CbwZE+ZLn2RProAxjGztsIwMfes/07j5nM7EYknc0AQuIDGNzts
eSjezg5+bvoZDQ39f49VjfDKV54ZD2hNaWOxyUafL48kE3COXiEiiyQSFuCDdg81JqrLQWJeHmlq
nrZPgu3j1INwVUVEfEl2b+0gNLFYMwItc8p4CJgn2aF+kDVJSk4TkvOvDOGYLC7dfEl9+JbX3JGZ
TbCNhXrHbs+ISs30VCd8wmVhJIFWBjBekclTdMDq3Cr3fs1lQOZZQkBDm1ZqlWv0fWWLsrbbCzBB
aG1RYsCJLy9DG1vQCVWSFn3yHbQ753ZJsF8x14M//kq7hbFRiSXROVVKZUPQDR5z1wn0IATNnkm6
PBgs5NzuMEAE2Cv3qRTcDRlX009Zy81z5b9GQrcHTZDBuwGHSZhDShnqJfoyuNvilZr1LGoVBkxs
R/AgkkhAaRrRhy8UIzZ3Bx851YtB2pvZCijW2TmjO80O0bFoxDUGT3Yht5UabV1TBcctf4ZJUJko
asfXF+jwbnmJ99axnG7EUtGvJ7fsLiM1iYFRNDVnbHs6Vs2rS9Nlm1ve8gTjA+JTTmihzpOdmH2w
7d3vGdnnSvyMD3x1Qkf+Jmc1G8BeJ+OS905JCyica8EhL8mxJbI/c1SEi0y1B6cb56QOTkZxa6UU
RRtwl+JMyt7Zqgh6UntXvw1MvM6QQPyrp50dmlbG2UD4Ew1MzBIAPlkbXcbFcjRKBu8qjLwO7QHF
SCnDRY5pnuaJHIoBAyvhjZaeDSILWTNAL9+965Z4tjGA1wwZ4gfgvZqXKblbZPJpBEBCFMRtv94Q
a9Wkj8Xn9/ly+dhtiVbGZ5gN91KxRNIVDgWJpyxxV9KlXt+jikZTXAxpiM7c4q7OYk3i/4qWrC6h
/6/h617UIkBuM7h59ebtVCjMtFRq8+NaEd+rGtqmTOmVAglXeDkPuMzJfpWa7Qak+nzhsAch9osv
TUZCidzz8ufM+HzeLaBD905s/mNiiDD4K2ztN+vsaqWTPGCmyghpBlw2JXFpek9v7xtNCQPinGrd
i/El3RvDLPTnWB9Q3IWTKr69FiI4ldcd42v1bIWkk9SFQ5A+6b4FJpD7ngPIwgdORndhAuuZ7UKO
Gv7ShhWF3SECQD9Zrvxtw+HMk9R5tg33RTK2l+hESDULeKoMwzyXkwy6YqbU+sOgFIVT7GduiUsV
SibmwqfGwcZ/4R6vUywYOn4X6cr1Aqhz/tmFD+lm2gqTbpC9MPVJD9cFIcLbw+QK/yCPlxTAp8cV
B6r4Q31b/IXN76wJyFz3F6XOf+znPstULcQGEunZuBJcEXtaVjZzECgmyqTuQ63ZR+/ECXRyQNMP
eDl6BdthGus3OcznV//+IBmuPnAA3cY8xJ0ivkolc2BRxPtIoJL3at8JywOyN8XMiHWECmYr9+Eh
z5pcZkTWddqOLr43rjWAuL3k8s2gkQP1eyc+ItK++tbXtRW25lKmnCaCAxCwBkPIEWbEovcwKpbw
PwAqolLHBk/4uzxqijgM9KXSfl2he96vJzrOQozOLs9z5CIBBReJyktw1BBy6ZdDFoPDYiY1i7TR
fo7lDz8QsnUhooN3AJlMsnlXPr8G6GRiG5UA4kSF3mT1DB/1Q+6nlbA/rulzp6G0D9dHeeWkbcuS
Pnb6T7lOq5nLpvfQ9vSLi6hT2KzJeNLwB78JQxM94pBhopP2UIpkTted5srynEkVpptkB+GVUryh
Q+vF567DtAFhiwVbhprg7vZyZpAfxbECeV36GiK3770a8gpEbLhb5GMFMKyNTk2EjKbtfHOVlFu9
xw1OnXdSs22LzEq1GPiIzDj48OErVLhjyMFoy+FIpNIH3Rm0OnhHoxP46HCI9ccQTDLauLiH3eY1
1QUyYEgiXoYL/fTQSBE46maX2OUz8+kdvXundMd7hk+/YUGKnWunrl2ZGtdn1ux6DsXzFSJxoeSc
UgT3TEDxQQZUs2k0cXarcmjFyQWzJq7co7aUvN8/XTjHJsiP9KAZOSym05z666gQaRbwY9cuzhmF
EoteZ/q0QnsdeIp48LSM3JFjgEQeC/xbVHAsfChjQN4jft+xPFV+qry6u2qyci0HdkGHSatK9T2X
6k1E7nUusNWALofLq3ZbDvEiqtscxGo9Tjk3zA7BDPRsYKVXe/wSiFZhEl5JJl3+fzIC/NAlmzrE
aX5WMDzBlM90DWdUvjrD0nVXAckTevEUuamxtWVoU2tzZCogmrwEkmiI3jKu1SYsvkZUOUz5iEpQ
/KCVFU1dLJVWOR9mbPxi5NFb5Qwrpd+uf5UhV018PePf2AXHlM3kTI5jraClAEMIilZWgpMXQ2Bj
EbmZchg0blfr9E2OoESGx5UG3ScVxgiVhoppw1vYD7RxQOMCoyLVxsdqB29KPJApfactUGBlGYd2
Z4BNazlvXRsWN/eZ1/jNAlSea0zzpPVMIvr8Hhw+uBbmZ4EZBpYyYfgWww9CJJC1qiq22+9TOPn9
FLnFFYTEq7WqbD2nc2kWmMOa/c5K7hVyxdCkpviDF+5kPSl68UPru/1Nl8SMaYvNwnArs9MpP5k8
JWH4OQEM4+Y7ADC2iqpC08TSz2Lx/yQUmN2kldItCD4BTon+Eb0fZOVDWQfLc9oOxkF0GPalXQs2
W5+JNRMufyDSOe1bgIXdXSVnc4EDAOTDGLmmwb3zU0vWQFW+D7dus3kcS28PT/lsUDMoIxBq2Sje
VJEwPog30IhBRHWnjplvFbeJNURq31e4cgKoq9KgYUqS035UCeFvR5JXKRLPxNI88fJBiRQKHvDt
5tN3KpISMo6uKJVR4CQH2vPTh3GF0Dn4ZCuAf/AqcxP9Lw01nwnpXCxRjy/A6UtyqC1w2QCu7WEF
/2N/9fg9BdaqjwdU8Rh2b2z8LyzJJSx1vQoFVnjH/e2xYTi/0NO8uEewNYgxTlraZ+tkhFOaKhzr
DjsSBLDA/hL2+oLaEIZSmYaZxFAzhTEXSs6xkdDeRuyorZorbAwLJD0i5eanZP1EAsPktouaPHSx
+tfZpfIXA26gFZmemgfDPiTkwRdJxzxyUkIahyURqZivSAzpQKNr0QyPXc726/f3D0qFPguXeqyL
3mVljUyMnpdToC7CUpdsRs9npo7rHfbCyrYbFEP2/NXGBMZwGoadZ7Ew5/LQg49qUSvF0bMITxrY
tPoeyZz0PzYq2gYfoNns8SUAxeaw45uEgPAdW0G51+pES3aPHKBn6d6Vwqr9fvtmahu7/dBeCqkA
PwveGG347lxkE8oqeDusejP9NR2EG7Po8fk31+I9BMr5PZGBWGCmSrlluQbdbENA6U5tDN0Y+aQ8
/lyS3vMF2eGa0nQLBoKxw9Y+pJv2+NjuqGxmhSPkOBWtW27xFaPZZIqS6CmScpupLu2trQ5gQ9an
c/o/UjUOgZZVlk1nBz4VslZ4S/PFVnTF7Pdr+u15FceEQNajwbLVT3K8FGpBW+skAgkM8v71CjIX
t2AguFPQZkx6nw7moGUZBX1VIvUvRW05ekcqAe5OOFctS+3xvVptsN2PVD2lO9o2z9OtAaanRRs8
w3XaCsT2Xco1cAc3nRPSjXpRDbsXsTdKH7fHxWeynVPNLAZXR2+vFOrZWlMt+NHyUsS98q/1pKav
e9PRgP+2MpZnAMrtVtnFNiSwW6mNNxiI9hx0Kp1nP6AjEOcTWMuEbAwHeSdl7q2aBnR0rGFbapO1
fyRZV2dOYHo5vt5rYoG1TrC8+ZcLYpmHsKWf+euNNqM9DUbJJD8DeWkb5bxxk1mS4awm8o3ShedN
IEROVsP2ee8az8n/MWwmqURrF0BS1LAiGizbZNBRh0szbupSV7d8i90xAUlt0Tv1s+4naRJaKSMK
3H5+3Sh+VwXRRaziKKekz7Pcdq3xzPe+tWEyVSKnfwkMRFJMorMl3hCq4om8A5tvmxmxltCov50L
U5IUfTyQOaGK0+8BsZWo76dr4xtTMjJ5CFsLD8Tst4tdxJky+cJVkuCWgD/X7zeIaS9LxVb1KLZr
rsoebceUZ6L/18n1Pmz/pOCRQDyOQWQb5rz2i3m0AFBLLPzvCCNeJigDZpoQaZr4DSz8JHNyi0BL
Yb1M48Ra0JqgfIfDmu10sAU5gEzVKxVReKiVSDuR94KmtFnSq2O25cpBvl47ZavZ4fscnkxCGFUq
6TNG2TZr6dALEaQD9xJWSYVSxDlkxdIn9qKQW8kJoqzpDCdTmS3ca10UzP2HFKMK0s+wPOSxB1OI
wuZ2kxD51EAye7E1hRBxR51ZzlZOvAmIqs6xpecYEtDyI8k/g0wRuRawG4oP0vBkCZrw1yoiqYVx
RYpVtwCipwes8PI1HQCMVykqx4uMDVXhZe1kmywrLJtQs4eD5TCoQPzLiP8FbT1FHagN08RCaCbc
nO7T+CUbtjAlzvPNexL1q0hsQrSdofmFbRMTlxsceaGbJh+ydbmowp4GqRGc/7OtY3WDSI9pdqvh
WGu1VSWV8bgGYfxvYuXPIaUtJODFNVlPcdmkZYMdMRerIaChvS3QXTwE+bcqVcjR+2KfivdIXJwb
8uY8PI3SG9fXOIUobr5WhbfNfJtBSHW7CpycTEQwY2z1ul/B4wH1KkoR07q9U/VR/C0vfCSevEi1
8X5ZbbkYvRlB0SitbI5hXp6PnSecXAXJxwsfHzZJNVkf0xu+MmRq8LDi3DeGduQ3MM6aSxiJKjBV
8IeHI0rrxoKIOO9hoZnDP+qiIR2kSGetTFoXNaXk0MUOZaABJUEvG2jfE93CgX9JHNGz0NmyjTHD
4MHj+Tanq4kiCD8IXVgkTMG/yDkoCR/Lo+guzn0F+0zysfGEZpbv3lizSfG37EMeCamSr+jyMS+7
8wICeZKWzjbMVwrE6a+ClnVr5uUrO0BrpcDAe1SvLS8yDzPu5CtzX33RueJN9MO2JOkbLfBV+wV3
fQ3W1s0LagmmL1rk5EMITwvV5QtuN9e3TzXSBhjFnWd+s0WlXGURZnY0XgFnuGCTwVfeblAFOr4k
w2D1n+saB/Ng6/khHFkvcVRcHkFlu4b+YW2815UPALchULOzXVRqZTfd9lR08eyiUzEF9xhDKYki
sSLAPpE+6IpTvGsbE8ITjRsbSnfWSnjiCUSIoEvd9tSfjRySpKQg32E3Tv5VXQDw2atGWXj3i/CR
WvtfjtA2FcaI25RRgxRJts2DR0oVPf4rwD/C5dzpZOHigy0H686CReHQ9GGWjVx+do1pkDwHAX9M
/kxWxW5EfPTOlLKDyOCt9wXKXc0/Y3Hj5LYGOMpy8xXDMRSI+Sn080MaocZz4hzeJMLTCHNO5ebr
G3DxZJmmQPcFZUmFXKkBX/fylaw6p28K/mAAskUHu6EnTbE+ib6Vlfd8z31IVL3xtc5T1uXnT9MB
wgcxl0A7hG4OENl+aw8umM7dFasywy3o28Vfc0Bz0dWjFyc3TeYPQA/wWLF9jsZ+DWU1xEHDR1BP
d3NuwguIqgcqgXb2U7yzLhLpcYu3Ajp4lJHTHUcUY8cnWSvbPy9s6wFve6oM/twp7zWVlQPjFbpD
RePbOvGAz0KMGtY1vjcVYPCqjZ7Mt7pdwRxjU02RleQyA/Pdkr15lT2NomfzSM585OTppUkJDuEz
0JxEiCelyDcbF/82+qNBBQeCeE881+FE3QZAJtd3scdbo3zj8W/VDXPB4rFiYkdTWWzcXcKqYslu
mNP7diS7R6njKOJwnb21GYaUCrYbtFV1bYDjunQV7H6QzWYbLL4ly/c2nTOCCe1KfOvlVtwZ49Xy
fySbHGaA1+XkmVmaIcy2/nD7Gm10KwHqydF7MlhZfRhZcvq5oTYULbrM6CHiQX/e2rBN8qEkxLnS
1N2k1jEPfWSQzy9P3VK3UdDDKqwAi3p9EGuPRS4qv/jOfQZlIdSWv4A23gKj2A1pxYgPXMfsW2aK
qUE5BggJFBRFelRlTXwkxafL+p6TQR2y31HQ8gNgqurRY3fFthChZy39WJh6V1mVl4hR27MPSGLa
G3c53TqiaFO5WK9tphrXwZ327EhO7N74c/Rzth/wiO4ozUbvuMbfqaBT2RwCk5mSU/FPWeUdfnJ2
R2qycWl1PAhhOQSen9G9LBm4rhrQ7rjzHdo/MHhKDgMrZny01z6ke5f5oR/zjjfjMaUMQr/+D8jQ
em/oVEpKABwifwMVF3LQmrJojw/DRWRNt3WgERAm4lNaZlWd6jPwWOB+IYnpi9QbzBUPtLlnzGlV
egpMa7HZ2Wuulty5Mz/vpPUU5HSkqW4rgtBhsnD5+LKZ79m5Z3iXED0/RN6zlOtSQZmuS2lfbnI5
SUkZxfo/4be1mhTfpwQPRRz/ofBGnEpw/6JJaSGZtuaVDYxcLsKXRo7ThRwpc/YIR32lXpfRVD7j
ao2bOI4bNUE0Kg+/P62W8S6aRRgLt8IZhlqwmipbumkA62banQP0NWzTXPzhY1psEwQxfVVOD0u9
9sWwZY2PMAd7NzjdSbgrN6/ON2kGbRx4ELH5iEF3zs1vCjW3uS6UALBhoiWKRh8TUCEYSmm1sIUh
6H70b4tD44LyJgoNO+ts55avhUafHfFrX3sKR5icriUJM5rzU0Bk+HRyXhCd9ZpXvBjHxl3MXSH0
rNRHG8FP+7iflMF10oNBtpZg7AdysB3h40GQO6tcJpTVynATxR3lPhu9til+SCggCpgH91anBIUU
zEmVBGDFz8UbR82XA5fVi0/VT9N8gVG9bfC43RPtxA1LZnsQ1MNMRk5wfoepfZmu36szVFYqi8qK
1sYr3XZhKq0V9Yd+NqjBufz5w9yP1To056N1bEwWRoZ+EFDPuMwEe1lyY0wJM/KnNwkWb1XcFw3m
XybRkjcjIPE4mXxFMLGwmRaupxBaQ0VaQ7WVv6MHIJnPNKbQIRUfq7b8L5vcFnJQa2tMfdJC1EJa
gxs/m2xiQw3I57Ler5qq4ZcugLBWYYOCDPOcFbMhQ/F3EJHdAET3H25hkDBgZbb/AULSoMcmuj6f
R/BE9BefS7MZqHXMQ8R0nrmU/saQp6MLFbRxQ12qNGQXrNicz/1wYSKAkyx0T27jvGDWPBPd+tZf
Kng6ciKkJ9fWosQt3syn0XeRzAynImsr95846MkHXVa4CbgBP4mRNn9LbXy3Xae7vUsnUj+ZXdPe
PRnG2hh5kgothHczLUymYO/2sjAuIhyMA3jCSa11S2K4PrejbHobfr6tVaQs6WuZBMboiyqIAFGk
mxNAJ+vU+ruFW64yOb2/QoE30HBYfZBiMOOJqBKKi4AEB8Vhq28ddKTWEuGghqAkfmQ16mHDuvWq
VokB9npsK947kUrCb9+zqbmGaTb3az1Y76+U/e5VMSU7gIOb4pKnTftvxkU39jWij/zd4kAkL/GS
meyuqmWK8CPI9GWNXmBQ5VDsZbIzbQgH3JAf0dE9pYc7XFnCB27kHGiP0nnYkF3l6GXMSulGQmns
xMcYl7XJWsg7qqLsClSyXOCTIsyiy6CH3GozRfI06+NJWghafE6HEasMhZmJf++Wo336jCpAqYn+
QKpmnV2hX4EcfQqWaYY7wLLgcftSB3p/qrQpk+Vh2N8YE5ijDnFACSdbez9yL12zydF74juObZpp
JhilX30X3E57BNcLvF53je01KVTN45cn+0Uz5AluZ/ptR0dLna3np9NgbktfzO9A2xv91MILN2QA
jZKbEs0eJLu+fXLXG2IM3vECP2JmWFQ2xlQjEeQ/qzeAeAtKHopJEfAASZi0PcZNc4jV09TWU4Rz
OwEGdo4hpYj43A+TQT5NerJh5YErAKwV8frhb3MY9nQg5a7m7wU4sg+uUC51dufBAyQGaMRSl+fI
QVg60+BN1IU+xaFbov4lEAV7Go4YXgNmkyz9I9dznkLpfSCVCzZKaoG2f49C2vV+VHJkt37Ru9Ul
sRQ22g/jZCdxQn4Plu9uN6TFa+j7zkYL9IyIWIcoO6kHqnXJKaCazLrT0VtAYpYShxy4rpx9xr4s
4s9T9VdJzwtW2uhPrhZ/lrQvl5gmDPoGHsK5weHx2A45WQwnCe2TXsKDS/AiUU7TvNq7rJQjFRZn
cEwgsbncwn8PCkRr60hWZoZwRebIV1qijESm6TrrkZm7gvC77LIF/mM7Evi1HV5Z0qgN/b2hBqmj
FIpp2zNDsksOFOgdSAFqPpWktteMNQ2TgQ4f+x+Lg85ATAwsZn4lD3MUWRA6IdDsQlrSYWt1aAZt
2NfXtq91KaFjklMG/E6s+2ZjReRMxCbZfFGxjbiL5GOt2Krj8LcYCTOEsfKIIEtZUgfkU1Go5Dh3
7mbZw8mgz1x0On+UHh/XUXZh4G11Q5tFSEcatQZ8cF708o5oyC8Mrz2+MWA42YPJCf2gQXXNJMkI
zfS0YwjpK/yD5P8pDv2Di7FW5Zp++O/RdGpO3LcKAF/0bCv4HyRHvxc1MOP6tntpIDdlzq2cFBpM
nXF/nDo3URndfcCiVOgCpXJmmaSTfjZMh1AfXPG8E1PjuoBg20ej5sEmibXx9fut+VK4JHNAiPP/
FpGWImHvwLKcK9ZOaLxGtexzj7LV5NAev0MjvQ1ZZn4/NYfWHbu0sR1WjfyjCiTggAtOfgKMXd7y
LIlWm6A8XyZXI1MDtOqTY1htTgB79hDfHH15fyRcGpU/gClDWm/kEqqr3C9mbL4WG+qpApf8JBMj
LjyQjznFjMtRl617z0xWrkZuVzFHiSyKvWfksIXyzErTMSEKHNBK/cH6g1hVTcnq3HWPVCWkZueo
WI0gCDXrZEwRjeBJSsDiJ8JRO5yw0TRRjgforEo22bBGeI4uTvRIqLcax2c1Cg9vpEt/r7TDI52p
PcbAxIrn8zQEZOMCCP9i8cggkYIgnRZOh8vIrYCfGmIFpeI+2s48JUV16VLGmWI3uhhzpW3+ixE3
IWUql/nfQTpykb5UKuaCczak8ltqnesd6fZ5VwXT24pyWBZcLtEonmYpOUZ3G5cdPdAKP7lRlkBw
CeFlBwNc+7YT7Igrn9CAnF3WyAI6EyzyMRrjDaPoZ40ol+mkA7BcKa3KmvdxW/q6po1mFwxVTP7w
+ajAc0ZH48vOPVtCfId6aFoTc956OoBthbJ9u0RndqOgA/O9YzlfSH5U1sQBvCshdnR/4CnWEZBj
fEETutLjCticYBE6hlQowwT9ZmS9TI2iOM2kDDdVsrnCWDUYJN82GYW7B5qw15z7lggCkorLJWmS
Ruk+KMWAL7/z9ovK7mUAek3pz1EhQ8XCCTOk1r7vr0j2eii15ytfYgrsvnzW4aROQqzf5OFR4kRM
hTyh7fqgGTPOQdDINqT2fL1+1Jzfd+41G5EvVB3f3FZnCGd4PGqUHJLz8ZFVAegqgkK/L2M24OlK
8Kyx8EpWEtilDvm+/h+VIfmebKknoPc0bf2emq/m36OP9BuWupSiczVhkkHQawwNZlbilN4XUc+h
tAsksJW/1lVoO9ozjK+nf095QmjAohB21m2a0tWM+98+uAzHnGXhNswUX2NkBkRR/B+FxMolmjS/
/aMx9clADEdyCIVFlwDYJ/WOnX3FpaA4pUZI0ls/ch7n6oLEtyjx+lsPN1JVpIgsH00kDYljO4fO
D8BQ/AQPy58lzgoN4eGnhG5wH+pyHc65c13JaiNnR0nbZc3SjjgbBweesFcx3giyAAMYyorB8br4
S3QXfqUpwwbCaD4BDb2oNRVAFYZQlwkr4MpG2Pdg/1Dl7LevFGW/7OCfuoAGWgtI/W5kSTPbFoFd
SKHGdgAD0JDtfA5+7gZPKRRoLWuNbVNX0SAH874MI3PqHwYzOrJUNt4py/1vc8t2PTVLBZH4j8k8
UFXn9dV3/RJDuJ5Qeupp5unPd948eLOKlF3W2704lwO1PPu0SpS7A6jPRDBEmF5ML3SqsumKaqsJ
IQ4RXo7V9HcSjImnaZxPr7To1nSjr/Q6HmCcvbN7ItBjT7p1hbfpjnwivLM6c7DngReMHHHHqF60
1FTE4/mBaA5O7yiuJSt8seHQrH/yKRr69QpgZvXq3/QfZvI+bMQfCc2lRqN/5pzZvKfhaB95RUmS
okrPjilYqDh30Vafekosphb+B84bv+7lXb7zau52LoUeZeBPCvaqj3S9hmrxL8Gdfgqd7NnCis5I
CdX4PfSYbbxMSFTpjvOwjV11bKEQmK4HYiwhAiF6Dj1WSlWav03L29ZUf5GiUcz+bwe7ygnFj1gm
UUg2RB3V3/NB+JCGITmPHDel2BrD9LcQVld6D5ilzYLjgnaQzfAPydlYkS4TwmdCUSo029XLO3lU
zTfsiJAw3eqi5qooBSHbtdQi8xjo+5qsLDutrkzTwPU59NVcpy1QabhwJlkslpC5CPbLfUIy7ci7
aZRbiWlh9cmJlMuM32wh5thyHicFUhWBI4s9H/zb5N+ZAYyaH8nTHk5IIY0qhmnKHXAmBhiuNxTV
Q1jX3HdOsi9E/RmfX/dHgkUF/FInDV5Z1g0pfbq2ALi338MBgLFAcFhlaoIFqOHTvY/s6oL4eVgP
kFgrFZ3EAi1ymrfQuo9J+k7ZnFK/WOgMKBjJs/XNvSCaSGjmYvmS2g67uCz8xXHSeiFOjFm3oulq
mKfUvfcWbSvdOhn+3aSF5BddjEHHabnnrSYzWzESpps7lwF33JRbKQRN0LIiIzlC9GkTv952jlG6
dLLW/fkW8LE7US8HHY0+TBqEh0Pm13c38dCSPrGyVezYt7BmKRgvQToOdVDFkULnWQobJhXrU0Rt
zoH9ahi91I/pUdRUX5cSdHhMY8jNdO9od2Y0S7rsySSPOKFR5UJrFsN4nomB9FjCMPEiYWglI/cw
ESc4LKMXMfe1TL/euJ+cfNigPJVf2WX61pacCGYXzj7dHcU8SyyR2WPk+34xwV5UEPIT3urgAEPD
Hi+teqlMhw36zEkQpeLnvog99J/ywRwDXlKigvJCdjSUBhH71pGqKXe3tXOyLxAZOxvlHWnHYbVO
ABHqPLWJA4Zja92Mu0crtXU3+jhmXdTI0moYb1WzzQCyP7nciE8vgxHjunLNd+aixsudR+JoYasH
J/+FoS1hbEa7E+Vvh5YsJ7qXio1TlvO2Ded/pvAtwX01pCStxzedWs/wlc0P+6xGHaRW6/A0lKFw
aq4oZz+BLo4zIR3CqhGlDx5K6NEBz/qW5zOPhMWsy8C21a+9om0UZktm2wsgWFV83YnZLnDRnQCf
jvS+JaB7xZynVahb72wM4szXhU6GiafWSz44ztJQnJZIA9PluImi4TQt1oJOmT84zZceaGj+ifMV
oeEgi94sY/JizqckEYVvIIDoETbUjF38Qf1deMBdnAVoUOk4mlF16/GfCAwO/0U+NE6s3zA/ewhq
u8rtolMJLscRGnXXkFTV2Jq5CRhxTFOqMkT58+IXRchbPacVU5NO5u5Qya34LEK+KP9DIAqsBblg
SF3spSdmevOjaoP0FZntd1qBtJPk+ExPAFiYUAdsTttxLo/eaZEcAU6wk8c6CRMfxJF1KZf6GMyA
HzKzWQzmsGV1zv/FI2yQ99CstYTmgOnWGr3NUxV6YIQDkzmGihmWu9mHXTsxWyQfe9YMm8Cm39b5
JfIac7BG9dKnaIDvVVfFc9D+ZVdELUejaMHKzT/BU3eVfvs9es1SYIOF1u8+K3BsZcgZawAT319Z
Y0YTQABz6bhG+QZ5YT1NKcL6BhDcuf+V04L7IimYBTm5ak0VyVotjazvS66MZ50kSQ54pUnlq/pQ
u9bBSXVu+9TgmIW39KQ2FHWq74WSYPG6km40uUaKHd7cDB3z0tCUubNY7/TpL8SjF3HsZ/EdMpBr
ftuhOVNhenZsOqYL6kwMd26omTY+5OHgJ5vVPe4RVUCA+5trfIHHAD9Ga0pk6zhh89YTO4I0NPyj
N4ljMnnzaz7L88+YWg1YvxMEi0lhGJY+Th5Ptic7yeXnS4X7XGrxGxtAQTHiGQ6E2yYwEG85oyWt
3ImFPTioSrHEE1Nrv+EYkMiJQ7ialfb5uqpRUMT0se+BLHGTX2DuYmyv05Ro0GztZUgNGSnmXMtC
VoJP8glYIj9POux9gy79C0UcdE2gPDJrhjGy8zhK+CoHNLP15s2CH/H/q/6i1cL30dHXg193CTJo
pXRCErfvg+wS3CgNeKrDsB9X1TO8/Rfzt65xLNlOKic8CNPVRUq4+NfrznP6z6J4HbP1Y8KhHBTL
rLtHEwGAQ+CBZ9qg0Fqr7+ATzeVV6qAZJsPB+nQJQsFZwFCJ68UveeDHdoGD0MirjrzEibnPzze0
FiDONrdlwGklPE98fVBJgxj2uhqxMmWdjiAVKOPODDHBK4ClyS1dIJbsgWpTncU2U3A+JeN946TD
IUfBX9ZWhVm8a0uvPH3SOAvzzBswP3r8gxqP72wUKUEIJIh78xWjhyKsdDo7Sx2kPeo2QGwif/8D
/Fm2u9fnT0pxUXHt1azb+t32VGTGGPN77a1kkeVrS5zcisqx7zkugmrG2Aye9cRxJbTJPXOjLD7r
SqJ2Mq/D+yhnU+3n2wHq+cvFYfzCib7KV5glbzEqiWe4/vRv0VDjlwoTS5h5ofexAZkpTErmJA0h
j07fp9wIkm/a8WgH8voW7iXRGefMmejDvYnSNQObKW928dP5fL3ZbcCOSoXigUvHLWRU+Yv58Czx
4wKG9YvfuwlQtgWJ/9mjcTlJ91UaZ76PZjIrTQhjgS9gGsTS8Dgd18/6bcy8xGYehD1RUOV1CTXo
SY6lmK2FrvAIDiT7dL4AiRcWoRQNC3wymaYCtiJMvg91WAnIXTEEwRtVqqAO/9it3mEPuwbu29uc
1JBsy91ngZ44gYq3uDOeU4MHxcdI0/BW1Ycetcwklkxx9frVjjDlTeJYAaQhgTRkTcLuLOqGy8B3
5LBnu4SNIE7q7z4iONlfWQ6LhXDdWJHjzPYxT27cmwr4mMH4f94BBhHYNgndluIL1NYlsKM6z21A
OQrYrfqjQg/K9QNQz5laW9TP93z7LpagwFbCAsSzxole010yMRRTL0jPcGuy0VhCci69jRsgvibi
lNaPRFuUKsPXOaKRdTj3ZP+itjoyIrm/bW6iY7RrMzWvaqTNo0OhvyQg0Dc17MuNEIXI2kh0iur5
laARHpdNA5aUdW5zsVxAgfs5Ey9j0BT9ci8Y0TW3SCCiXd2qmC4EevPuVLW01ebn7qbIt9+04OL3
WKPwAfCA19mnyY2FL1OTES2ckbMIqxowgQf2/gpVIzEmE9H6Bz56Ga9o9Gmg1RDRx1Xg69bTCJr+
m6dKxSgfWXdEbONIAM3GeUuc9QJ6lqwANGfTI4dplxC1EETLL9LuN2naIRboGsX8rWp/iU7oDxsG
tlLTW14yJx8MtlYCst55H0RtdX6t6IFQBkT9RYA3LmTZv0eVSSAzkNlYZfMTpBmzNB6EWQBLBFi1
34MqYymFQTGJKwXr5ymbwFu1X1ZYYjy4V9ccdAHCDoIz46V9Mm+C44zoRIdDYTY1Sf7UqYpWOzW0
gf/OMf16gTMmEI96mTLwA5omOKeAfoHQbKPDl6V/bcFp1B0Ud05TyNsuXywtNhO33XUFUiU7gaGQ
8m5Txzh2bbGFyDW9IuuHUe3qPdJ7nFwytw33odA00X3q0lmwn57VfnJRrEPfPoGn3+TTHvFLbK+Q
i9h7icVHYPaNrpWfLctQYOjLeXafh8wb57uSFn+uuIN4JjkzMKXfcCINSUY5MvML4ImKzV3ZdFB2
a0RTf5StSayBAsgJs4REKlkZlvQYfqC5zKu1xcFQDMgC/IDcGU4Umi2I4AIR1Sz3KY3g0HKTGlWs
mpLzcVyOeRJ8q1LUJg/Ep4UI90+I
`protect end_protected
