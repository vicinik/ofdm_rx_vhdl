��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�@�9ڇYc��E�}��;B$��9�=I�ĥ�}eߕbB�O$֍C�(_+ͣ��wa�E��ߦ�x̒�,V�Q,�%�w�d��ŭ8y���=S����L�|��{k��UF�v֦��}ba�ᯅ:��g����B,ܵ1�-� �pI2v��k���b��R.v��a��cH�u�J�AR4����c1�:��2�1�Bn��+PF�B�$�T��]�:$Q� tԄ�O�&�b��%?�����o�V?=�艃�H��#P8$���?ެU9���+WD�$�岫��3�>#���B���O{>��1Sg��[�������g�z��.d�/T��&_u�17� Q��4t��A(��?f��نZv�qs���J,��>t��s�)�]�l�>�,���1 4i�͚a��mk Em��ȯnNB\r�g瘢I�ʑ�'�M��/�.N���8�]��@�g#��;� �6�	=H��F��}��{ڢ�/�w�YOH��ǨO�l�7������e���<g�R�eýڔ;OC��R<f�K���G��8�*�/7��\�:��R��x#e30�W+�F��\P�'M	}���%�`*E�
{c�6*����ыjͬ��=�ͷ)i5J�h*�U��K˖+{+܁�6S ��N�'p�S9��a"�y���.�&	��pK����:a%���Lt!�oO��S�e�!�N/�b���z!����rp�s
io�_�	ôw=]Y��3oϰ���OaϢ��eNL/ծ�C�Ђ	<	.� 7�+o�� �����)j��F9��|z����C����"���D6f��,'��2�[J.$�e�[9��T�y��6pw)���-J����)F��زڌ����(|^�������Ȿ�RqՃ%��	Yо�K�{����.�`or�3�:�$�x7&:3G+<h��!Fh�_z@}�4s�˺I��=�=��b��S�3ו5rc�+O��0���*.5M�K��#AJ��CH�����c�I)��o�#��ɋet<D�:�6�Ac1+��0���g�?��e�[�Z�E�@��O)�A����37t�z�P��5���0�C[V�d�n���hi��Y��R�r�8_��Gik��	n�ّ�"��/@8	��[��>��m!�t'���o&�����]�9A��ŷ$L9��h>��L�b�=[� ��R�b�=E�b���d�e��*��qm� E,�cܙ�:*{2��[��Ͽ>�V�fC9�J���?�:�f��|�k@�TKqY~`_m�K�c[���B���"��>T�oi�����A�SI�v�wD]1�`�^W%ꟊ~�,yX�7�c���Q8�h�dŊ��� %�OQ����I��*h�n��/�l�s?�|2�n��|@A���3Z6[;����&B^0�y2���툵���-N�k"/�liR` ^��2[N�y��R]U�����ԩчD9�� �
^ִ�u��/��0w2����Cg�nG1�G��x���<�8�%7��>��}��׸�"g�R=EXұ�EܬЈ�.堙�
H�0��>���?��ܛ�>�Fj�+E�"i,�����?�Pv[;�:��À��˹�=29fME?*
yہh`yH!�"	w@A<^X�a��(�}��X���e����(�74�TH|޴lėeG�*�u%u�q�bLd���I=k1�n�+UA�F�d39���$~R����|>��4DD��,��L��>*�����[N�Ar#����+T0P `����tŹ_ӛ�%Vcx�S@�^{o�Eʕ��l��O9.�n�j~J?� �;w,���E7?���	���'#{2���.�C��{�jKl���P�.�,S�ю���'G& ���3��ܵ�/2�I"H�FY�c�p3�Y���_܃s��+jl�2�O�u/3��=�������� =X�(�l��+��8^/a�����j����]�ZU�Qw���?<��>�ؙtT\���W
�:"��U� �0@x~�~@o���f�P�!SĻ\�Zv��]7I�a�aWy:0��{�`9%�E#4 ����1��:ؼ��DH3?_� VCGx�7�M.D9ʼǭ���@"Łd�K���_�w���:O*�fB	�B��@/a�
&�!��B�9�!���ƭ�h���e`�p��Ë'���Y4y���J�s�X��B��!�z�3w9מ�s^XBu:4�ȖoVM:��6��:������Qf��r-dc_�%O�޽�9�ǣJ����&I�J۶����i@����Q]Cn�E]^OީS���l~rp�1�e��'�-���v��%<��P���O&���E�`J�81��� ��\���ĚHH�f1 0�.��S�'�w=#��^˕C�oʠE�j�A_���?�/N�$���[<G�N�O��)ӹ}n�C��<R��J�����\+}S�;r�~+٩FO�T(@83�(��zg�2T���b����� l�����K����4K�1_������ί^s����rBJ��U���I��b���\j[l�x7RGD,Vtːmi��qPK�5�+�) ��w%+��D�>�B�QĿ�y����TF�6��%���09ee�H4�<����Q��Ԥ���nM��0\ΥUyv��ʬ��c��h�Y��r��U-=���0�w�1%`b�\9���=g��S!\7���c1�h-3��"8�/�v�=, [�=�Z�:�i���������i�Eڬ�}xk��1�/��g�\����
uU�h��{^چO�z�����S��ϯ��>�Mt=30r��*Nr����x��.)��_��z�s��ѐ��dy�g��w��U�IϪX� C>(s>"�1|��zq�C{ޠ�e��W��Y}��-p�v/�X��̘p�*�����	瓫����͢R��B�l@�r���h���c����qv9�.�u?�N|�^��<�"�4|o�s��a��BL���U�JU#�T5E�
9@�<�v$Hxz���$O���Tw��hM���PL��Vi-�r.�g�	{�]{��à�Mژ �z�w����3���c�Q�i@#�J��p$�f����ړ�C��G���� GWL0��{L����B�������-�=j��g.��'��x%�^�=F(Z��MXl�D� ��W����nw���-�)؋��ŵ3'}5�x��M@�!�)�"q>�z
��������H[;$ʷ�A)쨇;!���t�UC�Eb~	��f8�Do�q�em�N�*����-�3g�c抇鶄��d�f�g�q�m%�>:�x�߽��*����c��	G�`��I������#��U�{�'��zI�9��냱ʗ�.{=A��W���X ;sӒ��r� tOYC�4)�{�I�?ѐ��~w
&���O�O)�ܯ~�<7;���}��n��l�j���a�LDy�Xg�ǃ�\��d�qf#[\2dß���uI���G�b$&�S�K~	C��K��#E13�P !s���2;����o�(7���bـ��*��m;�l�U�K� 
���"������q�(j2L�O״�L!e��ƺձ��;��6:�_H!N�_r�*]z�Wdͨ#E�lPP(�����<b��oxn�U�E����57��e�0�Xh`׍�~��7:&U��D��Z>��G��"��
6�D'�q�����*dv�3�iJ�\l���s��(�*��?�S*�Z����@u���A{}�>���p�=C�!Dz� �&s>�Ag������@����t���ҽk����ͭ�m��G�:����"�q[$aJ�uE��=/3I��&1���`��I�I�!'�L9�T㬋|�1iLH������>�[\u2Oy֝�9���M��v�y_?�WNA��T����~�|����]o�� �b��`�:e�盛^Q/��6g��~�=CZCV)-��l�&���S����&yF�&u9��~8�2��������f�̀���%��-9/��{��\t!��W*ҽ�� ��Lu>֧��,�^�r���{��5��5T�0���,��r�v��-���kZ��q�t�%����W;�ۚ�~� ��5���pÀ��\ ��M*5X�'A�2��y�����$�˔� ��O�<sF�L��ݖaY�@	꙱@�'!��IU!Mϝ/t�s7�ù=G��e����|}��cO\wx���5������Hk�8D���`i��R�g����Mp���1�sG��|�0��r��X�/����g�D%�=���x� ��,~ιF4��3H�m��"?�l����z/7 ���q��>3�?G������
��'��jozŀ�9ٷ����0*ܯ�o����X�=�J����Q���Ø�'�3$z^'c>�gu��:-�A���!7��8k{�H&�m�VܞM��',.'
|��7b���9vawxh�y9��#R,�h���B���)����)4H�r�,�u��f��Ôwup5�D�/?a۬[P�Uj�3��*Nehf�7�RO5���@ӤJ)��	yO }�R��|�3/��L��R<��w�� Y6e�,��T�v�yqL����}�o�0@h�}!��^1AH����Kl(�OO�{�8c��#�C����%����O!��JZz!�F��+�=_�Nd@�5��A����6I�XGI�L
����I%")��f!c[7���@�r_�%jd��%�U^�����\Rܔ��
~�_����:uj���e�����Y���~ ��*%��t��f�󂠹���w�ձ6ڸ��t���[oe�J��.��p�l���SdP���b��*�|s.D�j�6��L0?�Q���zǆM�R���׭��a������>�vKU�L�m�:Z�h�䑮�x�5n�@%V�Y���YC+����ݎ�Qb|��+�[���&�*���.mE�54�낛FA/�I������pe�����4J31sm�kJG7�F~���L�5��z^�o' ������2�y��;I�jw���$ֶ��7&����DB�pW��"O=�-x*�d�e���H��XA��.=����ų��O�Ϋ�;�����̻yn6��ŉO�q��
��v�����v²NG�q/��5��(��6���NJm!�^e�s���TBd[5��$$��W�Ӆ停�-Q��P��T-�~��w�g/H��a���E�U�\�j�	!Hv���Hw!�c�l��x]N�����*ut�P\z��^�3���I�R&��Oɾ5��]B�=c�  Q	��L}�I ~%����~�D���ܿ�$�B��5^��wڒo�(?f]s��#A3M���Ta��V��K'�h�'U��i�T���'.��r��E�q�0��=a?L3�.7"�zH�u,��+>z�ᎢZ1)�i}��Ba����u��Cr��Y<��Ȁ��.>�,J>ON���]zu�:�{0FSzJ>)��� �CgU}�A<~�s��r�0�=�t��B��߳7�n�W�xW�'Z�<��i�|�Q�*F$�䀀½���!T��\uσ��/ HǸ=�s�F"�s����E����t���|�S�!U���h1
_���d~k�;�!���:�)q�(޴u���n$A��>�]Z�/�G�x��3UQ!Z����G�������:E�,[v�#���sm;=��ȅ���kg�\���R���g=�ۓ��2V�d��W\7tu#!S��;*;]0�*�;�诔�p��~d ϐ��ٴ&brg%'��%��yqBs6I��)
U?��噍=���'�o�4`JjP25���j����V&ŁX�t8�J����'�c��2����z�r�_��3��$g���ٱ�x�Ϫ�d�SM�E90I�vǈ�3��'z�o=|�v�x�Ocjz)HEYP%f"�`n�@�n��`k�L`��v��Q�V�ۂ�d�+��_�ܣ�8K���eE@yMSх&�Ǔ�v_ڿ�Ѕuٜ��
0�byl[�w�K4�V�A<�/��PIP��-B}S�JM�`d�:�I��/�t�S3A�is,�ٵsl�ՙ*<Q�@L��g(���'nE���a��IN�B��vL�X��g�0e��-��.�PU�9�I0�
�a�'w$H�i7�
]Xebsi�m&BUEP�wB��Ϯ^ ̧nr����7\<�~��%��,����Ȣ�َ�����N�zg��(?V2���4�%%*_�j1LF��;��";��<n"}�a5T%��x�Ԍ:�fL�#@Gx�����\�")D�� xT�ԥ*�#bi.80fK
!��B�G�)̜�kp$�?��4C�A2�@d��j�7L�����+᳐�X]L����b*@�,P9£M`oL���0�&�%�oJLY�ܽ��-V�_�s*hm��Ex���J��������#qn�]�cH��R́�?}�H������G0�;����^��}*)��D|��K.�?�HҒёI���v���F���F}���?w���1�	�A@����d��yȥ����/^�r�Pi����'����v�jg����ϛ	l����-��-�b|>��m�[�a��p��UJ�*'�U�ِg��z&��%��L��/����'�_�jm��� A@c�Q�-T|�*���\]��+E�~����qI�aO8�B�7�s:��Dѵ�g<5*��i��H����)��i�bg�5�c����`��p��$q��Io�}õ�>8JɈ��pBr�҅�7�5 !C �}&q.��$b��&�XΗ�5��3�߳p�)�u�`���G��D��~�� �1G�$+�l1�����+���_*K]*
��e��2Gb���Pw�����hCf������@@C���.��Wk��=Ez���J��'i���
�w!��ͩA~�	��vp!F�8=!;����0�o��v�pt6��0r��6�d�s�� ^�g�Y�ȁC�ؿ<;Ts�a�{�ze�(F��nד���7��������)q���S��T.���r-���s�کRF�2/ulF�ō��mB���푎K3����b^�SN"���|Hc+&{R�w~�m�y���ؐ>Y��L�:�o^������p��H9�c�����:P	��.1ji5��#��e� ]q@,�k)J���{�����r<�T�� :���DX��y)Q-8�m�ف��������u��Ѣ�qď"����I�.�U	ل2c����1;�1��_2wsv�N����Qi�U5T��!bD���05�}�F�zN&5ʚ/F'��McT��H�J%�+q�j�g�YO���Z��`8=��S�ߋY5L���'x=���-��+�&����4�OT���it��掛`&���}��͐Ħ��Fn�B��
Xr1;�N&^����"�f��T�^ lo�ܿ��[X��t>G���N��_m�$W+�a
n �`�
��A!;�1�������Y�I���],{cZ:	g*u��lڻkŦ�2��p�&�(dy���l�Kv�P��H�?�C�--T����w��q�=�����q�AH��2w�f@����4��#L��ShM���4�=�^2��O-�B���?�3���XH�ߢ�v���
l�@���@o#�M5"o�S����X;U+�t���!�Ow���f�{c�bV����;ׅ� ��(��5��|X��h�R܍�4ј{f�+��Q ^�'].�r��R�y�/g�������K�3