// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
yNItg+tJVvGRWBK13o9QkvWxAS3G/JHdDiz+GQDGO5NhjtnFo0CHQRUZSO1zg1xCi39Z2QITekkj
vDX2PTpNoWJM5kjrBU958Klad+/suqfibu/rDGmtuavW+CEaLwMEZavrK7kO1c20bgir1tyoXZ9P
RrYHSrBTc5+LSEYCGLzmeVr1GvvEwEq3DwAgRGOnACkt7BBMOXQsfTFxLVkibdilEJQ/1FziC2ee
t4rQ6xkUDBVE4I9XUimgB7hX/xHpYYAzIp0pLD1to4Ve/l9yWzN5sMWrI/7V41Y6lHrN2mx4jAg6
f1ePbrJNgTvuhrNWdPh7Zvv6Mr1iPTi/nWuU/Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
mzHcY+KxNsyzg4aWmXCW8ENpVCFVr6eqbKyJuCvvCYGw8zF2dGddd/GywrSssiWKBBY7oHDijR7D
VFeFGLWrJTtW2/a5ahAZd6E3MmtUDHeRi4bfa49iW3He8voypSWu42HOVNvLgaxvP3apsffuqQX6
mpkEL36AkGelb6OCeWkVTL6W8zzfirD0izY0Q4LqvxhIR4x5IcAA33bGgjlAB0UDV9gLWrd9txVi
CbsVAMrFbGQCX8MSR9lBWrqZnNfDF7g71r8cvmkuRgmGt868Jcpp+GW1JGJTygYAS2NKOskVur4e
pIvQGihkxaLTAgLJY4mKL2e7SMxFawhvU40+QEWaVxg2sIsrcJ8SnVuW4iWWqtJsSoRq/W+4Nrex
2Rd4WvSutA0jgiGsZI80mAepVvj806+TrK/9tsBXBEce4w+i8AYPPY+68O1S3NaSa6uV0c1Xkbpw
oR2qMQXR0HfouqgExXie9TzNY7EbtAVlPALJ5dPLEj7nxu4ApqYuTgKR1JNXU4x28zrpw4DfS7LZ
iT68Z2hPjVy+M2epYVsI3BHhUwkqb6QLfLGwsLOROCyKOeQ2S6QMPJ9KCdWuFU5+e0nY5s1G6qnl
2Qo0Eod3Cd/LZ1mYYoGmbi3XEsWNTWuRP9nw7rIouWK8S6xA0ULDESjk572diq2cHxCGBgpLb2Jd
zJ8j9rnlRm/6fZdzv+7zrEWJECpsaRv8pcqh1zjIg0Es4NRf5YKfCn5miWJqoTJGWOW8b1Jn8j0T
bIFZMhlYSyAHzxbgP8xo0FYpVooy9fuvB/Yyt2GS0456FBLFc2cQ2y2XrjhTk5ut9WX9VyhIhHvi
UePai2rlWOP8BeSLNep2wO5nEqymgFR4jcgCYAuHvISpHnmAA1GwhaqKZ3GTW+YeKb1fOF4Hew/b
svlKnrqDQHQTIH7M6Gp8/mUfFXHZ/nOupWW9OSLGEgT8fBfaqy687i5rV4+mf1Wi2qeyK672VOva
2+q0776cM03pdIHwNDJGmc6+apEs8y+MiUlg6TAVGmeAFxDlUdHPl7x5TBJmm94o7nHoKhntfQ+v
CNuKbivzniC/XFjZriyQ0skvmgo8a45evRyebKqYV1vXHGsuG1OciYBVw+FA2rudW+xGYjvGzKrj
ZK4fGgaPK9WHGaF9/U2k3nbzf+ckI6QARS5h0RRA3QsR8we2a8j6qOA+GGRgVcyNGvaKXMc7JTXW
GmhO1HeUyag+jq4zJJSDLoaERsOgLFPteipGNq3tYJnKVgFJ6Tg3qCBYJuufS7hvmXC5kW4ljHwy
/lJ94IscY2+OgSXPMTIt1acBo596LVbFMrnCQUJrpXWQBS1I5rukItIsEMObypVmp/sLF+T8/qvy
0WIU1ykzT6VORZXHkyMKXUvt81Ae9Jz6zJd8Y9LW9HY0ZwW0EQ9pP/doX1dJbdjDeRB498nkoC7y
mvw6SDMePEbzG2Q3deJ5+il3jxMI9drHo20GJjad74rviQ7zpvgYTA34lHzejfz3vqt+Tx2gCqhn
U2SbPEpCy/gurhLm3UdJpyY0n0351tNJW0vU1xe38QYi/AwKaZbTd5VQNj8Bz4Gp+sXrseOQ8gEw
eyJb3AMPm79JJGt3V8o7VQDUa1S4d5BagdWWft6RFTsyoHXTsOE/SAq8TygAmHzYtKTvLPTEeDgF
P9Rd3YoP5YpKCaQvLPb8l2bjnzUcm/8iBwJJxbjnMOdVKSjpphQG+kc0LdqXc3ASztxXeOSLou+v
fAIpOQeILLCXlzGMTOIx0Lwds+JTS8GIVD6l2/7bKjsjHF5iklGT0LJwFgiOMJNW6Jhg56lcZ4H1
RDkymhWfqTIXjxaY4IVNf+vbV584EYL27e//LfygkOyY9uuBzqIEs1AGKzczyEO7kIFTdGIh4Iwp
LpuWdnO6TtufPef4SUi2GWU4IbcvEhzL3meXIqYw0Qqlu9vaJAHp8zk5dNIHKiT7/usoMhkpqFQi
c1S7TPCbZVB3oLlGs6KKrljx4TwWdew9jFHDdKNbEEGRPolj7PlWcLi2qt9pIl6CU4FNyo/N9s4r
CUZMWODnqYPKbEtPlO2aEsflWOJXgjQqJ5clj4MBoG8AZxaYNYzsCQZj0tAJ0WpIvVDgGs+Rz0jm
71OR1KPHngPkJpBDAKUuijyzdwFXA+cNEy1uvEzLL8nnBf9Adpr4Cq/ty319ialkOm1tDjK5qliJ
rQrhhK5KkdNCfcOL4VlO168EU31uy7UZ4aBbLQV56IhsAZt72dE66VVdAWUqhMC0F8lWNVpCeTU+
fjP2+QPtNKXLXSHu+rHjW18/yZL2N2/ZtdvDrO8dLMQXzh2KxVLGvczgXRWycKBrP5bW81pSLlgF
cI1/yKcsGXKccmymvokjLipT0Jaa+YQbqkSFP2LjWcpi6Ia3iWWgwgWLT63p6pyERPG7CzoeCAzt
Mcoj9Om/wlInGJr6sAHDDGD7gvxLw/hoTHssUepAqqRvralmaatS5eqACZPAGzGVlMzX7qqZihPo
7YI/Q170Uy5ZuCpVUqH9iKvyefTTzhsLvFjQrnh7LwyJJS9hF8tIhUqiK2TxbMk6IKLsElutWxSg
OJ7jx6soOtve+FIC7aQvaOmEHUK0aQMW4u36pXo6JkJ4PVxvIQX1DFXKdU4uc28pCYUKjvPXVRyP
B8zGJSXEtd6VwpjY8pbgQBbxvV/HLeb/hLKbqEw7Ib/N/EPM97m8K7CmkzBcLk382JMDJrBl2v/+
flrwk6qA5jYjf/cBxvZvLnwtOMRdR0GtaNCTjYRUJuP6//n//b9hBl4nY7vx8X3FbOc7v09h3bo6
25oGEcy9me4uZk1tdT1dwyOJ+OPyo7vaf1BW4wOvBRC+Yt0Dz6b+1wNjrWLBMVaAEwmvxHnirOg5
xpuFC6QeEEIZRQf91d0/0Bd0xjd+IEKRuej8JCxpqbM602zSGxNEbKdm2415erxKKvwTvyXDgt5q
tTi0qh1+R/4DcCoHd54xxWOOBYD+IpJ0UHzd6KrYQnNiUiMuUbtAhCj+StaEYaoE00PhAMKoGKni
EVgX1fnc5CvfBDbYQavzYSVCzdObLOUSOeJWM7s6JTyWpF+3jjsIxUNjUYvXl9MiGehGGCc3d7M7
IQ33BijUQxhgBOGrPRp9UXSZ9ogfKfxiGN6qK1TQRIP9/Wk1xqQY6mOYAWLKULXYx5khyfY60y50
1H1ETxpvN1Mla5ohYVbWQ2RBaZqeKk2jnUc6k+8Jr8RKoD/ZXVEG0WUhFDXuymDhqUKYwbcG1Y/7
55387hvWaZldPrQU9ULPTfYWVh52CrkaqwEDnLcfTAAQzIuVEGKO5Zeqj4nP2j71NHde4XC39m3D
8JJ5Pn1c5sYYe6cdr8l4X3+Uhbk8G8XnO801TBGNMAaH9YwDomxBVe8SsvAjKwXBa15Di2o+uBUJ
rNZtkl7MgV8lXChhz6uIOk6spRnfOYOIbG0sbac1Aa6KKsN3q9DfuXrtAtNqQ8da8G0sY5+Mzy/B
q5suLbg4kJeU79OgLzS8mT0zOWMwuAKHw6/bOcItU1IV8ngJer9pKBoakhShQDYL+g6yTYjnkRsb
CPcagW621TskbiQjIiZTFXyLb7j8xSqtb3mTR5mnIcloDofGf8yLxfcFp4VJBLa0C6kWDsodBPDl
liyMYSikAd7CAnWhU8WY6PlS/g7GC0ioHcQxgfBYqnvPLvfrrS69yY44Rc4/QbH4mSoV1ce1BmAG
mCSaeEYCEVgjhzkix+Z+NAUBtDRJrvL497G2tX/CSmglufl4p7Uq7IpM6OTM3e8snwcWWVE9li7+
MKA2CcP2L/J2GPja9tUlI+dBB93KULtccIfJDz8+8El+XB9x8Vn7UtZ7w9iNW1TRQF6tN8LxvT2J
EzIoHHBMLx+cGmPMgOL9ohYn+RXsLIBHs/cclEXbYTh3GSAqBso/zv6n6KWbtdlm1XVFT0DBguh/
J5LgOfoxcoVif3u+rjRNVahYkcoh1CVdLQ9NMvk1Kvlhi7xSUAMFy/1hGYXT2w1MBJl/mMa3a/ji
d7+HOGvhCwBBF286R0GF+KSExlCytoKRjS8FMt+POoWyhkCa6naII0wr+PVzQouvw+we1wZzL/2g
spoOmje1Qvn75ERbJ2HNDwwAVO6EaPJQTreDDEHoMUqQq9tKrGW75HKT+ylWdngAyIyYuDOxYs6r
XCHNXqtNv+O3qXnKxms2Vfkphig9vDMcAQ4CYK+lWn4Kq1+hKgK+kpeXuUjcqHO7lkdTThbNAqU1
RU1+vSjkSGulCZhnDu2cdPkjrFdRP75U791u6C9Zm49Gu7ZD7j5phzl+jx0CpJL1FliYE4m72BXU
n+mtUerhnB8w3PI/Ux5j6HErUO7+X1/8S3enF29n3zTsq7g8qITuBJ8kB4dOnZLUv9pzHEmv4Itm
EG524F8igQGEPlyVDGuWcmYtWNhx66rHfo3sprYQDkQyRLeRqze10uEv22osLa2c19HNvrNIFW9R
aTnTfRGHT6+RCqXZns5zt/rPylxCSoyBfp0V23IHl3Xwcc7Z2IPRlbN/wwal+VGkUHb1/H6kd6ID
URCpX6gLkZFFsHEwFmm0QfZUUR79u2yJQvDYaZsbtbsPd/Mc1rbFaBjaLVq/Yh9ra6JMmC0ZwLfc
EujW44TBU071GdaG868eSRr17WPaQjbdK/NkSje8zaoNJVZ4Yx+WWq/ort5GIUKnNNio99ScjPMP
M4WQCZa7CZiWjaVtoTJqElGEZTBsV6Zs8MC8PJTqUwhVyHxTfZH34/JxWtqhQ4H93X+Z91IttaWC
sXOEhUNNOINlmXT1sfLtoGdmjyo+YQak/WKJvMPCp75PvdN9+5TgQYhq85QTLveyeGkUSKQNsJzS
numXv9XJ2Okr5J868PI8ImKs30rEwP8muRshSApAAh2IwpqhE9UGYDMjk+8nprNrsp2FElL0vjrM
P1rVjfQ/DiuatNKtOMzA4OZHl7HPnEUgj6BMetnN++6l4RwgU2b/mfIOePrYPPx6arthM5ChQAgt
sxE1/9hiUYNvImOjbH2AB6oy+BL7TtPE+5sDN4D2ZNor+tFdIllMdwgVZr2XOVGLhkFjEr8MU8Qp
zxAYnQfnxJt36hkHyx4EOHo0AxwyBm9ZVBu6BKs8kddP2Eq7jwy6YcFzcEuyPsbrJLJeVlq+Dxws
B8XluGE2X/bNYaXwD21MDXBQLnprzqFImGyyFZH0hSt4KxECPC7VDXa7MBvx5FqbMmDj1Ugbfs9c
34evhqO8iWY0ZvS4mxsXBOtmIdA0MSORD1NdJ0cxfDB256UAbdLio7NpOPk2djcWqGXxIsADM8uE
IF5Pc9kF0SIyAgOWj1IsV2oCwHFYnao9S5MJkp/uxBXYmvHkqBf3Zv6LZFq1cp0fcjiCcP8zFK3R
nbIARujEN/uWjOi6bKeJKKg4wME1jFVtNNx3L1O58XE6YdzZnuCgIs4OgRjM3EWapbiSFlWaN0zs
rvxxGoTKa8M1+PZf1Jk6lhYOGy8PGrFP2dBdnCXHUeJVvBm/DP0PBr8PSz4yEMdukEkesVZXtKs+
zEH9pEnMLBCsxf3SriF8MujMpWAZW/NScMdyTC9xthAy29UbH11Ud1sR2HWHEZa3Glej6CDl31mA
PSAwdkH4zQ7iBKX/ateFZSvlITA1lLoHFweFhPmxJTGDT1sqospjFLTCVsL3Iq/hJ8GRDebKW2jF
Goxt585N+YJQ4rKiTbA/ex8TunnDKLuShPtzYKCo6UH5yXAKxh+MLcqBkRu6FNKMukovq5pG7bBX
4qBeY8ixdDvA8xVDLX1Kem+0kUWz0cjykJqu94qvLVFZs/QmzHLJE0FGGfXUp1juUkwo/3MuHoHT
DJt3M4/rXq2dwI3M1hqdUS8YNFW4+KxmeVMOtiVh+cF6FNRI6Gmj8orb9gVHVolCJ3nveri3ZTow
Pj/x+i7jf5HD3S8mVowWbMymyQoh22/VlgRNOzpSm/+sOhmOh2HlInuxepaumii8/J7f+NmTw5oy
9pJihKbFHuxhluAldkXe2Wmk9MbE5KBRkXZ+Nv+x8GWVQnZRgqlgh8s2cwJ1786+w2OITpfi2Mfr
XwA6CUpQSMuVwX/Pgito4O0oVBp36eoXQFN1qLL/Slx3/ZlogzFsdOnEarSSquI/yuy84IcQFJlG
na4qGkNAAmdEBxZ7UcKgmJX5wUK+qKYkz8NZxG3VksV4vOZw130xoeMIyhvfrbJI3c2cZQwSCT+I
Rp+/y3BU2xnqxZWjOISuhpbsmb1qwv+mKHppi786+hPvoRBd0sIXg6LQD7SdwS23zDUV+t/d3lLj
ZcnOUaWe5gKH/F2Ewt0z6RNZ9k0qO0Esoc4s744VhS+mNVFM/v6Q3Oc5BYhnyHdoiiLfpbZUjaUv
clI0GAoq4rk3MIAeJqzTm5F7afUlc0dfDBiiyGPZrjLxO41PHh+s7U5TcjB1YkC32eReBwuxssSg
6tZQCLHpD1Rp8hoa5ALAMnohHr8nj0DH7zUyw28zntYAATAoFSr28H8QqiJj0EueeywodA3WyQSH
K5+wpjSCkQVTe6SsDZn/vpzKPeFj1FxgOF8f/OWaP2OUtbDQVeFP3y3gmL29d4bzclYLG6ua7QfY
Cj7HZyXis4NM3zyldzPdPziQDh9JNWcBF5Od8gmomQu4hWMghPdkQoLG0zRfoVXxaMTHftwsUgEU
3983ogkZLS4IDpURJFYrs+qSGQyLzFNxPrXz1W9+6/7PsMzKBOpdQckeA1NnqWLEBQ9/5yfyqz6U
a7RYeQ1fdjqf/BJwSAC5oq9tbUX3sXiHh4httEeSlVV+2+XUOLXqUqsyko/03eYO0VXXB7YTGrtO
uBJLc7dejozCaDl9C0yrRmDjZi6jBCt98+7502j5A03E0YNIZS31NPicGKLXe9tOVi9oz15tz8fp
26r6I1eqAX5IFhO+Gp7LoJ3qXxl7Ua0U2M95/LP1qjf7i38aWMTPPjXy12FYQJmNYbEgDN91t4hH
E4UxWBY+wloyHd+tdkrtunnFKj4n7muwhhBUGkeTzQeu7T3rN1iqn0+xYjNj8gWykRHClkUTeOSm
OMfjgpVHZ42NwxWlBw1YX6Wxxf8/RftAtQyt23RbSiPoe9b0RaMrPXNZ3j9L4VVb1zU3TPG2Nue9
r66Lj4jubvS0f2knJs2J2Mskmn9UjbmaAsNY99AAULmJ4hXznJJHqErAbyCDQHc+PN7C5w5qmn0n
xxXiYSchZDn6AruwKFRZ+M5Dfe4MbQRkMddHrRW/aM2wSvbuVFpnGqCqjUi6m4NJ4dn2U8mjsd5m
R7dRo1/MAxhE80F8MXudq24znqTo95KZ27FNij1dqOEvS65kVQ14AZybRFAmdrJgicqFCMN/xMv0
eowVuXga8235vq+zsRYbqljtaTaVt1ngA/hGKTVFI6u8cG8w32zmPLQQ85reWTwvQvhBt5JhMKSC
0wDJkijcPQK/rEzOFjjL3MxybQ7w0z24J1XTVBNV8bJyfoTpRNLXdKQkGslZ/rYfZh7rfwIWKCfs
BO8u5GxQtbxwxzlRfelDahgC1k/YfZ6DBeHDqehx8CXFoVlWAI2MGfkZwiuInVlrGC4jwS4XBf/e
R0wih2C/jlVf662v5CHbzSJahtN7NM/M9HmKbzpsL6YGdImvOYogPZsE8ZIgFZnKySkFGrCV2B6i
7fwIcrZw244qGDr0m6+1gLU194JKWwBRCIWwyGcg/XrmTQptIzwuZivBPMkiF2hfW8Hxt5+pb5bE
VaKOr9RYCDVsoZXpT33RVkTsyWC2fNTw0cIRzZsdKm0xAaXb7QhwvCIFR5jbHVtYGBIC9yVSMOZS
ByhydRiyyjP8EnUGQzRE7mmI7w2A/ALwioLkwuzGWkcPGDeorDK9FIRhZwM2mJ84aCgKy61y73+E
nv21tN3lYZTMy8rWid9xhHbJbfU/zRqZ2r56K43xBkcCbkT9cLNMLPpljx5pEw1zNe1EzRbaxdNt
R/HrjdsZ9vXReeJFD9d/HvH3PNVrSJU6I5hhyDrZ6OI7nzFp4BN76zKjSRTi9hLaJ6W/EPTbb4kT
Bn2+JIuhlp1CNuQvKUrmW2wuzWCh8tUgfhr+63IM68cOEBQtTN8Uw3oylsYUsHGczb3hJy342jek
7bz0NH9VIfjGpzeD0XoFsrcpNMJ8HxG5Tu7IwpK2Nz4H3+xGcG3cuMD6MuxdWloD9XArha4bdPB+
O5QE2WGbh5ckDyzn/yg3vgRj/1jL8Qzk0uSR3uKBDEhTmWCUa+NwsXGgdX5xM8yCF+gHc22glgxB
pHP/IuNws3U2hFCpKfIMmLrBUyajZY8EOT3cRWu2/CKq3urXQiyK3hu4vxpmUzskmw0CDIx+HDKe
zlYKs1v4YRzPvYUhajEXaHhRut+CsYL9OAAj/jHnb2CDgJvmdg3oOGdmgYW/4Y0S6QyZYM/MOZ43
7tmH1KAWTEn1GbR7WpeZHcJ9w3yZrWxTu4Yx/+dR5JF1oOC41hSCTtnhzwwNrHkhKGjaXkHbJvdT
i7nF4GNfgPWtQjda2HitgJF0fvVGs4GmGDadDOw3IxBLHwvsxPA9kwqrQPvpwDbtA52waYK9Mqk1
TSpgYZ/zl+xYVlKMlzFF27eOaioq9gZL6lwOSSxL6aFhBIvNvVM949gTxJhEKCJD/YISsCelOzdz
xFCc2trwsL3BCDSYaT/x2qterlWQPNsji9Ny6yJMejezD9aaiitNXJSl4Z2O74GSYTYDHzZyT8fy
BQfds9wBeeQa7QzJtvkM5ewFjQBKQYDApLK1K+xClc0YfQDURgpxlIybDlwGFnhWbpzqIMgnejhM
4PAwtOARHagUhWsqWphAbIljnU+1XGbFnEpfgWylxppF0hLRst45rJkFZl/SiTK6bz3QXPdbhZVk
OzRuPk/4LSjJxhIJaFe/bnW8zXAHU4thSCepVXbrH4NTUG5tqFgbwpRFERTrp/cSgELPzzRUOO+6
fM6EXbJdDdufVDRMIUxlzNy/+GpfZPbFxO4/oYpXM2nvic/HsxG8W3SYoX3bm34gz+JrubRjmKci
1qIbjDnPmWWmeRlRFRs1obDUKKDsv8v7if25jX2y7uaK6AJAxqaqSLcWSdqkGUjXg3aHD8IulArB
3UmfYVWgLLFOa1UFf7MM46F230YF8crW5oFykJzxFj3KCn8A+jpcFW6G6mAcdgErqX/DwsacJaQ8
2QRR7LBAyoTeXy0oBM1pGemAwfp171KUQXUbP1U9CfLdtpIKWtY4zlKM56u4sbu88anzxR377+iB
xVzQRZG4HgvP1HH7xxEoDdotIpFhzZPMr4w1jl7jucCBjIC+HM5dfPzm053IxQMgZQePf3374qqZ
GvCGAv90n3UKBRMuFhPYlyQQPpYf973UikqsiBJkSa0r/1wXzj2ZQiM9kgsPxrC4Wk7fE/IpAyUD
Jp5Oibb4uHjpOObq+bN5DP3v9CJj1HW+ykIsLVETycWa0MlYrd0eYtQvmwbHgckSLANFO22LpCmS
rf6IIucnJl4UhlFVhKsho239cUat6xagO4IBr11Zq1WujnhXrZKWEqVijhXw3mIY047vJk2UkbiT
3/T/QB1wwdbqRv8m6w8rbSvG3U01L4I3cqzdBEcSX0eYHtHkVwBtfktjkfIeQU3R/tpavkUM6CmI
qePJhTizskyQenOqYERibiF2pg5K6kuJ09lvGRbqvJZmS6vQ4uaWxO4WkZOmVj5rq6gPi/9NQxSv
yaO+/A86DiX3gcpEp4NETSbXEWZQeygprBDOX4iguzhhsgup5/3D83hJenEfjRb/6JJgDpzKg6V0
hpSkP6kdQppWbxNOFGsI5Ov/R9QBRvRJYnGYGicjwxXxVNKYTTIGl/2gM6YmOelwugMaIybpVz9t
9T4VYdAE3ylvoZhV7xe8EAt9x8jLGy729kvx3ruospdK1oceAZ0hIpskqOCu4ek/mYwFOng+1tiI
p9CKlTENFl0zENcywQJXuDVecw+43tVMYJIZl9Nbr8y0KjYFu0N+8HN3/VzagskQ0pfaeXFj+8rZ
HL8+7pNaBIlYIFJJQ7ZeNN1fcjT4W79anDnGrooKaSKHzEKDzabSRIkrAm5BVj0dvJxdDOhZ0PyC
NFlfP97UY+kBCeNl0sf8T52UsNVoinouCggDW/8DMlO3qslE+9TA3uNg0uG6+5BA1JsgMpcUDVbv
xqE+VV1b3FVgqaDiQklsmujDClGrmNXCMs2is0ZV0vMHRzPVjOZRnq+1X4PdFSB5prVsXWxAuG/T
od/cDLoMW+xSl1yR1r76Y42ccdF6El9C4gYhdHIDYviju8mZYDG4CqLmlxQuk7UUrvZNSBwiORtV
QF0/3qW2F3QvSxmx/lp+6xlNNtmnibGsSEu8k5WtaRYiGsVpz77jr+fQsqSg4Z2Sw7nuCTAGKgjz
HKzicupZ9CfkQD2c3yt1waVpKsq+rDu99QBEjwF/StHoTKJoMj8V8iCslFWUVcb49KCJAEYPy1E6
Zi5z8qu0eqIxuBFnKX13PHeoEQ7czxiomaSRA8TI9k+QyB/yuYuN6o96rlx+hGF5tAijNlHEQE8R
0Lh0QfuXyYloA/IK/3Rt4xIpmlXzlrr6+HzoY1W6vbhw+YnY2lTS2M+zDvmTHe8KxX14od5hzBcq
kqDxhi0001RhNmn8nPeVaCYFaZb7S3PgtMqwlX6EBdXWeCZFYVd/rZ0VzVY+H9X0feZw1gYgMEKC
Vkc5sqPIPnxXrRtjTmhLcHsBZSFP47EH8ogME6i/tbG+8sP8vDeIGurCykZ1bQnpV1JJqqpxySFI
Dbkv1wxJ1wY9zNj+1xqjHkToNJ23hjCMz6lP39KjMvyc4n1/mrBWjM+ABYDxRAxbcZ3SQquLRh9I
OlBHU0inOibV84o86Y5LXptOjaGRFLV6TQtzApx6z7ycwMRW7UdZ/CDXTj1qwNbByw1l89uNUaHN
TQudQGMMfycnaK/SJI1it9+h8APS4cJagJL7G5Hy0DsNnj5jxfqRjRd02jsudFSqbrsfeAfxQ7Zs
oY+ygg80XAquNS2HpczxCmOuZddZDTfCK4FhMPDlMvfET8VvYKbKSeer2o8wLI5uZVUrXuQoBiBC
M7uu0jPAUz4DQ9WEqr2ysQpp0kCcnZ/RfOa8a6WSE2iYKsXtDM+ifRg89LfpezwYUbQjIzFZ2Ibg
C04B/xfuClzLplxGEHudiAvaNAYrxXnvYz/WQWJQXuScbuFJ14p81uLr3W1gGDmam2P8gMGQPzE5
1ZHX8IcC5c6K9Ti7QarL2hCdYoaVzd8TKS4lS6mremtUTmMN9HhLHIKzE31kGOyfThUmgkeu4uZd
5iw8Hhqr+o9lR5kWUgXH/gXQ745FNpB3Jx1uacDMPo64T8gh5RWbI31/e08ZcdVX+S2SGBvBWVqQ
IGKkdjW4dfYzMzMEuO7yGGmX1u1LmkeXqS3SWvGQHRfHrmjoDsOIy1lK4BgkJah+TJ3DC0znwKBN
DVjA/dNS3guaZEGGNUT9asi9mIl5qrbGchzVks5lzQpDVpMzTGsgQ1cIJ/qGX1xRR3vzoqVBJ5sB
/VRiYvz4I9FKZzT7PmBACqLOfOEuApkU8XsJwueH0lx3kMnSEzRjwEmu3BG1y91wQtSs4O9Dd1Zq
FLy7fITzIH4uE4UPUa3oIHohrjbuntHqP6Y7XcAWTHpC4xx51AzoItv2GyU37Zn5pJhV1ngT6EUV
HWO+o8peWqMSfPK0Lpwq8kJK/SsortqgF0P7YBwtassr/D8t34iBxOqmQ2yBG15VJydjg6xmIAn9
jARKBpfFiFdNem/QrHtYGx0uzWZrnsPBCFG5aU3foPK9mf0FiW9s+YdRsuHxqGXNMXTb7py/X0DC
HO++hqpYyHV+07j6r48yzGD3KnGCU5dWxbY10pDLS47ay/D5h+WbXAblETKVT/hPozHoRHEpBIUq
IlLkuI2YwEPQvaG3TG8bVZFOiK5sGgpQCTfAMgTIsL8mv+Yy27bWX5TiL6+rTL5n+TTpmKxQsgz8
EXMPrdk5ggfRme9ZYONvv5ccpRMOIZNrCIFuG8dWOioNqD4+qBR8Mgil17lnz6W1H/2o98/rDx3y
YxoiQ6BHtCZX2qaBlpa52XWNxJZ6HNPFkp+6g292ctt6waCzmSRHGWmzMExXzTQCeeJLc0EsqkQl
uUIk2xaAj6cz72VkaBIcRnfke9SymyUK2tdUeR2oWfbJUns8YgIAjfAaWgzSzkrDmVYnFhDBr0+g
estS0DVTvpkU7ecG213i6vk9GYW2CqvITBW7c6c2Uc6S2MmKBVl/L9E51EOl8NQF7gpNZ4CwxGtf
QR3MyWrMhc2Rh+EYMK3lIRGFnEu8bRaVE2xC9IhVsjEKsgf0zUhu7m0mR0mtpRbc1/ES2xT1xp7x
E8VCuLs5D3EG7q+a9IMi4KE0gGSISCSU9G6gyhYwHR9NkO9YdylblU79sGxaH3piiDUQQaeP9MCn
SAM7CMLFCF2ypw4wOLTCVfnoL/pbB6lINMvlNLRDU0/3uKlkq1EsezZDJyo1vwuxe2OQQk41Fz7w
cD4jc/EmhRDqyX9e6l0Lo9G5gMWxXUL0AjRWF7t6SZJL8qS5OYFOwyMGYqzOE2fQHT86ShZofFbR
D0cq6Xhd2xkRRen0qtjufytrZLcSiIRmGc4luulYZJt88I3J/7oc/HTcnSDzfkEngygF4ePl9zXh
ekHdx19g81+p01+LnFaOjL1WAPtIivmI3LDv1b+GFTI56QUY3IY0bLEvWWoc49wTD6jZ8hMokVLb
H3W5oHmscxZwLF66GiIjrOVXSwE0xsqZyMGGA4Rljedb6W22oJkSblCrS934SWPUnm+EjKpn4hGd
G1mN5y//79zrOK4yi/o6C87r6wn8jBdQIrErEnrqbVC0mYBgYzmEGOVlbMWYvbwi/KL4M/iIpfRZ
4PODBObV3/uLexFlib07z4Abeu0FpRTfR1dnsDGoB3E3CHeyDkpwdqh8GHg9fUmRekLslTs/lr5+
kIkbYVkZ95jhoOyMmhpop3uMLDJLAbzqeVbDANEoruhmGmXOJqPnBoVMaNmUwajMLY7AA0h2Sdi+
dHg+R3tNifIlQT6CpoM8qj2wf+hxRf2S+gN1IJv3ueXKzKCrABZSDf1mEydmDxrVXQEzEyZUvzDq
OBkCZHmUezFZxyCxLXfI903sb+IOUSq9Z+jqLZDpwrcdvVPl7A0ny8txJ5NgpvhTjoKW2kKLZrkx
c6zlbxS/vQs6ISFVD7wFzQMEg+Bf3NBFhLryr+zD2GiZfOcARhCONB696s5oa1nmgfBUbpy6VgTf
6sWlTWaqEUnxg++Opvf3O1F59uUyapyBWO3RPE2uhI8353k6NbgcBk9Zez+NqRRuXRtZRsAUNZwQ
lEyvvse5Istr9gM6ziPsnT+/NajDKHW1LTzQNkgGjq4t7vS2HKgfGCFlr1gKfJ5esKyDPR8h2exX
iS2F9QjRCfYAx21Ev7rMfqahUx2409MDU8ayOoAPDPRxWiBSsUL4TAsD8eIydSJnys/bRo7mhGud
wRN2VcW48AigEzCde08UiNBjfXj7zxnkhhI8Ihkc5HRiIl+xCIxF+TqEgKk06TWd9hsJLEiPGwv8
GDPXE+6e1OUcST9P0cp3+bjxx3qcyO+Tsizqjm1j7oGvl9Dt9DXvcFGEpy0rf5rXSIArqk44XTWd
DUUbjHWsItR7xRwgsFN7qlHUGg3oHrXqBpF1PQ6w3CH+Yw57okweR7yn6nVwB6yCk1VrAIXhnLnW
lPF+i5np/p9ZnMYyp6R3c0zxfZhlFFVhWUtDRzeQDOKle5pGGIJ3pMqD+7SKHX90m7kinjbbT/T2
nv/Bt2L5ho/WhP9nvRn0c4ocgSBi0K/1FaShmwIyVvpN8zRej0J1uIntdppW+HNbY0ZweFwYfAUb
K2GqF16rZC9YOsSRkRY5MkHL8p8+8+02v0bHbMc2RGLGuN5W2PcVZxU3pGz5kijxOnSvIKTbfwsH
Rm3AAygYQAVNji7q4gMARZ55BU3lK+dNGU3pLzqsu5mSMqBSbywYE0Aa8wSKIrbPXrkAgXeJ9d87
nu9Pd9V5/7z3RhNGaGkCQ7oZ2SPRwq+s5PTGkD/iO8HSvPI4FiJULq4dI544h5wFuQkL3YKGcEkn
7l6oMJ6WHfwrCGLSOuR4q4fBDN9FFTv+/gLcEsjhqqGdD9EVchjn4JvO0aSuwSFZ7bmRLr2plAbU
DQFSdAh5X0AUf5iGPM9xQPAPteeZ0CKEqg7MHRypBjLHMOEIAvfpsWgv2BMeUpLsBRl1EklnvonI
ueXckjxmjJnwnjPmAnTTKwZqxMlUnFFPy6B4zB0PPknz8EG7ARmMRmegR0SvapTVjSXBoax3mlBw
VhoYwKrJE3r4ISwIw6GW4Er1BSv4NeTp3Q/62bW/QEdW57agrQ80wkh0bOBz/B5AYodZNzN2WM4i
TR0KmgR9X0qDoVbo/kbD+jXrzQZ2AbAYC6m+FMYy0JlNQ+R4JernwhjfeVMMyr56Q1PJDDSCmXfi
+iCx2446PNctGUDyerGH5Dk2imU5vpcxiv9XoB7aYTTlvwhfDETCtfUq3Wato/Jp/wh05kO/08ut
9h1SRt2aKXPNF+jaLq13rzbGqUKfpvdgMMq8BvjfRMZ3EFUakw52GyEYtIoKIxXL148Xt4kHEyDh
mCAUjP8v/Bp2Ct17+nKXWvbuJfMMDFxZQs1IZqfoQBO01G8DSPNi/hxsM0X6XCHvNG57uQsFB2nZ
r2B6KOpCM6sfgkfcuhy8H6/niUqMSZ1Drkt0Xs4onP034KMOO4IRTeNCFGduxv8OnhtXIEiJ7Mgd
4rscbGE=
`pragma protect end_protected
