��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒������O� KX��g5�tEQn����d�{I]ٸ�xuT�Z��H������i*�y���`~�wn�-�z~c6�썂=6�j���a)�y��k�yH.$k�ѵR����&lOF�뾪� ^�x��dE��3m�������`��B-隃�-%i�MQ�f)9씰t����y-?�5�@
�t௰�_��U,�m``͔�\�s
|#�1��&��aq!��$�Ae��Rn�����18��rc�����z���%ӟ������֡��d��bV�?�%F��p�e��TrY�~RR�&"y �^(�p̥#xA9�Ff�Y�簏������~��󈙬.<��Y�i��-G�2�6Ǣ�1����	>���/��ڔ��������A�J�6����,�E�����#s�jjJ']L'�j�̧E�����@1w'�[Q;%�s�-�Ѿ!�� ��<�@_6K�15}-L�Z�:7T��o +C�H,��vK^���{���_�eI8�����W*�X�;�	kV���eZ��ar/c�R�L�Q����}y
�67�O{��W�v�O=��A��y����[�J��p�l]����J��Խ�#�L:��#"�^Ԧ�*��4��h��+�H/7���.�/�@���g(P��J%�?[q�w�X�d�m ��M�����e;'T�ľ��Y�`�.3N�����-�1 ��c_h��mY�쑱TG�:X�塱$���t��h�h$V&��Y�.���`�5�~�i�3H{��� WIZ������n﮶�����B�&���4�B�{a�C m[��9�D����J�	X��kҸ�b���'"`c[�<?�QYt+�����ʞ����L�BxL7M��5�e�ˁ�y�ⓋQ�i����TΎKφ����l�o��@�sб����ǉ�������1��#�Iy�p����Ճ,+�v(#n�Bҟ��lP�!n[�k]�蜴�������m��@��Bf~��<�&�x���	ӛ��4	J�7^�+�"x�C�ɟV�k�W��o�Dx΂��V�;|R�޽8�r��|."�*�E��ji��"�`mR.�|�)<Qm]����kn��[��p��^p��'���2,t�1���ϝ\ �p+�	�NZ���`�H������j�^��VS��ܽ�-[< �P�iF�D��g�Vd8�}̧!B٬GJ;�,tΊ���l���C�^@j��^��\�]�d;�.;tac�W�C`��;����!z��&�o�j-03�+��Z��`TlL,�UBo�G���8E	�k'3H۠h�YFu�F7��pM3�7��ՉY�e�mm?�9	
�H"<Rr�Vڨ��Y���)�+nV'��▎u���:�_�h�Cp�ڼaң�!��6n��d��[�;��3��i
t�Æh�*(`�{�H��!�����ުg�����#�帴\�� tn�`��p�t�PiM�}n��6n�&�/���E[L�C�Ů|�p���W!�5㱒	���V�8j��:`P[F��"v�'5�b�h�Ύ>	^�G�ݰ������enDÎ�
?�5�J>��D��0�L�Ѻ�nm�j*��İF�O2�2p��/���zHn���]�k�;��xM!~Jz!��[�w�J��B��m_s�5�w��i���u���Onk����ź���^�/K� �,��Tq<��Q�[%�`� LS���F5�W�Tc��� �K�t �����YdL��!6��>@��	�ۮ�߯�[͐��nFػR�ǹH3\�e���DT�gj��E��gٚ������_$��e��3
 xKv����>+���y���fB������)��?n���*�:������'<��|�i�-�����%�b�P[n��r��,xrt��?^��#7;����Ԥ���s���1��E;�Km�xZ�Pf[c�.#M(џ�{ĎLaˆ��ݳ�3u;;wZ��9�����al��b%ѣ#-ì>q�>�ė��'=��D�0n�k�����z�O�^�,|`^��m��w��h@2۰�Y���5��L� k.u�Д�A%��$��i��X3�jtҎ���K���8Dh�wiL乯�Y��Kw�!�~�Px��N�D��\f����W�" �t�
Ɂ�2�ym/`>�F�V7�"uho������X��v�ukY���e�P*
�#�ם�F6�D3�ǒ�Fu�Fm��LTg��p`q:���/Ǎ�q��ɒ�6�XA�~�.қ�׫,���	�K��8��S΄7�/�b&vg���g�T��+g��8���K�3r�(B��_�r�$�G	�9�c85%䭲c+�.�C'��\��1m����+��-j���p�u���	�,���F���u���>��ge1��nCk��(�ƴB�r)�|�����>��=�A���i����z� -���ʸ�e�f�׼�}��Z{�9��iq���vmچ'�¥X"Qw8R�}� #��Ai�Ng��Z�M|��	��Kp��ĭ�F��q-L�!�(;E�0�m*P���4RICG8�Ϋ�Gb (��A�3�O�'ч����i�x�d3#f�m�$~�G%ܖ�>h!rs��	\�{à�c��ވCҪ/�Wř(֨�ܕ��Ȧ�����9�|���< 
cX�Q����^���,�f�`|au�Yl�Ҵ��Z���x��)�!́�`��ݕ�k�7���4����m���Ƚ���(g_܂[��D@'���y����Y�8�<UE�b9�7����$M���S�݃�����B�6���f��.���R=9�ı�n��s�ν��w���Y3X�s�/]9ʹk{��ߔ~D����$L}�t�@a9��`�=�8�A���u��)݄����>�"Ng9�ˡ>��(�b4�^]�I5�H9�ݙXGlM�4Z�=(��c��#k:��=�o`�c^�̅��z����&%�W���9�7�U��j�KL^��q�U*@3�Ϗ�G���R��o���y,��������2G�Yi����'Q���ʂ3�4'AO�f�~�{Rke����!A����ת�3.=$�&Y�S�ֹ��U����~.����*�H�3ީ�p����n���T��[c�q9+���m������3=��A��t.�&�6��?f�!�p9�������?�W�����L����n�J�����?���J��i�8�V?��҂�I�������l�0�����zP�]R��|/��_�r��GH�pճH!eKK��lvO�p�j��m�5y���c©�Q��(H���Y]'Yf*�0M��CC���$����A/j:T����L5F���c��Q����X%o>E0�܂c�a��F��P^C� J��:��T(��&^��6ղ��V?g�C���ن�R�U��=`���m�8��^m,H���*f)���J�����%z�_�)����Vb(�U*�Y�N�TNy�O|��z�4d2m`)��da���P�X�Gvp&3$����&V���K�K�/�'_��bv;"^��#Aqf�5��U�6:Ԅ���\}�˷�	��%M�E��5�w��[�� ]_�ÕW�x���ǋh�m�6*K��AI2�����D4d�/E,�V�\��^]X�,O�ol��9��fda6��j$����'"��)�*�z<x^T��y�B�D6�B�����52N�3H���ٍ���Jڃ־�edy�J���ݩ: =�?G���8�ӵ�׍m��Y):��]]oH���f9�d*���X��\l�I��%��T�^�(@���#b��Y��m�xF�.�P.G�S�c(�n}����+�8h�;���4��.�m�s�j�˧���Nl"b��E,x��Rڐ�=/�}�*'�[�R�M����E����5ڴY�S�| �#�(%�����aΈ���$6p����	��d����#���~�92�U�Pj���P���~�m)��b-i$F�떅[��iݐU�P�JVO_&�w*j��Q��!Ʊ������ıD]74|B$�ְ��b���L4�V0q`��� �ћ��VD�Ƹ��|L���m�&�Sԥ��xy��l�,Z��	[!Dᥤir*���� "�&[���I^�l�̌ܛq���a,2��a�/9��>�Wغ��fV�k�څE��y׷��N�]U�YY��N���/n����p�k� � ��eN_b�z���Fw��Қ/TF�4͹9��˘��I[�/e9����-&�?sZ��f�����r�UY����]�x�D��֤��c g�2��4�<H�隰(k��l>UY���YY����Y$Ŝ��v�A3��u��؁�>�^��F5ڬ��j��ʴ�]|vD����P����$�M���Hѩha׋�b�4���k�O�Ax���!���5)DO�b|�K�^do��~�nvo����n�Y6�xe�J�L��&��F�v�q'gMt��D�'�k���n{:��2|����׵�ב��|�{�2f��S��F3X'&�� ����h���&���N咱22�s4������"jC2���*�pZ���#�r�'�"��u�<���;uǃ8�E��H?:۾�9f4n��)��|%��E#./��c���[$�
�
W�FJX�mP��*��z����d���t�k�=cm`σ�wsy�,�]�����_j`��f��=D�e�p��+�P�~U��	��iPA#4�n���ޔ���jC�$ �TƈO=�.?p�����@�z�<+� P+amۣ��VT:�{�H8�+M��#;�'�A
�^�g�}�A1T]0�J��̚�.�a���oy5<+�`x)xkٛ_ ޻ha����d^��YЧ���gr��� J�Ag8ӿ���%le�>�4e��X�s�5ޭ�$�0�<·]m��J8g����+�)�R!5;�l~��JT˒HV�����������w�M��U��� )*Xz�L��&��|�,��)u���/���p�^}�|	���os5��}�H�&�tF�*]��q.|N}?�s"G6��������T4�L���^���F��c�?Y�g<��(�OʎL�3F������HO�<.R&Ē߆ ��=Uh�3�.�3g�6r�V��?C��tSG2�Z;�3WD�ۥ�@��/.c���'�w��{���9���2�`њ�) ��]����s�	ZF^���9�*�$@ѧ�1��P�w�J�:8��%VE*Y�q或��ɿqaE��}u���W�1�����L�b�:X�}�h�ws�{z�n���~��B�{�O��^YX^"�������#���Q�PCL�J��q��$#a�$x�tMd"*�.ЌPL�������C���"��� ��{�8�q��t���ER���v��`<za�
�FV��d㐅�������Ur<߮��b����d�; ��0,����K�Bk��U�����CH���l��^F4'�$J�p��O�v����ִpڡ�A�b�ف
9�/J��= B�r �\ğ�
`��nB���O���<�<^����_�'�٤�G<:,��j�V8B��ka���Zm-$��^x}��$�&�O�P��jИ�J���Μ����0UJ��xe�_*Q-O����)(�|oJӹZg&�j���[�&ڦ�� &O8T��?=�e��5�3��n�8������\t��Y��Z`u��#�����,_��nt�5�y��Rv�RDy����\D�r�k����<p���a�$��8�s��',2�b ��	~Y���㛴��)�K��������}��j3�eb(���G�����c�>���E厊![�C-?� �a�Ԇz1V�5^�sa���$�FY�\2���D��o>��u(h�<0�C�ǧ�7��j�aA�ȶE=|��Z(���N��u���ˎ��`�W�	N]�yjQ#I�lTM\�7V�"ǍXFJM=���	�2��'�ݫ��+5^[��ċ��y�Yit�i(������B�|%�Z���߉��"�^�nS��GC@�i�	�dI�=/ ]TvX�x˶��r����Eќ>͜�bd�����%G���%�x�'Y<$��]���rj�/��9���B�|q>V��ت.�`�M�lv��B��p�U�!!�a�@�_X |v���1U!\e\i�S9!��7_�0Vٚ�Y;,��%�Z����CG��Qd�F�l5@@�-��f{xǔ|Lhz������'�/��}0��l�]fK���\ �ȵ��;US���zp<��]�H��g�cSU��K��������L�6��o��^��E�I���;��}+�%�
��o��+�V��9�7asPG���m>JK�U1}�_��b�f�2ʟ+�I��%]H��}.0��	#mWY��'�8y�-�;H�5����xc���7�I
�9a��%H���Iw�1�"��>7�m��en��/'{���k*D��dG������Eѹ�GǺj_��%�u��qK�h�~ϧ�Jou �-�E5yy�<>;��1��>Ѽ���O�q�N�EuA�H��]t���z&Gg�&�Z��l1.1�����Љ�-3nR�2i��)w��}P��P��r�{ܶ	��} �u�� �~���j����`;ĳ/	F� ��*�O�5E�
+E�ps�1�2��w�|o |����[���+��k���FA֟�P
�l�C)��"((AkUm���!ͽb�L������ĭ���g�s�����!1�[12_�XH1�!���=���T��z�f�q�J@�X��	��!�^�(�Z���Ud�4;�P�py��Gj�
>����-K2%����'V���Z�Jp��&টZ}�a�}u4�`�dsپT��M�4'���F��,�a��~�]���K��`�¶�bv��jA~Cr�(�A�q���F'P�rቢJKxt�Z<N���_��:eK�t�Ľ�� $IPą,��������XM��E0K���a�FOH��uo=�wh���8����`�0��(ǔ&�Ae=���G��{��ɽoG�';���ߠ��yy�{c�΋%��!ih��F�Q�H7=�:�CV&�B::1�x�ݡ
�)�� B4���[ބF�ڥ.Tl�̡�X?���D
݂x�����A��k
Q.�����5}�w�m��VShMq!y�-Z�@��ƾ��!��R��ݬ'?����c�<���
�}3� �k��43�.3۩�H�'����hw\�^��kWǈ�}����q��Q�XN*ղ�c����Zj�$�qH3�]�Am����%��{:�����N����G=���l��(�y8�>�"���v��V���ll�4����T� ��z1�{˱�a�2��BH~)>���$�fD���E���?���0<�A&����7�i`�	���^-��U���K���#�yQ<��ؽk���5+�,��
3?���K6P�4N�}2G�e���`1�+��� ���j�L~ODN%W8�Kb�R��I�F�#��X -㨄�@Xֿ/6��F��M��/��v*�_��f�d�R���#-�	z�:��v�b�@3��
�؏5�a�Hi��=�ى��&w������?�2���m��^$}���s�A
�^<7 /pq�G���W
�PNbPQ��n�kI^1~[U�T��LQ�+�Hu��]/���s��� ��
��/��xX�I��m�?gu��0c����{.� z>OaxSc�/�\Rh!`�k3�s�K1�n��-�-�͙Ql6w�|�љ
��v����<�dK��E)�xZ���NF��b-FzUĸ��(D�9=�|*��!�"2�ۻ]��7,RY��f�oDŸj�K[�0e��֫(m}� �����-\�q�n8�`�9�w9b�u�$�1��+�h�7#��uV��q�TC���č l>WP�Yp��;�`{�%'d���(fz=��'������`�����M�pl��bR��� ����wo�Ib��`5)�2;#�� c:@�R����8�󘲕��w� W|�@���J4Ϫh����#dy��Lh��xb�uC���.�9��s�9���lA52��&g>f�T)���l����ɰ�t�������S�Sٴ�Zܑ�k�x�*Y����4gI����3�t8���U�.�8��=���>��@{~_d{�1_I0CԺ�y�V�}oUj<��J��]!���e �6X�s��.tih�1�z/��Br5�h\Y^�}f�ʨƮ�&�93�/����@Z)ϦҒMe�R�*s#Z��?���e�~��|Ƕ�W*&���Y��۩�>Q6��eGoF04 w���v�0Lx�f纉�Cb?��)��V�@UY�D =�������"F3A��Ġ��[P���(��[Ao�4��p\�F}�۬�NW����J����I��ej8�]0��j�?a�5k��]̼�L�T k!���G����\�����6�D���t@���F�?�)��X���*��G�v_~�,�V�|��!�j�r��'�.�NS�c(Kq�>,3��\�@6,3�]�� ���W��N}g	�3��n����`cݽ/;D�n�l��������X �V�R��N�21���&BBC�~U���}�E~�r��W$�3�J�%�ڥ�L�,��x�c��G~��Dt�PX@:�U���:�A�H�#t�$���6K�Q��j�0�6I?�;h��I��#�m�J0Ҝ�Y��fd��*����&H�ur�Z�!$��	D�4���f����W�2{�п�%��t�G&�6��ý['��zA����B���Y��u]w%�<�7��2ZH��@����@�f(��W�ŵbm��Z�Kԯ¯�U���):	,�s�K�cc�*��V����<���L';���!P	�h�]:sŬ���1^�t�^~����H?��o�{������#�
-�Z��F�*���C��OtR��zD-'�b��,u�	"'��O.a\L��xMPa�� �	D���~W����h�� {��d��μU�h���w)�|�V!�-��)!m�;�������ڄ/��1$�������v}�ƌ_����|�]Қ)EG��������e~T��&��4-��$Ω�w\��,�u��}��+9Z�㑟0d�4�wX;c4$A�g)gV2K���y6)7���.F��R\�C�7��YP��ʙǸG�W��R�|u{�<�����q?�T�U�u���[@�Q/Ko��HC<#��D��"{�����0���˦L�[�/^���
a=��(����G��mݚ����a5�'2��$��hv��UeA	+��Ty�F'ۇ�h���P����}��XO��z){�-<9�A�3�"�"��|<��b�����D?L�K�/�/QS	�F��$��b��R��L���r��X��и�PY����=�MC:��Bï(�TI��
�q�n�ў��Ʋq��@e3���Gz��q}�D}�sxv4	-M�M�x�9�P�u�\��ck�T��y㞈+��$-wNZA�v�B45�:����[F��ÝҊr�+R�S�o݉��SW���	�lc�l�Na��A �'�躖�wLGSY�S�ܕٯ�S����������L��������%�L�u|��1{�
Z�N��u�����S3NOd#�-�x
��M�������-sS�%#i��8s����J�~�t��_��覨e �	�Q�U܂���q/��k�4	����Qo�w"�ܝ�qV�kv��u�|�a�X��	��0��)f]ص*U�\�:-M�
�E)��G�nR+�/�F��<��ϥ��@+���9!S���QRmA��g���[3j1ڊ�LA�X���8�u��,m#�h�q�C��k�n�2�
P71�|XD�[{w���ɜK�?ž�8a��Z�*d��yHaq��i�1��rnq9�-�#�0�?��rP.1���1QqB�s���F5��16o�;�����:17�Z��2b���:պE��e����ݛEd4y��p)磘S��'1�H�nUY���>����Yc�f�S�@Ȝx��H{Z�������$�횽�*�nz~K2�]A�GI�\�z}��s��+6��Ns/�ȝ�!soj�Qg� �9_ ���+SX�3�o���v^4EG�^!���E�а|o��ƕ�.J����t��o��#~��PoP �
�,�ѣ$���Sc�`*|�/��L��2�\?3	s���N���d =��M���8]S�w�'g�@CY)d��gA���#�jF��E��O�C\��≰�s����M��֙�Sd6JZ��k�55�]3�uQR��v�6ȭ;(!8`<����)�����;������`w�����geg��mf?�� ��ƖW�
�Z8�:=�@jN��AE 	��ּl���`��c�A��4��f��@ku����$=:�{a�:�g�bP83�}���x��Yh��m��Y�*%)���y��Z�n�Yk mL�%&ێ>�I��u�\j�Љ���!H��F���^������Bp=>�Jb��mr�p,5��Ƒ[�F��|��+����C~y�W[�T����G}����a;ʃ53�X|�t��\��<t�h�~�S?�Z����D���ƿ?����zvC�VZN��'Bz��[>���6�%�̭^�u�4��K3�pe}��%��4�T��Ʌ����nv"�B�fZ=�r �3�b������'ٿ6��`*��I6�
�B��gNɆ)dN�o�Q$�6̬�l��Bg,#�1��nzU	6��hS�`��1�`*,�ŸxAē�|��0��~I��!�xm�Nupar��9��T��H�+#��cY�Į}aG��s �lg} f��TY�K M�K.�I|��Zƍ3=�>�E��Ϯ��P�9���Y��N�T������$�;���>!���~!?��h����	�K-��@o�H����DZ�3�!Yks��,�O�+z�d�f�����*F6ce�|��j]�Y辈�o7����X�n�ec�8	񼔳~����D�����|��K�����,0���g]�N���wO����_�"<`�UWFZ=ћJս3��Mu-��^B\#~�1�:ё��^�x���(j_��>����I��)�H�t����ƚ>�d:�ࡏ�|��>ԩ�vZ�M|F�����|��U����,}���A<� J�Mi7�C�� @w��GeF�Tq�D�$�2"!8�R���<_\n�ZG�nA��BW{�P��3WB6fTF��$X~��J��9w*V��q*� x����C9ˏ�a��]�U�t�}1�}��gL&Z,C�����&��'�*��+v�n�)�,�	#����h+G�/��e���#���YUz�M�PR#N�Mw���$/6<����j:'{�>.�%Q���������74�Q�1��p�Y��T;�� ���.�?1����Yn$�E9��F{iFp���u�3�{�Sl+;=:���;�ʹ��j�\����^�G�����Ί�s,���^4U0�U���w|,pJmِ퐖����1��e����"�4�^n��MʯxI��;(	Ж�_~;�#R_���Qo
�8�D�)Q��s*MTD��YH���T1S��2������ـ�M`�����J��YJ�F�Sgd���K+Dz,�I.d���w!�`�E���_�^���R]`<>:��+�*����rxqP����"�4��IE��K��h@�f���p����s;{����PȬ�O��C��N��Y(hlO�PZ@ʄC�}���Xj�:�mkn�c3�ßĵKM"�4zp��G	���!腦{�a��� ��ț�b��&�)_�K�.�; �/Aվ'LQ�5��Q?�F��¸H�,dh�Œ4 �_�'_ru�R&�u4�F\�Lc#21~H�{D���Ц� �&F�k?����BV��1ct���5a�m�@U!�,��~A�O*�ѩ*Mbn4I�s�"_�x73��3 B
p_��i����X�<J���7C�����,WR�C�s�>&-���\�*W�Ͱ����O*����`�����A�>�c{�_��8�:�+W�#EBǠC	5bS�,7��1/�H�E-��4/�[�Gr�wh*'�G�t������wO�,٦��C�
D?�4����=��?��̴�����m'^I��l�5��N�0�J�Z<I�;�A|h���]�	����6$1�U85M�$��z� ��%�f�;z�LNÄ�f���I�Q@�j�pN�>)7�?P�y@TO��X��O�U��r:>�L�k����J\�4HY%9��6N���)�O���&���Ӊ7M,u^�k���8.AʏY)IDn�-]:�W�G�<.��>����#���Ti 3_K�I�{��/v	�K��Fe/���B33�oeX�C^�㌋"d��Jؓ��E��lE�P\�3"F�_���ȉ�0��b�w�!�����4�~&Aaǰ�����1<�?����0��f��c'PE�;�XCaѮ϶���Dh|�e�Vk��B�,�I��"�y��\�H��ˠ��Y����Ppg]��4h8�|m��;#c��ecBb�����'wA�/��'�]d�8�����=I��0�ީ���߶\�~I����R���JTܧ��y�Y ʷ�8��U�sۦ�opK��Ë�wqetm�kRY,">ʶPD$���=�m�c���9ċ]�ig��L9���>��=)'KP�x�$��&9߫�ǻ��s���{���l�0�w�:�s�\�chF�u�����wG���5|� 
>�2Y,�p��"�ιYL��)�����2���5	OTwr��ά�~��_����琊%�4��=Y�r���E����7��{��z[F�oX�*S�9�6��R�*��i�B�Ģ�enC>�E��өn�2y̋~)���W����MI�|�lϲ*/�q�� b�4}��s�~d��Б��(�'\�0b�1�g��cLJ]�5���'�]gNEϕ�U.�Xl4�%I����.��)|�,��܊�*��L�q�G1B�s��W�2�7ZF�g��B>���=�~���b�Ĳp�<1��$:J0$��"�m��a%Ug����#I���f��1�ڏ
��+���-��8�S�ލ S>}c&w�G!�:�0}�_��Ð
Т�7f垼'p+�������ҷ��0c���D�\���gr.�"�+�.�IV�.�Ri6D���=�ߵ�Ė���{z�n`5@4���h�DR��~��{(e�x���;��_ɯM�mT�#K"�Q�ζ~��避懛J�
+�� X��j����ϳ�5�yF>Q����7E�}"t:k}��i�P�~y1�8�î�Fg���eZv>jD���2>��',��O�����pg1����۰EhM�h�������宠��Q��'�G� �jK���T�(�{J_A-2���^�J�B�=�7Jk$� �����vQ�cLF�;v����fA�;W���F����l�$ۋ��v� )�%�����{lڻ��;�d�p5�ѯ�H�wjt��߃f�]���(	�0q'�H�kAI�ș?�{(��F��tQ�i�f`�������s��΅�)XЛ�}���Q�Ъ��|��X�AO,?cMB@`��ϣDMX���r�EVW�E����D�%9߿��+\���ѓć�����ȳ�Aj:��i|�ؼbq�t��8��<n�Vٵ��^cR�sch����5�o�
�����*CP��lŶ��f�=����l��αwTq��t&ځ�>J�5�&1ۗ}F[a:]HT���� �G(�ks�O�k��!W�b�
�e.T�h��t�e��6����L]��^�Rl��͔��/9���6���}{|��}>��>�����+��q@�:<�$;�ʭݮ�d%V�OfR=ZQ�}�#�Ad����Bj6�`S�h-{e��W�g�Y�R�!�t �Z4���,yd7O������ڿ��{�-�c�����Z�]΢0�!ņ����zQ�`XQں�����CP#w�g冄l+hT_�"��S��&U�Z�u���k���ڊ�X�j�6E%��k�ݶ��6C�_ۯ8���C��,�qt�r���%5�y��κ<�1����އ���ά{����6�i�x��@^8{9Z�]����#���aN_c�&?���t�#��y閗�ֿ4�?xڏ��]{%f���jߣ�U�܀ہ��+��bE$�����&&�^�~�����ֺp5�t<ӌkf:�S�>�̱��"�M�A�]�$5짶P$�"�:a ?G�rhӇd���߳��z���RH��<k#̓�l��]qN�P|
��������4��)�P�r���*"����R�����7�!"���,=fV!?��Ɇ�K�
(�G��?��*��騇8Xs$L:Fq�G��8pK�v]� ��]���(�zRA��8yPF�`���nyY�5���2�8\5�v�����}�˽*�����XH嘦��/�<���!��Ł��T|�p��l������<��ןqF ړC�@v�G81Z�F��Y����C������?Z�{Ȝz|�<�6�n�(W&��DY�uI�K�2$Ej<G�>���Izp~�WUa0�yZ��>>�(<��3䄎J�*���Pt-�k�z|�Y��*$}CI��������{'4�"���R#�j0�y:y(J{x�NƝj�.ű���&��[��O0��Ҫ������Ke�K�[��&L�VHtQ`�8�+i�@|�Lּ�R4�D�Q��N9R����p�_��M"�B�9K��Kt����iN4�o�P��/�ǧ�wXN�H��p(��I�
&���v�A����C��|���H�c�'/�|�ESn���a���k��\R��2�7/k}�&93D*k�����a�=3�9�y��b��@��\�͙Dߺ?I.�p"ܭ���d�*4��d��g�4!6e�ΔqJd"�-�z9�h��� ?��ϡJ�h]c�Y-_?�Q�M�~�OZu��Gz0��Ě�'X�@�T�CLo�'"w��Kɓ��i%6$��x�bB�\��O���[T��up�GP��v�Lu��� ��v 561�_8 ݄����3�:d~������+;����'j����Ă70�����9o��n�x��$N�� ���oF��'(t���ئ/���3D�o2T�=y0��Oq�Ga�gT�S�M!�wC|�g�6K��4�ly6|��$Jf�6�UH�L�����H�$�H;��NJ�=M�^֑E�8JE��}��,6Z�@��=���ٓ �_��"Pjt��y��� |gID
])^��rc�"%RA�Z��û��76�cۍB���;��+��*�똌�[u��7/��C�T�D�x�`��*
0���NDBl�=E�ކ��H� (k5iy6>�O�
�RM���cT���<����t���Ks{xMNzyM����O]�Z�&���s��e�jO��!T約�I�a/IYՓ��}h^R��]K��A=�aE %�x�*m�	~���`D�&�OZ�xWõ/w��r��\�0c�v��C��]%������l{G.f����'���w��q�ﭥH���!�J��|�{Q�-���5���W�g�K�C�n����F�F��h+�a�VMs��:��7�ْ��-p�T�qz�!Kl\�?Ll$Ӿ����o�/u�S��ŏ/��Q]Z���}�?��m����D=���|;�8PNl���Qm��V��>���BNA����Tj�J[�G�"�΂d�0ȥ=C�cH"�e�`�Hb��v
l5N����f��^�=YL���<\��ܭ�ܐq�ϳ�B��IY�w����͊��G�\/���֒gk�W��;���q�fu�_:he��k�>�7��������١���+ܚ�w�����K�Џ\�ђ��;F��	} &��H+^W��E�T5��M��R�a�_i�uE�O9��� )���˪����*/�B��F�yɖ���HDX�o�Kq�X�������� � ��@�?����7A��~H	Y9�{9��l���-R��x@�\�OE��qI.�YO�^�RP���W=2��-�{ET��c$��ZH��#����S�)*��Y=�7[�o�/���pO��R{�\r���*xͬ=���d�f}\|����Q�d\�r`y|�ݸm����-=�Yy�<��Z��/�x�*< ~_~H��3-4᯿[��}gd5Y��]�D$�pS�ϔ�߁���pŰQ��Y"u@�O��I�/b��eV/`�7L�_��@���	]u�K�Q�#d���>�Ŀ�K����Ɇ���Ά�[� �J�h��k�3�>A�ך6N�7�����䦖�/Z������լ��
��D��@�F�9K�����j�&r�k@u�#��������4���)�%0���"^1��}�fĀ�4BtO�~�o(ٱ�WLj�9�w=h��� a-���S*Q:^?��`����qJ��Q(E,�c��-+�:�&���M�L�O�V��µ��Y,��V�����X��'*#��鯧��|��v� ��ՌZv^S�ǂ���vp&�]�W��@�|{�"���{"���h7
kD����`u�
����"d�ϩ��Luǫ	�k���%�@ۚ�%fn(������o�y�/V�����c�������G_��G&�N�9�N2��`��T�m_B6tZ{c�!�@k)]f�/Wd�A�֥�³�iH��(�	��,H9�#,��WA`���?��&���J"�������ٹ?�2��dI����
��T�[w�:BԹ�T��-y�^�.3��B�Xq0f��GV�������W���S���R3�H��� �(PX�׈J=�I�Nm ��J�����_�"U�?����~(�&���{e���!�΀����:Ox�H�DIf/��/m�璌���k�OQ#�c=��/��sTY��IC���n��p�p�`���>�F���)�Ȥ�,����qȇ^�|�����U�e��qlNA)\wEWT(iPu%����w���_�P2�&!
tz%��9�5���U�"n�� �c��N0G����n�!$�9s�؅'����]M�WC��o^ʹ:�ʆ�K��Az�{�j�9��!������kL�"����0���7w��)�eQT"\&�� i�f1��KM1���`��Pڎ�c�BAӦR=џ��nJ�^��)2ɩ������JU�H��ь�6��0� _�Q6� �J�����N1į ��j�jU�$����DNjΆA�js�#?�����MY�/-�y��q��R}�p�J��=�-��r7�</�*9KͰ>Bs.�t�*��1K�b�c=�Kf�f9I4�R��;�z|N��/ehUZ�X�g�G�
(o�X��OW�@��2�XCF4)�#���+a�v��of�c�23�A�o������%��.i�KX��ҷ~�d��W�S/�@���s �Rr�v����[�n+��LkQ�H��u%��{v��E9!V��o�&��兂�������! ��Z�a��xl�t�t8F�_%��R)b�ԃ�,]�&�D zB{8���#�!H�N��v��O(n�B���,m�V��W���/ $���flx&8q��G�D��z��a�h@iV�t�Sܛ�̫ �S3�it�rK��A���rc�s�y�����G|z��\Y�ͮQ��.+�EI�g��(ӂr�a����B@sC�݄��U2�^%�TC⢬{t?��j��9�s�Br�)���@ 
��)��Wڸ�/p |����*��ݰӿ�=���þ����HD���c�Gǹ��_w�H6�{��2Z��AwE8X��.�O;��.�, t㣩�;#V4R0Ƞ�E�j�s�N�o.b�J�8��->��,V�!xz0���y���Ix�]����t�(�K��{V_�9_���R��eu[���f���K9\P���ތ�Ă��6Ő�tk��֭�F4tsD@ /��F�ƽ����j���O�&B��&�+�q�KR�������ІL)�i��ñ�0�}�fu5���
�f��}$v1�8u�Q�ɀ���C�%L���0�N�\a��W�?��e2�9��Ӥ�KtfԢ|��
 |�
�4L�������Lu���J��X�C��I�<�|$��I)T��7��AO0l}ɟUQÀM��T�@��D�"��'��Y��Pmr-���@�\3���%�h�m�ur��v�a�"�V��1���r�a͓.v�g���θ�5�/9�$?p*���~e+$��ѱ��&��	細�ҨH��UR����E�T�p�.���~�������������8����g]���M��@�;v~3�{a���Y7�)�3=e7�r��F�f�H��& �gdt���H�.�d,�.�Q;6kć��pV;$��"2�x}-F����Ӱ��dǚ֟cе��[)�ےL0ҝ�w^ճi���?= ���q�\����1<p�l9_�5�b��9�e�����dץ�ڥ�AN|���/