��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��[J���#��//��b?>�o9�T"灿|h�|��@nŌTu�L�ղ�4�B6���}���� z>�sWE�q('	aD��n��V���jG�g�#��'��s~�x�Kf��:80�Gk�P �2�y3�ª}��`e]齄qj�Y� �ގS7��ZI��r<�
Sd/����,W�m����'�C��ռ`h�����g��>A����v�z]�P�m��T&mpW�	��?_����ҁ�e"nD�����I'��T��'��j6�=�Ǟm�A�rT��~�A�U�k��<�a>��'0n�֏Y�@mB�Hg/�7""�<�j�ܻT��|�`Ь�%�[��"s�x��"e"zd�J	�,����A�2b�����+s��Ќo��ye�wt�"C�0��m�}<��o	��!i�rŮ�\"���u������:��$E̐b�eWCd�$oa�W���$�
c�?�6ɳ�N��*HP9r����O��w�jh��8Y4<���sy8`�"a���`�Z��6Uo����=������ߤp�\�8�~#��oi�l���eO�z��~P	q�G���ދ������6�1>t��"]�A�ߋ�Hv����sJ�:yMdJ���+�bž������^y<��,^�$�J%:�}�SB'uh�ɸ�_AT�-D�F2�PVF�IF�&�+�KX��U���f�l">/vx$�Y3�x�8�P`��#��LO9x����QI�]����<��E{�&:Xlvˆɨ��[
GXK��l��p��5�i�UE��������ᜠ9<R��yl�oy����$�ñ@3��EP�c�n�]P���o����B�Ml��O��;����9J�'�ank!�������l�.�b���t�k^>�+U|/&�:�w�U�S�����U0=C�<A�@_a���8����Z�H������`��J�5�Z�#m1!6�X�p}�GF�	E��q|2lo�������Q��=	���i��n��������8��B�����n�a\5�f?h���.�0�S+?��ot�`�ȩ���F�2:�e�����c~f	���� ��,�l�J.jq��r#uU
��j�a� LIځ��%[�8����̸�ɵ�~�)�[�[6ڌ�%lg{��L4�]o�����h������ָ��� �ɺ-kWÎ1���o����� ��N	��_E9��V׹ҐՂ�G(��I�V�mM$G  9�8���ilT�?�i3����V�L�n��(ML{m e������e.�����Tƒ�h 3�8���^<��q���:E��_=�s�GKn�IY�179Ȣ�|��r�H,�^�녡;��8��N��3�U6T|������8�r��L�Z��p����R�W������p�ڼ��Z��K9n��LN�@8�θ1(*�b����ľ��=�N��^���:~����uif�st�P�;��b��AK�"Q�^������Ԩ�Ey;��D���0QR%���λ��K�B�l=1slR���^#��ԉ�B<}�.�)��J�$-Q���}��j�% �d)�Y��/w��@����lo�̓��X&��h����ē��v�sE �%^y+uR}s���B��#u�E��M�����>�t��_�mQM��+��^Y��n�������$1�_�Q�t�$����G]�'�� ��r����w��ewƽ�'⻞E��D΀��
�{�����^�eB��o����L�X���Ë1�3��WyK�a�S`_gI9u��i�i��Ҽ3>fu�V���JH����`���Am	ʴAa�t�.|��k�/G����Zv'��fe�'�ī��#��Y�-�
�e��XLXqt٧�iA��M�OJL��rA!d3;��L2�l@���f�?YĿ36:9���#�e�">k�Y�R�=o�������]J�,�E�4���-*�~ǐB�2��\~��K���ܑ�aL׈�Ջ�a³\�F-��K�|dT_UL�9U	��M��W73�\���㬧�.�Z�jғWZ~؏�߃}�b_�w��g�O� ���^�q���)��K�צ�ף��3D���S���q�eh�'Q����}j�����Y�������G�ܤ��x�r�͝j��W-�P�o����w�__M�wP��/��q�X�Fy���҉���cf�Q����m=��9���xӒe3�����1��	W�����f�>yq�uo+<k�����Op�?c��g����X��w�U,�v�T薵s���"(����������'˳��-;��s������<�x�L�@g!���15C�NgĖ4t=�e�4BC$�G�4q�.�2��l�P$5�ɔ5��׵.���򖅼_��(�J�x��BrԬwU=$H$��2��Dc���ڃ����1��Y��`�o��W�M�{��xǥf����1-�`�a��)��	�[�_�ݼߗ2���3�O�{�����%����(8�(g�Bp��Ds�3c���m`[����M8L�|7�\��3�vj��>f��#.V�g^�~mĶq���g�Jv/a���".�%�K����R�Q,�?+W���$*�����4s$/�2�i��[�3���UQ������v��k���T�I�~<��j�FW��1n��f��F�Je�
�H|o�6\��}@�s��Xv��k h��"��]�O����=?�$ԛ7(6}	�+.Un�ꔜ��o�(���<e3Z�y"�lݡvH��<#֓dϕ=�ī#�Y�����=J�w�^4I�sfuq�fV]@��AT�����YGt�ZXtz��U���b9;��父�k�A�D�K��~��_oD=_۫5�}�֌�j��FJ���!��*��j;[}��m����z!�/,:U�S�_hf��usաʑ��d���L����g��UE�'���������V�Ҟ�qd�۱��$Z[H�w��5��ad�*x��M(b)U����aX�
�����,�b�yIp��}��ǌi�t{�r�s'�Յ �x�h�뭉�@���%�9�3p��s�����Y�ц)�Xx
�3C����}ٻ0�e�V�	Y�����X�1	��Ct��.�U`�R5��uմ�A����A��O Ҁ���,�������W�X:\v�J����sk瑕���$q��+����8d��)�T��d���3�ε{���Z��0NkbJ���W�0��OmN�hp������?4� �|�4"����2h>~'U6���.�Xi+?��!���S}e�Hp�7�U3�Cg��e|��|<ٶ���\:g���mXmP=����O�}oF��2cV��dVz�ҷ�T��+\,��scb�j��-�f��E��b@j���[O@�����UM��ɓ�\��.h��{B\N	�A��楠c�ڀ�'`&rT�VC�)<@ V��F3�%�~7�dX'�/�{㛎��3�4ؗ����A�L�I�@8����0��u?������$�Y�6�<L
�l58�sb���TIG"�Ӂ��7���0	�_��$\��Q�j�O ��lq��	�����<���ä6���@&��G�5B<���N܂׃O6��l����C՘:%�ԎDΗ�*������v7<��鸊�_<>�v;�Um�F����܂��8,.�E{����D�*��rG�Y�N�E�Y���{�*�"���:`�,/�����p��nj2��Sl��Qn /gtHPÏ{4�f߈�q(!��ݺ���.�u���j����e)����"!�e�/�ܣ�-$�#nϧ����R���r�����*:�mL�����z��Z\�]��A6̀"K�8�*'A0���7c5���10�~ �[֚�g5�T��x�M\@�Q��Rɗu��kܐn������5��D^̌��_������(c�W���+s����-��?����
�\PC�j
�k�!�g��"[��I}��4�;KzY4���SA�~�a����=�m�%Z�򆵋�� ^P͡�"P��`L9�Ę_����{��jH	��2r?��!�zK̩۪�0�I��P�|-��#�]�}��#�%���f	�&�$��߭>���~�n-��ME�v�W��T��C��XeP�mk�;�?�eK����X��� ��+�o�tw?��@�i�Å�g_9����#쌨��*�mz}��H��C�E�ſ_ �l�G̓�y�o�+�Q����K��C���#'��w~Ұ5A�8z%�59I~�],8yXaS�]�:5�O���֊?�4�����i��O @3�w��o^6��:;I{$JKwa4@������ �I���5�=}����P���(�9�ݮlø�Lw�dm�'cxn�xӂ*I�Ҿ 㛛ǯ����xhie�*��\�����=�� ��b������c�aY�����A"���?hP"� �U��K��Do����v5Ӥm��/��}��4��Ҹ��dl���9���U�Xtp���KD��.�Ӂ��|�p�C�)��"\\��Hr٩Q"���PM����S�)�Z.�p�)ri� �I���/��U��
�!��V#."�n	s��<�מ8m�vm$'�נr�0����V�3����Y��3�^^�-a�*R!i�	��p'Em�e�d��M�G�&]�S������|*Zt�m�����66Z�M�����ٺ��9K�V������A���UX*S��0LV��.��z�����5�D��RkU�u1L��GZ�	�֧,Z6dS��=��Rr���x��,�*b/��y =?������$i)KI`�0ցR\Pv�
�.Uu�}�$Gr5������&;ݡX��e�W�y�2��p�l�6�\Q_����p���U$~���!
����b_f�39EB���'t�Ɖ���[װ���u�ӊ�9�=�B�2.� �K0��D�5[Fo��ܻ{S����tY�p�:?��:�Z�:ĿUjC���$�C�4�K��\c!HAԓ[d����#D�F�T��!����/����c^8ZJb�J��Hn�
���U���蘥�C�)��jh-u(z�|ڞfr7�0�C�Y����C;4�A�Z�z��6E�� ����Qp�5%&��Dz��Zry�/���*�H��5EW�	��pleY*`�ʬ���>�R��iA�����;�����vŨ}�đ=8Eg����~5?�a M��!}�Oλ�¼Y}�B�,{Z;+O��2\ 61�J�ԇf��[,�7PV��N �����cr0�k��7�	�&������W����!�E�jM��Ħ��U	�(9�O0��ᐗ��=��4�s���;�`���5��j� �)�;��Vs��R_G���e���x��Т�Ĕ�B��ȭQ�?4��B�r��K|�'��c��Jv����ej*�&a}���HJ�7�`�$�S�� 9Q�|�d V�$��D�������rVp���t��ib�/*���7,N�B�;V�(_v��Ȇ=J�4���Odm�~SX=Ϸ�W/�?_�;ڢ����7��Gk����׺I����.��N�9��E�RD7������Z	p�,�i�ۉ�X������`��I�D��b����nn}���l�ޡ9���{���Q�ѡC�E�ѹ�/��%1�a����	샯� [�W�hn��)�HK֬������}bU�}Ҝ��K/�Y�B���fp�ΘZ'&��3b��k&`@�<.�P�Z����W � Y�������uC�\�`�.)�at��R�4���"��~5��[�$B�:������AO�~M]�C���Vǐ�!XNըB�6���z<\s��@R�G�����������6�}Q�Ћ��+�,v*0v	������@���JoJE⇣:jZ��Tf�+��})���xO$7Y�7��>�L�4��aU\nH�p�kvU���PJ��	DF�ܺ|�=�j^�1_(^��i���4�q���sr�����5������� ��N�;�[�3#������A]�ۦc�u�.&���?8?A�B{ �@>w��w�$���1�����b�=@���]��? n��Q3�d}'$�J���C��rS�ݕA%)&W��q��>8��PN�%!3�SZ�<H���E�����d
�O�I�@؇1}7���G�Dq?��P|]����.a���
��� �B�J(���UZ�����d�<�Ilg�P�2�?e���ʤ�T�w3j	ldŊT�*C6Z9��H��ok����|��c	rT�!����Kv~�xm�N��L�!�O��{�؋xP����9��yNd�>7��o:�	 We��^z��]	����a�z,N���.�!5p���mq��S��.�,��ۨ�E��-����%[��)�t�k�S�A��:�	@�
��K���M�*ޏ�?�-U������ϼ��e�J0=�<��V�ՖomM�^`cє昵�|��⽻�
5��l/���K�,��WU "�J3[¦W��������c�Q�z�Ϙ'����J=���}���
7�.)T��P%ʓ�+�M=\0�*E��a9
�/������ ��Q.φ�?�F*N�7J���ȗ]$"=�U�P{�%6��k�5h0D�s�t!5>�G�I�2�;(]<M��z$R�٣)ݞט�F�b��:[V��VK�
�9�Y͇�zm�d�Ԩ���-�A3LZ��7�?>�N�v;財��B���WDQ���e�(1��-}��;�Rf��6|�h��׆��I��w���.�l�+�v�Ѕ�UΧ�Ѭ?�	04�?��6V
/n�K_�]ã���Y���ޥ��fRCNWi��A�	|�B�@��"٨QdE� e��$th�{@�+ZO��8IK����ca7���<>�S��C��U������+�c��{^f/��т�*���X��k���S�f�z�2��LO�K�;��̆�="��C6��v�<��r�D�,b��UCt��]����|���Z�Er���`+�u��d�N�J%|�Ńp�B�_�HR��qL�<nQ��R�mw�̛f.�Ę@��r k��R���3��;�x�A�@2��9�f9��mQf'�V.�Źe�=���P���n9�Y.i�Fp2���6'	|D+��6c��
����w�4�1Hz�z�`]Ux��
��WX�7m��g�܋���%-��85n��C��<rU��m���%K9�#$u��CV$�H��R�#��+:* 
��D��R�U�8����^��SЩN'�����4�����Τj��zR�28&�O:�@A�m]���j[����!ӏn��=\󙑿���5(X�����`�1��T�%����M~p�P�|�t_/8���RF�|P�#�����6�]���~8�~�6���׬k�
�n������
��wK�vF~JD�K�
�oa}��l�^P�Oԓ1�q��������TTRV�������|t��K?�^Bh"�/e��<5Z*��(GTfN��z՟c�s9.Lj�Q���s���Tw����<��$������G|����^��=���a!Dk.#S�-��#w�����,0�[F�&2�V}�GdV,�}�f뛈�tFLM,7
�|'z/jLvhO\��;I�.�Y��x�ț��M���ٖ1\�QBP�bfB�E�pV�s��\��i��������<4�9`�Ot&�S��]}��eL��o�h:�����%ޮ|jj➴4u�~@Ƭ����'|�W��l��&��i+?�e��!13B�X��W_�Ġ�C���@:��NN�R����n��[6�+�v���v~v�}l��a���rYK(��BX���̡;ߒ*��)�0l{6��?iNP�JF)� ����(����<u�N>�H���R��s՛��^R�u�[m�tm/�H�FM� |���x�l�^�	�LO7�NQ�N	�i�"VUޭnv]1h��-]��x��P�Xᣮ���/'�8ۆ�x���7���ꑗZ����gh��U�D��#�JY$�[�N�4ag�P��u��Sd�������\��?�( |�D�o�ZyS_s>��ڭ ���ˠ3_M�cT��P���;�H��B��"1�ĕ��ڶ�(uS�a\���_�#�����_m���~uG!�P�b�����
�2��)˄�	�y�R�a����R+l"����(K��slm�^*]F������A�Aز[��������Ȍ��1B=/��QM�C�E�K�����h� �)��s��E�*دo��盚�
��_
�/1��E'	ÄW�I�O�����~��M�n-v�1/-�/�t0���)��O^3�1��hg�'��E�j��NʣlHA��Ʈ �����75;���R]��-"h>�C���E(���R�L��$/�%�)�=��G<�N�=�/�5*��>@br����S��t�l@9���[�.\ى�_���+�a)W�pٙML�-GV���-�8�;MֽC���ph�H��������D{��'1��%p����% N�'I+aoqR)��>���O�r2Z4F�"b���n�{����c'���!����<��h���@q
���q���J���~w�B��u��:b�CaTk�v�Z��Z��]�����L~cS� _��>���N�.4��A{xu�n����˅�V����p�;P>C�t�L�+=����P�0��A�5��G:��#&�Q�\��(��P��]{u����0Wy���� b�oc���R�N��퐀_�)�hˡ�Z������ƫ@�V�f5?�l��4I<��B�Oҋ��+�ip��_KD�ڶU���+ꗕ���&k��)7�i�
�p$^�c�8�6�W�U>�p�z�9P�A!�)���xIg��X������1�qnJ8��Q���9t��Bj&h�ER���G�Л3����{�����o�PJ���&��,��a�� ���&�p*�>�/utS_Ķ�_In���a�)w�0Ak��)�B���zlLP1��hۂ!����t��C��x��
!�+б�1KvI��w��F/����5��A��e��8�,���n�P�`_ah��ct�� s�ts��.�Lĭ�OHk��H�LZ6i�����
>։�o��E.Y!���2�d��j�j��w���U_�����������	�����6�lGS�#�g�Ԉ�u����V�uZb<�N��МD����כ��_��Q�F?�����=2ey�.$&���{�E� �y��gsLT,�-�3`�6e#���0'�Z��c>Y���D�4ҏ�p��Z���$0fE��2_����Ɓ/iy��|T�݃Μ�>�N�aE���Z4��7cc	��QH�qh�A�sbտDi��h�7��9�?P`����`�(�Bt�t�a;G���:��Pp�dx�,G!Yp���^��np�:^�J0"M%vX0c���G��F닗a���w���.	����I�q�_V�"e���@������KȨ��=S�p�~���1W^*�9|`Uile;�J������Q��M��2��C��Sgh����'蓆��k��zv:-k1��R��G1�S�����@�7�é��w�x�F��U�p�M%�sg�,U��&����	t8��$��K�@�U�M��+���RN��N��L�����H��3���,��֒1�12y
��·S�+S�cC%(t�aT⺚LO��Q�ܴ�io b�Jx�(��(a�r�ݟ+ݎ�M�K*��$>d�$ai,��3%aͨ�8R;�2�UU<�K���v"��/�oQ�A���z����D��u\|�������n��7��#cM��"n�l�R�f��4��Vf=��y���P��^�6�w)c���Ð�}',�������W����e����p�3K���N.Ly���!�e	�S@B���/�����~n��2�V�S���~5�[�up��(}�!+�D���:q�8�Hu0N6O�)P����= IVW��^W������ 3s�t�tL���̎2U����vk��IB����e�@��ֿ�q��>J�!V�ےV�?.5��d��90$��)�gR��tf����5�����GB^��LUxz16Οl*��΢����˩�)L�RH�u^���`��$X��H�V��=��.�xG�Dkm�U#��t���+i�j�ր���肝��Ͼ�	h�����)�2���4� �yH�G������Ox����Y�C��N�=��u1�|����/l�1����F[Z#���"�����55�XK�ou�gH��'~ �.�_*	ZX�(��KAݎ��
{}�M��B{NG���6Z����v��!=���}�f1����m;�RZ s0qǍ�],Cp0��D�Mf���d��i>^q�ɛ����8�4���KFY��uS����0[Y���E|���MS>�/҅��3�}W�~��)N��d�����OH!~�\e0sV4FS0a�۫��M��������l-*xO�X��7�,�:g ��HP%�ލZ[UMe�3��KW��)܅&U�̓��U�/��h��d���Mk{�[
���LK��3$F-�M*��MC/8������������>%k�@�^F��Ȏ�5����z�~�Ĺ$��㎜��N�<��*4���q�x^��f���wO5�1�1���� <--FI��M�H��M���r��K����WHޝĖ�������AO��L?�d�32��16HTFn)��ӻ�VN�Է��p#׌V���U�0�',��N�/m#�;�D�
,��,��[�#5��|���y���k<Fh���J	�Ǣ���pGb��2�Jk�+]oF'�:�����g�Y1!/i�/EC���x��W� �&'U�:�#����@x���c	r��$�y��E�o'}6����y�I!�U��D��8iʷ�F�OMVn�L�惼����-��d(�w`n������!	8Ђ��1%���8O�J+�����Vֿ�Ϥy�����w�df����.��x��D�'�]��Da\�0�B`���'č��Vk0��Cq��93 �Z��`l�&�;N���$�~eJsx��X'����=K�PK{�U�Je���w���VY�&�=��Q�+5��r)V/K�Bَ$ҙ�C|�" bח1��5<1�wc��,�tgd|��]�Xh���ܖ�a?2f�O�$LY�"-[q��1Z+�/�3��@����������8g�JkK��]��[���ֻ�#;#�wW+%� �#%O)�G���X�pz�_D5��L`|�S�6R�D��L�8wʢl�93ӵ'��T*��f�Pc�L}�C����í��?A� F��{
�$�i�(�Ѽb�N>�+��_�Û����C�É��ǐ5�ô��z4LB�g��V�?N�0�P
`u�߶��(�֮��X��-���������=��j���:{�p����	E��Y<�x3���,���BЗ��c8m�77�ĵ���C!VC
p�ϲ�����4%(Cz*�i%|�D�<�|��wї�ݕvM0�	k8[m�
�mYԸ�Kyv�q�^Pʠk���+��c.��x�Y�#y�ޫ��!L�6�sTc�w���v:}U~4Uv5�,+Ṟ���A�l��t����$%g�ݺr�Iˌ�zq��@x'}�n���c,��jܖc��ө��b��A�}k�ƍ3��y���
��@W�(Ʀu�?�EJ���TZ�ڳ��|���VNE�#���@o��u��(����-���1������n��嗃��/R�jf���%�˂���^`�=%�ln�����/�g��C��t;j��g���I9�R�c	�ܯ��p�,�����8e��)eܩDj�3/�	�����e��_��K|8�$vpF��?aЉ�� 6����7d��K��m�]�d�����齿�TdYh���5�@��`�-:���%#C�CS+E�#*�B?��h+�Z�4�мn��>�X��ffyص�O�)���|�R=pH�ӥ��/��U8��`u)2��$tR}n�#R�1��߄���.����*Y�\fd:��f�V^�y[?%S]�.3�͛߶�V�'H����6��&���4q1����,h��+7b����:"$�Uu=�2',��]33���0�����_�`��M%,.N�irSƕ����W@�Fh��韲�s��^[y՜�q���H10��-P��vq�y���y1��u��bK�����}?fQh����{eZzDG�N�pM#����HˁV�������X�,v>�Z����ԨG���ك��td�_Me��g�}�&rH(f���p��>����H݊���%U����l�T�����
s�1�,���^��B���q���8�G�5�K�;pԗUj ��r�mB��r�k�M�l����0N�`�Ȣ�To�m�9�Df�hC,GJ�� ���n�aU��[wMZ۠�c*ި��N�4̬�-0i;�@�@�{F
ˇC��,v�����|KQOB�����~���y�f�� &����n�&������/�&hxI��d�@��U���ϟ��鱰J�b�[6�?F,+�"*Ͳ��0�x����/�RY`�V�ʚ�{��1(M[�����8a��}.
>�����F����	�r�v�NG�%<@��Y�ȑ����$|��͑���m�s����
�j��z���F�Z-4a�y��l��jZ�S�78wb�-�7��{�#kPR*�A���'�>�>B�o`��0rm�9�!_�qH��i����$E�6�GB	p��뭭1�Cb��	�V9<����6���,`+�X�	Ϸ�'&s��D�X���de�
ѐ.(X�|?�3Z��, �D���э��,���\����:��;�bNS��&M�]��>���z��ՙ�W
L��n�}�m�7��ڈ��)�sN�k��	04�LBJôMH{</w�i��c�Y��2�d{�|����+����w�1=�g��j���Tm����j���|�6�4c�!��.JMt�}�nK?'@��+��1U����|5A`�����L��bf�;)���d�jo�G݊[&�7>WO&��J���Hv���"A9cb�25���,���b�*��o�$�����&�x�3�K����3��_�M�co��טg�r��R��~f���T�w�E�A��&	(��~��q��Z|@��.�;�	�&hR�[��H����g�$l[���etD��O0��+>�HlbX@Ư6F�m��m�q��㻑�ۛ����Q�F�`bkݤJUY*�� '��q�N	��N�ĩ|���s'��5���x/�7�3ި��w*�Z �҇h&����'�cl)�W�4�7�Pc�xXy����1$'9~�-�u�6`�܋�ּ≈��������5r��|?�a�������^G�i�"���?��T��ua>ħ�w���8�\�VU �Q���.�{>�*�@��a����sܞl�C��eU!C�R	Q�l��%��̴��� �@XB�D��fr -��$������`��v��
`�.�����h��������$d����mj��B5K+��,�N۬�}ÞPG�t&�;p&Y?�q�v!u�SdEC�"H�ˍ�ki��T���H����H���Z����i�Pc�[lA�O|��\�����S�x����fbe5�g���^#j4`l���0��`x�J
�W<,,��e=��3�#B���S@�w�/~v��~f�/�S�UM���1�ǌ��m��>�0���*M��u�F����A�����O6������R0b�$�bC���4!,�������(����W��zu�8nꯙ����x!I���,Wv/ud�We��kmRfѥI��II?�5��Q,]Tg�}�����I�ר0	` �?-|1�N;HC_XQGmD8�Gf(�Wg��������!⒑	�1������#����sk���͊\�� d�R���c%]�A�`|�qͽB�ic<Q���%�g�g��mK��m�?6�ݤy����F��2f����{���Rx!xn@�Z��}���ǲ4<��g �����K���*`��(���Fb�ĭs<�����Ksx%\TK���Ş�<��rB����r�R���'���D��R�ݙ�Z����PR&���ctE��e*qi��E �,pq�r`k�^�n�(��IB�Yd��U�v��H����+l�*U�U4���W������ %��.���(�聤����͢���m#���	LU�K珫��e��x�D�Ķ�F=��t��}�5ԏw����,j�&�1��g/������pd�"P笵9F��Ζ�p[%��KD0����a�7�D�m�lLb���ϔ�ņ~�C�<��U6)�fW���"���ن��k/��C�^i��h���`��rH�,GE}��L�{�o�8�ݷ�vJ>8���VֆmJ�Q��X۰�@Gc���B߄LG�7>堝?r��(ƞH8_�$��Ю��}i�1��R�ǳ����� ��]��W���OhI���9Z�=�<P����X��J�Ԡ���=I��^c� B�L�ac3n���bs{��u�n25�/��O+�"�Z����5F4=Q��I�>!�k��?�P[G��U"�̗n��G���FOC��e�������ݻE�� �%b:�ʔᢩE��fR�ia��N�%$���2�jJ^�eG�s�`��(D��6Ą'B���BdCy+�^j��8��3�.�׎}J�fv&9Kk>�"��V���G)�@���S5mԮ�����smO�B����"F��Ww19�i=���:��j����@~���R��wL�r�������18��"���y�b3�b���0,�祉!�m�)�~v�TIm*�К7Wٻ�f1�Y;�!�*�w����hv���Ɛ��̆�~)X	��#��й��2p�ܣUZtN(� �	�6x8��%h��o],�j ����%���,�"�U�/#Θ�$T>�)qG^��p��:
�OW�����
�Z哩��U?�o�p��	�$��ѻ���'9�����n\�T-b��9Q%�`t��8���#.fv��&-���Q��iqh�뺉g��1�o�� ���玣�E�y���BWED#}�cA�h����?��*�Uk��E=s���� ��D��Ȃ4*�6s?��Oō�\�����w��Qp�Z�F�$ eQL|��cCs�JߜH܌A��e�6�ۍ:�a�r��k�-h/��(��G>�Rk�E�[د�F�Ų~RU��}C�~X��U���U��i����:,�dH�^�w��/DD����:P U����0�c��sk'��Se�.Ҝ"F���q�Tc%=�l�A��	�PS�A�C��GN}�r�'"2�M}�m��(j�K�:8�����p���g����NM�.���Y��o�I�o�`�6mo0O�2�Ȱ��ǵ�m�Jк�.ƫC����ntH"�vZF��7LLͺv?5��)�\������R�]
�z��&]��4���an����v�6�����"4>�Vc�$�2V'���ڭf,�S�)�����2~W��r�s2{#�5h#�m�x]k���n`,�W��}m��ΖD����?�!lȰ�ǦEE�'��D:��1��剏,G?���p��Ll���zy����A:���rYu��(8���0��^�;L���=f�p�*Z�c"=�O�Ln/p���44|A##�Ђx�����	M�,bI�+M���ʻ.a�!1���m�B�{����}pS�x�͌@��tm�A<p5 �_�N3���`d��>����3�*�L�n5�^��2Q(�y�E��Be�/v��	�5����V�i����w-Ҹ�u A\+���d�9!��2��с����A�OJ�'��n��϶E4ϔ�Ͷ:�13������wBS/�M4�WtUؔ^����IE�IRA��^���yG&�U}(�sU�殉�и����d�ՉP��O`݄'S �h�A.���ܻ�����v�(3��-՜S��lZ���2��K�x��)��.>ϣ��!�DܢM!*	vmb��^ Kz� bWrA6�;Y�W'b��u|_l��Y�u�f��D��p�R`:݅.�)��M6��T���L��$���y���8l�i���R<� ���O"z"�o��=���Xї�
Z*�ZU������|7��'��J"G����Q��(���~�,�d7�dZ�(�"p��ZXY=�~�Ԏ�ӵf<�8������:KiT�,F��X���A���}���7ݙ�,�x��m�����E��P�^&e�L���/ǐy+�?�A5�zUx�Gl���1߉85����p�Z+V:X����9��r1�I��jU�	ͮ�!��]��f���Qa����r�hY��u>��u'C�q�K��$�eon@l��T(_�d�r�z۷�n�8g:����,��1D�f1#I❇�9�"���I�C�������j3O�}���OM��Ѩk�3���]ϓa����ū��}��*\y�^^pW�+݋�1��3e�b��"�����9a�����;�Ѩ�X<;��kc����J��`2�i���g��FB�7b�LJ�Qj�(��#8N��y65�D)P�0ݱ���'B�������JōV�'�8\��-,�����G�c`�L�|/�����0�B?��<Ɠ�8�/��&���G�)�u�XD��nD�>�!�����b����!>J����`�:c�|��G9��i�ŝ���oZ�*+�ZӾ�.Pߺ0�A��޳��و�(��
Eeah�H|�I\�a���a)��υ@�1K��~N�W7��4��63\l�K��<$|���^3�5�2x�	���}`q��m���D7���!ޖ�EOk����P/!�8�5l�ߐ�S��bF��?��11E�~���H2�w+��`�+�����AX �Q7�g\��nl�7*av�\�?���;��f�t�(�b@���a[��ɕ���N�0ja��!i����!!�x�6�]�m�_�� ��N��׆�]�+��6�X�ǆB6:�{�1+���=�|s�x��LD�+j��0T%�]Ӻ�grC�Y\�&�M��u�=5�Ā��͡�#���8��i�g"Ӭ�V0?@�g�©�	C2�������Q�یe�i�F]oT�<xA�k�h�溺�c���#z�Hx8�i&�)�2F�݉]�{s�}�l����E�o��h���~=H�7..t⡑vE���é�a4���oOj{y��&A��"o���B�_��}�4��\�1��M�F9���D�Ra{c���na�1�'|	"ka@'{�$��d�H/WO���-̸'�0����g�v;2���P֬W	�KB&nEFk˹ⷪ�<wD���3�;�*H�d��y// ����F�y��e��C~W�8�m�%i���]Z�d����Ns��bہ;eg���P�_V�����!�b}�;�5CS�]��K=���䇊*�'+}%k;'lE���7�If^�'h�� ZDn��Z��|9b|ζԌ�$v�J*.��|8�Zw:� �N����OTfԓ9;M��jY#����C�*��;�_���RK�=���K�rJ
��4�I�n9�Dw<0�mu#�7Z&Dv;�4�������wF��ԲhTt�LTJ
(��kz�o�Q2�����bM̜�RT�����\q�yx^ęio�)��n�a����4��o�₇�#Q�B��uK�Sm��R�P�'�^2H��״H.)�l�#���y����a�G��g�e�$�D���e��0�ҙ?mψ�<I��a3ڀ�n��t�}��r�6 �o���0Ș�!b�)�|Ń�)$�<��ȱ!K����)P�b+�D����-�e˨�_��T���;A�w��t6%jw(���F��T�1B3�0/Bqy��� ����'�- T���BQt�j�#/IJ��,N��W�a"�:ǲ�o�+�}�"�9�| l���)��&��p4@d+D�x�C9[&D��F��4�ڏ|�"�U�T��/�����Z!�`1�ƕ�?����8�h廐4��.E!�YÄ?��"�o)�y�Bf������κ,�&��GϢ��)M����d0"�;W�1 ks6�w��Jݍ%�3�9qlh�� �U2$�0jo��Vh65)�,�!'�����<�ַv��WfaMB�.�y��t���"���-m~��d@���+��I�:���î��g�(M)>����6W�_����8g7�:���t�b�4F�����)O�=Q�-Z��\UG5@�ޏ'{��w�EZ]d���T�\�P��� ��#3mw	�3`�J���xQ�S̊��E�5�j�,�R�<Ca�6i�ӭ�@<kXO���@�Ҕ�ڈ�ɵ�����/@f���j
D�1R�V$�+z�#�	�3q(>�C�>Zh)�����m&mD��W��
j._$�>��%�� ���-��͵�( �&��]�lh��A���Cp�eR�I��Q���C��rF�@�i��ۻ00�z(�\4�ݏ9y0�F�w�J���;7��cFB��=E��ndN���A�M��R%����b��d�"#!?�"��1�̨�4��i����	�o�#p�U���ռB�2
=� ��f��雊c�R��Ȣ�r�^s��p���_�Q-�T��k�!9�<}>Zt�鱗�b}��T-��4�0set~m�n|�m�z�q�@)+�~��乩z;q˵�=O�Zң��y��ɘ�����"��[7C	8K3h��i�dH�k��]��ac#6�D���ݶh���y�`ͬ�hr�/����Ym�tb���{**i��H�"�!f��9M�zG=��6�Vz�}��bF���F��-9�B�ɼ��#��9�6����n��]�`��o�4��������.�������$�W� ԵP��"��z[�歷r5���Z^s�@Jn��謼8��Px�
�L~�e7$f��!��Tز-rr�5�����[,;�z�ȗ]�"�#���=#>�]@-�Ԓ��m��G�EG�L]��g�\�|�=�yQm�+n�n�F�[�?��+���ޤ:?��i��p܅�k�G����uq;O3�+��Ǻ='U^cO�q.�DA*	�k"�ˌ�VF�!����d�Ω�733��:1�Y�1�����b��TQ
G�D��'��l 	�vh����덆��e���?DF���^9Fs$����aA�C�h�,Z��6f�I֓m�+���R�/F��O�o�
R�ʵ�@�+ ��c����ˋcw)Td�� H��pCh���o{/�b���t�vu�~�%N5+K�m�@�ZI�n�5�a�@a>
�Rn� �j����|��E�IwE`toɓX��h��;���r����
�%�B��/Y����Z���F�O��ER#?˽_��Ħ:ZU�����_7���2�N�u��`�g�Du�\N���1����;�,<������8�������*=6+D;��1\����'���	���ۿ�n����m���r����5����\��Un<j�HP���L�򣄊C�v�H��[#�#�bC����Y]%{ �a��d�Ca�Jd�Z�ՠf�Šl<Ap��w������Y��g�^~Q�v5����$��&��9�{1�j����j�'�bWE���rW��,�����%�%PS��	�@�(Z��~�F�:#�#��/i�O��w�2T���k�޳�}�V��Y�K��Y�s����=�<���l���p�1Q"����Bm��;�UB1��B	�)y��8r�E��֟��n�J͉ϸ|�8� ��K��,�1c�)��ip����~��A��C�V��.��< #ڴ�D��Pmv�	�x_�������������ϝ+mE�ɣ�%F��� ���V̴�
��A�p4�׊��4�J�kg����47�����MW��^$�D{�E�7��Hnx˱��N�������R�K�^w׈C<�o��)�w���U����b�E9�$��Nh9<�9w-�V��7�>sW�v~�EFD��U��X �gĤ���xvˆ�@�p��p�\�]�qF�Hu�'@�ˤW.JӦy=Fr��e�Q�����n�wz9j�{���M-�7�&�'��r�A'$M���IX�N��P�z�� �v�=l>:�NӋ�E�ڴZY=&��T�`Vf��߲K�k�_��Æ�\o�*�p�nE��E=������R\�#��*�'vSQ/m�͏GǱq9k��u�qaq����-I؆�1I�lB`���ع�O�7f�*��	�6��(M���q\��]�t@ٟ|������v�������W�������1��O ~�(�Y�����2�Mq�C��c�}W ��^��I�ER�snn�C$o�ZO�����aU����/���S��_Ua�
�'��+8�&��7|>!�����3�©�׮�˞
Ɛ��	G��1��x��;��M���uˀb �vtQLC��H�ȓQȉ,�=��_\����	:�}_k�l���/B��<����@�'K���8ֽ7�����m������}��4��(.����7�
����� ���lQ�v0�+�ء�{_]*m�`�.΢)ѱ�R���0t6�� �%7�#����^w7�Ǯ�qb�'2��^R?���Ɏ=�?���M�\���x?~e�����>��I����Ջ3`���i����e�5���0���{ֻ��֫���fc��X����*�B-%9el&��U�N�ed���q�*�޾�4?��y�e��,Yb�r����<�|���� ���6Rvn���j�+��e_������.�U�+�j��~����8��z��
a 16]��R��m�!ٽվL�u������m�=�q����
����@@A�A�w[mS$0� ��*�R��ݧ�7��J�Xu:d�1�H�d\p�j��e]�����.���{�b{ْ�KⒸ����n�_�	������8$�~mJ�J��r�b�5��W}$Q� Ҡ4�����4��f�[-FPHp�Ml��lv�6����$�%��!�#����S�X�%}���qt4�\
J���̈C<���.�n�
zQ�ͅ��@6M"��A�V��_�_,���T���w��աm��m��&5�0��SQ��zz��r�T|`@%�F������=w�dv�B�OO���yiM�}Cg�#�Lu�#���J� sj+�����ޟ /����^����b$C6d%��m��Q��T���q}&�s�~�2���*�{�Sޚc��O�pCs�VW�5�R q������3#�\c�����������  �S�ɖ�,�(P���h�yT��Y:���I�К�.�c	���A�t!�a�~������D�-��&3��j��?W��ų� ��y�ճQ���uƸ��E9^�?c� �vz]��t���5�s���==�������f�u�.����rJ�`2t��)�a�!�S8ؾ�f�I��*��2I�ё�z[ǯ�&tƑ���]C���
�p",ܝ��ƈ�C,�m�Ty�RsR���܁&`Ib�	h<�\������ ^{�B�?t��1R�2b�����V+��-Y�݉�,�t�TX���^ZW�(B+�#��;(�w�Xo���q�ojrpm4�;߱���K.�wrXny	�A!�׉nۓ����^�3� ��6:NF��̨�E��># ����Cα����O[�β?J BSsk�#�|<�|��x>f9�_��8����B.�]d�k�_�!�F$!!M�4�Ƌ�W�+z���ϰ��*��F=x�C�Ϫ���.	\��[Q�h鼞'������{�Ho�}����v�(��""��Q>zpx!L���Y��u���~�A�$f�u�XR���y"u���%oі��Qd�	�6�/u�Sgg��!�a4eݍ��VkU�2b���t���E���^͢EKț6^(u#��� FЦb�l�"�Rq�>(���S���c4�Czl��HL�V]���h��-�ڦ�|_T��ʗj��6&�K�,,G#�$�������zn:�쥈�n�=���L4�jl��x���ÿ�<��g����Gw&^'77sm^pv�����'�p��_�ݘ�^�j�Ct,`��Pk�0VE*��'�:*�����:'Zf�V^���k�8�b\Q�.�~��_U�c���o��%�߁|���]�`�P]����׷��fUH�L�VN���ջm;�+��+С���j�bn� Lc�������!�33��Ѐ� cf`�Ԥ98��R�����D�����_���˖-Â;��������9�.I*!�WHʝ��C�^�#He��\��C%��fe3�&��IY��Y ��U�Е�f�(�ܿ�J�=+�&�ΣX8y&Ln�\Fraf$�b�T�K�?�D9J�ˊ�t>j3�\fed�G���ѵ�P3�X�\�����}�� =�g�/U��F�u�P ����-`!�$[5?�x(o���A(�l�I�ȟ<�`�B��S�l�.,[��G�v�#i$Zc�~�U��x[ݴ�mϚ�}�;]Ҷ�H�Q\j��y��@x��5@�6j̋+��v!�������9�2B�"��Z�l$fx,�;���x�h�=�!���]/G��Q�!mfc.��T�0��-��R5e��ơ���op����#FB�U��ڸ'@G�Э�$�o��N&fM�ͫ}�������_Y��'�����-S ��	����7�S�xR+/�Ǘ��$�c� �{�/+����K�r�wo���r6���r>+u̞�H���I�ap$�Ř"��J��"U��:�t������Jh0�2N,��J��wZ B,�W�.T4�
�.c������e��Q�8W�0"y��9s2�^��+�H��&�������y�ew|~���p�4]�����C(?W���iK�d�8&f>:c�KM2�I��
�GE�������i%��\zm��\̡�����=�4��p����E� E�;�����w<�i$�:q��K,0��!<a�����9�ZF���TN��[�v�pCT��x3;m&���cff��g9�V��<�G�Q��Uz��S9b����&����ao�Ydr�)�.���� ���M��B1)��Ѹ>*A�Z>��Y�$��	+���|;���^�%��������f�B1�ϯ�F�4d��:�l���w3)Є��!��1�7�sJ�FN�>��u�~��e��:��*��i�M��D�ysm���u?���T��&�1�z߽(3r%��p�����Z�1z��k�5����8n/�]0�dᜬ�Y�(��(أ�J���T����~�1��
���w����]x�/�n�dO'��g����,����eӥ�Q�G��;)�����] D}�J��/�ۺ�R'v㦹j�.� ��w ���t����ܭ�!���t���E.a���W˅�t��s�4r����IÒ9�yOU��I�+��L��8�Ӽ�Vc7i��$�v�L]����_<�(oS�:�� �%��X�����=��5��d�w���b�/�q����o�jBr'�_}��m����.o-��^���kVV��h������,�����8,a@Ǭ�i}׋֔��a��ZY�X�٩@'�^��*檴#\N�+v*� �+���Ϯn� *���R�J	_�~�
�Hŧew����~�D�K�V�p�:Z��3-���m����nj��
'� wq�N�kd���Ȁ�7��/�����	�3��t�:1c���"Xj��h<���[�1iMPR��:�0�CQ���CP@�mb�V����ظ���#?Ě�]>���6(l`@�ct�Y�1��ϭ�R�:t٨���,���iɋ�Č�jq�_?�J��_�R�Õ`�����ޥY�a�:V�ee�a��)�Q8�?KN���q���]C[=&��F�*�k�|4�ۢ_��\���]��膇r�O2�a���@h	@���Iޖ���G�繦��Q��!����ߣwF�:\����cVƁ^��'���X��XW'��È��K���  5X����5�ZD�ٴ��N4�z�\~��
���i~�93#�=Q��Āp��b��������:�YQ�z�n>�'q�T2�c%i��jؐ�h4c^���j̀E��3�S�a=)#^a?\�}?%�l'������b<v�mS5�P֝'�؋�m��yay,�nv����Z-mAb���ۗ,��9>�{�
�{�ˌAE�E�ϸA�ak�^�h�6���ѩ��9/!�~����v�������&l~������T�m�b�1N#'i�xf��mV����s׬Pv,�;r_}|����K��`Atjǽ�߁��������]ڱ�z5��
(�����*��yg�n����*�S���e*EIL�^���v�[l�ګ�g[�n�6@WWދH�T~e$S�?�j��Dyen|�Wn&���8�ˣ��{I�J���sE�?���5B��Fo�IN�;���s-3��C��. �,|1@�*kI7�N�j	�L�_\���eC�z^�X�kŴUT��̟�7��
u6�[-<�߅,ޕ��m�?����H�_E�2_f�b-*� j��-�|l�t@��V�(�l����l�įXP*6��F�_S�]�n���'x��X\+���\�����)��!6|�(lO�;Q�K�|����0�o�J�c�BgU$�����ۏ�;_������Ĉ2?�+�OhV�0]lY[��$��� �������\���׃�'�У��1Wp�QzX�x�/' 
y5B��X]��K$�Z�ILH�[�R1L�[Ζ�P�5�B_�W�6����W��e��	IGՃ��d�4l�ҏ�W�����n�M�c($ZZ���ݮbk�}|���!.0�iY."�o�\��w��5��d�Yos%]�]7*����~x�Ұi��4�ʒ�y��O�7�������ad&�#%�±>;�=§�c6�n�kR�^ݸP3	a8���|�睐7��Z���fGlE���-Z���B�<�����K\����*7G`&hy:E��^���6C�{Y�����v�r&�=�̦��M����=t�bx�D�����: t�.������������\3���d\h�'Ż���4�
U�kK+<+�Zl�U�W�k2}^Ƈ#��QL�+{�0�|�~y�E�����TR����v5��=��HQt����Uj{���ߪ!�J�U)+��~�U��"��pm���{ͨ����>��B*��G �k��H�t+X%V���9#��e�K��&x�;�e�;��ԭ��|t�5u n�훋�.�ޫ��rl���m9��#yP�c��$ӤͽW�2Z��$�WX� $<��z@7� ��>ΓS�[}Ɗg ��X3p�Oe�]�Ŏ�#��XK���~QZ��pnW�"�a;>hD��r	5Pػ�tz�w����|7$�uKHԶ�����K�{��,��[Y YNr�\��_���5k��'(w���p��9U旣~�`�S��x�!�y�	c�h��hR�tt�M�wN��d	�@W�7�OO)	�˾}�2��E��+}�U�($�qV�ІԈ�jhboiw�=����)v���]���:����q�q�N1�Tm�AIO �;:�-I�gz6x<��xEd�>��}C�<����ͦ�b����ھ���MlG�w;��A�?�"��:�2C�n�Asq�䦐�ز3E�f���@^ث�Y�ubY�;b���,���5�S�J�LI&�늎^��p�}��;����(����o$]�¶up����� ����fC^f��(}G�=�������@:� �-�3�"m�h5���<�W��.�RG[�����{�/?H1b�p��))�63.��5UOHՒ����Tԣn�ŭ����<�𗝆?.b{W����`�@�lu��oX�o(���ԃn,nM��Cĥ^¬���'�Âe����޷�s�U����� w�4:�w�.�	p�ƨ1���ą���J�"�z�> f��Fa�Vh����c�ŨA2N��=��E�����~�֞��_ ��m~F��:���;������jZ^���^߲��{^#qXGE�M�C��Z��4-��-\�Z�&ĝ�GQ�<X���Z��N�Sƻ��xo6)�C_5n/�>��3��z-�P�9��nF[��s�o��ܕtd��i�hI-�x����ȿ�-q���)��yKuQ�FA�U�f��
gwOLB\���������КPbAݝ���7�ěU~�����$��eL�E�vKhЂ)�����*�c�Ab�ϺW��S(:��r�D3�7����$	z�( d%.�N�/-����~�;���5�s`�Im!&��gk�h?�g$ű3��$���!I� o��r]��w�~�hY�@��߲p/�54)픖s�ڇޟS��ɲ=���zͻ��G��ng���6��nA^������7&!�sbF�c�>˧�����p� �gz�z�2FP<�͹������b��~�<��6�|ʫ��8�Ԙc��6 #��� c��h�ݝլ���b��s��b���+�{���s�}hTk*��`_3s���v�b	�G&�=2�5��x�r�'V��kڱ�E⩰}1H<6F:�z3�q)���'�A�t�^�4�/���p��:?����W^�TD�to�v��5���$�U��Qv�w��"ͼ��*ȡ��3[�Q�~�0@Iz�|cO��8��������[���5G�	0���Ex�9�y8�/�l����~g\���-� +`)�=7áe5��ƍ�0��+�Y}��l	0�Y�Yb?��$̫E~�B�$�ɾ��8?��F�?����s�5�b6"��c.�uŔ��_H����3I5Gq�U���𼧵�&����s{q\����V�{��d� ��U����b���T��~�WC>Y� �s����A%�����8��e�����\'������i�<vXZj�1ʊ-��p�84(�iiW5_�Ae<�9r>*Y�����o
�z���c"�����h�����9���0�r�Z����	��l��s�k� �C��</��O�<�l��L�0�A��|�DT��v�=Γp�n��A}g݅�+A��:����1��%��b�����4�s��olfd-�\5G���R>9�`?މ26��f�
R���GI�N�V{ښI��+��=Y��~�k�g��k�t��$ƭ�[�#y�M�~w9���&��t;�-D)G���c��j���>rI��<�-�Y��[LF,�0sZ�L���L�2�/��H0\��4l"�5>��dC��� ��6p0S#UV�����������O�G��_d8c� �r����v"��
�^ց�X��L�UtCؼ����m�3����~`�!A���++zn!��=�3Sy|&[�o3!�BV��1D�'��b���}���=gF�2{4��`�W+Lvmy��?�M����^�8 [?Ji���A剨�����6��Z]<1lV��P�r�ߢ=p�X����|Ŭ��٫2�(�8���nFA���c�qcŽ.g�இG�S����љ�����S���8� ��
&��{K�.�~6/s�2�)�� �Mn[3Ӏ������o�'��4y�z��X� %�ݸ���t������K�+�0ή�q!��G����d,�c�c/$+��c��ա�ʪ�5�'*��m�>]�\���z"��3O�?D�	q�Jur3��r�ޠ��x�`o�3&ȸU�1�Q��"ǣ|���`�(�Z0[;� ������pu��:
ߴ
��~�>�^�`��m�O��?-7�~m�q���̕dp�fI�S��+!qυ��򥕗���Ӑ)�T|��%�G]iXy�Qq;��3a^`����y:����P��¾@�z�+&rVY^��X߲��]�)fQ5�􁢍1����G$�pnW��ah�z����2-�
va���]^-�=��Fj����n�����L�Q�p�K����ן!�e����Tj!��{�ʋ� ��iN3�t���H<�D� ��_�c����~m_�5^���1�5g�'�H�����-y�0�k��z�R�3�q%����iL�B�QxF�]�R�h���@��`��:���T�����C��&�B�ltǡH�8���,c�y�_�v��.[/P���v���W�6�~9��-H�k�>��^��.G=/h{�׶�D�c{����D��ն������y��9�Ⱥ�@�I�����Y��ư� ��	�ջiܬ�>}�m֦@0��af���#v��4(�=�{]3�}��Ttא�m8�;@p�ۃOW�!=�On-��j��%��J�r���װ��=��F- sO0qE���)m��5K�l��fu.����TiЛ��X��8K��|)R��gD�Ә����
���ʁ��锥�����FB`m�i=��q9��v��� ;$}�Ɗ{�vC�S�Q׈9��J�E�uz����O-����"�g�yu�-5ԧ2@?jUň,�1������K�b�EŰiqq�
�8頾�S�gѨ����� �͛C�y'�79Ԓ�����Z��ցs�Nc��fk��D�)9�G�z�2���|��49Z]�9&�=dS녨/������'��f��A�t�ȡ���:S��E�k[�a�2�C4�@����V�]K!����K��t*5^�E��U���y����V��נ��yMd����������M`�^��T.������?t�'W��w�7��iGQ�f ]A��|��T�v�vH�D��+n��2��C� �o3B+\q%��F�8y d�6�qt�Q}��{&KJ
KC��:����yx���<
:�e��w�bpy�R�{D��n<O� �f�|�m�:��G5�\��5�����W�����3���#\�ȒD�F	p%�w�-.P��d��JJYg!G߻�^5.0�^k����S�%p�R���Q����P���-��T��͆����B`�ܡ0fs�T䛣�^˭f�П�Yڧ���a���p�E咻>u�]�G��V���wW������g31^�!����WW���X
Z�|���돱��h�����W�d4�FXg� �����2�T��)<�S�Ox��ݦ��\����G�ϸ���� oj�Q\V|Cr����!H��Q#�D�j���G$˷c��������C	�x�B5�E1���!P���L��l);�D���g�l�F�*�=.0	F�_�5��u��ah�ȭ�H�]�\K�Տ�^�i]���R�X��^�;�w�6�7��SM���^#q$�������j�Α�rw'Xs�� '-�k!�)�ڴB��'��@ȐE�MX��t��0��-� k������������ޡ�J=�X���
OT�����|��I�`N�X�f��z���)A{���I:��}~��d.Y��:{����I�n\`#�pT��֐+��uA�'`�_�}�t�[�e��
;vL��񡳙pɲ�X}n���>�>.�Ԟ�ۛ�0��[Kw���P�9�¡^9I�R���ퟰ����I��$��K4>�OQ�m6?�\R���楳�"����6#����By2Rza����OᰯɎ��E�4��3��T���\��i<Pqd�l���Z�
���{��w�s�7_x�c��=�/W:FbL�9 �a����y�֭��dӵ!8$��QM��wt;�A E 4��*?�"�Q2V�Tk��č��a�3����G*�j{�_qVlyK۸W� L�!����JSE5��%k��k�+���"�<�u௽��S��dso��h!����)_�@��/����b3�����F�38���4�R_�._N��bF>n�=�����_�W���-(���F�;��@m�)�>��1�英ݾ�CzI�6��H*���2tD�I̬�Y�D��F�I[��T�１e��`xП=n!��fuח>��{/u�#g���iKff#�&0���ˢ�
�AR1���ጋ
7��Q=�sՏ�l���ͷ�$hʠ�vB��	n���D@n��+lr�y
�EkRc�$�L�R1���?~��tlz���6eN�r	!���Ǘ�I�9� ���8�X!u����yak�mW���q�w�|�G:`z#^3���$�bG~"��%��p��kA���:}�b�߷��˫�~����ӲT�p�̵�9^Ĩ��|O^�B�+iM� �@��`�0i݋��{J�/�H�x�8�&4�$z�y�siI�KFfC07��tظ����:�&���:{0t�['Iie�f�[�}����T}�@���G���ޱ��,*)G7��'�=�� �w�)�㤾�FKW�ws%����$��6�է�Ɠ/���PdC��|:���DWbA0YE0J�13���t��1w,p9[�{�Q���I���c˟��F�&�t�b�*�n��)t%�~I	oM�.^rm(��X�#xHsQ�ق��b�[U�v�o��, ��f��Kb�?x�ZY��P8�T��LW��'��Hs��R�v��A�׮�]���|�]�Ԓ^�=2^��ǃ��e$1��yK`�"�����%?X��nۗ!�\8G���x�|�|ٯ
N�:�;{³�P��~�7E�W�箮Q�b��V�:���d�DM�����m4/�&7�GފaC�]����������ʃ�����O�7��(hY+��;ԁ�� ��mPn��J����!��.�`)�S�p���Jj����g��*:SR��r��,L���-�Xf��~���:���i��F�-zW����52.^~O|�*�n �����m么	lI`�~��Gl����D8��@X�-(8�Ă���U&
�E����Bt3R���3SF֯���e�QB�j��˺��Iҧ]$r�0�s�������;n�f��֕2��{y݆���&�Z`���O��Ԙ���>��r_X����_�f����\���$$�������1�Lr97���?���{�(%��TU����$VM>���FE����9����.���"�K��`%�/`�G���ب1˾h�~���1�i���x�RW�TF�	��KP��_�n�l$�W���.y����qQ�Ԟ�j�:%i }�GD壸B+x:]�Q������F�z����Ԍ�ܳ���3�I���
��A�E�Q���������g��?�e��b"
�;*"d����6���	&D���"���/o����u��g�ʕ����1�OEz��y<��w�v���-dI=h���v!��_ ����.�����#��(�]�֭�Sk)�.����:�G&'�W�j�zC��C<|×�/N�����do6����SE��F,�֋xS��g�?��C�E���_��U�1�f{\g�]k;G��[W�Y8�^a�L�t3@}d�~:�Ne����_�r��TB��b��@~�+����JU�����n�g�ht� �"Nd� �`�(P��Qf!��!i�($| QXo�om�-��K�oG�J�z�D%�˝����I(XvG2�9#�$�]�~~Yp�N�[kv'�6(G�~Zkb:<�FM{�� �Rug��P�	�ֽ�C�m�B0v�~��miS�����mo�1P�m�" ��Q�ى�v؞V�t���i��G�q���݆i6A��'���PN���_�2�d�g\�~y�c� ���Ɓ4�:�n����;�/p_��)�� ���mPݚ>{t���Nd0�޼�i��l�����'D�ō��a<-�A�n�ͤ�j'��"~�gC�.�����v�C�$��[��K��?@	P]�Wc�!<Fo���v�!]�U�kPw,�h�qH(��#�>����I������g���{^DŁ�P�^��S�)�Ұ1t�351dcv��}�M�6b���K"��n�b@h�kqy��+P����#c�������]��>�Uz��&P��ugN�D��F0���K��C-��|�0�D�V��71��
���G�;�֜�ynPJ��-��Z�v.�cqf~�s���� 3�x�҇U��;���7-o�b�/g]��k��}{��a�rY�a��F5˞���p�G.�zo����6Cy�K�z�8�����{, ��y�C׽�sq�٩��զs����R?�|�=�j����K-X*	�,?Bm���0�q7Q�$Aw��,��X��P��B��i�s� فߴz����P�U*��܎�Z�n�Vg�2���/�S  Mvܚ�^���l��
A�4x.U (<�<?|����N��B�i���)3pzd�8�d
:�����W2![��C�xe�����[vˎ�/4���ʦk&ȶp2J�@��3��0 HSs�4��g�˵r7��5�����B�X?Z�<��=n1�i�������"�k(/u���ʼ�_��E� �Tq�N��*���r�pv�i��~��H��:��\��m���q�̢/���G!�8qu+�Q�e�KK'oBv�
�h8Kϱw�o�PTs��)�nF4�>]�;O]�Akj+ܖd�29�r/m���5L��6�$��Y�f�v�\D��Y����/�u~������N�Z\@��J{�E\|dWx��~~��;��Y%�r[���h����d�E�j����qM�kR	}cQ''�W�zU�'��
5����a6��K�f�z�4���G����F8J�wY'�^���g{Xb���͍VU�m�!STb�<+R�(_w,g�6I���̂�L��G:�|
������ƾMv��h���ʚ|�J*�%wlUL-�Ix��H=��Cٞip�����}=]HN�hS�7�74�� 2�g?�?���^�N�j�}�����eN��Y�M��2A�R��&ѓ�̉��B�Ymk��������d[+�����w�|���h�����)��y�r��	�0�p;��R�E���%��N��M���y�a���S�ܝ���'`�X��Ň�T�E�"l�NX�/�U�/^�a��?R�ʦg{k���z��a��VY슮>&����$����g���<w`/e���X%\]%�B���f�i�7�R2��m�y�U��u"��d��86�f
7$i��o��RDŐ��;ćD_�^��V9�S>�U�2IY�����C�J5�_���(�yڰ��Z��;v�n�"i����?j��E^�"f�N��Q��yj�e<?�Y���������ȵ��U+u4XRÕ�ܾ���?:Pxz��k
D>Xm�F�\n��%�<�Jj]Ef"�=lb�t��2�q4���Dm7��H5Kq�<���xEᵐ���R+�� "���� a���ۂ`cF>�p;Kͺ�O�ƒL��o|jP�5�>�dڕ�u�.*V?d6�c�,Z6~�*74c��5�0u�_~H�Q�k��Z��y�mM�l3�2�ױXZE�o�Lj�Nf(h*�V�{ x�'��� ��0G~�}v��u�����;y�b���M�(��*fL�Ʋr�w��W8��ބ$`(֢�m��ҖpNG�D�l�����pnB��9��B���e~߭�I��]�IV��?E�}x������H!��
�~|�|�-�7�C�üx m���������2���E� Ȥ�:�Ǆ�p������h����JO����%vp�%��%����@Gq�\d�?�W�qٺ��x��_~&�'d�ܫ�0�nCƠ]CmA!�\�؂ �ؔяF7�oL�AF\�A��� �,!�<���~O4��椑����&�_*�:��Z\0��eG����"<���[NZnA*NN��S�����x=f7��͇�r5�-V�x]�@�2!�o�}ͨ�YK�#RS���rH��%N��{�{���+�y"� wu�2�*8�:���.�pvo�+�'�H9�������P�:�B��{�^pZԢSa�G. ��:���R?�GmT��'K�<�}�>�%
��5Kl��hhIm:v��Z%��2�55��0�;ol���7y�W`�K�����n�r+~x��Ʈ�s��qfx�@F������5zoR~dy9S�'Lƈi�9�W��(����Վ���,n��6��h�FL�TԹ�Cc�(P�8)��W��<|caY7�r��͆Bȁ�-1��BJr�����o~lZB���=]ĐL�r��������Yn�yNa[K�A���̍���m֜��W��E$Z_NZ%/�77i����$��
��)�*�j7�>O`}?��u"�Qy�X�q�n��O�%��e�Y�k[�
 �.��rfu7]s��R��n��9ph������<�o'<� %������Xv�r��6�!aN��7��6�znMqKw������z��(kЌ�ܠ ��C~�Q���@⸤5��6��{���TE���$y��U�Q���������5�`\�"07 �W>*-W�ع���vmuz��|qp���1���&�@�V?�ًvU<�n�Z~q�f-�K�-s���:A/3Ϋ�B�X��㗥)�j�8�.���lȰ�([3�eܐ8W�L�����^J�i��ϭ[Z�v��Έ[��?��2k����Rʻ@����䯫$8F�d� �wns1i74�7�Tr�(@Qq0%��b�o�V��S��x��O���{ЪYk���F<�"dx�R�>�(�	Q[�[=f����j�Ҍ5�	�ыS4K��e�lVIk��rGݖ��=�c��ip��vc��ܪذ�L�A�'mo&B��R�_���Je�w[~)R��ϱI���.��o���N�`�[	OUY��JC�
��1�ȁ�pcxB��I��.%�җ��$�[��۷s�5Y�	�v�WskZ�����JBw:W�U��DHȁG�1߮gZ���T:�WZ�%��`�ʦ���R<o՞���i0�%%6E;7�����:�M%S�;fl�-�ł(�}�ݦ�gz���qd�rs��e���X��h�Հ����Jz̏I���P�A�~r���
vz�u�%����9�^����7].4ҷ�7������bo,�%�J�76U߁�<y䜯����=Ja�y���W>�m���F���������љ�S]<CG9R$�[Ԅ���G�5)���3�!�AXxd��Y_��΂�a89?q äX�%�O"(n9����$���Z:/�b��
CBZR�&<��"DR���t����^�D�5�d�K���+zä�p�����PX ��,uE�-��i��%�^�`�ف�������W[�5"��ƍ��r������?l��T>/��,���T�US�ܴ�j�9�y�� :����^�^��Xp����j���J5\m1z�و-�:ϡ �Ⓒ2|����~�R���a��C+�/W�^�!d
S���N���&��i'���e?�ʛC��W/bYs��/��S�|0 �d��%�%���"���c,+�2,�\��L�v9���H���Y����-� 2�D!KmM�)q��2��OIu6�˯���he�zs�.�T�.���r�?��͗�;�OLFF������7���J&@���C��MY��j��+�)+?z��Pw�7�_$w(�g2����Pd�[P��s�T�a� ��P������KH-�#��Q���<��;���Qҫ�w��A1�G��䖻Oof/~K�M��:_��#��Y�jX3_��_fBg7�� c騹�����܅���",���o\I����E 
Ty��@�jh��!�Y������0��~��O������lحR��'\�g�r7��^�iT��9�[5䆓���	�$H�+��Em�i]�1���v4:�W��D�X��9G���^Z�����!Z�6<������Qr�k�L}�@v-�=��W?o�GG�U��=�^��U,?�Bn�&?#���?m'u#gpf=�մ~����	)�;�1��Cs�����M��]8�L��s��8����qo��b�M�u	�V٫!l3��m<�FϷ��{{<�Oô� �)��l)[�W\��u/����Y�Z��{�!Q jH[y�h��b
%{qj�op��?�"?�<;��T�$�N$Ԓ-�
v���*1���}�G䊿)����5�諪��F�n���A��U�?Һ>��@.�;��� Z�P�8'��ʵ{<S6�d�!|i5�&��:8��pa��&38C��=&^a{���j�><`�6���[KB�u��܅�eS�Sa�M�bj��^� �'7�B�H���#���y��޼VrƲ#�w���n_�kn�u�r�
��:"7U��ѡ�T {[�m�<�|&�kL��'���;}Μ�j�M)�����Vyx�u�*�a���gQ���|�J]q��0�e]�l?�1�9X���8	g��Tnco�M�[���mCa���S��}R'�?����~y����@`�h���c
3�r�e��Q�٢�,�m��os��A�>�>eq��{[���O�����F�~�^�X`��̻+-�|���58
����.l�;�at��l����l�j9DtƎ���|��嬁Rщ
��^���N~�Ht�	�Q�T��;uSV��-"H����!S0�7ӍK����A�6�7�iה��6��.+d2�׈+�����k�0;��Y�z��;���G�۽�܊6Zd ;t"���7t(��
l�FN�q�r��z�5�v;.M�ѺTM�lo�R�Iqҿ�s{�����^A^�U!
��An������J���3z�N��N������M�J���8�m%j��"E4�}	f�Ku�V��������7l�q9�}F���ua����Rf-!��#�FjM~V��J�Ll��섘(#}v�^���p�| K�����,+�?��Z���X�L�
0��/Wa�6�`/:U8_�L��gM�,ɻ��nǈq+�H��e0 !��P\U k�����&�?9�
ڇjW. ���I�;�c쏳o�-�8�������#՚Q�dp��pwg_,@4i�=��Z��/y�*�r3� &p9(�(�O��=�0K��ik����a�Pk���4l�n�9�]�Oa�$�����~܍Xև��~X5}e���0)ƕ���}K+i����E\Re��F�;�0��m1�.��̾n2���[�����z1HGD#�k�>Ei�h�f_����U�(b�/k�@��f�]L�Ӕr�$&,�cA�9?�8�+�g.
���z]�n��VG�������T,��9A�]��_R�M�>]D�F��C'���[[Լ��
��x�^���������0��(������g����}x��}\�*Ҹ�]�Ȝ54�h~v��u��z&<�q�M���^�4�����׺�,�[�K
�IO�2��:�#E ����T��3��v�eW�Xm��<�2��zɼ��E�Ͻ�(��T��uW�鴳������T�]�� ���Qm��PZc]Y��=��`Uﺂ<Uu�k�q��KT8B��l�.|Jd_F���<�!����a�����Y��\>�9>�A*dGp�(o�*@�l�;��U<K7��D���,������߫�[��P����qȃw�e��&l�ʂd����/���B�'�[��#��|�Y�es�����`D?���A�w�	�!#�%��o�@�a	����O�L<VyxAºm4�B�y��:e0�" �Zp�EJ��7�S��tug����|A��Y5�Y��Н��J�So�|z�;�oO�� ���>le��u��%�*�5������~�BP8S<�#���a��]\MKR;��a��,��$
Ze�^����C,�M��[k�����;��O�q����pf��i;�oH��m��ʥ/^Aq�)m^��� j��+�}G�&�Ss��]G��,����5-T��(�mc����#����?��E1�bN���'����e#���Kr��y-�(����/a9�gb�&�LpA�r�$���4\�T�D*1�g���S��e�h�7d�a�8�K2U~נ�����Xc=��HNm��S�`��D�b�QE[���+�o2?��J��o�D�Й3@O�� ���C��>frJi=���wX�tۋ,���zAnNk���q�G?^C�@ؓa����E ��kF� c�;#���g�LU��ٽ'�G䉔���BaL����!l���	>r����y��Y���e�Ѭ���9uPN��,>����ܳ`���E��d�Y}Ѡ;�����|�hީ�K7�W�� �Qe��n�W���2y���ֿ��9��ʻ��d�23�.�̍tI��v��~��}�:�)v],��WH��EM������������G1��=@l�o�&��1��"�]l����A���]�����< G�F댘��C@N�;9�4ȡK�z�4O��뱋�������T��\�_��q�*P�0u(���vu��iH���@�9��M��Í)��5��R��ݜ͘�al�á,����G�t �W@����$��%����D�K���@���/zSH�+��,�ߖI��&d��|��c
{�!�P��|Mܻ��?F���悔�e7��'l0u�}W<=/ޛ�="���,�;�'s�B�#��I�т7��!�.z��T�ZG�{%��Cu��Y�^7�����}L�1dw��%���Kڦ���%�K��i���<���$�$��XI'�X��4��G��E�#�8Ek����╅�uS~�_)�<�?�"Zu����u۶���0D��T�}���o$���Nr[����)�8��U��Ӧ16��f��"u��7�1����U�s���f�W���+���QCA�fxB7�Q�e�kr=����%[y�rJ'�|���	s��I�P:��q.-���,��:k{��]n�;8��?L�qy;CO0u9��G��6�1Tf�?[��ծKᠴ@����ڥKDP��4�z���䜶�Z��r%e�(�����QdE�Jl�Mx�������f<`.�lx���?��=:�;�h�3V�vN-���m7pvLL����T��osɁ�O�$:Z�G>)�c���(�C�� ~թ���0����i�O-[�*Nۦ��ߵ��Ð`pJΟ8��d�/����#v�����+0�H,-̍:����?�M+��v�EǪ��,�L�&�վm=d�؛1��[���S몆��p�@�Y/M^�9b�#��P��?�p;.�z ͡�&҃ߦ�>�aB�;pH|�db\a��y����K9ֶ������U������_�!�=}z)���_2�L�L��%�:�=@.o��>J�����H�Tu]39L6FB�jA��#�O��9S��Ŏбi�y�X��e-]+���eW.�ܼ �DE�o4��������C5*}���������:3�S$�}1��G�ś��k�S� K�1̼/p5S+����~�q>��|�V:��W�.�`YO�ӟ�k%�B�::�:�����rxRW�7Z��~��h�����n��nم�~¸2�S'&^CUN�C��kf�ں|��Z��Ē/�K�e���Y�
AB?��&�B���#ݧR��񈷴���Hm,�1ȹ��$i# ��fay���pG��:�;�RU��Z{�E Hz�/WR�SI�\h�8ʕk�,[ם���8�Z|i=�����;[j�̆?���N`�_�m��]�V�B�F8^���3s��F/,�BQ(��ջ�l�EⰈa$ڜ_|��8j�-������M$��&�g
2���P0P��@r'�7Ғ��L���{���Y4Q;�j�V�>�4XA�S��XdaB&� F).W֑1ĸ�����F ?� �>C��[�#��~��7🴌9p����s�B�< �B!9È�	�8�g�4յU�'gߛ��ԥ,��>�n�TѸ��Qg������QL�?j0BBg�u�t���}�����ʮ�]�({U�匊d��%8%�1;ꥼ�t_9�4Q��Y��� 0&Kk6��Fwy^ =�w��ȓ?�s�_���C��RE���F�+�7�'��J�lt���F$�TFv��u�=�i ����k�󍝲��`��훺�%��p��� ��</v���_�m䙒&�Tq���Az$�7��d��׃˴}�{i�~xBS�p�T�q��樑��$��H�	n��m��wp�I	ɓ�#>��ފ�D�ߒi,'��/ל����.C�(����K9���ס�{���#�t���I"�i�@��G3
��������.*r����[9(]lM��E�Af ~�|�;
x,�qUo	��wL�I3��3�^�KJ7�c2>�2Ɖ��Z������\.��"�<�����0h��	,[b͘FD7R@�ܹ��P�S�#OV��'k���y����3�Є����Uz�e3�d�$�S��57S6-��l8�̹C�Y�H�2=��D�j��[��O'm2�X��Gߟ���}�
aAvf��ے��9�U5 �!&�b;TF)[�y���cE��6/m:�+R�W��	���-$6�A��[���I����B�*r?_bX ��kr=�1�=�\xj���:d�⚝yi;,���(Mn�<S$�&,�"W�1��X��Ƽ˱�@�A�F���J�j���rJo}���U�������A4u�8�9߂�6�#	�Z$��w\�&��ް����x�U�Z��{K?�f�D,{�.��V��Y�1>Q39?!Τ}���54����JR���#�ĥ�>.4��K_�ߤ�����^�����)ƹR !E[6�ܲ.s�G�X�? �i^�E�����_M�"����V#8����ò2���n;�4%�tF���*��`& uE�N��Q �Į��QQ��2��D87�qϔ�ֲ��|�e<�q�V7s��~�vD�{�:��Jrx����3�X��1d�W��5�n�a��������'�g�7� <	���?��G��`��>�}pp����RgOq�;�f�B��~��b�[����n�M%F�d_&*)86��`�6}d�L!q��!T�(e��Yq{W��V*e�E�o�Ik���F�oŃ�s���G4�4�����<n�u��@̑i�V�5E&s�h�@�eq���mĘF�����B ���Ә��EN�9��ɸE�Z� ˨�<�5j^f8��N�D�����x%!�A�8y�N!OGm)�d�~�^��� K�q(��8��	���um�,���\���ۤ�1�����0N��!2��W��zUB��=�Q��۾�:Ӻ�e/TF o~.I�M��E�Na���6���.��2ܧ� �7�:���s��6h�\�ݕ�+k�Q�C��C�@�j�E�7��58JѬT�)�Fщ^��`-9�:R#��l�yr6M�P�3Zh2�0�@Y��GW�iM��g5�2���Qf����yU�	J��t��;(�g&x���@�@?i����kz� �U�i��
���9��įk�Bv<�l*��xAY�0s�G��N�V����k:�;@�	��ظN�,���A*�n�u�%;~	�iA��I�p��m͆"R`�k��;x#)�j��6�κ:d�,�a��������x��io�lȚ�)[ku��K��c���ҹH�p�S�A%��1��"�˦Tj$r��b��6�o�Ɗ�3�j>��-aF��7���*?�3�2�I,�/��Lb.}ʆM������MH���	���Ѽ06Wp�@�����9U�H"rit�qV54֏���U,濻�`�r�6@D���Z �~X[v6�ڏ�p:�E��ߖcR��B�b,�����	�4�!
r���㯐[w�Z�e����9.#)��gnG@� �^�jLr�E��?o��)	��������m��}"�"�U��$�5��bOD�J2��%��Pl�co�4��N^��b���z��{;�Z�A�<\q��4s��G-
of,A���{WE��v��(�XٴE˗�s�g.�t'���k �[Ș�P�D������N��t���XHѩd��|:�?F5V�Y��>NhЏ��f)z`q�|Q�}�Ux6MC�d�Y����9�(����; �t����L��8�+,����lx�x���c�I���{C���\ �5 �y2�/��Q
�{�I�����ң��_�>R7�V����|��˂PI������	��Ŏ�l����#;����C��8�Hn�+��
�-��~2^�+W�@c�+��-,$0QB�`��Ks�	�'
dN�{�\��+�P��	jp���������%�G�a9���"V��S���Ǥr��ymd���)m��R���@P���#�yhR1D�ͦ���P%����'����_w@�5�&g�k :�,�As�?�e�6�+�t֟���`�5���V��wR�`�b��z��r��Y���e2k�;�n\*��V�[]粜�~Z�p7M���4�,5�:��a��ùEm�~(^]���O�8��%U"~Y���MW���:��d�i�&;C�d7=h����a5�f#)ӂmWЈ%��V�&;i���vz�VE�TA4�{���JI:>����P͋�*����c!�ѥ#��(bqT��4�]#�y�����V`��)�t����2:K��҇tlXչQqI0�=��ª�Kh�|�)�F	�����\���&���Bâ�4�g�p;�(�s;4I������_ xo(�:���lfE�=j}��?�ݘ~���N9ң U!�#Յ���P/Ѐ �M}9	\�ȱn�g�֐���� �n�0��d��i�i��樊'�L��Y&�Ĝl�J�!�Рv���`��MO��l®.|԰��x1��Y����օB{
�e:��F5�Vu�1�܉g�px5�
�=�'�r`�A�X\�pV��.���BZ��ct���Ԝ�s���H���xb�D�bAp�ԙ�SCH��� ��� X^i{�&�(;�ev�5.��}�0��2����ƶ���M�q�,���)���7O+#���*�2XV�P��-�v�v�;��p�G3�!�a�Y�&=*���\� ��b�(v�F�8j��ɸ��E��Gf��*�3�*a��_��Ij~��n�I�+���߉���خ����ؤM�/c�:U�K{I�s66� �/�������V!�VZ�%Ѱ�fD��s�O+g,�.�H"<_��%���Wjuw�r��VO�A����fB���	x#n3>�j�ȷ�T6���U����T�7�z�Z�a�!�\�]��%�Ki����{.$ϻ	��C�:��J��$HpM1欩8_��v��+~{�+��ξ�[),QE����X���԰��3��hZܢ�4�a�Ftl�c�W�u�W�������g��VFF$@ �Vp9�^��:�i��T����y==���c�8y>�)�ql�~΋��RQ�!�	���s�P-D�-b/_�L��Jr�_@"e$��v2��oTϴ�u�c
)�nx&�ㅻ�
m�p��A����PO�[����h�)��1"P����݆|+�`��I�y�d1��O�|WS��F��QL�C�r����b}��V���|�v��@�~'�D�$��\r � fn0��_<����È��e�: 	;Д*��19-UZ��$���C�JL!\or�[9��*9��<��̲F�ʹ65��Tx�MB���d}�Jȓu��W�;��W�S��GKʎ~����b��~3}~���+2���K��՟���Xg<�_����u����A۹�T?���G�:OW�v���.'-���?*�� ����GҀ\��Όs��F?)|���-@��E�k����(�� �t�&�ڐ$�'��΄��>�$��鯀��/}�f������!�~�m���~��f�'��
�g.��G_'rsxr�,2�@(��kxx�Oo�����$�E�I��T����C1��8�E�y�r����C�ѫ�3|r9r���	�#iiE�
O��׉J�=l�#ޓr;��[s�" �RO~�A[��m��n�ń�Mj�W,`��k0�z?z��<#y��i��W��(W��Ƚ�y�2��ezwvY���v'�1N��:v���G�@�S�Q 8���!�*P�Y�4�#�HJ��;�)���*�w<����-��ٶI�S !��}TX|�Ƴ3S��1��{UZ`wZ��
��}�O̱��)q�G?PyV�[�Pܯ�������C�c�~L9��,����#�[ ����,� �ۊ  $���Z�,
��gR�@��v;� ���������$�k�|��|A�.4J+K.J�|�冞��G̿�����0����Eo"��[�:��K�[��V�ʁ!�Q�I"R�/;_�I��zZ��C�5j̺��o�jme�&�G�sZOiu}Z�b�������8{rA�K��_Nm@�s�H7�hS\����T��B<>L��m񎨅@���5F����WaE�����Ҽ�G��	�X2�usQz�/!aa��x3�cT�|�jGi��NΙ�d�_�/�o5�$owbAk��E�_����:��P�孕�	�':�{��;�� �#i��8��}q�Z[�R�v�U,��Nc	�{��{Vo�{����?���N�և<=A�����#D�	\=Ӥ�
��,��Up�&�ءvS;�sq�c����K\N�쵌1����3����Z�����]o)�q��?�;T��d��e	��x
��J*�����|���w+�θ���4%��O�`1ǺJ�fu�0�T�n�	$�W_'�8�a�G���_Z-"n��2&���H*Y��\��F�I�� �$�b;,��3����);o��S"H�x�/���V��^~�PbN�O�;k	oD����P� ����?T��.�\�1�S����UN�'����geS$��G�+�IFq�>*��.I�	�7Y� S<�h�7�B	��[��Wn�{^�/R��9��y��|��i���̪V����o!d�B_U��N����P�ג��ڄ���B"C��J9��=�j"ZH��6�Y�Iܝi���BK��O�S'p���b���۩K
�;�ڇ�?3�\��Mq]"���.=��"��������p��ō��g���i.�U�T�n��N�2�}�*�	TT�y�I(�_L�/�foX����P��z� 

4�	;��$�8���أL����R/}��Y������[��s����u`��-�ob���|������*r�����E��T^��r:�����"V=
��޸���J.�h�:�(&�*]b���C�[M�J�Z�Cn�
Ժ�j`6�b�P�������j�qd�Kx�������(�9N���zk����,
�ǕSP�]<y�a�b���ת?��0#I�O݆fkB���0i�o�L����6��V��ۼp`����Y��&��C�i���4Sn^����˘6����	�ku�~4p�@��!������_�70O/vM�/iX�q�-r�[Ϣc�D�ί����Z�'�@�����n�M.�9�4t����+qkN &�3j��}�U�h�(��kJ�q�H�v0R�)䎊�~�4c�oO{ f[x�	'�g]�9���@�NP���W�v��fdR�()��}��(�ࣳpّ�
L�M����&�y��DUC��I�E'������ǲ� �Ŗ�ҏ�-�)Y[����J��q[�Bh֦e��woˠ��q�'���:�~��^�@��&P�>�7��7A�
��`���/�DA�s���{ǹ݌�k_%�y����5�&B�k��Q�R]�]���<$���*;	��ݸ�o���M�������Jc|ìH�P�;T��f�8���/�,��k�M��0Ӱ��79��T��D���l�V]n1H<��;]��3��s�7���-a�Le�,��gTe|{Qʅ��;k���Gl�T�%k�p�\��[�x�(t�.1}Pb��\˦Õ��R̚G^�`cL׽twM��+H����Dd�]��@��$2;KnU�mw ��*3����^�����ʼ���#O�ؕ
�%�+=��mA�dy�5F�f�����ȶ��Ǖ��ߝ,>��Kn�e�Ԙp�5]��Iގ�1o��N�B��A�R�@fk׊���"�>�u�`ķ�
���~���JO<�h��e̞.������4u�G��e �0r���Dj���+��׽�&�|oM�e��]���^�s�����ss��o퇟7�V��
�(\�XЏ[�+Z�.�+�sJ�:z��O1�E��]����aֱ�	��ir#�,�g����3{�!T#�<����g{����!\[K헍8�-7���rH�Ɏ|o|��(j���]�f��͌���H"��#H�Z�9����#��+�Md����
��/[ĢW:-'4���<��E�yx��,\8�7�d�c/�IK�'�4�T��l-(��/SD�헂aS��L�5�
߶��o����F@&���AU6�ӾS��X�U!x{%�x��;�xj�Ñ��J��+./�xl��ҍ�&V��eNy�n::���}pYǅ���x�����D��R��ׇ��p_z�}�kP�l�"��'-@#j�DL��P�L�Ρ�i��g�b�����������b�ߖ�$��i���'��^�/+��>�����^������9]��˷24j�Y4�J�U���~V}�V���ٮ<h���"��@�!T��m�o�D!���� �Uޢ�y9�P�o��<�4������z��	�]T�+l�`펧<�>%����y)&��[Ź2M�O������9����ϡ"���r �R-\l������ؕ�? 4rο:}b�)+P�;�	/�"�W���&�A{t�vO>l_Ѣ�J���N��Ȥ�k7�,-QA��2=�&v�㒇w�tb**�|��b�M�?�jx Wz�~���pru]�%:�p���� k��h�Ѩ��*4 �Y;<hÙ�5h5�a����L�4�l`�)&�Ne�/�#33�J��ϥ�$K�5C;�z��\,�r�7�������`19%�C��њ�%%Ҷ��]ɮק�۳��u ���8y R�O^T�[��7 w�ﱗ�6D�t%��~Y�l������ۨ����B,��v̲7��$0IW�����<L��N�U���|��DS�3R��C�c��RXT_���╃�#��"���*ρ���t���4
)1V��픋��c��4��!\�]�R�Q9�����:zxήD���̣ ]ٌt����9��|���N��x�W��x �ߙdD��&س<�~�"rҁ�o|3r�vD��T�a�'1��x�#P�K�V3�YW�I^��]�I�%~O�����a�>�R�A�O'$)�ѐ����8)��?ߕ6[�9>q�PF��I�Z�}��َ=XR"�[`�;�6��'9�ّ�v(�`��	h�|gK�D��\�vA��؏2*����������+�e�� IV���?��ԐK6�~�\���?��P����:ў��e<�fho�R�6#��:��R.�3�9�οQ��,6��\�^��u�XЕ�>�ϰ����M���Nش��Bq^ *��*
tݍ�Y-�%mh�������oɂE	��	g�\�^�ͥ��ݩ8;Q�m�|si�z�HƉ��c+8��U0�6Q�Gz��ڮ�R7�F���D������8P��lC0$q�X����~��Xe�:�k�[�Zk�aJ�I�}9�Y�a"��Nr��rtcg(��Y�wb}�w���o�ObT,�Ϸ�gņ�3��嚠�Pc�<;u˗��h	��)�ͺ���&�p3%�9R����X,&S���y"�ض����h�?��7�|U�a
��	$]Ip"���=rjoL��w{Av=��z��=�f��'<&�}g�bN%���ѳ��Ɨ�j��" Lmr������]�,q��:ꆀ�c	��F����йez���i��C���~5����?�8}Ñ���+�O@�h�Jv
�{�0��P��S8q
����T��/L���e��_�"��Èɟ��(��@���}��kV�k����*)��2e���+�$�����&|���2�x6�W*@��9�<���I�"}IsS,��v��L���pM5��d�����1K�BŻ�#(~QO���uBy�3U�D��-��f�}#�~I���)�N�%�~C�Wrll���Q."��*�}<��ǫ��JG]��s"JEI~k��X������85�R\�I�Tk���8����V9���.�1HDLL��A�E)���K	���P��-_X�����
�0�M�M�K:�F�ɗ���Z���|���8��86(�+�Ă����3�z��p�f�K���m��$�U��C�e�f�$[
%��Ŭև�j!h�[�Sŧ�A*$C�<e�GW��u.��cҽ4:���m�W�1�l�k�.}2��"N�>�P�]�=����;061W�/L[v�P���_��s�z�ܻ.���R�9�[�З0e��'�iyp�q��,uﱫ��[%�^A��@w��p%�������D����a.�UM�K�q�0H���A�-V3�hc��f^t�F�����{�.�Ԇ�g���G�'��U�Q�--K� �%L�h���y�-Vr>I���͞\む�ܩ�^i���Q.5"���(���+�7Ů
��	Qe3�5G� P�u�
z�'{�\<f>�]������η�D�πpJ�"��[��U�eخs�^�+K|{do�� �7�nl�&I��m6E�+J"�`��������?b�m�J���F��^�K]jrJ�.aL�G:0���Cbh��"�� �����B|��\z֭Bĵ�22���V�V�G�}�pI���qS�פT�;v&��ߨ��Ȯ�5H�����qdu9Ԝ�3�9��`�=#��A�.>����.�Q	�i�����"�I��~��xo��_+��}�{�����ߊ��E���j���MS�����qK��>�_(�ci������n\6�;Ki�;#� �/��9���@����p�Gz{(xIn܏:�_zs����R+����=��X�j��Z���F�mo�_-2*���ԑ��]�	K�j��1�5��܌	�79\�"��W��>גH_�Q��dD?>U=wZj@JU{��j�������7%V*]@xf���A�h��xߤ������#l�ⴉY�=#���UI���cF
>����e��w�����<x�4�z�-;B;��CSb,{|�Ԁ��/�LOb�q�5��[y�&.Y*v�_��F�0���{�.��l
g4�Y�
fj�8�	�B,�r�p�����`�Ý�����̐�D�w;��/Q�~O��u*k�wh�O�S밳@0AЙ�{���i\A�r�!`Y��~"g�>�1��/��?�'�ϰii�J��I��@O��/��wo���8�=&r�� ���w�a�L驘���q5�%hdhi�V��^@���O��d&�k�;����#�3���`�����}��w��_����Srö�g�&~FG�j���:5o��g"U�`Leu��}��#cl����S5�{ء�����N�H$#\v��w�B/V,X��f=�@���NM�:��i��KRy��ҽ�n���8���
$�졍��5;��1e'�����/�q�� v�Rc����l��ǚFBGIT��=Y!�/��$�JW�=#�y2��_Ú���2���u���m��y 3��^|�p�`Ea��c��r��!�C�k��M�-�c���)���k�G���'���G<�ߴ�u�Iڹ���QA�%�E7�u�.��.뇐��L�G��%����5
�1�˥��qB���ha���Du��ݦ��K����:��̻�'��F���;������n��(�����N��������.ac͖3=�b-���z{�d@��52�<��<bA�/�(��A ��G��d�"_����/Vޱ�Gt���}�.l4���,����Fp0�\(����=�~��f�a\ՙ���rNܞnT��IحNH�r1��D%,X�!�jx�ى^҇�U���A}3�;$�|���$9o
��?"�������X�I
���%�րC*�%BК���}�U&����ٺ� �k��L!�D2����ee�`���>���mgV�2~�#J`2q|����@����jw�9�*�ԨM�=��_�ю}qa��c\'C˗y[��SC�#�L�_���2!�I��$�,��!��uU8�s�/hEc�؅�R�қ�3$��7�5��ߊ�O�l���q�/��b0�Ɉ�3�Iq̉
�^k ���<��Q�%S�|	��)� 3h��b�t]t��k��R�b�y�n���8T����^���k��9�!��G�&�������:[�L����ܗ"<��c�t䘧���_�Eb�NOpns���]ټ�96u4w���?�ɷ�<�d迯	|�܁�BMv����ʠ����x'~���H�������-_sds���㰽�>%PȤ�#8T[���@�IGe>I_W6���	�]��u/mz��F����xq�Y;H����5=�������t|���\ p�E�6�Jq�d�����k�J!TC����`:a2��*F��z��<��)�é�����?�:�:>Ʉ�:] �}���Ql]��2M�X�!JVh� vJ�~����G8�X����+��00_+�*��ϣ�����a=���?����Á���9OJv�ɻ��&I��<�uM���f��TB�)(�k���e��j�p_f��e笠�ɴU*(1�z|E�C�զ?¥��ǻɺ�1�<4:���הl��Q�(�Kv�
�f��r�T�HN=�զ+Ƀ�ef��qh���+�@l�����Cx�U�Oxz�Fƿt���V<�h�:�Y�� �й6�VӇ�p��U"4�<�R���!U�4Q�L��^	Ԋs(�t�5����|��K�����E���1���,��NiUrTQ墪���)���ۿ��*�qw�_ESӢT4ܗQ�Ou�T9]��ɢ��,";���B�6ѽ%��暉���-�Y*Yh��g`����o�K�{�J���_�I� aK������:d��M5"�+D��U;)-P�N��p�G�@�4���2@c\. �0�r�IJ0(p��χn�Ǝ�d�̷H&8�\��;���T� �E�2!��K]ZI#Ł���/�M�����U#����c��;�?�4M���E�ȁ:fR���s+��T�'���Q�=;[���Y��!$�{cT?�Ղ��u0�u��q��'I���x�]�]'���(�ޤ�7����[�ol
���=F�9"��Wj�ڀ��T�.k\x:� �G:���&��2�A�׺��i�M@�;��$�͑S���WA��b����Xě�@W������vsё��P��{������Rާ'HϜ���0jx�r;�3�²8+����H( EoK��|L8IF��<ȟ�O��y�ϫ;����q����/t)��c�E$oSPo���Ρn�z��g������+���l;�OI5���6! HuG,�����W)�����rz �d�Ǎ3ԕE��>�q�.��P/t	F�1�BcH��Z���+(������fR���X���>s���l,�Z3����e_�ǸQ������+:�l���7U�b���W�'V�Q��� -��Ξ��bz����ޛE5WC�pq��6NC���4��-#"��B,jI��*I�3�#�  ��ډ'b����kn,���e�7Q��a�C���������)�S��.� b����"��ᵚ�&����7KQ݇	�B.6[�E6Jݟ$�/�F�SjБ˶�CD[>�E���2ֈk�A'޼��������0I	5R<��<v5���-�.���b����pwE5�>�|���>񓭖#^�jpo|;qYmR�@�J�ki��ў��$��E�����2���L6d6�_Y8KJxGhe��f�[ϔi	9��T��?l��^����|��<I+���At���"+5�l[���7�kk�I�Y��r��6P��:�W�$M�mǚ��4�}�-Ə�N�Kl�#�W��(�ը*�E�*���~z���u@͜��f CU��-G��G�U�|���/(�wʇ*�b��!��E��}^@T^�� ��P>״P��XyF��K����YZ!2�kS�.���'�\@љ�k=Q�e�D�Na�f���զ�d�%_03K�F����Y�O��W\�d�Q㖄�/� CK:tO^Ȕ�^�p����w��`
j'�E�/.�<V�<����������KR�����T�d�g�R8o{05A�w��~#�n��2�R�.�W1N���2?z�Z�J�QDw�^���wG{��<Xa�� l�߀�� �ک�XĜ��r������]���[��A��~g-+S�s)����F�Hf>s���7���_�e��M� U�|�)��id��^�D���`�Pn��6���5v���}��%��z<͡&�������
j89���~��]�@�?Ѹ!�A�IIm�FM6�W���<��=�{�� �&~�?O�}~� А��dd|a���i=9����;X�sa��cj����R��`��z`ZJ�9�N�f������1N�]������?���}N��
�b���m@�f~�7��,<>J��<�4O�̙z"3a݋���nx�WЃ=��?BUz�	�8-`%�FmbPL����4$Nx	>�K�d���(�a�Q5����Xȷ\/aQ)P�̳�(4潧1c9�Ɇ��+�u�n���%@���Z�
�g� �3��z�����e_BY*�1�3��QM���!�G<O�V�?�:y&]�o��19�Ɍ��5eN6������3r�tOOب�ݐ'�gg浱g:���.x�䱳�G�����u����PU�A���xg�����Hg#�'��^�dn+`����%}A�?Y�N�w[��'�<(ֵe�@J/��N���//��A��my��&��@�~#�ڌb�&�N[J'�t5��Q�¦��F���~@�Z2;�7}3%K����k�[<{8��aN���=�LU\�>���>=t(Kk#GS'�*(f����~�4�y@iy�p,O���%9�t.RwY�ˡ.#�!#�f�Jݎ��ύ����^�;���ݐh~/kghC,�!屼����,RD����<N�n)��ER:�G�v�,�7���>��+�{�j�ɤ���a��\�|��	�FJ�v���N������F�d���;b11ɫ���T��[y6�ހ;:�/Q�nGfs���v���?�]��T<HS�V}���zn�Ce�>QD!o�(������!��f]�J���b�����{��2��p��d�r[��a�vb���U[yZu���	�y�����d��v'��i8��7Jۗ+)a��9�X��C�$~J�����Ą�.���qQko��5L�p`���P�c֣P��v⡪tj����wm02��g�%Y���uM(K��$
�8�t�������`�0�$5���T�e��'�D)Ϸ 0Zg�B~t�.�0�.Rf�X�
S��)��h+ئKSV����K�I&�.�"@�~����O��37�ꠎ��3�`��(/��̇����^ �b���(�^M;����C���Fi���͍�ymM�1���9��JD��$�b=�i����+�M�[�C�Wg��,o��5���!�S8��~[*�(�ݖ �\�2'�~rڛC�D]e9ba6���Er~��:���� ;K�!��}�����$��ևhzM��'�V>R�d>�wP����>#%5?������/��e�O�-�K����g�E��T@�0'$�" :�d��*��&�_�ȷi������h@>�3P����k ����0���l3~wK�q+a)eI����S�Zx𛨤�("�JM)�
T?��K���y�}}�}�9xl1���q���EVj��~a>e�$&�k6R�-:�"��S�j�aR<�z2t����1 ����#!K�٨h2\�Ӿ�:j�t���\T��(X\�F���s(+��ߍ���Tƥ�aI�[R4h&���km���Ìl�L?1)�� ���ė�}�z��A�N^Q�-���YN*��e8]��"2F�GM�n�4�(ᛶ|�آ]s}tvW����1�D?@8�me���[4?+��~��B��MF��rY9��,�"5���J��rYVS:�.霬o�?\1Z��b�7�R�=2�W���s���Р'��3�݀ fM��̣흙iiJ���r��n]O�;�=�ӣ���Hg�]��N �~S�"[yK*o�Qd*A!q�@�u�����-��Y;�$���;���{�� '����b�醂�"3i�۵I���6��P�Ty(��@�X�|�X�Ut���"�x�O�k���R�q���A�i{Ę%V��7�`W|=��>z�F� �R��v�"yd��6h�.r�����	$�2|�}"��������bz�ɗ.�͝���1��ٺt���4���1x��v��OF�0ɒ3"�=cG�(^ ���$�1P�A�+|sb���wO�k�$�R�2���L��Z|b�;��9s�^�44�4M��,���!��,���e�:��N_�b���(��w"2���'�Gk �J�x�&��'EI[\�( �;�$�� ��T��l`r�*��;�3�4^����P�n�>�<�9:�VƩ���G��?0H�~��XH17�VE��L0>�m�$����j� �)���3u�^�l*
��G��Kqvm
�O6heX�c2=}&��
�Di"�nSZ�� ���L_Jv���f-a�$b�fg,��Wt?
{&���A��k���:z�J�v��O�ܨ�E7� )��)�K�������0Q�����o���y�ڹ��%lG�s¤�>$���ar��W>'��g0���P;��7�`n��pT���=+S�%hM�H lB�n��>UI�c �����۾����0���h'n�0Kkж`Υ;+<�{�v��v󻇭�;�����i)�ؓ}m����,��
��`�x�Ě[}[uo;nv�]��$��<=�Q���YF�ȸb�S�o�(oAK�W!���Z�����E����ڏV����WxX���[cۓ��2���ʟM�-ݔ��1c�
!D0�Yek4�����X�U�t��>ґS�F=�1�i���%lͬ�Q=$�9�M�E�O��>7�L� MI(�����@�sN;�����! }G�Ֆ�]&+��*����6ùt��n0Q������H���N쌂T���᠈�~P�r@�����V��oF������B웹0fY��U�)�.�b��`��b�����SC�l�[�e�r���ʛbF�t�.J��+�?cZr��v#��G� ����
���B C&�X\YJ���т_A�<�\����\�b6�h�����(��2��>|��h�	�����m$�-f#↜+,e�2���怰�c��v8�D֤|֫�I�#Eiq�����Q4�}��G�F-Ĭ�W3w^��@Ap&V�j��ֱ:�lGIE�h�/��9<62�5�;N�����s�0�����m�K3�մ
�������,�*�	/�TY`�]+Q���d���vt~Mk���OUb�@>+G;�@nf6�4]E`Y}�9�����OI�9���i�f
�&HYvW3��s������fQ�-��:7!�y��bM���F�x6cb��B���{�n鷶Ld#��~�/Aj���_�a ����0cӦw#*����߬�P�E��k����#O��Q��GaJZdY�wG������>b��n��4=«���@2��6Cv�����󖍔'�Ck��$g��B�ȣ��JD����ɹ�~����ZM`�Z�a���\)���W�J}�ϔja=;-�/L���	��@$o��'�T���g\�z�#�kj8�5��#�è1p����7:��E�������a�!{Dza˔�����d��Yu�z]�J_�����xe�/�KD����AN'����=@3o��rp���tK�3r%�jj��������V���������	D�'1�v>�Z�I6���ats���^�R���=�L(��`/�+E��2<�&`R�yc?���E��:WP���H&p5�J���IH3	�
���H�p�b5��./�|�T@e�� IYCtB{�����'�P\2S�`��_o��ɉ��Yn��_K�t��D) �b"gQ�ЬM���Zd�&�tŇ���i��T���bq��N����uv ��V�Y��X���Ƅ%��Kӆ�UE3R�Q�Z�>EZ9[BJ����?��A�td������L�:!��M=���֎����?"��՘%l6�\20��#
�,���X]R�*�{fby�>�UP��Z!]>�x����PN��Pע��؟$Gj��]����Iy�� u��AZ2��]aE�W�w���et��\^��_��:@�{�c���x��T"6=Z%�KCE��Ӿ1R NA�k=f��[(�~��wL0�1��w8B�WVh��Ui`�界`��"�����<ࡍOz�IQ�%A���|�Z�2�6wꎞ�����k<�A���C0��FX�yUm%wF�)qK\�s�|��,՛�I�]��]~Ч��{����S�R���+#�ן=r4籇Bw���O
��c�=D��p����7��i����'�W��z��H�0��gN-@�%�_��)�Py���m~Ṳc>6�����:=���&�2}Z���n�����^�H��1���`�<��9�N�X}{G
y���L~ق	��uM��V��4˭L5&d/�k^"gۙ-*o4���21��X9&ȴ`�@W��z��ȉ�G�C0f�'�]��-����Ke�i�;:�s�(������TJ̞��'�6������
x�o@��5�7,S��$�ˬ�����I,�t��Yq@�p{�M�� 	9���#=$'H����I͞��M���խ����O9��e���^�"�qV��4��Č�H��"���Ve���v7�ZӃ�����" `2��	 ��-�K�Z�y�x<O��hX�X�nvk.��S��Y>���Q�)6A&������eLt�K9lԃ��	��H��_Vʆl�;�R�K	�E�8��DE՗�D7;P�-���A���	o�ҸՠYz�s]2]�:Y��d��b��#�t��߈�E `��6�w�q��������@�v�n&q��L���G��6X�-><��ܤ�@X&����P��zC��Ǫ�:qv�SV�Rx�B�8<%d��I0*����0�Ʌ5[�v5eۃ)�����Д���M(w �6�wآ�7���
kk���M[��-���m�����i�.dǔ�t0b���ú]�{�*�M�9������Vq�l��&�l���8ŀw��t\Q��w�2���@{I	]�Tt��wL�b�;_���l��tS�>�/�%K)� }�����Dami��6a6@����õ�]���n�D��c��#����k�)68W�$���Q�&i� W�X1��8T�%ޜ�xFp��lD�,�,���l�T{����;7���p3ŕ��_����`�z��=�q��!�b\%ω:��è��D�0ۣp@��QC��/��@��/i֘?��
�â�F��!E5��*6�k3,tL�T�웫���AJ}U�^�A>�����Gؗ��i�E�H�����*0��e�A(9�����3|��r'/�x7i�
�$6Q��3��h&&[�XjS�Ī���l�=�yU��װ� ����S'�q��	������]���4�RxG��+����E�玶��C��{iw�ʚXR(㪰x#!�O4�m�$�� 0r#��9��C�k1K��R��ل�0�-�k �G��IQ�r˥�.zX��z�S�N�G��M�&J�2�
[��svv�lVMY'��E���R\����9%8�q��������Ǽ��_a�K�2!�]Q���醵���V��a�v���=��=�?+¥%�u����?����	��<���x������W�_$u�:wW�6 Br�y�~�����&�v��q9�?���-t����KTs`m���k�Qk.>|��
�
�f�@���&�}�bj�.q�	�3G;X�2�?:����Pй�O��j�57L�DL^�z��Ⱦ�,6N�r��Wy��)��	g����%r=*0��� ^�bW�]�Z|}��ɢ��R�+Z�0������~f�Q>s��N����'[6�}\1e�=�7�T��&�5���'�՘�",��/SrT�3�V�?�ʘ�����\
�3��a1N�cS)g���O4�ȡV�q���T��!�m��s��f�_���Z&��&:�FHK�H��x	�OK���"��5}2�bJq��������y�^����B�?4���'��]�ƀo�� ����j�[�#M+��c��6�2�Ked�욻Z�N1��AJF�0 r�	\㽆�@r��V����l׹�}�d���UD�p/Gժe��h����0>.�+S��A=VP5�+Ze$��a!��Д��z~���j����x� �2?�jm[�������I{��1&���<��M��������/6k��q����"����� Y��M�"��z_]窣�i����c�~��"g��֩�A5p����4��} �k����>���`�@���#4��ɺ�C]��S��m��L�������/�ʓBF��[�Og�D��L�x��FD��S���2��:9X�f8�N���բԐx��W�
�o�C�(g�HT�SuP��V�pIMDb!�'ٳ�v����t�EU��b�P�1��̇�+��7���k5�Sנ�F�2��ª��C�p,Um�6�E�B�t�';��C4I���L-$g�{=J�q�W�Wx���l1�7��_����DZ��-rū���������|d¦��ћ
�����~`���O!�$��&o��@���M��e�z�z0%����֙Z��;U0w��m$(߫Γ��hqu-E�n�g]�
�F��J���naP��Νxh��)2fOFy��;qvhB1�C��pM^E�z癸H�,h��g�'��4�e�����$e��J{�qBB�;yݺ��<H��eT�4�C-ݖ-R܉��Vr8G_zPc�?ZS<�B�������������BĴ�U�p����.ה]�Si{]����,��{u	�j���[7����e�4�����ˆj4��}���l����E��'�L�u��+�J���i�W.�p�,�-r~0�F8�u�@��I�F������(�r�,9C�Yz���0��`Q^�X��q�cc�(��D���~)o���r�2�C!o>�3�#�]�@OV�ꄴ���x���n��8��:%�f�.�O��d�brreJ�
�a4I �kv}H�q��E���s��� _�VC��1�yv/1$�f�I���Q�s�C�Hؤ^�+��.�O<��(��t0'�X�4�]�.�A���2��k������.r��b���nlI3��HZ��T����>�T�H�	;^��8�_�07s�c�Ӥ�g�:
k�D�\�|���L��{��L��|�4��Ј%";���*��!��DA`4ۥ��~4�j#~�%\h�&�gb���b�[�M�fY��/��>rW �Q��9p���n��V�N1	j���-��:�K`���t�a̟hr3,�z��><h�x_m5+஽��m2%Y����ttQ�(�1��rs��\Kc��B����'$j ?�Uj	pve=�F�u[�d���@C��'�VJ�A�~mI�ʶ�+*��r씨�:���FhdLa��Y��
�G��G���5L�v|C㊥�t�<=e��>!w��'C�D82 k�e<���ݸ��)_���vŰt䄃��LJ;�]N��v�y5ol���)�Q<�Qo���G`;2�h���r��:7R${�g�O����z[I(��%!x���%W����v��2�Z'�	�`j���T2z��a�Tf�\կ�2d=����n��6�"�K����T���?LOr��ṍ� }ǥҎ��&��fP��ѷݛ�ᰜ7/�s͓@�O<)�T�e��P����o���9n�81r=��0>�67[15��H��;��/g���C(�؁KY{{�H�,�A��F~@�J��W���l��c����L��Ң2���AgYвq��!���m�i}k�4W��ً�����O�Ϸ٪��q�C�Vh3�X�F7uSE���؂v�(�N��]M]�x"�ۉ�߇d�죭������lŲÊ�U�=~}������~��Ԙ�F�����>M��F��V<��S�ilS�%�?8��e����d�fY�݌�u�*؄n�=�
&��8P�%���z��>��p4ɓ���D�&EWaWN��Ƙ7��`@���GZ@��0*-7����@�DZM�q%�./x�ջ��C.e�+��{_�c��p.b�E0�1"��-�l}����A!O�{�N�0[i=]�2������,�N?=B��j�9�pj�..~���1?�iq��p�a�?�r5�fmK��C��� �*>�/���^���x�htew�
g��W�?�{cѧ�^�/c�d�SH�:�2�-��Ʉ#h5��]���ݏ8Ș��p�C�3�������Oe��%]�6�%J�f��G�e�(�SwAG/F����ͨ�1�|�4|�/�����"9��kzҶ|�#mcz���-=�c̯_�d	�����h[_����5�zbh����ʁ�����3x6ǚm}[�3"n;�]��~��ۊ��w~5=����[`M�;�\A���zӽ��"l5���eD��a��A�*�f��b���ǯ�
�/��Cu^YrR.s�R7�X
vb�1jSWwZ+�Zߑ�+"���R/��^�)�Rݟ�΍kE�f�)�������A��BB�\���B���e-��f�%�^Fg즉ձ�Ƒ�$�j���$<�K���^ɋ��.�i�����ڑ����4o��㘾��=0t�R��d��
�J�����x4�v��05���;��i��Ok�H`:W7ФI�.M����"�h��Q�;O)��36:@�rt9?��P�J$NK�C�
�^GN藽�ĨF9q�����	9�v3��D����+z��V���Y�H�/u���q�v!����WfR@�k���v��D.^�Ai�pie��l>�SD��\w2:>���x�I;ė
(D�*T�TS�d�<!��`�EՂi	�Ӷo ���c���s�K;mC�>?/5EA^~Q6���Ȑ�os�u�5���߻�`��E�T���ͩ$V�ь�n�v�#��O(�őE�������V��~b	���Q���,��b��O�(�����o���]�����	�Uo	��9B��E�7*gn�HI�$�j�	����� ���}�#n��B�Ys��pR���X���:�����'���bL�n�����:V׎>f���
��g�zt��n�z`���	mF�_��-
c��z6���s�_�����.[��dy�G�I���+u�*+ ��FE�s�'��P��A�Lo���r�)�*Bp�3H�Ũ��H1GR�ּ��r��0vƞ�*�5����� L�d=�=c��`T�[b�T �3GH�߹�^*�cjX�e�k+mm�8�Z.O�QJ���{���Irܫ4��`�B�>���`C~{$'	��XmG�lSA�O�d3�x���r��a�sk�b[H]V��|����|��n{�}��lz��tX��n���@.I�Gb�%db/����{���"����=�AZ����O��Ζ�
cs?k�O�.�I�V
��\E��k�ګډWE�S��Ǐ�"�Q���xB$��w�k��yih��D��9\*��VJ�=l=u�Մ�| �&��@H挹���[��ok2V{��(�j�����Y�����o)U�]����]G&X�eq7�tӏ�)R��V514V�/�X�U��G�K���Z�Y�v�?�	?n��G�1K0~W�7���{��3�r]�/ո��g�,L�
c9���/���\��A��[v
�۶ɦ�֭�9�zX^ʥ���a1�| P�ɢlu!�N�,%T	(?�� ��Ȭ8�æ�l�ā�po����}O�xHW�Y�?u����j�2���.ߤ��lyVc&�$����h��Yt�g	�Z8P��]E��ej�lw[� �s�ջ�10��i�ޔW����9/E=�Lﾈ��e���dg��j�aG��:^j#�`g;�$*�G��2<zF��=��+S�7���U���`�B���
��HJ��$��ss�Q��Ջn�y�<-�;�Da�
�	��9��k@�萘 �S�X`\�u�L�ʉ|�Uw���goD�Ƙ!>��ī��^��, _�K�kK����§2�f�I�=����D׵�\_)�iu"�<PM�ܽR�]�^�"��ҝٹ-�X��o-=�-�lZ<3J�sL9I�4*��j�R `���m]��������g�\�4r<~Km�i�(mpI��H���$+c�+M*�)A�Aʿ��)��g-яJۦ���e�����i���	�{��ŉ�ÔִMbr������{�����d����B�U�V��س�YGl�����y�1�<�����1?xϊ:�O��xe�M��#
�t=`�[��N�z�',��2�@�K~���$������ܺ��AQN
^��l���f��Ί[+�������Z�1N�Q�ưN���h�Q�R�WП��*�0f�k�GZj���Y�G>��,m_nׇ�%̜ YSDDћACM���u�0��{1��>CM�t�K�D}��9B�������j�5[��ѽ҈��"9%��|!]L 	�ǹ>�jS���
�5�>p[s'l �u������b�d]{�b<����y�8�F��x���w�(4x>^v�9fg�ХK�Lh����Y�뉾=ٯ�>d��߂�c����`�ŝ�X��F�+�mA����,�Dݧt�Z�꽖�c��*Gz�C����������� Kh��E7�kof��5o����abFR�Ip��A��SP\��<�M��=E��K�+�S����礧Ծ�XG��-���zy珗#�,�*+����L2��2EP���"P�iEe�q͹��N9�%��H+

(%iD&S-���jP�l��XW�E�₡���]7�^���Ń�nRM��z�����Z44�qP3��	F7r<H��"~X���W��]��#��.����3�8�
O�
2�ۺ�>퐭�{M�W��ޟ�ӧq>)������2����n��"9�L�Ȋ�*�1|#�R�z*2-��,鱗B��E�¥�9;n�=�%Ld,��1�5�}c8�I����љ�C��Qpv��4G�#wA��t�X!ɵ��W�c@��߇���ƃ�~��*Snxm��@�䵫�J���������&v"�@�n���A.$)�����/�~��������R�U����O�k���T`�Cw�<�\���]h�0}��"�*��)f� �p�d-��.��i3���m�WY����#������������+1I�F�tB{[�H.�0��Z8"��*�@	���d=t%P�h����)��+~'7g���l1�{��ʩ�7�Q\?t$��Bg�Z��q?uraH�_h�b�#�&/��i��|4<�,��!ƼXw��,�Z=1[fI*zS���+}9�Lh�T%W���H����ޯN�����L��'��b��ƆaZ69r��g����"�ѧh]�?���qO��NE��9�� �	��g��8��L���]���� �<�{=�.��'��{PR��\�[�8��J��a�#,��ȊN�9�&B�=?����-B��Rꕘ��~6�;b
�9*��S3���dvй�u$̀8~�׾�[�,1�t�[3�b�Lp[��NU��L�z����x,o蟄�,	�N�z��Vd��y/�͒߾����["�����s��tZ<�Z�NUv���ժ�t"w�[����My�5`b�j��^{�N��l��[y}ZC���s��j�h��C�����p��I�y��mi��a#��C���5T!J�M��Km'~聺Q_\�G�~&�h��⨑@�:���� ���u���0C��G����5Q��Db_H��0㶏���WREp��	Q�p��y�� �Ee�u���/M��^�$��DC�2��F@��4)I�ąw�ɣU��56��L��B$?���{x��'ߌd~o�ӫ� �p�A��!�� ��;c�dZ���e��m����G��9p֫s�	��
8���h�˃�pa-����!�G��i�a�r=8ՐW��;x̡���ήz����0����ԋ��&���'��}6؈F>2i�<݄�I��4����64�ۺx=#a�`#��{H���a>B&�6V�2���b��x�����d!�&��x�饭7Q�(B�(2�քooF�tG3���0��;�� ٨(�ځ�����
uA�����R��x�?�X�3�K�7X�dY�Ħ.�X������OK��'�����⺦�! Of����vٲ���N T�\�-І�-p�����;�ڳ�X�}n0/��'	vK60#�փ
���������Er)�^}���L�������c�6U��������~)
�������a@T�S�`T3\��o�e�'������:�Ar�Z��K�/��"�'Y��3�"�L�lJv�<��1��v�l�@�-n|0��Q��~Ja��q��5%�T���0W���
oO���2��N� ���E���]���g�T��e�A%�z�N/%�j��Az6��\���p�!�?��&Qrj\m����,ŋ�"(*�an#s"�];ݨ�5�|%i��k�Y6������r�-y�H#`������:u�?Я�84\��	8|?5��tRa}���Q����])� `��+��S&���i"�]kh�'�.����)yӰ��ե�B�9��ֿ5��M�9}�ѓ��x�� ��煩Zט����^�EAU+��"Dӂf�ƶٌif "l�$cn?�&I�Ŭ-7?��ƸL ,�4�x��ǧ�Zz������ʆ���4��U��B�� ��#�đ��~�]J��� � �/�͇�6ԭ�:>�/6��=�%w�����G�tT�``xbw�D�
0��� Үr<j��)�	�V�STw%x ٓV���pqq�$��!M�`�6�[����h�2>���>H��dD�� a���B��Q�^FL��c��!�k��
k��=�����k�A�nhp�����R���Ӣs���V\����W:��H�(�����U�lzr�UK��f���aG�{�=��n�u��u	�c1V�Ap�9�,�U�VHxȵ�H.2ox풒VWND�[���<�w~�վz�N �TQ;����T�YX[�|K�M	���s/�؃��hԚ�QD�~B�bO!ٗ����Ĩ��$�)�n6Q�&í
VJ���Gr.�уO>�]�Oq"x�x�=V���$�򵡮��k'å��]˯!O'C16�
 ?\X��0�{��]]�Jޭ����aE��w�����[K�Ԛ�F��sl &_��>B.�܃�pX,hIS�;L�7i��G0[�-��U�_f<�����M���P�3��-{ڌ���3���`%��¹:'�j�#f4�q����7p��:]������V���Ɩ����,��>ӄ|�&E�Ѥ�����
~�:fW���u=S.�s�/�7���Ŕ˴f3^�9!��:�ʒڮm����hY���G�O���rU=";>`L��"�˺�X��!A�Y����V�ou�I�2L
�����/1(�V�B���%}Ǚ`�d��}��͈�S��M#��Yމ����<�`4��WZ"�_���=���3*vG�ʙ�o�����lY��@�=U�{��,v_�Wc_��bZ�\�{������ؽ�5eY�&��4vJw��~�ن�Х�lM��f�ڋM��}��/����G(�@̽b��oɳ*�~A�c�ע�����OD���4�:6�\���݀p��ۋĥ��y����*t��v$�wx\�R�A��%k��>���9���δ8u�(�+�2̙P*�1l����
�/�O3S.%��
��!^���7졽3�1(���M�>���ݴ]�y}D�!�5��̲*��<�<���T���aJ�©8e��y��]�%C{c�%�"�>�ʦ���U�7��S=������3CfY�oOD�j<iVD(�"!�Z�-� KC,�g���>��!��2���B7}����a���9�$�.1��h����
�����w��ja`�����A&��zH|�Q<��h�A���H�9���	�Q�U-\t��#s �_������˅���q�6ECZ:��7B�������}*��� $������0��|aI�i_��խ�V�VA�}�x�����t�"qL�}s,��N�˯]z.z#,�?�GBn0a�Sx�`,gM�m�=�Ʋ�~�h�m�+*YM�����دOɦW~gn��X��C�әwm��=S�������9�@"� $kF�]h��ǌ�H[ 6�Ym飫Nݽ1}kZ�rJV�at�@�TcC(=�G��3�D��� o�r�{�+2^���$	Y�zas+����k"�rb��]#(yC�jz$����Q�{3�!�T��!�����h��ր�0�^"�S�6�Q�`�4Wc�Ý��[�˃�4dI��T~uV��q4b!�`��Nj�/S��L�[���?'ĩ�=y��%r���P&/>���:�Gzv���������}�ժ�{��0*P*��|����U)�AL�h�!.p��F_tm��#��]��E&[u���|*�!�������1&bj]��T<�m�;cn�R�aȽ��|)Q�=To��8���i��;�by������@|���ԭ�`_�1�q��5'爏�>wnG|������s>����N63o2z8v���EL)��j�$���x墾���/�k��A���d΁�9@I�O��g(�<��4���BF�����h0,�zte�)6rA�2M�-�R~$L�tTI4ͬ��#tfNH��I�m���;��^����z�B��?l�ݳS��W껓�&�D�G76��*�ǼF���t���I����C�p�|=m"˽�[4˴�*?�����AT'�C�(3��lhV�Y��=C�M٭~$:I�3�рKSN�����Ț l� v�ʎ:\o�'kUn���R����d����Z Yt�0����e��%WA��D��j���}��c�"+�K8$!�#�}�kQ&>��'h�~ʳ�YF�rg����L���$i�#;ߧ+E�{�%e?_^��%#;0���Αj风��*��(�v�h�Q��~�wn~�̅W�D_��1�O���MҺ9ǰ�Wo)�ۦtz&(Q����e��ۣ��v%��\��M£�_)�q�KNb��ݑ?�;����@����"�Fn�������a+ГA����$ ���7nhy�yՐ�M2��2�ʝh�U���a~�UF��K��}�"�a�S��3Rߣv_��s�i��Md�"O��rl/��Ium�ED�i۔~v]w]'��e��`+#�Ӡ7�M �����3�#��=��R�G�F�~��|�[���N~������36�q"�V`o#�ǒf�����5h	=.�M��ԑ`��>�N�W�F&�
m&�=4�'ئ�o��g��Z�
?'��Q�Xd���;x8%��� ��\��=¨�kQ.#1���\$*ʼ���B'|tYL�2���^�ѻ>����5J�k�yϊ���};�;��	��72]�eê�+��.2lB*bR���oW�a:�r�Q�"+�l�8ڦb#�R�k��cA�7Mģ�*�:��8�ם8�<6�1�`ퟃ��n��bvO��gݽ����I��l���6bbe��6��;�\���ݲN���!��Ѝgg��^"�\���m*"�E���_�p���!�v��0 ���4|Qa�;Tڪ�W1�Gz�޸��R�pCC���� 4\$��4�{��k�?u�#8Oɱ�y�FkGM\P{+q��Q�7z�9�lu�<�?c��i�,�z��Ai�����y�U购�~G]�L'�C�"0
���ѱA���mO��z17g?�+��� L��e�P2���n~����V��[����>������=�Ŭ�e����NfM2X��c����V%�ҽ�������ٳ+�� c�*�+�d���L�����^o�u[�1x�%�js��NPo��b�_cj`�DƫU'/�Q�u�d��f꥽U;C�G��� *���O�ז��Vh��uk�=�M�L"�F��[�9J��o%�a�Z����Jb/s,U���0���6V�GrJX~���f|��O�͛��T,$����]	�p}�<�ջ�V�ߖ:����ep���|j���GUVTϊ`Ѻ�ȝGd�tO�SGe��[��'s"��lh�RҘ#����?r���W��J�)���$oq���z&h�F����1����Dpx����Y;�K��������D��I\��u�i[V�A��=����b`W^$�� ��!4�8C���0�<3�}kM�Z���e���b��(�G����{q���Q(�2�.��J���gv1�O��^�ϓ�pE_��]��`C��PND�N�^�jY˓�iՙ0�g�L����E�dnOƈ��A-�U������BܒdO���N+���>�P�<��5�<�x]�ڔ���6��r����X���w�S�Y�Yܙ]���P__�U��%n�\���8aKw?@:G���k���ٖE_-����(������d-2��LN:�45�_��S }3��_�Y��+�vj�&al{����{����"�꒏�<�]S1��������z��f;	���\��7�/Bph	��S��o��QHoi<0��"��%�ĩ� 4�����@їp�Dn��o����r����������OF*������ܡ�L�����BL(-PCi<M����@f�^-KO,�q5�q՛�{�M�m����N�)#l7M���-���A�+�k���2i55a4�%��:�~b����	����,��E�3��i�B� �jaXZ������\;���A��Q�3����x���'߆�\w�V�YuJ\x�R; _q���-�bq<U�o9���y �sL� �󾙈�*�F�;��2�����L�����`I����9,�v���M�]�����f[�z�|N���~�e���1j�z����<�o��B�|ԉ�\�z��N�
�0}�5�5�7�qN����2i��A�̤�y$�9�_Q3E�J<����AcM	�4gE����q��:�Q��.��!�*���>0.�[�N_�K�|O�{��c�w���׊j�_>Θ,��F�S&�� ĸ���D_��;qW�Y�u� �:{��>�g�`N��3I���'�n".5�P]�� /�~*������"��K��H��e�\?:�@OHa� y?�;��t�{f�@���������E�f��P�=m��Ȝ���Ԉ�?�54�±�>��꤈)YO6�~�Wm�w�r3S�^c���Hj�h�>�ڒ3V���A���Xu�]�N�;���wɳp�k3Ӿ�]/����5�_�9:�����|�ѐxVcO�|��3^�e�!��Y�����f��@��]M���@��q�;�}�?7	E>u�3�fpW�C]� �8�g���-���o0��~�Ǝ��+�q���R�%g_r��$૔Yk:zdL�����W�Jt8�K�q�~���2�0���1۱T�]_����F�U��@�:��6#�����z���^�v������=�E�{�)�5��Ћ�ͮiۓg���������-�ƛ��a���;/a�b���Q�J
�M�&j���Te���Hɨܵ^6Z���:x&$�M!����h�HF�ɸ]ˁ��;���rM>x�-"�P`N��!]�JJ\�b�m,ʴ���NW��ɧ��]Cw����mчƨB��#(�K/!H#T,�y�A��3+�5N����<�p����O�4�.C��I���Vz��1U���3��,��be]�*m)������x�ϲ����'9�Z���I��wy�o�����w�{f��h�(��)M���WåqF�Ǫ��p�+Q����[ԎO�X8���^��:��K�o�Q��Q�4���Q�K�f�S zjS8i����"�-�T�n�U�v=C�9���o,I�Nw� m!��n�V|�:�0Y=.Ƙ���X�S|��؋�@ ���)G�xc�����V�>�NϫD�_g�-U�Od��&n��o_�Xą�# {[�,p�м���%����b�%�#��@_,����b.��T�k�2?�(�a���3�8��\�������8�*����!��>�N0ݖ�!��7�P�]�o�E�6�H&~s�U��%�f�� Y7V�.%���H�<i4���f�T�vᙋ�$�,ba WU���j�� �X>�����I����
Y��eqaE����5Xr3�ɩ�D,7��8�	_� ������z6G�qi�gqr���{C]g�kr������B8	���tdSCA8�0�UioY��D��"�1��<;O����Hl+��aڋ��.���׊�c}����}����/T��-'�����J;�GSX�'�E��<�=�I$8-*|`I��Ux�6� ";jb�
E��hc����Cq���a9(���#���Y�u�u�C�mET���f��ݶ�mSI278q?���� ��z�k���
���[�̹$U��t�p�C�������P�ћ����@a���c�ނ`a�����(=t��J��qf����6��3��;j�[���+̂����oa�w@\&�w�5�Ag��[�n"Q��3DPJ����uـs�p3���z#͓k�^������Fht=Z�UR#	�l&,�=�;�/��oB����`���JN������>"�����e	&���D#���#�볧��@���5��J.|��ʼ�O���*R�श#8��3����!d��E���y^��BL����R�n~���L^y��4��Q�xQ��qZ."Wͺ4z	2�<zk�� x�1�>]�و�`��IH�혙Q �<���:��YV�i�'�ڰ�:�~{�P�_W�'kͰ[��2��"rߠ���Nz˧_~RbRx4�M/�!ܾ"��!F��.�.5�&�do+r	�{�un-�r&�A�u2�]�3�X�&^�S��{��QhǨ��+�I�����g�[C�j4q2��j���0J/8M�j�7�om>��`B/-�{O�5��7����M�n¸�.
n�����4����ͧ����6kme߆юT�I{�OY�?�[l�3��UYu�4q��_������..��I�`�*0��~ƙr�?�%��d֎}�^]��詖����K����Q��jr��^Cє�ߦo��ˢ���l:d[�x��Ż(h���;��3>2׷�l۾|��r��IpZhH�&��s��Z~<�Pj88&Ï���/U,�6l]��b��BJr����;&+h{Z_����7�v�0��>�ba�0]A=Y��s�A6��h�J����#VE\ߛl��F�z�t&���Gd����[������3�z��ڑ�u�M:��y�ў���/�SQ5&Kg/g��x�%��<��$FI	#�<#g<���m>�,����c�
&��-1Ѥ~�O���Yd��mNl,j�8ȓ�f����H?�V������]�p�HL]��p��Q �8���{�>3Hޅ& x8�NQO�
t�eѾ���'5���R�J�sYq)���U�"����K ��obd�9N�i�d;O	�|B����'����)]q�C�m~�<����#|>��l/2\���2��-׫~=����bp f[�2��݋���dq��T���)I9"3 ��|�"�+�])e.�a36�,vZ����-�{�Rg5�(Hp��n&��V���M�UyQ`��E��n�æ�߭2��b�Se�?��B�\y�B�u������D3&$����(�I��׵ޔ�\�+�:/G2���z��zc7�tU|>6X\���ǻw�1Ìbj�2����ᦫ�����_�2 F�8�k🛬,/:�6o�x<u=Ϧ#FU@��^�K#tL�,U��<��mT8B��<���`u>W���̳�X��f:�N�Bw�؉%�^%�9��`+~Ӧ�YӰ�!d`���N�s�F�5�5�� �_3�����A,�`��eH$R�&�ʛ5?8�@������C�P��)�2Y�3F�J-��hw ��3p���û�}+'kFsD1Hs�Ĳ:-ҫ����~�~~� �\�!���$�הH��݁Pk�����`?�۲��?�m2��_�o��t����
��b���
�2 /D$����LY�S\ PH��w��:�}��w�>�՞y�ɏ�r��м~�b�Y_�ȳ7BX��d���� 6�K�PN�@%$�R�{8��]�p*�~���2K���WL�ѯ�I���9�B`�3�� X�vD�C��Z&=;�N� �����\�D��$YG�<\K��N,+)]��Y�8=Q:3^ʀB��'���C������l{&j�.�0s�vR��߉}g0Ɵ���{!k!^j8 mõ�[����C�{9�еuL�.2$~��M� ���t�f����Σ$���aM�Դ?�1��P�M����2����=����N�~��G�ٖ�n���Җe��Ҵ��e�eU�ac���W�& �a��_��vgx�WF3�W{�ȋ�^X��l��(_2��e�Og��<�"��Нt�dJh�A5�B��A��0R���z�R�Q���=?��y��5��t�'S�c�Y1yk�5��DZ��\5��G�9"�/�Hew(��m�
fn��ʙ9�[�ߒ�����s&����J�C�����Q�3L���Pv�޶~!<�M�MLR�r��4��>��	��*�u�a׽�o������X	���-8]�3�����ye�Y�\o�񆊓�I'����&\��T{��+�캊�Q����~�<�l��`?�����&������{k1�IT{�թ}Ɉh}$�<f7�*c�����ݕ@%j����Y��ݻI_� A��� W5B
��9�A�ؒd�/�>���������"�w��d�+,vW�K�C�i��D��(f§Ϋ���_zWB��} �I"��a���I�DK/����5���&~�<�Ɍ��Id4�d���*�H�I[o��A����ɨ����:�{\� �+��ڤ��5����̨�g�<+���]��H}��{雯bT�"����q��|��	�_�t�����UG��׸���m�I�*��6s�̵;)�qGi��{��+��d��p����q a����[�ǔi\��/���9�i���"9�t~{ q�pK՜;�`��{]�D)|��,�V�+0/��I��A8K���#�o�P �������_��z!?�[y4�A����zz��O��u��孟�z��$���ĸut>:�(�ߣ��߄IX�K�
��D
X=(x�J���c��r�����t����.VE7Na�p�a�Y,��[")�#P��	P����q��tU�)�\���Fi*��R���V��PV�U@ϻݳ	��qB3�U��>��rl��`e�r��ﭪ���\9���ĩ Mu%�G��x`J x�$�c��D0�S��㪪Q�=� ��:"W���w�!$��{u��~�|ϕ4��_��
�s>ԟb��u�d�eһ�b�d��7b�"AƑܿ��v���$SͰ��稆�D��������OP���z����>1�@��5>b�R�?R/�"�is�;_a�6?�w��*[���}h���۩�9�k��`4P`�
��kG疦�1j��*�n)��7����a���E�+p�"_��BK���0�(lao�)�*���9�����:D��x##��e?l��W"b�й��`��#�Z�2����,}����)�ホ7b7E)��8:�&`�bRc�=<��X�@��s�IA��Q>+$,$n�^��9�"��?�.8�*��p5��vH���ZW�Z�M�@x?����?Th~����M�^K5��t`�6%ߚ{�Hg+��b�-���P׋qk��Z�:��$u��+/�L�&��Do������E��j��,]���֌J��	y 5P��,�'�q��P7?���tϠdj�ƓM����?�z��E�Z!������	��R,��	T|JKw�wm`�d��G-a�<�j8&G����=*���[Hz�Ue��[8��sƨN���~K��%� ѥ?�*$�e�'��d9M)�=����n��!��OXn��V��è2O�F4Y7�~��^lA��]�#�����o�)�&v��>~���Gٌt�X� $O��V9.q+�0Kg�Ǯ�m*ס�I4��e�d���,�E8?M��T����vc%ya	��/uRA�����qs�d��sXK%��=��MT{	�7)���<-fp���f�?xɞ}g|>X��W9�q��u�$3W�-���A���t%|�1v�j2��+�H�\���+���ŝs��y��ԇk۬Gp�BRT�)�* ��{�U�g�[ghU�N�|�6�ݡ�e����|���g���gP�_����dt!P�9z�xЮj���E�)O�yi��S�����֦�9tF]�]�]^QP��L�����Ao M.q����;�'���.3 �)�����﹤���=AN��8��KDti�U]FK]B�ݎ�����|�ў�������L��mљ���/p����(�D��ѱ�=���Dd	�O�m�D�л�Qot����е;а �y}�a'���`_�P/>�q���4[eF�[��t@�`7���"��\�	�����A�_�`���D�����6ۻ.dc�5.-�(I����J��+�Q0H�5�l!%��-��9
I�R4<��D��zS{}���� ��I�_7����NI��OH(�@$fL�BJ1�D
�{K�����������Q-��Ĝ�ҲP���M�L��l�O��[R�)Ge*�}u�4`�@-l��e�<s>z�Ktt��J<�H�0X�*p!(x��Z���̏9_$>�����I����%}b!.�
��Q�q�9Gy���n|�+��h��G�H?�-��w�L��8ë�ʍ<ʨ %d��QȜ ���D-�vh8�g7�򓀔-;lq��1y/u�%N��g|ƭ�q�9Hc�������7������a�sW���=3�N���'����W���s�fMBZ{4.��X=�CT��Z#$!��N��d���<�l�R�+����~���ۢ�Bc�W�]LoU����&�Hի���(n�K<yv@���E�qe�j[cNB�&f_b�)h�Ԕ�����'�}�]�__d䕏u��U�B��n����+<���)�N�^ i#�Y�3�����:>c�VZ�Ԝ��}��>�@PY�1j�cf��@=�M���	�Y�Xh�c��u���ɵGF�T��di��wO�O�M,!MiD��B���~YE"U��ǥrr_p�"��&S�h$)����$b<����e�6�4�K��u��)n����Q("�	�FX=�]���gB\7&����$Ӆ@ǔ�j���<��>�`C&��%�j�x}w�vP�{D8��tM@ R1�O^��ʘS��z �=m�^�}6���Y��3�NTI&�'�K}�Ly�JN�>�Ǜ���*f��?_�Oӧc����H�
i��<XtzC6�qG�4l�ɵD�b���&tD0�7��t�]~[;�fcM'��W�V`���� 
輞#�9ʋA�n�%�ccgw9*��?�{
#d��S����Y'�e8T%��X��Q�%�9�th��A�JT9U��,��nuwXJƨ}�I1�k�Lm�v]bm��\�]xm N6�`��� J������*CT�LE'Ģ�kթ^�ug�9�ƭ��5�6�d���	�Ϧ��E�� �@}<��!���;]���t�'~�^R��cľ:7��b�f�}����S���N��í�P����C���(�_ϲ%�}qo�Y*�:%"<+!^��=Z���DΥ����J���Iy��_�1��_.�ǜ0ݺ9Ji0{����q��Ci��^�1}��oHB���*l!���(���$x1���� ���W�ut��7�
=6!�����3^zHxL+3��C��ǃ���=�.!z�S��<qzZ�|;�o$x7�W8D.ޔ�Ǧg[Q�fFD���5.�̨�w>�\��|~94!!�q-DU��/9��&���6�Ȥ�(��Ȯ�If�?��	9���ԅ̀���0�\e�l��n&�+v�;���P�*�UO�#^��bv�`O�L��yx�T��Y�b�d�eD'�`h�&[���c&W�b�S��|�ڨ�i�����4�t�w����H�i�Ѽ�1�I_n���;Bt:P>�ӊ��PYR/��X!�C�m�,�[�>E�1�o&��d�y˂|=� �=��;~:��p�S\�$Un{ui\��R*+�+�jo~�}���0���2~��B+��D,��c�,�r�2��s\�PT-»�E�EA��nbS�5����� �?Ω�'`?�K��7�/�o��/S=��a_X	X؋�~�f��������I�	���=�m��@�`Y�0�C�R�J�~)��� �Ŗ˳ <��������)���� H�8����?ƜHv�0�C�ם�k�
���>	���v��l�����(0��)�`�WZ� ��5i@l�k�Vk�_Z��i".������O<17l@��6��]حX{�M�Y_@�O�VN~0e��f6�֗n�ܰ/�6�O�����X4�f(0k�?�#.�t_�0�Ca	��NS|Jl�ӡqYЁAh�ƄH�?��I<t����/ d$��b�f��HB�?%���+)9O�r��/7�/�y�C��	�̻)�\7�<X|V�l���\��:�^�sD�� �Ꮱ�m ��6Z�Աl��y=��y����;��<P�~��q��Q8Z��;�rKi)��"Q	P�Jӹ�m)h��77�sK�������c��G�e9�t�����-�C�L�����| ��P�3U�����߲�F����h�s'Υjө��lA]E�\8���������Ƃ�����<�!8������6'�q��	V�&+�Ѯ�c|JǶK5���-®�H���e��ŏ�n,�^��:D�8�r� K�Br�fX�ʡne����(1̔(Fh��D��Z�T7'��+�$�=.�3a*� -����!��Psc�en!ۓ�����j1�,�vQ�3	M����«�������7-�2��x�����RL��<�M%���������T4�Z)����a���?,��v@���!��Fu�SI����c�eH�SvYD�1������׼�N���9Ĭ���צ��XI���DNz�I��q������� ���f9$�Կ8vΩ�"ىN�'`S-¾
Z���&'���gՂP<��C���U!�t���jyP������w�˹�J�6��?d�Q����N�55J��n��~��{y&���8Y���jih���ۉd����� �֬���-4�g�\��D�C�=O�q��9ڮ��g���C���:���_�9
_��z������m\��=��;��@���q8�����Kja^���б�"!R6՝�T%g����|�XM��a#aH���)#��p'ٲy�g��6p��b.�t�Xg����:`�V�U�M+M�AO)Rk��� ���d�E!��s�8��iР�m>����Mԏ�v+b��w��q������!��f�I�%�e�"գ�m���,�M�$}$G���4�a���oT�C�����%�w���N���P&�i �L�%'G�.��2t���^/��e�2�`Bt"6g[,�Kނ�\_�
��N�f?�� 7�{��(�UJ1D�,hJ�
 m,�4����.k
d�� z*s��/h�R+�|&B��|��5���*Q'�3�{�JNW�|�h�ډ���!�-|�I�3<�Oh��*t�q$L�fiz�ӻ����L�=N+7�ݑ�ʦ��-�֓+�O�=�Q����gy�-�j����\�����+��b��e��S��H�Y����@����4�E�^����G�(B|'�6�,9����{��4g
";a��ｎW�v�E�+�ໃOC�
��p��FLe����r`&���ʤY��#-��y�:���HML[ۄr�&f%�K��NK�%��ӣɤ� �Nj..�S�0��=;�}���[�8�!/@%����/���9zSg����[R�'"�pc�̆d��$(�+�1�n����=�����1�އ#�E�9�p�f
��z�@,LB�E�$O��ߎ-�Nk�G�Q�b>t#x����0'$S���{��`)��/��1C�OE�[�癮��Ib�X�dX�#*��J�qvI��B4P�|"���^�`��9�lL�8�v
�Wt*�Wy;4X���Bdl�"�8*��4��J��ʩ�;�&��+_5�iɂ���%�5k�"W(b��2ʶr��k�� ��xJ�[��N���5��zKF��%dj
9���N�|������>E�kְ��	��U�D�7�æ`Umٚ+�p�2;_�`P�;�,C{�m\���#!����߂�$�����Z2�쒀�oi�<85'���	���ni����{��R�f��_&�o�T'���^�n5v�5�[C��f	4|Ua<���Ď�#$W�I�wl+���{O�v{�F#�IDS&ApeM��{hz�cZ#�����"/���x*m��\͌[���mO�����1J��E�9��;��Í7�N�zy�O�øa�Lİ%�6�����X�y0}Fs�
|��i|'\1R /�Y�����h�8)p�m`��ֶw#H�h(�L_ p��}�{%^�q��Փsr�h8��^7�t�1�StLv�!+���I���ޖ6jh
�<�\|�d�S��c�q��w��sz�vK�M&�02ׯڶ*��s��g&�7
~1e����P�z����T��~b)sV>
 ���:��N������|�����2�¶�q�T������O2�ƀ����=��]�E�$�V�����Y¬+HdH�I^�K�k��(�e�+�Hx�{>�q��7�2�JXj��ŏW��%I.Y,��'��1I���@᝴�{��7K���
BI�C?�V]pҎ�a�b\����!%����s�U(�܋���򈃃�g�A.�����t&�f��9�O�{��N1!��ޣ���Y���nۜ'h�q'���lM�N>�t�	��/:��m�CIk����n��G�#?�h�O�j[)"j����^.�Vq�e��1Q��>3y��)�3baf����S{A\W�a���|&Pd�����Sh�J�b�E��;�6�=d�	���u�z�h�,�a؃�s0l�1�x�̝VEK�7�ؖ�cHe��E����u���+��/R���ѩ�׊+3j0�{�\v�5`f���r�6�����(HN&uR�����NB&Ĳ�I��1��Ġ�#C\`1�I�ݘ�NT1�H�b��1�rc�rw��M(��ܜ��2m&�3�E�2���̓�jS���S�1����7�Qw3i���C���@J$�NUXk:q6�\��jL+�(������� �W񝴳���ߐ��hQ�ay!����y7إ9�=V�H��b�`)��rG�d�Up,H��#��P��&��r��a �N6v���[g�a&�0�&��R�C�Ǎ���Kv*�f�HB��f�6W�c����m,�}ֵ�ɩdM�aP�����<���\��GB;�b]�psT =+�8�]<}���/B�i>ǎ"�X�QBA����F
~{1���l�d�cl�2p��;{Z���z������G�o4�3��@qo�mG<"B)�B��#��]�4Ը�yN�z��a�z�l�1&�f�Ǹ��F�NI�����NR�G����)y[�G��K�ةf˅��#�CJ[/"� b.!b#v�'���x6���ՙ`\q�(��|&��T-c�q�z�I%�y�8Izd���L�u�/֒B���Ż����oK���s��[-̵����������Y�4��+֚U�~�E���{c���2�g�,�/�H-�23D�.�.�6f|�J	[��%S�{�����{��Hc�Y�Ք���]8��3�$��P��!�^ꆥ|��Gn3�j��d�FYj��L������=�K�Ql�5����ߞ��\������F�<��d�94�A�OzKw���ϔT��%W؉����d��h<uӫ5պ�����(ݬn<�U X�a:y����d��J�Q�w�!��76w+ӦS�"�o��ne���M���l.ີw�p��-d˔���f��dͶ�#��9���������2p��	?��{1�7�G�|��;4���ʧL�z���V���*,���Z�E��=��:��}n�қ�	�:+�W��p���h��;n%���DJV���t�?+��2B$�{ܝ�Xԭ&��YZn��w7�iy+��ذ�#�E��#��zy���q�M��f�M��� 8GP�a��,)�%a����M�m�k��Vl%7���#�	~���
K�ߏ�*M��j"���a	��2���S~/��
^x*�%1p���k���K%�Wq�2�;�)cԣ��Hkz�y��b��tA���k��Opn�@�%Z��W+����E�����\8h)��/��G��ny}�V`j��"��7J���3*��	f:�F:�ɢ�i��{�N�%Ɣ�{8U�FԺ�G
�骥�]$�r67'7��o �"Fv'0ѿ#vE*m87��G����W�����ybV�4+����"��%��?w�ݔ�ȗ�ɧ�m���c�OiI�R_ַm����8�J��Ƭ�s�ơ�E���zw.C^�aݤ�@�-��������Z�`�̮��'���Me����(j7��J&�,��)V9�]�J����P�Rq��u_�,������5pؚc�]����e	�@%���9xh�sR b��^9�t��
�J��w9���'�k�￻Mt8��;������_۳өш�{W���c��B�|%Q�qXTC�/�4�s����R2���r>�#�����7���yM�F���p'�����@����*8ھ<��]2���io׎D^$X@S�n�aE� :ީp�0m��9�ȷ'^�:p�(�5Go啔z�����r��+{(ڕp�a�O�L8��_��r��"  pЋ�f�_V]�g�'�^��3]Љ��B��o��1��[�\f�rF�B�f刽uHMx���5G�'$H����!G��N�b�w��y�݈h���.�����Á>��+X�`���i�T�ۓ�4��CtGKn�Z�c�V�pIF/GV�W/��GӥF��Xjx�>�T����RC[^�V�C�-�F��;+�{�vs,�J��֜�^�~6��=��k4�IH�c_>��i�DM��d��%��?  �WF)>�K�����s(�1_���I/[��M3[�t��~��8���U���ߟ�5T�=�}��>MG ��}��y����Q�vP���bip�t�d�j2X	\K�1|��_��q�F� �;cT�y�m��ST��tٛ����G���r����� ŏ���E�J(�P�w*��v)�w���9cA���h	�� ���F��Ђ~Mʬ���92���橉>���s؀��;C:O�H6�D��2��`�7AT��I��u��qm f޿	\�~i/%X"�ye}��>Ѡ0������,�T�B��4���-ft��{n��f�/:&���ܘ4�Fc�z0*�Т�|G�[X>��E��,\"�*�^��jZ�h��}���\G(��R�8�Q�i+�*Ϊ�zZ�-��?�[W��*Suj��*}|�V�&K�����Yz6�-.�����׹�������v�?W^ OЎ����Ua$d]�)��Xq~.������Kob��颥���C�ܬ�����=����؛Ҫ��6���΀}��e�������"��I��S���B��Ë�	�g��ޡ���R1��k�w冝����㬡�1��ա���V�����34��6:�o`Y��{��F�vx�$��m�E@R\���q:��O���0-G�,����ld�B�?�>�T^V~r��	"���Y����.�����1�ܴ>�N��'��u�QYd@z�uڰ��be��݂e��O��q�.��1�I;��ԟ�5����#�$����"�ކ��Op��1��;�X�����Ǉ> �ʞL��w�56�d�����F{�M�H`��ԭ-Z��¡Q����9��4	���<���'���X@�BH�0��AMW�C�oq ���/��l���y���xFr7��	�r��qd�y
!���t���g��a�IBj����<�����R�MڻQ�v��\�H8�Ԋ��G��P��[B���5z�"�b��!�$�xPK��+莱r��Iɲ<�ir�޼��䲯����E
x���1d�k]�)+�j��Ҋ&[��*/bZ7�Q0���c��:�*ɉ$#E�.���#}%i��bvN�� (�-d��<Ʒ��0���Z��Ŕ=����D�;�,4�0���Tsn�j,ǞP��Ç��'�3�>\0�[��w��@�s���QI�i�$� ?U�͝��\�^�&˔���|�r>+[�py�}*�ܥ�{w �s+:��@e4����@12(�=LOz���yuF��4£�/�ӘG_V�]�E2��9��HH��� ]e���lї�ge<���5	b���6Kmc���<*2V�r�����Д��.�ж`�\���S�@%0�YQ�����T֨�1��ۈ4r>c4&S�-�nߖ8�O�����I߲Z)�Q��5F��/ W�E��/j��h�价��[6G
��9�W����m���m�G�Ƶ66?B�w�Տo�+������@c�g]20ѝB���1�)_$���S�-�Ęc�d����0iS�5Ǝ{�N�Vf�G���]��k�S|���:��/fK{ʰ/�Z��J�%3qH���l¡�zv�����Ɋ��=����J�"K���:����[�ݥ�AbyBG��:֛�X���b�v0/�� �&4�G	p%��Zk�"B�J����bB�> 2Mը�Ȥa*�zN0�[�^<�`��érR�8�WS4I�aP���"�	�7�|���6'$�uv���q������Oq�<sHj���B)�'��V8Le�Q�Q��x��RT��y'3��ډ*K�C�ƟJ�� E<�����b����x�5$ZZQ吮��h�к��(p�azb�rP끲	�JC�`��C����xZZ/�$V_���e�W�B�Jk��xV:y.H��u^hT9�����N��}:�S���6�,���1c��tr'��?J̝&38qs��<?ČZ!�o���amdq�	l����5l�V%j�S�M�X�,mK��w��2:�@�<*�Sܽk�5#^-�hV��FG��л�P
Yfs���&/�#��v�iC��T-��x�L������d�ޖ�-�U8��
 A�x�� �0�6�C �W�g�S�oQ� }���f���}S	��,�}�N!�Ց�j�L��M����BnGhs9]8n�� w��Y��P���AEa7��cT�>K~8�N�3����[RN;�����7Q̡o���|�!\�8��y9<W��*\SG3�4�� �(�j}�2�@�b�qn����F�_N۫�����T���=��t�!Z�9�:f�k7;O*�ƝZW���৫�;��g@;!�6#Q��yіp�^�Α&�R�� b;VŖҰݞ�H�M� �a�����@��C݁f��5��r��7�/V9Q���+����.���G�Ơ��wY%���LVΣ�+�oY���Q�(�.K����n�g�L�iJw�G����
�R�o��z����C w\�ve�.���Uq��)]V���*W�i��a�z��ܑp��꜎UsS����{.��NI����1�6����cI�jH��[��wAF�C��~R�.6,j{84D�X��e�x�:�QCR��� !�u���G�{�X���9QD��l������>��!z��XM[��P�FXb-#�^��z��eD��A]�����
��u�
8͵U��`�xڼMؒ@��c��C���|g�ؠ,�)ڍ:���P5؍���y+�=�a������p�_�m!ﺄ�}Z�i�<�$)t:X,su���1���VQ� <J�0�J���kс�0%ns�c�U�����0ڻ͐/z���q�S�ZM�)� �4���ԹЪ���������S1��{ۤ��$&ňQ���D�
�:����)꤮�t7}���:sU�����	�v�m�c[�Ĭp�MG��Zd�WB�T&&�����/nE����)EbJ�tp�]F�W@	G�R��/�T��������\1!7��@|O֭��Տm�t�/�Mc���c5~��0/mx�_K7��L�J��	oס�! k?�����R�:i�j4�R����t��po�JXb����U@u�JMѺ�ZWђ�da�~�3V�T��G�ᮻ�/e��zZ�0^[h�c�]3VÇ?ɜ�:�(���+����[;Ҙ�\A��n��e[�:�Cq�g�I����r����dB:�M*�s q��5Gѕw�~i�A�H���~%$�.4D�`D����;qB+15��I�ȴX������3���<�U�Qs�Iqj)P<b�*c�7��.mJ?=��k(�z�z���]'��p�ⵆ������|N���3�`Ȝ����I�P�q)8Hz0�=����(����i]`��k�y=ƶ�/�:�-0�d@H��#����Ǔ�M�E�(���@�L^Ky���3_
͜rm.���Hҧ�s��AD������2��t�x�x_�;q�C�3t�``�8

���S=�3A���ܕF�-�)�S,����PTޓ$��D9�$W�O 65�!�+}�yj��"�b��8���*�įgʩ����p@����x�\���V��*lo�L�RX��-QT��1[p��hbc�%r�un��Nz?u�O�V}:*uJ�*8d�)�~��D��{�I�����(av U�p+{?��}D�c|��,���u�w���X�ު}Y]����F1l=�+Rb�s�i]� �on��t��_9�񾋲fO�-#�����&2
�;ǎ	����Vc~���D*�:C)kJP�|���F�����ڻ?���4�Ǿʭ�ț�����/�w���u�^M�N�y{ŚU�����q����{��%S�dҞG���r[o��i��?!X���>�ԓ	��l��+=;�9�p�`�,P����?\&�u"�}�3�<�b�|? ���o��tN�{aԍB�d��<g�ѓG�|"������8>ƒ����X�,j�[�r�f�,�9��-!��I�#��������|?^lE�z
���AQ��c��c�&3��Yѩ��i0ࣴ�2J���:��Y��z˃w���t/&���9�Gh<6P�ք��W;��Չ˻�)LزfHf��d�e�W���s00��c����a��+5L�q����@�J�ځ�=���+�"0�ؼX�2��(�a���E�h:;
��2�J�Z�ͻx��G*�7�w��+��Rw�l��l�1UN2D=��*��i~�<�n��1���H��������Eb�[�3GV�EUZ��g"W̓�+d�5>)�S�F���ujW�sS�FN�N]�y0ϋ6,�k�|1�&Nj�u�����/��s6k�n�c��Gx'��=M���P����^��Lۮ�\,��c��7��]�s���4�U.��yӚ�W�vO�ޔ�^&O��
M��K��E8��y��;LD9��/�>3��x��=�:�*�K#�!HBHz�o�'a�`Gpy7T��bS��t��f��g��:��u����&��L��;��8w�y��W�^��*�{]U��a6�`�/��6��i΁,L�t
mB����_h��l�����:<[H~1�׉t�YC#�+R�H����TW�+�K~�U�o�$7�ڗ,��0��9��Oi�l�@/�ai�@V����JS�?oVl��p�\+��Ӵ1J�=�i��)fsr�2;��<�ns%1Z��ψUQ��=�����4�iF�(�QxT�+�R�G��y�׳g���0���ݸU��;e��?]��L��Lm���Ll*#
n��N�Ao��q��d�����=�	��58��/�A�j�n�M� #y���U���Я9b�2�}$.��w�b�T���Y3Euue��b�K��2Κ�P@q#��R0�
��6;8e��������}�٦�ϙG�_��`G���H>~�2R��s�U���V�w�}p�ZC�2y�P�a�RLM���J����b�i�� I[#��M΋� T�qb�%:_�rm���L�:�A['OWT�.Ǫ0Ia^<k���E���˪&���&|�6�̳�� I$��.43q��E�T��Y�A/a�;kN�"��|�+lW�8 ���*����r�>G�h����G���#n1��'j˸D�����C3��Z����0����qc7�A���Ȋ�I�Na��T��9�S�
8t"�)7�_|���ٳI���ُ�!��N�������slZ'(��C�s��y���q�x�ի;�e�XH�EiN�L���Q��?M@�	 �0��a�g`�G�q�
2����'r3��n���8�������ٺ���:=&�`=I�hɏjD�k����PQгt2�?%�M�L-1�BT��Ɠ)�No�dF��j��qh�N���r�mN��0:��,��H�Ȳ�(��M)�8\�4S\Wx��[x�OȒ�{�C�j��d�t�XD ���4���:՗�43	�����@:����p�@i׽��tU|�����&�Py��`�ޠ�5�ފ�-'�Ɉx�}��᫑��#ɦW��m)���ȩ/���b��u��9\���� �q��TQ��"ݩ�@�X:�F�2�������,��g��E���������#L:L��dAq>-_B�(��*�M텚��D����)�X�9/_pÆS��J7�߂��<��qŹ�dr���>�whB����ɜ{S��RU��"o8"�����An�Yf|�*PO5͖݋�y�?��%�N	%���G��1����+ݡW���-�y���'���� �TK
�C)Q`,"���ƣEDp��<?���noln�Xh�7��i��.Mȯ})�&w�������Q9��\�Ѷ�>}���J�єx�D7[�^�\֖�q���KҊ�АЄ�=��Xi*��Q���Y"�dW�=�ƹ-�;���]����X�g��_`�y|�A:K'?O5�aCH;p����	���C��Q=���_�b�^�ً+,p�2����瘝0�C�u���&�`F)|�HГd��N���]���7`�x
����K���c���g�����#���b�W��U^��,vp�O��%2����I��[��9r?8c��R�۫׾:V�}���	�B�Z�|$N�C.���.�\<�
��H����Ȭ���te�����<�WB<Ư�� ��I�H�k<m���9�y��M�784F�����4ȍ	Һ�{j�c|�m�L����PH��%���X7ա>�h�+�TG�ث�(٤٥�hKo?���x�6u��A]�<��!-���B`xt��l�18G��14\}r͋ᷤ
�KF���@N3�.�Q��Q�.Y��W�R�:
X�d}ݮ����@&n�v�i���P����'^U�>>��q�X)�>v���G����Buiʝ���=1H��Bω��{nu�Hw�����lk��l�PH��F�?��u`� �K����05cO��oj�`��ίa2�'���J׆�M����w��fca�
0��q�M�o.���w$�E"h~%��^���E��&K���ΐ�ºq�f���q:�Omt@�5c�v���!�1nİm�'�
����#-n�����oI���c��l�	@u8XB�OF� �:���>?��ߵn��\V�g�2�1��w"	!&�v�ł�5xt��kE���Rpx8#���`��2����0��
b'��{���ZaMM���3�[�EX=��5�K76ɬ'ۇO5Vٖv�>�LU9�+!�}t�N>�4�L�X����@e���?��ƚ���==��`;�S�L�e�-�ի��<|8e�����/���Ā�K0
��"�ɚ�ˠ�4������
�w��K��/������C �Y�w7�~����3��V��U f�WZ�kk�^~M�K�h��"˞J����&�_k������Q�4w���y����	u�c�r��p�:��?�� eC;�#�%{�\��� R�����D#l�d&u���Se�t*dᖈ�+�"����e��wUƈb
Y����2GF�*@֪އ�fM�C�HXb��r������:8�jj��n�*�V0�w�����A�a���,ur&N
����m1��W�`k��el����ƛ���Y4ȇSv�@<�v�A΢7�3��˸(�hn�Th�E�c4(��%_Fj�����m����������zK0nL�����Q;\%'_��t��y����ZGc���(�i/��E�Apk9�SFg߻Z�ӽ�JZ&/�W�V�A߭�5������e�f��_\������d�]5R���gjke��]_C��0ɀ�1G��l�b�F/���!�l*�(�*��[�F���.���1>�匣���.��ѡ{8�gn���%ɭ���i�E�]z�7���:ֱ������̞Ac��'�mw>�C�]p���sz�dŽ
�����C:�*M$
^�	�`#a�P��-��S�&UU���vkl�N��<X�
�J(w/�z��Wr�{���5n�<"�,�R��d/P�sk$��l>ӎ&PO�w�u\���(]����0�d�1��3���Jna���F�~�(f"{�֎�@�4����M���)EpG��7�a71�!������bQD��'3Ԓ��S�".L�M��+̞�1IX���b�$U�����o�mQ�[�u6����ٟ�d[��m9d���H��4z��*��}���uMIR�,q�'�
Asl�Zj��2�Ԟ+�����"&�`��t� ��0g⋁�ʃHl������wE���oA�X&�+�Td�0��5���9*5֘[�����4�f�&�%hTxɒG��K�Y�k�;p� �,tG��	�f}�6g��&/Jw��\�`���(��ݜ�f��4���¹����@�ŎC�P_1)�!
;����7��]��-�!e<�:w"�5����8:ER#��g��r�mK�"��PX�Zb#?�W@�/�����ʘwr0O��e��M�1�.D���}�*
��g<�i�e����.-�
j������� st��k\�v۸�����!|����@�S�kA�A|p�&E�&c�V�K����0)�Lx 	����t����:��oK�  ����x,;���h�7Wz��G����h�ː:�}y�n%
��x��������d	]����:�O��<jp]QҊ>$�]�6���G �xYu���TaOgĵMw~7����tzD Q��-��R`�<�.���=��/p�]�J<�7�t�����?+�Y��y��3��N�.*4z( �u1��ix.��%�r�lq�L�PB�En@����9.�p�w��}�	o��ܖ�7�fI?ݺM#�E�5O
m�v��C�Oz���R���ƅ:�����/Y��T�@�8��%���d�.���#�v�Y��`ڐ naq���"�����u5n�-��ad�;�☊}G��.�x�u���D7r����9�a��"�߱1��>��#S[�?��~xt���d���#�ȣ�?Q�&��٥h�Aɬ%$hwҼ��f���=	�;���8w��t�3Rs�W�.�E���RD�Xay&b3mW�d��� ���{I��e�;c_����DO`����Fc�6�C�|n�Q�X���	cYm�:&� � 	K@b���+p�"���_�\�}��ڵ���Sث���I �����1��<xw�t�0�t�0ֽy+�7��J�;�'��st￢-1?
����DE�wa W�`6���2oVւ��⵾��k�%�R&�S��_��w���H
 �����
7�j?��gC���&g��;��%���1S�� �<��`�5����#���I1�w�݁�Li䅗ouz� ���3�>-X�
���A�?�T!�oL��O����8'|`��{�?6�n�6\f�S�!��Zq���^ӆ�_}�l�<�A0����a�G'5sQ�KeG�S�]���A��Q����hn�x3����a��ttM��t'G|_���� �[�����ŭ������kh���y��O�Gj8þ��I�mZ| |��h�F���Na�N�h۪�"��'�u����g�	)+�
#����yj���]��b7��P@���I@p�^��d>jA���=a^!�B�����A"{ߖ�so#E�KA��&�Yz��b�F��V�+M��|�����cF{����`�\bg���[�-������J���"|�����V�\�t�vO�+�?�i�<���[�����~�[5n�u^�^&.�.�	��I��)�q��ɧ.L�{�y2%�'Uc���a�ޟ�f#��+��s�p�>����{H;a~��VQ�KK���l4�Iv��i�[�#=�b -���/��j�|f�CT+9��𸗚i&
V[ �8��b��^�a�؆!^�X[���x�6>�z�-��M���"���3{X�SH3�|����DktM�j+'��U�j�ձ��& ���
���}�s8t,���@�F
��<�@�5h'���D)^3y�+HCД m"�����z�9�~��[����|Ђ|WuDx�	 �L�����38��vQm�Un�b;��Z -�@�Xe��������Uu� 4&C
�{��o������2�>�h�Y�M�:��R`_��;2��D85�vi�v \�[www\7�9�O
of�Q�=�[��$���ĮG�!L�w�o�}ㆡ}�x���<�%�(����7�%�DD&�~F�����M
14y�?�/B�6z��t'���������:�K_Q���O~�j�b���K���Xj]��]��Әˣ(ݢv΀����$7Qxp���Ryz���gfX�)�5~��Z�� �0��̔&�ʚ���^�� P�`��4�I���G�t��I�u�z|@�[�ۯ{0;�cx ��ЭB�QD��,Џ�G�c3�׼��Db]Y�����x���}��1#��U@.Z�:�E, %����9\���hܵO����>@Z���!���C=�^'m2s��s���~�f�p.����)^iI��޻��*W��.6���Ă�h��wZ{�^�����m$���5����]΋��/�K� 0wǠ���A��W߫��3JVUgr\+Tz<��W!�?�����XKzn�Z`<�G[
��c�\��=ͩ��L�0a�>�G'X�!{��K�Qώ��۞ip�o[B~g�PK�|��1S:S������K��I���C%w6�n	`hh<A�����*BOK��P&�P������ir�5�#_!�A+�%��^g��(���I@���O�%�8z�+�6,^5�1���O�����$�����H�+B�Z� Ϸ�b��%;ߡ���\{d=f�a������oM{�L���G�U`�n-}l%�,�˧���լ@o[Qp��ܪ�}���ސʺ����Q{���8
'4a�-&���Z��y�Z�;.^$�~��K��Q��)����#�g� �@v�i#�y��i_lHdUZrNи�v]m��Bzo���"�*nw����0Ԏ4Nl�_-Vb.1������e]�PGlD���F�ey�'�N�B����틍����LA�(�{��4���LAǯ-=�
L��x~u���Ƒ�n��Bw�f%��r�e:���a2,O	��r?�`�M�i�Ecm@��Gp�:&�6q�%�ӶA#$��t b��7��/v����(y��}+�Be.�؍g@Ṹ wN]2�qo�1����� ��¹vĐ脻O8y��0�!}c�Ӡ	�X�//�,�F��XC��uX�@�R��̧߳�_P"Uƚ����AOk ʇ��y�AX4C{qI��O�S�D����7����f�xor��u�)�����.��2{�P4L��$�IJ�����A\�4`?G�(��)���8�������F�z$��"Jw�Gx��E׿��x�F�A����؂�Z�ouߔ^�'�e�F5�S����ܳ�#�� @0S˜n�H1���WA�3��j�dz�����x������&�7�G�{�mKy8ڴ����{P�-�qm�1����r�rޯR�s�=-(�q�u�Ɔ��0����0�c������ﻉ�U6��j��`O�]�ᔯ��9���' dT"��Yk2�ߣhek�w0>ZJ	�,�.�TJIX��]��>���\�b���]���5���[-���-65�ia�h�GF)��>��X</AoJ݋�a��1oK�Ǡ+a�z�$R��RB?�Z�k���2���%G�@�8�b�j�������Y"�0�?:V($?ףC���nk�w�+Q~�`;�9��_!���*�f��85��`�%k�n�/��G���TQ� PǊ���N6�z֝��BGR�gD�$�u�d:���.
T��|ʑ���F���`���@v���ǩL4!�C�2�XC��ޚ��M$z��9�|k"4:yi5\e�k�鱨�vZ��b�P�T��K}.���Qy^�$<�X�@Bߒ�B����Wh�y�>�,C(%�p�}�`��a��Z^�6�ҥ�@Y���҃_o(h�hk�o4	%	�M����w3��	�W�s����ҩ:�8^2o?�,�ԁ�ü61�xhX��Z2
�����tur���a�1�(�7�[�-u���2��ɦ�o๸�Vq���C�p_�L�[lw����Gզ��{�{�¯K��y.Vc��8!�)`X8�K�	����^�L�ϕR��ģ,K��렁k���RN��~&s޿�4i���P{b��d�O��Lِ�[7�tn?���˻WW��<�C"��`���c�V(!���e���Of`[\�*��o��j"k]�#�j)ͱ��5ȊO���vp�Q1j�)m�J71Rh�W�~���2U
�b���(V��%�r���ՙC��[@K�S���>�p����Xt���߹\H Ͼ@���w�����Py��H �mmw!����r�Uye�h�3qT2�~��8�9m�n���^8AfzႷ��C�\�GL/(i��H�
�wA��3�cW9ß���L��o�[n%ΰ�?����OjU�t9/�IA0%���0�i�]��h�gZ:����[����ٵ<ܼ2=j7�AyL-��ҳ�y���M�
fA��h�!�H%<��U2w_=�bD2D^��f_Z�IM(���,�V��[$�%��<�o�cQ)\��c�)%��mȡ�
�Ҥ��a
!&9��L}�n��*���Q��qR�vЯ�L�˷x���x���|�O�986M>����#�f:���D�	+�-�x�z�qE��pZ��hW�i����ح���pO��xq-G(��5e�bz�I! ]\�΍_{oJ'XT��4}�F�2���<�ahG�!��h��<6U��
����:nv�[ed�_��ۺ�?����XN���;�'#��t��bf[>: ��c�shM㷗�4yB��g������6>aU���`������>R�9}B�P�@��{��.�q�8RԂ����>���	�\ ��ϳ��c���uj����C:'�2Y��`{�)�������J>0_��N�E*Q��Vp��ҹ��*�ɺ:� d?uQ-(��(ix�6��̜��d���׶�H�Cv���I�Վ�K+Ԇ�p���{�	/�{��9��U�ѐ�T�Lv���6�]Y��f=�D��F�H4兑"�%؂Ĺ!���+�.��Z�q���釋��X��]byb���s�n�i  ����"��@ͤ8�	���0�|S���bt��.?✁�%����d�"Hr2^�0�h�Sx\��#N0 UN���ͥ����5P�Ѥ	��(�zԧ����a0��H���,���}D�
`�q��wQ�ް<��[�����pE�UGmT/
�����|��ԝ"�Z!��;K ^��S�)�0�-�iz��Dw�zM�����l��	�B���"�!��н��Dk�x�
�80��~K��ҿ��8�)%vv-$�
�^隙1�Ԋ�\��k�,ٍ����d�݅?��gM�ɖG��qh�V�L��20�`-r�j�i�;�����ަ�R�Ԉ�3�
��7����O�5=\�T\}NQ�z��\���/ϯ�U�&�D�"�Ñ�e*w%O��&�7%�m_��� �ʊ�Ż�L�+��V"�.� �UJ���?@����@ݡ�{/2'@�
O��T��i(I�BA�5��u]P�u')�����p��{d"�^��aI���(t��l�4aك�"���T�����֭��s�~9�t{�"\t��Su�����J@�|#�7���]��CagĪғ���4�nk�f	����ͻO>�㘙=�6�a�bx�Uo��PUiፀ!�E�����Gs$f@x��2���x=@OЇ��j��9E����8-	x(d�j��j;���cqd�����2�=���"Fu$/��j5�o����B5�_r4�/@2�`Ͻ�q�*RPT �$�