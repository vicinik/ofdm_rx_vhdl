��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P���1j"#X[ˎ���~�H����^c�x�����v�/E���_pþ��bɺ���8НRos�4�8ڂVW9#)��7�͔���t��r	�%�y�!��f��\c�鉚��P�p�����&Y^��Ǒ15���=�1�^}Vz0�����P)�i`��y:���O�A@Co���/�ڵ�?n ��77���������5��]q��8r�7�5���| =����tx�9�Պ`r����ʿ�>�wyM.h;��C@ N����Ɇyh:x@��?��l�[Ϸ��ݗ��sj�>cǨ
F���o�k\3;W?���܍��$���E5��}yh�:/g��6��EYّ�*���u��xd����R��2�&�ѯ�{�@�rȃò�k����qr�wh�ߊ�L:�F�j[���?|`��s�؟RjH���75\�KR@A _��<����w'(M�X�����J�ק���fŸ���s�g4`BT��d�	�Ad�tyCg����$:h��+GRU[<,qg�� ��L�,!Z,�?'����G AXQΉ�fN���FO���?�p��<��Bjr�'�}�� U5,�1�:�Wo"�nВO	z�����Q!�/�-�Cz�:U%�*Z��=bX�H�I�K��B"�U�@�:p�(g��s� �)����ьV�������DM�$�n���+S�R#3����	V{~A�}@����J�P|����~=A��1��������x�[G�)MX�w�Qc�%jۍq�`?�I�j�%c�aؙ��H��W'4~�01����֍�����L�rJqa�hF�uA813�S��KN�Z�tD�#����m��<xg<U���>���^V�É�.Fƅ`>8��SQ�O�����J5H*r �����LkwS2���m���폶<�ӒV$U��w*+�F�MS��ȫ>�bB�{d���.9c�z�.�wq_�̯i7�b-	Ԅq�|)��Ý���KP�g�����PɪN��"#T�W�� ��YH/����P𹻧�?l�� Ӂ��K
3��q3�!����;o��7��y���	@���� 8xL6��v0�1����:����ǈ������E�wb��������k�����<%m�c��+m�:�x�]
L!U��Z�*k�yc��	�\@�P��aq�������I��|��q�S���΂�Y|�'��@5Ӥ�h��#���\�t[��~"���*�P�+�k �D1���f�l5�Ӏ�I��#�lC"x�,Ÿ-���Ce���P�7[+3�H%7ӏ�>��B�F�Ez�pY�d^�g�4���pԮZ��T��š�)��!p�v��q� ��d��l:���Y!�<|��s�v<��ă���+[gn�L�����Ɲ0a�E�L���2�~ �C5ŗ�v�8�>R����闭B��-�U��1Z'[����F�� b"Oc�/����n�z`�bF�����ʷ�������=/�I.���\���O�� g�)3�Uh�c����I��U�饤䳈ՒG��d�����2��-�5#bSeGR����f��ok߇N~��{���4����r��A��=)�՝��O�S���R��)�um�'��T$�B����3�1.��^g'͚��s�������s��p���,/[�}��s������7�
-�:-^�k��Y�ސ��-=!������E�T���`��ݣxg��&�*/���>�_3�;�a���s�~�7�wj�� ��l�:��+ŕxl�.�l����1&���U�4��[�����!��V8ʝnD5��tb<�D�3�p�'�3{8"�/p(uς�d��!���s�kk�s����nf7�������W�8�I�G�p�R>z[��7KK~�YW+���N�D\��N�o��E79ԭ����`~	��U0�o�����ڧ3�|X'k٘S6Y��K���xv�l}I�&[!�úIB�k��`�G��fX�f�z瘦Ź`�?���k���GYq��	�a�lr�gc�����:�S{z�8g��-	�D����,�W'̒���mc�_O�:�~������@ML�zb��Ǽ���EP�!5��ս�>=���ᪿ'����ab�q�%2��f��:���&;Ԩ,�����7+Q�O�`7��v�]{��\CJ�.������yNay(m������@O���c�ܵv��	�p��e��ɴ�C�ʽBl�[�*��Sa����$ۄ�y�����8Э"g��A��'�\x4�	g5���l)�X���>����:�>�PaY�)H���4��?lV�G����Z-;���$�N!�_����SL���+�5�z�b��#/$?�t�n-����=�bX��$�����ԏr<�	�>e��'qb�'�~��Jx����Ώ���D�6!����H̜H�R;�@�u���M��a� X� j[��Q��n4�s��c��(*z���DB�|��S���TL�2�8�R��������7���i�z��X^��£*
5ن��.n�w�=��X��x�Dc�g�e� =q��x��s��x�B\\�*u���oz��F�Y�
Ut^f�1i�3���g!p�Y��m|rDAf���i|Z�wq�i�9&��DCL9�1M���m,b+���:ύ?�s>��)�?hNl���%uaI!�f"w4Y�.��B��8]��V|��
HQ?�����0�<h^L�ɠ׬v�V��?A�X��W�ܑf�s���İ��Œ$.4�NFs�����e���,��dc�N�Ѹ�H&n�3�/bA�������`.����~-pd �d
sT	F
kF�n��6�tj
��E1��&�$�J�G�LX�%=���j�D��yP�Z�cH�(z��8G9bDC�0ãDf�*5�6��d`�w$[��E"��W�޸k{��6���N�2
���Zl��`K[On]ĤNL���u����Q�w���S��i`Y&���o��mn���鲊�T]<��9�.44�i񆱠��������)E�.6ħ�q��&���V#�wd
F��(��������-C�=�"�Q��
W�dvy�.��3ɼf�����Y���&י���._�|�J;�<SP����V^�s�u�r������}*�2�rk�s�ғ^��~�	�yE` ������@d\��:�7!�ls�@�>��묂��q^ �����B�t}8I��slw��hU�@L�Ί��+�z��_yK,�p�!�B��;4�	� @*��t�� W���B��1�( ����&����N!"z�G������s;߻�m��o8V�ʰ��UE2��Cr#Nr�vB�1q�*5ǿ����+!�d�Q�{?���vߌ�@g�&OV���	� 䚟��R�=L_=pU.3�C�n6l���\貣i'�L�8͟��Q�>��"��[�z�j��	fI0kf�M��z⼡«�^�2,�r��3L�J��0�Uf�>������ygE;.�>�p��KJ�a�AǏƖ�"s7�=W���,����nf��g$��7)3>d���p�,y�6q��P�q�1i��k:>��p��eg�k^������hAÃR����	��T�O#Mr�頾��Y���l��Z��
f�����Z1%�*t|%vC�%���G{j��|x
�s�)�`:���z�G/�Qr�U?{9�q#��="@вa�����G!H�ٴ;c�B���iR��Eʧ��<8��N� ��c ���ZN���M?��y�b��pP��Wu�9��$�j�-��T}�-v.�]��l'�k*$g��`������3Gw@69P�p�GJ��.��4��˲C�� Ct��&�S0�2ݡ0��
ծ�j��>D����J��y$F@`�+U�}��z'mF���Ry/��@WZ�Qv�o�H�B��5l�O�w�32�k��� ͯ���*])d�Ł'J�u��Q.`C-J���"��4���%J�v�EX�5�l���܎�ϟ,�֛�s �M����P�e��M��ax}.�TW<W�~�@�sfݛ����p��#V�,��\X�٣�OKچ8���v�c�&�1��?�t�G�1.�#`�5�\�(�fu����`�Þ�I�5-�d����(BN Bj�jP�^K�����X�j��
�&fY� �m�BÍ,�=Z�刽0P��f�-w����FRD+�a��j�x��&�x�����{)+J����h��2�alS��w��tp�H�ӻ��`iv�=k��Z�ft�>��Pa�Z>^�gH�n�c���/�[x$�����U�	�r$J�'�>����si�0�v8�9q�on����!,k��A#W�=��p5��=��H���GD �Pr�7]�_#�aI�RX_]}Z�#P�O�>6A�w���-���S���c��4VΟ�㖎��אw�3���S�}��yXA�䤴>�<�$(�g�s�s3���|��OU<@)h��;���]�Klj�?+�=�T(cV�����jv�ݡ�wǘ����Һ��ק�"c�����2]I�,kѕ���f�u���v&i� ���]U�<�Z�݂�q�'�+dkSc�����=� ŵ�O��S��S0���{��f:_GKV@�<���P6-{�f���d���}R����c�cz�\h!���Gߒ���&F�A�Q=OC��gC?u��-܊mxRm������D���7��hD�f���ȇ�4C	�kn
Z��ʠ��Ⱥ����4��5���٥ �5�͟�m��f�ըL���3D�s�j]9j��mt�i��ۿ���9�v��z�y��?��Z'J"��B�@�^go�iR0#�r��,��3�,7t,`�GfB|9~b���҆�а�_#e�e�􆥕l.@�<<�'��|����0�[�3�Eң�n۹ {O>ky ^^?�hw� q3��g�&��ʦ�"�����~.S�r�b+�G�AYv�(,�����2%��yhwF(mˉL3� W�#�ae^"櫬��9y�DU�k�<�A�\Z~��?��A�z$e�(�K��<
�D=��Ebv�U��9W��P���U�q��o�%O<(�b��3_;||T_���e��YG`�$�͡�8.mH�Z��.����Hȷo�0��	�mw���1���Ȣ�=��/yl��������.�U���6�u��#��Џb�� �%~������F1��(0`
"��_O���b����)$I���?�Ife�i"w�FS�!�aQ_5�w�:�d�K�0x���%���Y��NH˜`
����S�-~�+q'ʳhRd@�V#�Vl�8�d.RH��
fwwAȁ��i��:7�����4 �D��Z������X��0�=z̑J
Z�:�I�8��cUq�����$�}��Ⱦsڶ�W��2��E�oT����+�0��b��[���������[���oJXs�rK��{���ւ�.n��6��;���n`:#f?6$�3�#v爆OLd�1���)ci��I��1k��t(�hB�Q7�C�]XM`��9�!��W�3j0&�:=Y�'*� ���:��&�<Ge��na9be�M/���1٣�� _W/�+G#o�q^��[�n��(D��m��1W�#s��}�x��Y�1Z�nG�2�?+�v�B)�7�P Xy���WI/�D�.�n]����~أ:��W��7�4������ܣۗo> ��9����{�4�v-�iw�9��(��/ô��GE���I�r��&�
>.S�ܸ%�7W��Q��D+���}�T�W�PT.Z���%dR.$:c�}J�W��n���˔��s�ʂ2��1���Zl/��'`���>|Lo4�;��<W�g4�MBI�2��s� a����g�y+�I�"�I�w2iD�(��Ua���i��������N{3k/?�־�Η�l+�0�ܪ��������%"!��w6�Em��5@�n�"����8�JB���ih�St&�&�*%��H�h�'��Dtr���L4�Ja�^C�*t� ;�I��r�M���q�K�<\!�>xX�Tv*?KAJpo8s�� X_��iב�R�Eyҵi�g*��p&�<5��f�g��䁴%=�8�$���_�.N; zz��D�N9�M8��e���!9u*�$�1�m�G3�a��J�`@;�4�7���M��F���'�5���f��]��$�>��S���+���S�U�k�DhִD��u�a��z�@��!�E�G�k�	e�Q����LSeϑ���3B�p���-å��	�a���X�܎��Т�T&���[fiX5C��eck1�IOHe�&a#8{�ڽ�>���:��8� �[�kh�w�u��{+<�(��C�ڴՑ�b���r���q��1""��`m��p܎����Tڌ�PV��(�[}PY�wJ�7�������yg��S[w��R������%b�#�}Z��,���c1w�'�N�=�h�B�65���83+Ru����;Ј�� �g��� 9Ș��|����`��:!5wP��)�h�/��Y�/N_��+���@�@R�>����e�⡢� 
����=��~(��c���;���05�<�V�����U�)�ʂ��TV4І�+��]��,�9.|�����2�J�ؠ�+�ܼ����J��%S��F^W>C�2�� �@�`z`eW�Y�������d����b��l���ڪSxG䳻�eFrUM e�t��_�,�`c�u��ѽJ{�/A�.dz�5�+B��������j����/�+&��)�B�z����06�[*mN�%A%'�;�$��P�W�M�F\Eq�,1�F�5�D�>>�V�#g"���<�Qx�<OM�7��%觼������8�.y"�s`6fx<3��A��N�n�+J�h��_�5ѝ���쮲޶E�l����,;�O{6[Z�*��v��-�c��?jL�2�]�'�׈2��f�t,�A���p�268bbetUi(nQ!>�Ȱ��3�ʋ�$[�&b��e���Y`{��b���+����IZ����Ӫz��7�!�j\�;��:�����a^}aws���t��\g�C��:c?�ָ|)���/=Ȱ}a�	�Z��ܝۂ��X��sz��cTInB�C ���*�x�M�c@q,��bz�o�ȥ.#L�����Z�>;���c�3i
i��W���p��)tN���u��Q�^6�6�(����a�ѣq#4� E�Y��r �%�`�D0!�ƛ>%h�
�з��!�ͩj���܅�d����	!]�\a�9ن+	�f`x�t�����'�"�ѓR�� ��@��ݸ���c��;}�
�qU���Д�f6�U�n���;�㉠�䴙�����~(� u��^�/�i�AS���](�԰�13d�w7�=�W��nZW�o+31�Z�s:P�dHfȋ
�!"v��H�GO�&�-nP�I�w�O�u;��_��4��d����1����;��E����Vw�/\���{���v%$m<���#f�_��.c��sj�K�Y� �2�a9VeSD;�������_�ߜ��&9��Bݭc���������כ���>@ſ�ep� �B�#*u�:����G�VM�/����\���-�1�V�X�9l�Z�Q!OAW��fÓS�������q�����=��� ��,�M�)��}̑^�=�]���K��p0cX�TFF^�O�V8�y��dy\���LI�}P��QB�ֵ� GBԺJ��O���訾#ȣ�-�dː����L8�7#��X��;�����4t�[1��*���z�M�(!+��a$���,�F*�`5�n9�k�v�$��v�z��*V>u��1�:�����.*!an�n�6VRoס�����B*�m�d=��%�ʦաy�2�` k�JHI�=�,�Ɔ����k�4��f7"�
1�1�'�eug\c
�2O"T�cSw�
	��Ԓm ~��p��N;�S�;