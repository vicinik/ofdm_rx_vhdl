��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��Pޕi�sݟbC��i3|T�8{S���TzG���j=�m
	Iy5�ShV�Q� �������c���g�nzn�h�?�N.l&�����
1G�p��s�E۔�](����Ǹ�1���0��K������b);l+�iH� �I���jR���V��k�alT�t� �����X3��K�!��D�蔠��P4�4a�,9�T��v�|�_A�v�:��j���A�o.�X�{7�*,,�R���aՑ8R�&laK9����jr$mO�F"����kc[�����9�t6iy���vb)�NzEl�VC�2{��Cłs�s�,�ܮɌ�-_�$��-= L�
�A��������T�)��˧�;�в�kF�i/�)t �QV�ATt�e
�2�S��pv��<eT�G�F����ɚj���p�_��:~j���R��fy(�D��W����l>,Tiw�j��ٞ'*�����>h��ܱƉ0u��Ly3T���\�'WT�
)kbˏ��Oe��N� '�ԍ.[o��`	y9�W�z�%kG׹+�t����Q�b=IJ���td�#��$��Xt��bّבCR�_j��G�4'�iH/*��1�7����Q!,��B�K�����G�����MD�3�]Zx������VbF�����(�F���̀
�t�����D����U�䬣�Z`k ���=����	�:�6�G�#Z�m]���R:�X��ra0��m�����U���\��K���%�EΨ��_�\��O��Ƥ����3����_B-���=rx��Y�n���E.��L��'8QEK��IϹ��RX��rbr;���&�
*��F7��0
�����"�V���X��������˘Zihb�?��I�^7�س:��n`7����6�:X3C3Kb!q`���4��Z�Đ�< ]�
�՞��Р)�	^h
��"
���-Qz�D���{G�喙_.b��I�z�"ȑZ�%��u " ���M������\-ӎT�'�,b����5HuQ�7P�V���Ns�R="�Y���Ý�'a�<f�3���k��4�K�X���uZ��-l4$r��v�S	����ҽ��C}U'�V)P�\M�h��6Eo��2,6��qz�^��S�` ؈N-�l��د�1h�\�uC*�V�R}@�˟�c?�N���J���nE�j6Uަs[lm=J?����z��V��,~�1�����(ۚr��1�ܕC'�;b������\��3 VW�����3Jz4���+AY����e�W��k7���Eϻ���Ԣ5՜�_,e�/��i> L����,����8ԑ����|)�z�q�c����٢����Sc�Gf>��ɚ��H8���ɋ����o��6�������.�1j&��A�D�H!���ҝ/��!15j�<�:[����СwW�X� �� �c����gL�i�woy'�.�$��G ���; Q��.��"[)-D��MV�*�swX�0)����� �=&��x�����6N�3_T{Eh�+^��Z[`���hsa�v^����oy;����7�|���e��C��C��6I:���1��=�Y�(>�PFd�����%�����{Ӗg\�9?q����s�x[��$T!�A�����=N�-�r�|�J��P�SO�(
)��4�^@7a�������c�ؓ%򄳟�O�&�@%euJ�aĕN�/'���`/X����b�vZp���{[K��^_��"1,�åYn�ғ�D����1�JLY�W8�V�:�pn�'5��˪���Mi��e]a$S�A`��Z�|�X�U��O�C�����D�������c��\��?�v!�,�Ґ�����iH>U���]5��Y��F��1O���<ʗ�H)�5��P�I�D��Cv��37�U:�����I��HB|�`��g�k-���k�d��$<���%��*���o}��&�DO��&E��X2X����N�L<��D��aH<�WLB}6rVD���'j匇wJe���T��ԧ7��wl�/��N{Wm?�����>��ծ{��(�Md�����P��n�[:�n53w����9۫���L���
I�Μ��+N���v�.r�+�k\�x5:�q�Q���}�+�0TT5���HЌ��\0���'`�CeQ���t�ٓ��^+/W������q�ﱤ+\��g�5U!*7�v���&{����X��>��%�͚�ܗڠ:�͑�X���ה��4_��P���E���Hu�CC��+�m^g!�r鶐��0p�C�)x�>)�)Em2
�jLb:�5�i�.��879!߯��m�l���2ϖsN�<]Q���d2����Q���KV3�=�.�o�^�&�}�b՛-^}�p���(t;�q'�%Ƀ�����%��"V���⛲Eۈ^:ܖ�y�(�u�M1����'�/�X5�ڒ!�2D�,U��6v��).p�"_��:bl��핖H���~<F��璆��Ͽ�m�]ɜ8��|�Ņ����$�m���{_o�����?��|sV�Ti��5��Q������28� ������q�r�2���`���_�o��������Hs�\B5x@�Y-����\�)�1�f���M�$0��?*򺛁�����v6E��������[P���h��Ĩ��]�"�ܷb߂�'�O����O�Z"��x�<��$� ��8<�b�'�Pۉ0XS��DoO��$r�g&�V�x&��B�y��!Oc%Ԩ�u[j�͕�c~T�a8 ���qT�c�{?r8����az�Uen��mN��mC�=iJz��K��1>��,8(���%�ù�p�#tOIO*�k.k��K%��t%���Iw�r�����@Y�T?{�"\��{X8C�Z�]}��lh�'���K�JD��)�*��y��S3��8��MG��Ӊ����=�a����h��X��0Cn0�f����� D������^���YO~o��S�L�l:��gu�_┼�r��)�a��o�,8�L�%&�D&5��;���[��	�������IS]�^.#]N>T^�;͉�s�y��}�Ѽ�4��b�0 7w5�$�뿤xRď}r�S��u����2Ѿr̽T1�x�� ��E*�U]aw���R2:	ƙ����� ���I��
:O�t]0V픋�?~~
�{���\�ȵX���G�+!+Z�Q#��	3.���Ω**]�}2�Y\$�K�R����s
:á�ey�p�Z�&R�x�9
U�~0�2#� �Kkԅ�g���Ȝc�`������C��Z*_<���,���S!���^Q�c<8�kzqp\�c�n�?:��{��ΟI:v�W�t9�����9M�T.�1
���L�4�&?�A�',�Y-�Jv��E@M��;���d4��ن�i�Ɏ������\\!f� �{���HJf���n�EAq?��S�����|�&��EN�0֒3Go����'���=\�$ͮ�j �8�x՜�y��͛nV�2�&��۟��.�1IC{�6��Bic_�eu�lyV��� �,�����^�rr9�E;؋��y��kDŢ*��"�q��rZ���▔HY���]*��k�?����_С����+�1u2"�/&!V}"����Q�[z�%�jR���@7n^3��t�X@��܁$���{׏����r�)H�(=���C���f/��n����BM��� ����.���m�.��]V�7~2����|��<SCj*�vt�E���G���F���(-f��Xjw"�%M�Ex4�z{O�1
E2�6�s� �P*%�i�	�&P�=�C�گ��#r�<�}��Mt�k\N;]bv�A{\��$_��.��`��x��ݱO����2���V����m�S��o�}��	&�M7-���Ho���>,M6ev>����r�[Gfm��X�{�ѩ�آHOS㰁;�nx��ՖY���K���뜩�~~�m��H���'	�i��E8EA_?s�m;�]R�lW���/t�7B)�n�bAO�Ȟ������+B�2C��9Rp���7����gʖ���"-�Uᦼ\����r3KB1~Hd^���}V���"��>�	��pע���8�.��������\�U4�=��S�0G\	f]Gt2�+)�������1��Dp����B=5�q6�/�a}F}f���LpC�v苢*G&��һK���&��
��[���(Rc����p�BL��
n%�n�����ȣu�;��P�]1���Y��c��'K���Y�E��kP)��;�J�ɼ����:��nQ�rZ�*�qFJ�
�N� �}W�l���y>�T]��"@6Պ7�)q�}�;4g�D���۩�|�<�xZ�d��;�Mu?�ӄ?|��:<~��4w�6��	�dI؍3O/p ^$d�q�2�O�"	�����V���P#e3���%�K�Hڤ���hfx�"-��Q<������ů�>^��Rᶡ9�8�_D�p���9�V9ַVS��p��.�?�Sޣ|G�7/U��F#-=L|7��"�,�ik��H�&�YW���@�5B��h�h�Ɉk���t���G�T���*u	
a���oɎ+n�j��[_x�b�|�TЂHrje�U�p0=%I����_�Gã�µ	byA?��U�G���R�f�E��#����=������+��ْ&]����V2�,Bd�f%n]3m�60pPy��$��(�9�;�_�?tsn0�ʶYT�[�b����Hg�9^��^���!\���G�6'˷�~�D����y���1`L�[�w��6"U~��۷��>�b��nR�<�8�u]��1���z'�A��]�Z;9e�8�<� �����nD1:kɽ-�;&>bڛg�Q�Muo�tBC��~�m���F�B8��qI���02FYI�IL���4�����s-*�Fx���Y�kJ?�x;R���U��)*���K�f���3,��$ (�/�[�Ac,�.�2�=�����@t���O-�����6 ��#��*���^��o��Mkl�"���6خ�w��i�_��*�/ �ʖF�հ.O4,����Ͳ�ƍr�Q�ݕG�����LW�dt)��)��������-��#��s�������H����b�͕�B���N�fsNҜ�@��kG���;�%\��%���Gy�B��؀ZzV�d�@�3˪ˤ��/����D�&ٔ�[v�_培��,Y�����a����?�̾��h�D( "[1����]D��$�̷�q��7������*���R��l�+U�j�?cfI'��3���2�c��o��6�If�W(}®���4���9'���D�� U/(�)����?-�3�^�F�{IŸ:H ��f�ʇM��l��eD�����V��2�U�����s���:l�#G�]y`��کs��O	+��[+�7�����#�F�y����=�P|ڝ61������?�n��%sM�t�g�T���8(�U�~����5�>U�U���	���fD_!���z�?�͜�d|�Z:q15�q��j5J>y��i��$�$�*?��D�ڜ�1@�E�*~�b��Zޚ�h(z���ʍ�X)�>�u���k*3��Zs{�g?�cs����V�@NhE��5�Uhሎn��*��e>Z'���U'�͔���L�����@��>�>���]Ņ�77�*�e�|s�M�	t2)�)U;���ptQ":l��9b )�����(q�=V���ܙ�[S���j`�#�HB���Դ����*`���{��?�3�Մ��m%�ì�&<r_6���gb�x���Sb�NZڕ�f`ùx�r�������^>�\XT� pC&�H��J@�+��rD$>��3����YĒ�92P
���8y�Ή���$�z��h�g�{�f���J!I;ے�I�
y���x�ڑ��`K�7vA�u��NO*�zQ��i�ٗ�>F4�,�#�ǧ2�ʄ��S�V(����.��p�?�/dLt%�$�.'�ɟl�W�?أ]Q�_UYD<���G����o��h*I
8�<=���(��яT��&���n��7���K#3Ό"c��yj����J���0��v��+|��A�Y�ڪ�J��_� 51�V�u�J�K�ݙ�nh)�&���E!S-���;�J�y6 �s�uJ?#}��7���{���tf
� S�h�K�f��XO�r/j�ؚn���f�-+��a�[�l�Hy0���2�`�ן�AO����#�6QR�I��Ǚ�Wo+S�v
	=�ۯ��/�sFw���c�xHW�����>+%�v��A����m��tB��)Ops��gJ���n&�\
i�qI�����>A�M���d�m��o��C�؇p.��7��vE�g3�>�q���c#�������ʘnb�S�|�= �{���F�竪x7ၠ��G[��C�$���2�0����,˓1��M�O�,8��������3A�i~�̙�^J�9*1�\ �4i�v��}0$��y�R<]Ď����o����6uh%B �J� ����s�����a���T��tt�Dc�`PzGܕ9��T�D��Wɫ�Ė�`�,����t�d��Y�����n8�PnV;����Jc���~U8\�A�uk���)�;��=�	�9�o�'S;ԫ�0��.)��Zl�u�+O\B��!n+sq??$S'�]`�o�4����thǪ�h��'u���N���He��M��LR�2��'��}���6%S�W����Pv&0X¯@�a�ˇi/�_+���$�(
�L�FE���5�����C8&��|�!��������)_�͆�5���M���(���i2�3̟
�J��@%�ិƷ=��x�c*i�	��r�A塢9]"\
���n�P/\F�i�I64�g��q���]�7�[�m�~�v��(�M٥��>g��i���^J
) ř�9e��D���i]P	+B-5Cd�����l4�fB�|��k����"���NQ�PF��pk!�(h�>�<p$�a�I#�OR(�	��][<����[k� ��5�(d$��2�16�떙���{���&�C�S\��`-��Gڠ<�U����~}�kiäD�7;AonF,I�1Ϡ�~ `
�����nnqZH%ٽh~Ƨp�nz������4�#s��{I����2Vq3��bHPث��0Xk��U���[��Η�VD�v����f
b$��W'j��K��rq?h��g�������F#�����Bǃw�� 	`S��	31^8-�{?�3�+h��5-r����DO�.��L��z��>v��m3�_�^P�0��R���E���uq��zjjXѕ��-	bљ:M�4*�d�{����'�v.2˷�+,Ǯ��!��%r����r� Y��m{N1����FЗĉZ��G�n��.�t@P����8J.���h(b��_��+���x���R��9x$�k��U��Tv��U :j4˵���0���c����*��i,�=���/�A �S��}*(.I���T����	��l��eMm�.C
V�- �!-M��ö���تm!w�PkL�F�û)���MA�я���ݠ/h���aH	�g>/@G��������Y(R�5�y� ���7�zy� �eu۸Q|M��r��2ɖ󥆘�
����˧�����  =��Hrf��\5�1/a���&q�}F���"���	.���"��
�?�=��uN�p���ꉀO�͞.�Y�׺��Y�j0�I[�r|�Г��֭o�^��%��f�FGX��F��1.��)�2b�;@n/(����#��Ʋ$�����v��U���C���~�����o����2��k�|U$#�w��@����56�����q��qӳ�qꐮ�p����{|�~0�5����Y�ݙ�^�s`3��� �n^m��d6�B��y_��7bR�M	�7b�w��G,#8x��%C�4�]�f�%S�����t3q�I��AX�Bt�Hҋ�Z��h%?�U($�ԒI��˗|��i�a�F��"���׾�ܷ��`��Ri6դK����i�:W��W81�!�_KBc����^v��)�C��P�i�� �f>�$�3��]�hȜ�P�+��[?B^.x���9P:�N=�Mns���?�G�s���=�}e��\�	�VQ;�*���.gu��g7[8��ӂOO\2}��o�:qćx�YX���t0��'��VՔ[N9V}H6���� P��	ڐ�9Y9��4�TG ��UG`[4ߩ�Q������v���Ef񫶦�������.����8WO^�����C��l���8��RҘR�Sre�ٔA�x-�a�<g���;���4l)���=������2��C�ӷ�~D)��7r�Z���D~�_���ပ:���yb��H"��� �X�A��㷡�v�+43�3�LM��A`���ρ-w]s3h�����M�(�j�|���h�W�ގ8��G<����%h��'�Z.��l������g�E��v�|&E��J<E��&�}��R=׳��K[g]o
^�r��c�P	���6���]s���>�VZ��\��S�t�$b��!2)��=��01��޻>���Ο�m�BA�o8t�0q+��=	U��*}b8��$�0�N*���'�3%�k��F������@��H��R�m�l�k�)�%౅��t�MLy
�