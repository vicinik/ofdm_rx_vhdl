��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7�����������	$��BR/�`�f����=|o�hN�<Q��^0Fx{!o �<v��	 �[���y1�E�Tڅ7I'��7�'^#��́��y�'�a�� O�KEʇ�m����@��=P%#3��(M8���p'����U*9�����J��Zm�;�}j8X)��Ӗ]?yMm����mN.������j��p�]�H��%Xg5Ԥ*�X���9y�J���\���7{�f���]V���^+�F��6��?k	5�H��9�<���w�at��a�oA[3�r�QA���R'�`R�^�鷃07���)ص2����d�\�跮�:�˄�	
�bqMBܭ D�"V}5y5�"9�|,�K�T�҇�'�.# O�&N`�]�סO"�xN%���u�Fcj���{}��$1b�ƚvy䏏m��D]E��"�}�\���A���n!J�}��	�_7�_���Fwo�v	N��9��C��*� �������ZhH�FIZ��L\���U"�����VL�Ȭ�)�C ��Ā���+��1���D�R ��MU��j��IU���N؉>EBɫ$ޮz�Di�!#������{���Q��ol��!���|?�b�.��_m��9��_1�<ϼz)�I9���O̪3dP_WkC��if�Lo�F�E�sjh����օ�����n}���]Er^���'\�����f��uӁ)�-��d��u��s:u����\M�psD������T�6 ��@�wq�5� @�O���M�IpF��F�����T��Ce$z���	,(>�/��ȋ0J.A�����Yv~Y�%�;�Ҡ�b5P�-��_��<�}�f_-����Nf�'�~�?_op�ȊŀP:+�ѐ��>�ep��Ď�s*�˫������VՋ�C�;A�g�F=W�/;��(6Pl�m�y�{c���6I{���^:pt�jE��9.�H�M�,#�RJJe%�=�c�3�H"�����%tcǒ�зTقA{��:��̥S��Q�;���02���>�s�̲�,�O��b��~�'�9����<��]���x���^y�IeFY�-��4�M�i�Tk���8[.{Ј�a�vL
(n���^=`���5C�b�1I�B���L�gI �:b�kyqXV�
[��4.+�����hM~azA�DV�����Z��5Q�ub{ދ6{���%���a��FY��OyP'�A��x�Vzk�ͤ}�$��t�ϊ�#�GԒ���)�#�e��粉�����7������`�W$�*�<�8k}�B̋��A��A��`.�I�6���ê�H_�IP]x��^GӶXLHr1z}$�<�B̤�v��
����~�5q{�S������r�U������*V�~�W�;R������~]4X�{8���}S�4vT>�F�C�X^����%m�����6C�d�Yx�(!c6!@Qr�k�뮀�S�B�~�h�S�_d���xf]T l���=0�����i�����`r��1�n3�xSS`H��O�'�)��>m,�:����N�n{�1�Ӵ�Պ�6�������<�L�I��gm�u5xG�"m� �&�F�Ѐ@��L��ȋ�W�����A�Z����܎)BF���WU��$?��PQN6�5�p�y�L;�=�Ԛ'�M��߭����J�NrzZ�r��`�>�����-N��Goo�ܽ\�7��Lo<��O�4�W�����K�>m�.��7���=6F�z�佘���b1���ս��S�� ��pe��!	m�(L��!s��q7�AD��9�Nkh�ҋ�{��n��T}�]�(3�V�)��b�-�̪�F��q��|�E�M���0�6���o^��ip۝d�"Y!�Q��.15�?
'Pp��b���-�b">|�c�����G������b��zx삷�^n@���>��N7/��s�_��i�#c��(��|������)I�#*���%�9�q������w�G;�lQ��u�)3I���n�pl���/f�������/�2,g�C�T�s�WN���<A��o�O��gN���8�m!s�� ��X����5�����JZ�X_TU�(3L�'���2M�)�̩��6��{��"��%�y�Rg�sp�?�;�����[���'��2mQ�vU'�ے$*x��0FP�/!�⢄�&����0��# �^��͆�	}R�9�j��<����WW��3��^N��,�	E��O���D�zƫ[��Aw��3^����C7�m�6����p�p�9��J��6�7���S�B��5��+@�h�&��������D�l/��Y\,�w���'ԣ349��]|����7M\
jG�K��6����6$z&=�"�e=�#��Y����x�K �QW�]g�Y�W{Д['&��6��Ϫ�D���J7����V����6G�4�Y�K�N�oo�|N`b����������(ߧG?���5q��ȪZ��m9����=OJPJ4�����瘓�c#J��̶'kX|�wc��j�{7�D��M�Z�o�h1Y�	�.�Њ5�%�D����qk��J�9h���6Q!��@g�;CB�p2)���ReH��<��-���r�1"{�2�4�!�'-"����!�wĄ���)���njؖ�Z�&7�#����!��е;t`)С�	y/'�툼Jl���/��"�Ě-��Y~���r9��߰<��?6hW��VE��?a�U�䄔s���{�bvp���cl����[��BMq��O��|�u@n\�BZ�H��~Z**#T�����v1��.�\Q�f&�JX�:��b�y|2��Wdj+�m�+����̘ݟ��+�H�4��b5����w�2����>Q%�7�+CJ٦8��v3�?���gLDWW�=tGm����FJ��S���`f]��9���*������4䛎�� ��ʶ��9�U@������WL��*� Z>��<��uů�tk��Nǻ%->�EG��BP<3DRZq}ydw��ώ���&����i�wu��x)P�(����L|k*��;���|IjA�g!iX��,��o�F�
Ϩ��O�@�EC�	��x�	!@8�Pd��ė�i�~�Z����rM��T��@ҷ\���g݂�tS����@��o�[<��o#��$����yT��h{:y=L1Ic�60�e,��AL1:�&��}I�#��{\�z4��ZF�کC��:B�<�:�zk��G�)��	H��e��������0�Ԉh|ʖfOi�	��8%����M����|F�����_�a����0��u<�*e6�཮'n�7��	�E2�d�<�LXsm����lR�{vX�)_E���(��6������T��~��p�<j8w�ic�熙=+gC^YW#�ݫ���|�����H��|��+�׏�M��}����!Y��1(|�B���>�f��i��vc#��hY]�ZJ�0�M	m ?J�e\��N���T]t�J���_��x�qG���ɺW��u�^vl4��
�?N�y����e��8���g������2_G�q
l���Å��!$j$�
V���\'8$���e��T��g���Q�aZ��H� ���Ax��P���_g�f�l*���E"��!>��Sf�Ճ��?dm��Ge�E�A'nD�X��u�O�G]O5�z�_�9��:�)p��ɇN� ��Zi\��
�<g�K�z�&s��U������l�<��+ld��>�u��ƙ�OkƬ��zθ��VZg��8y؛	���v��J�A�)�?��w�%�����Y�L���ykd���D�_T��MW�ۆòJ=�p̞)���@b@��¡�QP�Ȩ6p����-���3�^�s�9̟h�@],�F�~��ǒ)�%\�y�Fr�zO!�3.�
O��ԍ \tf�Ej8�y��`��J�?�^?v�4�naٹ����0�{��Rv�pS���klQY 4ȯ���"���`6��鉿����U�dk��w�*wUt�	J����2���L���:��4B������S;v�dh(LN�Em�'����D�[G=��~��U�պ�-Tp�A��QnqMK�x�i�z�lϰ��G��Zm���3D/obK?7���D�6��hd��u<A9�z�����Ʋ�Ӗ*�=h����"(��R�71�B*�H��D�Y���Gq^)li�Hڦ���o>�}�����$+��h�@Y�9�g����r�������䤝��Z+czt�eYb�T��b�)���PHv�j�o�ee����l����dJ�`�I���e-�r�Z�]�̫}�p)Ѹ�Hȴ���K�~�}3 ܷ�zN�:T�Œ�^�K�AX��T���G�*���50�6� '���`�k���s	wi��wq^����}�.�*�p��#`���·�B@K>N�<𜱈�(�y{�c����?z�{8���l�13��e�����~�b��B�~�
(��ｼ9��}���Ŗi�x��,�F�M���!c���5]���W���<��-���t��q��K�?��=��2�;��iRJ%��(�:�Yi�M�&�s���x���?�Y�5 m�hOX�76�O��-���X)3���ʂ��=%��c�%��t�u�F����g����@A���R;���>���#��~o ~"Y^�����ES��OtqJ���V�#7�!�-u3�Iw�sA��Ճ�#K�����yɂ_0������ک]�p�P�FB�����2�Ȫy%�fW��
D��Χ�k!.���Է�����&)��m�����)�	�[ا�N�>ݱ+�|�w+�5@)~)�t��7��P��rW3(ڗf�4U��85�z<�� |Hi�zK�����%.P�᫟2�(�;~�i	��z%����x�ЍC;]��s��l�&��~�4��ͣ����%�f�h���8�#,��}
��]��;ޏ�g�c��c�4��^�^ň�S��)�Z�ULr7��S� 	6)���l�H\qv��-��S�q4��U�Ty{!�<�k�3��
C����_�|`0*��!�Q�)]+vpz�_]~�AqRͰJ5#4�$QX�3&M�\�ey������+��wE@jX�E��ē蟠n-���R5oW��t�:3�Ef�k�_��^�1���c"_�n��Yx	�>��'�=ڸ��9���t���`
q-��Y0���N"�O���x�%+�ڱ�S�n]4Vʅ9pZ8�d0� �B�`���Cw�p�5��/2��^M����.����0��wN��K�C@�K��}[3^$L;�&8%"��S��B�4�b.��>�ut�ܹ
�⢽?�,�����;��!"��� 4��b�W�7���v(��f�I5�[4r�O�c��d��7	�k������D3�T��,��ԕ��;;^ �r%���=̂,N
� ~V��g��	s:=�%-Z<>��F��âȢl���#f�4�b�{��?'��:�h��P8�3���A��������l��O𑏹R�%_��=5L&���O�#�>�UI^�Ĥ�FR�[r�L�K�p���Qa��G��-�jcD 9��� �TQ���M���Q��J���+2-]AW�~���X��P�~�#xe%�/)�3��k�5j�Qq!6��W�M8�C����Z����O!��i=�Cŋsw��GД��|k��DW!�\xy2��e�s,�[��"z�Z���#8	@�z�4�Q��'W��qYi#��8�����S��S��Ŋ����c�jH$�{���sY�����_���H 71^H��~�t��:c���EI�*�~0�PfU�K�Uܩ��/���՜7� ��fw�ߔe�pX!I2ęB�c�Mq5&�?8�		Z���W��8�V,�ŝ�d��e�z'�0�1�����Nl���{�@l�e*�5o9Mf�Ӧ�q�T��!бx����\����eC�UL��W�`���� >t��2�<���bbλ���a^j�j'�[����|�v�ȁ}�G%�>�a�<�(c�}<��RRM2K�%�|;&,�(o�AA5�Į!b��}��#��"+�C�Y�l��w����V(�u7
@�[��\&RX��A�S|�;�+���t���pPp�5Bf�W���ٙ�H�&t�K��΂�����vs0��xhY{Zӯ�1-�I�_A���
fҡRc #a㾢:�V�ы[_-�����}�yT�������\>�"B��]�I��9&)�v�S�����.�AM��:<����3�P��1��km* �L7wQ+��mM_�J�WZcqL�������} ^���}q�>�ـI�-%��ϱތ��{����!>"�W�(R���եu��#k1}\�jw�D���$����*��Ś����B�\/�4��p@~ce�ٚ#漟������sWǅL�Ow��H/��-�JK�Z����7��6��*ew88?{�Ǒ�ɐ6�r���밶iV���gn�������N�G�KO �B��� A�b���CmE+]V:t+��j�M�')L=��� E�L����+��Ⱦԃ� ����6�Z�+4+�K�a��n�oɷ"�t��� X��-�`�V`���Cd��`\�	LBCH9b��~�c�f(@}+��}3x�����S�t��?�{k��'~3��6Y�
s;�=��Qt3Q�μ�H˓��؊�|N1J�5x0"B9u������T|Ѡ�''�O�O?&��g�wG�M{�����=�<�A)>�E�;_|�~���6m�V/�wR��L�ln�6I|6��\# ��sŸT4��������������μ44:D���X������[-g��@�3�O@�_�[������ߟ��'�9���!_ ���U���qK���������q��f��j+�)��ú|:5��w;��j�O���³�/:H�!�d��ځ��� A�u�`���Fc��y��?�C���ំ�=�����"�ӝ����I�\����)-	�_*�xxk�$|����9X�&�ہE�E-E._��U�y���_܉�d
���D��$~/�L�ZjOLL�I9�<^ p����h<9"O}���Q����#��ȉ��*69�cRB�Fش�D��»#��?l˶Ű��^�x�\�B�#8�%�;����� �2�L�a�EI���h
*�$5�TT�g,��@�6��K�2�z�3����#�?�E��<�Z�t;�V�fH����֌u��!��#v��Jla��l�[<�l�y=���k#+ :r����i!�s�X�Q<9}pc�T��@ޟR���+o�q@}>��^�j��*jFH��\R�����{۔~��{�VK�<�&X��o��������J���C.ւ�x�YJ�s��(��@B�f���r�
�@q1�/�2��0�S�P��:��.�ķ�w�(�qD�K҆�OfP��z��N��Br*�<�T"ػ[)��,CuV��u3�E�9�s�S��Ғ�q�R��#ϖhX���V��1d���������}f�	�g��*�]0�����'o�����d<B�g(��Re4��pbx��4�{�B�<X���s�LV7�;��ުYנik��)���VZ��\�ېq�#�#��ik	kK����l���������N���:�0���L�6Q:L�æӞ�H1�Bq�䒢�oL!A�W0&�za����s<�N�gE-�I��[�V�HJ���|��~ܢ$M�b(�&���W�V+Tv5E-��?L��r��*;M�v /�H��WH�$��9q�wJ�o9w�i5�p-�C̕&�n�Ѕ0A���WWk$=��'�����}�K[62�PEFё
�|KZ&�����-E�h��c�R�.$��<Bl��~��|�~�W���Z��ܙ�����%_��Y����r�+�2�b��l��,p��q��V�Txu�<�4f?6cTJ�T���$Rvsa:��NX:�rӻ�=r{��-y>4��$k'~�d�<��A"��a��X1
1����C�/��Җ{e@����!w�-����] :��nT��x�k���sQ����	��;|�W"�G��0�8}%��� o/�a�P�;�d�[I����-��~�͵�6�Y:�� ΢ɶbG�٩nS�EV:�Y��f�>�9���`���KP�0��ҷ�ou��s"���@�V�^�qw�����=7�2-���b^͂>�T-ܐ6^�_��(��F�ı����#����y6�}�f�p�!����a�'�M��Z��7�f�3gX+:I�wȠ��5�6����>Pل6nd�M�����oj�D1�D�TP�-���F�#Y��02���l��ۼ hH���^�n��/��e� `mpޔ�'��@��w=���.f`Ź�Ao�FQ��-�}N�z�GCY���L��s]Q?�.I��PO��v��}Ma�ZwK�C����]_),/�WxȆ$�[s�{��^+o��S�Y?ߋ��j'.�Tͧ���V%pv�S��! ���Yk~��o���j�iObpn�773T���ͷ_}�58����M���5
�o%�E�r��Wj֙��_� �A� �N:TGՆ�e5�c �����`T�?ap!`@rI���ʣ�.��S] eq�c���-DO�\��8Uǰgx����߷Z�h�+g����86	飵;�g�v���i!`�������c�&�v~���yz�|~p����:9Bu>��5�����8EIrU��g}i��󛫒t~ఓ�H��z�sƓޙ@�a���&=]�$1�8���t�:r�Z�+d�LW�*H�=(�"[:�8�q�مO�
�%�d��Ѳ�S�Y���������Tpץ�1{�>��D�k%�H����X;d�2���[�@�,��3KA��D��K!8�n��
��f=�>"L�!P���D�Yo����|��ݍV����v�V��	�:���kb|�dƎv�Pa��_{όӻ��kN�tQ��P�q���� nޒ#.4F �I�SqL/��� �1
?�H�3(
`@���rh'�~8\�MA5|�ٞ��^u���X��e�6b2Ԇ�@�����~}lV&N��y;$���u�NS��bW� )���k�b)o���&���Z��X�A�'U�Zi�]�����)H�/��U�t×�g��o=��r�Ԉ�\ն"f|�>�Y���95`�6�'�3�-�o����*�_���-�J��L	Cs�7d�@��%��qD���]�/I���r�G��Vm��1U�x0ġ��9T-�&�������Ǭ��4�Z,���W�Pbt�� �V(�������`ć��Q!r���p�L��P�O��FCl\}d7����yK}�	i�I��4sV}�W���9:�ǫ�JM1U��_��ar���&J"p[Kٝ��J�-A���0F�f(�����x��kM�����0x�K���%W,�*�4؜pR�*Xw���������m�?�OL�D��-�B�?(D�o��c�be]fpJ��a�Շ�&�-���i�gfl��`,��僱�V9�\@�E�5��9����C5:�b8��5#a]>�ZH�!���S��@�$�Ke����L����2�[=�@�ш1�Fƀߟ�u�'n�Ry<3���1��퇵����e�fr6��`O�9�������K0gѦL���,c���iC���j>݈= �P�+V��/k�$>��q��#;�� }I�r�ڽx�q
j��1m�����ũ6���!yc�}�s�	���\�L�K�G����2�|> MS
$ǺA���^��6�7�54����;p��J"�=�4gQO����-UL*Ri+AD-��{�9/��f��WEhBS� i��r����(OAR�4^�"_|���#|�E";�R:�~ؾ�m��(C�?��C>�Pv���
��o���S<�9�7���}ǸT���ܟ[��k�[=%Z��3�-h`b��y�
R��v�ĩ�� ��Q�\�1��yPE��*%���sd����X��w���m E�C�4)-�a��z.`]���:r����^o�b+��
�V���r�'&�|u�M��{�V�+��=�A�	��+M�p଴�S�5X���T�Yp�=�`�oN�4�4�\K�^n�ғ��_�I��w[�J��l���|���{K�~��2�`:���-'~AZ���������mi�>�1{�&DZR�|x������	'F�膑�C�z�u�JV����-:t�.V�/I?����؜Mv<��W��Y$�.��H��t�c{;m�g�K��=���x�Fk#�x�(���`�P]Wz�VG�B@�I>�����U�J��(��I~<�I6}m���,%�e�c�_Z4���$�T������T�)�������5�K^�5�IR�*���bN��=^j�kC�I(�F���SO®��n?f��N�ßK#�J�ǫ�5��`�Ez,vD���W�
��u#x���\gQ�n4���4�;����ǋ�'w�U�."&}��d��A,n�R���Իi�+���;����@ .�������Vyl5�$@>f��2\���.����ԝ����~"��;霾O���&�S��\/x�ႇʝ�{�t�2��Ў����B�v�Y;�4��1
�vs^M	�>$Y�:Eg۠�	͎g ����M[c�~xo���6�O��CdĺP�;��\�����W6
f=C䅮Иz��"�3��L�;¢�3��=��|B�Id��g����ņ0T�EM��E�5�$�FN���]�J�D����[��ɚ����;���.=�S\ª��"es�6�G�0��]�8�q�ύ=YIuc���Mq,���b��Ӣ>�6w�r17o��Uӭ�Du����Ҧ))u ݝ����x����N�Ќ6Ly�!3>h��1W��`�"�Tw�mX���a��_��n��R�WpUlD6����+���&�R`b�3�����2���9f�f��6�E���I����dN���G�>���GYG�OȨ��2/SU���O��L�����噜�$!B��6�t0��+�æ$�D���;���w��������q�'v�7�K1���Cq��v�v����P�@Ƴ&�5����g��#�e�XC�VM���f�$U?Bs#;��O��#i�(b���D���n(����D�	܈�y7e�N��Jr��9����R�͸A�#^����f ��Sj��?�]�{/O��W�zm��TG��v^�g����\~O���������4�7�m'��1/N�/Ě��%�WD�d��#��_"LW���v�o��YY�*�v���3��͖]���Ϸj���k��(FU]�tf��x��g�遞R���>Z}��[�!����9�԰a*���k�il��9ܗ�F&Y�\E1�h�N�K7{d���Já��H��D���#�@lt����ja�e���3�aN���\r���/��x�lj�=�����d&%�@Yhin � <�}dwђ��S��Q�X�g����ۡQ�+㸉�"î��vi�p�P��:��'���К��<�	Jl���� ��-���N��pY[(���Z?��F�W��]]l�����E��]�R�VN x� �hc�R�d#���Ө&��V�t���r��	��&��rT��4���q�t�8���"�����N0m���ݾX\r��)�Y�ί���"W;4d����0���4�aA^��K�y��썟H�nۆ�U8�m9hh*�W�-]4��S'��T<���\�_��?�'k�O��f�gm���#�V����7�b�^���T{�����3��Mܔr�Q�6� �e��	��p��y=���.x����DW�����os�ٖ:���D5s	7j� �ȏ�����t�a�w��� /��Ԓ3��/L����H|#���r@��Z�Pc��%��2^��"��֊��r���L.2rXp�yt��x�ݛ�kP��� ꩘��0ñ��@�CT��36�<S/�M����#�Ԧ��[��zȲ^#�,5�2xNۍ	�L<���e$�qT���[�ު��å�n�`ݓ����oB��=�9��e(�憈R�E"��Ӊ��� �52�԰�Ԯ�q�7쨙$�S�r;�;W ���q�{]���t��9�Ge5���k��h���(Ϭ]<�y*��[܉T���t~ u��ٕ��w?�s���D�׶$h��Fd�D����ؚӵ�*Q��14!9����Cۥt��L360�hGc��ȋU�l	�,��1Hd�g�#]����f��f���	���@�1p����K�����)��ʉ����+<�*�	@�	��Q���i���MU*�FʞTu'܍8�&7HQ�JB�q�a�����KRi�퉡r	�ސ8S�����Cgk��n� 's_K�a�����s�ۥ$���+�^^Auj�Ԟ�7�0�O��C��+Hzi�q�-�%X[�m�S�OkZܦ�Jf��<������7#n"��M8 D�I�b�見�c��������� ����ؿ!9���	���>y�51����XM��(��H֟�pM3:f�ϖ����z�6,��ۏ�,GI��L�Lw=h#�56��u'/�ϯ���m՟'2�b�SY2c4B�݈ɔ� hj��� ��ʴK.��Ɣ�d�b����"H�
��A������5�ȱ�S*x�~��c"�qB"���ːfo8s���ʍ�6�܆|�$�~��$�T��4��$�(ӌ�����b�X�)i�W�4�{�`6}c��=���'�����;z�A����z�z��%���`}��(�����/#������t��+s�u�V-x�	
@�4x�q�@EH�Ii�
��P�[�iL�4f��7q��ֈ���T�&���R�c�P�K��b��ܾW=^�	1�B��V��\�~2z�R���&�����V~�D%s��;ӟ�а@o$���[�*]@@��^H�����4E�-�j:;Tc51�����њri�I��y�T#>rDVb8뗛xHMH�[,�� �7�Qe�4��˩?�"P���{���١�k殜��R�Av�iNj-Vc)�Sve�D���]*p��oJL��Fi������M�|7����xY�9�O8Ԯ�XJa�K*�٪gՆ5&��5���S�������o����JFZn]F��m�D��W�W8��%A�ɹ�:-�k��ݵ�;?�*E�X+���x>�<QDs*܂�F=J�r�n���қ^�%ye''e	S�f��,�Yک\Q��VB���#�CE�؈�1)�4HD�[q�_�{�g�1M%8hᶯ+7�e��SIfN�Q ����T򰊌�2=Q{���ȐVp�ۙ�(i���2ƚ�&p:�M�)��Lw��3ނ�ك��l�(x��4'�VI��~y`�
�(��21�W9��jFkT����G�[�YĽ�J������o�_�˞K!|�̫xq'����S%��'�[�JX���� o�7weM�`�+�/oBL��j��M :bݼ54�����:���6�O�R\y��Jnz/��;ʥ߽M��Y;��qz�f�-��-��Q=:v�f�$�]�;�`G�4S3�F&�qX";\є�:�'��Z�&P�]ݿL��5ۈ6��~G0�y�/\?�%F�p���w�EFK�UNzq�
��+֗i�]����ė6��G@�A����a���<������84�U�*��)s�#������(	#(c{���>�����W,C\��Uov��~�^�]���I��L�TN�y�X�n&�	Z���!�d�2S�}�D�{�����0=Kb�]��OQiU
����<F�	�d�Y�F����5C��l�!���rW������ӳ����)w�����s�S$6np+�e���%�yrׯ
l|�D.�rA��e�4s�Vq�4]x<�N��7�y�]$ۤ��ٸ�N[���/R. W�N�eB5�<����������\Z�O5�Y��8W9���GYO�$�Z��r]6�+
�g����I�N�Tx�x#H^p=�'�R1R5U���|�lD�;��#8�BД��=�>,<R8���6��!��QBF��}8�����(�\�ܐ�@_��~w�f��-=F ,��))����d���Ĵ���)�o�� Ȱ�^�n�MB�sԪyV<A�yj
F�WQY�|�x��Tl��&K��f�Qs�6X"hb��Z��t����u��S����4Hw�#��t�f��Zc����B���"�lV��e�[�l���k�,�u�{��m�D���eT]�Xtט��h�K.�"�����<��Vu����@[]����8MϔV�S�7���!�v^��Y:��'B=��i�~K������n�K���<���D�V���mҎ{�\���aI�%�Ay��ⷍ��L&���p�|�m!:ԑW�|�ʸ�O�y����M��&��N��Z�a�(^�	s��
�&5�	����I��BQ����x�Z��8v�H���s��e3@�GL}_�J�_��X�F�I5/��r��ֳp������$M��"�@1d�)��툟�"TV�pz���|;]V'�y�c/�P�D�Xg�����{��ۆ�ItO	��������,l��F�8 �P�EJ�^c�{:*��;|uL���f uj3���\:�>�4_"�o���Q{x�c��r�j��E�#�<����};v�o�O�齂 �X;��/2��*
��P��;h|^�2�.�N#$�$ڕX��$V=�'N_�/ �0LS� �����V�u>�种��u���0Y`�遮���uP�j\Z`���Et|WƭD<�O�A���Ԋl��[SgW�3�"J���!�\}ˋ��FZ5�i��������[!���G��Uϵ�5��R�,`�x�K�6�Y1�e�g���tf��p	jG���ҹ��jO��x�ݽ�g��/J��$����S�f��m�K���F��df)�Г�t�%�*^O7s��GV�q_Kd���H�~�1�ȫ��<a�&A-�x�&�0N����N_����ml�'��C�+��:�ǿ��v�f䲂����)Ӣ8��'4���}MƜ�"x���<�Y�$K�|`��e�򛲧����-��!���r��Wp�lW���H�a?��B[=�h\J}�͌%����B��v��#���\,C�ܧ�����oi�,|�p��B���F��Xr�ҳ���*AZ�m��͕��l���9��A��1�!�����#��s�����w
�R�8b�a�u@"��(̿"&j\�� k:'�*4��s�y������7 
, �&.ѐ2	�g4���˱m�������&� :^dMQ/į�{B�֫�;����k��@>큓E,��g���XB��t7{
���5,<M�����k9�KN��Ae��yl^ٍ�g�3���m��^^�%�����^l怘S��1���l�n��R��um�c� �����^�w�]����J�^��q78W���qT��ū재p�h�%>Y��k"��>�7+�q/>����x�!;�9����SB��|W/iuֹ[�S:h���[�hO :'���� 5u>η��k���$����O��뻖����:�@Sm5�ͬ�W����}6�]��AMe-�R}!LN��(��:ƇJ�,Ar��m��W��H&��mu���OྡྷV�[B��/92t9{z	�7��@��ֈC�s�"�޸���J��p�!��`�ƥ7�b�4�A�:��� �}�B���卾">���|e_l�ޜ0�-`D��A�9C��J�tz9`�Nw#U�~��\�I��2�DЪ;��]��ᴣi�G�J`�+��uk���C�BflTLR�~��� ��x$�v��YZ�N6>���BpZ6|ֵ��LR$?(���8����@�5���I]�����
�?ž�ᐞ��cF�(�ڏ�0��:?�[x����e�/��.��gn]
I��4��řn��D�Q�ʅ$?��6��S�bH~m�bt  jh�#~��{��t�d3�݇��B���U�7��;7��<����#a�����Z�!|̅!(�'He�9�~ `>�
��g ΃��5"����1������u���k�!m��E2��{���A�f͸)[m�↤��ُ?��|�D�(C���y���۝�_A9E��	d��u8X//M@M�o�(}�S�-1�"U��T~���PA�b-����[�yp��O���,8�ؔ�ӆ%${_����Ѿl�y�+>���c��`s�Ģ���,�)�_���#�#��-8�v���ЌtQ�\
00c��<MP�1�6,��-�%���f��aɯ"��}�W]���Z��s�j�
Tyj���&�}`~��O���nc�͖L�$��h��[+Z�u����]0�����'�v��Ǣ]�N��c�)�� ��?ߌ�K�ne�;E����M��U^��h�# D�W���y��W�|xӟ��E�y�ny�D� �����f`rS������� 6&�=
k�hO�%�H��5�H��ID�0h\�_��j}�r�`�������/Ka���a�J�����=����P�߾mZ<��3�P]� +�?^T�|�m'���������7AG�������5�I['���ʌ5]�Z�(���-<�R�w�|i
�Q�	������)F�O'j�쮲�A��(��n/]
������జy��0
�{�r�@+V�4�Mf���	�#�o�{�0[c%�q��\w�<�쀑����^o&�Q��T�+;��!�ϨO3�cxU}��8�H�O"��p-p�C��������7�{�@e��?۷���h���x&���[���:	�mM����:1�f�MXȧ�K4���ǐ6'3%�G�'?��-�O��<]BH~o?]�mU�ZJt�����(�H+|!Wd�G��X®����FZ`NL�&��>.�Q��p���u�9�"#��)x�?�@jj�͢���b�K�Ve�LC2kՆ�������r��W�|�?8_`�ǘɠ���%�M�/�@<_�0����@�}n�hT*�O&c}�fhs ����b޹��o��{l�	���� ���֦���,�5J���>�qJ̛J�Kf�;�X�8�h�����/���bn�-B���g]Q�{08۸p�X)��'�.�W�覆�\����=:H\�^,��@�)-HB�Kei᤻ZZ�|���"�A$+5��6kҒj�XGrN�7ԬJ�oI
��� �!�>��o�b޵�,�V{�������v�� >G�����M����=��.�Kk��a��|��|�X���~fbz��3cT���\!>��F���Btw��l�c�E>��\ӹ���6l����/�����/�ԣ�>�̌4u'#��s�(�1{/
�֙"��5�y�����wu�S��,��'s=>�d�7�����I�U�[^�S�5J�Z���ZW��I�;��
 ���puN%O1	>m���=�"�����!��<��rY���L�ƣY�Pi3TK�s��MX��3��JVI�	�fd�j(�?��m�CG��*�F�Lb����5�ƆOr9s1j.�N�T�d�h��Z'���0����װj��^ ��J4LeH\e+�z�u�a*Ek��˓��gi���	��+���`��M`�"^�v�>殠�*��|��XH�qu���	�����2�.�Yaw��z���U)��w��M�"�C^ug����E��o��E�=�fO�*QV�ZM��
�g�3#��'o)�o���;T?��~�C0b���T��Ӡ�2��ˆe�Q]�W����3$�fI�h�%a���Q�Y�?������f�n��Y��oI�����FW�g�Ƽd��'D���%��Ӆ���L������U�D@B�|��B���Mr�W�\eH�S���Y�-��j�K��>RN�U�B�Q��T~)�ݢ��-��?zňj��q^�¯wK誺��`�'�~J�O�-z(�o��������ҳBLꑂ�|�ٜX5h�VG�3 �o�v�x�)F!����#�ir|=�"jؐ��#�r��ѥ�:Nzц)xA}������HJ>�x���Ю����t���r%\ۂ��@�h2{�]nRl�6,��;�~�D���
��X	<N<��lͲ�dl)/3�&�Q���L��IԒf�B�p�K�=D��d�Y��n6�t�ǝ��0,�֛��AS��I��I*�Mqt���Of�px�hq�XJ3t@B��{��d�˞��h\�N�6�6��*Z^�\+�=���5'�i#�柴�\�cLBگ)�Jć��=8�<.����V�%��/�*��	eX���$t�)�Z6]d�~-2�?�D}L;-\Ae���ȓ��L�Oy���=�7m�]Q�Y?�ա�������yO���^й�N�]�@�m���#И4�p�&�v8�kǀM��qy��T�e}��ۘ%�o}�c3�g,6�M�Kɑ��՘�|��^qӃ�
;������@ |j���hHm	ԯY�{��	��3��U�r�qn�=@Pc�c�_ ����c�f+�G:�(��VT�����%�\(9� ���#j	�(�,��&
�0~�a�u�s�a�A-�/ Z5���z�qX����ǜ)�G��`A��jZ%�S]GƉ6���m��m�ޒ��B�Z��/�=�=M5'4�8��r���~��Vd-J#��HI͒&,���A�b�a�VeB�c���<��mA��p�Tl��Sp��<��v����?j�0��~����J�d�N��t�#����3�$w�'������V��䉛��4$LJ�9AV}�U�H��P͵B�Z��tb^�$�`{�P��={P�04܋�npm���+��BFРq�A�FzH���H݌�z�~�������vu�f���X���IE�:�u69��=���%���o��>⊴���p�_���{́&�6������Utn�kȳkV����CMiR�D��҅c�^r����Z�,�J�W��
�9�Wg������H�W�A*PI~�]�*ѱ��)	L�E,�U�~��ڹ�P JA��D�PW�E�w����a���g��,��t���(Aw��c�qq�u	�NU���YJ�=����V&�!����ޞ�WБ*:��]��F\��y���b=:]߉3f�pn ��Bl��4� �������u�J�\����b�%D��3�g�S =��)/���Dȏ˟�B�:=�{q��)��@��6.5_��s�@v^���~�;�
X"�>j(+����������/VPR2��;�]�'��LH@��P�3��_�ĽV�ߘ�� �T�Zd�����%�������3��HS@|��8�׉���?����0wYC$w^�.պ ��Ju�[>�8ҷ_�ډ�e{(ǻ���+�u��mٍ��2���I�[/.WN�/���86��&ެU�}A#�f���s��s�y�Ua�N"���C��v��VwK[ﱦ5 �*.=nc6awQ������ZF��O�H	&f�+�i�������g�@��	P�(d���7���C�.;�
���6	���g OJ�̘�<�H�?�_e�&�\��!s9�a��-�}br��͘��f�BĠW�Lh��k4ţ�4(�O���:,-�PE����4�X�X��Q��2�4��NL���%B���b�,�5� 
�ȋ!}�ª�Q��:W�o���^[L�H�|�&���6���<oVp����)Ϥ�x�m�LV��1��9�U5x��� ��g�r�	QƻL�`��e�����P}V�O�!'M �d:���'��*!id�cj����L�D+a
�Gy%�~7i�f�۹��[��5BUVt.(j�`<D��\�>G%2�lۈ;4|��J�P����'9{��SHv�"�r/|S~����d����:_t��_��Śq��l�7F���<D����C���0_oC�B��	��p%c��}1gp	��=���3%p��?Gx<�Rϴ��vLB�~c��B��x�k��v:�P�$"�1����}'z��"�x�,\�D��>\&� �����$��'�Н4�p6����2OK"���G�0�3nN�wFN[���q���!���WN�)~�v�]��cl�iޙ���)[�E��q���ʡ��\O�9M��y9@�Mr}�'7� �̑R`�hm�H�T^��}�a�
�w�k��2��U�ڤ^0���Hs	E|��Y�h����y�M\zx�:o��=0�o�r��J�8�ԣ.����[��w�cћ,��7e�-���y���d�QKt��'-	V��x� YD{zŘ0g��[�/�+qV�iny�ߎπ� �lH9��T��Dý�(1�>F��3T�Y��/̒a��������+�-**�w��8o��A'=偸���Y83ݠ6�q��ꇴ2���!OS3Z��N�eH�Z-������$Ԃ6���Ҧ6"�|�h���`���c�����蓹s�GV�i�M��U�~�*�nei��k�����ӧ�z�3��ϑ�1��+E;I���:������C�!
�CgE�2`��hG���ƶ���\��dF�7w=�ܑ�Y�4�-�b�*���b �۩���ȷ�*�pI�xj(8���O/#���Ͽ'�����$9��cZ��*G����>,P�px���H��֭e1&����S�)��$Q���T�!���3�Wz��_�y,��>ޭS���Lj�9�c�����QR+b*&��.�7!��\�Md�rM�*;���^r�6��/�{8�s?b�{
kI,m<9�MP&�Na�����H&~dXL/�a��H��QڼI���΁�������I�'_�0�Y5��@�(a.x�h�W4P�@�ij�i�[�E��3��!���5U� 3�Z��=���S�]ʑC�6����i��1b�f��BF�k���n�o7����&! �4����k$��� |s]/�<lw�sĊ1��u�5�L�1f�" {^"�E�]�`��[�
]���	U <m���E�LzL�������F��l��jj#����"��k�ky�2#��~M����?�]5���E�b�Ցkt3���Qn���0�f|3�cƊA�L�fn�]�����_�V�A���wTr�+nϘ"��eŏ�k�X�Q��������Ϸ�?���}�j���<吐�@��%�O�wVri磵s���)_��+aTRҊ�8���&C��2-Tm���6�go��}}���k0�y	i��H:I��Qh#�s�\�p#;$[��s}��̗����d�$�A����߱�n�k��V�:ȡ�`�?V�6�����b2���/��f�N�M>��R�՘�G�P��p0�x����[�O�G��o�[�N�2��B��O��4��W9�5�u����Ӗ���2��N�yc�&?�s(��Qe���?�̈�lԋ���:�?9��4t%�kI�fj��	S��BA,�uD�R}�D��7Rxm]&��ޕ���2OZ��U�ƩbI*��Z,v��4'nHd�W�c��.Q޸�Ű�̗^���z'��:�h��i���ͅ��v����s�8Zm�#\M�6���k �-�ߠ��>׊`�Z���Z*�	S��G%����5Qv�ɶ�v*#cQ��d�,���ϓ� @�|��KfL�\�;�u��w7��2�������?2	Y���;���j�q
*~�t�f#���4����>�qa���gF�}u7��>@��AO�����ڝ1��K]y+C�,�x=��n�(E��I����Kl��+!�xt��-<Zʺ���N�=|I;�Ld���^ā+�,Z©��_C���FDi��L�φh�>��\�+����}l0��Y��zNu|�wr?@x�[Ή߯d^i�e ۧ,bOh��@ `�[l`���(�#p��+�J^�g'�GV�5�L.�*�E�M��B��9��\2�H��|y�~��
OlЮ2\1
эڔ�#�3���,�����9��<�d�Rj�	���Vm��#��R�=+�M�n,���P��dzb�2��~$�Y`)�%z��ÔDJq
��5�a��pf�H�T�(��3ӌ3)�?�B��7g���δz��ȟJ�`���~��b4mYq�O�h�: &���{�*���־OVn��~_[����/�:��6���l���k�O%�g�c�ڽ��$<������i�(>�j��y+U�Vf���:-����+m�����X�:�<b��" ����b"�<��v��e�!uO0����D§��T�x� ��4���+�z�s��H���2��X�^�q�7g2,�Z/܊)�3�h��,]?R�����'Χ���j��|�J�J��}D��n������#}v_�����6�9&�#&%8P���l�a%^ep^r�NM_CS�䥔�W}#�=2��,���i�L���*�~�N�'�����(+-�A8
�U��{�Z���i�&�8�!wZn��K �ir��pEL��
|o ���İl�sa���`�t�?-�ɄT�XY�Oj9+�\H�M�f�m�ɺ�Q�.�k�0Igp��3�{+����x�dw���C�Ў���ZF�GȒ�p���!��WWBn��?8LɮjZ��҅N���$��k�#�$
܌I��z��0\�'��B�H�������;
��>���ɂ{���ѣ&�|��5K��>����-Qq�C4�V,[_�i��O�R#���Xְ�F���k?���qc��`"�:	x����s���z�����k��&�1>�rwT��-j�lLR�b�S!���*�]�g*�-�k���y+���u��eծUW�(��HǨ��ˢ�b��įW�������W��;�|u��y�\7vt���P�z�ˠ O��q��l�����
,���S4qO�b��(�3�к��_֨f��(��u�&=��KGŃT�JjW���5x� ��VC�ժ|N�����T4'�C瞮k)�(�'�	�w,��I�Q����	ج�����|�<>��X�26�4c�����s%=�����k-.�A>wi���jN\_],JV)��)�:�X�z��l:^�����I~���͊xA5� r��{������@�Ei9:��ZE(%�C��R)m9q4q��	f�4.����u,�Xѳ��{�xU������i�}��Z�H�{�cV?���1�`�����ξk�t���ŚɌ��Ý���r��ol��� g����� �����h�k��`�t�ю��l7���̏���c1Mz���A�`���k[?��G�%�$��6�}*�%���7k��}��c��i��o
`,ѹY��9/wqzN����;\���v����(� $àM���H+��7_��Q����h�,����k�b��������<(,P��VE�?��Fżq�[���ᘒ`���.�.�����̨�.#U5Vl[�<��#�e�Wb��2�����[RN�bP�(H3��ϧ2�3uǂ/Y�n1`���&u��|J�/.٬�x��_O��VI"�Nԟڴ˄v�
���N����&^0�VBz+U�[�8�Z8��i7�i���baʜD�B:>?1�~Q;dVϮG�A���k	!��CqR&:ZcPuѴ�5F*�z���u��V�Mi!���V����s�Ɍ��d_zP���P.��	�Ǯ%�)��;S(�x'�U|w�S��$�1�dMё,��kEr-Y��b��C�R0/[��zC}�x��)ĝÔ8����?�fd��8�5[�3 D�o�Az�w;|�	j?�9�9��͵~$��ݭLޡ��9{
�*��_�O�a'�c����}��9��mI�"�>/b��~e�L-�!0�Q�aԀ�u'����J�����?��n�%�)<;l��,�KϤܓ]�WU�u��f�m�� =��(aL����[H���6���I��Z��-x<��D_8TB�.����;��2�SEMWyC�P�iUYO��A)�CO�6��-�k>��*�aG����	�(��h�"'!؉/�j}S��(+We�,�� �=�h4=>6�B�J�b_����v������Cn���`A���G�Ƒ�'�h���'���J�_܆ם�4\}]բB�r�����>�9�鄖�M�n�3k:*�
�^BA����gK�C����^�J���P�����"�<M�q���h5��w�`��Ͷ�̟�!ōG3�>^*~�i���&Fa7�F;�{�-��m �9�<�|I���b���K
�â��2��F'�j(,���?g�<F	5��O�އV���O^.x���^�>WV�{"��x�
	�{��qE�`(��N���}e��u	�>i	f�5���|��`�7�4-��ë�5Tj�HQ�SD�Zzv�=��o-�׋��^-x���wܡ�Z��G�-�5�F2ʹ�S�"���&D�f"����%���V����^��lD��_��u�P�%ia���J��/:�ZwA���7:po^v�I܆���1%���=u;xVǅ��\��^#P5�ð�:Q�;W8O5���uu �!#��(MҖ�\䘽9n�o4���[�iՓgC(d,��S���KZqs	,�C�3�T����~�ҳ��l�{^1�sB���l,�dB�1�t�Ұ��� ϴʑ����%�f4�_��L�_T	�]K�5�� o.O�4E��$��y�4;��R\�1߽i䍰$�
m��?u��3�v�x9A]�c�2��N��L%P_�����ج���O��#�s�h�����/��땔����,��"ǰ��.�I:�&<��)q	�*H`�(�������Jc��2n���'��9m_)��ry����J��
�H��^���m�	�[�?s'��"�mv�6ϧ
���	�]j%k�m�F8�"���ՒJc�ߵv�����?��/¥���W]�ġ{�o�m;�O��/�+��eè�}p��B����(��U��J�����e�JYF�z�]����u/���=�N��û��
�����M(z;�9L���6���������e^��Y���;��ih�@���gXB-c3����Q&���RZ*!� j	lG�J|;����I�G��	�I���PҥOo*VQ_�!~�
�}>A��9�{Ӫ�O��,;w�'����l�>*��"{c�L�{9,��n2�9�Y��l�ãı �f��:kJ�|&,���!b-1\C7��"�A�Q��9�:��%��?^���:[��\���%�W�/�4���vu�.�(C��=�7GҿE�K-��%�?̮+����0����RY�v�O�:�jS�c���a�4�r|�R�R�<����m,����?��xT�8�V8�j���J�;�M��X�2R^)�E3%Bլ��x:.Ӈ��o���X(i��؁:���I���-�n�p�\>���OAL� �\j�x�F~�Q��5��Xz�?+Z�kEE �Kq-�}f,I���R=h�׮:���g�ʩw�l�]������} ���HͼQ�j�*	s^}��/펭��I1Y��Hg��^�� �����/E��z��%�/��٪x���iR�z����z�m�Y3���/2�.W�B������5�12d>��?��s_�<n�����{J�R�_-�2=ɏtɡ�2l�� D3!a�4gj�l��m���q9���R`���X�.w�I:fG��}�ߖ�����������^G����@��F'����G�͠�^h�->���o�3�'�B�ۖо`�JٯW����x�v�t)��w�[2��	ФE=�8��|3󪢤�'�_$�\I����=g����~��q�t�����4��rΜ�ErY*8EF����v��;���#a��tV��p�\�u���L���O1���r�q~���o���n1b���B�7vFSV�ҭ?�� ��9Rv �.���[��ֹ����l�E�l�yY-����J�WeDU�R(0����3�}��'P}�Jra��3�r��X��B�E_E,O=PW
3?z�hp�,�|J%�t5�hƴe��QZK�XQ���P6P9o9�-�$���m�It��6�m��K�i"�+x��gtOT��:B%�D4�Z�����և(��u��a��\78�C���ro����]O�X�}lc�'4q8Q�0�ph�'�E.��b���#�#�Gn�YL���g)�=�WR���JEE�2x�U�ǎ�~�p�M�T��`;��͗�6�H�������mp*:����CLn(HMnM��w*��n���Z�92�N����
4n�"�u+;��tƙ^�n\�7M�`�;����$PE�͇D��^�D�F�k���� F�i_8Fԃ`?pA���-�R���yO����/���PŌ4G�~axD½� �ߪ�D����
㉎�@��ص�4��f��������P�V֟RM;�t.�#ª�����}T|�w����M��bHw&�v�C:CN��� ����N�����y�/��y�+w�|�z��}$ԭY�xq����\o��B|�q�0xp�[���#��]9!�y�����Bƥ�!��a��~,�D��4��(�T��2F�]�Z>�>[:�`�I���?C�ؼ*q���2#AMuqь��Dn��q5�:���͋���a��Jm��>,q@�%0��DzP��P���m^�g��s@a�hk��E����� l����\����EAHҀ�K�$�%�Đ痣�(1}��ײ<�D����G���'�(5�.��	yaG
q����.,��R�y�_=o��:��#�XVFvFg��z�����G�[D'U��u4��2���)B{9��)��,�## Gꞝ�ҟ��a	��q�H�{��og5/F��&]�x�V4�����G-�;��ӑܷ�~hf�(��	
�u�%�k�!�'^]R[ׄ&�.� �%5�fX�Fa�Yl���V��e�x �L��`#V�r;s%�GۮY��/]�}�F���,�)N 'W]F���l�*!�
W�	�˰'��p�l��ց��<��H��BX�P�.�ϐ���bY��,��rE�u��MB����XB��X!"����ލ��VsZ���eI_���ѯ�*+`N��?����w����
��Ï��0�蘆1�5�JT�9�ހk�_�$��҂#6z�0��0��@���V� |��錘@�N�T�)���Q<VU�L]�e��~P�X�>�NZ&
�E_+���	o<H���ޜ�lK�\E�@/k��ٺ~��i��>'��n�R&�k&�����p��-c	ӂ~q�Ŷ;Xr�$�\2Ұ	��TzU�]��A>kW�N�ˈ�O�@ׂ���Sӏx'�`K+�.��ȿ���/�b�-껈�QTj���q��)+Ȏ�� �˪jm?
������T(�Y�4���x%Ć�I2��?X��ߤR��^լ`ឝ,����$�an�i�7+��Â��������������.x�����`i��m��$�9$�T��Fm=�s�W�5`O��df�d8�P�	-�"�W�׍L���R���됰H�^�G���=���ƥ��r��b}eƠ��n�M{b`P	{h�*�=d�\�mFYLS�^�N������"�ΠZ?��ƌ��H�Ǎ0�	�a86����o��P^���Ϧ��a�rѢ!8��vVO��r�����	(���(��>�þ�ăJ6��c�\��Ţyj{Hp�W�
���Q���e��>Z��J@>X���v�ez1���B�a�h���R�]�5ܙ�����/d��7w˽ި�X�������o�Ԑ�k���[ҠT���Z����	��K�S�8�m_V#,�3�G��t#S�lb�;�7 �+@�%,?0}����/��Sv��g��U&h�L�;�t��%����^�(�A8�ިE��U|rx���S����8�gS�d�Z�(F�Y�J��f���V�j�B����3/ԙ�=ʹ80�YՎ���v��2|QZ�Y�L�������8>z�R�
��`_��~�}��M|��.+���sX}70��aIK���c�S��
tw���Z�Si��h��h5?G��)l�loJHvHd.�d�P"#�{���1�CG+�%Fe}=H��h~���C�rEY�ۂ�������Ȱ����W�X��0�S�+R�k�D�R0O���c>&��1[R@��
Y`���� k�0~tn��DE��и�(0=�blQ�&�e�?�Q��8�� M�ώ��v&e-���&X5�ݑ3(��Ґ$�������G�k;�i�Af�aZ����Rz~����m�W�χ��O�vՙ��J�+���(\i0���������C�h�1v#B0�u
���^k��rp���fX�WJ�ʶ��L��(���q\OB�JkYѓ���T�IvT��V�|���ȍ�o��N(c򜸿3�o��M�3��I���e�Ұ�z
�l5cv#���VXSDSv��e�=�s�05���z\�^9�I�'m5t4�q�>~빗����I�k���g���VMK�I���I�ҳ�j#�R��r�` (���/`jE��|T$9�L�F�֠):hE>��viz#����<�� ������i���[���4�� 8�7�=ݣ����L�ՙ�5G��,�ߖ��`��=�/��jp$2c�8����rW"�#t�����Or�j*e3	�4v*zD�r suU�6�`��-,�4�ֆ ��c�]g`{��Hq��O������/@'��D3�V'Q���s�W��Yp]��a��B4oP��r����iӷ��d��&�X$̓��A�m�c!ڷ��vjLK�˗�՚4^]5P(�_��R�P֖����o>���	t�� !��~�ƺ�_Kw[��
1��*|��˖c��[2��l�~�����'�5B-��l�ǖd�H$�+�3��/�Y�T�4�)�	��`�G�?�Z���,�Tl�;G1r�f�$[8F�f|F<�E��W9�76 ���'e;C� O�"-��5�_���� I�q��,����-.LQ��-�!r.#��1��1P�Q���!!&��Vـ��>�
��s�����e��xW�8h`��d�f�0��ݢbH�=�:�m�'��M�Dv�7��V�y�@Ƿ�Ԣ��ܘ�/\r���O6,? ���/� ����#N�|b ��g�jǞ�ͯ��׎� @��bH%D)��rT4���@�� �$K���7Y�ս���ՠ
�b�+vI�~vX{|+^{�w���)�^��y�\�V�,N�c���MI�1�>�Nֹk�����YJ$e� l�L<"�PZ�i���=��e D`i웣�!Q�L�q2�?I(���pB���+br-H�.I��헹�.��V�ϐh`��<t��oM� aa<�.s�ȃ���9
�<�>7U��Bw6x������pf�+��o�@��vY?�Z� w�
l�̿����=_��5щ��@�}L@����rY��l�[�~����M�I�m���n��)����3�ٍ{t�Mt��;Ш�>xA_��4-���5�����hO��s����m����&� @x�#Oa�f�4�>�>��N�?��U����/ BɥG�Y�O퐹3��S%����h7؃��4�IS�|��7tkQ-�`�������OB�|yo��)W��]�0�,l��z��K���s��_��a��B�9������$&'eJ��^M�x��J��&k�^��xc�eTHH�xb1t��x��ʋ~פ���ٖ�OB��No�NV�E=TΛ�c�A�0%��ǜ��rsi�H�[gS�~[�ߊ�Ԭ%�٩;�reȻ��@�)ta��=���\:̝�9���bs��)9������F� �����vV���V���V�����虜W-X\1�l�zi"� �}h;\d�������㋙���7�"�P4��h�Մ��u����	H�S{0��Gw9� �c�7zDfC���Sb��׫v�|���[@��3gm	)sp"��3�yRO�I�&����v�m.��ʨe<2@�u��V��O�v$�MI�k�E�m�enk�?�(����9}�f���{�"��
��ܐ����&`F��s8́���c�+���c��G�i�)�w��-y�Q-H��VJ�Wq��E^̒q��3�!uY�u]��팗��7J�_ecaˇ����='�2k/�*��r	���O�F� �΋�BG&�I�cu�v0�q�E��*�2��6�3�X���s0��Up�8��~v��g�# gv�S�O�J>w ׸�5�ha��^3++�>/P:H�^g�� V��GR���%���/��Z���q��yN���V�]
��#9$WԞZN�-hY��8u$��?+��YK9�`�Y�E��gqY}����uι�2�艢�߿W:uӓ������b�������ʑ�(R,8+��V�����J/@��iv�[ ��K&���X0������]��	\��ј�
b���J��Ȅl��8}�5mk�LOO*�͙�o?�t��R)���53e��Y�p�$@D�9���[l1iWE����Zh)N�*.�w��,����De<Q�m�ʚOa7�}b����*�N6����!��+��Yz�W�ph5I��l�uk�V>�nu�֛/<�Ya6u�X�A
`��x���k�	��9�lW�"ٙ�"�X�b������{�]
,�@��N�Ha���e��k&j���e��FND~H�9��W��0pn:�(�u�d�0v�R�M�Kʱ���%M�5�vݙ��87pZs�P���,��8���IqriP�Q�}��0o>���r
3�m���f��ɐ���vZ���xO�(MCS<�S�����#�a�l7fS��M!�QAl<D�1�+g�^���%ǴXt]{�x(���N�~�	��L����V~�O9����0�������*�y>�ټ3N��E��DzB�������s��v�w��:��-�\��%�pȨ6z@@��G��I��+��f�9�|JtgK�%e����o1�Y�a�%��SfB�J7���m3�<j�u2��4�E���#FY����r�?�=Q���m�3��u 1�x" �ݍ2��?�W	��~�ƙK�
�YYK��=�?���b�3rgMg2�L�Y�	��[N�ae�3⸞�/#����=��q�f�r�ٍ�*	lup���ۙ�-��l�@ ���o7��z���Π3kK\��k~��a5��h%��ֱ�"�38 �D�y3Ph�aԲ��.��7,�E,�'�m�����x���$8\��򱓎h$~/&�kv%X8�'����l�,y�0^�Q���ye���T�O7��Z ����X肙�1�ݠ�`��̟�7_����w*N��$�2��|��q^�5^F9׿��&��=������5"�M 7	΁V�mik-�����C~wyAM ��+ᯓ��!��PQ�x�.���Z�L��4���������lƄ������IX3�y�ӕ��+�>��3���#.Y�'+��i�_=�`�B �����R���4����\6M�$;^��#$Ǥ�[)d2XL��09̢��9t�y���&�FC�:�ݐ@�_���NH�*�^B�,);�S��	ħ1�5�@oX�q�'X.�� 裞��n����eL�PZ ec:Dd)M��7:���{B~Kp\�~C�����H�z�׶j�|�<���4��YB	�{(b�ς�����x%ճC���M��*hP�**,��Du��3����ٳ[�r �a�W�[���Fm���T�D(g�O	�F�
�Y�Ni�����l�+�>B�g3Q���s$r%�?k���E���~��򥊫�e99;�M�׹K>�`�ko�߳���];\zCI��\Vi��~!���!ju]����~�h��穜a���L�c��ɾ�i��轫ӱX�ǛZ�9@ue�������~�̄��?A~�����;X9u�{_i��A ��w<K� �16,g{��Մ��������6�m6�Jㆳ���5X�ˀ0q׳�K��
��V�T<�#Atɦ��ځ�?A�{�=
ߕF��
(�K�&�9�/*�[)�
�D<���P�'��vٌ������P>�Cl"@�s��G�S�ڢ�@��~wi���e)�?4ԃ$.��{-��8M��-}�Wi;��Y�t8�#��L	�:뿄�.>��?ۯ�:H����f��ir�s��|��w1nh�^U�_R�ϓ%&ս��v�����c��8�f�+��|a"ˢ�Z�=sq2N��S!x%Ú(r�g��r
���z*�'|o��j�љK{�=�|�5;=�W�nDE��G�8�᠓j�e5�I���"9A�'X@N9��$��hzb�z���@�H�PS�ϐ	��4��5rU�M�2B����\��;�ga�u�k��xJ9B��6'���(\ڵ�BG��LY�FJ<��>����I�)�6��C���>�
ե_��0Zէ�(������e ���w(��1�UD��%W�,�
Ȋ�����'�y���	箦��Q�i�	�t�=�>���^��z�8��M��!X��`�tQ�1�����o>З��R��C�2gZ���~ŵ�1��K�����i��:�['�ɨ��O�rM�ֿ�=�z�U+�Fl��Y�	�3O��p6�J���M/��STΛQ
	��P�rv������5�p���lg[3 L$�^t�G%L���Ti�tb�j%����CN��6�z�u�x�2�f�(#z%�iB�9���!�_�XG��O��*9�}�dʮ�?��[���i��T��G�+9c����}��4�y[.7tP7	�NAJU��<m�'��� ���(z�EƇhQ����߁z6i`eBh�Mf5 ���|�I᳸g.��(��'sT�RYJl��S~1��Fy]3@�iУ��ϟ��Z:�::�Y�'���>�C�b�b���R�S�W��穁�P�'��v\���uP��O"8�>��l��x��Ӕ�.�s@�������!��3�2r�~�g�3�V-�1e�|����~�ʴ��m�7+/�j kE:��4,�pu��g���wz�:���ђ�O�i5��:nh�7{ƚb{��"���
�I�҄6ם�+���=�Z�G�fkIL��<A{��"h��vN�j}�h�$��C��ok%d6H�8�J؃w��!�����@{��;þLJ울�M�$� f���D�D��5в�˹�:�QԹ��0��f+�z*婜R ��I'���*�"u��DL�b����RD�4ߕ�z�1� !3	�ǝ,�������Nl ����T@�,0���>5��"ږM����q�
��t����n��T'��4�1�d&���t���9'���sܦ 6oy":x�U��)hxl�j����A�i��[��t|�;�Y[uUaS�^,�0n�����}�U1&��x�`�:됥�h�̖oo�H+_BVтf����fH����T\Z��������y`S'��H��L$�,�� ���P�p����2�%gq�XA�Ю�*��A�;��#�P*X�̡�H%KMc��i|��'.<كA8�J8.Fy�j�[�>�FQ�����jm�\}
-Sm#�J֑T�
0�&��Ou��)Y�I:�s��{��Z�U�2����'��c����H>M�k9�h��wY[ ��Hct��z��@0}��Z�ޘʈ�^�g1��`mI����r�@�z�hӸ��Bp͟THo��v�4�߹[-%�`��$�6E�;�Sޛ.���;#���V�u��I��pHMGQ�!�=�y�.�k3�m[��͍�} u�6�xI��l�������Z(�c'߇��)��D���*����k�f�S�!4%y���������,���?+B�M���9���gL�I��l���W5��a��Rp�
�7>�]�9Vu�A���%$���VK��/������N����и �U��xSlWMB,6�e� :���hTW�C�j��R���fz����i����#���'���1�3f��bl�݁��r�����iT����>�>�|�?���~�K��q�lª�$�/�U��ȷ��O��Ǉ)9�&t����C�e_ �2�N��4���r%GYT� \cl��FP�V�Z���(���$���%�~�	�F�X���Q+�_b�y��mՔW1���m��B_:�r�*rS�g�-j:�hL�k�tn�W,�!���t�xEU:���1��Һ�K�N��+V<{�/�t�rt��!S��إ�h�}��K��;�S�����{0��!���Ӥ @�.�U�Y��LyʞN� ��dxW3D�4o�� Y�!��Y�$��	nS+�Np��C��zQ۔&�N�; O
c$�g�>&_q�M�ڋk�yo�Hn��>N~3[�9�X�XΠ�,�,'����%��g��K�0[y<8Ѫ��ľ�p�Y;SP�L.;���
�������!�A_��mZ�M<Xȶj���e����x&ư�)��8=��`w��E��'"^�{���~�c�x*L��5t�cZ�Z��Z���E�Z[R �;�k;t� yT9U�Xe� �e�:Ӎ ېbn��/�B�HZ�-!ϷړV>��	���!���#��g��pИ��dጼj�C09�Gc*���p��k�2[��Z���c��u�!^4�)�gl���O��lK+l
�K�Bu��Iv�k�ƴ�P��% Z�( b�����Nsڦ|�6
E�Ԕ,c{�s���:bf͂�]���jI�px�Ϩ��8�Q���enl�Py��AAl1�,���]�Ob�Y4v��`ʪ�x��;��xY�U}J*��&�	Sl���M�+���,�j:LG�ˍ��g�E��Yt�hu�r��rr	m*���"S>��]�ꁁ����}q���ח\l��N�v�I�so�^��h�B�1���t}�L�t��v���&t���I�e�g6ж``l�.8�/���K�w�b7�����Tm��}���<1����z��)z��F�rS���_<z�3�U����1��ZE�:=y�cCR��~��,�[c��O��*l�[](=��?��[�Y���jRL:�&�X��� �KIL-yT�!�E��DD]�+�\�:y�nٗ��@�pc�������wK����i�%�m�}P�咃)q�%������|��N�h?؃�k��5���[�=|�lHɕG����8�3ZY��,-�����=����%����yA�E:F	`���(㸰I�.�YC�D��,N���WXK3�9rkt�7��77��v����Fd��YC�) 	������.\�k`3�6vZ�|��ݟ@�D�tZo�[;C(�&�J��4�P2S&hF� Pg�I��X�'�z^�<"X��&�Z�
��\�r+A/?�,;��Rb�� ��;�=}��c� h��\�VJ��ӿ~��T'-��i�����8�ݼE̴5{Z�A�:
D�Ņ�(h��"���b:��Eu�S��l��<B���r~�9P��a�V��,��R)Ff���"��6_t���:Dו��:��I'�������
��h����+��U�=���H	������	�s0�9�D;�(�"{C�e�,�;������ȏ�.����Ϣ��SH����(���:U���t��z�@ڱ��4p��Njjw��$�����W9�7��ޕɃ����c��Hj�y��ᐧ��I�h5�H�~�#h�g�~(�������YV��2/�?���0��KG[v�r�x��V�S�������$��w�ѕal
�r�J�m�R���I/�_��V���v{ҘRM�Z��A����(<�9�璂�� �{h!�싥^��.�� C�͗��ei�h��E�R����0���-��u�L�b�o364�^��-6�����ЃV���	 5���Y� ��dL�" @�|�ظ�����R��|���P�ꤼ)�8���#�����|۬mp�A5҇/���Rz���&�C�#�S=�cɝn�1��_;*������RJ�4�+�(�H���Q�Z;����8�N���Xp=)�$ L����m� n *���'I6u�?b�����V�Ve퓳�7�q�&�8���O`R1��%���5M�'������W&�Po"�h1�܉|Z��
$�b³�l���	3%F�d��R@l��$��1+�Ԏ� �� �1�S��!h���ll���:b"������Kw M/=����n7Z1�=��ZF!j�Ğ�Y�=���h�H��JAqyT���AX��������F�s]�xϣX�.C03�Jix��ݖ�d��A��0/�T+�`P�u�^�<LyȄBL\��?I_Qb]*��$)���r��"��[�tW}H���|����[��Z�3G	�O(��0�b[C|8����>Ӧ����xϻ��-�܀��U�v���aTDf���}[� 1���+j�N�hN=��������[�*0��;I�A�	�=.i�C�$+�k"���H\Ŋ����BN����]�.�����9�� -ϠzY4a�d��C؉�L�\S�n�TsƐ�K���N. ��^�|�IE{u�l�Y�/N��������B�Pp*#ȚW�xi�Ǩ�i`?=&\u��=!ר��Eq��$��>�a�
'��Ѹ�ڡ�n�Cu<؊q�/�۱d����u���@6 a,�]7�à�j1���ӿDV�jFR�L��:�M68�e?���ǋ�,���)	���Y@ଈ�ޏ�_}�V��Y�z��v�7�����g͌�'�p���٭_4'�)�JYxY�9~���*�¹��^�p��&��[����#�h%z�&�$J���x��_�P�N�kԜEyoKm�������RVrkl�MN5�T��D�(��߬������׋^׬?.�b�Tx	H�_7���X
����A*o�E������&�И��6'}�����n�4)-.��O��2��3���0�걂�r�e�v�`C�y1'�fy�U����g��eݍ�z�/s܄�)���ݖ�gp����i�ˁV�<�b��;ҩm��e���-�Ս܈��t�����������l�H]���4���r�J9f����/ޱ85�PGM0nR'�R��N�x�hDH&����F�$9�T)��[�y��-��AZ��>ݠX�F*���4�L5�F<T9i�L��5�:�˵9*���(�~7�B�tC<�1�s��-��s��tTXi���;���56z����B��
�b������op�y���˼	 ��XC��ˤ5���́\g*����#�Jf��t|�̽�T�-To��i���j.C�/�q��R��H�˪���s$��Y��`F��\����Ҕ�����B����q.H��OR]p���>��_8J�F��i���u��o�]{���4�

~��'�����mG�*X@���S'���U*K�4XV�	�|���p�D2�PkMT�D��2B����O;ů�v!��;�ۇ�5Nz�h25�=w򻚄'A��N�9�>d�p*tʰ�>
ps?B-9����9 ��p4/U�$��,L���Z|8�Q�?ޞf�	�T'����q'���}��E��t���3�}f���wr�U`�W_��/Id�:�K0rD1�J�$=/Ǯ��·�j��kg�/�s�pvF<��X� �^n��,�~�%��G7&Wf������� g/�-_�WH�L�5گ�?�*�ȚLH[��¼/�ħ�'A��j�S
R�������\.P6b�����(� ;H ���r��$,6q�c��0�C�{�#Z����nif� �`���}��V�'�>A�@Ma��0������Hk0�L�����s�[u2e��W蟣��/P�m�]�8�9v',���N�|Y#4��;�3.�����2_���<�VBiGQ`����V�$��tF��+6u֏>���G���Z�����H��J�լ=\�4D���Ox�q��+��Vɜ��X��ס�e?��Zq��ϕ)�L�T ,�]�O�!��q:�܋u �\��WH��@��{ry�k8�Ahҹ�y�B���d@��j���E ���ddF�>WyR�9ƴ@�o��@�� �V�����d��^+��J"`��~�b� D�V���i���1�J�OY�d���`�qMy�������S$vwu)�2�n��o.�q>1U2��[̰��H�����Ʒ��v$}ޛ��p�&h���<�_G]|��;�1�[�A�r3�DE�p(��均���*�;W�E���\e�3� ����QG� I�J��kBC��{�h�`K\,��n�1�/�x��nl�^�3/6r��F-�0rk�V�&O��~1���nͮ����k�v�L�=��F�Z�{�" �HJ��P��������7)�E6Z=q�TRT�M����ê嗵s��9¯��%$�h�ѳ���9B_o��?�t��r/m��F+4��s����ZvL�ծkG��4
�R���xev f�ΰ���D;n�!��{�^�6H�m�����D�&��_E�5���Y�\ EB�*3j�X��V���e�T��i�E.Z���MS!Z�,�u�gj�K�I��m[����D'�3���<̨.a��l�Q��@R��0�r$�Ú�,8�Oni�oE�?IH[��g"-��CU�՞b1Y����m�^	L��3,�ʆ)�D�`�Kc^-5#pZ
=��c�c�я���AE����Q�@9$���#�Z,�`I]cm;�.'�����7�m���ZA�J
dt�Ͳ#Mry���}��~��eK.���4����7O��(f�Q��/"���%j=����4o>����U8C	��c�y�YΔ�� R�S�uG��1�ޅM�쭡->�S6xe�(z�=���Ȭ�	�vK�:lӄ���D�����	����[9A�Y�v_"Z(y��A�e�<I����x�s'��b��	����KT��,�ҹ͞���s�Z[gl��2�;�����G�n^��"�X#Lc��0�Zb�ˠ%��=ׇ\�Hm��\i�f�J�d�ӳ3��Y=�x��I^!6Tn��2����b�o�b9GG�GY��hO��������R�ÌZ1��_�Hqש�20��2j��_��s��A�|�71p��
�aˁ������/}Ҹ��T��@�Zaz��;��$�e��C]��$q�}U�g��ZZC��f-� ���	��LV�Z�<{RdR%��z��3N[�IrZ����q�|8eS��m����%�հvT�ܿ�e�ކv��M�A��������M��@kg���D �Lv��پV����g��%�1t�f�^�d�&�آ�E����t�*%�Nl�4П��+�_�䠱������7�@���!���8�,�\zO��+�Ky9����Q�<�����y�ǯ�4����]e�2����J���<ĆNtޓ\%fĕ,�*��C�	U��HVc�4��}�%c@^�Q�T:���Hl�=JG��gcp)�%��Nkh,��a�'Y+�;��:`�7"�<Ok�D��W��bkr�zJ���*�I�V�PŃ�I)�Z
�S�y��l��c�j��'�:���;"�8��5�O&�Q�	���	�� R}��cJ�e�y������1ϟ_�f��I���h}�C��ü��O�i&���lI��!���棊.� >�Åi|K�ʸ�_=<������2liخC$D���˘���k��5wX��)@*V����	7)ˣ��u�v�l�ָ&��)7�LA�*����u ��gzw��gZO:Ƅe
t�e��l�(M�,w��]a�L�S�fr[�~䱄\ؤ�Tm 	��:ܳ���8S����9��8Ҩ��p���O_	C��03�d ��LTU?E�7a.�+��A{|��M�_���E�F�ޮ�9f��)S�ߜ� �����)��gb���C�/���sG$�=�it��F�B���-����eY�}ˏ�		N�z4�r�+�m����ײ������p2)Q�p�0���6����s��Wcy�`��'K�5�\���m��$��ֱ�ц��ӏ������w���i�c��Gf�:�����.�7"�#W?�n�p�цD�vb�)]Oi֡{ӷ\9ūx���(���N���s��1P��Y[��T�"u����ҞU�A�U!��M�: ���5y��(����������u�W��K�(Er4��ցH1�n~��Mo�an5��"n��t����V~4�#�yD!V2+�9����E�0i�?��`a�Yq˖S1�/����:����N�oP�@Gy�Q������r�� zF�o���.C3���v��'w?�r�iD��ZM�n�O�쥭���	�`Z�h�i�����3?�j������bU�"L;T��4�T`���{������<5�SbS��a�pR梃�꾠��$���?�◂hn��328�4/)��1̎�c�X�E� �Y}0-�n���>8rJ�3��Jn���$B��1-�FJ]v}����� 7<�d�d��%�r�x�
�TzKq2����8?��B��� �1=�pN���UG�h�Z��m2�7�S����;��t]%�Tĩ|���¹������!�jb�V6�o��{�����%7� �y�9�ėlÎ�(�bp��L��c��HMP���M�l^��������"� ������\�\���!�TLdwE�#|�_��Zѩ�������3m-�N�U��tV^9Aa�8L�ٰ�$]�&~��r�������_�{����z��q	�J��}8}�y� ���f!�o+��B�QG�7�sl�ށJK���s.��Kd��+i;P{$��~WA��R���Sc �Ƽ�=Fs_��� s��,;x_��y�z��;�s
��:�yS6eBa����6�f=;��j�����	C`�q���'=,M����Ѵ%�����;v�V��{P䙔?�G�-?�u>�,���eѬd��46�7Ƭ�LY|����͟M�h�y�Q����ǀ4	�$�Cu0r:���.��kX2+sX"�]��|�>D�4y6Kl<}V\^i���"*��Oqj��Z��3��B���]���RR�N@ve�dY &%V��F+zm�,<�r0��phG,=�
�ȃU{��L�[�c7S"�)�>�C��s)#Eke���;x������A�R�-���,}\x�+���;!zB��C�c�kqÂ�1|榗�r�?�R��Ɨ�;�~7�i���z{K0o� ����i	�љ2�����t�{�.�`mj�H�8I��l@��-׆Ww����i�u�B 	ܵFþv�LVz��d�2a�y���YA�pSN�PѢN ����f��x���#�!�: �mZ�Fԙas��_�?���=_M�r^�v���i�p���l���R�,�N~ky�Z������^��]�!>�>��3?h3d�mM�h��u���� ��ΰ�K�c䐹�^S��GskXxϿ�5� � 1C�T'�%\����m"�~��;��i[��ҕ�,�����>���<�/�G��j���G��j�b�Z,�ِ0n#����.l�h�[�JeЍ�s{�`뛭����ǯ��瘶�s./ͭ�	CK�Rjv�Iu+�3�nc7=�:�`�aր2�~[u�!��[�x�(-�@���l��8E�Z�qٰ���L��li	��Ye1f:���gu�����+�]z�y;�u�NP2�m�Q,�g@+���2�L��M�
TL'˶G0��ME�$����F�Дtՙ�
F�bx��o����mH���S\�Kp��Ȗ�[F��A��{[�N�7@${��vF�x�d>�^��K��T��@��
K7*؍��7_�Vm����jdh⃺C��Ж;*� �ߍ�dzx9�T<����H��se���G��V��=)[J��,�$��Pø]yݛbJ�b�Yk�5^���V9����x*��<b����ז���\R�H�Tt�P�r�>n�ԉ�)�x�t�_��x��S�)�1��"���]v�
e������޼���z>e&�I���u86�)|���%�!���tXw�+11XC��;�0�����,%l��56 �)y�n�Y�'d6�-�9���	kj�z���m�x.�|6|���(Ri�k*��(���xBs{i��{�Ƿ��a�vu+�w>]7��k��ͫ�@%Z�����4!:m��B��N�=2�l���R�75,�����PՋ͚�$���)��/p���E����g���x��
���~�m���c�z�B9��n�=�gY6
���PIkZR�5s�f�+-���}E�6���мZ
���S�e
��lt���,~�ܬ�e�o��<͠�jTsz��.�F0{��a����&���_#�X���׵K�܍��n\Zqp��rڀ�G7(g�A�R:J AzQI�M?�c����-k6��ȯǢ7�e[�x=7����w7	��~KW�^u
�U�cy���n�?���
^�����@��N��Wzb�X���]�W
ͥ SB��D����c�UT .��M�E���áXP��"�$�Rz�ƌ6���l��ٳ���b�/!�^�
���$O�t�����VH�br�4�Ui�w$D|�1U��c,��%�2��97ݠ���M����y�y9b�s��N�g�WBC�Q��u���#���f���,��QZ	�!�s'�q~�B��0l��AN�1�sY�+YX�k���>�t�Y��^Y�ϒ��o�@g}�3�[A�}��Ќ�Pn��k�P��Ăe����N�R3]����/�@@4����uZ!6/dD���Y�7RL�Z�h�ɭp�����~_`��O'����xR;E���քԆ̸;Q�=��_/� 3v!��̵a��y9�0��a ���.�t�Ϡ��EU)���X��B�b2Y����Ձ�\�Y�q�{�e��b���a`�@���I����"C���p_��N����:Yk��d���a��6T̑�2P�
z�Ty�m�� ������h�QD�:_]����P}����5DI>t^-�AS�U�0@lB/(�
�$��3�gIއk�ۻ�#�c�����[��! �E~{mS��5�O��5�D���V���v�G`��-��7�T{3pje>��YZ�x�f!�SQĺ�ϭP ��Q%=�Yr�C�MW�'Ɔ*[�|"I�x
4L��L ��%�w��.�k��h�&�ėh����os���)Aw�K8<6U�uǣU��aʔ��"�"E�{��\��Q�m����#Į ��9�=�������SZ�j�nj�J~�M?	|dۇ����a�W��8?��j��A��r>��@k[��B@t���vA�vB0� �)�b&�Jҭ|��x�kF,밼e��X_za	2Gx����ɔ'�k��v�-/�uP��/�Iy%РY|��Rw�)���m'b|�w�����ᯇQ��w����ŇJ,!�`YК��f�h|2��g�.T���Wk���_)��B�����3[��܈x��z�i�_Л�n��U?�n��'��1����7�7v3��휭<�}�"h�L_g�+5��{Z ?�WH�Ο7!5�w[���3���O�V�S��R��ј��L��u���ީ$}�ҫ@���d�����.��>���t�Z�����	j����
���K�x8(H���T���0HMƿ��
���ZG���+��O..����:��S!��D`�!��-���K�"J����\j��;ov.����ŐJ+G��\��R8�#��ܸ�O�����( @�T9�^?�Z���r%�|�|��枻?"1og!���C8� �)����k]扈�L�V.z�4�ؘT����yۍ׀�C�jy)��&:|�n�@��T�׃�M�-g����>pFbFn�A.�,��� �:�75�
�G��:�б�g�1�'� ���+frf8�� � �1�ևӺt�%Oz<B�(S�cN#�G����8��]��P٬�{��j	��p5������u֦���':�=Ǜ�С�9�����	ӒN�g��1$q�������^wq��B�s�`����"y?�a�C?��#���Ag��*��].��r��3�#n@ ��W�Y�3��$�N�;{��T� E�I{Y�:�+zi���oK2L~�� �<��ߔC���1i��C"-=;7{6��$N��@�y�]l��f�����y=d%xҍ��ȁSz�=#r�C8*����T�Y�0���YM��?
V����D¼P�	�tE�@�"ī�����b���;-~���ʾ����&�lU\(����p�	&[ �y�ܳ~�ȱ�eG葨��_�gL��п2l����rY�7����M��ی4)��mAEA	'��Y ����U�������?�=y},iڗ'�5��ՠ^f�4��h,h�\(�"J����n7�t�4�n+�}��!��%.�q��7_�\AҎ�H�*�^7�1�&��-v��f�!����DZ&�&�(�)M��b�
i���%Ƭ�x*�D�B��L�)�X����WD&av��G�\����7X(��Vi���3]btbZ
J�xX��V蛩�g.n=�߫*~bc-�����2�������lf�#dr�tO�N��`�9h�����`���r)�O��f#�U�<�+��sf��Mb�*
 �xo5]�=k��=B�Ŵ�J�t�@{vj� it�}�
8�<Ш=���w�x=b�@n�_�Vĭv���3<��^�r�5g����/�k H"�"	��X�(/2��`m����2-Z��_����^�6�}��!7��D�|�|
�A�U6I�w]v_Y�H�Z�M���8 ��*��k:���i�q%p�Ť�V\VS�	쒸���*)��� ����X�X	w�Ud~����`ɻ�WW���+�����d��׊T�y�[�c�z��j���SB�΂�x�@9)
�kɰU:������������M,�t�$5�T��E���)�}���,qDy��6u9��m%d����1b�:��]��Wj��(�ʒ	�2��:w���u�9�G"���OmQ��V4Z����[�χG{�B�-�3�R�w��*v��
�|�
�(��fm��7+4����Js}J�B.]]�40�U�D�����oL@K���a�BAK D$��Y;��Û�8|��+��b͡9
a��w���nZo�d����kz�:�Mru9�n�ٚ�S6KaO�ҩ�Z�.�&�)����I�2�}[�/�%�G��nރ����ܥc�$�t�l{;�F#2Z���鉀W�X�Ћ32���K�~X�ާ�"%�x�siAN�P�c�z8vwƺܑ����u��7������/�t������:�m�ϧ��k�������b� e��a�r��B�p�Dii�̑�*Y���
U+�thI�Ն}�& U���G6��<Yj���=Sᣵ�R��-��L��f�,�n�u�-�`�X]h�����n�M����2:����!&�A�58vؽj ��@�	���!2��+o����N�f��䭆��s�P�����9�F�Qt7�Pb�/��D<��L�`�Д����<�%~+��L\�_#Fp��&r��K�V�?q�{�9�=
�bMR�J��{*�e�$���6����9��C˅4�x��6,��W��"��4pE�:�����7�Q6���t;D��l�݉�"԰����\xQ,��؏px��@���DF��V/S����LZ��-�4 +��������O+�O�g`�5g;�� ;�P�E]���Rr&ωR���������N�q+Y�S�
.zd��G���Q�R�VDѳ;;n8~o��6�.���Av�5���s"Gz�wpX.{ ʷ7�6�a�+B����$Wu��T�c�����V��ڼ���͒�O{b���M���;ݦґ��>�Z!��S�Ik��ۻ����YB�m��%M��^�̖=�+��,�^�G�~����x/���8+Wş5$\�^��$��k�|<��n]|%/��:Y��)���z��a�ӗ���X�Ӊ=0f��s����_�ht�`�Dȶ����j�B�G�mwˈ���C�aZ@�`g�A퓸&|R��"T�ͭGa`<A��腒 ץ,s�C*-
B��^�$�S��*�	**@c���N�DS}��4��r��L���+�Գ�G��,���w�L
`����O�C0�|���QkU��^"�q�92�
\	���g�H�#T��4ژ9�W�H��ci:����r�q401��|��)=�^tkj�M*��yq	�dy�V�t��P�y$z\|����D��0�n@���}�^�p)�9�>K�[����	�4���M4Q�yحP���/.��奯닁����x�d�*��vCyKU�Y'3����j�5D�XJ��{H�
*&0�wIո�yml+��y��ꥒ����"a�Ym+#�G_����:�m�4b˘��ʕ��-��M#��>��"`�������45֬^�n�
��,ui�و$������\YF���A�G�������T�jy=(�=�1�9��5�����jf,�Z@���l����Y�bb+ѽ{�\l��D+�\!�(E��۰��e�+S)D/�s��s���m��́i�9``�r�u��z6X���1��`�8P����׬2�|�d���;��Թ��cx&������4  ���K��X����6���Z��s6�Ln8��ti��[B[�J��Sj@4�� 5�g>���M���^�]�B�OG����}������O��b��_��r�M�9Æ�i��.d�^�m������
W�#�t�)�)Y� pƗ��}�w��E��)R��*�jϵo����8y���6G^�Gҹ�]��7�j�p���Gx�3��Mx_���!���1>nk�����(����W.� ����iό} �:��.���[�d��|�%����O^ ��)�XG='���F�mԲb��:����I��u��U�5�G���벯/��#�7zrG>S?L�'�a^�V�����M�-��K�D�Y�-��P�N �oH]��针�FІ��1W�kw7M�T.��`Ճ8Ƿ�]k���S���\��c��Z�3f�s�	,ٓ~ANu'�ķo�s1)�r�[ْP�jk �����[g�#�0т]�_2�]�$�H%If馠8�v*�!3LUD�?�����Pkr��~a�<������>�E�#sCV�U��)\߬aO�1����'�
\�]�솃2�{jx��@u-�|'��(k|$P���pAӝDH}�l��#��e���x���Ԫ��Z�*u����U�&�y
 ����Q��i�wd���4.�YΫE�.G�G����pn�y�� pty	�k�G#�/G�f�M�Qи�f���Tc�;i4� GH�L����G��Ñih�^�]�~md�~��fw��Q_j�/T�!5�$�z�B��[^��]A��կ��hY�Ф~��]���|�	� �O�m�ZO�|e���[8-(�7�������^�m$����d�8Q{\�7D5aUX@���\/�mg����7� a}���i��+�� �	��ӥ�w
'�f�B�D�e>�V�x���'�Cd	7�;I�˿%~���R��68�~ӷH�o@������;V��Mt��>���A���̪$����Q$~�M���[{֮�Z+����?}��⟭](��P�"l9���~?@~����d��\�Nz�@�`zx��v�,ؗi�85�&�٘��5�P�7��1�x`��p?߻��.إ�^_�� �yM�8r�����<㿹E��'�]��o�f0ܟQ0*���X�?e��7�hF��"�^B椳���Q�;���J م'z �W�� �Q�kJ��ғ/%cX�q+6�	�MӒ���n5�K��h�w��\te�$ZsZ޴�v�oy�JV$Ո��\k:� :�b�UR=��QiQl�%�G+�O����p��㎲�÷Pמv�#��+�y}�Ą��E�>��o�����H#� ��\��8%��ɂS��rJ��*3�*�ã�=��6?9?���ׁl��?�X�G!qz�/�"�A&�L�M����`�&�1��xMSt��*�ٸē. ҷ���������U1м ��EZ���	c �����B�����r^^��-����r	�T�31�Bb��$E1���GI���ZW��2�x\r\��\s����jC�B[���v.2��Y��x��Y%oI{�UF��/:����쥮im��F�,/*��?�3��z�%�ɻ\�������K9H\%=��n�Lb�B�g�MpF��RB��V�0Y���9���29Ѓ]�nD�ui$uv�O�JX�	�ʷ�&��j9�ܮF��A�V�
呵�PD�D30^����� �De�{��SÊJ��?V�d7G��z�lf���
�m�L��%Y�١P�Fn)#W�GN����?�+�Q2y�v�h�6C`R�>�A��Iw�DY�(�~�^��=�󦞀�Z71 ��H�)O/����Ib�� p��A{�Ú�#�!W	�(�!�5�g㵷�?�Z8RU��	�l����8�Q��C<�n����T�PV؂�%��/�[0Ŋ:��>~1�3����TF�`���y�_�xeI��Ɖ.,��_�qɲ>�%�=���!e�z���R��U�V�-�KN���?i W��>�� ��6:.ZZsJ8��ӎ���Ϟs��G4�Ԙ���A.d2����!_�����G;7K��j��0���#�~! �X+(c��K(}W�����\���X��1�
LH�Xg
�����(cP U;-,-�
���s�@Ъu��a��!��/3օ�}p�iʊ�i���48��D!��w�W��X��|��Nun���/�"���v.
����(}���#6~,�_� rg�4u�r�h�R0s����g�\b�f�mu`�Ѽ�l;d�4؁��-�uXD�'>�kJ�`�g;+�j ��ǌM��옗 �$Y� ����({��#���W0Ou\]�e%	ѝ�Ԃb��yÊm2U��4���բ��K��'�aj,��"2~����"�DdZ��X$b�nN��TI�_k�}�֏ɣ���z�ɚ�����B1��i�n�2�m��D��>[�^�9��q.A,b��*g��T�B��3�6�)ȉ���PzZ'�QQ��!m�u?�칊�%�&���ُ��d+=�zi5N�qG�R�H�5Es��O��:��M!v���wL��zd�G��X��ޔ7�%��}���Ӵ�^��!'��a�jX�.Ԏ$5��F���;�rԶL�����SL�MS��z��z�Z;Ǉң�'�J=���S ���}�P��ZԃageK,^~�-�pp�(t�͂<���[�Q,��������Iʓ��x�+�BF��4]�XO�]h8o���.G)m�.W2����\rO�yĔp8x������ ؽ-D$�:ru*5��k4v};/��qIx�[DK1��xV �t_�>	���±���"�@)��4�Ӥ��ZA.���#_TH
�5��9�PZ�w�-�HH[%[�{��Ś,?=\�~3����g��.MIE#
�n_,5��}y;��5��k��3�o���p����[��4G,�*,�C5Wz��~>P�Y+ox*
B�B
ٿ�c��a7�ch��>����@�q����PA�g�2*��_q)�N!�H�����&������j�����9��7�>dnvX�|��6�U6jp�c_.�j6�i���u�{��u$�k*�F��Fc<�&�au�c r����^�o�h�CȐ©.���mN�>���"*>�Y�Q��[�̃է�e���5��c;��E��X��mC!�k1{�u�-��c�I���ZMA,�G�vWhh���ǟ^^�h<;ڏ\����4;�ߦ��ȑ�;d`�	Y�K�pGc� ,]��kO�xq\�����C�~�A���~�g	�E�t�+�/łu�������h��`]��
� Ԫ1"���Lv�������vO�X(�S�(9��
�8Hh�@�ڼ�B�se�S�UR�5�5�6���L�Y�����OHJ9g���a�Si
SԳ�b�m�Z�������ܞ#Vi��7c��rĩ>��D�p�L�m�Yv�q��T�$���Ld䄁ӄ�f��h~�<y�uM6��2�A<L�R�Չx��\�bCyc�^�'�I0���.�
