-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ri8Vg1ZKtW5qMzH2HxAKb+BfOC0ecJ6Hk1ghJgzaXXDSp+wDfAhkxu5cbEEhZbxXCIa0FUE9noLk
kStMkIdpfyYW9joB/CiulOTBbNlqPK0n23mxIGaSXRSDzIx8klsm6Wr2pDhnNGfFrVwu03GsVW77
Ty9qMQ+qJM7LDV+ZwRA9tlxJ/MwgjLVxEmi/d219lEVpfZvXVHSJNbS2cx8Cj/iTtmgxtdVKGwGA
KMVC1Ks3Iej96pEFbL4O+oyFTXjsYGwRKtZdiCu9tSV3Jywoe0RWClFtJ4QZqdDU4afkliBonrfB
1y+oV8KMk9hrh2o1CePCuzwkOW1FwocE9KCiIQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 124960)
`protect data_block
Wg5Ouw8uV5MYQ6zWypfyF2oWjc/VtSuHhHJhnFHkfhBdSG8AAar2NrXs2QqYQq2A8rOZ7k1O9kyr
UxrjS5gOs3D5XE6+I/lb4mBkVkrJpLms2r69inH9IQrBTOUGFTbAbd1gwdjNdjrxTaVWI62yowv9
loMSsHu1IxB+72AjwPEP9zMfh7Jnco2CM/Rz9xGVwKbriIJv2BOqzkrfG0J1rHdWKtxnDeLZXZgK
2GpcSuCoCkVeZ2flAAeE4F1KUnxry2cFhoGhIchH+LQn1zxc5KdqL9jPR9DoZ7u2yperJsxkFik4
kezrfDAyDmJVgKcohclckgD66MWFiGD1dUamyGfAqZhXe9YOu0JEAKcgAZ/VTIX/BGK5wNh/y4mC
HGonXTT+MXG7nZ7V67M3ZlkmEJxR/yJ3O6rdQVBWEv29i4IrGVvbdfzCCwO90oQ+IzseW3Ld+/sF
TLeagPhoKmW3nmzpOj1yxens7kNjZu60hKDgROxBELUkOJAOoYcJqYkXzuybm6MMI6UIsMT6/nZK
FVGUbgQ3FFcO0BaNR3E3ZDZ7gVe0kLQULwQ9ZdnSdxXqjtfIGNJ1m1wwjYUPVZEJ3AW34MvH0l9E
3jGSLqcjj1hqFGwFdbQwp9zcYd75lxyzghRLMrdWhjLNZivroqEgQlb15dIHhcUX/qlmdU/D3Auh
4EFhMdAB7uiKcZ+5inJlj1VS6zOMBWY5M1RvN/CACVMIVZVTrpz11ZHPfBAI+QJJ0dk8AeasILIW
ZC/1Xlz6NZbgEk7rWb5K6TpODxgR+wMZCsQUrvxEpiFsrjZUWqIO/znGpZR+MubukFKGUZixgVN7
Uz0T73dPOCB3Fv5Lysr4FlAVwyH/dZshI34nmB9z83VKZPpIEEVJGTZO3TqJ4DDxt4wJwfKmTRtu
WtGGcNroSYLrLb1cJml+NsYjbmOZOwREMqJl4HZ8O65HafJOnDU0sw3jkcbmPfURbbgOz75EA2L3
qJ9YSZsUYwplznQ19bw+bLLvbJYPTTOQzESNsOmMXgsEPAJJYtW5Nu6uYjN6RLVjz3ku8GsrivpW
NZVRick+00MhSe6AXbK3Fpy0KDrWa0pIRv8Ag4CpEdSHCDiBCh9qEeGQRV0ny/2G/le4FlGpYfzo
k4qvH2MU7LbpN33N9IhY63So8MAxyGPLkvxgRdeOQSKaY4tw168AJl+Er3uePWTSxdAJ+BqVWFdg
N5glfCxOA5q+bUTFsWyUmT7lGLgFLpXcFT9ln3Pu6dUnSmZ375kZD3tYTconxx6++/UlCRjcABCX
Xqc78cRF4pISbWYMJXCUuD8hEU1W6eGiIJGXuaEhW28DmI5NFiAk2BN40RsG0S8XmOvryqkI1zp1
0g1u/6nSnCzLYeT9zTJfWjz2vq1GihotjlLl8dJQKhrphC9FYtdq7jkhpFYPzVu0RklpPp2ytLB/
l2EM5X1h5DGRJrsIcvmNaOKdsw7OoSr6ymvCOGfaAtPXAp8A3pgkCYAGENjqV0gLstD7QsGPtcxq
SpyH1OU6Mrc0CaFGxQw+Z8ZiaxWxRbFDimbW69WVFmeVCZ9zskceijRCfw4qZc3BwZmSbWfjJuCy
DsAzXVIiTtqZLY8yoviw9xIrKCklRMg6dqb0v398pL+fCBSQYTsUZbdtzuyWZ9FLZNrdyXUqE3+i
uyyCZVRl/ggToJDkyu2kf/3En8rl8Sw1/il82py9+TspKKCCTPxAmTSvy0s26oRssv2wk4n907Q6
Y/l4LqMIAW220L6PzWV2imG4pYU60xtQqxV7ZQwVM421PR3CF1Rfqhs2Z9KXa2rarcY5FHHpaRhE
tcfrY7FbrenYzKm37hIgE6cZNhXzp2VjINsvgLFzE2IwabXgpIsoQDQZgMI3zighCWCLEbidta3H
bnpGqYDV35JTuCJykuBQSU27jZpefSCmSx+AO3a1kJFDIkp0rC95uPwjDCQl4RkEc0Pw9vXAOCzf
l7d9Ej3dyHGXAKr/ReF4YkM2c51ywq+74ke1+ceyH1mOZSl8195EGbyVlRkBDMRfXacwio0cRhXm
pC6fD4cov875v0Ig9aXgJMLfd+ptgcu+ja3DtBDR2gD+RTXtoAY9Sr+q9fl1eX2auA7aruAvQ4uY
mciJSnjMZV1KCk06E3xeM5aEaDr475IdAV3aSmM37dZnaAgiVspaKe2uD0OZjpMu39/+Cv0NaHze
V3GApBzurMRUOmagL6/2kj3C6e+MjoZtfFMZ+XFDMy3llpodFN1HVrf1JBoJejI4ibrDMLREV2dR
fawM8Us7/IwQ0AW9pz4+viRud9YO7IH8n9Ncv6lD0hHOSwYrMygd2vT9TfNsSYkHgtpucZibt2Xi
8eQYZjcBQT5Fz4NQoPfqlA4TogzgzNdGeqZHvjsgCtWhYtCfbkUo2iTQo08klwtzZTsMm1pgd6L/
jbPNqm1rgEK4PCA+p9qfu3OFuuGWKA3Twc2ePQTtRmMNm0lFWbjGzUiD+32zdMKb9En1I3xmcR5Z
fDvwvGnhacl5CRcn5+QbByYwWtsBPDjgdt7cg39LKsqyT9aSe1hMd2mTt15gB8hbFi0oiEyyEAFB
GIXCN00sObMpH0i4qsOGZgDkANuxzeIq1Xrsjpayu7oNx8ZiOYYt4bUAadkNhNeNMP+OPiT+zt3H
HZVTvlE7sogeKBrZ/NafVVL0HCtykfQY6+dbOAJgGqlPdLl9moRiD8cE27kU2oIxfYoH383jU20D
usVLz5MJhl/y7JhsggTDQi8tjGmfReLjbEzHctLyRQHUNLGquk9MTrvBPeSDOBT883gs2zGOHtZN
velqr91KLUtUoosxwBmFoGUMRK07Wf4M0o5nKkHOesEK9Zdt4CTPWe9cboCgiaJGvSOD47cs4q69
PTews6SlOj+i+Dt+B2Ww7K08r8tipHxj3Ukw4qzuhmPy9j9OXaq2jj3LswRYOYMjImjTqWx+dbMN
8VrVH6KifvtggvLfHj/8QnH0dS3IofexEF+UN0XFK61/WacExMwwbqEl5eAx/IpBYBZ3yrJ58wBk
6IFCES5Q08qV/FvcDiDW1v+XJ+McfkfnTidgKW9/jgnGOfQAbP995tOHfxYdKLxtAnRPUbI23oWI
13rm+LdW5kMaO4pyqykMiwIcB8LlfPGGT0mtat+x5+qK22ptmBOPkJgSdoYTI0UQyUAQ1TZs2zel
xVUbD5P0FS1VOtoc4+UOLCrXvPYQO88jPUm+zQKVb5mPYj7+mE6LwiB1pMKGEwExcyjLe0RpQKSs
nlzFlYxxSz3Q3Wk/yBKHx1L6Dz+UIIuOlMMFPVN+sTR64IN4pfHY5FIy03EhYWYAR0cb56R3HSyw
UJwZuUDcdCYo/OITz79K8uEFZzyEJbRKNv7v/VTnf2tPMJkknzKwfeMCSkFgkdaApEC8mLTBXLpN
h+xNnv1xprm4RG9+DyUukt9j0yWjBdMlhEEZYdW0gJoO9A3NCsoMzTUYdAtcwwYxKQgsd7P1suRq
aaeWCcqD3NJ7yJvFUpYwhbHHp4OX5cYs69LbyTSfwQkoMGp7iOCj19Aq69mtPvXWJq4A/Zhic17E
5ttH1wukMa3IZJCyzmY1HZY9drxHas4sCJJ2EB3k2Ze/J+y7uorZoZ/5qligtV2jb2EU6Q+VqeOG
Ufuf6XEuQJVF/ZhRTONC8UzdYNmTeHHmfjD1Rlm9xtiLhYi1U7T5wncgtotPMIqT7IKSaWKxRbC4
VNah1rJEuimR6JV8py6Q6Y2w8mttV4HQGOtLcOWnk2nbX+x0VrDhO81mfxOQEPXLiwWOhJuNhykW
o4aA1pxzO4HMNrh7HdyDb7Egg7KTFs28+ZCj8I7NqBYgVk82sAfGh7BVoUbOyhKiB8dA+Q6ITtos
xB3W7w1nTNdL2XK4wNKy5u3SOTuIYqNpgBbTojsB2cOXxaqG+bk0k4YKgUVnKgnPnafEA02w3oP5
QDvofiHc8ZbLzBhxVE12ziFUiwm8ES4XPYp7DUsuSI5Uazoaq2Ezs4ohJDtp/78a8OexKoCpLpDO
w8RTe6rr6hbH6jf2aSQXKR/CqaGRd9jW3UFVSiXeWo3br96xqNyfkroS3u7aGpkGEzGPmLyUHNqX
NUNcsHYFaIBVR2wmGgsJp7+NtQSwPnasxJSWwxlG3EFBD1xt6cK8Rf9Apoi1sjjewGLx0dlRU1XR
JVorTG+23QNae1nC2D9MKW0Z5RL8nJQbv342F4vk3zukJAOuU1A5IRcMaUlSB6rbO7eeI6BaHhtm
L+SKE35NlGaSWSSnokB2/8nONG8sb6Xjt121WPKOh4aiMee/vcamFz887f+HQe1jqDtmkMVcu2pm
8AAlDvzsfpxVvmC5Edrgar2jVhow6b17XM6jB+fQO0FqmyfLcHVJXarcaDs1h/m2/8Jf26LrQViS
16/uKhwfAMVpl5a+/7giuSBzxlccBo9SzPzL3zVyEyuJ/S88TRkCj1Dpzv6r9Q2TMQm+CI0+XAi7
8DZ5w+HgVqwo3teBaoNNmkUNSdv9N3cfpOnrhKBkU3YzJ7sNZzIXqfFK10xOltsnkHzlUtseYJYZ
pg7fVsHGmFZ5brIaXv7ksYB8TlgQUosHtANdI4EFC1IyaDkHaMmZHvLgyins/HFFiz0Sn4HPahuM
IVXVJTSod1FligG1IwwwT54NkzIR0TfqzidtLqvUu0IO1rNvMYWLZKin6Gj4rWDtsQBFGAgMOxdG
TOIc3O5kXZHlinnxmOwXXZIHEbB71elQgn6lTinq227uVElxA00UQJwAbESp0bqXGMWaQFcUVNtj
DBX2/Hxu7m5kgH72ulUt6CiUjlPvKLatTDBS7IuOdmmYAYniAyA9VvIgoZlD+8goYYUpeLCfHWT6
ja8pmeNnhQImlYR4TTMky8bgWgjcPobfX4F1cU/3ccu22jFvindUxn7qQm2cnrhJmzdUls9JTJNk
uOrFLsmBBoZaLFRYo/j4UXgCVwgr4mivPEz3yr2IiHDcnhdJ221uMBmzH+dRW0LueZt2SduVW1ft
EdcNnJAEoWK3utmv/z83lZU8A5HVPDcc8Zm+vlaz+boguP5WZP7F6uGnlSrmDAqkgC97nOVXUI6v
taevI3LCa8hbm7Cgr57QvngI2ztwuAE4oleYnPvHhseClBc0Z0wNgD0pUFhsOrVV+ewSp/SuZibU
cpP7zrRUIjey1QjRdeXcdmhkHDr2yzAKk5mx4zpie9lvDNC49xgnwCh7hXBxyS1ZwWiD4RgnO3SB
wDF8bCKNtislwn/Pjq4JGuullUu0xovUz51qXFsVZzZgkvFkQ4Tm7RJFxlgljthRpnn4jvQqKqLL
2Yf2+4/K5X78+p71Q7Dyz5MCwPxzKSdy0gsUbv9V1cVqag+/vWOjPWfk/aBC9FyIGYmnwEah+YPB
gJvIXQKs/+8IR3QD9dO6tku4l2E+ZJ5a9s/0/lmaN9Tp7q08sBQfTWwfzmfB/oQ8fqXk1LkINMnb
Gu3J5esv5JEcxHxcCRrKe0/PF2tCeSuuGTql9l8QR8TjNfncsAka/49ESp/LRcG+gndKihOX1P6H
tMVIkiZxE1hp3qlZu6NJ1GloEf5YtkqXKeMastJkMM3ThLeuY3vQ64lXQrC5hw6ZDH/zAhjrZmEF
h5bloDZEcIeA8R2eYFBEJGbcd7ZSR018Rm5PZ0ofWbabiXAx9dT5gY3T0LcbxFrLE3Pljkreq7+y
lhUyqQ7HkfIvxOK0W0r/WR72JhxqLkooW2YVV8qqQVDMCi7rkO73pSt3jkWSGc5pzLaVFwbp/a/1
x6STcemJmGpjP39o74dylgzEnxYmLjesmwTroNEr0wj5Z2RcWkDKoaQ/UioIwLddewE/+T2VxKDb
RwcDiQzdZyGGkXJYTtxjVKhiQudfDnM0pGl7I7Okov480/yRlwHdMKVssENshd/3eBvGvJ9g/SYz
9IFxZRGBSaBuHt9Pyc9ZzwhRXDW21DZSnH8I5TCBJKkdZlWIcBh5wPe0hmr1lisDoMym/z6gQF7q
w8cVIiBPBw1pAKG1ESH9KKI4y4D1no9fi4R04SD4pa5OAmdq2UOacxP2VILzsWDkXOctmxMwFu8j
rwnYKW/3XNaH7gr0JW8Lk8kvDSjBMI8qfaRzC3EKK21MF307Cx8PhKaT54+fyqopkqBj5mpOKG+d
xIJZGKc2BpY4dP13A/sru7izpX+XeaThOiMN++69PVYdVFwYxycFpReisapncEO+lGxmr2Nriu8b
lW6pnfSbH1H2fdkHTlXbnf9fdWQ+5vPaZ+NdcxmUnGHKqN5D14w9n0iUPI8TcOCBvcGy1dDxUJSu
0mJPRDtxAkZp1jGuTOzzFEm7apK8wD9i8lE41eQsDRyQ6orqS4t2MxgH6JYv2iwOBY1Fp5zEYUXf
CP7/LEoLUeHVFmIragXsZSVImkAkBSm9Rs4vvexXIk6urL0va5ogMTXd5mAZHJjwGLyYpTWV5mUU
QD3+LyJtSJGmEDel9UTc7dcpCtAwJ9GcdsIW/UWHbCTG3k5p/OacoWvbMC6aIiHchYon+E/BQSEy
5NFaDzowbXsQ+cyJdi8G1DbnVTq3Izh2cm3fCpPuwb8C8DfjUQJP3mxHNuDW/qeeQ1t1R2Vingtj
Iv8NOX+uGFn4/COUVX8v+ZNFngSgw2fFR5BCN2wHBUPEJDG/Pzg5HJ219v2HRiasupNDmrLE7wP8
XnizYsDp+ROufY7d3TXQJXT4xyys0zv/6vk+hVchOkau5INnp7UHZmKr/5waYnhX7Ak4siDJZ9vU
dnZnetqpOUlCToUyuV0ksO0X1MP7dM3u3hcvNPcWv4QX8h4lXZfyDgt6EqgTk+JFbtRD6JnI1Ft5
y+8PTRABw7+hGx6Vr2jk0XUx5WgfIULCpKYWke29m2BtMJWhXlwHesF5GdTUkA8E5A/pPEH9ASzV
Vh3yvAVr61RRRmF0Nq3HaSCG6i1jLKeDBMPxxZ8HwLH8rr7DdWn0xtuV1SDvQiLuJL9eV8/iFU2a
xA1ZmMMftYSu1Pm5POQq99DDqapIsrdSCokKjFagg/5Zq0M5qImyLhBJ+oVIgO/BAPGGomgHWSZm
KmW+nlOPXM7yZ/GFqXYCQYUiR+EDP/MTAoydfV5mAUPBaOf67WZoTTEyzrvNCS43cD72uv9kYnyE
U2YxtBHavy98O+x2nF9VEkTkGunEnQ37JMIq1Zcd2Gm18/zQhyB9RjBS7KfQzEl7HPSHG8PAgf4h
SwuYo0kioXxDLE2TuuTZHqhD4SR///TSi7E2bTETusYSJmB4ofCZn9+mpSDexPtUMVznclyUWNAi
TOU/wktvz/5VRlTNEQqmfJ/BGMF+hIhF5XBi5pPgYsHSPDXDnCoXCt34Wph6ceDSPIeo6IzORVKl
cQhoKsixYvvr09ZhIP66OYHg7vzGJDJ+AwyWEhSnU/WQkKPuh0Tk4bEb/VT544rOxObifON8n86+
5+p8lVcnxV3LWImIXShuKD5KP0AcddVvR8zPLqAIesjJ2Pl4lYudVFORB0tEffoDSjNo/DAgJdxg
8yq01gMNycbWAuVS3MSt29IyfYd/ZAQwFMTF0ub/GeS9FQ/MKe9rFLekWA7OFs3M8Vs9+etg+vGj
jd0rmFAkBTFKpNegcEwgLFZBwvZ+XRyeYZfrw4D883a8u9WIt4mm2h878cHAV616w+CAU57DHI++
1AwK0mwP7RxeBFAkiSB9vFnCulx699LULuf3XMTxjBUbFgP+ph8eDyWd069uyB7Z8T6c9CPgmxtK
BW2JVaxDkR8QByLUHdRQ9FqYVki+pQ0WZK7mpIQKImFVmaSwgdOpeogyEP1XmLUh7bysaXREPY8Y
DlU0eNs6oHPn5YkFNg1OqQBLhkTHMCYdaIrjCWq4X5yVoarWoKpZALQT+XihD+O+qtYz+IPx3Xjp
FrgYgnDxNPIynfk98REuYZLXYy2GXY3KxnC941jWEUyEWrtvLaclPPMvyF0oBMc9H20hxs1nSh9k
NJYTCFwil+OXtC84mtsycQjfGGXN0j14PH+2+0n3su7FGiB46+Lh6Kkpo/qQH4qOh+l3ObS0jjf4
r34lzWDdNpimNTecXb+htOZiFnDjLl4ZE2mlMD1Ck9f7YxvPs9qVGfN1+Nln3frgbIW6sHHdZaQ3
MvJpqZ95shKxWIC8dXfPDsXu3JPlc4OOsSi1mIOODHCFJs6/+dxcuFR3RfD3+EX0VjaL2F81YZ/O
4oJOX6yGEJn0p4eWgyrmuQOBzD0dL0OiEDa4xAAhqlVQIRvWTENrTPfYtkjdvRg9HfTcRZ2d51cv
WWkqaH8rfJnyOxnDRi6B5pZhVKjbcaXiG0SejeZ+tL7kLNwk/1Cmm9+Em0uL2y9mZ3sPxdCO1gFE
jZjyiLGGq36gC9D2/uBmwkN3kyANKpf6Z1XugxNYpDrwiPGCJfiPGjXCmYfHV7Nk0yxtskbNH9NZ
2W9lqzxMNt+MeAbZuQ+UEPc581aZnGjDNORb28S5pnkVrR7ufcdxa0C7aVy6cfSDnSrJDTanxycM
gB6yWsoSpYi4N3UklbtDh4rnzE5PyIwecK/o0+QmLdM5btm+3Hs4QyfdIVJQjjcQZ68j/B6VxDQu
TTCMhuXSWdF26kIEUQddENJft/aCL62SyIQz6yzVeHnZ+9nhsVmbRQAsqlZA072NIfC78FLcwBRb
vZSTAxnnBirVDpqM8z2r/aCx/phHP9v3kj0Dearx1qMXIdfXOrdWrVzDFesPmSVwF5wjq/uo5+ER
qWFOgNNII1jytCRYj5CtxtkGcFzUuPtjJ93RLF+DPaYq6Ds9gp1NYEPphFyAURllbyAzba0+IkAt
4VZw7bk4FROWgqKKK5r5DmDNNZavhOpKImZ812/8E9GwaUexXT2eNOmNmREUIdvls6c03wOyfQEG
362rmpjrbyPY6tDusMEKCvvo7+EiZFeNzYdSqtmUDxu4D5SbYTaVSkwyRyP3N2I0NBPhNl1rhn4P
gyqHS0RgiCx6D5oSewtq4vkPRIIec3XLmSgGh9sOLdx5PgqNNGnxr5EEMvh+xbcHDqz8zimL2lPO
okdtxNHwhiBgZfI7r2QQTU0Cr0vfQNkoWprA/E9u6e464t+nwJgM7ixtFg1pqjpNFIAI9owwpxNZ
70PQSq4BfJYSgdhduyLyEbe6qHDCEXQAhckIroFXP89Vh37ThU9uwaJvYXNrlXNgWia1aUo8DWq1
wfx3bzG/PRMQEKnRH06ahVR/9edaTb5FMriFMYfCXh90YE5aoXOrJJ5WsUbNhlg3g+L8FUlQO4SM
x9xoHUZoXGZnBpCvQzRUvSAUMXFVmskKOIRuqw0tUScOMaowmuD2J3BOOgbWv9zGgdW8LpQFDxoW
Iu/0P5uY7zYhUG2e94YiVBwuD7OSFstgqrPSUwTI4TjODkIgfvvjxkcnRfNLKU2N2mubbbJWhnKT
dokYS1slL7Rz7PrKWp6+tSO5B3pjanL6NsJYp9qcosJTMt0MJssbTMMykY9Yt+PxHJBSIClkijMd
wWZjHA7lwvxKHl9W43s/01nyE4m2b1P1LhzXs5iEBQt+oZ3HHYrwRqMd2NcsNIfnXSxmhPRH1m7v
zt3LkKbKOO1ekKEcMbbIJVzOquJAt7ret2bQvOSqGEwAl7ZoJADQUJxjo6xN8+bNsgm185p6t2o6
KaSfqdqWEysuVI2C6JiLJHvDOhjKWIcr0NVcNIpinIbtsF2jV3nOGmoPLcClCpLKP+MJJlHKI5u+
gbgSTzupTnQlRUuYDxupVy2HZ7n9MyM6+wz+uLaeM7fvoDLzgZvwv9TR83skbBzJtwLG3JHUYHin
mkOa9F6aBVxf8+qhVVEiyExf7afKILVb7Jgl2f/W3SPN9PK4qcqVZ1tiTuV5PyLbezmcdZhtvD+M
4r+j7xD85foo2amaO/7hrHROK0eycrxbwu6E8ZQj2Jht7fi4qKwASrfGPzJLMHZZJvkMFKKkYZu3
Tw3OqtsKWxY5GuR1GKGnAq1UcQXjLNeSk0voQ094ghMVrnpipPz0OkqWnRLnfrpa/ZFcSxW0V1+e
Lzq26sR53jH0iyhzhspsA8Y8DBto/3oWY3NX9CAWXsv2OgLxXm9M+kG6cvPLT2AsXiGkRnU/vMeq
/2bk6fRCYnqU2TeDgSWibkaW1Nqdqgf5T/oD6RCr+6CYNTcej+6XDL2HkUfdraVuD9S2Raqc0QTU
15gJl+OYNIkB5A6cCkB28baPb6nPlKaDT0FMlZ2BuTzfWcYtYDrgHeuiwhGvjR8Lc/rRnT4Jr7dw
ghhsivlx4alBU8UmdGDgTABw6NY7ggNIk+l6sD1XiGLTbGKf0IwFa6FWkJA61b6De1d3Mhx/NE7N
LKW+1tnysYyzTG6HpbaVqbKzWS6B5NCgDN28VjPQbiBcam2MCwxZHZF7ZaG62okEdg1e4TA+oxgT
l2RVR1ntRi2I1jLJJSOeSn/srUOzhBb+Fqb9m5iQgZjNBNk6ITOpAfkFTAeE44AhAiB+c+yrQDek
NZQxr5YyM35kys8PNcd5Tr1rz84WdkgZn0BciN7gqJHk40uYAfdtA/4ViWnk46cn71fTOm1kEJ1b
ljL7hh6pNx+7UT0D4xIH1nR8NShnlTcALk6jEV83AHKhEaKWLUIBN7/iK9MbsCzgwLPQ/2htbo40
JqvhMTbwxIxSpZ/LXTZ/Q7jMFFllXm2gyQrry1rue3yGAjwldcgp1dBT4fSDLgaDBBYB4BqpyJ+w
9a0ELsfOBpOfFLPlFm9ajnB3907sZk0/3iDrunHZ5d71Hr/GHXkoHVTZ8iAWguQ1plCXOBdPU4AP
AgpBKSZwjnv2yB5u9FV4OQcmKpIRcmZzRha1kHcsKfGz2uZgwbBmY9jaBiCDR2cLFjmVZLpTwpAS
+xo7SLtFGGTCiUUoV8Ef8E9FaFGg9h2+FoaHon5yVL/U+RAlsg0fQ3FKgTMC3zJb4yimrQm96BqN
8ZHiEzh/Yjiu3edm4P/E4JoK7Wu4lBI1Y00uwZLUAXUNqEkcW3BdiwgqfwPA/K/rMXSxZiHqJZx6
j52FphBVORik1IkiYPkRCtz8XtMmGF6O1Hd+hgT9ndJpOMHuNWpLZ+MrTplKsR6jh6qY8JYcX6i9
rVYhUreFEP7UDTCnDriHUe7s2nELPaTtGp0sNudrjpItSsF6KrcHujsN7cefriRedFd6vFl/hE7k
nj5lOS94FbgAtMwMXRAyJ8rpCufu2pN0r+QE2eKyAAquykxEhrT5ofBnYXcppZAK151viMzmR/MF
DE0uktrHTUL1igHLGhju4DzBRVH3omn8KJPlFzFwIiNIP0HZ+mltNW4rwPngxhkbMkdVmBAtAaRi
63fMrWzK26cLaav7as8vuFMBRZz47TXlvDMTMTdxMhd0cq98flDP5F6oFMABACBck2kmcTf2iq6B
qkjfE2MDgNdRSX2C9o3Ces2716hD1Z/qT4cK/1MTWnxN09yu9v0NyHbUPVHhYsMXMJB266twOwOX
wDXnX+EWeM1cgds0DA5dCTKgYYwrFhWrsrzFtsqpH1SBjcZVbZASRZi+2aD0fuVh5pqn00Ht+Gh+
pDgMe+mmBKSw4/IJSvxK7g42jn57O41ZNHdXGnyMZYH8tzWUy5H0MFP0yv0wwkkNbUroZpAWYkzJ
uMEdn0RlPIe5Xm+1hQds7U9/FjnM7NlGNgM7bm8plepkBZHyUJNMzCufYlfY95th/e2OJEL+UKYJ
E7unKrT7aTE/5/rK0UvZGZlQG/MjavJx2t/D3I1+cNURT5hO84RcRXXJBG2y6cFulgQNCT5mPrlj
ujrLT7AXxmvh745GKKAUxdtY3pPoI/KAM6Z4cQFRPk1UDJCtX/Zl7R70l2Shlzr0m6kKD+32AUu2
SPUK1jkVf81ztGHpRGJ6stp0scSXylajEOabtI1Lo08yGHLoj6D7qUZs23qme/WwQ9PI2KUA45UF
ZZfCtABdfydklvLs4OSdHoDaAyac4C6UZNEAyhQf76OE4RsCXqEeocDCUKCCZv0eKXd1V5HRHgsG
vUs1X9tC6VvDq2P/p2x2K13RAzaYmANJyoHXc78w1IOTqo7N4zVU1804RbVCqHjh59eQTEKYf04h
yO+po60TQfCzb+HMC99bJ45T1GKNfazvkc2/gQus81Ncqw3eC7hhmfGobeHSpMJbcChAm122JK83
nKTy+rvGwTA9EXYSIKLZcoN0dLcwEakhOEHlRCdfJGTb56SRXW+CO2lkcRWnIrRi8nKJHlMiDl33
pBu3zbfAsalaB7RmS/s7dHiB0ReWkS+Pk0QIPe+JUtDQIKFNN5BLXK0Goq7WMir6bvcEZRlmyYcq
IXgrar2YQTw/gTjpgXxrIeJA6PntZasfLaceHbZ22O5tSCjUIt6/h6bFHIeYPu51jPQBGwxkozdP
E2Bm4+daJ9NXAilDshi3xTqaCg044kphBDw2srewJTZJW5cDKvSlJFPSbC//0IOu302Gprt1/Vxf
q/XjpZwzQSoF7bUEqDkVhRZIcKcPXxjy8YMu7UrxGyxWI0vCLqbbRlE/YDQFvE/JIkVWXCVA4oG8
DbEpFNOnGVBLJVXnyGfYePgbF9celQC97wYp+II0kaj6qhCe86y9KOCoG50oEuXa2bMzZMTZopOi
/jpm43uMA3Cy/vCBWRFxaLu+j2ovsJvHD/wsaAe7GWi9Mt8+FfGqLhjtawaqC65qvzDmTfHkpBA9
wiVBDyTsohlD9HkeWdg29EkWihiG1K5ZIDhwdiBPbUTQVPJTDl8v0LDGobFimVnfYS5fAAAr8YUM
g254UNoWtZi3ZZCoWLU/MnD0tqj+X08Kc89sATYFvWzr+sobbZhstCBTX3fEgVn+R5dshx/pMrih
dsWvZ4HLPq4uogY7iGxqMrd99jXVkh0o+DSzgDMnFYQ57nt7Mc5G9brYXcsQ42cbyTtleHsHQl+G
h/HqcRcmccYTMbOmCLSyOkmkls6+63Ho87l4oSjwq2WtdzjHey/A0rm6vh3Rv/U+RK7ShrlXQwFm
15lN27/GJxD4XEcpHprvy6JYXgWt4NlfWawdcV0X7JpJcRvTQc/fBKScJN7ExUW10AmP0N9iNDv+
Ykfvsb3hxILfp8fsNSdHxegBmSq0vUKDn21hIOWne6Fm74he+1T4oD9CjC6vu+8CgtCdfizNj9lS
OuVVqTqkaCam4pJp0g2weHHYwVNSuhZMxrJWm1g0yyjTLkXtA1JsFSGlISdY5JUdts9DcYmEaEGd
fWCLmeuleFf//1mBzbxxmc2LboIOsvLC6TCVu+0VvV4knQWfhfJQD/IaFpc/7LFZR1+8s2B2YDAg
1QE7vxtz6DfNhzm6McuRAJGv2N7p7Uim6mJAgVS9UMJLod7/XtVYw5YZfdvKdxhuydiwv3cHzW5d
gI5Fs8Ngy8PdoiZGmOko0FlRkCubtsTwn4RgSn+BgFRJKqIERLuASIoorPOs/DrZVE6b/qMaxY2x
GhfBhndtQ5oGfvSpy17vKznxHuMGF90Oni7syIiUIlJwh+Tv+vomwvbEtNFF90QNRwBAwWLa2jqr
Q3K4XprlYaThJfcHJ55mVkRhdguZwe5HE/SXpKXQxSIzLbdY4T9UFESPJXqPyqnEScreHEHdU+1e
HQVpw7Bf+gNqOMAJvXh6El8uEGHbyGg4zoMxR/zNq84Czwt+gSU91kv3BmxJYZ8IaU6U4+vVUn3Q
AMhja/lIs67mvxmC4POSr6B2fDk44Q5wr/yzWfmDi75c0Q1KhIRVftISOI4T8vr5e0s0nIEKsFc1
jizKNzo/Fv/++W97LXFL1ETNmj1r1DZDuIfqM97BL5l77gyhzWziwB0qIBO8+AOEd8o0KGOpy3L4
xi3nqpGjwcG61Rl8va/IyHiOn23/uz5mrHzdiUnVIlBDCSUrUzfq5oyrTqAxpT4J0peoR0YcbRbE
83P8InhAQYFviB+sABiTPrq9FVkdPzp+cdzh7wbHjw80nlOkuleZ4KZJBHoEOjKBvrNWYp2OP41C
XNorzjM3/ee7a0nPV9AcBE4AWO1jLYSeMsIHq5oqxddQRfgcrBI94mk86l1U3GI7O1yrjzQrEhJM
UN4EQYeCcaxildCnYI9b4VIqIdiEv8kFCyAFLN0SRl1FepNyFL/7g3YnWN7i5rQE0d0suuIN0eWN
5haopKKnUhIjLWZ0bQ7vso/ANx2GYYQqMnjxDitlrm011EH/6FHheX1FXkclvDU3hs/82xwtjWtS
vKzKYAC33r6nYQZLAaMJowPqicu0rjjRYx9qd88GLsPKtdW8dh4ISPdnmt5DwNjptywXbMxggSkX
XhNhgeqD0b8GkeQMfeq+N1uPondBJ5ROJsGi/QNoT7tpowmuFndY4h+grN1AglO36jclyuhL9TQg
2mSFr151uTu6TeUIIKOYSgkG/mq79x/lmtphcGrUxPc0bA4ZZKVx0Pl+qxxdgCmxpAMRxg5q32FV
64G6SDZ399IF/DPbl9DFzfElSBbDxcm/Cp0uMYhEL94miXSm0DS9Y67zUcJzm3YZo14JmXK+zGlL
sj0kjw8SHGJ27W5BquS8zrvd4AKES3zHLrnmG88tCzM/dm6uGkBtC/twjSd+UdRcVJAQ1izXmtnl
lJ+wKaN9zCnD5x3rxxikv4I9m7x3zH6XDQzMFMdvD5wBLQpo1+sw/HcN8Jw6BM3mdGkp3V9E+Cl9
sRe5XH0xI1QdzTUZI14TwYBuuIGcTMHV8S+SAS9i4Ocax1UfAxMZhraSoV7gISw2RGEqjBPMWSK+
09aZMAqefwr3AqKbPRUcgLmnHpxJkrPDOjYhF3H0DEo9RxAQdufzgQlzvezPyHcQ1vPSa8Twgg6+
1zudRq3manXWVwkjab1E/4Spg/h0qHS9AHSxyBMPNzeo/SYEMeRDGlFjroBxGIbvMBgSuEnzGG0h
VosVpxuEAYsACslC0Kt+iJ4/HmFZKDojqK1QLm5FtlWxgwh7KNCIDk2AhitrTK7A24Cab6GOSbun
NF78psW+pEYsgnrdK7XHnY9+t4t/kCFUClwg4dfoVU7cpUUfLFTIKQDuYQq4CFl6v4ZwHlHhTKU5
Dea01aneFWb8nR0NrAtqX4wNHPL5kyhlPOvTHszdrMYZ30IzY4T1OR7MZhdqiyAenBbSDGnzb1UA
zraCkiUJ+MbC9WxHFnQB9l/W6XFOJgqypX8fnt6hXDtd98+anjkHBJTpOkUdfd8WBzj7awhSsSkL
DD6zbeUTm7c1ywRJlRFI9FVohnqYg5WKD7AiWkgjIJcsDlONK8dAbPKbPxMOJEhJaBxWzZKyhZ5I
1Y8/OgCOcSSGimcAzezGaug8mCwOosBE1hMiWwqpFmRiaOqO4ZyXAkKdG3B/kfVLUlZBwDJPSVUQ
H63KvN07ZhvJDIMyESe+Vt4FLIAC9+F5tATqtVpkDaord9c8yxXUxr6mzA6Pt6+cFXvXRf/gdD9c
3DZT+cMOm4UZpb+HbFhsrFnMv9+H0j53dNFdKrsKhYOuwbgNi2783Mcscye5DPLnFc4m7oKMDRfG
LWK1G5WTeaDBCz/LVhErYtvu1FzAX/UA6t2zyI5MwoYMVdv7a618Lc1hTUx0/cPIH2+Pdo+lwIrt
OKpsQ+WZzzdIsnZ4LUvAneO5Nva50RlYUHjMSOZGn2kY9MsRUSxwfFbalm2VCmDA22mv44Jr4LMM
3eKOwtmrheS4B0jjo5MOKxqeGh2g1KUcsUP1EWNpYFnQSEmDwa0QxT+5e3Tic0biKquHqrEyUk36
BmmUHvrOVLORSN0PPW0s8DoPNhd9qKQvan+6X87Gg7h1xBB10Ux4+UCv4p8h0T+TlRet5zYPWEu5
r9HmSrlqhDrOejPQbPNHs8P4oI5bzmvcA8qqA59gwO7W5KbLG3Ic0+FuN8idTnmgo761AzRfts9M
g1A9B8eVbYNzPhRbVAkzTDLd6cW8fP2EwvFObsrPF/OBdfcaF00ZR/5yp6CD8exqFkrhdxE027fT
WofOilI1Tixe2D2hoGCYsILGLp/7RCiTeZnnVBq66IFakG+o9zfJvhmZeVwz//ujaMK3rQHycxYw
VOt7EbmVILljt1lZed4CmiDoIgp8wMs7R7O0eqGb3r1TnZChwu52WFTrrIYCgYkaeJkTcO016OS7
cktdYYQRZGNzBIlQg/zmYmG/M4bGMambKssqYgiB3shN1BZt2F2ziJ63p6jqmhNy/G/rVDnLoGL7
mNk8df7F2NqPQHpRNUI3hSg/nVhYqrG44D6p1cO9TSBMLKsKvvraSo9S7+rkLA8HnDBuq1YGNVKc
drr80n1DKU4yCrCwKg2P3wKTv0Y0w0DtD1BPB7PGBLvbuKXZZdY/2VvIZs4xSoFXph8avWTAkFrE
LVXdQKO3Cx7XHSmvWnDHPEiP2InyFlhvG5cdgzmEDlTbfCDhpYbF6c64wKuLt8BZj/dJsp5vdXw+
puIWqeYe4p4No0L5LUAdXbu926FGhVnufoRI2UfG7BgQUNhyLf0R0xZW6TSVoWog6W8M0POM0WDS
DAV4z2cJbkwwQ3t3+szt4017xyBm6j4k5g202itQK9HMP0bm8+N6QDOe3J50ZvIAHXgasll+j6hj
ax4YR8PtDmIeJprtbJ4dvXzs5Yl3FcZuyG7gkNd4ByHRi8Ak/ZBgX9Idv386ihMnY7mApEEyzm+L
0AzI80aq4qoSTcTrp7GXDfXx+ALpaceWtHHjQXLu05UyT47Ik1WPXEBgtgkCI48MhRUW5l4WAYWk
NP3hX2dCyVnwKCBtNoLQ6sOQ2fJQ8y65TWYajTXeOHRboI9n/k5g+2pxiGca9XxEcCC/bWvAkqhU
ks2eXZKnDsfg2ziUQB30e0Rvbx0Xh9jn4EXceZUs9fuXED3Lft7XCAyO6tgGqUXWE6Hx0ovnKRo/
ll5dJ6G+RoDB2+TLklJDgPZglY4zcEpEt3sZMOH9iVKWVlrPazA8di8iRdWOa869aUZarEuHW6/s
JXWEJwwrbJjjXbsrNyEZCz8tMKRbygwvguE4uLDsAjB9D8kMnFszIbWcIEbtNFSaQSe9QmYz/1YU
FLYEeZp1Fa6HZcNjhbvuX7RVMw1HkepzuE9Ws31Era+YJwvDLPfVYQbCzLxHL9KwiAt5AlUYd6GY
S0z3gUfqbQWigsJN4bK/T7P8+r+jM7zlfZt1cpE99aRHulXYtwWeYYrUEyMee3HyyvoQcB4nqZiz
IeedchLVdszTWYr4hF+ukSIZ0ZFbaMbTJXVUyMIhZzNPRkdyAKRRSWS8H+zh+Sfyq/bkHV5PH6tx
OHLLlf1v6PhDVUkMnsb1qwveNNvYrHIUihTYDeMqjjXbLqaDGwAApK4xa8O3x1HyksaQ2RlhCt0n
0tAgqhWykawH/1DPfJFy9KbJMzn80rU20cj6Air7DFv7vtoXegyOpN/nXTRa+TGYRO193t4XG++K
DW0l7+LPv4WUEym6eL23vjCSPuvwbYMsvQRkdd6eXRP65np0+YydO7h125AteKIFogEC1oZz/5Ku
ZDqPRgROD8cpuhfuqa0OBt5PrHXUr2UdAeRSZm3whco5KcqitBN4pXmCHAxFq8c8KMsUMzl+6y+i
ZsYS/AH9ITchXmC/5DwQ0V5Fi7yxu2wPLTSHuFRR2vCClHCs4s2MKsh7lQuiQRRop/2gI71DoMKZ
BpvIaf3M2694pQHMb6nI0vA/MZ+Bithfey6AtpY13E7x53opr0pskID1qkJDmwUGdZyQ0yqL0yLm
R0pgO+/3H962KADDaBByGygwDx2fA1okTYVl+96iVYeYZNZAykWS3dFlBma6o76FGQZJVdtByxo8
B9pJnH6dtYEuz66O91vehOYDMTNpLL0oeyPlvfoQfaIVv5O9gGardo8xQJe7D9AOA0TYgMq2slXy
lpkFbwAa5V0XhwL7dr9Tck3TTD8542qKBzvyMjt1yeeNFSw8MVrX3b/1NlccPh0Ly6abFtriurKG
cyA1NpmiqaompIeaAlymC62ReU5e14DssBicxF0BUeM34fTMEh3b8WOMyJCnZFzkxbwNLRd06aN6
oGdGco6jRO/3z/IY1FPQkNsQuh53XSMVvx9uBHp9Xnxjc8ZWyEEVTjQgyP44djMZ9FHsp0VQiGvN
xSmKu9sP4GNSKGYLELBUPO9R7ffZxlAzNYZXXGVSfabkMIJ07bHPwJf7UrkM8+LfFq9SOLVeh3hz
VH9WJA9fgVUejiPi6Q+6/zUYg/HpjpY8D+2e6D0E9KnGNvk7oGU7ybTMHy6ROIwhRWPzDfRkp72C
x8oJlZsPXMiLWuEp231TBPA7iEYOqqxqMLY3dseWM4+d9wI5f4QEJwRy08YlQf3Y/g7NokPuM19M
ITP8zGeFoBtuO/LbTW9kbMwRiplWRXmbysQABgpBwbVe1PKdltJgsqhkr3LVUSfDgQ8Kp9Ij3nM2
ameW8qJQ7VrfHFEHddP9lVO/J8JOANfCyJQhzJwpVcuwO8nY/QUXcf2v3PKR8x0precnqhs6I0ol
WL1JWOvpkhsNPlbud6QynSmf33bZyrI7jT5W9nrDs4R6bCzhArVgDgYffqN1ACanz7lz2ouemV39
7JwHJj9RYSqX9NMUJIFN7eLsLAE+Z17JDS354CcJsemf2asvemTHQ/Id0dL4FVigJuXJN5WfU3mh
H03uh85K9GNbtWiMI/GJ8Uyp0iIpT/UKjnEpw9zciGWNA82nWoCtL+RYWYHpVIv+oLIW9NJUKwo5
tDpGA9UkZ4GX/HsXW+GaUFCZ3OPvj1ymUwhRJPjAo2RprkGoC+ATUYc6WmtUcT9pmxElDW9/fWSk
Gi0yOJhCyCnjFh1dm7x4quD9ZS1GPGNzoJ7xK7LBbfCEQP8DPolPaRtjmL3yHjw1fED7mLRhVnVY
kZz1GeurQiaGT2T2juBzeXtliDvqzl/DSsebvQd2Ae8QVnIszZcazS4qSFP8RK7UiB5QlMAUfosw
o+KZrB9J19gOeKHtjWY8zev6+bdfoIaf5Ae9f1d6RplqrKhbpxuZ0N0oNDOGvw7N0brz7u7WqO0w
3FWqlf1uEkngJfDnt0OI2+pl3sG9tJ4oLyXMgJJzXMNBGtdVN2cIPZylfDmvChtRlD5YtHgyaZCn
Bc7A4aznHsRRnSOH8cCS0UAoWwg8XRCyUgsTbMPgBvgaHpGwJu+e32GZ+aAAMAKilpaKP6P2ZE5T
lsr3dKKszbGbHIVMB+JkW3J8nc3UBRlOgvSX+HZQMIy86IYisroRRgRrMepQe9x4xw3whjkeZn5c
mSlCWhYaVOlMpLo9S3U9hAIM01/AYrMHLVZgEH51/ztP4C5SYvm+eEfZv01rLwJZr1+Rw7ENjESi
K+cClCtTW/+ll4+HEjfPG5/ZCZv45OD0YJlQeL3QT2XPri7Mo01YOvi9Fq4xxuBP2MPw60NksmaI
BOd9h3VyVNLb+NqGMauv19mHs82Vgvq/CicdqORNYHPMjGa3QnI82+x5dUOXqLPa1apq8zh2vrgf
7ZmQ7n4ko0FmtFomxfI5BtgPArZuDMfhoTviNtAFpQpIwWuQ3Wa08PDoQXlbzFsIR6GKyVcl39hC
w7FQsmgu1eZnTVvQQbmP3kQXik1wVJ+RCJOQJiRbfXq7tjcAwXCGglqchbcmfTKdOzHxZXovgQDE
unV6kJ2Kf86AA4nlHOOgKH+8raRE4Hq7nWXhQgluOeEEIz9lU3aZtgf9OEhhA9DG9sSi1ZtQfmKd
Aa3Nq5oyb3NH+8DjfTaMgriq8ftEdYmIPnuujSmh/Qd4G0zv7EWod2YTG06ypMX1WnS/Jpr/GQDs
hVhcCTyKOBWFn1rCOnW1mM5rZdE5lPK1LI2Q9bcae1PGBnqt59Hl8UaKa5w2mt4WLPbj41X8ilgk
jg2hIuhRI0IdZsN9GLxHm/UAJtULB7h4I/9EHxI62sgspO8Zi3W6f4alL2c2uQAJA8fq8++TqcST
hubv1t2dhuiULoz4j1VfdnVCRhfb/gatRvmhxwL3JT+sfcEuDLiBi8YNepbuO4A54Sa2eAF+npQg
vuNKyH1FnM7QhVHllaUpk6Q8PzPfTdZl7iFU++sWgvLo3QuAEvZHz+HnfcK09Jgh1V6i0H+0RGeP
HEoeyo3uXTw+pL1HPi54zj2xpGckt6ADsnariSzzL5E0P0tB6WEQUkr0r7QDBeaihopkFtK6Qnlb
+7SSqM9tx5wCLdLXFLLA20E3kxv14euCEPNS6tLapxxK0LKdvnyucRZl9dx4/wABH7t+CPlBz4lH
EK7MfK1Gi7K4vPW1jFR9qi3GFQmEwWbK9d/zCZt4XBNE3odsyQC4OHIKI6cFNV/IAlylb1h3wbtA
Udf2RBY7w/UkD3iVB/tR5YXdvx9Az2Ell4JxrRUR4rnR4CW2BB4fcOSqF+fwdu4xKpdXZ690By/q
9jVyUPPAyJRCH+v8yNYS5ohi2dASMJgMEkjmZU4HndtBF63qOaIKoZIeRVcSxPBW2EJf/5e2+GfZ
+9NGYGb6P4a3NkznkE/dreisHc4jQ3KD8U+yEG9EK+rfQErh4HNawgGLYeXqncZrSJ8ktcW0MDJz
so4tDy56tJSrTDpLzgNTRqn0QH0/MNgKK5zZBBt5VL0Wbn39Kvo3fcQwG4TePkZk8SOufCfY/uhh
hUQCHNa7unl6LFXjy0LO8N3/8jH8GC4UlfkOl+upy8qPm28axsjoAXzUq4SCOac1jTRt34ST9j2m
UUDl+VhG2Ei0+TEwhjMTu3aAZhYEHaXF787XNY/Wh/FQiq4Qj7NbiICXCNtwTkkbjcWwD5aLBl8D
c6HNeLwIBYDfsN3nHuK8DBWCK/8a9OE6eOgTSUKNoE5nUFzFGhYIvG6mBUHrmbkrKqQPXRWUOGn2
hRXqGZJemrt1j44Eu3LxoVDD+6z6FxqWkgz2RZviXlkq63yAd++J9+2mutE2i5nntQ6FfMfJWshl
Xf6f9kh0ruELMpzhggEnWdZrfjvUwDO30/RkqtlZdMrfTGd6O5vLKg6qlizhiIKqTxjBnCJgAiyF
HiY09cZm6Od7VJ1W5/mITq1amT0OCy8q+q4BixFJhGpN5N1qvJUujPQdg4z/rMNeF/9s92PX6OTs
MGLw0k88rYbIHFDzkcPM5++AW7WJG79EhmEez9tH+QVecwpS683qHNq6/HKooWfKCoCQboDcc1tO
JqtpcPVK1gc7WPBXp1zYpws//WBYdIRvEAofUgvwrrlsxMDB6CEaK42ehEr2XcVM7PIUmAWL+yJU
K9TC4nWN1iN+lTSuO/elkVvgCU5O7uu8YWaTTb2eV5wd7cSEP2DmMU6vfxzkTQNPN7tO+ws5WIlU
w8L5reT7LvRDZHEhNftNpTG+huGR0PVy8EyIAuheBC1HhWSYKvd7dCtBZmAuhI9h+LkG+4zslLIk
tzlc96e+i5xpmj9oz8V+mxcT790Oxca18VT+a7hIb3utzhyZd6TVUFK+/xurhrBVeGXilOEFk1sG
xgX5Eyt6yYb3B+sL/hlNXJEiKTTzHVa/ulUmzPd7U8J79+mK2SmuFBeWDSf7vedUoyv4/qLh0+8B
Fv4+nSU4rwoxmXYFx6iFI2TqUI3g6EUA2WFNHfP+ZKjt48Wov7EBSsuWJ46eQYSV6XaUgS8Zdyu3
gMaFjZPD9CISMMZfnzn7iZhLCiOPQYT9Nep375KJlG7f7ByKjXUn7TDciXObsGXtVCR8ftYOSPCQ
+oyseMcS9hkx8nC/me9y2l1uUs8dEr1HrAvB5De23++ZuZdBTDknR3aWhW8En6AbrOKpmhDx9Ebd
1VSjTotACS7L8wjDsHiv86e07sfMyzHasA4l8ZmbY3sV7kNAsGR0w7nUhfvampjxSO2IwEhIooaS
Y1FidqzjLdt70KK7m9QjRlS8k9svY8tJ7R5l6amLSrW9FtWl9H1FBcD9hHQIbcy58/pDjpZtZDIv
31MauGD/jI38/Hd7WxY7HPpVo1tQDPNPLLWDtU/k52vNuECJMo5GEUdUqn5PbDi/Mws7sgdOG1zj
+PeNDEqDIHrVLt1srJ8HENkwjuJbYNG2IysJ7WY8gxC+xhMnYybW87i14QX7SabRuFo2SD7xJ6kN
8UUjGYojPcaf5CE1QM4kPfw85m/N2JrH1ULeKj/fE99tflxuEfqwXfasIoGldHRDk23UClrBO2rX
dQiXz6LKZTOBFVRWKGHoffWeCbshdALK+JaAnlWJwCFAiCVwxQ4iIBkNq7G4s5yd1WCv2ktmT7Iz
gV7R0l9XIxtCFiI2/03n1W40p1gV6bHEyu9n2HdlKEOBAzZ4WQEgZZM8G2Q5j7Adpyjgie/rCBOk
szPoV2RdR3iovZBntaR7WlfPEbNFgpOY0Nvv2MyaYutEPnZZXZLMLhpXEUqpxJ1N62J1a94QUG06
SDADsC+OUBEKsP7g9osP0ac4kSP4sLc85LpfNEefEdue2fPTaT6zn6xzPELICHBhY0csFrDhXALX
rDLMscItuNgP5CHzWmLwpkk8mLl7TZvb2LRvjcqoLEqLviqs/Na6Qh6Ax2bqyP3Ts9wcZ+acQSSu
djnNtL2jKnLBRgoYiteNxL4dHwMC4txdkmlenX0I251Q5skLUooMf+A9cZTHL9tPLlMF5KJBBeaY
+FT/iN0qEE88TXtU/443uy5r8dG3oWbKLBva1SYyGrfMTralGf9tVWCM/bpbEqEhW91I1t6cRGx+
eLpxzU9HpR2AxmJMS83JWPYSV8BqBrzv0nuf80DrZBzqjwXeRRf+0QxD2N+FUgZBcZfkCb96mg2U
7e2TDhiztkP4sl6zTmOADetHHuEy2n+G9AfIPklEzXKyyhjBlSlKimrfDtNSDVWin2md0tB/5VLL
ZPEwUAk8ol0QUqs6VYVT8PgeKIppf7dVZku9bmbebBcoxm7jfeASZH5Uc+YQeTk0qC7GLKKHnTtn
JxTA0qNKhDNXl6/+A65YTWhlpB+QrZbKMxfoM0hWDHCr36AchkxKXlO8QHWBzZwbcTpVHpmnIYvP
T8Pj9wbbuFqmRZvNFWl5AIJ+ZxUxgj81aaKb/XsuXpxa3c7CdZNiEdGEQi0I+JzQ7uboct/zmlG+
fZWATeGXv5C2piFlPRADwoDyu29Gi5H1rfpQO8nzeaYMg02TgtFLQ6XF1txAvyuVyfpu5rMnF8yd
PdnxklSy/kq3uWT+gPknpW2j4kE5SmJa0R5ElH3XzSuUgVFLnGKX+bVbwEaC+Ob6EtBFWFc0ii69
OO/HBulX5WNuBBOwTjTVzeFBhH4RUzSg5lvbXQmAoM5kencPb1WXNIAHmcAI5bw3R21YscyBx+yq
b+QTSfCDSQTWDLsDuQAd2dPqwW/R+9BEpdoZmSh6ikXGeAATuMOeBbQeQI4i2x539xp5dcT2had6
KQ5sKcF8Vd9WuhCZ2aNGIzS+Y5WXPWTjpL4QH3oY3bHQbmOwWKSMDRyS+wTkk2lSBj/pEDM65yss
zvnwH/HiwyBsd3cW4uuebrhoPJspjHNw1PRtWBjJNyMRY6GXujT1UzDyPPWR7yNWqSIp93WAFuS0
/rET1VxjuZ/l9Xkb3+zoMfPFd/bnXdwjecZ3rEpKQq6uBKh3RADZ0eU1ycwa9jVodGfRmWeksFJb
xOtENJydvVIAvMqt9Vgh7lF/yC69kQt2wNfnI5dmooT31eMAQuLCFQQMdWDcrZ4rdInOUCCNHOHu
2UvUsrYxuimY9sdzsWDhRRNS7tInX6RYAD61qqNkIpd0oX6gKSkvhf6Mq+a9qFchqhSTgnaEavFy
ku+PatT9EPzSSCW1z6frkBH4TllaDH5cwNtQY2htM6E5kx0GfApaKu+3cH3stuk4B2xqISL+amm7
s3xqDpnAz8yhHjNz4Y9ZcvouFEco2W3swcmW471TwfdZzwzDZbWmiLyg1sBxg4EQHmZ5MPdAnr93
Z1HAnSTLzFbDZ37XKLLTDNzpn2c5/aSod5C0yRi15Oq5zV+mvpSO9K4e5k9PxoFTx0fzteNviH9r
CgyYqZ2w0Y0UNypI8AfHB+hocRmviqi9Ra1XsNQe7j+8FPpcsqr8IyVaMr7FpYnyVBOoFp/L5WCc
3bWiKoN/ElmAzoMCni6mxrlfGJ93nkfyWUp6BWQvIgFVi2P5GXBGyeyl0uJ6/QQvy/IaviovmiLN
IAdc+T2k7bfF2ZOrssQ8NAWmQCLD2XlQr9HNMVIP7U8L1jhAB8WwuVqZdzLR6ZqxaCUL3Jo6/4uV
RTeZJla/MJ97LtwrKzWcQTmHd3yk/j1altjdHUIuj3DL+7X+wVwa6YeL3SUBfvO8WIjCN7GEvMHy
F6VWCZiAGdNw3q02ZcUTB/qKZfPwcIEGCcAY2cDYK6QPFpT+hNQp7O5CJpMnOtA+cjwg4auiWBha
+KVEvju2gDS6MJ0VTe7C3Lz42FEoOHmZHUwjuAYuDJ8nhLRl+hDPqITqzqZ+OHtMmTbdtKcVtBzq
Rk7UbDWj92fd4JljD7oxkm0yvEmb3+9rAdsC2YfG7/LQ4G17PS3AFaxfjouANtPnnAHv/hNK5rDe
8st34YdyN8W+l9VGCDad9+fnZa/sEid+WY3eXYYhfgjs3tziV58mEqDnwZnoPn25ji3CqL0coIBD
fMCsHwn+UIm0yjekYZN8ZlBGDjA1eIXORq2lJ2ZwORXGDs1DgmSy6L5ctZccd9qMiH49MYLBfbYn
Y2IllPmj0nKXjynNAkO50wSn5Tja7CfGAh65rfnRLmcYHr8ILms24nyu91Yu5KUW6cBa6cNLL44M
KjPsjv4ExqTQPBp9TmKE1x7kQaX4mPtKWM7AqdUKtwRKPmvGhpvgfQ9OQcfyI43bs+idqD+pf7Sx
hK9ehA51lo49YgVqg9+D7y7h52TpA8wzVK8n0g60n/BlQQKJDnKNld9LKnbdt1yBQ4NIth+18V7o
2USapUvJzxvZSjrSo5xmgnqF/ISOEkaNpFA5OQDDH3XGB47LuJVK6NSgfDbaoDsKPnvbph+E1Ue6
oIKu/yYhuMyjRMbuZSnoQMfgv9N1TxXzJ03zMA80utDEGPHDVnG8Cy8BcA0uC6pShDlvowE0hQkh
L47qHny3anC4qUpUAD551DDGqMhqpooKCEmt0h7iPSvaIpmuiFL+V6/ErGV4km2YziHrUfJaLNnZ
O9spJwHMIL6Ueajwk472Vl0C/es0U7kBZhQEbrQhJL/u/uTuoGYFohQKxiIGMSyujnfVozSwYz8p
jAor+5sTajEdhzZEIsQs+5UJ1/iMZH/Y0MZagUhOjIAE3PnI7FLYjxb5+L4zC082c5T2RZbrU8cd
+eTNWZx+ZkIcxHeX90WRmLTZAipIsB3I6azZPcitbmAxYek26P/2wUuv640yE9zfLfIKDHrbiDW6
NYfp+HG78lB/oLNnPYIbgVnjZ+EbG5x+1VLF58vFjPUv/nrTjzjarqFs/SJzr9AiRsgi3weuvVGl
gyE0SyLMr5WPLcxFpit6+lSP6JVdz4BEjSfvVqfA4bgeuKJ2J20mALyzccNwdo5WQXeikl7K4CfH
onMR/SJ8cmHjvg42IoYMgqw73v2esMFih84Rwy+LXoF3RETR8XhClvMzJvrQvWClbyxawwax00pr
Dnen5uscXaBXLFtIPlIbRDrXNmfOZB4XgXUPhfFLg/dFXADqfSklJ+LvduqU/V0V7NnYsxFYy5rw
G1xa8PYpUwKCaA2qCEZ06UDrQKrhopkx9sNIJN3dirrAjAodTMwNIzFkTyQKPLWH8fGYwZXX7o1p
nHuSBBujQlQ2uVmjw5zPgOntYO3297bpADxW/i0tuy1VKVJYEazSUVkNEtqa8xfmo8WUP9eGwhkn
/5NHhinafGsU9MfpspBvrpnzWC+aLdxifbcgpeN8sqNOykKq8Vz2CWhJHFTerazWocXzoT4WCL26
QDUUW2EpYBz8VixsIV6oy7assTr82iKOmoAdfllb6ZhyiX9AExypGCSBfyDLs8gliRGJpCbUvAGr
NkJ9dkjZ59rORnPn/ASKmFJl+w0F73q+ZIaZnbd4LS28f9V7+AVGec1wtXFoZuLkCtkD/mnkDqdx
J3YBIm881UnH+Wstxc+Wr8K3pB+9H4pbZpXAFFOQu08iSANQ8jmOOQflZc9ohsyjYKBUU5InZbF5
vHgL0Ox1QDUGHn4h/5EHRQDI/bmnyAj0rPDqALXzKdO2nku+VN9677bDhJ+ktLn3RglGdwDpHSMP
AD+qGD3DsO+/7/peKSynoxQO4woo/ecX0fBa3vCrKoLXb5MoaJUYO0Y9DJRIxWeRUWLkxb5aWDBH
0SAO/sxP2jIzOGA6p3LO/6a6RvlsqjEUd3GN34xvQ+i8jd7Lkobvq/5LZE3kUOYMjwHIlufhA/w0
gmkpBXkLIBssHEtbvW4EfodjztHnx4F/eB1CcBSnHe/dq8upzh+92Wksr17hqPJlL7eNXo1CyuVd
4mxcMx10aWooy2d8LDJY7oXxCupW4gWTlaDXf4p/wDmmWE72VWyO95a6qT5hRo+at42L9nn1FyuY
CVVEKAAAfHUH/Y9PR4xXTf757ousjvrLK6wotg6rNBAckaKhyp6Cg8HGQStjsnGRuRNRJc1nLucr
NRJqonxhicc85mak8Kjwy+fNHqrnu/F7CrjlUutTIWpbbd6cBVU85dq/ih+qYiiM1VLoW+zm6ImK
+AhK4fFaL6Wd2cqB6SvcweNX5wWpKr2TnvcGt8KGuskWjzoAW2D62XwWfSpmOLQWMjAT4ddJFr8V
cg0Tfpfu8YPH2jypvX4Zmx89DY6Eb3WiNRgzTeV+aLMmE/IYpeezb9VPuU3gQJxJdgBUW6gydJRD
I+2cy/YI8SX47lya2SupG5GphetwPDrEzHlxZvvmukTbLIJ0NzryXlx9zuhtNqQ/lr2tZdf/Derw
MNqH9fRltyv+IX9+OBEwJpB3d5j50/4EZ9D0LruYwG7EKhs1CnQheTC996O4SlbcJ/QW8H61EPgx
jewHX3WX8GHyR7dF5OAfcs6GIDBMjYFLZ5Xc+o1uIpUF+mUVHUdTHR5aaqN6BAh25ATkT5rnczXP
ZXUC0YvMy3j9R5UUyXEogOhyIkedDlIyslMXvAOd/0ZbD846/8G8tlIZ61KA888hEupGPlC6SEr0
O+29w+esE5i++BUoAc15b/tuZgz9gYmVZMNBP833bZh46Ut2fjMAjbMa2lmGDcTeYCwTcoKpvXwR
Jtgd7cCGOXdZ7hpcifIolYCZmNcWSGayIyC9JBG3E+MjcVkBPAabtKKeqiUkw4qZg655tQYf/LYs
wTFkarFxlWiSqez0aB4nlp0C+Bb4Piy23ltXJAp4PX26O4inwpUHUXAk9j5at3UvLO+I+Zomd8xh
Ks9krzGfKhcd2jvSz9fvoO9XPZys9qWeNFxIzDM2MOZWZzqeK0TAK/tlVCY3QQMc9M+jnobzR3dn
YVaOez+aEw3iuWxWGrri32KQpi3SYRsdVVBKjsgQrtN5gWCOyArmLP+2m/yAJ6SVPfddxtCyVsZ4
K27YBwsITMnuEfkr2FETz702EBLJ1Ney0FO5NkK8P9hZvto4mHRYFLXhKTPzwXjHi6wXgi6zp9bs
Oo5nts9me+4k/D3anP4BXHShGc/GLT9MCzfNizI0LPtsr8Gk4bZB9pZ8F15fesZjKEQjG0L3jOfB
uLUAVxKB8MAGtEcuJwULdI1/6ZsITBYVmsvyTcDIWNlpCpmfZtaSI7QLvC71I/KUklWZBNKBPEZj
eM/XAvXuvqYInbTvJm0U76UodzNUff82H//QfhlsHuo0QwwJoYADOeDyAw44ssw57Hth3RdkuCpF
RcU7mayzBRTChmBBM5+oVzaSRawJS7e2wSI68sXAYJ4PP0fB/PpFnMntY7k7Xz5/5y145E3gV0Ii
jde2RVvYAF96QHR+0R06g/oTt041j8pJGE254kiE7sNblktN0Aa+88kfZQIWx3R/y8b2PZ+lCRjB
BG3QFKfVsDKzi4O/SJATZOn6Qf+2jhl1XD7VMGAkR5vR/lXEU18O+yWk6LhBFIKo6W5pcuJQOn2x
TLIw5woNUwvu8ZRzACa/txn0m26UprnlhFZbmAdyjUZ5vdLPLWIr/9t8pwLog1iIHa86zDscPcAZ
KoVOMw3WYpsGzJNGADDqr6Mb+L64t66vIx9kzIutgwc9NqAuuPJr1FcTGhJ+G7kggLwx4otXXc4G
RD+OK2M8Z9kg3tCkwlIyTDd3iS2C9KMsiBzxg16Rgjtop/tn2oQstyhkiHCbbW9GAwmKBRIdryuL
fQWT427OD4obzY3zwt9R3ELk6cTInmua4DI4+DGvyxihq08oZqQFdzIxvjWvAOifJyONCkqy+h1i
PwFTeIoX0v/cBHZHbNLM+u7/fWE3a2CCsHqstlSD0Uiv7lVAD/p2TKP2myFsN+m5FvSgsxgjyotQ
yliN8TMqgTU5Qju5TvRfvX5KuQD6d/5p+dyLtl2fUgGZdV1gJyYOI+vcO+tsoG9JfCOsO4RiZ/7+
SMJkrHXmQPO/JirZnlVOqNYZUgdbtb+gdBpJt4DDlF6hzejxukNsPOEFf9AarYc0tj1rD/D72x/X
AGghdVIktI6dwLada4cdVIKsPzIZR9uiCEAMhqaa87m0VkBO1pj/1EAy+5o2hrrLItSe6OiUg7Zj
S4LeK5IyBs/8t1uSED9GzzVszXfLDO0pGoWXgtDllv+X5VOx3se5W/oXu+WCG2Rlbu/KIbmPwLl1
gepe/QfvkNXpc7ceQFO96r4DD3rVFODIlWWgN0qszqmTiZ0HgSmxHgA1eO3aRATRGr5aCup4yRzT
1ZdzszbD39kccdHM+Fg3pic0d4mcLAjlY+OW/0YqgooGs4FYbrY7HmR0swsAwdLYqP3pjFHdwQjj
DerxiMbw7d06d2OU8TEXWircOYnAxvovaip03AIF9X75lEPF/LXR89e3L6hL1m0yFnX9yNaq7REh
hheVRKLXjOwydLyV6TDNImy/SSnOoe/kq4WQfAMyaEmxRDQoD2SyXt8JcoR18ShhBPh5UsfP1Duo
tHMcvMw1h9dkhI9OvZG1uOgJjeuxlXS1sgMqhzI2h4JMmXsecb5yBXkXxJGdbSbMxwuyEvfQpaPz
3ZISvHM8cjqwtKlD9XriOZveK6Jhx3UvAPfPZvf8dNGvfVn6bvUwal5GZgFmLsaeagYW86Dbh/ss
VDk6w/goV6hM29pVqeuwOY4A9cKBOFmckMkWQ2zh/F1TviXsgcyO9iCjyc3Tv4b3fQdpGtm0lqjB
J5OQy5mhEvIBjHBmT0AhHIPt7RG8UoVHrSuTC84Nihow0QJZmA8qp75EwpF5H19ZO6Kj/HRARf8A
aqur2s0wCWWOVo3sCxwpWZ9ktm6hTP7m4k3VVlZmmusOrYGU9fhjppQI5qaoXn5MNRuUIHv9uqRw
ncwoOfFKNYQ9q3cbDQ4COON6XOOutfYdRX+AROtA3CCLEnVzIuKntNBGE6FdQ2L2IQiAxPRs/b3J
aGxbZo8MqI7KwJIRezcr3C+0J/wnEeP90VGG1NqWTSntoYtczOYnqO/ULuTcsAHHXDaHEERihZtE
R8YstVHMEEyJJYbOWjOFm4rQXU2+oSoMCYvAmcGfSY7ozSSz4ZErTfKd/taVqwrGdicM0kNw4j3z
1W0PEO6a9AhpNddgRBfG6i+bGU6aNtDwJUXjwIUnztpnAL353D6FlkF5HSVPzmr43E4uInd+VSaX
/wPTNZYGs9uZCHvKtRk6LNbxWJ16El5M4oqI6jhZvfKBy5WmUwTvAKmO5uxP3vCRpgRJr3Z7/QD+
NWnN6KhqgBwcSP8nMECIlhhxXbwngqoMa+ot3N/kWg9llNaDpqAYz5Pn45zzf8x7MlQikub6196H
co/3kS3ZUg9qriLvQ79BCUkrYG8mnN1Jv3RXnauY/eofn3+RMs5ViSeJ2/U9B80UWQShwH0PVjFI
ksNfdWq3xmEEOStBR7SM4PcEOaXskArpVzQTjEGYCSvKiDoQ7MZ7L0rna735RmKVhOVjXCCM6hiZ
m0H2kRz2xeNHUtbvKooJKltPkkZCMZn+iATpq9ALVT4SabcWkWYhFHlWp0FHxaeG44CyN0IEVocL
TQsQ9GZbL+n++8fQk/HxcZJoYtQ3v+SfByd6V4Ren0szH3lg4+hNZfPnhPM69i3wHro6Pbcdz6Ye
Dk5ccLMy7I4metXhojuWCvxrCpQItYbo55YyF+Ksbf2nI71JN82V+LSHE7Iu769yw30+5e+pSVkd
1Qulup6T0oSCtl7dTxtYgzM5USGg/gVRHvuC9FtMNXMIMjDNXOFwIpR4BKKCwhaRZ3r0fc3g6xFg
73an2VFuqchmEhGLzpO0F3A+3b7jjyAugp3Q/KGXTVNzLBD/iu5oHtGF6T+UEHBHFXAFnWNDRayP
1zujWyV/pqSNMUuVmsDbrUjvNsN4ny6thTJrf9UzvU6LVCy9zBNkHomtgqZDWG2PhkY3gSTXiSbU
C27SaMLz8u4I2pL9CWCB0+BD5KOjqvnGBPnMBtDggAYOPpgHvPvcyFyS0R/2+l4kkK0qDIiONSMD
CHSPlFXbkSEpXC2fyS+hBIr0ha8oE/Kjz10J7eweStYBxbGILi6VxYpV6INGUhhWwhSpvSaAP1TD
17aQqiRjeTIMY7jGIc3YGt1ny1ltQy/CUAExDh7LRRmDHMMSxY0RwXZ+WgSOAXhItJD6WPyXv4FJ
Cg1mO4Su9BDpdNWjqvZSyKJ/0y3SfB47o4J8TNjuf12vM7dET29X9aGGtw2ZghS7EBfNAgnuw8rX
4GI+Q3I63FiqwDzSoyO4tzFir2rZdJlTBJZcrkT65bDJEsjN5Q5y77YnOnu9jIaiU3HTmzHM/Ulh
vy3aZ8qjd8wJfilrVUJJUdJ49l5Ilo+YKaahTF9bYbX0T7/vWHHbLBi7h6BbkrFRjHXj6AkNT/uF
xqJZK1bEkA8Z5gyqbr9oJW/7AlZy5yRwSGcKHEPAVGM16YNh3dq4qL4/r9NdChTF9UNMErXQXi1k
nBmKxLOK5FXBJBgTyOoHCAw9zA+JRk75fFVkEfWL32JKO8bwApa6WY1JsqM31G7tSkI+foy25tq2
a8oxqNKwlYRxQx6CPfvz3Irnm4Tl55h5DRT2B3lCo8P7yXwun9c6amZ/H2ylgDFSjm7pqXbANh3f
5/RO1dq2vnnNamkE6tvxrFRsopIRCroLzMdwKvVW+K2eo0PisUPXlyT7d/MAUAFedW8tsVRFC8rk
Z96+AanxbZR+Wi8GSdTHO/sTTzFVY/8iz0IQYZoHutaXxRTCD2dlXyUG36srxA/sJRtA64g5AZYv
EZi4qQt9OP1k7ErIb+ZmejLk3CVaMb5QuJ9psbnXezFgtxQI0PgH0igVjH+8O66Cg5TSnijBb72C
5bckxK+Ts4XzVUfD9/ZJcMzEFSiq6k3rlRIgWL+/BholK+ecA7aVACmdmrXlJBgiKyUfkEcPr856
uU6jLsGDD7jVbhFA6OuYq30xmhbTF+POASB58FLF0QBDm4EWerDc0GWpZvQyJpABNLw3tYrmvCIH
YZen7EkGUE3KRjjiKLGJJzQZHBQlviWiQKZVB4muxqER07PtpQxhQXOXx11iU2JRq14cNfXirwXC
1ydiImRaL1njS6GkzaZg9g8eEerHwcWNG4mQTlPHPLKOYJ08UcXVgBOgsHuHrqaED5tA0bXQVoxX
ynpv3z0ROEvXXm+MOdyqo5GRpqmyVni3Oeq0w47qT/2f0L6V+H329KY0QMrn4VmzIoN1gxbtUcXO
N4ZU7H0Ul5pc3pPTbhoiPZ0SrgWh++uNIU82Nn/FEGfThyXB+dmxRActmh0PDm/0B108PR1jpyIC
+qVrGbQWn5oWvRHQfNIAt03xTilot3/uz03OViFkaR5QvFFTfbAjAMu5XVZOyzODZllqh7Qy37mx
ky8EbDmuHuK7SAuOqZ/rnbTso/7ahzFjR/HcQ1YsyTPH5wRzzelDxaKL2vSFxb4t9e7UkV+J8o73
jpaArvrNH/Qo/Lqe4+/jCxttIh21J4j4cbnFih2oLoWhogfiGS8AwtFc7okPWnFwLeIQtSuUN7yF
pp3ne0S4LSnTLHb3fCRUy6qruYbDwSp3Sro8FombKbnsNEE7biKDT8hVtqV/Asjq9sMr1YWnyVr6
/jEeWKqDzGFQiePQu+zeuaBJNtwvXWkHfDCzrlVIy6m+J6niz7F/pCVKWqdzglSkCpzEZdqadGoJ
7MvZl7Ts2cDtADYX1WRjhqtg4DjP116+h2/9YqNLhATdQZ5HdPkeAUfCjrbe2OeEL1H7rzlW5BgW
SmNrVfl4Ug1y+vC8JwGXG+yohKl+FlYJdGQOR+QTfqyjUuudPWE+HogFGx2pdW4RqULphYupxLWc
iOegbylOYK3CDFtj0fUYn+ND0YpS1pNh/DlLoEEwCAYYtI/dVn9iuV8Rj+kyGh7H2k9EVw0c393I
GW1/lrcW/m1T+1jGUTQIQePFhLsWkxhiqxbycHueT2p91mBjD9+zyum8Zmqo/RGEKOnH+WfloAIf
FlQb+ewj5IOXzKa0WMZt8ZE6H+K0sjmv9OfLjVi7LuKCk/bIMAXVFeOBRWNlYymMl/6VWMSvWNZX
TZTE7iGsDIu2qtMtAW2ebkTgtBzrqaOk/OA2ADLxAaT/hZcJMz9xk45vAq89E5A383YIkbUgYwMH
xif8eCDUy/j7El1P//c4/CF3+E3hZ6YblCnyUdR5urKtc8eNX7GIl6QO0m91yj2pNEX+kVvOezoZ
4nW1mHn6/3VUmlF/G3EG+gdYuXOeyRZ2A08yklAdyyHvbLkIEMs4bH2JLfV8kl00iQ8WJzmlUaXn
wa7XQcgeTULoCHak2+bT55O3RRlqEZNdq3CwxNQrsCqvL2Z6XyoAvncJu93U/J7x5/eczc4WtNCt
waRxkt0RiPErELXgI4wtkPaHomRXdsVlqJJPmY7UMu5mrVa8DSoL/Ftpzu0RSUyDBVtuRTgk6A3V
hpFo7CqhwhQHUxZjsoD1hmtPy9JMpMqPJ02s2d+5Cvo9rSYnrYMh7fDPIb46rtJUoZNtitxogrL5
rVflrCiwjXrRAROpk68nhZsAnCmMxdDjSS6j1zytPuHLe9aeRsPaejNZQ9eZz2uK/quocO0iJfXU
yNIOpnMRGazXNWaAguvvOlR5QPLG7h3+dLAJZZ1hSK4W5yh+CzvNTWBopmYN4mCXvozJ1aalu+C6
WCos41lKMF+LUr4sTtNJQxu0yhSetImvjtBYl4OW5Rz0wh/0R380eyR173UTUg41KplycdFNEgHm
e43lmUghrUv6R3utrLPkCr9ndZuYHcpeLJYP8KEdc46ewyqfw1f6kPviwJwKo/ZtPi6u0460WP/g
gjfRF/nWlGuvQbT7ITql5AdUFrABiywxwhfTySH4Ibaikywh+L1o673ZNIi+9OBJhp4BNahYYe39
tBb3AwNq2XZIIhWSPk6Q5qXuiXAe/p8J2W4/VS8v/haNs3dt6qPrBl/pdmfGboX/k4E1FiRkuk0T
CTFmmX/mpuWk1jJeGEogWxnyb7KjASYdj9l0wi4Vd6tfSAPvB4/34wvipzvlMcJCv9YkVyUtHanb
r5h3H5FySB+hozKc7MFN9A/fX86LXa1rxxfURZqcpBpqO/JZZAJIweoYZgp/BBir3ccEdmTqgspi
cddmjXd4a8Zl+1ldBOcG3P7KA2fr22IO4nfgENH0bXU1mXFTImkZwOQw1UROIm5OupbGzqLfB7yU
gu28ObMKZiOl5u2V7a9SGWBjkGXmFAq6RomxakY+VPLx+di5tt6OhEVxy9DRKtfQUXm0lPRkOXXQ
tqjy2FUfzW2Y4/OAuWkx7eoYcie6N7zXD7RcL53EXf/JZRseHcjeADlQojVhIR99NoOyWOT8y5zq
PhrKr16vrQcY3abzk5W87Q6gnrV4rCk7LJrFjc9RSYf8aivsC5f6EDQMN1PP4sT3E6Z6W4F2UWbe
qbchyXPQ3sQJS6RvkXskYGbR6i7XCej66H9JrSTqa4mOLuvUfjw4quwioCDMYzJUot68ZkL37F+S
CMi9dgHxBx2IQzZkjruQ32F84V3HaQ5nCnu4N0pO4h2anCggbPMDa2Gc93ahgY/tIEen319vMGZQ
LYED/+45Vu9dMI2x79uK8LI9GpHsyVtxxThxnRPulltDloRG/lh9cD6V+KI2EWgAuwPNjTMvfpHN
ioF1+30HdCruFYglcX/i1dz+KuWqrH1AbugcXmCEi9M+gFnvQxEt5JBdfeqO+lsHh0ylIB43VhYY
HJBNUOb3yU4vT2R5TSUl7vJeHhDYigoWGjKbkmB9hUlxaJRsvEnIIYH6HGKHFaF1T13+3KL0VhjZ
m5dttR/uWe/TyZCtZc26qdkgaqi5idWtGqeLsXsIYt/9KuIRoBL6kHv3SyamuXN+GrVphRnySZO3
hDAGVbZo1ZuSHcWOUmcVMJbnjv2oo7ZfaeNbWrSawqPr+r9DN9LUl0iFlbb9sEmHnrJUUh28ktbo
yw7fozasjePZfi3063gQlUc40mJynAMAH8B1V7sWziV7mh9Ik363rxa4/RrYc6xWc4Pcw8BXLh9t
ZQvxvzZ2Sd4U/75VQW8w4M4DpAFvBMM0AnKXQLMpxCxALVdenGUWWPz0Hu0RtBvAINFamgWafF9A
5RwUsnWXzlO4aBAsm7lZop88ArZ8+ekux8Hs+0U0aieHJgHHAoR4QO4Br774jAoeYLBjPtsaf9J/
XWv+RWetbcDL+iyG1vUy18QjLRjhh+h8OeJ2oOfxmrxYtSvD+ALRIj5WnZiYgYy0DDLy45iF6PNr
Cm9/bWj34XgoEOeVkyVOGN3t7ii7stG3t4PnnXF1jzA/VJtkB5lM4U+QfLBWW8ssGg1JNykqyVIR
lAX5o4CWb3Q+yLJfM9C3XaZoF0AYvglgyn8YMPspuHAXgPiuo1AoDEIpu+5pM4ze7NSl6mK/K114
lMwA6hKPjQjKJMm8xE/kSibHe6owm9ZIM3zjEIUffFtNV8ffnTkS7ijbGBya3JJwx2d9DDnlAwCp
u2dTsJxJDbme6V2eLu2sJo8RFrpU6/Z4I5udQdeEBD9iVnR4vJvX4NPeoTVxA8R+nZNZjVyBNH0o
9q5b7zznycCm7Uqbn66KkKGKUT05S8Qm3DlykWARX+VgCfJqbh0V8sXlPH12xql7s+cioAaLaQW8
pBn7wm2w5pThZbpFsLiWopDWTyHTHmhBEEdQdRk1zDTifSaZ62M9VoygSb/+VyMptVWjmR59QwE2
EO96kajDJwNA0jIZwU59mAhWKu2DFlnIVuBiWqpoEDlRYxw8EFetI327/xit6Pc5RxMQZKbbYPfF
8eTNZ134NN5zw3UTDSGmHP5pgQhSpmaKh+OZM1hJrpnXWFI+u6lb+Mz8Jc8YQqQbUQ/WE/lEtnX6
YVb5CNO10IjlPZCbpH+vYlNPpoVw7WmHwyG+lvSLS7sRXcxOQs7fqZ7LMP8JL69H0JiOv0SqMt2j
gtNSe7QtRP25WOqoRyrAZRS3Q0e1SmvDiy2m+kouUOXfRoB0YmbgIP1P7FJ/050Le3XGmXFWqY2Y
PDzwRqBZsNvzYmMb9n07XDUcF/9K3ekRD0+oCr8OzbUZqVJrSFBzx9+Jm+NABan0hFQK2ddJKnSX
cYe6qauAnS0/E2fI5E8zzCyCstZs0pNxXoUdIpoI84kqwMGbQxjY18sAkhbBu3p4B2ZA7giZTAtC
Phd1ZepWQEOhleDQZGmyoHjMOBAYtUYOZTXBLMcqr3+tS5jzV55rZ45Zsb2DSX49/EaetrE3tR50
1oOtc4N26O5KnjDOMbMGL7oOb6xrerB3h14yV9kZmazQdMnU+86Nm8roVEwuAP/jEJunrhJbPwHW
vCgip3OqjRNAYNqf68VfhcvTuLQ9OO46cYVuASWA5RLiEfTI2x5Z/3TsQQLPTCwzUzK51Fll0wRo
zhnivQH09rFJuLgKkyS7OV8T8WmZ/lbnK0CqfLAFRLViVM9jaPLiE2au/tBW3ywZySzn0NwPwM3t
CpAAYNNDPSTt2oJ6SJ1qKxob/58EUNVBRBOQCCuPp/kwmljTtd+kko/NZ7Sxvn1OgYbH8EcOtqF9
aKBwmdPrRIB3TzNDnqL/ezhEMZxWBfRiBWlnI79yscmLK4ExBfJvJtIyx8ySwMcIaawA+q6AH+wU
TLVYtUBQ6AwQD+FYhJ4QgZV69A/Jx03f33PBFvP3v64RsrVdM1gPMkpx9FdFds1DfTZNBDJ0ZcCs
lWH4VrSC+tyHkMnOeFPcCQynByBpshZv8RUd6LDXkc5hDkogE6zwRDeZs8HW3JuhZ7btlLxrYkMv
uYTsVqGDjERa0MICf/G3ApRHmgIPiL01/CcJwh3jDuWGTOm6/N/SmzGG+O9Gikr2ZKKEzO9UFSs7
gAVdt6QoqdIQfKcPH3VoQk8kMEq6v3ss/zMCI2zyThlMiLtrwtQpGDjY2adPbl+hjnjgJpKZwjEJ
EKYvEsUtJ6SKzhw7wMvZE0ok0KgEuto4Q3iiMvzyQTSygvKAxvzRYvIahB8LSB3IO4v2sT97JwMK
CAYaNWgQc38n+4CfAz6aqzxutvMVSCW9iJkYO+Gmrt/H+wXhT/Qcz5qYYApaH2lQOQtd8QMxBCik
L+N/zcq4KLuxLuYpAv8CKvK0z/7+DAwD3c1nzlILFRBUSeswX7itycGEZhmbv8KPMiZndhMsuWW+
gIn5yHtZ1HvjLZ6Hgs9QrlXPZ6ynisX8v8R7N63600aSwYlNCyWD/WF7QNT8I47xL1aliAmEUvAH
hcjlNt0g33J2wdCH9SHT4b9LwyN29+LpbQBxS14TpVFwUrssaKb/doKNFzGyWZQ+OzOU4MyjRSUg
6NQMDtD1IHyGFi5qq4LO1KM4Vjj99TIdXvtT7MweLxegx0mb0HKTI8DBt1LTLNeqvaRXuUY0bn0l
lwpvgU0QZ/8Yif6Ix4FlO0nC+qwWKT6mL+MsW0pQBsF0QuS63K5xFAlG3+4FYHki2GOj16PUGrN0
RFOV8eJWupCbgPcsxT/deFQexcscPX+W3VNAf9a9ipoubPXz1MkWB+/sKSRc/MS6fRekEYvZOony
PLmryQzJjH0b0+MJ/uFRTb6HvHFD3euDCLaccriq24h49eXR8MoItZYgZcYk5M1lThW6HxDrNE2m
2aesRr5wTktjR7g8yQSoNo4O9OMZSmlq3cXF7GOo2GuFFOB0HmLxnZRCGoKV2YlKiuoEFKP6waDs
TzHvYjkPeLaliNacdg4+kG4pD/OB8GDxYF3gKrbhMPYVm76uIx3YM3K1ukuYWxxSNYzNnnYZt0/J
gTJu48K7GVm2RHPVJ4NYTxiN/og8FWuJOIWzkkchZY/XzCVYTQl8Vx825UY636PmSBJ5+WeYs+hx
ppIdiYE8WvQdwPAWqZlINQ9lReNxPJtaTCfIz14HuOjjr4Byd9079GLwoBwuA7F7obuchsUu6fbj
hUuNxFfaUNH5JZEpjVTSv7LsD8uViqLXtiHC23NQ7PqdfktMqkO16ga2lAbeoJMRvdjuwcnAo8pw
KeAOv11UbNlQDAnPcOCzTkWbQAtV1DkSR6MbyHfdMHMw4HhKhTmCHqENxaPPVkdlCpppyzdQEryq
E8JKM9MAQ657A6nm1bWIwwRy4aeRLPKahj56hW00L66U+f6Jp9a2fE3QSDaY4mJMlHk1w0pFEkmc
ejPsBIDGZ6S/vi850wEM9hFV0rYkUQeFvFKPVhlfM2DS8SihB797Qt8qFA+gyWbUFoCwSNO0vEDU
czVsBmY8x/sTrVRcE5vfsPxAmXfCEgrvoeLE4i3rNZRuWrnthPOOV/r3NcdE3jazb+XLx8KghjDx
Rf0JMT8D8dVhQCNmfTwZi0qFJ7j4a5oJFOJYqSF3VE9ghkJF4dfwgcNrgAPv9evDTwobXiq78S9a
hfaPWHgGszaMNp7RU7u98yqFivVlxJZ8AXgR6OPtPXfCSarSCerUgSQHY0kUtt6agLrgzI7oJ7ZW
+OGXq4zD9c30NTl5np8c1U/nuFx35g0DV0ITCfN1JOL1S4haFE4irPFbWhanqc74/uy6+emHtRBZ
zEvz9d5vpBgNJgj9xicFXkMHsJKqTQbtkgULbqsi3d8LkDQtWzdNOBPVTFePzhTmgqOaxJgJhw3P
CB4edAAkoxYZAwgEZ9x3ycrtJSn8RJ+hwQv4vm6TFvniQM5dYE0P/uAo8E/TXB4kCoBQ/7j3+XJM
RUwsxV4aO9bT7VOevaBYbv6fcCIQwsKfpawIUBVPqTliN0yVn3wlYfOg/gmhnSnt11CqK6srGV41
MCIP68lujXgL4NNdbngiIH75arNDnXtWkzgNaZ3J/Kga/ekaPfCjJsNkyyXimBD3f9+XBv+MOnSS
pLQV2Xa493qab3DbdF0WubJn2CfSUYNuwFxJ5DtSTYxcJRaEcAHUgHrwECQGXzFZdM7YV3X9QGiQ
u+RDxDGTPngi+dy+3ETnZUGQJisSxPFf+sAGwXI/hHO1Xwvr2qnfuEuCmDVDX4RbNciaMIzo1fsL
Qpx4xMxi/RFAPZpGc/G4L/qcB7HJe1lx0SqxoG/YnrbE9+nf4bL56NRYoNYTOHQzMasOMnlfzHHR
Eydbl+VBv7erXk1HA0ybd60w2CxIQQvvoygQ1X8xB5uwaczx4JbcpZVrExspn6N4N0fg0F3veYjo
CUYRaPgrMnrAtuA5fGBchOLA3wt5o6+laFOgP1/dsMP4X0jtXqMdQqxfSNfe7WYqArHMavkdyK3h
5fJSXtl3g7OKkIcstCVffJspgqFgXtXvhpXAlEOYb1yb2opBV8ZUuNs3k7+HGry8zyNWGhEivkik
tGM39GzrUAQcaQQWrWmoYxETXd/YoYFp8lfGRmIMkft7Mw9x/RP/hTqa51h8G5+vmiQ3P+CtTkR6
fiXxyUHbo3IfxhsuH2Ln2oMhI+3vgaGBjU3e7KCnuRQNZJbk8cD8bt9yNpQvThdHChivF8gDzVRI
QPzXybaR9vhFwaLjwP2McockbBFRr0ixIOByObjMje6eugYgFsPN7MdUy/FC7HU4rL/1HGmHAAdI
GRDh6FFSYM7RwAc6C004VJ2cfCC6pAadYHHk7PHRe7tftcZFUio9ET7KuXh3I/0nWD8/MvGl8kLG
e27DThybMTuSzdC55Lc5BFqxsrENHkqTU9AKH//BD5bqUbAdOL2kePGT7QmqMZBEFfzmvCxxguwa
qWLJSZnXvZuvCULJk8ndLoXoL0JEiOITQH1jT+eRY3Fio0LHDWvnPZkorCNAAuWC12AezYGOl2AY
tYxXE2J24kIFU5fo5IyAfi/i5YfloEGrQQEJWKucO8d8TYtqve/YFpNzDAtlKOqUMjB/orVHWkp3
lRDV07L41HrQiHuLzPRcFF53SiqTlzzL6CtnQRd+fVJKLxRJYJ+5sJBYoBu1YNr57rMHnc8PEcxT
q3JS+OSBj6jqQJ/OIBkcn1Gn1tABkG31DPCQMcc7I6DJWc/5Y/Vep86gcFMWzKYcc40JvPjCRclw
A66dbw3dh14Svx45ONlGI4dwWenIF9oAmkvS6k4N28XGY51KNQkP03MvjqvLbdIFegeSB/f0IXaM
SrtfkEq6Bo6izPVsK0C/8XOnuVDOsKI25MhuFHDQrdVRr1uCuCIwkEP8xcblMBEaiVzjf0l6loBI
k0TNyaNDxCePfbLVPykEerH/6xw6IIIpgxI56NT2JsuQspmOf8L0b9OQVqz9h2/2MiCndfHyVdch
mOO0QUFPvoJc3Qu3mERJWt3qnaCjl/Sbg34OhpRMN39H/uyr3fcp9kkXkay4/XeDOInvDeJAV5/A
bIm5ejHpQcB83i4JW1DqKAiA0XBQhX6MG8oPE2pfLileM+3Qq7p88hJhqHEHdoPUNPq4iLX2U/7U
ScVQ8j97gSEdnnP6NRYdx2AhHpT8SGx3/EgZeBU5JAM4XYkFoCt7rKERxlMKV7p1hiJZf0PR5Q2m
DJvEs+hyy4pGbsanQ36FpfSijiCzseH1xFSZv/y+DPaJH3vTxqDTk+5vExQrha0Od0/nBh9677Zb
AeL723ghnNZiuUzgqBhiqlrCecqmneyihdDpexMCoUaTEO0nmVbH7JLYNArzeLxK94S60VRAOaYR
DQy2Lkcw7zEiSWvWLDgoF9MyG8L0fYQJNQgwZXp/bJOl0OqrH5MCaGH6joVSNGZ5qczB9yXE8rGw
83qhMQP9l2wzf7ZanX0pxHR6dderxB3QIqe/3M9y800c+n/uik+uzAWu0QtH5tp9pXP9Tictokb6
pB1i4EmSK2xzIj2EXIQD96VONMBSwxE/dUKePIr4BxOZM9AdcvHtxuuYxb00wYQbsRNThligmJdw
Ec/GC1ewXuiIYXZ6Fs9v+F+eJ5ulsgzdA6twWFPsnQpXEHy/Tm2/5RYuIt8T2odolAG2+IW1GD4X
Pjyi0+sBr24SBbnB0UswYzrDUlb5sFl7qsiOfYwb+OJUn/Fp1cis6hFgXru77nV6tyTRMAJh+M3R
r7cDj59cXGhzM9PtqtW7nkQJUcvWD3DYVEdnApS8n4IjhplrLfULLWvzw8XxVGiOYphyT7du8apt
4ZemMq9aCXXy+lJuGsAt8ostGTbDG8OURUPj26f5/8VZOLJdo9hUOTMpaN23uwlcwv4x+R6S7pPU
uu5SabB8IbUZsrIQ/N6I0suRu5TaB5n07ZIACcrMdjVGTB1vUaZiSflwe7u0gaSN8YWb3KD9VlUw
M9Sj6I3njgCx8OH7mt9rGBusKI/Z9aw6iGzfRxLOzhvv+Z62bQ4LDZIx+bcHg8A+TSlZZT+SuIJS
+h1iblXzsTYVMQt5EhQ0c4w2LPQUEKF+K42uenRT9SMOiGZnDnA3IGAJ8JuYL8q8B8V0J7i+sQub
I2UNeb5PMikzKx7Xz4heBS27dVtUQzIUnWKE+h5r+Weqywp4SsHSZIdSIwdBVT44urK4i6D1eVs8
q3srfz3+4kg4A5awe8xJb26BrAPMH9YV5QuQ7WIsMmdmB0jKvfNHbeUVhEIpK4OVoXbrmhpKLnt5
yjaRjxgzY1X7EVxNEobhoPlu5IomTzaR03NXZaYeaoeOIbTT+j95G95F1W8CHHCoOthWWnqSA7u0
co2Ir9MME11M77jzWnEgUCloyR2NSEKFUxjJDXRX8SFbY2G7TYCBssf7uVXVGC3oOGMUzkRAz6Z9
a7YjoJoRQXmbReumNVNbPQo4tTKg/4DeIxr5dA9LlDxqNnOujP3QbhlaBYwYUXcKxW5k5/+UWe02
5Fu1TmCeKGmdfgrESufy4/N94mxDdLvjixXrzKsl0nbFEpBnhWfLhE7llB+QFDwXoVAF5SdusgP7
MdjAteNHpgYYu9wB8NDWjm0VqUehE/qc54kJfTny16FqOfhS7vNDK/d0/mXjuLljFx1Q22TOHbIa
MSAxq90wSgWj6o9VfrjA1dI72QyCqs11WDPpmVE+r+1RfCkcJAbqdj0jwYCbJhFoXHiFgVXk8hhX
9WzHsiLuSbPAAPGjJK3GZc/48KS+O7Rehn1NPrP+Dm1HgxH8FiG68cWQIjxofwUbHVeDB5MwV3/s
SV5yexzGQwvX8NkhOHUa90Mf5s304BkeAc3DbSs5HfiTaGyYeroLPxpQVEXnScxgJ2cSnirZnk9f
hobZlUy/pUhkKdfXskvqgr9/nhAgmDg58W1MMCJX9s5dnJdS5yfNn0AgA9/+P8QUqeYzefCag4L9
eEJYD4l9BRUjereIFoDlx1AeghXROEvkwrIxmmBY0e5kalgKiPprfNGk9yasQHrQtIeKr1IIQwXd
ab+CPiGdz+ZDplWkfvOYasm9/1oHQmUBsmeJyVqa8W7vOylnqCbesZfALuBtkslGcggV69cq03mm
dIrnndP239UQozAgqdFKJMn8iHuB4rdJRJHelAg4jUjJvGNWGrQNdl7ueyNwAi59t6vfPhVYXq9M
72J5j4EkYWUwxzasq8vUPmCI+MKb1mtkDlsyO8pdY8IZJwxG0Xl+9VWtQN7XhaacHX1++jbYnb7o
0K5R0n/bAjNO+jjS2Mr8EkoZdqRdqhU2+HBEazWLz4dHNfJDem17ShgAgWumDy0kXyZFa8v5V9hD
Tkjja8BxbFo0XzCbzuiSv/NOAizmFl2rB9x4WOOX6kfO/1Kov8x1GnyOT4QlBoGYokYuyrizqa/R
vCFfoN6ePIr5Oo3PnU2eo4jvIX/dElv4k44WA3o+aMmq1jXmk7xolHF0kFVodOWR/GMrnD/z1PXP
541oWDhBZ6EAItIY9lypttFsSWTDYocHIvQcjh464OtJqjSvKcJh+T0SsHsQ8CBT/AOIjwCdjmiS
JDlaybv+E0SP1n/Aci6ShJtVGzx4xOmxfWFn+ag0JzWHt2WS2JXTrtnAuV2tDzY2b//x7ig/a+2Q
rptdqra9q+VksTcjiFCdnPiA3tFy1qAmZP0FrwZaWul20WGykfzpNAZUG24YkO6/juwVS3uAhlHq
/sV0EIEN94BSL8eFlKAEyK5RLWkGC+xtN53PZK3nThqUmZa8mnNY7n1I7N6dKt4hFxUA36hZ3aqF
K+pRFBuX6wmHYoboZw8BKVj0AwTD/XPjfvPW9UAynhqDKA4Mbc6aKj+7e2XqMnPbE2/AvfOXzCPI
DV9JVedjZTx4S2yG/ecj1SkaetLs9sVaDESN9bHdcD+ueIxBykr4XLF1s1G01CefwSg8w0zTOKZh
LtQh1NBczyk3qms8uOWAymL3M3rTwfMzxhSdfjaskoqSMz1hw5i3FCr2x8O3yfzI3LtWkrL275/8
j6yxmfX362K03Vo2zBlXnnjE5qb/iPQNc7eLZ0JEWh6YSjI/nObxLnkrwKJe4t/7Xn6ynapWg4va
HH0jvsmHSOOp5K3mwrtC9YGiC2wxhqQSHr96+/WSMjoxz6k4mA/KZw2hQjA5Dm4SyZSACm82T12V
VO/HKm5VJ7HeljtiH5mnuXTNLGFZnNrxHmC2Nnr/UhzH74gZSMJzCs3U1lytlgFc7opcQxDZDo63
5uMuDsNzETMvMcuOOsICuyY7VmsH4izD4cdSjvh/C0H4ljmI7xkJIVDdNTfLdHQMXCQVEHUmNbqr
tV9v0lvoe5WC1MfIamDWDfgrXO/jMPIF7Wt1YYpmqNg3SYFeKcfu/mguL9vSsKydxxA2rJONyytz
LttDw50X98RiMiVoKXQWy3btyU+oGtuo71m1SSf0IrHXKod5ghh/5goqkdANEr5B66NWBxwe1lkF
5yDvAMVOdRVvAD9YRW5cmuxZ61p4JKx+egW1gvouDbMQ1apk3QjvPKXJcgeH9A37rienhCULz1A8
Hm6p5vSGatAcdxOx5b7rWsKRDuVXiIYCyIo/qajOToiY9tpCvnVTwK1F+FpHn0jK3PiLA7fmCJtX
A0969sYmouFMAZpQuFOKS/eRtFwI2tQraefaA7pfnETOkMV7gxF+Ney9pkNGgBdEZG3Ru+RVp9Of
IKP9/rWb+gnSGdhxFMj9eNFkcqZdA+0v5hSJSsOIawJhbE5rxgAL8fcNAYrGweR/H5Eb4ygDUUXh
szhsCP1Bod5VaUhv67ZsgHk1ByNecLBm1Jc7Ph1jGgVgcMWiLf0orHOQRn9FN/gaO+cpyEhaAv50
zqLaVpji+y7WauTiChLxrxX5XSQHx/cRK6JN4dtoua4hHyPkuNMkDkQixFIPbwXCouRZ9qzWeW86
lojdQOvqugUcwPtxe9K6aveQEmUNXOHxHHPcccyXoU1vvhmZuLhfJQNRO2OkKyvrlLgUit3Sm1Q9
J0ZSLO8elYJTxB67VlAIuxMZ52Rj6HUZG1Xkm7zYC6uzsbl2sSSRXFkzyZtq9889xdjaSeoDqehd
np5yo/8IlmFo1l227BBOdWwxtrl0ugWLEjDNS9k8kT6oolPrgwgbH3pB3yMK1sM5ttPStxrkvTTd
P0YzJgRPJjcb8ADFqAfjmR2xyW4Itc/XCegG3AXcZnE973MPsrLq/FMBOikjWMu9b2DkRQfWV0Py
73l6lRqNcqyb7kufovBe7ww7sPlTKzi8ZLMeUeRNza+psvwGizHOgGOVz7gtYX9Pt5BFt1F1aH6q
qa9HaCybKV+b2Ey4WK4BU1IN8NFD9nKQPFmJGtjXKF+DBY4DK1G0Ozr//sRnVQOag5iD/emzVWCq
+Uzne9A2YbKqlFSsJxiGDQAjMCz5Iqt8U8AkDJTmJVc5Jbwymt3XbRnXuMu2kQAkOrVDWX3ed5zp
kbRg3VF9Talw6FO6m9WZUQnypv1t6FoeBBcsL1Wp03dR+iKFjxahk7au+8V4GZtNra5Udn09+CKB
Cn3u4qCGcq9maXCd6jsbiC/PkPnnk8GeZWBShR1AJmh0mX2N+48pbxQqjWLUAXqhkpEz2gCV0JkB
ZN5ApgHKi1xDpe/xLkmwmAb1ZSaD4LG+Odl+A8iaVC9g7BmxTjh54VzTwewRl7fzgoW3z3aLCrgm
fJF3/NPTT2c1oTmH1Jqsz+ca6YcNAa7zhsv4E2bPvCFhWdSIbwT4qJ7Jzl+Uei5xGjgndv32C7eK
Ab7R6R+EjfZLwMLfzMGHKNDyQ8p6n+nA7ng3i+xPejZ5mzPiyGvo0lL0r3gU3Mg/sXJ5HoTCQzsn
0ysWGSoMgHQpQ3xNmJeBXuqs0Dyz+0lm0i6oj0Xo2RlNXW88lRFP2Rhc1TItEEE0WB4kKHLnG9PA
bfTpf2+u1V59PYIGlxrnFpJaCHyaJEyr0sZM2hlbJkuVmsg/5E9YOD0mypFuvsFNZ5nAuBhJDDia
DOxKpDdt3Ca00mKT2n8UgaB1RxDcNLabIBT1Odf172enUYenZCPAZJdDuVPbgDiYS6Q29cgwZ0FF
MBQDvN5lfHWNrfqkD1OxsahSdnNtVrVx/7HXLj+I+zbSdoNWCs9sC01qmpgv8mcId+vNw6dPxGkc
eAukkkKIFgnb2zndzKOEx6brMKl+oxW37aZV2a2FKYdLWhyz2ArEC9ds5vlPqTsKa2xrvmIN6fR6
spoC9Xu23cgFmxVSK2aSMflvNb6bvJqadm+oC9aCunqAVEQAkesQhf8YOUcEMFfxiafeYhh4U6WA
gW8Q3d1bkPC+Kq/+lTxF51T3d6p3+BWsPe7ahTFFOgZd758DYl4v+1NLuM3hsgO0Ob8nDxgtlDHg
jqRup1FJPS9j5yTM/bgPWgiyl6URBeso7MuC2lMKMWXwzrEFTte3SYXtAnB8y0bgshd+osZQYzwD
XrWsf9tUmjT4TaXNYEssOVe7BNg8CNCpuumASA4KCouxwpOkhXJxnEulbJN7pPqgMdq51Z+D68iL
mX5VA1dJ7FUoyIRJv9P1HUGySfZkRmE7qhv+J+DQOb4P/ovS6N8LO7wrsKzcCrj8AR1wImh/0fud
BYikuPgXj5IgjW5VTBWbNaH0D+QV2IbcmaygYaK514cdd8WzRh1nLezYwJ0ayonEph6EVRw+u5RR
m9QK/c0+nOcsPrWICYZNVRdvNbLefYejQf8F2wgK9Vd52ydt3jJc2BTVUBpO9TiwAKVdHzTUEi/i
M/Lw14hhZGSHHVySpXrBnDJlOB069AAxFhSxOeSC8NuvEnIvvbDQ6warWhYcyDTN5FQvsxt50nx4
+GQSo8oWJDLmc5OIw2O19EJ1QvZQlmizKfUuh73uuemA6nmoC1kB3FXYO56p6OSwGBm3mHh3fIGo
Ym+8tlLj3zVlAQvJRzOFo5t7GMsrIDSlF1IQAZuQyH1MJeqUvFosdHyLuqfblsmyjo2C0wlQuBGC
qEe3tB7TPTspCEw45Gjqjl9ZgDvPLgNDQswojVhvhr6UjpG1DbArSXAHCD8PdjXA9EAToOs5DqaI
73IJTY5ztni1hGKEb4pTiurECkBvj4kSKkKwr8F4aaKS+8KXPmi/eDQQ6oNrqJuFYATsiL8syFvU
P5XjAynFALB0f/Yui/cYmw7syIt0EgnLW+1cVo2X+HtAhNvoIRo70nr74orj+iCjFcKseY/8K6IC
wmB0tytQOLqbQctfXetzygsgA7Xu3XZxRb3AnaHAw5KSBaTaKirw/onc4HUHGcMcoOJkUiLBdDnr
SC6uLSyu5L6EBYwCfbpax4qCQNoRWemboOGantSGhwkdOwTN5t+TfyVP33dMz4ELYgJjOWVkfJml
XtEX4DKASDOVgGhX0ylpcLBvgUcgbGLVXaUcKVUHyzKNODOnfTudjo7hArV3pSCWHuXB/ox51v4o
WQKyvrYFXX+L87JmiTuzxABXM1sxb6EA1L1m/pGy3WQyQ63cMa63aPWdJ6iDOJ1EFkgeJXWa7XwB
ZMlbHN2yGvVIwQtGNkW2awGAtpJJ+7YPq39aZzkve/XzoMS2GpWxKwigVyPonaVznTD7ahE93YbJ
/eMrkYOVbG1KCrqmKrmO+eVK2wAimlhvEslh02QmZStKtcpbEF8sdJd0JLfTViPEb+9LsdoRZrNM
MRrLrs3JEd7Znql9QnMbApmQUDglZEgsrR+GQCfUWOJkpw90UNZJnHhsql2nEqWgw/FVPsJl8/I/
AmvWymYVuaeBI3j0CoycCFhAlU8rsOLSYGdEVw4/MbIyS9Ni4LYIyYklD8bWTZBiF9PPSjyxGJ2r
e8lMsROMDHO8mOStkxp+eveeua4X4AnMnjuO6VmffhbJ624JWeMuEizOVkNN3C3RZRj9cye/KxqW
0cmffLzHR/S8QhzHMDjDFzJH6Ld21SlTJk9rAJ7TwMfZH2eiQzV7M5DVTemqEsoX4pdD+zRiZDm/
/wuOkDW36gubY2Y9FJSpFle02rd0ZATW0S+xr+fsX540zkSaihUPgz1qFi7wd7jn1XnXI8TvLKEN
sl65deAI4HjwUpUsvu5zHIa3pKsBjkT33M6dmxGs/pBdjR+yP5uZSIumCpfDU7AWgJEUZ+EMLHPs
fFO18IkbmTgaEUWxcDGdDaPQnVilW3+W5GrEMkC2MbzzCKj8ZVNAmRFC7aqH8PbdObvSnvx764li
mukzUjIYSy34tk5+tFfSxEBBrz3k1NXpWPNfFpzLHPVZUQLtj8vSR9BzhE3AOy1aTiP08pjsZg+F
0GbA9uAHn9WPNikLbDusvow4WduS0dU7KNlqkdzzygq8Odxx6j9oBQe7PUiC2CrIiY1BpPMYExTa
u7b56+8tzcz8GU2dSWb9DIgGsCJ1FOmXXOXisXSN5ML8xV9GfR5siRcE2AgVxyMVYxCvNaO2u2Nq
763b0sYbZR0cb50d6DaxO3691vcifkyYBiC5uTL/vWxGNu1CnvCAwHzArn38rC2FOsELALyMiD/L
KCXfrfBd/wURSyuOuKu5DIJRv9k4LNhU0ylYiyMK3dtNgB6jt5v+1YEVBk1dEzxYxWaIeaAhIeyJ
S+sVkx7xNtF/9SYbtH940Rc9BOShFHPAsqySmyJQSSg29J0koFe+XuMGpgOpIlvp1bMrzs6ebYC9
7uVk8b/H6EeMg1q3A3uEEWtUx8P62lISCtTrpe0OVeBmuUDJ/Jfwe5It1Vut8jZ7OaINKxTLJYgH
0OkMSzGocLn82Nn120JgNxII4DRetn8nQDA0eNX3jKHE12Wk/Bx18p2ODGdWpGJp8NVPk46pUWzb
U39um765G13VFR633/C/l+ml8gdOD2gb0rzJld5cAuXRWfflBLl86lYRKb4hlHU4xblE6YsPCbWn
8kH1ujk95/ipnvsVlGUPcyOhTGnK/9nCiRhz+kTP65xEYkzddNR/1CyHfpCIob6kFLov4zZdl0bh
cyRGqhmPahHKhkOVfgDr+g6Iv9+GjZydDS8R0QuyH28YRcBA1QxjBz2CkGmisWCG660z8A/QMcyU
nx8b5N3caMNYqTbtR8nQE4uT0TbWOwy/kevBA7HQPvWR8mXKC99aRRF7KI4Kn/AbbxoNavBUqeIv
CRXbzb1DP6qUp9bqD0Gxm61GR7clEO1V6W9FL06XwZIorr5WFYkRfRQ51A7z04jEVDDqOtO0Zx5W
yTwL3mdO5xevXvTi7YwfkLmt9zQ8v+lWwnR2mF0MPf4aBmp2rq/GwR4mn1dLKUEuvZ5Qp7VZZRoQ
djXHYKjDEJ/Sw4+9kanWj/wrdSuOw8MQnNngYYYuP0po2eaECxpifSUY40kq/XmowSh/wdmft84S
kcGK4uXR+zUk5Fgz3sNQ9eWPxUWrUUUEjDzr5UyMGNtetKWv1KY12k3hMBmUeYxdfpZWFBJ04T3A
8egV7rfdwrXecpKykY7CsNeffstDmeyTpr9Ky67J81zDtkRYO4ftgNDqwxKaDfTJdl8ZIKAhueiS
3niJ3HFmVbnOk/AvkXj2JJLOLI1kPv8v3z/CcW/cGU0mxOVHO4ETw8ZvEp181n1MOmAOjXQxLHVo
aKzkxBVFM2a4CyoLjLsgIRasSw9cociTmsO9nkpJowimBDdA1bQYh8E/lpNg4bW+tcpREV708EBH
m3GMIOrrCeAXQZsQ9PYd7EwZcvuk9Ank2hIc7VyrQyIqhz41mNCcRc5YlQglewPzmAAxVByINpOz
P09tB5kWv3iu89baFSKbTtj3sfrcTTHi1D4VFVrDyfWlr6NWoMZYd5V0ZFA1q/KvboROi4mtZ0pG
7p4xt8Zk9/YGnCvDKidvGPoBlJxZ90uru1rviM42FEc21imwIHpX61/tdZH8UUE+knCu0K+nBk9c
zGjgv+HL//lmdrf99C7e9/E2OT82+6Fzft3O/4dCH5+12XWnydsQT8Yzr4fBJrX2bmYmRplsrBKi
lIIzgDcF47/404YMcO6EKGcES/m3iIW2gJ6z5PTZCV2BIRuae3VAuXzo/3Uthp6LYS6AHkaCeS7x
DIIoQ5vpSKN63PfFVHX9GuwxaxvjpXPAlkv3WsoGhkr4xZs/B0aJKiW+gZ5EpmaVCTWcmG9w6v1L
i/yXxpV1fC1RK1jwV6dLYdd2E0QNq+kis1GyTVdnsCatF/7CF8xrwL4z3mzkZavKsyUbByekcrxB
vPD38nu8xCbs4SUJKXWrHoPd0IbyMudkG/aEOl+mN+85oQcbR+SgJrkmiSXkpnwXRtBgbfzWjT0k
K9+QS2v4pIaVo7PccKMY5nrA4qstGEy7yBsGm/zTk5shaTR2/fWWwBnLFvRXHEuy/78b3CHLRZBn
c2FTJzwK90/x6LE6ucEzMMXM2ghSIOtbbqfVYekuPr+Jm7ofj8XPoYhoxTPuTW6m626+Y5FWJu4C
jBlCjY9J3HMaN/xW1hYFPAZ5bIearNAxcZ/qmrDgUR8U6+AZu42N6T3fkxg9DcyVMu7Kg9yPMwxI
342uBbql80WdONqbO0XrmBSMGGPJFJQgKg0lEvPG+9dSScGZtrEwIN114q0R9A2AAV75menjlOeZ
IlJmabs6JIM8KRVLx12hBCKWLyfst1qCJv0PAJO85BGXdWL/Ivu1ygeeVjySwEtubf7I2ylaWPGq
Q0hvfGSlTfPpjWuEACdxht6f41sqi6hOUakj7tydcBaTTmDN19yyJTPkm+hcCW8MT3Q+lvTXjrDf
XVDqhwEk3+6tSLEss2Iaxr+s4HtOpIN6VE5O/e1wSswN4N0vmXfdWRu2RBzBfgt4x/T3Xwf7OV4E
TLx8pMxLvW0YxDQCKeNRFvhBWZv50cAVOu1V3Cu3A/xQ4QoLfXQnz1636L2eYFlZaONoB8NdoeDd
9kMuKvPVdc+1+IixxPPWKGpnrHpD7E8BHrWLnNiPATykHMNeIsfmYaN9UgUCD93pzuZ5FrJcsvOX
g8D3TzqmhsaX+MaE6rJTOMLAt+VideD78d+2/5mKvzo1iyauO1peLPDAICatAib3DNjjPyvOVo7x
MJqx4+83N3URzjBcNn8q7Nr1vPS1bdCLkLW3B6VTolg90MKpjC1mXA5h5OAoWiZkOrvtqTfB9Iyg
4YQ+4fYF3pUqyphpQF0dHYddve9RMAXYubP5DcNbeS8+vqD9NSzjRScOkyHULJqyE7UFfwwMwsGG
JmIg8cXlnOzdDnrdEeNejNolWGWdzbd+zR0EmCadkk3pubcRjT1YrSkacY78bSUkQFK0faleHFC6
EIQOls3IY0jFXsBDEJfn3I+Aqm6Oiqr1E1zMWujC7sYgtcvQfkmW0JHelR3iKoeBHJCjimSxHhKc
9W/zfQfmB8ABJVVLMTN9AkHB2CSivAyU4rlGhky06O24vJNbE/W3NECveh4wkFAnpYEJjK5ouyeJ
w1SLw1POA/mu1c+8zbzhz7rLg/7SlN7nWwPzkLWNXr+qP6sD4+UueFBdhIsEbOskaX5wZ6CNYDzS
FV+AYZqfBy7hRVqAje3zIaHNPJcAox6bjPnbdk7q+5/93Zvd19Gja0F/q5yT7C5i8M97dUWhTmsa
QfFskmWxnf00hzvIb8p2IWPbBR/S4IlJb5Ztcb7/NMFSM7x2oNv5rZrwhqrooxrAyJ3NtE4huvgg
pe2RXh2+cFa23rpf9WwMx3ScyOYPa7ed0MibPoAxapv8+4/tDeheXSvxeCA1fD1WvgYvA2e4valV
JhoqRNkSAaDsbO+1ubX3g7pgpWgCPGdPt0PGtev6GKFdI2bu9e1JJJwGqrsdSRSyD1mV7NVUnmih
XzLVLllIvgrGwriJMNofxtqS6ho0W0WzlX3+bnYwbD1zQx+Jb2OuCSSEaOfc0F2vApZqu5yaNoUk
fR9wOO8XMADcSoye7ljOajPvwz7XphT+gdtHO61QEtL5zLfLOe5QnMnLCIU98IfG9RX/xK+1EKnG
s44D7J13bUwqxPe4bMAFq/rADTrMl2uBZJzEEjfFuKFVRwoKIwrXYDrPqGUcg8lpoygAZzYaKlKM
IMzOnQo4xWj4Wr3ryWeGGO1ktNET3S7o+9YHqntkBqbyB879xNBEtTLMN8WmxTDYtqDTK5LH5nwc
Jce13yEghDHBQ6Ni5qY1+RpPiHsXm77wHjDeyTWjg+Fqc73NPtaxneuHXCeKutNKeZlpXwZQr3Sl
MXbQfiRXpQBSnqTlFZp76ckMQEcu5OSGWZ50tLkVqZSqFnRrkmKAtBL5g14Bta/hsNHnlx+jNY4U
6aNmDD+3ExF1NXVj4mamKu4Lz3X/Shrsk1vWJTX0HQrr2Hek+NLcATTwDpcOgavlTCeCsNDCBRph
5H6UvWhkVbXfcjIzqjndiwEc/YuNamBWG2PLfcghFiQJpQjTtWYNQweJlkAcZ30r5Rk8iRAyULNx
f18mnvsIYSAmJOKk+6us1tpycvbcLKZFj+S04XzKcXcQdiczC4oe8NX/bWOJaZ+YLOcZrfvnzNYx
kspk3LLs3p1TRMIfvkdj/sbvmKUlESb6youJ+0In2u4TDj6F1+nX1TsmTiSMVVCyTgkSGM5NQGSR
7qafsX+vpREmJaS/mjpWKbRNXd8BH4Vc/GxWqe0CcRNHt57iqYPntfkiNCG+B+3pkGoO3sKtq7AI
ShLKrAOqD+ZVFV/FHcl0tECTLKgKvOwlZPPV1hA3xr/8ywMcJWOUyKw/rSgT/gZ0oGIkUdFRf9Mt
LZNWVkNLBZVWQXAXkWR0azpLTA5OE9ZsCtTqWdp8qTDRDoRkkQoJPt7JZHFd5rv+m5t1WB769w+V
kgCbKqMdFF6ibN3otpBkrKFnA/me1WGncKzzO+31cBmhYbK/ztur9aNXTO2uR1VG7N7uw/7DQwpO
ZTf+rE/frwEPnlzTDr0SDoFFQEGSSp2BRZ1qZZfruYIUp9D6ZuCxPOl3X0VpdaIxHLB8eTKk3N3W
kLkquD/4KNoyShhuP7S837sMHlW3fmT7RCMOjNPQL8r9wLlYQMFdWUY3V9snfOsFoqgT4Aqic+bs
xNZH9zE/dn5DYClQey2788P3C7x1nCbuba/3in23BUpgvI91wdbWKhmey+1HFt6Ny+eKy3ApGd/W
XZMuvgGvDTvB9iQ+RYbQM/kuEBDGpbf3w0MvEkgFVJWD7GmHy4P63bTsstkRLxgpzgjjLxeftXLn
X6fnc+gz3aAfmY/9KQLh7lozOptHMZhje7k0+QukH9fDrYm7LusycXcqqfQTk0Sky1I7xTpeQSAr
CVopDkzOAii14kwPtjZGy6AGkJx6mI1yjdaB8hYvSenddRONds4XpuFnFoyqGq8x5vPng6dKvHDN
CU+8b2JH0Vqstu3jc2ujTiODU/2E8i9IG0FfA8IZEXwGbwFA/dvSNBASyvERJ0mMxsCpCpWAX/hl
DRwaSNblsVeoJKZ4squyMotbE7rWJmE3YoDdJEINJVIVrFiU/ccWzz/lahwPZdh7u5dhqY7ohN4Y
WA8amOVXC+t2yjiyha7nTzk5ZMaVQZ7tOMr4AQ34BW4IZ6FdRZ/FuPVKqwwuq8RFxrj3Og2sNnjN
tF0lnOZN//xZ5BQEgnCAiaj1hhr1J4JKO+k6Rkbx8aOlwb1e0o7clO7xoLyLleqVEgTACQwZuEFU
FTAxX1GBcSnN+xtHXLTAttsl6g/AU8xCz7c2qzz9EauchKgJKfu/GJDy2Kj0AdjlYRPYAkYHztFu
c677Mfzl10955JjkoXgzoq/+IlOMkmhZqcQCLMOWm1YZHaSM/tznj+2WaltJzEq3Fbg8z59eSgFO
nfMKuXQYzax3Mo4Oje7usaCRvF7yjcoNOM0o2j0OELmpRC6jaGcKtgkljYhqT0jiA3Wg860KCaRd
9wU3YrLsGDmQz7ceiZ1Ikcw+06xv9UysGIcwtZAz6dQUi+DazNYAM7ELx8f05FwcDF7kyuNMDmdj
qmMhmCGV6KYlpO+m9p73l1CjuoNmoR3XRG72CXe+bHqDXQeFX6ft+saIaUibOBjTrNm9xnMENVLp
Auu4/qASwzixeIEAmrsFwCRSaW+M5h5yegglaJHdC7T+maAKmYS/TSetQz0vB4m5Pu5KpJppWFHh
igMwePUJ5DDBQ948TRPk0zfrlfZrE9dIZXE8c5sHjE2XgjuSQpFWzcl/2flwiX8vTzImRAMFfTr7
TZDDnI076958JHDa4LqAlmrwE6tNa5XDQhHON0YT3qveenOLWFf8ZYz1py5QMQIhDXclVYfJGUaE
csHY2emyxzAANdPUNg2zcBJ/RfCr7Qa1IhB1RNWOiKzzFdq3V1pCClMobjIXcVB9MlnPbXEfixno
L+KlJ1gVh6XiMmbDF0Dmrr4bbpZ2hbekXuM7ll53fkoTD0aM5nWUl8F0etpjsb5R5It4g0nb+mUw
r+Ah13jKM4rgGDo9YyHJ7YGcm40me6qmfJbkmiQ05gbzPHUF18P+E3J0jwKUbWYq6qAaKJuEsb4q
4Ow7Nt9oXCGp9i2dunhnl0rrSIZQtxwQia4wCHxjYTBbtj34zrfjFSCexoR+RdlF109fJ7Nq9eA0
0jfCjJeMsPVXB4qw5gJkVfJ3ytmFwY6YRMLZy+iz99kNrhP1UGWZei6NYQE05aDRXqpJQKPe+X4C
6xX/DjLrUADlACqx+4jL3gMo7TJEH1ne0Cr2Mdoozz/iQd5TCQ4QIh45XKRBXvXShdISAWNxwXgJ
/KGd7vnNLqBIe6K0sgdWB9Wgm0OMtPfghQH03Kbg0bUEySKSPA9QtpLMfPZkWd99ldhMqaU3pJ1h
daga2IAl/miPjbY0BW3QIdU0Z1BwWADa4AqbZRhANv2oYpGPM1tc11CYjaorUmvcnIRanEPMU5fV
yeGtrrAivchOpZ96XU9rdHX2svbNJYoZyjDJhY58MI7sNm0FuvrVWfsKl5bsK8RV5P9ssAens2xY
CWUhjoCmF6GioLfCydj5wBi+x7ZcZ61JAF0RdYppQeCpPpsTOtMF5IFnRCnt89lacmW6ocbrJ/PX
FNxJtlDt98wBrTashx0ObpeBYhe7HUMs7RTuCnQFOs0hKif4Lp5HqsP085wuUn1EUWLRR26JbjHN
mkr9dafKWyAChdIj24OhreYTFS+oyWyJ4TDoxaubp/RNnQ/ynyXsADX8nkf1/SVPuB6el6XuH+QP
rH0R6e8qTpycttQAsA3IQLX9Ek9dL7r+c2nz5T6faUP55UzyQuJdbs1kQLJ8RPX+ze97zDbb1UCx
ptWH4qD+vlrkQf1bnekj1nOAeA6KmSjszeAcnJbLocgpYVO3feNMuZIm0UllMtty5kdyTvnz3V+0
sKiNMu+ttM97uhW9KHp8HU9Y6PVIFBBDQOKGmq0qZiAGD/YESb2aHqh98Kak+X1zcQOMI6irMwbF
rtcnlub+CWGVpcrEB/I4NOi/TjZegXOfBVqjD4ZF9x2nYfvgsipktF2hbwg9ZuReMItAEypH4h/L
RvodfkmKG4AZpnOmcNLLC6egsxlqC/K7oIMtoHrKqhGMDjCphhndXp+9AEgRybl0QmdFotwUfGeI
EkrOZtf+cU6tFqgKTrgZYW/vifE3GooMt1JGkBJKOl7CpQR5B/4pCCPOICyUmQmgnXUcOFhicFNG
cG9mUc4jyEh/mUsXUoWlM6U3mlQAVIb8a74unJgsz+3gQZAB/2BThNG++kfCk3P68CAeIUgRQJx3
celq/YVdRV/OEUZAIbjzOuzk8EteTbTdWKQJ6+5wbhSGqsjCBzSySno+7d0kEymM1NrKFgTIbHxQ
beaqrNBZ4xqtkDbnY2g8jWdSXSxDa/U2rG3NXJWTaQkINipd3+AXWProt9FcvA1MQk4CtffxlDSf
4c3gi/rwHOQhxDD8p8hLv7iDbGWWepny6n5X+N9V3IWlrqhtUbivTaQza+JxAP6H7y7Jz2On58gE
3WGZ71Ph96jNmhTCdcVjSoc9XYPDYE/xqcEkoh7e/Qy2cyIy10mRPUljMenSeBgbHwsKlISDGs3W
wzDBQXWzk2MWc9vTa6AKHED1qzaMIYSWm3+tfqJUJr3JBN1mo/evfhbXwhn9CbhW+Fb4w8pwBo8Y
Buzf5wPZ0W3+xtwyXDHoNW0rM2PCtYexBmZR1/cGlSPP+OaILDDnnDER86tCKoqCySeHSj5k1Wp5
yDwyxbcKeqrqEWx+XZZowBOoPzTwxvbVmphcM6YQQ65bT6xsRhZQLGI8aPUFsvhtSYB2t+ILuo8g
7DtddkhGApqyx9ll/MjED/53u5AiYSGQxAHmgFNcFausEfFoadiL0lLJ8hlZfCxq+UHYu36OUaYb
Cdjf4UlTxQjTPmtNXFrNLUUkUgJr6NdW14KIYEkLLYZ6uSKvctLt3Dqm1MmdQkFBY6rm2kjZPvjC
MbuooKlLYCt6FTuLNjcsyA9DwfUb9aQ87+fHOuTdIB0yT8QpXbXWanLo4o4Hu0UEyb5TOSTf2AX/
EcHKsiYZ/hIQ7ubiwRpf2oi7S//DtvsM76awGsRhdPMrplicRIcNxJw9cO7vwrulwZg/HJ6Og2ST
6SwVwHj+VoMqxEW4Zw67QTXYdQxiJgl/nIOPhtRIJLbO7y1RoudiCUAjh4qUH58PLDipdnbHymsZ
s9GPGTuGTvNoQNdv7UWr+hmbR7EyL+8bMSmaSuY61AHI+554ZhNv/ZsEYXfG7BLRiCKXk+psBFwH
R1GoAa3cWU+b8aMLp+lRm4uZiJkvozxM2jtvJuvltj1AepU3QPMeBxD6b03mb08mdvryTt9vxPYd
AiU6wxI5coowR1DcVyhB1UK+lXobxmZOFZcIxiBbGjQiegI7Z+qfjM/lb1qCVC9KEcfOSEiVrFO4
DQA3o3xqIzNIl8COI9N3a0YSiNJcSSH/EFqgqlLhUQaCx33ixmA/6zSWTbohRC1PTYOKlzA5m5Kh
USDaNHO3kGb/rP0LqjPqHP3qkqVb+uY2utvXv0HhvyPNXK0kHMNRNmJhhQaQJWS1+xZXfLktjYks
LasnLEO1j5RtzoDUaU+6gVrrPvuwUPYX62vACh/BbHRJYsfKxWxdRr//1LjNHsb0C7xRFAaKRvVY
wMxST9Yv1/S34gou8JVzjw2ANFyMYfT7w/dPCDHDK4AYV5R+8WBqHIUB3DPzsy+T6sVTy3oXGo/9
1vMu2eVRF3uGnULjxSZz+WKvNJDxvDKfqoiRPO6C6YYDZtcq3MUy4j3vXGcfIdQ6RIvBoH4XuQB+
2SBqnjb3SN2Pd9f//mVVCQBTwzxw1v76IffZNUCR9tVndyIVeCcAq/nj0A0Gq3kSY1dchwIAqiWU
El64Z9h3UuJSq9R1XQkfbs6TTwYQd6CpDwGKL+JVqjKxopYwtWXO3HwGsV8NIN4Zf/mXiLU3oSNY
XppQMRh8MkQwRhQeNYWc/tXuRO9RvXmOyB0o4p5QS7WFUxDSCFgMDQkgaF1QRrZnFiOS6iDzvltN
ebRgCjxJmfeHmgPFprVmWjGeQugclv/VQ2NruU2GdRmXlc0t2TZiIUqldooTeSqka3MalXe/uUi3
75FvO6R5lMq5kayOjSrPH6jwqJpz/aHTfFnRmadUB5hMoyYRJN6H7obFpYnEOK+8BVckFiNThGvx
xssFLM/8KcB8vPkTcIkXhd0T7HDr1uaB3P/M/k3d+WtUfyTPftli0llMHQJ/u2z6yf5Qy2oXzilp
Lnc72AmTCQkv8yjR+QGpXEVhV/iwa3GQlCFkW47SfAEiOsDIF1t4VhJxHBI326oMzPYWsXsnAxNR
0vcte2wkL9QlyPxC/y5GfrSvJs4xnIcXpMk0cLgv4LntSCc84eB6lXWpuhxBtgWmD/sKloRceIae
UsPyRaF3FyMRCqIdJkMaUnv7TrtDdO2fdhrIa0XY2u5JQa78ZP84nUAnpGUALik0+CzI6P+f75Pu
uPEbhSJPQOk9tGmy6to6vRwQ0NmdF2C7qInlpOTNLEcDkfmslr0rv4FMlL1KKO5uvnv7NMj6RIaC
IcN44uUdwywDgao1xTdZMADsk1mPsCgVkYsOOLAkZw9ZXR9AfhUVqTd5ljBEU1G3/DjNt6wQqVZO
WeQ0ltNhaxSar8Gp6jEEy3FcVS6QjYSpfFLMwNdnNWgbfTwVH/kdePu8vnxsqofixixth+UGsnuy
+76cNIM9KwGyeU5xmRqev2z+Ml5oPNK/x54qq1U0724h6kqyH5P0vKcvJds5xdJEMRWa02aOKUQ8
gOnRcOuRAhzjf3c8gPbvIApQzlA6+APzqXLJeiu5BvrVjV03xCprRx+Dg+343bFSlYvIq6uENkuL
4Kes0y76Ucr1hu6myn0GB3OY2gSh7/yiIhBHlxcexljX2M2q+dAkPle8KiPNn3QvR4aO8rB06+Nj
ggzaJgTtc8i6ry7BlXRwxUkQw94ohGdeW1BeeoxrU77FpjPDIiHn5JHa0yfGwY3JoBifgfmwenfU
4TBPPpq9ABVGFHnHqy77ygpQdsrjtZodS8de20r4nYfasX9vbMVnTdie0IxpxDapXsty7I7iV+G1
t5nu2wwFsmLQycQ4yKWCXUChfVWyGdoAwySFos/o0Olb+753srTxJqHl6zgwAcUTHiV/zCNVqlA1
/Fubw1ZVlmSbPe+M4WWbvbCxgIrlniNBrw4w65lg3oYK0hMsWg6eomCKe+X5gj9W7OYCs+Yl/Rw2
dHLCP6sbF6xiPwJvXVJPy2rZ3zRNNJBmfNbkIKIFbP0mp3QyBm1FhNFEoOkB/nAGGU/mAbTsaRRh
NUr7mw5E+x+MkvROyOnddbBIcA37lekWz4jFNPLoWS59KCPzbpsxPUnWai4z8c97aiCEFwLlgbee
6okKeOdkl8snGhpvBRIwOIkToNKcLeImjpZSqWZppZQwYF4ZWY7vIezOZoD68ONTpkBE+ArdHA/l
waeez4/85lcz4547DvocKEaBrvwbKCPR9yofIPmneg0fBV8iHFWkUB0PkpgxooSd4fQcXj685nXN
hzVs/GjpAbrOn9iGHmWSOtjaQbYwhUCJzNOmYUP1O1Uy5KT6R2ssYsordltXT2bBH1kWv7s7SuQO
7FBFutOmIrD5eE2S0ZvhAJ2qJ0ebYRV39OCICR3PRWewJCMNdR3Gml5VIYu2ClYJmx1bvIm6ftwv
8GXpvD0a0+XkzOMMcpC70hWnaG3sKz5VQvth1/Q2qt0E0fSC+/fXygND1Zrz3z7BQ4ROFdftj1+8
8kW0hnBiq3AQlYXZLgQlJQJowSUydW0li1OeDo/iVZpiOsfCz/8x421TNqVmVoombAsYSJFYRCA1
lawvLeQzI46jzoDAE2avKxJX2mbvSoMDMhJZZOcOsDjd1iwig32jw0JTEu2bIgZbFF2nGkSNPq1W
QJAe5N0YRnv1b8GcJV12q0PFojZcmYZHKUA42ir8Z9CAJSnS/1GW8pZkD3E3oyKUtJrjJNBnCATn
sWBK7yUK6rTmvvdfWtOezjlWjwx3I8oaMrH81YgLXG6nnML+GxGwPWfxbWE+4N67G92JUcs/F46E
6806PF/p1GZRSTB5856ToY6X5XmJ+4mvn/yT7hVK2z0kXhOUvALBe6in0cuhjERPGfZKRiDJXGuD
aZpENnKJZjBymjVOh7K3pOhhtBxB9B7q7GMqjqcG8L93c4zaQAdGXJ6EQZYfUK45RmkccDdzLl7t
7ZmtyvQInf+/rZImXto/9igkwROCVfr1WdBWfsDKPzOthm6worxTKXQvNIyEQheC1w1dqq+RTdfG
82XS1UMCyu4qJTuHjAFzTUvFW1/PmVvHbG95UWIgZecOxJIvi96fP9VEMjfznB3n+74lZ/wfw7bP
9IKfq5LsMgsPBvz21q/ZreEkk550B5p67g53Vhr0M50viYsS5JQIZyPqpXV/12TphxBP4QNAwj5K
vCr3fR7B8xOI5VpzhpsfFRcuvn9r5Vly5xWAVqhRNwp2BjF1KB45xqiH7aJAyQ7Mzl/r4sTHla8l
okQTkHFz0w5tVnQ2m8n3nfjwDyEUaimmvJDM0AVSPUVfg6OTS79ykLnSQNaq+v9SzWP8qJTCDnEp
g27tVKnMHXkWJv+a80WF3ITOBmmxN4SCSJ0jK684tcH+GLd13G7SltRE4AeYCH/1iyzlsjxZGHTM
TROV5XJx/0CQFF+X9BnwBNxYZtShJaknJPswJ6DK7KHrytFDIivZOI3b38gndAwMAcS5rdEPT9x9
uvBNHzzhmgi5N3rlU/aoy5lciJ2SQRODcHtbuMEuO6BwUP17xFrdT0ZkOPB2eCKbpqhlfVMTIhjY
JGhM9xc2cdPwtYFO7vabHn36qXTiXVXq6+HmTnseo7Gs3T9m6FuMTgbXhflA+wjY2sIGQd9t/9Ae
bKf7NpmI8Etdc71TtBXfVhkmk2TKptEy4JaU4zmiWfRjqQv2U1E1swfij6TquFfNiYT0fBY+3xaH
E/S+OLiDXWYI+ZvaeJhsC4/gYd3/noY9aIhnJXsmbxjISPy+ZZoX6M9BW5vi1dpyrsagfw7RsuU8
eET3hU5sivfVHj3HNHdn+fjT/2BuWmDNVsPiwqscUmdjUE8Izg1LLqEc0g/+1wQzjdWgmIwn6j88
+mdNp9xKRj1JHbefBMggDtbxdKd3KCUHiswtv9TjPnTs5/SsImacAUX3E/4xKGiTk3OFYJgQJw1H
6JyrYR2G9eUcVvzEoUJj7IW3Bbt25Ia7k+s2+vvIxnRrkNWN4KYEXrIMmFS41XZNn88iaAWFhDGi
7bPMAgF707XkDBzQZIx3hrbAVO9OcQ2SkjqEZKtf1U85xsHfMLLLCAtDaEIFInRFo/y76DOy1nSp
X09DbUQvAZ0wXC+qSmmpZU5VhFLMH8ULJmo6FhQabHoxS8EkDuruvsNjAwhth2Dm2GVG9njLQTaU
ap+fldVUMSi01MhCxLl1YBtkYxtTDy0o2jsUZHxIqKCQBy7tEVZyBULKlJstXElQFAWuwKgnGjiP
eXX6efKWIBM9/+MpRATq6ePMax4oG/2tFJivilOGMIUPNeT/FGwNrV8NKxAOTTiCKIxWJdHqjZmm
WsBmck2rzt1pmL0aBt7fP3+AfVkgjWmrjQjkR++xpMskByTlwnZikmHlseQPswH1O+NGGIGy9F0V
9165204yu9zu4abAkxCkkb3HW/SI8q156nnPx50oBpOYPLB5y9Q103iDDHNb8fDUPArMmjqRKXwO
IXiUU/8D0+8Yrjisq3mbYpsSN1O2KwPh1BVYMCczRx29eaK6PckkMhvTZwEfsDN6RkRHtFtoqbzp
plyqP+jtIH/CDfCEZkJMPj+50ppS4QllixjCoCC+o2xB/Jy9SDVq9FIf0w6ZJQRAe0L3uopR87tG
yRZ/YK+oWnbsHlWtuAOfJ/Lc6UeittrGRcvF7oc12WYlRI8IJqDNiWaGghFZ2HTeqxD3K73RGEhb
kVW2BY8eaMNCewMBegxiFxomnNCPp1gR6d4s8DHWnq51NUY6dop2081ir2iQmNzfIHJx/bObAgKp
2ggh6OwtKpJxUVAw+VCKqNlRP2H+Eaa++SbdHkHo3Hg6GP/j8TWtz8n5pao5ELej3KkX7Vohsyi5
0RlMacUXGxht4VBXz6QmZ45ixpjgEFZGp9zDO4nj/p2dqym0QQyV/eXuDsSHX8OmC3UKWB2TZ7so
bhQwI7jFcIxYqikA/ojuG4kC4Dn078FUhlx1H+1AplCrn4TQ/DKIInk9XmgFtPK5xQIbNHX9mZkd
A5daw9QxwcPe8JSFDwyKqSftqbPonwB+h7wytypK/1yMfrbnJ5X88M6QobLyxaRZkyZffb2wJ/A1
H4+vVMVDI6Vhv+9726eWLYpdbREbN47Bfx1AtijSo8UoMdkKJfTP1TotJKik241spEZqAyFuYeb+
GqDQNnAi7hN4bY1DCmLqUuQQ5/zlZf1uNtuhkrz/Atr+3CAcqXz1HhwHzNOR+aEjP7fhLl75bdbE
R02sWpgu3iwHZZ6QVq/DjTS/NQSAtjOa9HRVOS8YUnVn8IWtb0Z4aEZbdZracf4um/BLIV38aHfZ
TBhzYB6mdsfI1Bs+z2fdIvHygWW8d+Y3JQCCNWOAF8oOVnN+eVnd1gkkDz7pzyP2tdmXokCqKNVV
bMFs8Y0mo4cJlDXrc1bU65hj0Vq1CNKoMRoMSnWEP7kjk5HYWKYeR6rriZQy7fXFSWoLVvtLTWCm
Xd5UIyKjwkl8GnMt9JYn+BXecvQ2qSkkeJ8JjRYqQunUTL0hE7eDZgf8+gLx71/ajAH0/47iUFgB
0jmIdoXZTeR/dancld1OiY8s9yXRd7w8Uy6sjOjD1GOXHmcZO0pPbUH2S0mzMkvmE5MAZ4pLz2nt
xnKaYJ9NIdk9rcB9vzbXITtg79wKaVADXZrg9uVo4M/2A0Y2BkzgYFicm+BMlzkIZK2cmbAcTNQC
Sa1/5BTCGkMvzs2zFOdi2aWAx89dG8ZP83vOXxLdyLxO0rlEnGP6SCRf9bLM22D1zZ/VKXbuAMen
IrQuo8qVbDBwFvYEnahrVrrl2VEElRJeOedleU5D5xt/n81aJEj6z5os5RwOgsKx/5DntbpuC0gY
wqnU7CCBqi+k9QoOb9mrXs8SIES+/GgZOdQy6tYreWHfqtIINDYz658C38QW5R/HP6XJtn1S+YjA
y8QmaCyASgPfFOI3AFW4afSxeAXU+/0MLQX/Lz5D+6W/7WGqQnh7/COtjAeTbzV1zJchkgpp58jk
gPjC31ieqCOeZ9Vgbcer+RArQ9PQQCw+h7RACxDemY8YxgwpQtAN3Ef3+fsAyTxYTABjOnaMnWiz
B5eAiHod4hoXr25y4I714npVETTP+mJrHG8+5zk41EKMVYUytvAk9zqGhjoyzbOZv5kjVlK/j5/D
TkLyO6D3UO7V40yfc2D6WldUWhvHTtJf+UI6vmcj3vbx+vrLPYpbiWUYU5Dk1QrNI6+Y24M2xpwg
CJLq+f7viUPEQs2HsaoMXrq8VNrYgduJrTq47nrIV+eG3Fw7Gu4k7xGi9ewoIFCznvK/jLavGdPN
9gSs43ekQAA+qia+hNBCCv5VrBEPQWJM0oBNPwPaUx+8fh65/WSPXobatEw4s8Xs/JAC9zv/nA6H
iYcf6Sj+CTLwYR9tf9wTgA2ifp2fjlPAMWRJcRidVIFaAd1W77ZcyJbzIwl8jrMztlHXGspYMnEz
Ab1mIZ2Of+ns6VSReF6Z1wXVSEKRALWKnHNn0xFWmm5t4YDe07n4e4xj/+9M+xXHnTljWsUEtOO8
nmWIQpE9/fyjNDBBzSx7KUMNXUhmolexydH7cFCWfdmiDuxpqhScsPXSsRBoyxfcazP9E2X9vdPq
JbNO4Vd7X85NaTb5Nt9LKfwcL7m8JwvjRFBmJ1XQUGbD/MRQa7wfuw5foud4DGzNfF17tFoLyNqB
/OgTosEeds10LJ9c8Gv9lf0+hZcXUT23qJEPyUOJNu4Sh8va0rb+JXpGiJy7lrvLS8DXInx64OLM
hOBRdGtbzwvNIpJruixdxwUFEwofVfaQBr5xCIEn0C0WR9KX/jYDlq3C2VBV7EyPKIp6tbSfeR3g
ies22ve3nD82r+IldAZLg1mwVsfbHkG3+gVeLSB+e41CpSZFWKogjmaEJu2+zeZ374zZbkRk1thm
H+C4TqpnHkueCue1Fk05u9KmQplrhfimQGQqBCw2k+CJ2H/R510ahf1HwRYfstAQfSUvchVS6bZP
Y8waMcxZ3Iag/8mBN4gZa+VH1i2PsSmOArJTgLvde1KgZSuK5jCEpV2Esam1EjHjzlQ6J4pVZDNb
JPxFe34OlnPNMcpy6QiJ93IwPQO7OPs6DX4DTDCgdtZkodXRVKZqCYuxKT2YEl+iVRMVyoVbQcSH
m8Swg69JmZUYRoaPNHX2w3WzPiV6ee0uxl8WpUGseeBYlHEPnxgi0k8vIjy8Pul6pGIfhydPzjTz
08qsY+RU66tb0nnHXnCnJypw2Tx8vKNtVX972htFYuMNVmazlZJe/j7HN4c5sCv/1QgGKijUoHYZ
Up9R12iuMaWP7u5oWzeFE0XlfWBHj6kTFRo/oSHsGdQfloCZFivuCqzqFzwUoIdTcdiv1Uh4O0uT
wck5bty/QoUCR/WnySDnL1jZcG1K5xuj7QmL6v2bZXFaKGZjiNh+6FT2d54e5HJRWQ12PPxkxYWF
WFet28XRGtqy0QuRHl3Q8P5OunDNb1V9E68SQz7YSJxpMMoxlv1ItyFizBFIdEmE/r9U8sPuqz2+
Z6ogqDkTJ2iP9tR0EwRoO/MjlDJ1wvMd6pX8vm8eR//ovFFD7PmKjwTitUfSYBWhAKK+HGKFOgDt
HDnvg5AxPt7Ksb55MetkNAvIFGFvXelHJVcoWylOId/OkbXgcMcEruamLhhoAFj02bOOlCEroeqO
tNhdwCQAJA6Ci+E9OIrVqNMsKvNyGs+sh3pyWNHg6b7yWAIh+LeQKLXGoglz0IYKUDGlZ1uH/UAx
2mRMGiHb0jyfbNJEGAU8phyph7AG5VbpUa124rQ+ZshQrhoKpsi37y4NyR0tTJE4UBFm3wFVoRcH
QH5piRCFH58uhowtzLeCy2NJhOD03nPbZ8feM9lMnMnkTNfd+wK9eSiCvks8jJagmn37dpxLOIkc
fbMGT6rnBMHqoXRy9SxtJduYj6ie29m5CNzk4cKTFn5tlLwk7oJ/yVejeFdLWVSCD5t2egHr39CB
7PSyr1hx9EMNtCEw4AJ5b9wD1EReZtewR+tk/54b8uLT/v6iqR7/0kLKNhm3eivJUBxJ18phYtx2
OarfJ7+ijfbY5KAJfrd2CZeLaOye7RL+LR+0nCMVCaxMhEeRes7Ts4N/J4lDHc8kSe0+o00VgORG
KaJ2nDdjYAOZWJvJupKYliZ9SnAceSXhOfmm+/vsS1/aAlYb895reUWxqa5OC51roC+7ZCmppWaM
fpCIeWaBdozqO17+jZZgVvqfFuvuw32gJTDgCvP/7HZh2XiX56rErG3sS1nQuobNpiAr3c92slTS
9QgEclSydBZhfECv5yt0530TUS3p5mEoaiqWMamcAYYHddviGfPo1qRamNvZ9odGgJZItI+ht/gM
Q9BOyEUjX6HcDv+Qyj1EaMCGm6kZ9C0kolRTgyimWnVlO6Y6OtJxvFbDJeQO/SX/UMCGMfzOREVK
j1R5E1l6DmnQTdYkBYorHfZ9KZaAMmQsZxpUQrKdHsJwAiED8VvcDKhBMy/ch9FO7mliCtotMqxK
XdSu4nOvTQwejusxUV8r+OmBGMZm3s+fbtTmSNuFtxdhj1SqKZlWYASNvo2ejhyeNmfOkGG+vHJP
gISaPof/Uz8iccVAUGUZixuPtCZiqRs6ziOPisTdaTaChM2SWG9rrSj90qGHIRoQJk27PPmeYjIQ
s0ldbXsOstsJoa2kTeTKhJjlqnWtNkpkOmsa22Q1yNfXzA/aBFYVHfHS0j3hFeGvQhicgfuzpT2J
EriNMh9TVlzTJ/gWDi28nAwYf7q55dLzeWU25LnSt6l/dvcw9MsPmiSRtVIcZ90BnID4KgbbsBTS
84KxqiEteS0mfvrrF4GaXIhWydv/6JVsrnHydIuN/4McXVgxVOjQYgoDMA01Rh7cUnWSo10UWVZ4
4XUqStkPs4PvLh+oUSqCUmXExbVmKfQh7bskcc/2ph0zL+F9rw7n4+9oK8Jf7lnqWL2ED6OU+iAk
gjQ6zaW52Bcey5sdsLcG4MGbFciAkLXWfCU5pANVryWO9hupbkoQHcDplqaHkBHG40UvHKls2otn
fb5hp6lJeTstjSwTW1qQw9bIc8DUYMwXY1kTgKOil7OjEuqKEM/pKlFfKv1GFPkCsUWSW2c7PXBk
kCM9T7N2QEv16qc5cQxqBGU727Hh7azX2+c5dbxr6sXDZoiTMoI474ZNAyAAILAROoq1dn/JOd7d
0T9ywovbt0GctZq+UoYzaB1mGNEDosrxYQ1yR5V+DwlW+v193RXj3VDMuqEz/ZF8DizpQGyz/oEP
GNm70+eec3JetLttmuILu0IDVC/SttRUU5kzvk2d82VlHn0LfmsYQw78/zjciHf7FugoHN45SZEV
aWQbmoZt0kG3N/4F2eUaPiX9600U7q6AhlyYIubBnHEIfjmA7eaw2i5HOZs/b2M7ORJGJx4S0bea
TtZ5fD38pK7/lJhNhCD7OV7oY0kGmMkd1dtPh6IH8WFK7+gsfIkiiA/Qpd00Q9GouCIa4b2PoU+h
M6Bz43cm0w2qOrPhuQDVzn9+XLpxFWLH7FFxkJexAoJ45wMNpVqVAUC6x/DNUeN3vL+D4mI2LhRr
xVKXKYx8ShRB0FWYNMf7JrlE7dfVWl1KHWXzBXsiFXXBZeQxFnTYeWYgdBWaX1/RsT73bZi6aFhc
wpoX56jnj5ixfOvd9rz25+JVwuR4HW38h2FkCtyhKT+uCd4N+ktSI5/0XdquvXVARrKIU4mQ1q1G
NJwKsuuKvJmb6PeDHopom1LRFaplQD5yKwqC+Ljf61/VZbNAY2NVd56YBWaOE5gzXcNymdoAgUws
5viKUUqFk0dV+quG8ZUF6UPDciws66s0FKiUF+L3/USAsz6eseUtNGEoEfjBhJCkh7dK7GcH7Bd2
6C7o7f/BgWLNzlKSucL1DS3/bTnoeVO6nwWyn+sN0jLrEHsJ2tF+aZej3u4h/yzvUUrnV0m+enQj
cCnCaqdcLwKl/wF1FpujtDCfFA2HP8DFwi1jwyInLtWlbpvBl08Yi59NX1IYg1Q3Dt7nCpfISzYq
zZH07VrCbV1zfv39xV+DcilwkrJ9fYW84DxoZvzmOMGCPOBKo0D5PxKQ6pvJjKWpy100z3qRMD1P
BHAe8yFlFeImNYSX8iLlC67bIkvGA4ac3bUeL/RoojGVmkMrrJ7OXzagBM12zCCCG/DKwqtYdhOt
/hv9QfapYzlv5bqmbn4qlFQa9sa/ekhh/NyS+SEDJVmXKyGjZ5DGbbQ6vOeUZE8CuvITcjYh73/4
yDUjoyfWK8fCzKAQlwiBksQPJB0AHjGo9tzg2ysZ7lzm0v9QIa5JO3gyEOz6eZP2Mmdl11V+wclP
s5qhODO8JxTIFvFG65Kibds3jYlGIBFg33l/WhVBcOO6RMezlBdwh0G4nLvzy8TfIcTXKzulryWJ
pwCtZvUvwyuE5+U7P08bC8Sjhb6FnrE7Jo90o7acokq+kkKhdzz0jBB7gKdlfjDVa4Tt1LMgX5wj
u34sr4TWyeVPmEK/Yoz04SeRnGflHy0rj9sj3KJgJRWiiK8PpHvIofXuUsuM+Al/QalLkjkvAR+H
lceBXI0mqzii6LcjTmcIKEDflOV+eQECsOMK2EbtTYdu9MjmpqJr9jSqf38hh6V3uEwmZ5cEHrFh
HhqL9GlYk0AVL0WsMf4JehST26omeLBmYZDJ3vdHoJS7YiJ+F99NMMs6ohDtYcVD6ZRyv2ibyWN7
+EqyBYwI95xzv81J7IBv41tmilOZ+nO2h473TffG0xprkToWFrRCz9L0JMMOXfrUuSlFAfD002fG
psLNRpvrXwV9IsZSLGDG3LLPqZtS5sSXd8EV7Kl26sTIn6cl6jt0NZn7STgANWY8a+hPiYHoVTCi
sTihv57i43JT3hCJzPX9LID725WaUvyqdhG59prCKzhUOB0XtuimFPR3QGi1mxDt4IpBPe2D1nec
PFhOg8Fpz07XSb9rm0glEvUZ+aNegc4RabwscByB04gNPuhXBURjtIfQD7Y4/EjFLj8ncy1Xn6O2
OQaQ405zTzPhr+1EyHOGqwpBB1LX/VtQ3YTBBddraGD0ZLFgHRVQrV8U6QpioDdhEsP9Bk9fdZ5g
W+7S/CHKl0A0M0WTVT0FcyeXUFNqk3ZI459oOMN8VCoMnfc4NwXQHKmfRxIqAxTi/nU3YwCTpcvL
jHfpF1fWmjesXzWwMqS0g2FaTUDxX5ipAnK4m2EiQlUaWmF+BgNpAjKvedJTwy25BiA7wDBgocRC
GEZQ5gIQxswOUqL49oV0wCP2LXWidr1YkqNtyDGSq5UUyufqdLJOJjPjvX1/vYy9Fh4XVXq0K/Yp
YMaST9yPhB6f55jC8rWvPUI9YM2n0w1tCmnVwAM1HFdvNQcviJpHEflcjWICIv4Gjvl3frBVyreO
iUhfXgtSJXo0l2draCfQCDIuvDt8iwiC9QC/CcuyrAOiQIYWu7b7wzRMhmLIHJYg2IkHkkcUcqDx
maxL/0HI8Jb/iuz4Yf36O+TYj0VonheEvLmCGyEU7TEKdE3DldXkjVKO8Z83HjnoztfVGZjBfjyN
gB05e7E29Tmpf001NlMzAV9Jf4UWEqjMKx/8pcQ3+EY+XOeDFaYgvwla/SHP+CDP1JBrUbWOmAB+
VeW3bqDRGXXitpIerico+RaiJubd9Z2Pmd9drdEjL2hLYsDbkgxGUk5DlVDBn3Hy02JsAOiUBE8A
Whvfp0xLBx7Bs6yZc/M1wdGrwqX8nLSqmhfyL/FK5FsYX3y+w6fLoVumdlTE/yqgbu1DxSnAwnIi
Yc0fIdZ4qBMu8Eylv8cJ/WCGVI3JRz1SsWiq6cJHFbj6tP2hPhypwGtLaizuBNywDy8H/zvNSKLs
2DFe2hjovuLh82VxX/2N5oRUVtl7Wmz8PLAGQxV0V/LGFvqUUpXR24ArINGRABpx8LiODN7Hvafe
a4eH0gb0VG/iyHFxWnUnewg0miTPBMDW0fgPz4YuAlvwfd2dKx8RWMj7H4IdSKmHPkl6vmFUVCDR
XYiXm8wSYlFmuzYfsnBSc+zwuBwlyDvwa+hTT17vab6gXOw1HUimELy8K08eGM+KOP330ZuU6o9y
pfYJDajWYHUOp0leadZfoZoG+CFK6G0/utTFTpt+ai0RwJKcAd1fVVJShInYJwG7XtCCDipqn+zQ
rt6KYJ5bJXe4tXhi1Ubk3Rs9ywhbfSF+T+B8s3Igvs62i19k/ZMFKoWZLFXw9Z6h4oFmS24Q670J
3yDBv200owGDJF/DSvUnBuEltrO/ozqIydAQXASvfolP9fydryNMtr+1fAO+yDUt0yIe/uR8O41S
xLOHirvpptTDX6Y/IdUdkVvDaYU7TCLenYWmZ4ePsQYn9i/1orxYaVyP1taxbAXYsB5jyzIGbgCf
G3NbNbzjz3djhc2lnPdoNlkTWh/KBrwCgRXHxTXsusrY24G4WbbMEzFA7mU82E+kGlQ+p4jp8F2H
9/5EPZYfnIfg/g6Q5pUrFBtKmEdjlgHL+6O9e6K/WnbXGVshIxSzQWxpqKSxRTTgeDZg2g8LZw+T
g9FSK30Xk8lPS/MLu5lkrbKeqkmyCyTf5lwmkhGvX0c1SbE/V22Kh3Rx6znO62N1Osxi2gQN3GNh
y5FmLJKrYVQwYcFOalD/KytZOMwh7We+ne9F8d1uqVD4/R28/Jqy4bx+XF7G4JDG/pAoBbGFCtC9
maA3FFTADdbyfLRCV7qCqzlYiJMGk97l1xsqy/zN8bQeisi/74UTG6P0EPj/+jnZXc7smeSVI9p0
oa42N/I1TVV4xgugAqjyVuJIP++Uk+vGPvVToIFSRasAJIT6NlQVuwqZ2/qkuT0gQKYjK6XifT/I
Y1+x8uTMTQ5I9/+MVYNE4bRs0O6eJH0+5ihGe7CzO2ra/rDOxUaokiIzIQgCvxqjEIGuVXAx0QXP
f8VBuWhmgaG2wqc/vXkpHCCrqHAUV2mlq+wPj0LdMT8L5Fv5u95BtMdHxNgRcSHgY1vnFtmsEjiI
SxhFkPDQxyEuh8dwIqfLCzOrs2D8i1rmREDdVntkiNhpSQbwBXTUmqrN1Fe5GAzKB765wXPLSi1L
ic9lTWuh+tvgwiYoGAAR3QpxHoerAk60v7zMXID3+FV2tzBySV1BKLXzZvaJ0j21CS6jgI+NTKDH
n8Yau8Ljs/SwvqdErSoqlzJ5/KvL4piAhaICH6foxy919n16gF5pHJ5aSBmoJ1EqucpVHucXSTNR
gQLMReuSRTyumG9rMh8ljeC0rLvoRyFSlJ6tMD/oRAeOIZLD2hjHasZsk08euZW2XkvgGAIpUvV6
LQpxD3LGZdPWijiXukX3dmut4TqBP+bS3HDJdyiRjLaN1tCk0P2NmLaUV1vFVwGNhpZyrca/MInn
AINtehm2kNFngy+2p58TDWn0W+XAJ20Q6GR5uxV6OXJR7NovYLK/TsWL3GS3jZcuowFmoND8VMfw
Wyzu6KjTqlSGE7xLS1qAnE0R7W5J24v7oUHvmf0pGtiz/OYS5ABuA5hSROw1s09r97qafRvvl5bs
Nq2CPCMhJXvY0qnz4joebEGwNZyFugYYIFqIwTqM906vhyR5n0Der8d+nDeP0p0JypDYL/hMhltu
lcL10wc4EA/xFIdROwGluEymFwB9+D6NGmpccanzf/5AWLuDNoyJiVnaHcrnHxHXIOkO/y4rC1/b
5LHKC/DcpeG4HGh9pl4VEwS++bsrAGzjdqAf+g2uoIBCrkk2HLbSmhEKji6wY0tcXtJBV9BgWfxA
fwnALpC8qhPHQoIwvODlTzG88qHsNwfTvSvPJH6n9OemTU6A+M5cAzzv2WxY9BqOMiCusxNedxl0
TJ8d29fEgNl+lpsXYEgzDtEKzm6XVm3KR7OyInPjfwpJezsqfZiqHhBSLZXkxuyG0I7/pRiz6QHP
gUDpcvKV/E8tdZovrpq8XTVTJAeph3M3RepHUsMVFZp+DBahGW7GxINfihbVldfWDSqrMhs3mqZ0
VAK80QxtJrZ6/v+H3Tlfj+Bp1tcRb96epcQfPFWfKzKzSXdesmC7PKsfROyvFkiNR5YGg1somHgV
pDEaOYElGTX+CJGa31BZPGwN8LEGG5AR8wz9AwBi/U24NERBhgo4cJIP/2hcv2p7fqP3aQ8z7XLL
i76KWcDgladT8qlCrLYbuvuHDo8gNuClRVxlgj+1XXl8o4qbt9y5cWcrjLMhETBNHYZZ2OoT+m61
lcGtjgipcJ+f2+isA2ov1jRL6CJjnedprfT77IfL09WOcQAuk/nr0f9NUX4e74gFKjZSXnTdb2hX
vaT5CrWSqQEhnYsow9vOnzg1lmiE58kimIrorvbL8kxteeyYSDW1fQomEWmhyHtPOIQT3v/0BCgl
zLL6G5kX8UdGqJxZN85ituoVJ5U89U/CLXPAMQ1bctp9kz58//AU9eMNi8t8udBJB8ItA5S2GCvn
/W8/Aw4Tr4ribjGR5rHZZopHcfam5GkOjW3DnFyjAalJErpN4S9rtr6EKWwx/jlMkvTtseOf7jX1
CXT9TaxPA3Gz2e238ulIS3xde2gxBMqD60DeXcZZ4IlLmd3GN+CYM2RzGY/ejKmw9qLPtg5a/+HG
LRYyIil79o8igS2g2ugmcgxDCK3oT0UkMvO2nSz9Lk3ODDoumr660Wr2ggJwjdoUYgxAiKGrBROz
E7504v8uT6zSZIrgN0ZOEnmt/J82zI9720jo+WTERBpFSP9HpYjfmkcloau7MSnlevW0WhiuV4j2
W+ItaQIS1ccMUONGgjJD16rKAh02PcR81grzP7NKmICI90bTlGQ+/oEnZnRYnfsGAwS66OaIiqdU
+CBEqw0iLltc9fIUJh14+fJcHNeTbZZ+B9SUcDipu9YRD6+EOE/aCAbtE35TcNWMrdsQM0DavJay
lskPofumyl7z8CpfnKB7z7bZMLheMqmgM42qpT4DxC/5B0EN9I5gLMljJhKch/+USsm/kmYq5660
GnH2tvea41W9pc/vFwJF28Yka9Jfd/F88+aBy8dWCpb9T6v+jvJ5Mcq8kCmPWlZDN7lq1qcO2YEt
e8m5xasq/jHdn+u99hoTwqf7huFosOLX0eYkSiox+KLRe8MHZD/8QJB8k/q91KFswFY+KcdtGKvw
RkSEUmxsElO+zsL3YD8Ag/t+xUAlOLBoV4LpTFmo9yx8q35k8ligBPJw04k7BFTjU0nbK6nZdug9
EDGMINmtorcOlfu/tVH/J4QW4o4ei9TZFUORZq9JfZkvXCDt2ISwFWOCfRHpIft4SVipjWBUptkt
vxjP+hRMY0k4M7cR4V+M1xXpmOSZCqnPzg16ZPihnQsJhYLqCaJgVa0YuFxwLkM+7uaudaagLWIC
ajnOthrvWzWxHA1f2bs26AdGo7WVCpoTmBT+EkNuWDD0qCIhbszSm12Qp2YyR1+15eNNhxd4mw3E
4+j+XskGLFb0UlGMSfegHTNZrNnkDx0z2LS1pxVHIN1Ezoz2htwRrAMmnIQ2F23hThX6RKBbMgJ+
Uizojw9Eo/42RpBwOnfRXgfI/GBr11libaWvKTOlHCZxte/HdedRRyiEqQProfR3yacwE36M/vor
5cnZTXerB/OAuJ2ImWXw1mIwNS21GAQVPmzErluvBudbPcPuyYfaiKzMPcUBMFGQFBaSgMc1ae0N
OwMYZQWJqD1WA1kgw/VcyJE9cbB+0yPMIZqzsI3VMZFBcAr1gEOUH3RwTsB6kZfKHxxRdI5O68KI
BQgtDTZLjokk4Gm4lnRK46CeTbXr6J+c747Dt4HXgXVwCwoExYTJzG4tUuWLtxAZIfxwRYAm4HhK
14biiXOr0ENsuaqDN69wnR/n87OsEoSu5Q2BEAGS0G7bBDvYtHZvOzZ4sBfR0tZtRjNMc4hv7//N
dRkZPDI9c1JKDAsLi9g9v1fQqg932KAkMzyXGM0x7mZxfAEJqNorz845t6PMgP4IGjeVBzji71WE
dRarvobsM7qLlrlogiXyVYn+CwI16jylsCrqvygY695ywglJX8TtcBRh8AszR5pG9YHHIKMQe3Yl
w+dOy7aOYkvD5SOL7ydSXq6Pu8vLzY/HrxjKjy/vCPGtbvmB8B/d0jj9xKi8utV/ag5KybR/SJnj
koQzriM2EXnD2UWcMh4ZFjGVHxaNLNq/x9fxi34NaJq+PqvCAbPqBjANmvYBNDyQDmWtyQj4YZEU
yk+ByrfryKJ1a3a6yMzL2TxFAQJ8LTiPDGPwVe0vJzAGcpHmBsQHZDgD6sas6wdZLnCrtxJZJlAR
tslkuV8PMoPTMK2Ln9wtXfqJg/Y8m8O6pxC2vGn0tzS65wevF5vhjmWVYBS4nxkGd5u3iZEUMFvP
xzCWzm866Vaz80JqrrvIF5CiyZnbr+SKR+x3ky6ZC5GWoCXIh4cDfec1p1a+1fc0WfT7aw0hfo6O
8lACMdl/tSe4WBRjCbWgH4XbGJE57psPIgxYGOmaSs66uqu3lrAbOGIx9ZawclHq4mfyG2aytng5
NE5QJvKJ3Jtfl6BD+Wfhho5FvBydLXB5OKgQllviw+aY0UscX6tZH8aFNYa/uPM2NSELrY/Dt/2H
kkKq3XzQfVHUw0d+ArVa6KH1VPIyAV/AWM95VZ35bFw/o7SjjeLgAmmZJ5JUVc3QYkWVdG5UtOsp
JhJPf6R0ikGGN9sf3qy283sxKLAwMxqWBj+e+21n+CAqmoBrZk/5xYVlM8BZ3kztfMoj91uezO+J
6q/FmDolXb0pM4qqOogVpsxxcJu5wF3lZiAWpn1RfpC1qftoQgQ2W0iEhrZS/+EL1EiGl5ZOhETd
ZUg9e2WO/3JPWlF0BwVzJ2JwcS288igOtK/4OsQSfpYd/amGUlOYfzIVXYVavDXQgZGeME3PtumU
Cnu+m8CMgOZ8i3KyuG1OK8qckghAzD1k6Hcz/366iUkLxQ/f4654zw5ddu76liqtbjQ8bqUdL858
m7HmvNwx7WRxWqgy1yHJjpyA51k5yvd4K+Gcia4+bSqtjmh3jADs5b1OW6lLx5u4kOazOiqZzOdT
y9zI1P0y04vE/sHTqVnIc2U61NOiaV1VI7tPAkypr3WSmeBGY40n6dYq743uNMGweaa/PK2Dfsid
5ptwcreut+HtAIS3Vu5+rXmQdYiPRaznik6QqbwxOOKm42HLeAzq2EQxZd7i/PoESF7cZpF7MzZG
CpLXxj0Fkfw0UZdXx8JiJmxX58w83k2SOdUOdodl4N6avoqz6GZWOPapc9Q6BdsrPT/0XunG8tla
+gMWTkzdvvSsxJd8D2nBpTB4qO+XVG/bHfvXUEAhg8ngq0spTX8ow1OPqjJOWh2XiTAt9voo1Vvj
+Hp98MvYTipFcqt/7ixABFZo4OELRBO1ni5lKOWp6q6AMtAs/+BEAYN+wld7H4QOOOEIZSRUeD/P
HeRhSvMJ/4nBtfKc8RbgykGILXJlDOP0jhRwAzmHjSopSo+tDdnuv+N51QGDM+ARAeEOzLOJg9AH
XwxDYdWt7Km27p4zq3+K2LM91u7vgtFDf58sTF3VUIN68i+tvxlqrcj+rhAkYC8Sm6qZANU3axsW
U6IlqWu67RrnBEt8/N/YnsMKR5Daod1s+A22cj2pYcSI1jUSzgup85lZAHXwOwUDn1OAqsxXuEqm
8wEKatZISSCSTa+tr6UO7hCLT7bFO5PutufB38W7JXIU3u9q9iUqAUi5sxJXMtV1L2y7wzug2Q2d
I5AcLDa9+RlQgLcad4v5YH0NZ0hQ6RrDkjvlX4RrzXOrCF0JY2nOqcvkJUk3PGsbABOohZkiUK3t
KSV4J4HWffiR2k3bzgMAYYqy5vs6bVsYmBcR9V7//oWVZMLhBFz4eAxr9VpRIWZ8Bw97ySVfboYW
d5coJm2NLy62aAiczF1t/ahA+0Um8QoRkszlXHsb6EKFMxEA2v9sAdbTH/OasH+nvPWCddWmqoz/
UP9Tvfjw6cguPAuJj3L6aMH2MGW816+ebCEvjZzGQi0XGUE5x1g+JjFIZ05Hi4u5teXDXcTgYELa
rWe1Ey2yjwsVoHt65x4Cel86hOoj4fDFqlpk+Z2gqbJPNbH+IMij+kcmTeiC1QOut6tsNDk9OBXz
4hYRtIz55e7abZWhov3/Zid3bsYoh/AUnU3TU09wM4hSBvn2cDs0BIeOoQnM6nK5EKEBWlMLj0He
ni9hC+HYppTbagAdPuXLg3bW0YByfTEd9QMyQ1kUVDB+jspl1jhR1uFdKtTGg6K1XRawYnUMNAOE
/6o6ZaW6L9qBvfRpfYijacXJ6xOR36PvKI1Ou8CxVuEJn7XF3U9LUeKzWcpAeR7vKwE3MrH5nqeg
dQ4dhm+QjfYKkZdq9t6BB6dzoQKRTqjYJ0y2pCS/P+rxwaFGFHetHsfgTpd4wo1w4KC+50ID9DLO
WJImXwVJm00YP9hm6pIvpHndJ8Lo/p+Mfdl2nDKuXmaueR7/afMypvlpkOvP1AQL48Fz4cKo4rZu
n+398IWHEbZJPgPPDI9J4wmCkUOShFS0qEY4k3NyFHxe079Zk1JiUvvLZiXRJsZgkjmcmxRbQAIj
NYkQB9dxJ2CU4CoEwSRF0nfuR12Ele8OQxo1k+jaahVDd7XdDayJ9Oc8wqWP/IOHsPDFwSjfthjk
a/hv6G+prqmdxnEyHxxejmCr6cFATemeew+lr2Y7VhVnz5TVgTzZd3WLd6CPrUUVeu2zlfCJ9Lp6
VlLMuanQLTyPS0yAiZ/Jj0KObv5SnHET4ozS4X+e3ja9FPrTvq6SGSrSws2D+cycOC3qQ6PHMeAS
80epUOUx5NdW8vBxHdDgn0/TrzEUU/Awu3egbkdly29Zwbpb4fbwGQWeRcI+tvvwJaHvXdfV/MCp
6XkbVDuf6i6t+j3tNNRF2kik2nB3AKRyoQunClKPQzAQ8MUl2qQNMC4uzoWDJkaThUXWE6MvifVT
ukOXtreNF6dddIw69+iT2Z4BCv0smxPPEcvQnGxq+CIrduVDPgwsNsm6XuSITaRwsM1rfMacz9Jm
CPlxVOKfeo45V8K7gL3FzfJHQXuwOdg7ovCYOB2Em95uJDahvoG7qtPIxPKt28GHSVtqBZ76Xp5J
k9q/qPawlajEXP7h1razwwN/Jpo0inK4z6v9ekBdxF27/T8A/93y2AmzxjQc7DTvHjyAez1iDg8A
5/APb+ioYEET63lOLDHz888Sk6PvbWvuWSaVWTlW0lq4krUR1fLqYe19MQkKWngvir0ZG2cvBFuK
o6c3UnLlLnrCxI9sXmmgz9wVaOm7Xy47eKTk8PAjgM7XY+XrEeCCVdpAb3+F3Ii60p0mq8IAJJds
t6SOg5NgYnbIxAbX5Ov3/JY8kVPi1/l9K/Pr/Ey04uAu+W+j4V7Ylvz1V4/JlHh7pm03OJN+WVfL
J41wlcRZg1JKScSGW4m6fuw8q1UJMoKOIR3nKVYJAa9VvneM4lLfYsjdV1zdh5nPldzIGvMNZDbN
ksYQY7pd37gW7RxqjB0WJQuGdalVEKqsU8/hJL1qA5HVWPWzWINI1GX14D94lP6OeGLVAo+2ju75
W1ncScLJHtoMsz8R118KocQLj3SNGjZqWdVbAg68n1UrkUox/eFI3rNLuP0wCkswtUBABT2vDSda
m349VnHPdaWVZXbzLzsUVBwld+9VQqF94Jcb/ys+t6ybbIVOJiyWjwUl5dcPFxXHNKPucV5lkeHX
kIb32Fuzk1HJ+2rphBoG6eGGbl/w9RyCYMfmLrzlV7KTmCbZrC6KiGy5OeJkXoVt01xSkb+LwHNb
JiqdUKEcHlBh1k65pNon/SnJdsu2Li8GTDdIy2CTlNH23XoAj8+pAibeEZ8+iO9DnjxDVBspDD7b
FqP/uxRvEdwxVEMAzJfrvxn2Z+FPQ2qjRl0UHBG0e7+sMjg4iRmyoOJZkh7Y6pgA/nDmSWLOPKt2
e9f/2y8WEvaCfEqVnEcCoSD/lbjmBTdoy6uFL/0ssPfIUn56Df7eeIeh+63rCALFwcDztD7o+XLo
ECFQSZTXVaRC/dcfRXpc2EERCUi3H1ogvHjwAGf7uuT0b40fkjw9vKO2gOpJg7DLk22NnqrdRk0k
fzoGRoaVbaKj5Lky+jfjwXSA/ZyhNxSpGHGxtJwePAFZ48t0CDywg61aeN0aBWFND16SxSGva/Av
FdzBrj+98HGWR/8DdaRvBDN30XLuUzIB+6hWhorDSZE8YrAQ+ciGVDL1NKpGt/twb8DUDqNQXumJ
vHBYUoVGWN1ePXb43228Qdp5xgs/d97SxWwGJp0Wtgtpsg7lIwgrH5FgPC3utWtMLMr2qz+h7rbP
v5mxo8zQ+ZTXCcMfV/vEGzPRK970AnqMRHFS+YE5+bXYai4gaMvZCWhXtK54SHjkMHBVpwdhFnDH
n4xkHndhoNJpbprGxQHBeu7Cx9mLl57HuYbMpD/EG66vT6QZi5rt/v33W5tSf02YNBFGO9AoWsMx
nTg11y7NYMYecedisCuK7eFd1tJR4cLDDuYYo8XqXTWImRrd1jHeaymHU/0sGT8VBTB2KEUavLKG
b3CAvg8/6/yC3+sTpyWadvWxmvQSYefyoBuXJrDJbk4qg/0m7lcJbDNcw+7OfA3yeiQE2FZEMXPu
ZPW+ljzyIjSeUyqjuDNv+KYsaCvplmp2Vo2pvnrrcBz9t988lbPz6/ybvZAi/rl4Cfgt0Kyw6GuH
tx6HYq6tGUYDGmX+HfYUQZzZGIOxRLzab87fkPl/rRbHK3K/bn8AYg66O/rFitbjwZLJiarFrIVb
rbawbxwoAW5zU9Ge6fgx1Jz+SlsiivKQcP45gmY9eHfFSAzsjBFGDBXL83JzwtDFEosTbIlz/0Rt
f5te+7N6JZGNchkPAt/kUM+s8RyA/g/ie4a+vAP4oTRLPNSscD8KXA29lj9YtuG2w92r5BdnusgZ
koVk3JrnozGeW7D7YrWjkWIWzU+Ib9rt1TTt6TKtIQb/SW2Rc4dMq0CeWREH7gO5PTzkR/UjOnwt
oxeiE6GJrFh/Ex8+sE8JV+E4LydJVO9cowZkY+64r6JjfXi1wbGdwRtnVW5kr4Wnt+MYfG6ie6Ti
oQeKU14b5XYiXDuEATmmvBprI99MDOOW3lCf/DDhST3/T3AIDAj83HYG2NqoloczPmEdThjtFngU
yAEJ1MqA24nQA3RKOaZYKU7Jt3h6ETWly/bFG3e3oln7H9X/YHaSmSTRlLMpU4/GRgzewM3x9otB
FsZVPhf9jn5vimm0JA3gkRfGedudRjlU9jjDZWRL1FdOskF1396hUN7nEgX5D5cWeGOrxLuWA4Uy
T2086PtobUU1xwqGbkdo2oBzC+q14aCdag2AUuykkoMz3wkWiPRXKBnEPGwI+eCUxC0zYvfHLpir
wDG7Yi7VGM0LK6sp/FlGWATNii7g8MniuZGWaI1BKH0Akgf5Cyrlbds0TvEjv1VQ5AleDQFDUe5E
JD6Cp8z+1lrpz37S0KALpgVbvoQk1j9MWdcHxZBkcl/1hLFw087fjWPsoSmgrQwAGW0NGQ3d/Rpc
Fe5jKmRs7RB1WMCbw/o5o22vApF8vyhEtzqx1n/be+U4/FDSDQrhjdMTOXYEyxcXLg1slwnAUhLt
aUDhQd7b4BEhiObJsi+JoXOZkVXojDkwTpSMSlIAg96Br1U2Dw+WKYMGdFIxuU6XhapZut5I4mMh
KS1t8zluRANMBLmuwl3beUpNipx0gttPau66ZHez8t1mf/lYwfQcK/yZT5HJ0bpKUp36LXwdxRv7
F2u02KtW0yJO6H110xTo5Hfx5ztE22g64iDXR70Dqu7doYad6QCQQ+ZrpTNJfy8lgudgCrocKOVA
MKEjCvUxA7Qc9iPxOXCbWCeF/+ovHXWYf5Z0MNOyIX5Izp02MFRj3Uc451k4cfRsKPt7+hqVNPiX
D7IGpGL5p6VpXZtIJCcX+CxuniD5YsDjs1S6gxVphGanl9PBYQ9MUca8sdD8BsxcSnly6Nk8cOZt
v3seS4uMWeYfnaxkxLk4UjU4uupI/1GEcVd3bIewzfZoEuHXIohrpPtsffLMAb2aG+0o0ICNsacT
HbxRG0c1rWwWZyjTo/f5j3wOdD7F4/OOn37b9di4/0f/Iu0KPaJRWLPLoFiLbNI9e32GHHIKpmmo
Z3R1zDUhd0gpzb5H8fszBEKhX6/HzP8UP6Tp1xtQxPyBGJgptyzTOgjcelm8Wcy/BXXiRhSWc8W6
67CFUKVULiwZqjwcwHCMvBK7g7v02ti8Hn2vuTfvIlCfUwDzOS4KOsq3FmWdNZ7HE5jl565aSgmS
Uk9IWCCjzHD8B32i1R0E60FVCHFbbVszq1vgRZn0ii9nTMiWx/rh8Y4vS8zV0hFum2ukTKmEatYG
WWsX6Bch7zeweCPQNgMFdcxl7PDlCBnfcdkCVEerK5O/bxU/eHOMLziFPVLuHXNbm+QzVAIYj2Jc
rpAdSVdTZ3qiYwelcIH49XjyVW1W7FOi+h7lKKhw19lhsZWdL/cKpVBsVesHR1Doo0u6p8+SXgHk
ryyIicoXcfGyxU0yY2ZSqCh4UhftijHlcyW50tehJEOA7Gaz2XhT9ShM9ZanES4tqRQjYge/r5jg
jGsPYlworclA5/e5u3Kv6W2bIZ0U8UJXA+HZ94bPb555P1ZKxFm7SDSzCSa+K+y+M0Q1Jtfty1cg
oznpqQtMrdsmT7gkEcVq9zW8mFx1piZ5w/YdtWGp8H42mTLmVKvbc6xqUjwpjM+0ABAdTwHk/WAY
b6V1uyY43b6exsVePJzui/9o8y0UoZ6mJKMI1mK8SNcp31efnoB90fc7uFo/t8QI7iq7rXZGBxjX
cRmH4KEzvdE6z6fevan6UrDYtdqTuVkNT9gLxI1I8hpb9GRpofOoQcZLCeCnymQuDlKr+2r0OfWW
qIWM4vngaoIKyezwkgvhj9zx0QJW1/HpOeRJBWtz+CF/1ooeJrAPhg6/ShlVhZPy8LJdQlzKk9mF
WAKSIVbe8rirDS+iyPB44Jf/5r+c3c28hT2cnhsgDHiqkdfyw6MaNGSKGe8gZqE/CIxbSXeXZILN
qKTYZgNSXeKG6mHtALN3vJcX/hHI9zefFoOfuQo49/JNj0XbfP6X7UXSdMiJS+tYHIwY6ak8gw3r
CudyDlASowwCpv1r/md/oYsbbH2k7h7iDtIo5PBpVsQOaEFlDcM8oDr2lKkoJ5TVUYN8zU/jxR0z
CKj0lzCKLD34pHPCu9UEbZDAFMvlXKhf/COVrExk0U1E3++PwetsUPZHC1JTr9U67irLNs6N/zXc
TKv0kkmbtS+T+c8DmW2/LKkIFL0WzyOd6ktV6YEOSLEQXNGo3OW5D8mJPIhbQwfVWzUSHMJ8loH/
AKCRRuR9ivk5qlzjwjd0p1fghsD2p4RuhP08THnZH7N+/kQbThzCj6WPhb/1gbPM1H3ezqU4p5pU
bHbaTSv4n7DZ/JRf1HB+G3qs6hrbwbCMAb/KFpkgQifzSK8wNi0ciQOw75kwDEX0rdTvlKyrwW97
JkpoxlwhfIjreB47XmS5HeJIArLx9Xkhzks0uybmkxDseCa5Mp6ZUHDRqKz9QSElvmLxtdZcbdw9
HfSj8Rj0Rf71RZ4BZkAknHmN2JoYPGmpqbqdAdeIyiueCqagrzfkFBpqJFfnGI7YlDYshF8t47yx
Vi0eD2drMTSJuB/mPq1ANoXTeuUKoYqp7gLdss7K3SbhHQlLupNreHiksgh2VKg5b5EOvh+RevW6
4S8IHVxopXbjXe2Uoe1VrhVO7FWaLYgymb73TowuphqQczs/GyzOIlUEvwK36H6j/MfynFOolb/6
ppHHZ26Mhy3mZ0vx4vqA+P2DOrZoS9NdLzRqkOtMpjQ6WmWRv9u2Ye6giLpSkqvSJ2UNCYj22QuA
EQcKMle/9QrDMaw48asgOYda6NgimAV1piE0QOwM6SdpBHS5991GtN+2HQGqIZr+RBlzZmh+hjC7
UmEMj96//bonCOynouG28B6cAjzcfl6u8wISMm3kABkenLapygPs2EKV3jQhmBMufdPt1fx43I9f
hmER7s+7CrKI0bAxnNoTwonEKOamF3Ko3pp5XF/MNPttgeWkDviXPVNrrjKcjy6hv6PuUxhHQxWU
wD8y6mgcz9py0dalxc5RfbpwCacjlbBKq0B4lkkCAp0DinYyoWECW2HnUyn1A3aLBYz+3FrKZs3k
vtjROMZYpW8VcGCPl7YSu13XyJEogDWem8usNRX2PxuMkewNmXMtqymZ1ivQEEG+ImnOwl2pFsRL
++LDgPV/PLu0HY7xEPAZlVhkLuhKhmDHhoyiMQ4MggZZOHzcAMWmL5IRJnNTLAJx+i3nUvl5JyBh
RNGqrblBQPTdqvlItb9wEueBpy0xlBKEjBkq9tOylLxl7IsooF6vquAO7IBpc0LCZf+QLYuDUwQU
jfXw73bhToVdn5RkNeI1fSkgN7X1+sNF1aRHBO9+VEzgs08JmqUMo3/CZ0VVUq0WDMW6idhcea8B
Qiigr1mDH30ClYejS6BeIKSHb6eej/yubTt2cQhkMWg/3lxZfIzuPm7yaVm5wDLQEoPHky49eVEw
CX9+BjcLna4Ww+BvcZxMl9AUHSPLqNTtwp63y423FGd0+MWIbI4pxDIFMy3K4oE8FKg7YmgmibqD
QYJgZg7noEln1p4zhxG/DHPbeh3TQHuMgE00A+0Yur+6YTmkexQUbZ/9+qP/KYA3wguBsVxh+ZGn
MB2xo8Yik7uDZwxJzs7ESMv63GQKeyC/6BenV87KK6AKIovL23aabyBG7NHBk74XYqheMlsKxWZn
2LDw91fFdSYxUVc0WCezcdCQ+pDXXLGq8G65XLH3w81gmgwhT+RR5eruCFyRLoz1g83nqceSr13o
j6otg6dt4fOX1hE8ihFcUWdfFhBpEbawnj0cGQR4j6EZe1KhXMJ6AuJ5qJdWK1H6zOfchvtbOrzP
d0PGvJshBKUI/Fhg2JZTVoCyu6G2FJ5xrZSHGjC9ifetdcwrZ9hHCiZBU1fd78FXHfij//bkLfg7
2jjBS4AaJbFgDLp2hvfOEYYiK7NnqyQb7WXXm5l1fZBMR3UlpjsDfCzHacSkvzY6xdKXFEZS0fqI
7tRSfZhbR6KgXTJLhWlAbz6kWUaEJ1MGrEdUW1RVw8tfejO3e9Zvos71CN95PfNAdOM+I5CHEVAz
mvb+9CMfxDba+lu1jz4op0MxLwv9CUkekbAPMVYkgIZpeFQ3usdxAdY9b/kYxFn6PQgPgPZ5zLVB
lIV2Lj39lXnF9pakNyezVeEDyf58P26dEKmaPq8JGqihWxnWlmsnKvJI8LSrOTQIUu83Kf0DeGqV
Rd5M0FXV9Ul4YQjKnppEXHZHbdYUPVupZk3dtoAqj8Sn/vE0PigPub34Nix5jMPKYtJnn2Y9eZip
7JQrbQZDUgP8ciAuS1YVXWjrWDDTo1B+5nxclBDHp5RWfwNcM8dV1imHfPOG0RxcTF6YlohuujiA
xyr7DtlF20XiDuBl3YZlSS0wAb641bucRSVe+ZIfCck5Jvt52wQ5j42uiAwoUMpbD/sQPXLOlVS6
ZWDFY/Yb9SZXd9IK/U1Y1/wFBah63ETPN01Tjr5AmUs8oi4r4TFYofrW5XX5VW3eJYOMRAdH1jZd
NktlOTbG01Jp5Xf7YEeaLAcsHtpD4JOrvTJudsgVqHqeClCdwHbuje/VK8gwwbyJwanPYhTpzKlj
Awpor8RWLVDP7fxlaYHDhqyePO2QfnZgDbdac3aVCkOS/S9+yMiOpvfoT4oF2gPAWBOhNjBEya3+
d/XWtCP72GbG8GnmMCkygvjRye1KLG/7gMVOTOkLyGAmzyd8LbdqV2K/sV5UwJ+aSq8wLFTVzbib
WlMiyzr2T6Fa1RnSX56lh0fG+qWW0vrjvE3ql+xaWLeyufqek5SiybsJ3OSrv4PUsZaOp+m314U6
RF3Hq0A4BIGDiSxi1YLpfiaEZLjlpZu66ghf/a5j7//Gv9AGujLrbwAx+mwOChoP6jLIfAwe8NfH
7eIGfGcLrdaGxgyfqCJWI+scYlR8hF+8g5HvCcEGyRfdAZVfEiI2RtZnTnKkq5rcO1Ei8Zi/QJop
3/ld7HhrgXmU5pJGYRhwnHyzwt/+khhvM8NsXv+FirRg9mPhS8vmdcltBt+90cQ8xK/wLvJ66A0L
DicqDWrsQEXKRXu1iXXV1ykXI4BwMJDZ4+bQXmqmsfmy6AVhZT3Av2QggIaIqe1PgW+09oQf0lFL
Riem6rG+skIwXxIyCdewOuEgXZ2LAf67fEfwJaSiq1AhBs/4V9/VybF6Bymfl7AZ5r9a7JZ0KvME
Sw8LQ716ZwcgnlwvMejsCaNTq53hpObv0bNHp7U90FW0tb1GB0QXotMQa4DJOQ2goHSQdvs+GogY
fht/GG/R5tVzEiv6hFU6M0AbMNmCCiN9AYS44aLQhifB1JxsvC54C6XkB4/0FzHtMMuiT6hN9CYs
SGIimA4XwC/sX5ofxMqBSaEOppxzWyBLpKNDGM8fjko6IM/Q5FK1A9IKjWKqoa/bjdJTKlLlsWci
hEpm0JPkpwnVpHd6BuAjJbQRl0QKQxS7XWPNIrIPTvtsWcS4/+5VzYnIyNLq/NQC2ZiqsNtXZpye
Gaicd92gRS9dC+x/zMmKSPFbLmO9tB39KjjHpU3TTuHoVZWCrSPvxW6a6cefjtKFaFNFADiuTNut
ACubgNakuYNKvQ7LuBnijIrTLWgD0+9wWNjtO8Xjb0yDpbBY+bDUz+6DT42pg4RRzYH0FHNi2AYj
U7QwQ887ZpUqzqfCzv7kJHuIQBtPVUcPYwlWKkj/kU0O6m8seGCz+Mkj0SUShFYK5ABOu40SYc2F
BihfqAmkuCOrL8AuQR4rsQGueuAw1UZhaQpCl2W2BLm2ekCtUK9voL2TQzeoNHD2y0zoGmPVk3bw
p89wn4YjbbGSv2gAs948T54ivwons0h6lXcQJ81wvogEOjoQ0tIgTrNEFi5DfhkMjxnid6CXuJXq
gWy3ZwZphL9MhhVGlVX4qamGh/BPRIplgHk7FJ/0IJJGjers0yV5hQBU2RLM+eexCsI+TnlQXEsT
5rqfD7R2KQ+aUPU8bHWluTARLdibWS5nFR6zeMgoHWUomu+iM5fBSObTcSGFS3ZukpTmLx0PhrP7
M6I/sWp+mHoMwMt+HkYLsOhvpkVDRJqjvy3VHnIVwNuGdbx2hF30S3KsA6uGkM43bvxo0WSFvhf7
SGZlMGfYujMSexxf9d7jw1gXC+QAQaS4eZuITsNd/IAvvWNQrRsQlMibBNwkYrgVya9nBkAifAYX
qGOchZRVgUkOqhufUL7dvVIK1Jb4e4/IKPYpzzXWliwyXf9WPKmth2RYDg3370YYf8mmwWGvReok
/7aq4HduRlmIfYioZrswUJBIIBrR+zEgjQ7LLLizEJ/meRCB+Fu0EFHmrnn2GH0BQQqMPj3sawFV
T1C/neRGWk92OpH189aOZH9iY0UUi7RjOAYRowlp2P2+KmuFP2fdL4NC3Q04fZ+G87G/lqbux0Vx
RuInyEnbV85jdQA/f1lbIVW+wOPrjjpcx7/Ehe4par7X0SkSNvAD+FvEKr0nWHjWjsAbK9+syiAX
Gqeo0w+5POZJjB0AdzImE/Zlco+lwdYna62z4L+KFwuM0VRsRLOlX5XZcf4Y79F+mWgOT9AjpVlp
61v1p6Hg5IdOcAi76RhI1SfhgUSUKs1VxJcebTZfBlwSYS3m9tIIN2H++8qizDsoBRLcrGjmCjcD
E2ki+vf4OmgbtwVeF7Ulitga0Rw/qtF+mBhVf6B24pEmENZd3FeivRTMfM/qiXUpvH1I4YA80HjM
jJRWhRb4fMlUnG5QJtJL2amrE+raX0oiF12NrcjkGp4V0D4Kc+q/MuVMULfxjo8Kmo1BGwr/my18
BlqjwkiXG0Za5OH46xbdpVBjVNRWmB97vKdPBatLQpIH2htpWGX375txeAXcsn8A2Oltff2hNXag
BuB0BfP4PPOsE8HB05rGcx3amljT59qSPLBWbnKckSit43eCTJWEz74RaUL27fpz7SOeCcafwD4/
ujGIzwFfIMy8pfs4rn6Wmh5ewr2cBuh25AW3Mtw+R0Y/bRRJZzPSod4L7wYdWzEPonuhe1bPSsW3
MmXWk6UUp32sLwngm03YpGvkxqVu2ATqpukTw3CyoGhFQbA2LB2Q09I+nuDqSA218C88RKPYEduY
5/S1BUuxpT7AFKts4cW3P0YTRKdMcLmJwcg6qfuvQQ3CdnlSEVT4z78pnIEBJQwCQ1VuLoBl98Ll
ywWnAKOpP2/ef12NQ2mqF7Q/dsF99p7/QzLTKjcwRRfj29PBTQp/Fo4BYsi89ALmILNJP6/WiONP
aOTf3N/a4Jh+3iL09dIYaIXIy8Io7Q6OSn2Ai73upGSvfAT0TkwIfqbyamcdVXLv+oBwBHoUfUct
MHucX1eAP2J25C6P+1vk90QEfJHmQv9J/6tuqNJMl+1VWrOMJrfvmfVohPpU8cRibFnVo/VCC3ac
63dB39FlTF2nicX5UPtHCIgJBCHXShG0QogKYiotQtb3WLPmTwZBoc540lxfcjizPcWUj76evwpy
0yy+TXNIY3RrWBB3mKdcy9ECYNgYA/iyBho5u5+CDDnBY6pmdC+73AJ756yXEyftHhDNHJcqLbMZ
f8I62B/d3wvX+/n482mkC81IppAEtbMFTW9e+ASoosuBXwhpE6KgnuedvOPaOJ3eg7+Xx7WMrIt3
3bzTifQ3xO8Y4cfSlOlQllmE17GIVPJQIwmy3Tpxn9ZjRFLMvQ1YHZmkT4XtPgHDDWNfMS6YM2QG
UhFYlLFsfsQwiTlaM7YQfhxpGKYnyHbBMusD1NQk2BRX2EUgOh8eiBtDQX/6pT+RitNdMaA6gvAz
GnorohDSKxgwaX06ZAHeArjRKsG2dYQ+amTBzdeTKpSDOMDstiQwjJFjoSZCa4Slw7nPwkqs/l0G
SMWSEf1Wy9FQUSHXS+aVdJg4+aT8pMYBY2qQqTddbtiI8Shb4TBuzmFqxPQQj/2ipDoF/ZO+acBo
sR4AJ9i36Vh6HcWAeMsqBO9XFl4JL7LlP/SgRoUxYCFzb1NVN+9Nd96bno48Yg0f/5R74n6MiBtF
viOPZxlnFPkMlFVfmutC32KlY+TTergxdX5e7mEkL9tUwBuZSf9QvVcd/FOeLmeYz7d0pl0GDADr
BYoaxp3vqPwuwwhrKniMGlBc6jEo5hEhkb8ylDOtsEfvVygotr5i3HKUgD29kZC0XGhBJ5L4cFa6
NDzitL7S3nlJweGliHdgKdWrpxpYPNYKAIUky5rpAh8tAiAb6xVe1wx7wtBxp/3CqBzZUaItJUEZ
fPiEgHjkE9xUNQu4KE9G7IxLNQgGgrR8/dZ3BxoX1FvP4NI+33npRRI7qYKshql/THQpEAefD7Oo
wEHsggFKQjdwV9ML19IFukyfkA7562fFEKUSIdcEOSLtDAczXG2rIhgdDxwBSUhgtQWlv+2SPsRF
BtiIbW/Ar1YqWJBD99Jb8y5KNKa8DqeeP3KqRv+XhHRcDfjMm8iey1AQ03TImkgSR1N2ybbHK/f7
Jk+TEzBzKx0NZnm42ni1Yqz0fmDg89mda22s3RAEPJ+mFBfyRYroB12JrsYMLekv8eDwhJ0eC0SH
uxOJOzeStEyc47hio4wYhwYAc9raJnk8yTu0rNqLxtFCa/4a9gopBSb1s3Y7vSmxtiQBDXGwjf+s
+OaqhF2N/Uw1HGGqHZanAvl/NtHrt8gKNG5bHPNCukUy5khjr9dW6YW+hODKPEi8S+2c+Mdp5flx
5QLoykTVZZJMPzoaTOch58QG4kgVjIG1ZmWnrTDZmixk15aVkryz1UxdQdbcfsWqoc+rUmLXYXfv
474EjLJ0SM/ZEdizeaEDq4JrdVBZeq6hSPGeGbGco88JAMLMxvINq89+7+8ObPxfr3IlIeck9Weq
pL/Ol5YPcvmyZPH2mt8nYhdTH/JqpK0BAy+UTj3jIb6Xs55hxiM7WpAxKHTUMqxXvDDtstVqpesb
yspXvu+g9bEeSPaWfFkbRCNQoyc58D0X1t+6cPNP7TBX05gfkpWzKOcY6N3fr+p5zDn5IWySWFgp
ULELLLr4a86dTACaozdv+oK76uuPGlxDT4UMG+OJtJdPvnYYY5HPZG2meLElzgYlCOB6F2bcy7FO
vnteyP32jym18+AKq7KqxPWPiEziwYL3q9SZT2w2yUL2j9sf1T4IN6RAo1Y362Xvb4FTZ2bdVwuI
qayrcIpLKVTTyVtFqeAzsvujR2XrktmQCtJfI4rtPd/jzreZ+z/5BiJOF/hq+LPfId4gfX+1weey
TBQ9p/Rb9uUj5ZasTholQt4E9xOB1Bj3BOOZiz4T9TSzdz0xEi7KN3iAAfgfQ6LMqDVKGNNJb4rv
M3S4zGQEpNnejDfhGhcc8Jv53PZMdj01sS8e3fy+5otaKZezVF9AIK/x+VRCdqCt/hzqpLCVUnJ0
W7Kf0OrRQ3QHKPkkQSW5Ez9edWOegYczMt9hH0jnc+KJu3lbz4pI7IOSruduyEe+daqDBQEXYrMQ
8nEK9v16PU5fRbVFaa2mIpNtfUp5TYDTwYwgMHTJCAqcuKKYPEo65EdMhVvtsIBvkTBJyOTfCybs
o2C0kdZP3PLZ5jWO2YQJEIr6iZEMMGAH3x+DgcX+xhg/ONk+eXXvb4JAZ0SDQdTeAhqvrfzy06b0
k98OQ+dn+8Zslk7JPjeH4ZE2wCbuLOaLHnQ3nEwKHFI3Z7Y7ZgBv8xOrrcEMqKv5tcKKehsfTT87
rgJz+aCKHA99W0P+gAAdUsZ+AKCZElewJaheICLm0RJyVQdJiKtq3EgUlQdnDCH07mLqt5ihxL2H
rd6z0qdRhGeCVMCPxGSebvC43bjUxdOAblbMX5QHdXXtk7TCkyFB8RaE3qF1UEW6m4k4ohXAN2I7
B8AbOa+T3WzoYZdkz7taQ0tuXzBfLxdQNkR62LU/W9YItEhR7g3FmM1/rVDF0RkxYxDorEBmDugX
1naDy5HkALaAHNSk+DpcQXHxxMvl4YbfKWPrJfrHP9cAoeAWPwiBK5m9wxtY+rHuEOiFiK6sBk5k
174POTwGsG8kjGedmNAOvu3p7gqz9vV1kkPBE80AvvgthWXBhPfZsfqQGvDgUZflnD6+VDH7reM0
QXxaToo4Tu9j5+nWnNFlBfi0/2Z+XYD4NKxfO55O6dyWwdo5MT3+wkgkshVOxJ2++ySG/f0xaQbK
Frx3Yy0H0LVTr8G5t/YiL8I3mFM4JPTkxNn4nzu05wV/APERz9aDAF4mwkac4dmQLn46SnWNTHMq
lPPaH3Yy9HRGFXjKmxRx/7rU0UIkua4M+aeMCkSsC7Z1MjIKoblpI+y3RlySSUSsy+865oZFJdLK
K1CD4WEtiRnZDIEBzhxp6Kss3sapZsR+K5WNL7XhxQypAh0Ux77exd/WV/JTkhFfq+bkkvZ5mxkp
dhAdUNxKjBRjsBsT3nIgMdJTB8gnZwwDL3sKM5RJh09oPruGzi0MvR8ey/sr1TjVe87qH6inX4+Y
kdibj8MKeonregPMYiEJGp4vpKczltKUIZ9SIqA0Px1CulldQd7kvJraWPA2Jv0agb6PSy6DchkX
oyhbzBOYclgqM5HR4tMqnjVyaU6IKtFS4hy5rdQXiGcG8Sv/MxK327nGqt5jpNAQdrX1MJCg4AfB
9R0yb66LO9I3AyiTdR2yr6rsJ5ndtUWdrtxXBmPY7CDM12Nj//F58L5NqyXDReLRV10LaSkNe2jY
7U1n8C+rRtBmdmjlgmm0D7x8UNKD/qUT8bsccw160NXWaTkq1V897hrivlSOBku06XVPCJ69FXJV
EoUg2E/8UosADUhTHZGCGKu9oIY2YzDUtKn1+an/5OKv9WwcXMkCwoM74eKbkN9vcmwWC6noTFfE
Z2BoqBPtyoKlnPxEqPDZrMnzljlobhMK8ZXlcQXkyAatxLZOHUFgSfoigNn6vsCuJyFLF/f6scsb
1g9kIts1XS6cZ1/iwj+fdrzO3ySDF0g6VVQ4/GbsqBA5tpaFnmzXkzP7KjTvNkDawytIXkuoute8
+s+lS2Al0mxJLLlB/3L8VFuXlJx2CfTb63DQEbVl7+iLWNxD4w2xhh+YfSXfGS+VhZUW/5/jXx8i
RQSREBOaTij+RdiMPpHvA4dt2Bmjgy9GBHsH1BAhbIWLZOlr1Q7BreHBwi5zNLm0oqphVh2y3w+7
ha6Fs9snabOqJm6E+KtrN3nKAefjA9LN85hUr7w5GcYFGdqForM0Omq9X6QiHENhYM5aoCQBzPgk
fvj9NSRTd0ws8U9zW/MwVf6Gd58irCgCtuWUizTRqzdkmllCaXdvADQ5CAHklRaHG8dpZ8YgUKuI
dsVn0+F4YhV+FZGlPRFi1bMojkwk5I0/1ppvHV8/Fy4BQskXHqr1m9nJf4StZsOHd+yMAwM4+QOQ
uifC9lWHPrFqy7x8IzEHLIgTFDx9A9xzh1S3nKxb4T17Ys80o+93YQz9ng5IoDQzlf0uWs+vY9fC
kQmGfEdJtl1Gr79h125/KMOvegLjvxqEv6Se4gHgUzLOxRuP5XkemVg21eFVRIsPL2KDyuPMORpo
DNugkMGsy/pZ2NM0VMXDiJI6zDrVuuwc06sbHmfSEvhZc2AvYKl5slvxFoJ/JC2P+Hjzwf8IyGZj
p8+NdOyjG5xUQXTOEs/wH9OP7GdFCFFq5GHqN/A1CfODaKSvmcANmUQvNy1ZigFfSi5s8AXDJ2Y9
iECKwyEYLs/i7r+41tb9BA5tyvxGwpqNKE3xkxq+wETj5ojE/wcuEOq86LavPCW75oqBzUfzEIKY
Gs1YxPqEYZj42hlA6Wqw2dKtaJyzxzTLeJ1kcAZuUyNKUx4JuF8M0MxujdP0z+QKHJZzrsPkdMoV
cdG+9qQQ40yASPCEiD5TxwqGpgiHB9JtZeM5nfHQrhWHbum4j3DKxA42NQlA7D9nuBxrTF7uIfpX
KS7LxLgaMTvmuU/EZYS4otYcfbjcxB+LVuSa5uGvKjsFsRRjgE0FPaS0H5ny6iYoUea1Y9PzNqNC
mMm9G4QsOEe3d3oSOW1+V9VC3Fy1+3B54UA55Yh5lgqkS7/7kC2oCjRWrWim82gIJL7wE+I2KKTY
0dA47m/HUTSZdsX4k3J3xsOp5j2xvMk25KUXjmE4cK7FmKmak87sVUCGM0w6kYat5y/MGSlOw9Cf
rcxwxrKxVgalVz5Srbfb6VJAMgO8we+/zU6uW3RP3bGqdqhie3z9imFNeqWp7VVqziPDxRuDIrWu
hbxacD2QwpZAm0vjTWf31vQU9DAdriM9SzHMzQjqUsBfBNRkOEENoqE4CegvMTnFIuQPZIyXJ8AO
MKoBcWaP1yXj3hqKWjxSSdBDQ3EnAr+NUuko4kGEZj013SbZjVZHpWerd0TP7RRbtwMWJA6EDm7d
Dpc6a5frC+6nh0yL5YzQPlSum5daYVa9n4eRvLKBbFPJcyM9v2XLgDRJfOHfPeaxkctYTEjzfsA0
cDqySrSaCXYBdt0hP9yX6V64HAob5RAZBWQgmTfi1EBNJ7Onb0XFRgMup7uKsKHDowsZO+LpjSEz
VXEUbWoRVBlIVfULoxGThDQE3mqLimaEYZtSR/Q05C34p9pRcyVpt8BGiC+O289RZZ7wpXzIyMTG
J0yVkr1Ky+SlPs8OEzJ0U07/nNfZ0ViUCMDJ+Cd/vuv8qGiYhaRvFkfl6FYl8y3RM7uDQ7yqgCNk
TVmOQFjcjAOeoMOjiJ5U64Wm55JWAJBRHQ0c+Ji+O2dR5qon1hd50K7S3cKNQpmCKGH75p4WdH5S
FA9yypKNeIKblQBCjaoYImox3lzp5V2ggwuB32BmPWoyLzVISAaw+6kMSIOkCknfaAtemwaQ8JrM
TjgQxWpfb1VdWoHDt5ppTQeNDhgUFYsUto2/3LxoFwA+OEHtEonNHApVXMl9rVjEic99CJoupLQu
rvmBmt6SSbIQx6Q63Ta9npCcxtE7+DuxvyDTi6InRLQqLkyw1g4CmM75lq/Tn4Wo7HKbHJXMG2N7
0FCdSHnkykeZ+DNXnjnGz0nLoX63ae9Rf/a527wBcQTg2l15f4XCoKMPpD3acuGfeiSAT1pnVxQp
OtWG5b7uo87Usvd7muAeXsyI71FB8R31ssOJzI3rtZO9Azlh00q3MneXPrO2AZU8Bv50t6PTOqRd
E7jTv+w9I/SPK8L7TsWsXbRPoYKaNIxGjwqZGnc7x8M0hiysJKl3gXcUi2DNpKMxvacl2moeclVF
aVro9zMU6/zpIVjllwskwtRELJIVyIvDLV4Jk6isdOUdYCFBQqVBxtBDxrTOmr4VNqZoq/23i8Zw
IawxTf7NSZcxZAtBb7GszxqewskzrRgS/gFNz24xRuacKba2OneiBfPdugahrYclyp2qRbowNNkQ
GwBqGYaxKTb+uBczO7xaQPa/o6ErCsIRpBZazB6SkmhD4eM8taAC+QYOMJhPiQ7PUEHo5hpy+w2Z
wvp6kynwDt/XAdf1WgP+/SeMhwIBjXGFp6lm4PyRojf15KrJ34sFlOrL7SwvlTKuufelS17zC9Ds
kc+/SgVLayE9/ibB1DgYxkzT3X/g97YNU4VvOPFWw0KY5RGuoDyhsMUsqd3XTASkPhGKLYPfACtR
NCHCtgFSfV5d/kJ1sLxKQPBPHD+vmjTJmqRQEsAyMjG8p5E4m2c8nIquuVq/T9dKEKPFTYDHDWU9
W/BphAi6UYgJkncO84kLC5hCZiBkMUTxIXRPFqMokyqP+1soQFGibxDaYLybRzEyIgGg/criEFZj
gNFGQ7kPVVGP3NNUhnJSXMJj/VJsz9W9fpqbBWhud3zVAU7noY2+f98AZyEJJ/7vG+Y0hDiVyYAs
83A4/dG6SSKUjLq9a8mdd4qKd+xK8AMiPj5RO1xJbf0eXSdl2BO760ikwUqkLzqAxY+t+hRFZD9s
z9AQZh8NzM8xwjcZLygIm6L/KKvF5rz+6n6UrfiwFN1RQ8krmj8ERLE5ndjkkPS78kzd2SjYyg7b
7eO6dmKs/Hn3IipX7aCSTUcxg6qCVXpm48BzBgpEAnGhAQfERlu+hGoBwOYmaZLFtZQrWIWH3/pB
Bb2Z7zwVmUfzu8y0vnNqdcTGYSoUxqgzNUC9pC7+m8bU6FWF13oR7qEiYRECDTw8h4IDKQzCcUuf
/AQ/fRFPTrx1jRDA7rKNXeVkk6yT7XlmqCgZwkAxDJcG6nps38TI6f1KfoJTVxpRFDtIgvmRbgJ8
8ywXfFwLsPD+WSO4BQMWU1oULoTVEjsiWl0QNBZ0bNOSUTDtaMoZW2nyTDF8NgDeWq0krKjx/pHK
zEvgzAmcW81OnvFgJFX9RLxBiKMliBMcJR9BiH0/3+wIjBrlYhnBxKRtnGUIQGaRssxJo1SfJqo5
oVInOU1xvEdVbY27VgEOnsr1RTfMg3HIWYRx21hOcuWkXGABbnAcWWhyC9vrEXzt3L0fwZZT9CLN
sypUrzeCkRBHZD6wixBXdjRDfU8b3dbu4goOc35lr3CBEYY5DfZgvJ2GmhR6a514vU57C2S4Vd9W
Rmf0bDYbmCtpxkdAmZmG6T/GbTK3PfpKdGIpB+cuZpyXw/xmFY19T40BDMy2U0vDLBuQfyjlp49X
qr1EUK2J3DR6QR6KeNgTpkagueNE2p65WhNwIWZkZG1lvlsf4PDtiWsTueZLvXrCv5eS7fKtNZog
8YLpOwLiemMjbEmrvqdpNUGCiNCwS4z3jjCGeP0rPU4zSSJmdA2CtbaMg05wcv9jFYkWIpeqV5OO
rKpEumSoRsNFXsbHClP7cwPsBXa9W2SASIwPFjRK7Ys4pAmNysHf4jg/mEuFtwj/5GTcRcJEzfUH
kBj6vNB7HwPmatPlc9Fgzm1Gzkc+Pv4YeV5rOrCZRCTESypSZuVto8gntAfHfZq10Dp3lAlDUWvl
bxBLw5h3iELPQvZYw7dTZOAyTqiDofNRE680m6vH5dkEWia5JFfl8Ak+cgQ3wd3+fKjxfIMW4eXZ
j/LHUs5EWBVjt+hOJCfAsRkWh6u6n/7zo1rAMLCHRNps2QdyE3CT6OfBly2lAUMbapAFFOSxGqOP
XMGfM+g9S4gen5G6KyvD0XmwOqYHKb00XOSN7YwgwbyoFBJ5/GqyxMEeTSoeGXv6naNu++6Vht+R
ctHEIi0WRSiMM8ESrw+JQEWS2QMZWt4+eyKV4liDIZhqNvTndxSekMmEoWadNL8JtcsaRN4F+Q0E
9mL9FxoeUS1nygaeFX50lv7YkG1VBADLGXdcU1OgsPfwDd3XGt4tBBXeM+o+Z5RAS/fuET1B6/1u
SPOFwtYr9NgXMnz4P5qNKXBe2q3Fa5XuxJ0IqgJqszvkqndKOE/h6Wx91WctntL4bcvyxXCYfJ5O
rwbsJPhOsTez/m0d3Z/VPS4wFtWqUyppxOdEpdwn2KGmUcjT96D6+IVWM6ozCbwIv5NknKiSNCuE
3jHhOKuSmwPPmszH7yI74k2KKEHkcJPMilhZdLW/NSoN185MoWQZLQkF7LhoT1ptD3twORcniuTC
rmZl77d7x/IuiFIxEcT/T9PAPr7Ebvecm3s2mJtXHYMMJ99sI/N0k3FO2TOj38C2zHQF2lcMsm8f
gc+8VaFXiREUGRCrAmNOtv+7t9uy9XvhhwTzbWzMSTzg/YUrIBw9S0ImOPe5oQoJH5ZbqQzs8hVN
lnLYTDRMFGp/BcQ4ZkTvXWDafmAO+o9QgYePkRVqUkQh+lEZXnbbUmrax+YHXd0i4lmEy0dRAnoa
ybZcNAGI2rPdB/KTBrhww9qBRZdH9xpAY0cWHEI9PmpKy59cRSBu9VUKNXsWQjbY/9Ul9+pbgmr6
1m1E6dcBY9Pa5uQubjJlUuwu8yGlyJKUdDNEEVscQDVKhJJZtG62pE9T1XdRpx095JUdo6zbnFAc
NBJbSYBy1VT61fNeu+RM15O5q8fAcau1SDa7LwcvBOd2cKjPR8M4I9jMMGMeIYZeFNrUJgDT6uJU
SolBwpdSbwNb24DuzDZl2Te0eBDMcUD3p230HL3J2OE0glpLT1fQrGeYxSV/q8UPbGO0e5jEZuoy
gRrg9BISNFHNnXpQOXt5erpIeUiGYwBEXN5yBiAA5oK/jNBWfEH1ofHPfT1WIouYhWgLV07rGKLy
C/ShsEpl4O2QfymlQZpTulSczlv+TPIummpKLXG//NrawaPclABYCGE4Ep0sdrm52EGtZeW43QtG
N0BNEies66dZg5v/eJR7T3+IvRa0qxMZewjAZ3hA4VKFX5yrPmJTh/Y2Z0N7IY5lrzK5fDSd7cr1
XwyyO7dKZ37v9zM/s6xK+7jB/FGPdX1T9JuVM4hNcacobPlBE58eWfBD+Sz786byKLdYDcFIoG3i
O1AAm02Z4Va4CJNo+zg3FPmIlkqiNti0aHXGhAwVxnyoq6l6M1uVPTJxhx4uj3mjveBnTQAmU6b1
NIBwRU93O8N2u23l7/wGKm3iDlMWciGOAFdWsVl8P2/SPrVDBhcnltjkRTtZnfji419on8AB7XVP
7qMn0NJydJBlDAQCQOJ93H2jAaag8pflMT+OLlxexClS2LcRNGXyKN5iHGxXejimQjfEy6DvOMvg
VtxKx4B2ExwwCGE3SlczbbaE5EXaXdliUaemJ8/7Iia5paUO9o2tOBIxoGvtn9X6S9gGjk40Dgxq
RMOKQ6r06U8T7TmbhGV4of4+vxEuPC/+UWPEIDGtVyv6Kc4Ps3abggvPPcsfEZawEXsUBkTS4V+O
P+zxWVR9ak5jMWcGNbX31NaqJ+RWoJBmbbfbvH5jLUnza+y/zE2T+zWy/ab/l3Zk/Gvl56UUl8eN
e6Q8OPIxzLtv/MpkbMd+IvgxrR8njAo7+2DpEK+UsjkhsH+AcEqo+Ux2NXy6GJAE+vzHWdo08sCE
jYtmRzOer5g8w+AfTaXAWpjCWXmtZnkH14GDpQmbpgTRQiQ9mopXXa+YWrXcZaamKRnb8UwktJek
NsBOttTqLmdi9wBKpFLRZQv8fdhb0rscWEFHRG5wE/jZ7w7Om8jxxr+piIvqF4gzJWOEW0R8R8Z9
xGSrpKjkbWmXEgQplgUaVK99n4Etl8x7WdTM6AYwYMDJPoNexr2jwkd7YozurmIalYJEaFI86O44
2JHqz2ucCIQvhWeqxXW0PT4dHb1wbHPOQVyS9ub8HRP8avMmUJikwzkOzWJUtgJ9KhpMEySyhLp1
mBTzS0UjRN9enVybQ4V1yG4WqTe7pg+aA2X6XWHC9t+f0tz+1lFQEolzTk2sFTf4W4jIAomox8So
/8M2maU+Rz/9GyZ9CElbJwOSqPi2MTy43iRWECPXgKHk2XiIpMyiwwCt9Db4kpuhOzgY7XIdNnOw
l8EcYM8t9OuFA60Rz1KzYhlJ2tGKiaTlakonMDUranqjw1ztSWiDHY3ELBaXct/zEnuLuFeXbcm7
IzbThwNh07+7GPjvc5H98VY9t/Jyss2Aa/9apbeTivrUMv60NDHCaUHcdeDt7Wg9LH89d3dKC8EH
cIfEK9Wld3qBrxvhrSDTwpHSzlWY7T7MXQ4q5CP2SAvuZ814qYPtNmmMNEwJXYIxTazozJ51LRKy
BPe57DdDDj3RHxkwpPv3+X2/q8C2INKGORxeG0+DAMDqqFCtvhJSK1p/c+PHyyT8O3cNhO8Cjmyv
IfE6tmqlw2QXUkJ32MYmiyfLfwvvxuFLwbKw+EZD5Rh5w6X/Bfm1psyRFYmImsKBoLPlHuXApWdj
cTRvXq4+gMA+cIlahoBRoK3z+GRmy7SPNbIJLjbcGl9g9IeSH0DBE+wPkpCNzkxpNR6HG91kwhvg
XLsqcbmtX42cg+FaFiYtoETDrE8EbOqwXupq1y/wti7bZ2b1iDmytjUUs1GtduXnspfhfGoeduH4
RXxrUwFqUt58hacnqXQYfLME0WYNTg7f9U9FOrmv7nXrxdhnupuQvOcIqYRxAJHZ7dW1tlcNj9m1
+Nv3izo2DHIZNFgHHF7J+j3lutIAAwPb4n1RTT5rsYzml0orvGX1Qj/qtD24kDYHXwXklHtPRFLD
nXZHOKb4W7/3vzgTSGqjTnmEMwMEMqGInbEHbJBv8p8cMpSisXnfyVYpwrLcXxSMnca9mZKSEGUJ
syCzuZ/nWnC/jhSIi7uwOVIxj6uShkgBQRiyOyTUMfdKiG2Vl7Mo4y+1OFT6qG0HnSEjUG8OjHGQ
B5gBjQt40k3wuzGAiea9YJWEX6EvFCvuGryZnQnMDfnCEQhJ1yvwnAdZVcCltFed3z7B7JQ7pn6z
V8Jwhg3mAYfLywlRT+5sqwuU3ZnvTptw+wIFkmIvtEywoJee8JihtLUJgl0S4XX1mggWfbUhzPu2
2XJ3hoR8HLw0gc/fm2rukc/BiqDi+f9MZvlwLBVZRX82fQGPJe+fK4Vgvjzf0bUkc5COkQLkZQXK
VE7YBig5lWofOUJJHJVNfEDVeM6g/jjL6BGA4yX9UEP3xb77wMJtJ32brkogV1z8Mjz7RJD95b1m
D1zuhdq8yIdT8+pHPPiTjXaL4XjZHCPkdHobMgDIlwlR4odjQ7rkpUPmxnF/BQPcnH9myjG6A6ug
5z8Oyki/Q7sY85SDtlX1EIIHxQLn6MqEnV/LibnBoHxjfUUAsJkM76zmUH9C4nZSsh3C9oY9csQ/
fyVu0mUXopn3j/cX0uahUxSKZW0vmILMBABsSnvZaPe8vB7EsqMD9up9AL26h4Nhh3nMki8R/lyL
3+JmsG7cfyCMdlAEpjycKcRw2M8jmnATMCn3yl+W/N6A1ZdlZZA/0qYz5Del+3+RzW0ySz98vdx0
wbq+ffYvNhwctMkm85W5F3BuyMdTxaCYXwG6j26Af8utR/GDs7ZEGjQRKzFuGFAf/h4nVcubeimo
g8eoGiA/NZECE3dUiyk9cH/r+Jn+oI6ZHga9v07q2eXPzyFBNoLNYcvbrXZgXLF5NSWKja95qzcq
xuygLqR33O36LjxOtVP/arSMZL3oWKBP6/oQnsTe676sS7XUPZGp16v8YJFfaZQhMXm3WHGsZ643
41T1sg4pdoRliJ4LNuK7hGnI1yo34d7BWNCQzG4tY9dYQr3OaK+6ZOQdF/fB01vpQGnZZou2X1N9
U+5OedtNL5J2F1CLtLXYqh/QAh3lexcW5GCAadywf/MW5YTAvb96cDDw8+rvNvi0z/lAc6DXeMD/
GO43OpcB7/MO1uDpeYntQxXBPpnp2mjBMuVFnTqdau1bxY1X58wOfRrTEBaSovj5bYCRz82GKbUb
Y2X/MKbo74pXi0EPYZB1ddA4oT7MIYCq3D/73opJrVDBjvZOnUIik/ZfBQEoFw5qK/KIo0/03cuj
CiN0LgrJ76EcqInPZ1mmQhtDXFkrt1SJn2HbV/b9T4x8zVjnJ6W2YSnOp8x9fHyoINBfsFc42AFi
Op80hsTUCEFGg1RY2748Dkcx6UXDwqwN5Ida3ohx5FlekazlDeRu85896Dok+7r/68/0NkD013p1
dLfY1LP78/piUo67hBaY2+k72jNYdNgS2+pjSZbfO9+DRPWItTxBxRvWUOZ+JGXEYW3xs1/kKfi+
VifZQYYjQVMt9ODgqwS4xOjw8ILsJC0MQkcglYZDpkCdmx4THpsSkttRSP+sdFBogSaoKEB15M1e
KwNdTwpve46nEFG7Vuq5e+PNUyKvPn095rK/k+D/woBT7Rwo6thG/LrhL/8bkU3MXiQSHs4WZ7ni
kqPFbM8aG5ILDKCGq5DCXg6aWUbrpYscQj66dEM31qLUu+KmRzbQuHei1WZS/l25SiqcjQ1HZDt4
B6pJg1yD1jtQNisTa9y6igMWIQVUlh18O/lj+a5mZ3E9xqqknwDGbtMCMjNgKoMOJ0vtiJouaPjX
alYmMJjsS1kZKcXqYh07jbQT+LWXwtSCBDbJhAP1cMxAaUFvj5HIdpfxt44TfdqDR/eUbmU5o/dM
IVEv11UN1tvRy0j7kYBJfElPsDv9u7vBYUUeS8+BpTlwOpemdT5AlyB+JPml5fbT1I5DKtmnIFUB
mAtLBsmoj3Nsl/9glFgw8si6VnRrO6zoBwTihEhA3OG5+cNW6bB676T0rThOHQwS/+yarH3hBuQH
sW3YqUknCl9x8sxG9EAGp2ydX+5woiO9ALT8PbFuvMpHrbDX0TdBLsO5wzmZf3bCBQ3TM8JANX1T
aVDwxJVwx/5cZoqrI4ZWexws3VQZqah74lT/n4kYvpklPVh8anrwUWrVWMg451Mj51LhPdY/U84A
qIcHIkyuK5MUhOwQUsOKK4Eh0OBi3DXjggJtq5xhMjK1MOZbRcBXa7MU/HSs4T9fzx2u5GafCxrr
DbPkZmYd3sEPtKN7+OYhrmd1C80MQRrMT2S1dk4J4z/HqZcvvr5+uaPnt8fKsvwgxKr0m8eJHo0m
zRQH+IrzrJeHTVF5ZEDn9ZLpX/uebsKnNSzbEGDXwPUK5liFC8pec8a3nAYnUY0oKI+ZzZUZk783
yJP3w8tH4cWsQGpYTQzr5ftv9vO96kTtiGos99G21kvvOT2rAUj+lvvPdcpsPHBK5N/B1ulvzosU
OWUzuZ+gcAsmRpBP0VffAKMcxkD0l03ZXimZdRoJ4cbyLtYSdQ9oBqwEAcBSPz6Hbg1YkgLDNdMS
oCkjz1HwM+jt3kbIWwdH3MPiILAqumemz6oOdpMf5HkqJ+1RXXGSmWTIQU1Fnn4gt05sT/8WmKrq
udE/92VxRZVBcoE/can+ojCtvpy2Fuw4lapDJR3PHOKTTNyZKuIR5kG0I/aDUrB9RqTKjwz+QKG5
sXdi3k22/f3UFoCasBPhogtA3Sx1YKLJsP5APbjBKHVwvjzYAy8Q1ZQxZvxtT7/ZjNW/S54g204/
B8JM6qPhkrqAFfRtdXXWb3XCG1hdTd40yW2wlhWglwaT0r9NM/8Wy3eZfBcX+TRLb4zGTa1JFJOM
K51iEtfN6ykTsXPPU5LYdCr6s+PFExEpq4hCdyoRPrR3z0HQdJqECDDtRFVKWldX04pE8xcZ0Zw4
DmCcFDwvGVI1aTzJzf5h4/BIgM9JotAThJ17gi/fOeTJ21lRbROwDHRJ2Kg0vL9/GyTkl8BmYlQ/
GTn8f7WkstALffOmosu29OK0IFfUDoKCpYuhETkn3C05PFv3Oqy4gjKIlwvGB98/4bTiOQFoX3d+
EWZg9Ue37vPKDgwWbFp140v43jSeNoAYxJc2W+53M+x4OeORfUrzN82Iy5KV8PgjiQF51OJRxEo1
D8jfNd1YspXTdlWTLKC5UP1EIff+aOQtBJNetXVPziUGVkU8aorPwpZdAL6cWZxUYD/btm05NlE0
LxL7u5wi9mLPfP1qcYnFK5e40SVT457qQ+CCSu+kT7CdCxWNj+/aCg/Ypl2wPCFrUS/xR7cuBR8n
u2wrKp2U0ox2C3rW1jntlovkkKgBiorZ/rwbkleQAWGAnUKQglYgOaDI5GkA/iT0ycAXSqPq0vql
jqJyJOU+driYxqXbcPJf8Sj27sEnrXGUTnNWYepQ/wdtADec4MUBxj6qloJFCL52niAs+qiNtNNt
k2B592LG9lz86zyv3+rxm05VggHmDcnrDRn/iEO/aS38ks3dbSDbVyo6Ca6PCjMmcl0uXKYibcLM
nDCcMXKIAIvHfZ7NkYQSJDZPQXjW1Nfs1NxRDTM6CPnw78X3PMTJwH/9xkwyl57k9lV+F1iSqyyT
gRG0ksbm7bZmSR2WOrHpMsV3sW+Bz1XCYnl/guiOwTHtKU/HYI1bUP2kas9rpXTg5z3746RYqM43
apeVC99zEf4Gh9KUXGKo81tjhXbeYSE/P+OQc0ECn6rFb06LaaaMgACdKo050Tqt5rynuNMOcdP6
rPlE5qIo6PX05oRd3ECVPA7DtFZGRaFr/3E1cvb46rhytqJnu935TvD3CbD2I02Adg6nVpN3r+HV
qglGlmr2SloRUSdsXdM7FLkLKIOvEmoB3BLMyTT4AVGObYzjUg2/MBPKrQZrXh3h/+nEtQdlYaeK
Z0urb2Ge5GvECatmcrYE4MjW42L/yoX6HRLvSBnjHFj6DVltx39jo373rcOLdh2l/JMQ1hfBZUcw
hoT9rfD8LIJNwJKLGzVznHo2Ug53bwhDCQCO4OHf/xs9wSTrgcN+qleT6vrCXqphJzxnSyNxxkSa
CD/PNnCU0b34CiJYPDaoF2v2VtcPl6K+gWXSLrIy7GsKEw2lZ6rQyTXOzzh663IAKhbXhZRsOWcz
x9/XXBsx4CstQBcEcmSmvD1g5LbuJDKmbQ4L/hqvjUZfMqHMZHNY8gLlzOTdW0FQh0UyAqpznZQe
YxRaUAJHjWslXOjTfn/udXnGG3vZBTfvOUA2anxEuf9vyHR9war/X4ELHCYM4FGYl+SZlCVPIRI+
umJkD+vOK/sVLeClzHPZ7u9saVexf/9FDzffTQKQ+NaQqniDx7oab+kKBCOh1QS6LobCRDxPpdVw
VBbGrCCgsY+954Q4IY9iSDdYSFL8+mst9p4TUGHz2P2I6aVVRpMhc3x0XOjg8d2ibkGauE0GrXvQ
EYJZDq+OTpXEmCEMyEjnqnqhh918DKYUspzx75zrgrsJ7voJcolgJwDMmqyWUif3CCR8RTKILrwv
LVX+9PLhsj7tSlUVUIelhncfyvLOJ2k9enB/fjS/9+J3W4eaiOAIISd73tkcngjz3qFWyJRHvwW4
gC+0Io2VbAJwYek1A1wxSZyID7lN67/6pXhsbRjk5eXg87n7yd3BJbKFF6MNgL/PE/T/zifLC0Us
JydAq+oNGN3guZCiin8SRounTJYif7+TBhTwcpdbjU3uVdlRxyn6KlC8t9uG6dt9Z7up3wafaDBy
ljuI5ng2XOdAGRyNVomXaUEIoYXHnlxyxH8nx6A0BpXbZAhLXU+eUtEt/aJ89GcFtCzRn01NT1at
KEvwdzGMzckqiOTkSIp9FEr6DZdFvQTnu5HxO6J4Nr3jaKw2Oc/wdJrju5HbEdpJMXSkTUPLe5qW
H8bwM6NV7d8pyDhamFDOTOLvVg4oNzLaJJXbCesAI/BMziTT9Ci2JxkTBTOmC8DszWd5VFC5WNLd
tRtzJUSYGoJ7dMERtx/tLMOx87sY8uxwkCtLxts4AstcNB97QxLBDsfYAfpI3IQTdgMaKDBk2k/4
h2oxx7uuXGM5uYfWYs/iHZq0p5gfX2oaoElLbB8OY/drjRAxuOxrSAU+wd3/hvqyB/stBGj8L3k3
cValYUXXOPSNophnQVMNff0PWzJWuItK0tA1baCcMzZyBfKi4r1g0afwBn4U+HzsH6pxgJIwiuCH
q3/ZRp+kC0WTLPdhEdWrgnSlr3GMIGMDTi8W8MIq+P0QLRs/ELKt3qHd2Rm4ujMItrr1trXuZyDL
l2k+FxfnOv8GukBzoovckAyKO/0bbJ7QOgqO1heH8y0B3CLKnb03u+rV9FNtjbxQNmPHfNMVqY7p
eUnW/gg6g7TvIWBaN8OVhnsJUyJ2Liw42eypAQ6NaIropUpxF9JM7ChYjqpwuKhjOBaBMJyq/tyw
dn/pOBaD+B8+HIe9tABlypcxxep4ELJSrZLeJiNBiw5nRIsuWTILRSS8GVtX7lMHcw0ufyzIwb/G
Dh0EUQrgXhYL8ovWTrzDOlNDnAlIcrtn/1rdN8+ocVYH3fqHDq3buf32sjliAcRVmtkqmTCOX4Kd
7C2l8aATssIrAZCo1EvKWh7yxnICR966jyW8KRtZ05AqD6bGCvZU8HUCCcEwgJXN8H6fwaxO5kwG
eiUMfbiy3HMskd5XJwulUVZb+6Dv1EwZNQ1nVOKMGHtXZe3DITRhSM2BM3gVlKEf+qxv6rckPpfo
9muJXTWZ4No8cvEx6qyE6zoT7D43vwvl2YB+1wPpzTLrjoeBnRe28Ba7R0tctPbP1e69UXKiQ82z
6O0TJ9LZVr62EUIblef1g+gLPe4YOmoenDJ16pkzWCbDrrnpzhzd9QBEcu8gFsAc7DXFFKMSULhR
4Aaz9g9roWBzwrVWiQ3eUKHngToLndyofHswmScsFT3GiVdrhFHkUWeTGkLtXm2vCgN/appwGOSv
PRcs4lOBTyFnH+oo+Lr7XIpClHYPRWg7Fz0YU/w8dv2ERMRqMAyZAHS6IeBheb/IRUbKie6c23oW
nm4P5cE0EmQ0i4ENg2BTu5h5iu7xfDyKc9bk/UmGjrywFsBJvMtiQtLLC08XjnC17Wnr50/1s7g+
UmfNDvJm2c1QtcuSzTK1vDX7aHXCpj0jAM0jplJQMjYD7ISWOKyNGyos1CvGVL9fKsMa5IC0IIoV
f3vvy+luZ/F7hi7YyuE8dbN6YYsCvCXVFzZU7dwcWrRqPoMvakmduE+P2/YtUy3emZJckWA2gvM8
bsoElgaejmPaJ1oFRl81kvBXTVpXhwueoeExd/9Y6ghHzbB28zEPJXMIxNes36egTmyVCHnGiA6x
EVPFL5v/BYmYT8AQJr9njbSsIZEqyl905vXdkCfsjBkFWnuC4fiEWrEGiNqspAx/Fbt/ot8S9vii
Hmrkm6eZYAgliD5RvBkF5ZeQin9nNvYt1vqOWcRLCfI8zwCU3FP/4PfbI99MZxjqrXRAnXgZ0PR0
AVpA5ecERYo9on3Z8LCZ1z/8tkwtG8G4VpgHBDjQpyfX3fxqGTdhWV33ja2LCo6RQylYP5eJ9X0h
PmPyYVuZk1ZICBmbc9nTHJyjK0FHHXZc2sH402ZcXz9ktrlr08rpFB6EwfVw/uGhVjEPnzOTJMgp
JMNg9825hH4hjN2hpxvk46neA9kjsY9oLadOaaQpMDfwa4qk43m2mEkk+Mz2HM6Wbx2M/yHX8vAj
cUhfIOiwsvoUAaC+uEJEBhLTYCngNZtO8rwrp36Ex0197Ceba7JpICuiUwlyYuxEtCSI+zIc1uN4
tdiE9vDTCX1xeCUa8AsyQ79NJMvn6oBj8vr8WWIhPd/0/oXSFfrokgp+CIpIK6T6+w/VUeWKq1Fx
kHx4sxeP5RQwItlmF3NWM3+7aCdFbOFLAapo4q8ryVaJmavGE39622sli+1Wl2ftbpdqXbpuGP01
Nz4HGUYG6Oua6CfYXr90wm/meynzFhHk0HMGIfLuOPYOFxroR+lXwzFIh+fHMLlmAX6bWsTO+XI+
EfIptP2WbI3ghBgqmpRtLqe7bDIj+oFARaouplJAZIHl11IGWxqChGsxGh9x7BrUjmnIPb3Ose32
Euaz9SbjI4//qOmJaUWMG8uK/SCSTP1vGLVbGj82e0EQ77mc1KmyYJwmAhRIRBdg6BwxYmlUCUD9
9rLFvxijox5NyV3dyJPQnFs4sB7twWWIQt8G4+6frkFAW+661YQoT9AogDPOcKvH0J/NQoTXjPpy
Ar3QcH8+GyO3uGPrUy5KZaUg4FIq6VT21PURpUEVBuH5w5nsR3stLnwDhDFv0F5CN5oOaVHU+bRy
eC21ECrvBN5BSV0KJfu06cOjr0ehr5hcXLTVng46ATpQj/ZWMtygJBQ6ErnM/ckUsZd7vVmixasm
v1lyq88voRglK0h/KoiRLPFR/5I4J9U0O1NiOGs5f1wFMF29Ww8oQbwMxe4PqDdIWm4eHbrVNgRe
37C2yABr3xYRnVK2OX0VxK0G4qjf1Zn0q5iH47kq3lvwhM5FW+KJt+jZB3IRDQu7oIBQrLycnGL5
tzTeIRxzXxBBIj8dUuLQ5GskZEnmx00suqdhFyuZqbgXteEXE4yARcGgF34x07FxHTmN3/Rc7uaR
3gLZDP/648Pn/iK+KM/bVTpwe42EzW9woCFCOrZqRusecSui2eZf0jeU/AiDTa8pqFBBAcnglOYd
Gv/JhkMXMUYvpohKk9UU1S6sK7PY1t+6js0qx/2MqmfK0DfZ4g2kq6dJI1jn6ygZLcmq6UXCKJd/
amd8hlhtXNcOOrhUkTKfz3UTla83Pa8d9xCq9CDmW5PhCll7Qs1xk81yne/LgGc0pfUA9zbpVauR
ccL6FVq+A0ZMMmNWUqUDpo/Xc8n4uZS/534dwwSwb3S0fmfUqfcuGeorGLJsXe+HMedJOtILyKSd
W97j5JjW0a+ewUwMpYb9Ql1hOrCnaRxZ4Bh5I4mCRCHlZnNf0QIGcst7A8yuw6cYRzD263qDzBv/
IpR9YMoMb/9UWWstSqpcSsYlneJufNU17xd/W7mgSYVUyqdRqCxrqUzqlviFPiC5BirHMh5gSNEf
JbXbAKihyA7e60sc0v+E2QgJvNnAeJtqURjh1kbKBuhTiJ/xb0uQtoAzoAt41qFMXlo4YEzSQ6EC
0GUdb4Z5IRttC3cH+wagFQreX/a8/LiyDAt/V/1IcNL3vWCl5KWI79drEg1STClSTGdiJvUx38WK
utWUMfkQ8TTAoetnt5yubERRAlyoDh+86tg4srEzb2EWCcdDKP3H/daIsgzwxjPmKO0GprLQ2nN6
1c1FJA5VkbsRUXMg+MDNuDb/BLyh8xXwhb6fmnYtEDW+jkt9PuKeokJ7u18j47cF859NkMwH6kXs
Hqbur9tls/hqC8En6wJW+4qr+QJ9B96Hh57NMc8mCZsPlbtUBQMzUpspOwEKPc/u5U/FmAsgRBsr
pDzocxd2Mxn3BukShaoBcuXnQLU91N/jzFUHNhICSsyasZRAjS4s5lJQMek6OgKMeMdeRwou7qO6
TxLLmuwvoHi3pJPLd3Cr66+no6TsrevBtgxqnwkeXaAGrLaEXx8jlqbVP+gJMbI6rbSFBbQormfF
EoL5y4+EEjL8PqyjB8q1/ve1ajkVHpBZ/bI5yVN1SNXc6qpkoOCgmMWltTDZAZBwD56x/dmJeZSH
n84/LjNabLv3F7msefL8fFDDq6PlESy0OLB1o0R5VSwGzEcttydzjNiUj210x81V0O15rVwLVoxs
ojGiti8ctUG/hYDltvzrvO+S5G6zwY+g05WuU+FN+5gAhLUpKRkyVaHELuMgtVBf5IdtjPeAZtPm
JOQXhNeG6beOrIcEwgyUm0cKJHKpIOk5xqFpA17kKwSxd/6EjBcV8yXLVcB81l4F1QjL7tRTxdow
CwnSwgkfFRYrE0blo7CKjVEUHzSpx3LtLTswU+bw6/dD6lmrnrCIL6JUYOnrfrdh94BgQPN812qh
CDLu02Oj8spx+ZxF2fhW5qWVAACTQjc1pkU08A46UWWv/vKFqDcfcpFbMG7cRrPlWD2QzFX7xOX2
G2iTwSlrAcSzCAhZKde5dW/komn2KAjYNtLqdhAKmwvpE5Nk3oOvjsfCxMC5LNaRrMVAkHyRIsId
fl1vhjOzsxzUXI7G/a1SNH6kVtNlmareNyNF3/766iXh9y+mh/LH49Q2hIwaARK6GxCHcvcIstYh
eJf2PAj1VeIWfHkVod9/mhKsSQkbkiMChR++ViLgkuaLJAKYjNdToaCA9Z548L5BQ/FirKbvu6GP
JHlYc6i1zKs2Wv8vQyNEoOIf/CRDRQmWAWQ9hXX6JNHJay4+ou7PyQq/LM1xj8cEfn93qttqluld
V6IuW4QQ0v6zAJe1K3FeMFc3OG4jEK7qA/ZwkBiHJSv+G6ezrj9zVdxWw8deKupy2R4A62EiKp5F
Vc038OFgsX+PBCSW9clMkFMK1DPES7Bs0Nla/kutUv817i/ric0E+9Gqzkv+WjdmFOtxLYFoJHJJ
+UdCzydCEC87E9XGPm8Tvwd85WzTszMG/NUF1n6FYCUr3innpwTx4Mja40egv79sXtG0ozy0O3UY
W0JGImT0cdhfSeqxglB2bGayXX2t5O7is7sH4n1oFEGd+ILifWYvw6riZRXXE8HQGI2zCGRUu3CM
SgZkWGSUwNQv9F8cNMNWWivcl9V2CXQU0+LLu7NuuqBRQQjnoBvINl17s+SrNARfNZeVlVIPahQq
wPv7P+xYbPXuJyfDMep1cSmzUxkU4c92tQ2WZUkT/GQoCq/cMKXkpKsmyB7ppa5BwVLRePStjgb4
qtVGjO8HvXngrZEaHvYAWUVSrhwr1UC769Ec4MJJPbOOvAweMINXeIw+4ll4Lbpgqu1WXzBgoRJG
RU2m42Pnyg3cRQfnJi6ygKbTMHenQiZLJpmvZWlmieaKfxAsi912LM2uWn7ddxLOSyr3XK4pA41l
Ydde8Z2uu88CN6skq5D48BKki7u9nJzAtUzeqPWyVnIbmfSQ8Kx4vARbj/1U+NNPL2eszvu3hVCd
vNXYXpWC3VPV6H1oWyEpgO1djpuslWgrgEpY2SbHxdp+q4EUlGlTzqDhPAqYSAKJc49F/77/4VC5
k24tfG4IwWeCXz/mIQo1V29/jx18AQ2HJaAXcGITRdNxwX7TfncOK+ToW/Ag4SvV1+G2gs0U6TmN
XRkFeI3xenpwni9VuPdXYAVJnwSpE1lyvK712KX++NHfQmAUGO+XkLgu293/9yD+6Ywz/+yIvkLX
AHe4byRW9ypQ/6RNRtomlA5KN8RNnEu3SI8YZqG0UCB6TXfVhKKhSrFUwQqmEA2Epj1SEYXVIVKG
hE4XCa9zRYot/VDgYuzbO/mhrE525veVmdu7VxMr8+aOmn2Nw2kUVOZBlwDx/807e0a+2FLoeE50
uzCLtg6HsiUm+dyWGGtgxkFg2zgSxXtA2+wJCuM+RwH5nBu5/bhq73CKULdaUlx38dY5DCAHVXg1
o2F02nAlr3MPTCg/VeOrWP+J8yFEV7sH8r1tC9QKHHoXyMK3yu1qs/q+GP/mE6UAs90grtwXbzDu
tlGhuft3EInG/TtZbL7IcENB2gqDWeC0CH5fYwbMntdPJNtBnYZoCAQwlbf/oYJzVeYJzD/si2Gr
zBoBQRmCsHWs9A4DE/+SpEMaqo85zK7faSB8/63yGa5jEUBR+A7kC5eKHjgwVz5SRRocMJeI/cUw
+JfefXL2z417ZJb9JsRwIKYiZpndSuf62JGmOipgxPwWl557RJ0E1FW0rRLIFmFpd3EUD73XZMLd
SrzxqSsxy9EafjeHBjWWRUHArwBB9ITJoozREoK9Rx+A1tJAdP+T9sonX8Nhe62vh8Tm2ij+7haw
Vv0t2kdRhq4/wSlx/nsCX6ZfoESF66E+HaFJUZNEIq9jBtLj33cqDZy/jCMgx/FwPjOufhLJyIvM
7IESr43d6k81wOcPbOjIToHmbI1HUszW0my7RpQ0ig7LVnBFt0Xg83qpKAUFWshgU3HWXqlErlp7
+Ln77CMWJeAd8W/FYPin7oqHGRNRL42zqCpu5NZIUkrutY13NGMo4YgbP/+OpGWb0OB977LGD+RB
4L/2QNw2BMfN7bd6MC4KH2QNMn0VwkDnkeKwNflCRd6kwrGR9fLmZ/6nmw8nf15HHd+2jATqoRdA
R5p596B7zncOOaDflcDenIasNsP5/1NRske+njXTbozDUs9k4GKEW5O/VWhY3c7cXkcM4sTABqtZ
ICfpAPWABuj7bBClHJCh5AH3mbgPgRxbwwJw5qSpjk3+o/UNIixdgdkbe1pBopgPThSTLgDTc8PF
QXLY2l4rFOenOJCWCrAOvGbtN6caYyZGzCiaR+IGtEmW/srg64VXw1zxS8VsSW2j98SO2D+8iRxa
Dr4XMC6OWtPqgeRYIx8keWmcVT6wbhyFasJ79uQfmd1ucaS58/Wy6wZLM1kuQyvNSswlWR49zhVQ
iC1Oo+bXSLobz0tGmFuv3fivxxF9Q9xZde/GGbe1tsbJJawe5qtmE5Svm8sEcG7O+2RZiwJMXGAz
525wHDLqoWlgQcZ54YY1mwJLqxlLK/OadD3mghkbMLnDEqXY+tkZ/Isu4R6ir6eSPFdIz6akBE0P
tCLrjPK7Jp70mwf+C3sXx8pn4R7+I013dT+piOpiGvk3XegiTpm1TgdJ3Duw9ive4k8R9qlznzbQ
NZCB1sq2DXOGVZMvXdARMwj7nOnEM2mBMXq+/+4Gb76E2sKtVLJorBGav1WrnEmAxTTwQMxCMl5r
lYE/8ANJ73+DGWOj/owsMLHZTGenh3DckgTjVZZH+NXv5h3EETL+gmWckjF/hBa9ltUslPsgNF2/
vmLGv844Z5b2SBZ0TaSSeYZcFWkieT/jtF5AjYHOQAw1RQuI4BAv6zZbYV805ZfHFhDDVpk5ey5o
Z8+Tiu1xw68KgPNMBipnJj8GdFi6jiQQ+kGdCkSgbtA8hxmUIGnskJk7RIVj4ykSlsWdenGAY6rP
yEN0Ix9MysxPLP75NnGnwPPh0wXZmosLGC4YeKy9rLrAsQ3Ja0KOsZHcIQ/vzZn+giTv+ItIg7q3
IV/U5QjxOdSC7yc+7gJHXLcsoyQn9kDYp5jx/As4URMam7leQjN5RiFG+BYH5kGXTuVlAyqS3GNh
hS3zTSHnttKlb1/xcNy3OWGKkHhfMpmNT7TR14Nq0RCWE8952qTPfU3K0A96ve9ZMavss7XHjSGW
jezhiZpdMOwu90TDzvrfV9zYtnvA2w8dFt2Jz343fNQVAMS1GT3EFvyOuyL+vAkSyF7Ube5RClJB
bThilggbJV09ieVvQkq9RFAlxhf0RvljQZsSVO31IDvAjYgQcUiEvZdgchbJ+Ecewb33rKYle/SE
xtmm3tnZNa97USxXs8nSjCCDRF9ksRDTpl/778S67PpzKI3Ejg4igTOY+OV44CIAvVp+uW9j2hPS
1HTOStFLl3+CBjB01Gq1QB1c95zZP4BnQlTKPcmPIF6OFoevzMxqEjUcmWAhxJAhAvOYo7pPDmZ5
nwwlccodWcJikYGVxA1Y2aF1RZ9MSviF57neEjDAyWPtuL/yFYpl/sYqXTaqZ1uTC9BXMhn+ePNi
MJJ0IYKRVlvBZDciNOJnwHgpJiOfPhjn85DaM/8fud/BLJnKBTsJC7ScGngKzmMjf4pGMuBopNxu
SPJqPSMRbZ7mv5blW1Nx+DzPBCQ9xp+OQ+yvmWZM7tC6DpfYf2FWjKMn1yJuUnWGZUxIl7YCUa5t
FNfClrN/0W0aBbQNFSu90guCyLcpTmjMci8hdkjgduEqDco9MrYdy9H+cR0yk3Z55vjh2zdQknsx
CNsH8nxm3vEYaWukI9tMF8VfiLPOTPy9u9AuHFytoeuVt16mtOIQqEyAPgwviRNOyDn4RsiqgqDn
ZA4gtMhT2+a8lvFIi6JZ2pU1TZiuHKuBPLgkIhSsSIc1piJsW5BOyyA318Mw20leRPlVpc27c0U7
wiWJS5F/bH8+4693cs87H/oCSibwxnqw3hUCGIj9XuINS8B3OaeeV6DqK0Rtk9e5M+frUxXGD+aA
0gQUwHNaSJ7uz3g7z/Tv2PCoQk8eP9XoHRIUxqgwMr3KAjH1wjYl37rSz68JeX31IqMnfIyiRE8k
s65X2uj3i+hqgSvmeMkpsJyL3XglHbZzBIUiGbhOr5JXT9q50gn4PlCz0HnHY0szuj1lBJOWVWUJ
Dd8omRNmfO/mA4O3YWWFj2NdXD7Zqvacppw3EBaCf+5mVA7zpJE9C8FcxL5LoLavLy0BkphiyJcL
8W19THeO+qNEo2pD9u6VpEisOrJSRbkYBeuuzmyr8sENzc+D/6mOXXPcyA/lBqd5sPJ8lCOlFuzB
+Fz15XuS3uh3BeWT0NpfP9rDMPld2fiqw5CClmSiv5KD+LY7mMcws9Uip4rGASSYzH8mT9mjOJQ1
wcbJC2Isci5IqBCu/gGWFdTtVNwujZpBwPX0mHDc1z4mD/jxcn3m7zD6B/aC3Yve9RZft4X+b+fH
sYBUvDr160dNLk45PhzAXxTAyI9zctb05DqZJ73HA8QvK1pQp8gNrDw6qQNd2baAoqeIpahvl2nF
Kgb/FZGVR95Dk2DvdREXVHunQ1rv+QYyBfQjUmDQ/hzYZTOAg8W8Cy1sqfagGm4GYQebvsyT4acK
5S4K0mIpVmDA5D8NvedUoqcDbnl5DKhHL082PsduPojPA8X2sDtLkLvOZFG6F54R1ffY3txspOK3
z+8vitVbWhQMo6jv/+ORYvu9H4LnB1cY4OYTacgyPtwzD5yvqcqGGd0RwuUfSsFbUaIuckJl9kis
aH9DBQuobj7y4+r+CGsteTtSp/pCAdi8AR90TAcz/juEZmXgw6w+2Hb49/4s50z0vVgmPWpG7nMt
9j9VbSBblbQWMyMYARJlsHDev40t6GjNnAtYhojd+M6so2JgRHOgeI2oRkX5vUe62Hjzy+MzsJg3
N4gpXh1xLxIQ2MJSmT7f9yYyIJNRO5UcNMejc7kIMK8rD92xQApoL54ddnwlygDcuR9Iv6g5Abah
txPn0GaxI+mU2UQu42swiUuI8eXio8AYrPw8cCKCShEWqv48VLWS7mFz+rE/nJT/RBYd6WNu5qsZ
HC2TkC2MPYMqHZ2cvB+3pvngpo3df04qzI62AjOLLLiHXi9fQKAPiZUAarINzpbEtRBGNT7IQJ3U
KWJuUjF1MX9g+TRSOriqXTEQJyw1vVU7LQT7WamH5xsUhNkX8VFAl5bY2wyBj6k5hjGhdaPE809+
zqeCnm1rUUAZd+Wk+BIPxkNIBtsick2GjTUi4ICDhjxiT7aWc8goUcwD5vp4gK7l6Sqb60kZ3tUD
1TW3kdhjw8w/wERRc+8A//21ET1XAT1TOsaof9Xttf3Zg7cZsMG0QesRWVBpBjw6Qts4kOGqeuLO
Oz26y6X92xDw6hynuZlCY9YOQTQX0ftGht0TIILN81Ae13qpbHSvb+4Vtnu/sNqy6IepOHdbNz5h
uPcB1dTlVokdyBZznfW9A2kxMMTLK0wuIBLOV2pdFy3sxoIlvdO5T+JEPrCpIZNaJ5q4XW85RzMX
QYoRRHJFs864KN9NoPvTsXRcPA4iRqHlCa11eJnSeEgVjIQjVLdwTn4oiM4X8jcdqXnMAC9Owp9A
mhA5pobRJEHkEG3Isj4TdODT5mq16uDxk+bJl2dvQzbhRKenyUKc0OGhB+ITajQ03zsUsQN5l9Ad
CY/Sy3EMyuEz6EFcEC7VURzylwkw6jGC/BaxZNewJmq7IYMv6m8sBlmzCOtDdcMUL0mrHWEXsqEL
k5EDXFm+Ul91ARWE8D7/VTvVdSiKqmuDulUoZHvZavW/wnPHt0WPCiGoYB9wNHhyglfGrsUXjoZa
qPHJjspDAA0IJuU/Rp6nE6dye1hjxIyS964al+Akp9HzqyzEhmarWA7jxPIDJU86L3+FKwKCfWjT
Ib6EUI2SHnJz0e8I1fnOTp1hFwaFrPIGYcYjeQM6tgn2nf63dUlrk2wcjpE1nDxcGEkMdYHCDrGV
rYsmkuVBcvmDVKsRnLaYOgAdV0n8UWSpdxRTgUyfTUljjfgMEodM9ITIXkKmnYumg49F0q1DgRxS
ukPDrTXWThFetVfLLzun2ryv74zrvmtM/3skDK6Xebshjyq75Ra7hQ8QrcRkybGap4v3dkN4z8oK
Zi1kbyG5vCyUx5zIULAbJJe2HGV80tueof/xNxSX82Z/d8i1+OgHulm0znVq+ZCSb4F7aRkGA0DY
AzoQNbPBR26kqYKPDjFtnoBCcUEs+dByXafmus7mIYJXWaPNHwhNOHZk/lSHNJQc+wVkKqdRFPHx
9feJxqc1efpHhY6qqWiOAq0oJKqfcS4aM+YlLCbKWkg0O4E0axR9yBhNeyxWVLPXIn+gZszA4NrG
dcxMUkoR5HID97gWpy/k5oGpEpIN5zhh0mPxRAtwpbvnJTDx6/rih9PFAQKY0iiCRqdQ4e1N7grq
vvmp9HEolwYIajpa1VTLawWjbshER8G9uFH/tM0ruKAM35lXiMQpf0W0JfVN0BmatRalOniGxuFb
D10Z1gYmNY61gtjhwEg3mL78qTUpzwmHJH7u8jSIadatgNInxqkrzKA/Lyc3ezSi//R12tDlgPn4
j7otJ0wwANPJ4qBKZMszzTV3sFbrOCUF0tugbRPQe2NnOgXR2EhcXrWSxwxda52HW+F0xGzr/dsT
41WROPyFutVCfO5ghaETol+1OCqy96KQlv4H+wH8rDAkEEGz3+s8/DBKpWEcsDuD2Jx9TQpdz6Mu
HrClDYJOYPey0zizdhjloOVz9DGkp0szYvDs0yWDPwukZpb8btJEtbH+GD8/xN2B6+zYybwbEvaZ
E8JNe/b29e9kuj6PZ0XThbOVX2jGDhqvTVzuWBixUxWEjufvxsvFK/l6tuAHY0iqlepVmjWRBkf0
l96q8w2iDGxgW1iSDlLXyplcrOgdnrtWidgHwggCLAPSvuGXqw563W7oLE8TjDL3IJkC5G4HjKAy
uNAxnviZ/7vfDr+GzUb/SmSw0D3Av4v0YbQe0Nk9NKSDP2oqrVzrU0xQPgCiC7+MyANF7Kz29fJI
xfsI0HcvxY+Akov7DNRIDsL8C8hpaqM21zdNCbdzvGu0FQhGeuI+0JKywfLj1mwdN12yIFSjIgv8
XoVxRlvoO6geH9BWEHdWy6k1eWuQFQrUslYrQGUbp9ETGeTpOxG9SCzHnkgJx5tPUppoO3Qj3cG1
pw9d3JDYeBMh68xV5sFfJ6HHAUtDinKZBOJBoI+LqnFNdZeMKQGZZbzhLiPgtW/m3bG1VzdJtFVi
ssF0bLFBudGtxepiJhkecCGM1I1Hdm3P0rKcY3I0lq34Y4AhZJo5lTriBpA4kedJ0Mg4e5A5j1t1
Zr1oNCIFQBE+XUoSpMslxG+Bdu0P/B2z9GjpeFzYq115qDNGuHlAvYX6dqNTgx0NCfv/MM5hU8Wn
T8QHwWjYUlkR/dgBeVostNN7nMvZ6rsYReWp/j1kqW5T861PEncTo2EijE65Gk+f3yqiCJ86tbmS
1heVcGH+f4WWeJ8K25pkVJZfFQ2mGXTvKahqETDtV/thIhHBf08SXz5YfEVIPUgOh4h7whOMiDnt
yrc7tEjsNaycRC/+XVX1T+d8BOlES/HV/BwSpCybfixFzFbaZJ6+A96fH5LMwBXYC5rx/pX7YCtV
o5OHIwOGmxJ91yRwWRi5eSw5FAZ6h0MY02NvdunSVDsOHpwuXz5Yv3C/3N60hOgeW5/nOgMnDFf4
i3YPkbzTi52RCvTs7QXFdKJRC5Vv13DYpUqIBryUmfSwrWN/9VxOsPZWAI6Wjm6ruw1O2gh7dDqp
u9Q1gv/jlXakErGGo1ZVJVu5kRx3QVLvxb3VgRmhM9KUTH4aSCZ1lc+eEJU22WcRgiwmD5mRBVBe
Nud8f8wkrlchTYCeQWIIE5iUphSt0rfgMqvwkv3C95bDRiBogDrctRrbQly/+s4TwcGnw95hpjVL
t59hqfDUteKYITEFnvno1qYuSnPHoGAr+P9bC/6y5wOVdUuadExpqU6IjksByFy+bdJ2Gx2mWWx5
2LaKCZ8KCwYdW3OijR89mRKEnARFuvlGc1q9+ZQVIAHuxhUuwkwHTRw+jqgiPLfO0uL3vZx3GaXm
1XytFuroqtVNxLVJjGJOLrWfnE5+6vNrzDQ+I3RjeNCsYh8o3EZDO1xy6MJGEHNpjF+2hfIx2MRJ
+6HyBdmB3Ev1WlT9uRq32kSO2FeqWKVC+N9SMN5XQB/P61ooW/XgPxwTAiQTh3sogmdJ87x+PTtZ
yP+RZcr56MI3hbevkC/zaMhkQBafPUzwO52FJ+i+9DpROAMGnn/RkIEpn4+yv/mUB4w0deuAHtgp
VdtP0z4wTn1gn8r4nZburyh7ZeqXtdsYI57CPAkNA8yWp2M/OkCXlW8W22LnbLe2HwWYDCsg3V59
O+ScytsrKWTQkT3r/1zw5asaWw31xgHkaiSkH50oPA07/Q+Dvtdz0vumsr/sITO3m4y3quKnqohx
8lRwdytmhGHkcJbDO+maT6wFLTB3WMwzW8E0Wf6ZbNKZxdiBqnYuT30A1KeJ5LJcRu3l8YZsICho
MDLbiUqqKlukrqKZee6rOqD++mDj3xQD79kOiNvQ33Y8eOKNsGztMrbzX7oGtNQNlh8nZJBetr7H
76nEqHgrEYZYWQWYe7KS9gs4N8sB+crrHdJ/ABspgLgPIdnDTE3a2vSnaqZZi5VpEwaqOYbhyXsN
DF353MLfQNcXloInO+sXrO27ntIBTwoEgAzpz9vWTeXkVP7KoVdVwA7bkFqtsZKwzyNtlLDIqLbD
0czGy0k2wcSgA8kE0XdsAH5ULN2sNt/p/RsFnd6qdfUMnoWWFG4oNQ+7rMJz77uFGpy42uw9PI8l
VflVnXb5j9qv6c1BZJ0DA3E+hE5s/pCctpScgKxwXLvStixJyZ4r5o55mgwDigZ+e1wTh7YgeCts
a6t6eU4uRaITfedRI4Q2Paso3nWz1tL3z6MlKklvaPjeIDHu5yPxNcSwuae7j/dwfXXq54zrtXNA
yPcSdJyciIcBJ4ct9gJj73LZadBYFSQZ/QTyW1DNDur0yl1fe83ydD8KtxO14CQkzlmG6d0MKw8k
Ea0k3aQxQiIWhKhYMRpEeU0A7WvSnfXW3k11pjG5PX7HHJqYOr2FiLN28d846z4EamgWWaZ4itc9
9T8QA/bBMsNALvEgXU5/5N+ysG8PrdFV9Nad8rtXS+L3teDT+cGmmR0HmSDd8hs8ocqXmynCesP4
DPzOSdvx6uCwiuDq2o5kEHhLTJoEGY15IQrVEkv50fSMMu45v7gpl6y1xOoGknby9pUtSBInyyAl
7IvITZRX70bXh8nJcI72Gy6UpWLhXYxgwv5B27EYWQABcrluHwQ6F84YdH4JkhAEkt2knZlP+tH/
tQeA4y4MbJSbhEGZcoWdwhbD17KPcxP6BkKIMWo+6WYvLpDQHf2ZekPhsKNMxVeaKOb0PPX7PzbL
XYRmJcc3MIXbSvrh+rZWPzWXlTyHYy4+qZ8m/QOqcJiey6rz7OkMpNrqYkr5D+698irmHFVE76VY
2L39TYIx6ZPRFFjDcCNfNoK7ilY41476mjoU4IVq/DVijonvsDfLRkOUqYqAtGqq6vc761UF+AKj
nt8HEWgGhPzMhG1HsLV9lU56ybXOcVu3Zmsh4KseVlijw0jpz3qMZ4LnLVstI1ecW4Gxm1SbqV6T
5T9kiqTO5r/RHc2ZlQqr5bqC/bJ0dSOjoGVmGKq2atFVK16Vy1YzyKEuiFJaiRcS35vR65Dyy+Jh
U+p/LSPE7/AkzfYrBHR9tNr7QBkOUzwRsNzJ3Iz/LpnAynEAIUhizm6f1VzOAURcd5Rio+o0KUMM
3XxX6epqhZe5mgDi4DN0CQO9LBsWvnJwHfHnSI1rpS9q/KoosVD3WbWpLtnSsSCEx86VqIFMsyN4
Vg+hzdq3sZPrG8R2ToQBu3EM4vGuS2HEnMqYOEKrBwxgpa1tEoM/ZW1soMSiEkdKwPqZfXB/fcG1
zPgVU1D/rcJV6Hd6dDa5L5Mk755bbHx446HEh1BvVEXf6DMRzxFbN9XTb5SQ3QYxe6BGYmKG7/c5
g3/UA0ktryA/r5ZyX5fylj9W7fOLLcakyO2duWpw3GB0oFXG1Ue1qu/CZort9ZRzNx4T0q38ZLCI
kopthW5XxVBqrChOhBpGRSSKAm3c6ZvIWEp7M1LfVY4dqPcuzqU/7CZO41x7VfuPIUej2i7/b7WW
Udoi64tctXtm+FVy4akMOLSJdKpcDtCqH67fuV1lL0hPborCNLNNSRud5mWjD3OxBgjGed0GZ77r
XIXyhCAzVv7JA2v7XvlW9jbbNgTD1CE1xPlFJav2aFiB9iOSRmaKjuW4mIgOdEHdY15ry5ZHMMyD
mSHiAXZ4saB1oJiEThX9blgScIN1k2vEj2xE/tEnDMJYiisK3RdthMtoz4IzI13vcZxY3tuiWmL9
g9VL0WF9WMSnxkVBavAaegQ45rdnNgIx6K4wrFskPvaPfhqnh8kWYu2vU+Btm7U4gAJXJRlFVmQF
EiCZsYiLlYDdaapjApCkwlsWhjCXjs7349x8MClISIiwGTYCI47NMfLeWJJoCTlCtpqc4LroU9hh
x/3axwdvYXTv83lOLKQ9dQt5nwufvzYuqgnkoT9dRn7Wsbv5WXZK2YE+veiH0/ZXgMCp8ZnAwIy4
FY8JAqaPda5d3xxoIf1tJnXZF5eyovQ/uiziimeSbwbZq8PyfMGyg+ig7pbl9zrfb+fmgKxe8dz7
W7mjmHO9Xlg2IFvzNRgRkI2xRtC9hz9KsSgjeJ0zk3bW5SrhPxL9f8L84BNXLFPf11I5R/TCtt9w
xxFN7Zn3KYowupJNvKpYP1xJIs93Pjn1/vNZTX9IPmKBorzhb84mu8BGD0T1uVBkZ1Utbw+e5X2m
qtGxwgbXGPJU+YAufzmJ0R3SMqzdvIyaWwNyCbESQzksvTPSf0VVImx1ToeRk150qQ/OwhoOJGB6
9DYGVcXSX2RUyFOdfQBc/23B2oCwAwceSdaixvD3QoJ0rU9aO4xBEGS/bgB5aYJX/Q9gIstJaVMw
dpjgnPzk0OBlzo6oItNMD0RCf18IVCyjfHVVMpSouVq9Bf2keiPEsSYIX9UYswrweWFdyD6s4Mhy
3dcd1SESvAVt2/T6r4FnklphUXRJiHEZ1crAejVgVvR76Pm6LxQD1LLrMCbHLReMxen/n696znOx
xUDDcmHkJmBD+T2CIxgs1jLXjYRsQvdH8YmZxMOzWYPt2vycOfOb7B6Oy0IENpGDWFnEGTVsIkHs
MRq8btN4M3OCBHIQjPOXmwsyS7MIL+kb5xX1XTHMKKryPlfibwiz9tuf54VZs8zn2A8mBS0yIOtr
Fqf7K6Kd07kdl1EfMcqAmLsOcqNJvReVzrBBk0knsna4dC2GhYJnpneLcoGBsDHdHbIUCrG4i7Gy
d2AGs7D2ax3GuZpDitSzV3HKWP7oElYYobPBeDlNnA2xuTE+cKplOaNjoBbnaK16Oo1U29smRL0s
KpaaCkFZcqtaZxPxXBY276v2ZrhNdqaLodhZTA+o2aQxkx5/KMYPdUVGok5XG402C4Nblzsx/Gs0
NB285HMhKFRriu1LzWSMGruAUVRrgOdiHaiuYB64Y3Ni8X8oGyY+C+wPCqFPVXprdzF+X7fS+Dys
cXQtSW0G0bF44O1OBXLMl2FB3D3ZbDs+F6GjxDBqbd/NOimKkDaroFYexbeFIZRqO2KKb75AAOyG
IfHm60VdtPjdVswDHpaRF7rVLFqDcHV9MZGhm1wGTNpA+fMKPCBXwp6YzRBTwiw4xPl9s+ixDDMS
Ar/tDmmn8pjqKMLwe/paXKlkLZFAXaAnvdw2eklMc3lCMXHF5bpEimZn3ZL3lzfuTIL8e6i5zM9b
wAOeFTcD78i90Gyp4Z50k55KPDe5YriqbZFgvZohvLtfa0eAPPOzw6IXVVdPqgNt/1MmzWDMeT7v
SyrAXtBLjLUlvZXUFK4fQTaiB0zPi6nhc3hjdi045Ke1I8J+awUHGRkdOHCPenqigUT+23DmCAc7
wwgZWoCmXnqT1a0AF/KOmbEAQeDBS2CzdZaHVm/bpV/G8Ycbzn5/eihLoYfjrsh8sE1wYyFULLmQ
c9WfCjB8EOyIVPdnKhEWmvt0EszY0n+nnnVTR8dC0N5LcgPuintw4dYe/CsWzPbDw59iY0hFoNq6
C+rrIUYG6Zkn65KLUohpbcl+T4epVE5uWMp2f70R3j5bBfvy3H8+WsI7YFN8jaBmT882J7FvCOBM
rkVewGLkwZ1vuNH4CSp64dAlavcVY1/Mx4PJYoJPtnqnfPiSi13dx6RGaWMqpFeppLVrYwf4cIME
Z7dONEyxgaDlmH0oPXde3ESQ3WMCH6ofYtuYF8enWi/iDNs21OtRfkWOqgX52DFirmA70RjOznhA
V6f38n+EdIsUI/H4jgSqjf9lijaxkS7Xw+/FxZYe5fp6z6WRYtWzU45QDiOD6uEZUOt1u7wG3itV
yMqMxCIxVJwFcSDSiWGLBvVqU008e2gMgbhUAj3zn45JQFYKiMBu3HD3cw/R0XOIAvQ84NyoeGlC
2A8WUbKVLp9djZplPfFfKiYtYvBoLRLES9ArKm1m3PJ1+yW1PVAqYCODKtosgyhDAA3qC5zLMgN7
I9HrsaWliNj8dsUwd3DYvKFfPwiQUlUzsG8HqiVDS4ko14aiPhdhSTZ/8CFjQTIvHi3AwDioBI60
rQnRB09N2F8vRuSFnLaVRWM3qH8MCRlqTB36Ya92mAX/E+zv6yOa7doVGG7QV/XBBX8uqgq7azne
vvIUbxPHQJJED7bfLGICVPPDMbvnsLNKZ9DVFR7meaThDwLTicQ5GbIp2WrQZnep5g1Rf70x3LAW
KTK7QsE3ZIQAokiGQAanqpBtmVm3+l+aUZZZCNIP5xahCPSJa3HuFQ+Q4fkusGtln39KB55+5PY8
tm7yXah6iKa4Bdnq6UaGPRcmDMd1h8kG7dhP1zUxcQlorXfRfPt60/eW7ByJfu70TarPUvs0XaWM
ADN9Oh40skVQ+25DMSMpfW3/JhOHCRN3FXvNb9xkA/DUlzMUx59g+DkhnlFOzt30Pmtd1I+y8bDP
0q8e0ZaBddU+rwd9gR3bBz9Fh8bUl0UdurVpyTzBw+OzGpRaomSAvwex+XXFC1k+i4irOy18lMQ4
xCnmhjwIpq20C0rQuGMbFxNrtqwf5x3AKZvJQkzI6LNHiXetwEb+RAAD/EoREYL85xTWrA0XgkY1
1hJLLC/GebiBnfRgJVf5fNvK1oeHTn+vGksZs16YEeiHrV5oHLNEdjtee/6Jx7BF80ZdQYrqVKIq
eDf8INkeAno6DeAmbaZTiOgny5UZ8LlG/9ODjRRcglokbqX4+d7HdXWCMNRiuz4PhAq89ntTkSCI
LMR/giQLoWY4hGk3tEuZdALr1zD+GdoJ/tFNc6hgfs+DkGkzisnpW50kuHIH/IxgZiPxRxtXBLfv
iNwiQ3AlkHfCVQYyPu//wxkp7yYA2zQ2mS5lpkMLB8zYY0n3GxX3ExW7S5c7oZ5CmaHlS5SzeEXF
Zo79qJYwIKqLbaiEdBmw/979JtJpTGmv+xvVRn6YfHWQk5oaG0oDlTkNfkscrWpOh/5FbmftWyAP
CcdQ2rARoFRSGHZrKelPghtYsubbRi7AvT4AJcVuq4drsAW8N+V1EPLd9gl4YtRXDGCsFgpvsAOk
zLbw2ltuS3z24yKKBV246Y5Fki3WySOoGZE/RkMSzQwVuNFbNeWifw9tMPC6teKWdX98wb7jTQ7y
vcdLKykR/4QA3GdPvlHNI8TWJXkGuKvsEkmJDOmaYpNUijjsPqFD2VuB0JVjlap8EowXuR3zefJr
jnjz4W5rVPIEGsFV2TEx4JBGh17tu2zOt2aKUeN62DZkyROVVpBxB7BFR7grUJWfTnfBofNY9T7l
/yGf21Iqh+/BBq7/U/Y95bOU3uVDUxxwt1UP9Bfp1rSsNYp8iVVNlUtspIqHV6z/KCECux9wsJlO
EvR91Bp/iYxj3DUVBVLViAyVY6u4QDF29SmNS9S3q9Q3Kpx4mmh7VBo5JO9UtcrG6y+/UbQTFnpR
Va1IhlNhspgUjk9KrDpLOm9Mrfp73uporQnJNnBe3X7sXDgkXICWYr530ZEDgebTpSRnQJsROoSq
CSIxLkqyZKtSG78hhE1xVnq0tErjQjx2qL4ZhiuKrSZVdZwvjmBdDIG9nZJcjkSQ3V+IUyqN6I8C
9cQtEdMUVj4VJkEzHKNc4kisGCUkJlLLOAMFjD8gKBoI4T5/IvS1s52JXeaIu2VfuoSHula7mSQ6
vPuv5pBM9aMkEZxcUcI1e8PrprQrUyTjxoA7k88yQ2LAxhncwh8l6LmsLIYx4csEIJykyo5YdT22
VoleVpqtcm9qBRcZGYKzTr6NTQ+dZU05GPbVdlhNZvhFpYfr0AXEXx227aPtjSMVxKAF5dIFygmf
qdK8Qe9kWHdv3gd8sr22fros+2tHVsK6oyCksPCMZzpCkrTwbYgIMFv3GEAfDu3Gvs7rkgxbarx5
ybvWvSRgp4c+Zon+PIBPgeab4+cEpnVvyNUaHUx/uFxSWfb0WJ0dcBZe4a7UbPCBdIF7fkZEAmmZ
gW2tgZRTZcZS1+wxDPzZ26omrhw1k4WtUwXbuzHCwVvYqZSoNexhdCR/i2LHcHZeZbYNrBVtQ3b7
RdPZ8Rfj/JRx2f9F8n1ZPKUvwMkViAWuswLxrrl+rLLlJKKRkgw0vwRl2MxqipGqcm3nVvGS8H3M
Gx/IVxLXLwEG0yNbViMOzy2yg6+Wsrh+iEitW/O4RcE9Rk6wFx5dJMVeVSHROI1I+noOaLvIDZb4
feCccuGyMfvxW5IReGQxmaQ7Akt68u6mFpomle8/j3fZkg7xCGty9zv/qTBOQGgUe7kAE1hw3QkP
HVgbtwAjeZStEGZHOGKR6qYOp/OevyGyVU9CJDQ5b8/NUsDKn6atT5wQpNFIFXc5MNw4JmsriTv/
SXou3M2ukQJ/n+H4qLvswha6U1j0FNMuARz4/wo4tFybYBbYyapBUssVrLZK1schKzp2mA/b7x5D
7Y9HOmKFkn4YEnRtyut5UTaqqgsI8ZMerJFRIYpkusiqZSbe7BbHU1Q4ZbFQEIxDu4MNWOBM0IY5
mleslvniwndaD50Sib+GJWk8ujcEhdsbtIU3JJ3sPsvahKWBYBSPogNjqaLaTsV+rLtHpZrg6rtl
mnbJEmO95blu+0B+EL95AdJ7h6q8XupT1y7qYZfzpuNtGIsW43r1KBKj9N277GUNl0A2P5TutNsL
iU0KkW29l9wZTPh5OG2J1zSvWmoX5eeGoEcSvJdjhcgrWneabHtMSfR+o0dj7YHIaySwxdWKnRbr
Z4g/ZICTNxewVgzRn5CGAp9OxjCuW8WsNecofriuGpVa1KEBv9d2TCC5snHtZurelBuf2AaYeVSd
TAuUU85NrXeEs6r4g1Omj3ZZaxeV9jQoh5v0W6pBUPV/a0YE2s5kmCyKSpbZHKAshZ3ORy6lQQSi
UvdWhv+UnIKl9nhC8PtKBLrgbo9bPubbJqGQ6OwxtMHbnygntGQgQEbfaqo98oElTffUieSKnaNR
xTqo+yy0SIx+vVv73sNrUoOnwjvNnxY1njDV5kNcA8SBvSrNCRjHeB8eRPxA0rP2Ad8K/e/Fp6f2
S4F1Y1t1CKVLxd4AhG0fTGeoQQ9AzEGTrniNMV68bzLKmSKpZTvar/0bzh+JFGSEu7CuMBDOk+/O
GN3dv0ywjc0F5Mal7IkYNeqG9Q2KI/yZe3IOeOS4rwJ2YrN3fyw7DOZn2uvnIWqXp5IWMSizXgCv
/D/7IVwBym4f2KkjEPGBDDHSS1x9ZdzWuYJL4cinu3ZksVbdpKjoc9Zp4gh7xUVacwamhGObFKBH
3xwxF9q7gVqvim0/i0zl6xVaGbWHOfmeBBVTCUQjxjOB1iWvMjunA6tkacs+FiPtKnuoTdXhXMP3
OnaWEXWAmb1yC2foYqf45ulsRAjG9ZRQJWiNDQX102Eqp7YCZe6fNhtlHejYp4L2Sv75l8kwIIdf
lPUnYiCfhUQWkglXKPdJ3qVxClw6rMwd2nkHVgG2aaos9R7Wu4AJLIuEx37fzDejb8/KM3AmYC2q
fZUIZxS+xuIVmDeIFikCw06t7ktNnTgNbKX1HNk+t7pynbyxXUfxTmCKLn8bfS4WeHWcbnkzw8jY
1s1eL35WRhJYg/hD4UTg441o/gVGTtH2fKJc/QhoxY1rWJFjoIncJW9+ms8sx3ANf1w9oRom1lap
2OFadQYWTjQdU8b/nORyufE4r/Ao923wFwL/wSJeNfozJxO3AHq6u1mZJ2KHRUBwfBsftx4x+vEm
58+gsVhLRTwdPV965SCkcuxL1G4GCrIT31fGBcseBM1JlN58Wn3e1iC3cys22kYhCASR8vpcnzEo
LMZ6Hxmvr7onNc0iheMH7owRbqV9AEWxbsZFmnwJTGdHmDEKOSE/ith58lPgrNlVXL4dY+5fpvsC
gg/lqxT9ijzC3p8Nt34TVP48fv3fjSP5LfH5/xT1LeWM+zylp0pqr8D43ogZhckwpmfRUzM8gLjL
f/IMIF6EZqdohC/jlFoxg12YftUfxbJWtT8znkqnjBWAHeZpyV41OjA5lhav2ywpkxh5qsEaTWip
BDQnQ9vnBvE5hlVasphdS6K+J8E7AqcLhkGGND2g5IH42fS8tM6BWR0Yuu+vkkG0hcd4ES4ZJzZ6
x6rDsf60BgMfSJP3pe+rh2VG59Ird9aglNdIzuSGH4lJ16h66R6Kw5ilgpYgspM7F402H6mbCzOp
WdHjJcQrHZgyGEZrLZHD1AWherPSD5HnIh1P2IE0mAWdEXw3Jc51XI9jBy743szWAeDL28l5WlFo
Dbj9TiyvsGbourpFc2FAajfuUAb6didzy5ST7XW7qdxy4eDioFoU/Bcy/60rkIA2Msa8Npy58YnM
ER+BtDtgZWov8KXftj5M9rYEyvLUBTUNNhBlMbtiE8mhnliIZ9Nls8ZoEdoFT3f7EFQUHBktH5Ez
dldUgb7QvbwTJKpID/Jzi0JSZvK9757OeBgEI5D8que5yfG4K0rtgmZBj5V2r81E8qL/kys5Im/R
fd3DIPYqYAimSrNbZeBTSdJi/HKi6AznCenk5dhMoL6m01jNAELcxy+eyRF5GV2F7yRmh/9nS8YF
aTL0s3b6M3V3QoZ/77qtu/TnqEnbPDhgqfeP1iyEpOgY2/U/TddWCFTf/TOmTkFC9W4iVjhuRyCd
D942J9fxwVFqg1Lhe0rusY42cTPkY4vZXLO8zLzKPpT+CLR/IiRKhAwbGu/eX6sE94/ot1eBxoF1
8IQugTOGr/va3cMtGw3YejCoJXqyjK5ApDHUO1Kmj30pQggPAEdMpYj4S8UjJUbQ8icDvQevqmlS
4/tMVrTTRyAhULs4psSF0LXOBTNpY1sWwQovzWEWibFIGa478RtLcUrC7rPa2Ry+DDO7IUsl5Y9t
NLjSFkW8ik95j1sX8AFITUWAeAksgnEbX+kUfCVEnqep46MZgdmyZuzNgSnpBE6FRyZwqALCf7le
OSUwdZ1FAE4zXzuLC8BaRoOBD/aQmoeKjNr4t2eq/7zqPFFG726dBf2tVhvAMGoJGf36HRtxMig3
/BaScD5iBODClZkWhYj7lJpUMXt8siS0s9fvRT8BBNklvAVI8c+YFEJMk0vM7/IFRym46mlXBPIe
O2SlCm0GdycCQMWXVpm/lhriuAp4GDiv0qddrdUEgErL/uBql8jI53ip5GLj508Z5zsft/2ZWKiP
hEN8Ab7Mlrib1oDKQWfOXTCL3bW72NARAhnV1OUDWsimI0xBOhhrzR2/2a4/hZo1JIDEh2Jxg3Ss
47+JI/ODpwtIkStnLq1R2+QIWTTvtZcZiMaVn02d4ecUnrHCMfuHU0270GqhTbmAmPmXZ+SAiNTq
4WMelq+1uXlQ7gMVrCxAcHdboBAE1H/YYhaoq/smIg6Q3219E2FZarzKl8U2+vo7w3zVAiMvZ/VQ
afPpWwtJqv/7s463ZKgID34qIkuw6yGGL6Th8Ist7Yaq7/SNVUtdlQ/PiDqV4pTUvzlqLxetDtnG
/xZP2Ateeg1ghrz4KWFKcw5wJkOK6pqsap/12T6a7nP942RtfeCdMmVrhhFJfhmW2l6HHugotjtN
K6lzDAVZgc/hMX32IdRVRQD2ISSLRMvor+x5GJPgdvZd/v6E0jlTioyyAcs6H0j/D+8YrZQJt46L
eT4T+eEY3rcH7SlcV4M6kStkcx6cR7HRG5XDNNhNLmvTinwgyfQzkL1XoIwWjM/lOea3ipMJbLEU
p+WXys/EscERX6FQcEWA3J12UWWcZvUeP39+Z+NNyqU25B308WMGSSEnbiV0GlH5uO8/Baekc5oj
Gxqb4vW14Vhy50o+UYTnWvkMsnZ/mW6EdSXSI5Khuy2ToJXhbrN9MlcuSf+BQ3JjFgvenygwNk6Y
mscdOUEL2AT6VoC3Qf3F4lh4ab+k6uSz9ms+ygvq+jsvgWv8owPL4ZDOM0/Agw4beNit4gizKGbp
WExnCNN36i5ThtSUlGNtZE09L+9y2NnDVMW8D1ZIVT3Phfzza4C8kgeoshLfhat5ykAfKiOYNMQ4
yWAj1ick5MRQGnE+9kKhf2iBGxgBx40Q/Ti15+okZZhJnsWNyVVZOf+cVnWQyiQOHXoyw4N1gi+M
qBF0/i0Ok+r11VRl65R4iLliP1Pzb9ID+P1MyXjqol4467eYxkaVzRS+6e4jRp0teIVbumAbMsc4
Fc+YY4rACV+LgtdqAz5dWRH7nw/gDG7rRgb7JRpixwu1G+hbmwh3jpfo9EFVg+gkZjqkU3UO5faM
Psu1q/wHpKTS3jN0E24ixWmo2l9hYgrBGmdYNFQ7/qu5XtXz6fp32++I/mJ8bruviBLxCKi5Ka1c
wPu2nqFXPKQAUTyvNuYRz6Gb/WygOV8M7S55aNXRzqvNTwoeW71v/mBJEZhHMQrEgVjZfiEfbvxr
fNABBZIOtYdTQMGlq3Yj0o+Le2fRy2s6bHChMvJYSrGoCS8vStKEDaV078qM7v+dJfJKYzRmB+8K
WjZy8zjSx4IpYqkgpbGu0BvbFykk79oG+1avdmTfch5zV0vlx8xBec3DGuAXCgszAjvEcct75smV
itCharwWg9e51QIj0NhsWtARbhFM1iDh6XHW01gYk2PFXe0ifioaIL5ejcI/ApBm+ADRgOnDxZi8
3Muxtl/oAO8K/jazGGLclB5RfWgjfZEvXTQS2+c5ZPHwCkI9eOTG++gjknolVQgT0R21di9Dk1P/
U7Rn8eGnpRrhg7XeofQQ5Wj0RJUIn5z2Jhzl58mXLqByLq+vJB5aSM5toRIvIpD9kRK1sMcPl6tx
+m9zPfv8DCd7a2AzIh2CMA7MzATAakwdTU8aEgBPwCa4Sung3lAq32Lo6CV1yto2hN2mVLMhhHeY
zB5SfqYFhhKUbD4pvkt1VSSqWo7CuDjr3OtMPoWOlaqyCxQns9aU9K3jhn4ynbVv9glswkyl63ej
fZ0MY+G+CWP5+526ZmZoJzdcOdInGaD8DYpzAZFBbOVNInDyh1wIVm/tE3Sugnw7UCLElDnF1vt6
p5znxaXR8xs98rPjbSSGB3oD7rt+/cqtsAq1NFmpW26eSVGLHSn4y0Kus2IWFIC1vy/qq7bM8zaL
kzsh6hh9ZvnMlNhlV66cM72Hrnd8RI2YSrfC/f6bjVesOZ0kqSN2eoigczV6IagE1ffXgTdvdSrB
w9yd8464GERWHm7S0Np9OAMztZMJ/aH2TcSpLD1vcHHvsapjsFu0lxh96AAFg00bDyGj9B6wJ1+A
XextKJHWYqCCk+56NUwMippHeUD59+oT2xF1qxkO9GbLIuGI49i/H3k+izEnvUXUFk+C9BerClR+
tM6bM++cSuPiasgeM8orBpRD3DDPad/yMLXuy0bZ/dCfksKOM/Q6lppgkdHpRaKJWHpHl/VfirYN
6L06e/aHqd3okp0SuObxQlzWUrIGTPZfjGiXfYUNC+qDLM/UiBmOVxXH9ZJZtY8JZ0sJmQaM3dWc
P1nW1gVJubXwfy6yQaCQV9HH5SGCZPSaVwOEEXCtWIWmNjGz0FC+XcAD4YyAdWSE9p2OCnUsW0tq
IlIyM3COCvNIqqtwr94B+8kYj2ZpkgeXwy66DplXI80jNkewakN5xqoydCawK/CRo1+zhzRlLuAt
kCNJInchS0be1SBTqlEMiwl58e7jG8ogHC6hfV4QjcYKrVw4TT9TAnF+E8jIpKMKcB3x9yPMOg6b
h6AQDcKWKnJlk8SZ0m55iPFiOif+54aV/NlmYfSiSO7iPONuDP2YYnFE4PtEm2Jfry+KHTIkSQi4
Xsezm95PgwYPfEuxVTFngKFmJuWt5giolipGw1A59qySfOV160we4QF9P1DdFj2engs04cbF7zg8
zQIHgx3JK8skm3l5AxobHSD8FEwloIoO2RFruCbxwZlriXcNxfICctFVDAZrXGS2kyjf1Clz0oRw
V100ThQ+WNNZBZbSWZKphJxk+//D3xUP+jnH2LCIiFaJ3yREiP3eIVazsW/Hcf2lPBykicqvFJaa
+lANkQ6TaI4391RD1Q1gDR7PakmJJ5axjFwgHXg/2NE6LyljG4R1pbQ8E9RaBZ8xWO8DepvZhUY3
jSWskHtuLu+OVfimi4ym2JHDVs8foODknSW3w/lhqgT29mOdloh9wHm1zKk48RqbPsVI8GL5JjXS
t8QO958ejhux3VAmheYtkj/EbHabrhXj4Y5Zox/14QC7IhUlmwMEIUeEFrI9dkV7qKiJ+0rL9sFr
P7hDpxIcI2jvHTaPg7nAC3mUkwXMgwDCl36SQGlTnKWvjSGUy7tTp0lKqOV4qZv8Nsxf4fgHtWrJ
kKA+5AsRCk83ZlYaiwIYSAdm/TFQ5VShErjIP4cmF3tZOja9IOQVSY7AS/VqsopLfh/qTMXYgWWF
bchgy/QzH+pm+m7aGkDuym2KQo8yqeQtiSTOQwaX/UvIBVAZi0vBIV9LhoizlTXwV517oza7/nYR
W/+r8bilXpr9DspvrhAbYW9guVb08sN6GfHIRcC2eVCyFDVnqAjVa5/1+GqjlnGCt+yfzeSBtQBb
+Gle/uf8vhaHm3l/8leb6pT3dOAQLVIU4nbh8j6de5SIe5ObGhZs2HuF7Q23zEqb7/aWbvks9xMC
ERIeV9axNuJuw0kDT5uYQP/B515cuazVdvz5DYBkXp+pCuwQtJdCATL3RzvbaSf0APgTmj4P2pdf
ouTfmiIwynuUmPSKOzREr/OqnC8CuRQuPGRpyMzk15fegyrmLbRBMd7USXe9nAHH0ttVruSkYzkZ
jwh1j+/FukywVdZioCDdfASrpSy1yWQyMEMrEhv+Czy2PTj4NiCPCbLz/S1QZijkWZWokEO6GZQY
C9hCZb7ol0GG5Ds8dUbYoas/GIt870V9eR9lSzUtkjI2nsojKx351+eWspLLiHZ4q3gJdS8K8Q/I
B6CKwHaYQVJpYgZAEBClOCf609oN6X6TYL7MSc98Ycg4sVAIRmwxHFtcxav1yn959fT6mVg2JLIZ
0nDvYZA77JRg4E1sEJ8NkAuZUWQwZuEOrEDaLlLhlo2go0jzFLpfFzjUkGNaFnHtOTmCsH0DTOTS
vxK529m35k5M2Z55ci0StldvsHjMWwD7e80q0EADfcJOABhIn+jr0HSxDYCrcYjU4YCSpo/tk4oL
Vzp/0KPTI2OI+Zm7aANjk1waJAdvemdIrmltLswa18aOQ+0o4jtjgu8j5tv8PQbKxVJTzaVm3Rov
mti9X6cYUf/77OxjaolI3qAwF+jKE1x0Udm5oIJqFCA2Tlrrh1aif8Owxxi6njUwNLMh89A+z8Ic
1r0OPEtiEZDtcozh7pg13u1HAzW0nx+PD+TCWS6TdnBKn892h+SaIYQ+Xdd7wnaRyxOmTxpuRBnT
qDOBVJPWNoYRrnZESmyuf0BMIWHsOMq4ArzrjWME9eR0xwd2EhqYwjMFFCA2KEIklmJj94noinQh
D8zRLEXE2/bPrLEaeW8wPPQDDBN3z45ckm+unUNLRZmEgto6uYO4C5jkaBPD8cxFPH0IDxzZnBj4
RUS2reS+ElvUwaEbp95RhtKdL9xOveZeuE1hMjYCbaqWB25J9uV5wfMF/TPvyfuQKEwjQS9BUBOX
yONUyFnfC5VnfMg0r+6niIYs7dOcNtnRY7ZmN39YdNRLc2dXkphMjs6lQYdeT7/EKhGJ1BpEDPh5
TOrmt48sIOCTu0O8BfcCTG7vZ/d08VMh8GsEc9rT2tEw2bGZZ6N/X5hf/l1184nc6JFKMnF3A+9M
vCKX7jLSBaXScY+WQzViblFhO90zKfUo6DPcBgBfSsSVhbPBptN5X+3HV/EqrC/GLzaSZltn6BrV
1xgMfPRisKXzBzm9VnE17utwyvEtZ3oTsApzHP3kq1HIR0tSlkawV2wphu7C5U2o534AQuMWb1oD
LsJdvNMhyLaxsKrCA6/bm678likJ4JwapXNn5f1v9UnrhtAgB3KBCEV9YQo66Vt0MIqRPQzWh/Sk
uSwocyB2+IgRt9At6MqqzsNrWIQ7vq7mFwAXd1JkNGw1GF9eRbbW0rChNm8vgUUwhKkgv8RG2mvY
+q3+2/Aq7cBajILOKgwN4+TJm252zZh5iARyOem0veov78Iya9bOf5H+7sSUVqxLg6MwHjct/Oee
3cEkZ7h/T42rWcMie1ggqY4lVOUjRLCRQe9T1wY/6JtjAlKK3Lzm3tqX1MQNtRXqszlxleVrBzSH
fD85kVAKMjyrdD+qlEIWUpZhPM4UIsfOQGtNR6aFomL+t8zdNtkILUl9YySMA0XI+iG4l+xcpsFF
Muxj7GsFGbPgPQL6MSM7GEltSB7OR61KyCf++HYk8d0c4o+BchChnZaV7X03wexGUfvDUzapJBfs
JUGDJ++tZTQkcbuXvun06D6817IZTX6sOCbgFFNIOuKuUkBs0E6qhme6YyEs6FpOEvON4Dvsd9aq
hYDOHemWeVPHyOIz27ygz4TzJ25V3lZgzytD+/a9OPwBbYdSfjA0QizPW+HADJ5Vdk3imujChUwP
3IggPC3usLmsHHGiJieYK59khT/H7AnLNBQcJFqfpPakqThX3tbn3nuWyEpE5QnPctZ1OsqPa5JQ
cez02FURMxoUeplpssBKzD7ntAX8/2fotQB5bbVYNcV/Qf/dHj3y5lDDI+WtEmdOCS3aL3TCsFJ+
hduLTMqDSM1dLebQs8SyKfGDVdpkK2bERKuqBE68bP+A5tNcvTx9krC+XE/sg2dDaPUsRRDerdVc
BVSaZhjRfJ47v/6/bNATNnAr/MHOhLAgeIwewATkltPRG1P6Ryk1jJlr7+83WHl3CSbtPkMx9wWF
zYCcfPwXzw+3a3GP0EB4RkxU1A2WCf7zjopat0f4OlO7xYgilkTI93ggAt5D6lmbXobFgrGEZg8f
71AyD31woNalv/s7MnrHzc3vFvzhDKB/OAVxg/TgVhhLZdMxT7v/xKRc6yhfJro/YcnclH8/x78K
2MsWRiMEbYdru1edsFIYUEg8I68ZqZZxYfBFIhSXHBCD5wx3igewTDtUXvkKS4q7zuCMoMDD7qqS
smKtGvE6SxZtVjErFEnaQhp6hfpgdfKnLTifSUTbnfR0bp0/OForgr21AmWZZxdckB8+h3llOGrY
UnI7asOylkX3wYudIklKqks1oIqOlqerVBk2MRtBlL6sINe1RTijBQB2ab7td9tLFc+a/C/GpiR/
+LoHwXO4weXVjoOvnWXsDndwH9nD0UmhsL5uzHChhXv7ehgos7GTEdxJdzUUT1x0uexb6C/buOiP
PHYIN4Pl479RfqOZNy2+YHuMijybTA7Eca17ACWWvq6uw4pu5tBQV0UKZ0yI9w3vafTDI+Ih0WYB
j32ScwWBkLCnEg2VO+2MFlBahJ2YyJtP0VaQjyKUwD93VCeCkF1PCkp0y/lZ6EEBvTYZpLtBZ5aS
ydRKL3ke5nO7wJFNa9b3fuS7CzvASwmIpwhBPpQIS4FBamLfXYvBRIjCFHUxsOlAkJ5tqPhL2BcA
iVHy62vXcqiivczaoNFhk7G7zxzUFZScmUpLwNEsKcZOFlRbT94rFLgXiTt9imfuIydz1smTMzbL
IZ3I/JhRGSEy5buNuQ9HtPbTVm+1WlfWVfDlYEl2cpjS9k2ITbCRlft0Jjihix5RFSgiKVpgg3yY
q7biMpxFzTE0INg4v3XpNjYaTGuLnE6UinHPnt9+BQtkkKE5YaSX/j51bNGjW74+b4qC1f+kfqux
i9O5oeOXIZ3RKMVb9xRTiVYZfe0Z8/cH5slatJxfqJ9JneIO00MNvxxSDRdbxYTIWDy5ZzBFQZsU
Q/nBbzH7JI/+/Hl+gSv8HseUIBRo2ymbM3v9OSD1KFbVA8R1gzZ2ETTeRuIPvCkcEZ17UO6EkjeH
GEw5QFqre2f/8zr5UYFBLrpi2xnybSMTFoTrRuf6sn5tHq7fP9hYjUGpKnH7BllgLuNLNAkX1Ehc
c8TWEUaT0kDAUViwF99g9rn3KMJS+fP6J3qxB5voEYDyk06XGeZ5bmMu+Lo/aWGlG+DYUCimZ/Sv
opA2dk+ind/OUeqjk7yzwiIdxQY1exSTFOVKtopqM4KHPNnFAonEYrsPa8pExfEBVxdd6u/ss71L
HxDHyq5rxh2/10msTTt5XHn7Sr/3OsiLkLK0chnUSFB714QCulbsbEASTW+8+3AUe1pjazQ+p5TR
Mn0741If9YPQxCxt5Ho280z0/JuuySBdP4C6HcEoNXx/u27fmqqWJ1oHVXEvQLHnc+9bV2Ds9E+n
ME1RAIIbeUuQ7s65yPOIxES8gkWVeqd0D96kRuIC+RiUDTCWTSkiH6t36YwY0ZxkCjzGzJuKgT1K
JMvqE0Jdv57HE9mOkIaWql78AFMjIaa0qvnq8lOy52C6HLJW5RdrbcW465M5ESyEl3jI4ZRDei92
JJs5VKKmecMNaRXJGIUtqVuBpSlGhvnuX14RTw++KMbsFUTyZXTOqv2hFw4ad5UbmvHwwAF7PxNU
ahiIVQ4YvT2C5XiAh9LqQMxHPoY6voe3OAwUGwCEruYXl7Z1YfH1+bFE6IaFcqUVZeKQZUTRN471
K2uM82iVwiRZ6J8BqDVMsPJZrgAYrXyF6yO8SKyRDD+64zAReHNhC2mBWpWmnAk+uzQODBHTvteg
TAGs2DD6nXkYex5kKkfshZgD+O12X3+872wkHGMMp68+o/5DR67nEiwMA0J6fOtknSyf/5QvCGB9
O+VMPbIJnBcu6qgiETkjZVEL2WsQhHfWWUk7kyatfhRX2d8w+yBzCKiARyvkzGgKYa415aRD/Cwq
MVXO1HdBHdXK8OQmPSBqu6rQvTeJgF7BpIkGUosC8NhiR/DS7mskaJsKNIdK8fuqmuxrcQlTbXs1
wzC+1rRpDy5OHpmnNV+IhEH6Qfugn/Q7EN1HbSfDOl+s8wtjwpj8HBxAgvlYJprXqzT+D4wcpj00
r7HqC0aFPaC6SpZdQoT/QLiDrTYBfql8ekAK25+OTp0AYuXb8XLX3dN53M7FzlpK8n6luJiONZKN
JKGR6WaH/Dl0P0dSAy4bqua0fQNHWykA5H6/jK6CAb/diTV4Wp3S+2lKHHYQMlGFO3uFk6bHxTGY
sJ1tykamuGBCbrhBcxh3GRoKbmXgQ/CY4IM0Zj/a83j0WMVMimIG/4eCF8U3r8Y2gpqp+BTnRjJa
vQbYS6RO8E2vojfBF9G6te9AN1tgw2hRVCBq/C568nAKfHIrZs84RvWwQrkjUdsh/uoK9rZmjBtF
/fve4DlFjpizxNtPO1m9OlA8FQHoMuJcinB5HOuJUfrwhlOebZX4bBrI29F5iUv7yJ+tWMQopDmw
OHQQvkWDZRtS9NpYNs5F8DHefIbDY4oc2MMhCTQfX4kmim7f7jcUQkziyQdfRZfDIx55prtB0oQO
ZAeMWfesAR3U4ERCvy+yQKFsRcoiQKDNXsK0O6VjsExlqDzXw6svShC6k/+4dA82fcxTNeudx33T
ZRPTiQilDd+9l84Nym2Vo6HYcrH3fuQ5WQRTP8AKHT3sZjrhY4s9Qvcw6F3RbXj9W15laZYQLcKk
qUU9RB5QVwPC+nhaeX5FMuGA3sS52YkMxyayTHd48op8VByXw9Bk5T4zbkU/P8XkeCgXnsrYy85r
RwpWW1Kn7jNyEUJx69A5gEEBUucR2a/Wl/TiBYIZhRJvnZHODnVaFH0+fLOGvZs7Mf1Z3DgrBotU
nxDLTsSglFfLuxWizqNoBIjQ7iS3lNHkxYEilX9VOav1S2cWvxowYQaOCms9NEemo4mWooC2CVfK
gkx2dDekNc0YVdEKfUiVyk+6uJ1M+HcWeBh0GFz6UZLUjtJGU6q6VDSKGholcl2brAcUDYr+LqQX
TrAeXmxi8T4zd7eZlIlnSi4HGYnJUNRkfXknLO2Nzb5x25RG2r223tKqXJJSl2VC5FPGwNIBskXt
DBOz1IufZGtbR4Tw8T2NsB9NoE6J03DNdSeqsb+l+/VqVpZvVJWxMQJIr9eSboAGaCmFDT4wbkMx
533xgvFvOV1i1iNqloZFqbYvEclMb2qDJrmaY6GA7wGY6bXIQvolwcCqanGhDOMHOjb1MZTdxTWB
YAegMSl/+z7h2JGuv/W8Zvq+ZUBHWUqQRbndJr7/EqeIFYFFgoEqaUBAbn4Kun+yMoov9yUjlpeF
432cxHyLIZkkFKm22u4XPdOCqLre2VXI4Jnfnox9iGh3XOXifaJj1UIXm02WVy06WsNae9XlO/5l
trcy3bVJ2Eg/OuLcuXZzI5C9fK+Sf5zfrJa0yFrHrXLZ4H3fqJwFhusfTCqElWgp/lHeFgdWgu27
F25pR6EY+hMKtmeHGdihmTGP/4J1J3nF+m5NA8sKPdosAXzdERNTZKSd/iM73T2/g8u+GEXUl/am
sKYwjg56+54DZD/UGUiIjbCvyqwHv1B28X83gxX+v9ZiD2jWe+DQkKeOhsyBwm4tQ3E2zzoWkWb6
Yz6PNSQj52wsAgM5hYOB7hK9R3jg7VD88nuwKqcmLgI9OVPWuOIIif/5I80nslOq2H348n5krNYV
thEnRTBmgZcUnJ7uvR3FOKz9JZV0ctHKcG86+m56NIFuokgYO0WRmjDI6lUVMzdpKPF43K4gJJ5J
lJGsRN6+tghhThDfz5SZDEFDM30wGp9bNIQR81aPwDViTcgcjRx/NYDqCYOqboHJ7BMDQGT2oTvN
0snimk1brnRHn6idBTECORO/yeYoL9e7dP8elyMyOoa4vXqWSuPgm3N+3G0VNtS3IUwpmSnWscU7
bnB5LZTTDLgoHMtFEo8r7uTEb+je4bg6+rD4sZkSjIpTV/DnJh5E2uEAk2FM15Fp+ua+l0TcpNEg
JCtPp+pyNlnhvResj01faQACYHKSapghlbliXdFZY99I0yu4Btvcy/nDzGqSwaby7gTDY3a/UgB0
87goRL6LmWAXrUo6NpzdKT7V9JacC+ka7AisgWVwmfIyz3OpsrQFn3CsIJtba5S4gSlOEmJPOVr6
fBHcC76EFWSNML3lbGFHn/H+5EX4t0tJPPBntND1GNDNGBZPa+Xm1pBgL79iTkGZLSE4YSCGyxKX
RxF2D0JIw2ylbg+FVFYz7OPAzopRqJtjgtKbF7Ee0vQUGjBCnbmokd34ysUTLJU1a4acT+RcTwlI
SEkT/jCynqKAtUTMTpUsA4re/pxAyQ+L5xjvJS8AKXKF7kOIEbSjLEqV2Oq9J664wkoXCd4Yx8ua
A8yTUI3PomwZzGh1wZ3eHISw6PEFLf6/0BmjnWaja6gsueXoCH14XtiP5Fc5CrtaifSesDIM4quQ
aJj2OqV8hGs11fkNvqbrd/V0p78ihdj8ttRfj66eHtoHISr0AyIJREyD/qjIbBYo1ACLJi85FFem
/CuaHpGWK+W7/wCTjwz3PzmASoglkgpoZwXn8LUBLMxq3vQf0bgoKuGXlbbUW2KjqZJ6Q9iDC44x
Pm95wnVdcgcCfBUf+OdptMNDgsq5+lw8afRDzZFbA/q3crLyhUxUbcLSrOwNFVyr7Vo+BupQ8wID
cme6nq+NYDR8dskVwp//VIQ7k+u+U9nCLU9YmZSi45X4Ytwe9qvaI8FVVCtqCMHVBy/VkQaK77ZB
Fx1gyQS6ARjssIJ3T2EkKJlEGOPAdVa+jlJLO0XW2WXIXeZ4TQkVD8okSM2MlurJe5jz/AlYLBvY
9DHf/eACeiArpuxD2ESQqyydwp7aVuEcP688oBCl1qABbm9tHU7h8HJgxPRQy1EfKxVwwzyzB3tD
gvKBjE8fedR4G7vyp5TrLsr6D5H6R/LAjqmz6+wMRx9nxy9eii4+lSbiGdASxtbtAI2b70CsnTJo
I1QaCBz1jxdppol4JHBqf9GLrwFh8QsZV2JeUMTM5WjUweDrDzTTj1xBM7+raRGMrU0gGP0kaeVA
Rjf0nz5LoE0DLTMT05RcbQctgmbr7dB3vZRJLZQsAbt0+dIcRBHEtqwAUf00yiREqI6Cqwjn9Btx
zw1zBAZtTjZ81UWV0sulOuEMwWEwdomGPXujnpjevhlAQscXEECopaG1qv08ATvl9ifKsPrF9hPS
66+UWTeHo501tlO/uXgLp3KSDSAkrsEl7p0UUMTAjT8sgO1vBy2jltEIMSt0ko40nQD1wIBLhWuz
nvUtQqhvdKuVZNCqR4CF9sgrEIA4AdiRu3gJm9CNF3JGEPoVu3IpTs9eSLH+Wt/Pdz5dKp7j2qJO
dbq7JkhjLjTcjqypQoPLB0JWTwISDJoLKFTbjiXDKhXwRe9b6v0FZ+gyZ7yk9wHK2dJEyCStRxe1
aYKCI9v93gjy6KHfjz3f+iJ5LByplpiGB7XlkBKiDFC7KjIFhna3u4v+CC5VE03GGT7V04yfBw9o
PKIHWX2LDBz43uOB1oHXu1EnZM66F0GAaNmlhIwxMxc2bOVg4dFCfsr6f5di1zHIfvvLSjY8Fxhd
9AofBoMf2ig3LnkouVc03zazx0uihFZ9mFYkndeeQltc45WQS2N2RrGOPX27O2xtkGdUj5642FFm
DoKE4Mp/NL7ZSZgCEZlqp3qJafWOHZuF9WJYtlIR4PLoi0G7zSGferOFeUEV4YNnvSa+5jNzHcuD
rXud3ogordrMadNngg9D92as20/RqxEJ5pStkXUTJhZHU3GNFAxBJ+ibxDmyeMu+LaotQ0gjpE1F
2bczsANOS+HayNs+Y+VJnQfgkiFJcXels4p9vmG9vK4z7K0G6VMkYLiYjAtU0WU18SEWXmcHp+x3
hzBF9zWdxfLSZnglE0+GBY//j6mspQ2hMsUGFmmqZKYklxDbagYi9MNLAAGXDW2UapkDVhKOQbTB
MW/BYRkcTcpwyVC3lcGJz4LYtXjbNz9/mC5JaLoyPKglGM8YsqK1x9NwUPKJX3eRwSrnS+ZwvXc5
wdLFSBv0JyhSwODuY6HeuXwPG7IDDqc+69UWdTMWfd2cSpAcWV+cORflvt5YJbG+xmimT8r+XWP0
Q3rOC9G31efYYRilgRrSflS7x8oJVGOmAVYTYDxNqc4w0glN1WYOceD838AfGu2GBOc0ljYqUV60
+1Maygq3xFpdv+tOrFnSmo9AAyxWMxtrHlry52h/WyOW6O4O0j4x5AbxjbR/1JBQ4SC/C9uafGzf
Eyp7Qy0yVGRgjXbpcVnY//j1CSZZwon1n8iQIoWxQYd9b7eqJZ71XAaC3ookc9Ik52nVtreJw1qx
wTiMi228jyBhvCY3bD5o97xgM3FrTHrfnsaTW7zNx9fOGfAXwLwZEzntyaI/3e+ZFxicLs1rnDZY
z1OG86k1sZrLLo/OrcXelhgpLAAIQe1vC6uvLetQ5XId052YiNiM0X++klOjFsFwMFrm+E/8c1xY
IdnZKxdSnxnv8HyS2Pn0oww6DcBK/NFleSO9RtmEXRxpBBR6JHsnkwqbls3gLqiq/47zoU6gZGtR
nMyvuBOyLA0S1+5lC/7YijpopFnxWCEep/6VnFcRot0WYUDm++aRDYKnsQddr4UjxGocsSRep0NC
Ir/HSymnensMnIuiygQJFfgUS5wof9KmCz668VWcVrKCbPbJYBWgrHsu9Q9+Sfe0W5bkSIT7ET4V
6jJlsCEwpxrCJAr0NR21aNslwX44/ZufaH6yKtDrq6J0p15oRtRQOvakl63jvgdoTI/wh0B9aCAJ
qyPCPU0Bv3eGjTdGUagx3JbY6pSe9hYsouIcd+DbULAyej60wrsgY7ELjy0cM9V0S45SZQommM/s
Z77W/I1vhiDSI+ZQQwqIG31aDKcvHhdMMu7rnHeUOF0bwDFgUaU/Tu+3dKjgBysy/HX1qnsmdAj5
xM4eeQzXxckM1j5vHG/2q5+XiJeeqJ1bdIj8y0ttx73c0I65T5AzgL12SePr/ZOxJR9IJNIGNBy1
aO3fCuAJS23u/9bKg5YNiMAKy71JDcYcWtGmcoE+JV54rfpzP4paPAQj3nogMRoJKHiBG0+iu9G8
xBSBxDQW4K2WwnudjrwqMi26zkWid5SmkRXT/ijpneXsr+toufNV09NSAolIpFZ7lKIcCWLVSPF5
tBEVNoyHc6MF4ikeXkLy7N8diunfdL6nXyk/yD+ad9yQsvHYm97AGga9XAYob8FyKRiFfhpsJ23c
KaS02ijtW0kAPuoIoDAUhcw2Ks+NG5COQ0zUD4KRvfWtdSrZTWre48WzpvPiCfejovjYbT5c2Y1a
8yMwPwiWecEX1DLbMmbpTqGNV0xxhljLog5H7O2cyNU0wdzcJbe7Lap+V24f99wG/Xya+b+emwDB
U4d6nR4f3LQDU/71TX+fbkEFI1XbM/BSu1pbJamqSIIW+lOPuqWfKeEkv84EknG/VoZtMJhhS49H
1aTBTi9/+i7FBiSpjpHtGZvbE5uUNGyqmXKgQgct6SRHBALAdyoM5gWcWhBN6H4dZrCpxm2SUUH9
rgukY9D3sqc6sE28VD+Y/i4Nw/3d4Lu5metJ0ZqSrmYrNtZRqjfuELjxy9SRQ44qw5DfCo+rB5FZ
SWCSrmrs9VSVF+vHBtLEVev85cTmpw2ZfGGpQjpDkYLfvrH9KSlnbLTDPd3sM+hOMPMXWVWtKMBb
mtGFbKdSqUtvODikwkpF7jSY7MMpdnMp9+xvKrmRDTzBnbmjbeZSAG+ABzedfgXp71mY36/Otpoq
DJbynJism1z2XCVLOhtr8WstvGdTpRhIONp2UWBRhLh5afypcrx9M2G4z84YDNz8WgOGrLbqksW8
AVq0pqDaxfof47HF2WXeFYKAjrHqnshp5C+hYob8dSp6gFmHF0Snh+29z4w+WNRGIbUdYiVo4JQJ
cmwbRohypBAmmur7J/n3mAJUWtO9zIgs7SZys85nwoQAU9qvNzRJCWwNSgemRarRr9yhmA3Dtfvn
p/m7xRIdLdOWl9n0erGE7F7dBRXZiWqotFGsGgi7Db8rfNq7wl8nKY2XQFcNslwcCCFSskLLQZQO
+Z0sVU4YL+yHFxrmduSpsAom4AZqaVMTTpmdXM5QpuDvrwBCgfDn7Q3tOVHh0kwtrv3rbHQIuTDx
m6d9M/CjqX+/7YeyIV/VJ/Gs2Aq+Mql4JNxPSHAEN2bIl7v7kOBALw0xMn6PuzmCHlWJkv7MZABj
4OZ1rZVjpY43s+qhqMvlfLtJygzi3pCoZsOKaZRHVBOOdL6Ch2bC8CByz6wYgt3UK4cvUuMJwWce
aKjFJJUDO72GF9KZl0Smja2nJ6KZDIFRjQMhZRZPTU+hNpmzgCrcOJAAgz2/B6V75cjYh85UnKHt
Xfu3hCJabsHgur120AAQ6+F50dfWJ/Pp/AMuBKHxZsZXZaHV7IYy6bRzianyihO1NNjF0ciLYOuB
FU5Elbb8go1dPH8v3maognA+UoXc7hYArwnhcl8EqAeHRZOl2Nrt/08Hbv5d9rpI7tRBL7iuCffD
ErO9JIKGoHXkdTakRTx1xBsIyfrnpNxxGpeoBHIssWLOTfHOHvrE7NHH1QNU2SyPUxmnjsMq9U0E
9plrVG8TXFVCCf30oWXcEBBLaWIFL7taBbQuU9yRQZeuiHm5nA+VDddqhi3TxGRc1JqEeZzp8XLe
9WEO3ErLCvqCZsL9k9DuvDCwukazhK7H01GeLHQ//S3eOzqNkpcfJGua2B6EQ7Ylz1nRYM7b2vTm
hfAOLMWZMSpPhe8F7SY49AGwXaGuyclATegJxp6yCeCaM6MCqG/FeUGk+gUide0k+PdzECaNy6op
J2YeZTuBm4OTlSlH9b9bMrM5qxaSwblzQs6gGy25SIxaKwFq/OWwEK9W0BPelsmFzaoD9luXEGcG
hNB53Mnu3bf7UhLey1uFOl64JFowXfm7Rzx/gUsuV5k9Wzy4yNTX4DYwOpnAwj7fIvWLLdy7EYPL
JHpTciC4t2UhxQJEYTCgAFPE8+1fWK0I82aN1G2UQYkaABK02+dqf3C2nFGTxk2T9b1pTnHZYAFp
gKyNckP6SJxXZmBMGjY7xKV57lQk7otDvq9xS8QYGeTPHU8WP4hdsMn/JdfPqIwYv6E6EXZOc4kd
fWCelfrjZ6E1mo4a7wRJ+UedcXNs944MQzZd7AoFCz/Hch3vGDNuxZdcrw4naWHVCfcup8HQuSZ6
rKRBynvBdXUET1mKRWLwv7Tm6HjgGdNV3ourdL+/2sAVCzT80DqrinoA/SxaPZHu5I6wUhYTC5fa
Hx3Kt7R+xXyf3mxORga/pRT7Gh6bfNPeIaCTqwKc36jKkPclzJqFBeIqRXTlJUhmruwR32bBTny1
lsjGlwpLU7r1Ac0sK5SigQf2Nr/k71aygkviSFHHP1KuIpaHvkelPEIljFtvPR6GkoGeFNaYNRfu
F+DUf65vkSrMHenjgt8ntJuiHv+VFg9ob2RLX9IaRFDzQix0aBZ9+qRg05YZSIXq8CtCLEJuX11d
z0SFS6xDGP10CwiHzIz2pJ65uCikjVe74E3DnWLAnNlUPVh1x2ae3kyI2RwrtNw1mL+MxxYorL7/
JcOuGG9KXm2g870OTc9XqUyy8xkwhTq+jvGtGMGrjqD8hefVH3zK6kcZKbKUgHFldP8MRt2qYAlM
hvvYlug9JbMosJYYcd80+aK0RVWrVEGmvrqfsHKb3R3ycB2g+kIksh+WmuHOJhcSbNInTmbXE7Fg
cnQvLwFVxgdDEx0xzA7lEZG31tdRnBx9gjwnn8w0I0YOOsdg79nb1djp/bbUbH5auGhqaoJf/i0E
UnUOZ8HV4FvPElfp/l+YJiZTA1CRWe7DdoWhvLnHZqT4W9uJ6JpAic5OrEg95a8T9cyf7vaRLM4n
nQOT55ywEAzU2FQk5Eoa3PsngMAo4i4AaRBM6ebOfA051J04WpLtxI3H+exabzr77/9ZGg1uId3m
ejoKI7VlM8CXbSRn6zrL3z1Lu0w3DnC8qJqFxrVVcHzCLOMsTfiPSJ3Vpo31rklaPGgdOPcBygkC
hqhy27dycWNy5lm/HB0f9ZRoYE+k5Oy7MWVqX9q9D1yjuo8LjGj0uscpD9rIASahLbx++UTYUqzo
+rFXDjAOT7YDtIBZkKslvfLf9CcfKcyCsqX52u+rLktEcGssST5jVS5TLPKOvx8SAcyARdnarJJ1
PtaS5TY3JyAwNq/Y6gzkXT/f2VgHDcB0ml04zkocVi/CXpBnLO09zwqg/FOcCZiRwlA5WOiBFJlq
/zfZcmsxJglM2kTzI+xfwWEJrlzOdbZIBmASGAIxYYAziJpWq9EPuB3F5GjWaTdaPRiub24ldS7A
RD1HOtcLVEOYw0AcR8R5p+i6lqtnk8h29BL2PjYrOxWe2olci5AW/Ouc3nfKSWnWGP3danWVUNIJ
uAw4Snkk71E8Yjli5viq+LL0SbTrUHrFVuVa9cSXbGohpVIQraEbcewrbAbOq1oL0A+kQxkITGCx
pyiE2b1J6Cpd6szFZdTlFLwskqTd4VKgiw2SP/P34MFpFKs3rRgfixtVrEBNNWRYKZRzjTbN5tWX
yFPAruDu3yJ8CwuBO2n+ypfhppC+zXkarvqJ8RMyupVRx2oX85ZKhB9dO89ejFwiTIkcAKQgLci3
g4cyDfugcNbZ7TGOMBKa8x+SLMtC2SYF9cOlSklXFOnX++45nWmj4Jf5o2Rj/bKgjBvYUPPlwJSU
BMu0/b1VGoYYAseN92Yl0iWxygt5Yhznzt9Gc2/IgCmhSM/jGGRE51KOZMqmykgwIprQKUE38GPX
fsG86AeQG+tPv+l8qPY6NvAJaBgJRQTZkRsKW36QnYXk+/sQIpA9eBTSyaB1uMpGFttzB7zDk83q
sRJUHKdb1W71EIzlAiad7PUfzySs2zyNtR/0+DKBxIPxKPlWkTW437alynA7X+dDx/umjfRUN+av
laxOLnAuZjrWCFO3tIkiv6CKfw3utn1+m+xeYZsOE5S1gOBOHxLYTrXUwiyFk60DYF0EdsufMrgb
nW3cdJb7QfrScQicV2zQB+no4oQZsibsZekHR2Ee1m/MjkRQWNYRwAeNnt6IllVmhbIWnQsC1Zwd
lVBbisv4f5XZ6n/H4c0wGJnFQ45HX2GNUEE/UPI/SQPR7LLqvmHA/jKxyOzuDCP+SaSC5lCeZYzf
4RYpSp0diAam1CXD8x3EHzQR8RTU/pOwX1ABFdsYZiDE5EJdu+FAQec9Kg88frzsQNvdwJuEcR+/
RkYQP2rd5RGTxJ7ZfxVvkhu/oYU9w5izvdNV0xFlJxSEELW6nwC1/d8PIXnmDpyIW9ogcwKYdNc9
vWcbT2MXR1TKZEr0WvdcB8GW1bzFZAXBjpCuj6A/ea1ecwcbeyw4N6RmgFRx2u07uss+PmZ+FGOC
VgBxIC5doQt++FRPLeHyaQCsk4urffnCiDF9eBwegVqamuh2CoCSYU+pxSprVUL5n3PlX2SR20R5
+dvKyaPpET4hGL8xJY43W49pjfAAaW9SpvGM1ktN6b7MnnDuP7E0PhDWVIoLO2t5xiOvs0YYgxLr
z0MW+1yK3evwOSrLZW1OVNm9m7vRjuDDblRU2rfubmfQXGkX3SYgyHedThq6SbKd+gYQMi2j7viW
6cgD2EXyc9b+8Q/ieaRLlWNeRLRFgpFsMYhsxu448Y0dYnvUu16MG6YicR1s7eL7fKnOwLLVA/Yb
9EB4+aqi7Jc0h6aUs2LWg5lIP3kbUzEBZYnTxuVGXkHZOUYcPZ+kFP0Zx2b/12JL4lMLGK5MP6co
5JOJNMzAbOtndleD5IXak3mdi4y25lT0k8IZMnMFZsMrt3SqLUYg0MR2plrHccywS0bfW0WaaDtA
GzcuO2+ASd+lQmy4Ldktod1VPrRDsGr1u+jPBoa3t3CQ6TKAot9v15Cq7DAAAYgOaBRD9R55kb1R
BtpyC0RjO8R3CyGnzzuvC948dkDWt/bG5Ode53KL0TJPLzhf4WOROEmgxmxup+JL7mgZma8MEkQy
v1E82DNcYd4h9XQVTbzVffnNXIMbEr8uy33GhQ9KefP1Qner2yURWSRN7tBzH1d1b5CepTGL92+7
F98+fjRbscOm7Hp3/Pxfk1pF1w2KXUSQAu2uod7Lm8iOWIf6jE1QrtpHx45rkvvBkPgCNYwS3NdC
ZUkS5HYaaI2B6rq3YWZM/P+sD6a2UUCzDIu8uRf25ObrkbTb0jDqVQjJBD2vDVsxGn4W6xYWhkRq
98Cz/kKjOlIQCE04cMhcGyN8o4C+xcJHQrKbT89BgbIw1AZnrb8dE5Ix/qLaCcwE3wq1veyf5m1K
1LIbzTLKygIkpFZKIW94Z80VkFPM2HEDqd4E8qa7dgNUaxX+Dajo0XuK+ipum03PHySZQqgLrZb9
wVQuncWFud3DGG75D5PgPHURV3SFVs9kfj4AFZfTP6msPGiizkOR9dsKzQnHCo+OrtUYk1+fju+C
pcNjcjW1oEkiaCfsKh9kt/vNRkEELpW+wNRS4Fzsm5jkQmrTYtvD2O+JFAiwnH5zOb+bUnDGBqF6
Sv/O0LJmqMZ/Fxy5wt/byGU349xtbFKRWQeFq/spPY9yurf00RCcZyPNzA4nTeTGKjj1ITuOgBAu
1I9bQHEYbxrdn1ke2OA02rCr8CQkhtGmvfwtzGhkuDZEI/tL3Zm3g2K2IOuJuEnHn1ZsnXkjWyol
6s2Mf9lRicyI3n9b2n0lcBbgY/mAXzNrhwNaDJS6nn0eRF8vf7q9vry+jWTWnVIT8DVglycguz8o
QcrqOT+ONZWY1l0WHGnNdXPQHo/vaGT2rhMDtnySXLgCEvh0GTJIAGxUgDgBh1qRiRZrtVStIlaa
sIyhpm24D5Fvt9MXnpL/P/ePw8R5gYJj3NwFZiS/lkCzQKvJlmkkYd8W3UOncyW8M+2TisxxFBB6
ekmCaknmd0rsO3mG5VsY+m3CrLWt1Yey53RjPeGsk+k9+Te+QvjnoH0avqzVwseUR3C4UwQx7Td7
37gJg6W9F/U5krLHhbDTcIj+wjrD36YLfPfWvBGSdgED5D4xSsUbhupV4/8QJ7ymRuVJjd3TUDHs
gi1zRweHv82LW0bNcgGXYGhNNF0ScvUkscNziPXNYX+oZPhd0UOjnnKRT88+t7hyZmOyzlh1Mo9I
i5Hua35rkfUZePT5UjbqUB0wbh2N65o2GZ2PDuhvUBl9JgczddjOEDeLJHu6tZX1WqcQnKkAntgj
Wt/4IsO6wOQU86OlwIF3Wssv8n8FLVv9kfHJfyMhYh6c3wQbft2sH2YjbUtu+j/SqYchTYB4qQ8X
nP8KmJV+f5nSpYlfWJw7zTLxOIbD4ANKhDmTFgvRyFKtHkUhVKSiAV/U3Tqo2Y3jntYbmfPBiUpy
qy6/psATWdDee70D+yKPDpOMMH6CdTuTcbWS7sISL4ExnpnWfzBvXYChqTkRV/BKTr1SqnQ5sDU4
OGLFleoYYIcK0mUiEpC/0Ns8eLjp8U6jQWtEnOFEQZ+vtEuCqbZ/Lt4cZ0KVKRlnCu21a/55SPOk
1KWRfl90tR0FEnpwzQx0ixVUhtz2KE1vFUzuoUtd6+rEHaKmNf+4JAkIXN95GYrzn//xwyBrGryc
DczwKHOjUDhnYsDEr/ymJ+IcZ9crUNXegG+HATzTeu59Zka2WRIHy7jTqD52B09/Ys3mCx/7mRze
bAh1E2SkkCrymiMdS2B7OfUhdNejnY0W0Ic7bAbLFsOJldWvVC6LDrXfEZ95qvVB4TAOaNyYpCrb
yCP7nwSOKTo1Iu32N15VDxQtcme1/F469cQ5it4rpKtqm8GVthco7Si+9Mew+yzJrV7qoHuP5eVK
QQPxbYZ3flfl7qNetiaetH4Qld+irGPKKWNkEdXpfYFaiAjNmInbn3RDXGSI2iT0OkN6s1meuP05
McV2uwzQE2MaZ5wWM4AzZl27Z9NxOOyq8BuUxTxOcORuuEOnVIEY8CsDM4+zL1iaDNfIUON4QOaQ
CSnQrpL5oJvoQqrbqD0OB+n/sKdMlsPaqSPIFO94vstCqwkSLSHsNDr/Cp72ExTYQzunmdwl20Mb
tZVuTppw+6QIsRkO3Uabo1PtdcPisOeutFxMK8SrbAXT47tUgCghTNTodo/ccaVHFnYuWPh1tlKD
sc5esTkBv22Z6nHk3lB2t23FG1eqzzGjyzyFTG+EpmKAyjjxRhnhkLgZ3IE+kuxOjW96vqaVg4Xs
8pUExq/5MgQg647Hynyv9dwirQ2rdFT6emCvb2M2MK1hd9kR3J5YPeP2Z0KBbYazX5etGDWgqFky
MOXACLAypyeenrbAsNIWuq+y4IHlBVNHecn2aZXZWdqsCyNneXp0ZSWal310UdD8J1ktX2Z7/xa4
YfJJPFYj8BG75dF51hwh+Esv7vg3Cv+QUiuBlDzXTkB39E1bpbapMgrIEfHNUUe3cbKY22O3faj8
fYtsXzwzMR7ln+jXWDtuxEPwaj785hcMh2FmvX1L1egd0ua98C6nqyKo4jlvQzR8AHc/FJnVesdF
BMmbNv42g+6IQ2igm2+erU84ODTSOi5bdVJBlpsQBsN/2sau+bSRhgTo5HJ906RFocKxOc1SN31R
QXIk6JgHE0YvrOV9opALQncDml4nKjSXszXhu6Q9tOigTSO7PI4rC9iVKBWfgnGXSlVq4pEPIG/M
cvUeW+MW1lIF2R5A6ZoCukh9S5nW3cNqDXE1H2YU43KhBUXRTjn5TTntJCkBG3vqiVlwmPU0sTbR
lW5Lm2CYTpuUNv3sCeq26YuLYLaNtePMEUwww3187JyZiCHCb8VGmso7acEoJka98+9msgaI5RMb
ecwuaiDCd0/lQ/4AgiCrhvhxmg/lfNDsPw3YaTYsHDDko1ZCTx8BCgLwkdjWsyJjUMcTOv60iTN+
6pa0nARQKGAqVx624ZyLmDBv9/orT+C/I7PGaP8JWIUnIlSXbwsqAmJnXvabP/rEx/XJO9VILNVx
Ue2qu7gQHGteZZzQCUVcJxpnGMlxy2WnlJSpmLsbfMbwqK+jjYBfc2SfHhNF4XefcKP+tK4zGxk3
OxiVuS7XAVOoz/LmC3pBCeT1aFbM3/nsl2F4NnhNpUXj2dVU7VuV97UQu8zFKPRrGDyPSDMlTqw1
cO20UITvlgyltVuHUda7KylgQrB1KQIDUagnnled80etLgGz4442Ty9DIS6tj9O+mkMakMCxWvhq
fZDlzPQRHPLVS3JRs3yKJTMa0fQt5hchBIQhReWY+ugt2bdhd9fC8YotMLpsja50aGm2khzjJCE/
CmQTlfGccP2DNJJTe/m6uxjR+VKGGSoJt67EqWBf5OqDwiI87pjCeP9Gdjzo5ZATsa9S05MFAH5K
wxH1DZy89fNzb+kdb52QQv7Dhw9Vz2Zv/LSReDlHmwG7fHQfXEsF/2RCTZslMSB03UKvHMwuBKwp
Ri6qEpF9E8MQsvnTA6L6we2o8txDnoORqsIKNPcUOVTQu5KWNa2GnteE/13gltQu1fLP3OJeEgwM
bYwynWZk2F/FK+wo6ZgIDfktAabNWtMXcXNyIgN+NKq+nZndRWkSTPceF7XSuu/qZoOU84RO597n
d3YAF7X35FdLAAfGDGG34XeD8HQhxq60kEWLytLIwdbRwWRjmTGWSlYFOJyG3Om1Z69YYfvjUUGv
mvnm5WyFxtuZGhpQcJy/569l9nXKTk7ZwNZhjPYObspCsKT/j1HpaYmSwUlX8dcx2KPoqjnz4FTV
fr2c+SJfDIx+OzhjyNztQHbNIh1oVyADBoyKyl2hyVUqRI0ugJE/kxwwypAykRFirythsH3ovfRf
J0AhlNa47Llk3QNzQ+A8a4agnso1wt1DaPOO+hvVo+uzV+CtQ+B9dYRnXeJDzuTdjblfMxhtvFhH
iL9R4P64YCze0Qxda7R9CoIKovaKXrw4nlA21JR+Jkjp9eVRDDxM4uWjDYvWpN/YZSZQZ7NdLdMl
DbOF90xPbaCYuyQjwF8ILssTqcuOQdvROc1moSyNosPEFd54e8qwWyakgMDaLuCVvn9mygkVOE1J
P9ZsyNaUlI0BWp3fGQtVkZCx2OCOa/SDeGJdQHztnuf5xCZsl0QbLjb6geQFIgPy/H4dje43Bjci
vftSN89aL1+c7Pd8yYhnLrK7comhLBlYF9Ae+gx0+NU+sAW0L1nLy3NcT+rGJu9HQ2svYjF1eohN
JAdnTzyb/+MGkNllBLXPPKvUfnDjlGN6JzrrKJpJjUjw512SQZiBAetZDtRXY2mITepPdtH34QMb
yZVtZymGkh2CqqvXSPFssHMIGPkglpkWRcf9/eEilju8gQy1z7rmRwg2/FSqGObrJyEzshnJ1rxT
+81bIdPiAxt2hqmReeCuFzQbfT89iZkMFfGNQKuYpm3wKNGPIqn5k7k0ro6TsJFsuuoa2gjKvdBT
mxT3rNO5LXJmLmE+kOR8dBN7Duo22ts/3lWvpugnyl1M/TGNXz02wmzj9emhb8xMJalhNLxPH+LR
+q4+KpifERVVR2JKSNpMYD/trS70aAxR8oxw/d0/2o4y192QRBhrCAxIDvz/aWWQcbrBhkDoyRUZ
0XFMstfbdpgDfh2jnPHfZajOGsjL3YZeb+b+4Rp9BSm5+eH7H2yl94gtR4/POleIf2owGDPZFFo6
4glsBxLpqkkm2tlcwwQMxnO1C22pWyFYYixAO1rEqsb8bNw/xOmVRwZ2KSq94KM5rQE9W3Vz0JZh
F9SHEfOgUnTbZUflEccy1wRkLtBu1ijGaRfUZmjXrEtp4GEIA15cwOurojeaz8cloeD7qfAUo7Jy
ZzqvJM5pQwhBuehol8ni/ZFvvblWFEWXW1qZz3kcrfWaTBKarvSOeCOwOEHB5O/ZYDFEbebAYAQu
jN6ym4hi8rJl/04C75jE71WmdErt4JESRfXMKxh16W03e/ppxY1xF50AWbbhnXHaq08cwT9b/iTE
UosItUBCOw4sH+MTbIrlU1ZBArGS2xxIoshbjh2nPRHTGbzDRfrB+ouiKmMhfZYbg3rHNmQdLWGA
FhCCF8drM0AEwrA5Z44VcFjky6KTjEnwQrc7+KgTp23zzcetv2lgDihq6HhmXMp/D4klGZkqeT8W
larM/HTrTKPj0swrsf01MuZihj93AhFtE1lsgHMXOMKd83SRhHH8pPlrKmJfNkrKGakVHg/Vzz+2
ansEv8uRCfyol35rAv7qRnBBSfzu3pidr0BALHDBo93O9JePJ4zID500gpcuPVmCzP4pM9KXMTdS
eYGYcF3CZRvaDa4mcoAeLyd4QqcwjwsH7YLtI+2pF1kYY5c6vRDfxL+hb+a8wT0a3K9L75FdXmQf
0evSQhwpT2b7ZSbKxzOY3HrbHMUvbpYnkdFwjcMYo72Ju4bypTjUZxbzDW8J5huggHFIfMEi+8WD
uI7hQcr/+/R3m01V67sj7zJi5/ira5GpJEXPcA7o9+xL4c/pQEQKQ+HEpuGoD36Izly/ezIR19EG
sU8JnWbeY2LWR+268z0dLyqexgh9Op9FUoaf7UXRs428xnPY67C1fjaBuNqSQY8gmM0VFJxiBTX2
7ueJX4wRGzBvSYRYTMLSAc0qJKK9an2+fPw5dIYgqlndE5uTVMKZPs3Ybx+CAeb8KuQOYgvE+UcG
Jl4GwrFTVUNDY2/0rtbCKagmtT7vkSuZ/RNo1xoVATpdweXlZgmuCnMMi6fYIol8VTsZMcepUF2V
bUvvIl/p2TPVzR7fXGKDXrQmqvGhLDT6JLW8XOXvCMbwfCfR1rD8AIBPNplH/5wxURryYLfrn30N
LsJpnWDou7fhKbG8z8YDNR4VDSFpac54V9Wde29YyfP3/9qK/IbFDZuYp7DJt46iqzCkodFOgsQM
FvGk5ardHEg1X+X+JW6z0uhvv4Y4IDgQdFPXDyS3ADI8tcBEUgmvEE4OitjhH3NnUL7K3wbMXAjM
fo/0MKqtpDLEN9cFATp+kA0nHo0t7ls/MWjFKbCxKwncfO3bg5EFMft6iOW3HnIHehApbXBGllcx
FfYYTufvG+QONI2vkmG6JaP86DXUtFxnhTDKUqAA6XuTAFvcHEvAHNct8vVwYy37RyGN309HcPcS
I98aOttILXG3/eLp2izpC9R7gzWi/23Nssgug680A0pliKy1zo9eRIJoKqzqRsQ76esd2jwavtny
T8tDBlIPkoDHI5JnVueVQpN6r2oXt20t+PmUf8CiOva7cPru+/MkEA5gKaInB8qVkVceAJQXNEik
fh3nURVpfLdNEIEkV6s0hHJm/FXhEJJTGp1Ybl+ADkkecUQJyZ+SV8/xaFmg3ysXlop1Pht7GL3r
V3syG+MVY5lh0/KAuQJhHY38xW0lV05oRk6UfmqK4h8AdUH2F1423xnhWiGTUntTBKOaGtb86bUR
ODi+kVBTdBH3lpaEk6PxmILrCZezZyXt1f/tX2GTjJ4TeUOnM8aNKBNHGDioczgjvXyz7QriLYO8
asDW4sLXPQ019CrI7ky+OKihwIMruowUA7FFXuL5A9EBsplPHq+UPmJ7hOW0gm6XlmiFXDCK2w3A
1CVgsRbI+mRaXKVfIqZJABEXMXGXTnH3OD+9JFTN6NgplytsdVRdx2Z6qT/jeB1CKa+6Th0fYCNz
uKYZgR1Ugwl+Zo0TirrgUgzzv4RLONLpg7Nb8iXQuMOMccs4ExaFZDhs/lGZIu9nDJl7Des3QYPg
b8DIXK7txW2pzOoxuc5iPcPcz1TYEk4I1/3uq+DztwNacevmmuwVFksqPiwxjxXVfUWhYekjNb84
RtLflNu/mDbONBbOeIEP1ElYaVORW9Zndde76hIevp5o/OaBrPWcuESTz/r+4XVFZj68RJ6NsAoz
/8cRcnTrlkOjHtJ5DHEhfV8kAya+DlQqhqYWrJ/WdOUVzRNUK2U2G/VGtcZCc0AWMKZqCBL1tWl/
ccctwXn+nSbEXEmTbx8rJdnOpLiU7Z8jnA1dKfMSpx7sGbr+6KZfGW4mQU+cT7B75xty9oXVZiZB
wgB//9vCGyI+Kqnk2mS6gqWyoIC4fHAhU10A1jJbhBAtTH/22i2HAR/gu6Smig7xS32IPFhkJoUx
X/QMp310k3HUlVqcd7gTrifiMDEsdhSnx2i3pBykjxY/ZYesFqPZsueEqosHGlWOLoF3Mx/PPApE
c/syX6TnLmK3bvltD4Z+1y5tzwlFC/bYYYNmQ0e9b2SUqO4iJh6SOZXo82Qx0XJ/jf9mIiXdxvna
N3Dm/+X/EiNOP5/rjZnZwUgTrj1MRmquaJw0sI/zAIZVJ3QLg0HpllG2OOmGSEbH7ylJ6d9wQi+J
IL2txwxFjMsoOCtwxzZInBefTzbLVd2RhWDN80R/Zy8Wrb8vG7Y7oeeCA2DO03SqMlfXn6nFlQxt
rIUtgZG/Q9/fBnkEwgUQXvDVwcaGi48MOuaJElUwz5ym+e7ho73ABQ49GxTy7ezsdtuBZhjzdyXs
6GYa+ibGacE0Ziq9xlg3bUXbLSXqWthnPos/k5MQOC9Yv7htRLm2MSxbEHNZ+CNorCz1zmh+O+2O
Kb0Y4uzsS8hIIj7x6AXZg3sCROqr0EyTy/Dn1OXG27Ad7rs3WjAce1J1SI9S/gqNveyCepyhFcli
xLWazErgbBK4WMinrugI52Q/rVCkmqg9N3WwY7FOO/8YUhQF65hpQ4neq99QnyM1bxXPS2+kf22G
xSGmrSCDlFfO8mCxb8UmNBEdGCw2nicXY2IH2cuj+0AD/WD2xf9lQ1+EGx7x25xTdLyVrc1xpy3B
k6II3ODZu/QneDBHsY951cUiGRL024/Qn1VWgsG89dsf/hud69kJPPPx1gRyPjjetr1EQILqK3Ob
6d7rPYQK4uqV6gU0z4H0TUIlayBmes+UpQ4QjgTohMVC0CyrWms30yhNbrgg8cOfhqrlHihkd/L6
eZgiaI07ZcZlgsMN77EVdbzk1DjTZYBph7/aTpfTci9wobcGx4d7iXwVqtSOmoSKC0tekD8aVGjP
Q0Lue/53T/meszBLoMXzQD8O+52fvWgQ4OdwCONtpT6FkGrnNwtWxvZs1h9RYdSYvilWt/Msa0FU
GdZkpYD7gjyOGivex004/sS+tFP0VSbr6tHYX6QiwxmQDurbMFN7Om8D0kJmMpFCe06gRD0FzBU+
E3kEdDGgYF21folnKzoZFK30NNFOt7d3t8f46uKuVtKRjsVuBA7VH7V8Qdh2RjYJ3VasCZPTcjUf
2noJ8CerZu1zKjxEKiT7m2oGYu7CW7FQW+jVrlS0nSeRmiVCV445coyB3mA/a3eyB3tqUtQFM9Cj
tp25iArwlSCiea+Q6dL9tXzR7iMwBPl8jhAicAiXeO5/QnZu9MbTAR15Kc/RffXwbohgY9OuVDAw
FwkNEzNy0Ar6eULmKMQ6+wrEqN7D3WbEf88lqvTrvH3dlVqmz++Z5LeMG+mInnxWs0bABAf5/WOg
RX78TagxPzDItVF9rJoKEFG6auINmtrR3fr23xmiTZ0n4NY0nLau6EWQY4etXxhqjtPvafSDJ+V2
ydiMb3Ngf9PWmOLW8Iz4WLYHEg/IhQ2XavUxyDjx5VxqeolB8u1PMZdYepDd3K4O94EEtEGUGIrI
9RxMWXl6OWIn9jOUi7StgNxAbFH1BFnEP5a3hUi4vkgnY9PQ0k9iJ4PqLwbj8lOPS4K2E27Yq5Qc
jsrDI6MGHLd6ym7xQ1AXgPd4iWIY02NGSACjt6bDriNeg+VySLOphTHKm7KwliQKUdnZKw4hj5TD
HOOSkS3YYgyBl7me7+8r2kTDbxE1bbORV/O1FdvuVr6WzfxLh9sp8HhCWqkxp2LTXry//qJfisNc
VNM9frpZNoUIASmkTBHDzO4JC6DxUbnEk+qsuFOj27IJMv8wx6CXj4PwLeoh2RKtNjrFnRPMgb8T
KMcw4WG3O4h8Qi3JPiBOwup1TQefT231IwBSUaA3FfTP6xguWWKfJ6W8S3Wfp+NwCL2QHJDMTjbw
vqls0ryBDA7S6sSIKddAWz0/bPrsZijXDna4hGywd/i0RKjA7i5eH8cd41c0sXxA2eQ/d+4ZqMbj
TeA1l18R/V71GK+dUMoRw2jP3Gzts0YqqIkBpTQAP0bCPPLmpRhzhsAjg/ImA4Rvov1tivHYbj0T
JjnJXag8u+yC5mnyXDoXvlkgNMQkmPeQZBW+W6NrDPvu/eiutZUTnn4K7csxYMdumpUWNPRuYQ+R
JTZgAIa2rhFOtoKMqB6n3ap7c1H3aeTcb3RxldUPceZUqYC95x7vdZNy+4UkIHqvCazyQUqhZbfd
SNKuANUqJtcLziLk4B+M4Wz4IabXLARTOLWfzAERHpmRUq1MZ6iSZ8nvcV7WfhwesgbTreis56+u
uVXDXu7NVwJpeo43GSmAIGIh+Sp+GRaH403aCHZGU9z1qt9YN9Qtjev3JOfqRmMW5sJD8zQKImib
E1HsCWkZqwo0hyKhiuqGLg5yDjkPlMVabdAh4sIZPOhWpkmI7wZHIji3qmGqE9SeUebIG6f4xw7m
5pH3TeGM3FtJMD/X2a8RWA60U86kNZc3EvBIxfnptlIthEKB/NgoiX4pCcZCa2Tj0aDeJUjN0b2h
oP0ExWygZmoY1oIib8foYNzmBFlx4FBcbGfBkt7XNBrGMP6L0UOP4Owl0qfYOE16SUC2W25Sbw3t
I/1tEsFjzDQOK8EaGWWEBhsjEu/lZAR0EKPnqrhv457tgL3siA+vYu66hIe0saYhY7EvLXN1UoSg
4L6sb83e+RQ37egMEbXFUmASIrvSElA1O5J0fYsgW24GDvcq5GVIa+PyXjfgQWOeEnYPuP3Wm8Yb
MQcfe2JVPuTCxh9h3moZCC5zvCN97D/eabgjZTE4vLLEMFDpcTRBE1wa/K1alh7GMe55KDdQT5kv
wRJE0FgcJGf3+rsy1/THUXaOlJBN1fKko/J86RuRo6VU/dbswkWK31UrVgjE9hiavUsFqqphRUlD
LclPpZoWXXrSE4AH7qWVXn/hPu0+PHr5NfAaOMLtNX5Gg+u01HCNNlO9KTIM75q/HFJJ09p4iy3W
fjYQPVDKkbVPgrajCJcJpgBbbK5jTWX+TUnyBFXMtO2wBoNKWX7STW0BAGt4sw69LWlaNQ2ao+QM
frwXlP38kJYUzyrTeoAFMgdwjtd40GkqYtuWh2FWsKZbHKveKGWEh+uSFInh+oqH3hzx3qGV9Zs9
ScCOaZwZR4OXwkGzl0FDpXrx4n/oY9tiNybYBK0m9EPOM0JFXt8Ggyb5uYYniGGyM/wpiDAZIx7K
Lr4hXA7uQckhOocW9n2PxuKZOTbv2UENX1ehxhrKWSTcOSVEmC0cGatlHbx9kRGJJtCwsreObM/D
qYPEo8EZ/6vww6fRoCITM4B+hGwOqLNoWUKbYwuQzWFYso08UkW2dZH7grfh08p3S9dmDA9PhjeV
mk9TUm+WkcaX2bTwFRn8Y2/aQFqIO/4ZnKWX6Rw2L97Wzhr0tBbDBNmvCQFlSuMfiTOjTcweFkfj
Hltg75HdrDn0OSXh3RgfluEhDO71cEOLxVb4LBWEo1v8yrOz6P96oAZID5ob7pHCrd+YwT4j9/3E
HOX727KaKv5DnKqx0HOOvdAoJFeVXapu11iqr332VX9LORnXRZVyjXNePyytz7/7oNpJ9V7HhtY5
ASaWEcxVHMriwSCz6OkONWpUuRSUss+cnDyUQR5V9/kPU0gNEdc5OruVpioO1GMOfheX4eh6L2uG
n/Bw2g1PLloUt9LxthaD702vsg5hsmqWZWnrz/5OSCt3MrbZExT9FEpdS7R/sPIhmX2fbrRhX8JI
sDNzyvFvxLEhneuYerJZ3CVu46JRdEiDqGajNZvh5GkLeYkjPtKNgXdCjbUrJiXTFzApwTYFyFTF
qfuF/IELrGJGkcQ5zA4U0XrSeLep5jqxtSEgSFiSYDOzA1EB4J2akxBruRTUdJM9EhomhocdTPhy
pGSb8lnncE5NAfEsMOtzuQTqclQK8kat0jdrRfaZ0Dc0jgaEJjgXXupOPk8pte1kPq2OcjVdPk6I
WIxigAGCEOkyHQ2v4TdmWZclJewhvfOShAPsAzmIwaV+vl70+wxdEwjKSkBXhp62IwJjMxlwq/g2
BWmcfEQ9YpDiaU2sRwtOPDklN6PnXZUdeHJ6rTRpNU+qrDFFkHV4ESDUYtGfK9/Aa9a/7yKaCzZD
5UYOGw4p9wnqiE+MgSA4EFbY36R9a1i7GXlIbNR1UoAX8MniCWuMgXtkDjJTVeNoT2oQitZbcNk/
NZ7rhH5Vm3r3d3m/OWvbXz25lVbfc+BFtCHXi5M11+4lasCJXLeXOUHSodHOX2huey+4JZVlp5af
Tt+6R6UBFInpiOp8Ht3+mPBvWhkCneAIqhAFSWRzvU2NPTFDH9iZyHTS6ifDffAlFvQrwodOrn8r
o2fa3oZvE/XLJhotwI4bbg+VlpF9dfKXf5SO/fp3hFf7N8Euw516Bam+EAohXKCDhEb1s6qPlrrP
liCwQSHsVAzvqqUeux0Y1LNhrtGmRSQs9x+ZMrlPd9C7nhZjgfir0XX8AwZxntqpjeEF/lG9C3kX
hpBhJMOmwZNyERfNxKi+HfghXDnWIttCw5eGNmV3sWpqHSvbjOrl5+FoikXprfNHRUoH1AJqDurI
05WIUlWbQ9e2mISugG8nBWHV4jm+9dIrcJztykRQBtXPSME56YZ6T43T5B9seuI4NyM2IINCD62p
o8oKQQmyeHvjR8KFtcjgTmwncmAqn3zhtLSIdB3tu18ysE5Fct/5KOmttALCl5aEh53+SN+Kckn+
Z41fTLQrAc1Ga324xSGmnP04wFqCna4BLXAiPqs6OU93RnI/DCjr6HKEtiZDAYPcNSJa94M+X4aP
zkFZTpjkVNwBJrGOaHi0u1xHt0Yv9sAIAJhZ6wnwmBcuePeyC3NZF47Rypv0U7n2AGDX+JZoj/iN
4IyVUT8dotc879d+cQhMlh74j751xFO3fj9scqDiNMLr/jl3SJUFtnZxchovUfVJKBbFTuHHOM9M
10qgX4qYhOjwJW6l7vlJhWKEZOqookrdLItBsXfI4NhqzV5MZ0MSQlUtTMSjAMQCnKpdZPH9TRtd
Hd6mcPMLAN5QWCV/8DYpyfvkS7sicinlThJrrXNU2ficLgRqUHzAPYFnpN5maT+7kVFdNXLBXpkn
O15v70KKWH8/D9nvWjvxKaUXmgb3TkZfBTseAzn265TISa0VrJQXwgRLzXgmUYavwe4RWd1FSzgj
RMIX6OTvDyGArZQyVkuljntdTSrkcaQpF1EDX9jVrpOtcxVo1mhIq2a87Wku2Gth4W0EgoSVjEw8
JTH7tICNFdED3qSaurb+geApyQaX/SGmrdPyCYpkf1cQd44Eh2oIQTL+zJ0wO8jdZs10gVBBI/F9
FtUpzhYlitpYoHw1+d4OGpfTaVfMNfWisr2rcWOdjfNhFo+56f4RzzDk2Q+xg+ChlDfzpKOuvsH8
OGLVatbMCAwlWRrDsK3fWP0igqRmZ2usb0WdOnR8Nza5s6AScMOVkdYmQcAWGcRA2yTs9iRbN+9l
/ZD9QFtx6olJpLRwWI33Gk22Mk2XlLlt+iq51KoMb+IdbD3kuCXuCDntA3YeNf4nICM3op5eUiWG
Rg7bnMt3N9/WpUsofV8esV+STop0ilECmC6nt9VjYDFm6PQJd6JIS0LRK4vx6YKEB30BCyVSOjbI
niiN5FbDuNwDcxdKt93qtzEYyIMO4ygHmyeTGwWCaROFNpAmThjAKGDVrr2alEsT3vrg/k+bfMzY
eVT4SI5KG9jWLxEzydit6/6uIFLp8NB9LidtMRkEfnPmMuKZHjmvTUKtoghwq6VwX7LV/a+E0rqr
ULoV3NdVdNaKcXcqDlMgJ7aUFzK21nRk1hfVekiDz6ln4kH1CqwClMzg1SRtmXyf08ROg/B2d04J
ecNgLzFu1ygUfmgwy1jRpu+g3UJn4fBnoU+T5jOc2Uvk6Pusey97q7HIXSDm75s+72lzdhenkZq9
AQHMzWE8a6NmKGQmX0R2khKa1AMLVcv13z/O2aHGF4wBpwrpFYKlTT4oTz1yggwy/loajrZVWbox
5qWikzRuc+awYk2eCZnwnvS/nzQxZzYXqFHwi2ZoOaKoSLxMwr68d88hK4P6fhPIz0Cd4Sua5N0s
k8FpzxqPBkb1K89c09wsFLBVsKkghVBIeS66lJUT0RhcTkC2B/5Ou8QKAeYG7JwhVG9lmA4fLnpQ
JqByOJf3Y2pk46s4l1U58uYLwDrR5kSwwz/1O/zdizpoBCCjfPv/eXe0XOzl81sO07/rX1rDTNSG
JxDm/9zWKReEy1N9gsAGyOz+L8W5N7HLqTNeeiqYEqGg71NcU5MIwiN416cI6oAjcDoN+M8oerzr
7Q3n28Dhj7VDKfLGAX5AfIAHaJZHaNHRdQ8eFtupi0u4O/VlvKUMjKKr5oo+pgcyNCHbZrz643N9
t4hURcq55q6cW1HFRBoCJwvLDDHOiFY/2NqRI4uTqEQ8V4qF+nQ5C8bsskVHvmk/5G1cbS078ttZ
jFBCYgKGsgqDYW4EWpqe9UOTmRKk9fhvW9s9gHFGxFSRflPytEZT7nm2f+ANBK+YEuD5s4M4NGlc
86eXPkiAM+5d4IN52VXVl4EprpHgrcI9WN/yrIbdo/+mPpI45z8P8CTjfcUAFfxPTiaFqEtslkBD
4e7dgB++H+OhTzEzHNM5YrzOSinMcCOG2thzNycwP62QbyuMqmD11Z7NYsaA5ixnic6KDp/z7P83
4f6Eb/KTxtcWrGYxgu7+1X7hg8mUNkPIyaZPCioVOO/4lP93x84MIPlnOI4+PC2XnGMvtL+8sWF3
SqH0TTVu9s813/khq7YSMLuC+SfB509cmJw5GpnAJMetqPbcIHq3qFRAY83Y1FtE/Rhn7aLPzpQL
Vibs0vdPFhc+We2sUpPlge0BmZrS5bPWu0iz8Nzxhz8ftlTMfWQ+bY5+1S7ZWA6fS1hRE7GTMC4s
fHDmaKQZcCKi1FaN6/1OcfMETBf7m+ZAbCP+MW8wZfRK6Wr5ETDbyEdutt5GpiKOXyXiTg6gOAwI
LZ539bWFQZMPAogPDrXaHMWMWCs5ZukZ4hfb57MVpIEF7+ihoKkfMIyeYCdqSEkC4ww5+e5PYRag
J08+BKU2ns1rinfztvjBg+Paa5sy5ZB1xNgToKc6yKV7Pbv759nQ/h/z6AG36Wlg5EqJEz+z8cRK
XLMPc6cHaIyBfUSMgs4VvL1RuIJFNHqiL7xGK/TRbH82Oj1ZpmM2d8TPZaOJnqyUKThFATfxR1Bi
mVWixaDZKlIx56yZwzSn9dG+TXOWRkQ8d7mcU5d+R7zZB3EJLYvrCnmSaFWlfXHg20MQPJfd2c+S
oNNF71hm+6UL+W+G0TfF7ngmuh/TrS26jZ4NwwawWjZsh2zEXDR/HB4s9QJF0VZWxv54UNNIbMfR
I96AC/cYLITDFjrcVQoXRDe22HqVu8Z2Ihg2e7KQhni7i6PL1zddieFJaV1adHoX699wg/9B2gIZ
uMBZIm5HxfXsYUhDN4FyhTjOOJ4FOAhFBJOd7jybNjVt3mmV7/r0BC5wWnz5jbgCt8Jj4A4h/20z
gOcwZnfYENVjwUgZEFDDoYc29lUNNwFRYGvH2IWldXEW3dJ8UpRUWcJsMYFY/4QkM6E6O9It0NsS
FpGlPTMlSIb5m59d8aLePftdQqCXjcGGnQWGX/vWC/9OZDVbVudcPOEJNNF9sTe45M8oNCIYHHLD
jNemoiN0+0054isZPTL5R9VtsBBVZ88C38WmW/mkAhjL+ZOA2ovb/qf/IBvYXmzjRj/c5VTh5CKL
JsrU4QpbaOOuxT7z8LRlmh4np11ZZkd8YvfOADI1Gqr5q5qROcb4INtnHouV2+zHyqPi/GG2Vvud
CefeVLE5DvDuFNNSNA68WYPHLkrXEzpUfv/RUcnQt4bO5HgpuZe/5c9BnFEE/mCDWGmYCISQSamp
0o74h0kbBtkBzxfEC3ulmE2y7gilp+AI6D/kmigcSwwz9/WD5D//Iiszzp0BaUA/O8aww4zKAGic
PI76Bvyi00bU0xHQ7MmMr98ZmLeiuZ3F8qTyTaZ/s0r5WI1ofa4AUkNdPuDCTB4ATEqDv6WQZN0d
zeLmmsyp5clFT8tqbF5pQGfgiR+8Lmh1/kFdzZWSNj1/3xMDPUJ1foL7aF+Rf1qvqTU2ENGdMdwV
Xc6dQ93Kjoj+K2dkkEmwrocNkfIXVbEHB7V6VRIHkWb+FIUo2UGqZvUEAaza5RHyI44j9+NR82Fb
Lq3tsadq6farfiHVUa0qm+vg7Py3CLYrtjua6xozByhPzfpNWhj1avbV8VuEhIKk/iZ8rK6Vq/j6
LAFF7HVx1W+WwFI0VxJuO0j3gLY4987T0+iB16Xfwy9FiFOXFsbMo0l2z8Lz9+aSsrF1k2nK9N/g
AiGhT9npBs2U2GBGaPToFkzU/jIgjk11JylmR7DCJ8zdC94ddpGaz7G0orxKzzKy+Xlg86G5Yuq3
nXTqAqU2J/Rv+U/TffTz60UmfHivSsqAVB+734UlEFad96pBkkAKJQJqdcvePOjd30EylmTHf0Om
IJlxkbjln2LaMRivLFmrqdmiAV9CtHbPMGPRkGE9jFdkU7Czg5odZ1Sx5qcye3dOB4E19sq9Tlec
kJa+ADVXuHPUkjxtCV3dUz3omViNx5yixfi45y1fuIZJyDjmHu65q/8xFQyCLnNKTsxkJF3687Nt
qDal3NKedN0QzHDoiQqJxa1B6Vvdwv5jglhl0phtpjK9CRrvIndsa9WKXT5zm4GY3F1YUFQSqYed
sccwWnE8VutBcmg6vG3a9PidXEvqY3RhKF20hWITRxYl+5dJFYIXAGyFh4SeFNuHtXDFEL0mbihh
cRiHwyWrvApGhzxKJ+9+hR3FYQuyPZrsief6P5U8WOHScCsS8FBSoVk2Ho5H1n/gefb07EGuylCi
/jgBuezD0oDX6K3NNCVKlYORzM59/1Q46sEvlTQ9udyzHggcH8Ci8aO1wW/AV1LMtFeyxeZ7wsMJ
tW/fr+VANTmNu6KlX8l2s7bn0YmIG+EzLjE8hnQdo7dS+OmeQZMWZ2e/ozTYgtQsfkiuEFaEqarY
AnWD5xFxBppDn+qsssRPnkRloIy64A9p9AiWftG01mV4j3nFA4zZKYcQ1LMOuEHUxz1lzxlIne/F
y+swhxUgfZepGws2eXE3ZVs0DeorzEXhbD18p9TqUM99wMAb3KvJA8QxWb2uu5upYghyJQcrJB6K
UqHpdVf5k/7HxX2IrbSA69DfkxUIiWdzyfelpiQxti/lbnRXcyZ7eTKCSziTrkrCGz1Uv8GZ1hoo
b0YzcqBMJjtq57xSHSJDykAy1gl8HqhmBSN8h9tZRqlVyDo+7TCYPZ6BwZHnYoiJdl3+1us161b/
qoT5g+gqOuWEeNRkcblufGvY54AU4CJQ/F/OaHocmdd1InwxGOjGBy7H2qgiNgtQ6vIDof71XLDB
q29ti5mTzd5ICf/uh3J98irGfYhUvMcGDW1xxnfe1O3U6dsr5OzgVO9jCscHafFxCOv83qz2XnCL
SuvD784dllj9C0aHaZcbCKYPY1hNBiHeamnAoS8UMqYiWpkzM85d9ej+MBzJal9WwCWLd7q1shJu
whsi64oZAIvgtNzndYciPQsLXYdW8DVZ9ZBfSDcFW2P/0Xx5VLp1OuS2T9HhcxWM/YKEfsV+joV4
SGX7mxpEAcM58r+ESLqppcUOzUWTaOy9jc34kBrSxHDhF2A7HhxC1pcTKi0gRzdaExrkco00JKmC
4r1FDI7VovelvYaH/7X4gDdx48FdaKk0iEMe1GHBnowlD1E5aShlnSAVU3o8PdItS805By/aqj8u
AMFRKBAicwV8czAdhZzPARWzOtgfEs+6Mm+yU9hxMEIV60o7fPnYl6FjcPgrOoBY6a0SNlnesBrw
Rc1NvRSQjerAs3Hn8Dw/kgN2EUWyAJZwAfk4a8GaldZ6zNwx8Tfc4N6j7v93WJkqkxwjCQw/XGbj
kQFBLSlb6/EqBiqG8wYY1Kbwh8xPq4pt9Tv8ZzxWY1ssbZsq5/TPX6Z2XnS4wwsgcqudD7uubYhc
Zk/hbhM+/5QdtWG5450dSvJvQ8PnHdb8mHlmVU4Cdd4BwFJ+lUQcDRt8iZtNznbTPdX0M3knAees
XRQp/74Tn5K4Tu0cThfwyNWmRMC4joHLspOHtEQs+j8ZMP9xwr7Jy1wbEX/PnGV+Tta4Yq3AvjZw
eCIMDjCiYArhikadCd5HNeApC+oEdic76sCSAt3AY+VMDRXLBOZDhbp1nQvT7X1lJAEJGAD7vzfB
I4oYoM0ZqqDw+FeXF1CKeMT4mfxaEKxgBBO9p+UNUOE/9ppRVwWdzx1JmWFR09pwW1IDSIiOa58i
ywhfnAiIaE5p9/Ju2Lg6UmJcNAr765BFKqT40JXZBKKNF2tlYDsuKDKAXLbDoybx/9f+DGBiExZE
2ZkQ4m2jlqgGD2buRIcEEbktMsfV9j5eWjCL6uV6UHVhoq/guLAr+fZfpeP8wyKeLKMd32N8cwAb
OkV/yJBRUjShiqkaY3jmTwGvaKFD/JHhEKa05f0QFQwDHO1pObm21ANXYtlE70AFWuwLWeUpGLVn
SvbzmERGDhCQkanUWAf+q09w/sA0zvIphBdlMPq5c0JsmdbK+7fkti/7sE4tUbb/jrVpewLuXqr5
BIOnfxGlflDLuLsIcSwsxI3nK0ty4jGhUjxthBfyi9UEg9GaatseS58DIDt0JNhQKNYRCgXSIMlo
9Eu2F7BpHhbTIV7N1a271KQ1vnVs65xC1Ht+X4vlN4VjNO8wO2pFSlvz8YjOgIvj1bJhse4U/ds0
vPTznCOijGAw7MvYabI7b4m0rXJoiIkMyKakkUemQXUfCp/5QqLLRBguIcoe5WmwwsPehAHTDJ9p
AAymaOTVTAlkeLpRWGCJqPSZ5aUGJo3mpcYXPafbS71b4wryWAhkckSufA9/ybO7RApM6AIrrWYR
m8dC3+C6cb0buQwp7/x3FuhQPNBudZ8LXgUAnHlEYXzdF5OzI1X/6968tSxlvAfBZx2gaQmU5gPE
KrcbEeQocoy5/M5mXoGwcoHUxRZ+3NuYA0JnjFZM/zGlvDAbgOGhv+HBfhHy7caeyZemqCKpXUz/
q5HL7D4Sz+Hyf01jZuiGdI0mS8XTLJIxBpJ61x5jpfZJ9sTYdKgDnmkjw8qF0hklE0/L4NoP3vu+
hwnzr7FIYiZ2KjU9HDfz82vDvwFMOOTO9M+Edzla1HULeMMaBuU3b1JfC31Duizwh9L6lNomFdyV
X2GynUnQUYz72zSUmsjG0lVyB/OLZLrGOkYJDxIAJDaQbkQwVWH7E/d6oHWMsOSmdci91w7uCs2Y
l5d/lDUqBcxNydbIULmxQnGULnoMl20/iiCqx3VRaQJ8Bo8zBnB2pcg1g4SHzBFJcCdZCFVS1UsS
mfJ2SNGfst8C8qls9/8IYxhgs4QM3ugpYJxSrwccG1AHICZzyV4BWaXcAHo1NyOnlOP92RsQ5BK+
Hl/tDva0IdFFU4lp8898bQwkcYOnkj2YZTFJ0qEaPLDDFZdYJBUjNwwUeOB1hLttTYleslDUFCg9
fN5UoKuQ2yBi50FqP+IHRtAP4xNFqsAluk84+mgtINiDAPJv6st1I9spcKjIjzW89xusq9AVCLPl
bneEBPQ9x4ToMZmNs4jzBdET3Grodn39w8QaTvIPz3EHS7KWuiK1yys2JApbyKTNKbWj9uGlBNt3
cYlMgsAjngyFokCBZfdByYJlpbeYNxrXujFsgFy0gn6MPSKiU6crLN3U7a45e4rb0IE38a7FPVLo
VNjUbawyKpF/udXYITVMbVztdEqAxbxUskME261+8TDG0TramPsNhZ08b4jEzH8x4eTR0D/nUlzr
P5cdQCWOLQ0qURQGTxFHSQeIkX46pE6TcJHWU3Lj1HDUOzdII3IslsL4EZ3kuRmzvS3st8nC3xtI
U/YE9mlBqEjfn0T8heDmZSmeL5t7uxEfPpGVajfTm3h8mANeJZ+l/afWK4DuCtq8VkAl818a5eEL
j6+4Z8f5Xjrkhwl7UlHOQmTVx3jwWPt0JAOQj65VpJkd/NOClyXNtkkz3GbnmwajD2YmhXr0Ninw
ON7p/uCaA6u1H+b1uIClArCi9CTLEEo8W7++eUfnjTKQv5P8J455KDFuSrhOZ/ZqL/DiqDsk3d4/
4fdGgSScxY3x6MehbvtVuSZoPMLKS4xCW15PdWRnLfpuvJFXSPvUb+FNAbFm2uSqYNQSZB11b5pr
3aPhSUuANikfWsA2rHoI5II6to3QmzPGjSw2XdMvfaOISkXNGFngdOsY1/6HNmYblN0Z0M1uyEm+
PPr5H/jyK2RzFCISOczWNf0A5yD+Kp3TIZyy1SyLht+f/j0ceFsWbd2jnuFePaYe4rVBuytJjdda
+XBJJ/vKlXsCR/9eUpf4kRRNP2KyhKVEtF8o4+7FeB4LyFCINtzF1k6D4SnRa3amMZrEe+NwoNfg
xhHzBEjHG2fBEG+JEfE0BKoClhxN4UrWvZDm4YLt0WaA1opaAAOzkarBPRWXxxJvR7vhO/pc1CuA
S34Kc87YGJUSO8hAF+neMsyTgnNGZOtCw3tBA/Q2wbEGLE69joDa15KOfxjUfX/YPVEKGOWzzFR9
jQoOEOLvwZ7HUVPIShgdMgZXQzRPxfGKcNqT6DLcmJrWIrQB3vK6y5VTRVGa4QGUXBkGJlYEm+oo
9bm3eTj5s7kZHQp2/GiddMpzJQUVh16ViD8cMwmbgk1bJwdx7UBI4ud70DvSkzXhYxaojZo3PAA6
jTYjZUO51UWv8joq+eUIm4W6mJmqsagWfvexMR/TfPWNyf32SrZILeKoBZuRz9SWHeeMJX8xWMh+
rCP2zvHTmAO6rWUxP4rWOhtujGeXF5hRQ9awMEeDYMKNLKlM6pLLJgP/g12GLJfRxTBQ+tJkBH4v
0tKsx2T+DDEcG5KOVzGSA2UtHJEI8T8zB2YCLM6MyXnvhvK6AzLollyBatYX+7YUWX0ErG7aU3DZ
VWpFBLvve4boIhc16JwxtPKzS3bgyKSkNTRPaaEKl0RKDSX9um5x13fRoh4L/M0Ff3nPtUzxsWtj
ib9AlYOQ1x3KpVTQN07/pGAvxnqIDrZbxxwCjZ1BdqtOp9FSgmtJzKOV6tAE5v3TPEVGasM5nu7C
I83HOiGPf8aN7rGxEWQ6JwmWzT+D7t84c+xM0ib0nt7PWFI2iyQ48cJpsTEcV41xG9zq703HVCz4
OhvERRPFYuhjz/xDF4oU7IAUnNyINLAxClQ8MFGzn5m7HyfXYkikQ2HbqsWrM5oFhGIJ76hIZoYU
W3p78PjN8gP3hJ9W9X+d/Cap0ZOEvBnsz+RefVo64bhBvICs7IYAy+HG/ZRaoqGNiYcHi2NbFfI7
Z5CQ35vveul/nhjmC/X89MLV1Y2d7CDN1nJ77k8VDnLGfVzq3n78xc5ClPRdPVHdbZEXVW1uN3Se
lr7f+xN1ei8RNPxHeJrc3w4ibKKRS2IaXGs3ZGz3sszJXCC+OFwjxQEjbPjJaeoTtvHsaGL1c9GO
V7Q64lvYHvttgXnMylacn7pU+eRr+HfwBn4YNhaDqq7I24Wwq4SP0SyZVSkFoOQXz1EuFhSgdi/v
sZKtlkbeI9M0O2PZnaMkDOweWThCO3blQ/oryc9Nt3f1uMi49WFyoFu53uP6cxGWrNC6A4icCRqZ
vSHpKVygyLJ5ByjH2kcQhcuLjvb4aNKKO9YoAgYq+/zaJeK/VT2Ku7REY/qwRsKua7y7/bC35kA/
1UjXRPPNnPeSOi+OwfJAFZoeSUfQaLM7w3xzVXmtybZHvv+z83MUEfoCDNGTB/5PEOwZDiW8GcsA
fcQhPXovqD121dydjfiFfjjpuY4yNZ3gSJ6m6ZUfERl6IlIWRh72qmSkK/UT6AwR9fpzN89tAxZ/
8KsyiXJJNnNcblbj0Zn53RLAmhU1Hm+Kmj96BbUklT/qmtNVPCF+/xLvZlDqkGjPMz+OAucP5yg1
/lpV7C9yqWKBbBsw8xma0COazGVY88DmbvzDk3BJjmJj4tD1klSywXa6KQmSHPR5jq7OUMCBTuWx
xlo8STPD2lzDPxm1JMnXBeUo15p97rNOiZmkQGt+eAhauxJUitOdoxOMz+hrTYQ0ipJ3TPn5rC4e
9+Sms2WxdwBKdI+xBpgttkfAyLnqDO5NX5I0TSDcqO7UerlIAuGOVpwmuZjiIWHu4sac5aJK65Kn
xcsXdxe2GYK2znX5QOYbafEhABDDX8iGCUQFgj5rv3wxXj46qHXKni3H7xgONI0vyeQ6yJVRnzDy
Dp70DNQijC79UjejeRvOxvtTBUIUa9IAMTMokiAmIZY8i8NF6A9q3OcuHqEhARWCW5awQKBhIWpm
tkL6uGr8WdjO9OO639Lrbd61GEhiW86g+2V6i0tnwc5E1PuNiUKalE2nThWKJ63TByjzkjeS/nLx
qTno9zBlAAjNW+shjGIWL3WPLrTqiSLszZRL0NuwIKlsb/kxY/2A+zNuZbgU0aGfW29V7+MUy5C9
wMe0f9ccleJYtOuSrSKa0B3upBI2T4P7JYTVr/bFuRMfzX6IZx+RwksTJU9KrXcQO3Z5SY+hZbMW
QZRgcjdo6pOzabvRVXeAdFyF/99BwzwaXdP+1v8UO5G6l7llaE+LJoE6ceRcwlCVUDKNeLLmQ7hA
Em3q/G0gpa5J3NPYBtu41Jw4TgUQwB/oZlPg++CMX9iQn5xKMZb7TdrE6PFMdNyJWsc01zQvyw7L
HdaxSfC/7l6jsK6tM9W4doy0x8laxQ9Zjln2pBaZd3zV2b03gNipswUmH7mzRNjjNHQji9gIehl6
6HF7r9zrigtgqdLrbpuCm+4xuGOXZRql9OhgIKxh7jEdqc2rVMIPq+Ce28iUARWpOuOsm3wbLAbu
ujECuI7R8Hmtjpw2/72tJ8GIqwMj2U4ouzlOiRNOufCZgDeOqjQ1C/rz4UosQ89zwOkuOVJwQxyJ
MBeAJmQNWem9YhaYTjFEgGiWZQQmmu+JjbTQWH4mmWz8aVRH9PfGwZd3bm1z8ApbJFq45vK+D8Rh
gKLkR2qXOep93X3dOWXmDkuVDdwzZIngFlZz26czLjwLeSmpP/fqKMUsDWbMqZuZnfEvnI4oMr4b
xTRHC3V0j+PJOIM8rkJl8CWafXTPlf6KBums0RZGIyy/+0moxWDoHSV4wWSVUveSwxl7H2DFtXls
Vi43J9BPXdG9JbK9kfllH23VO5P5s3GasjnYZMZzyPC/3qyy0tqJl026QJ4iuKNY5lXuxL9xizVd
EHZ58ezed1Zfuxdm39QnXJJnfYQE6e3vxbHGgxUFJn7BTNJU1KgBzBGou3+IuFwg44tVCR1kpwWz
PFRimjeOJyx3t8YCTmn6kytRyLAHoWL0lB0uVymp8fyOojMFZUuMA2tQiskRBDuPiaZ1AInwSrco
YOjHjV/laE2MWiu8LzwhPWkY9Lw1yA8tSWoANafXikZeTvC81xgS8ly6zZERSK+WGHq+IqNxaSW+
5TX0U5OSUrvkYN8A4r5MqYe0oP2nK75uEdBc/jbJb07o+v4948KDFDMHSDzv/zR4/xZPFyy6/qg8
IA0U1WMs2lRMKjfoJgkeuXd8Y7vnnKIbSUUNEBmph5pEh6g2/E7t0DabdNNP1L6AI3VKjdNIYcek
PgN1YWfbEAcyZQpCK3XWayyVNW2lm9vyWfMfJXKuKlCW6sK03NN4DfYw4KEyBIyZhCh9MyQmO+sC
axCra8Z/7mtnmVK4uBZOjExAu3di2Tno7nLrWMr03pUKRELsGa4vJrv18CvfzWVy4EF/zR4B4Tct
KnLDQCoShcYB294JdZnGeov2mMypp9sdND/8JuCVOi0TzN/ZVo8Yi/cmUVGIb35BnoOCnLt99WTh
ME6ODS3G5NuLvSgZXGxB2SO0wX+Yo4vyPsSyxMS4aKrVmZ4/JRUf4c+XmZZp46Tck4KKUZxYMQ5s
ASVoA8x9Gq9vm4Gn4qpRGw0GF3q3MZdLvc47N/TNSCEmAg7fPIG1Bz2wlO6+Es/yrXMh8ajPoUnd
qyrNraKVZ0PPitWsO8xtBBiyDFlX5xWj+58aE5uvkjUJHCdeM+gGYe00UERFTIf0bgnud24iuipk
R7TXvWqCLAsX4sJ2P0C3JbyO8uS33AYxfjEKSxgxeblXe3sFtlz2AFnKxHSMmbZISspAsHKJjzqJ
e2iphSqFKRBJMmsNAMwff7ip0r6mvMQ/eJ0h/FBaNgWipg6vYSYx4sZvxMgYW+e1vSTBWDuYXFK0
TenD1juNsl46NtX6MHfDkLWQW/pKVcThJjJYJUg99D4dPcdSNb2R6Bjc9tMsGaGGpt8B0oWB1Wah
0biopsy3hYSH9nXBEqWm6tBrQ/fu5IuultGSBVMk7U601/MxRWJh4B4USaqiGxh24h+mg40O26wu
Hia5Z3xrVHW57KvXnjRZZwhf1ZqCfY+o11VN+GurFNOSPocbhk7rNDOFe/SmdGbdtEBsIzfH011b
d2wmY0FjS31GDM42Fq+RhKTbtMlw5N73kM2mQ4UgGQpa3Mx3pWPp9jrAlwRec0I8t2qdLEO3Qbs7
/SglqLERdFa5fZOoBU8XLDwg5EvlTUw47dQDgH+FXVLLuVMo6IxdTcOJfktbkFFp0Q89dhfKJ4jT
fGYJgcv+s4nSxu290v3/XBmnoQLkQsjAv1zH8hvbMvtf+stKAqWSKf/ptFkWx4TXWFrhsheCggyO
X9+hxbjgc2655+4Fuam9cD49D9lOXDnmT7wW0zcmaYphw+yBdXy8yzO3qzPO8CGme/i/Lw6H12qJ
zb4UzmldQtvQAS281QkFUxkLmakdB7NL9HkXL1LaOmFhAsLW8sjW8ym/7PWbOFS/kWBQnPet6Ykc
kBx3RQZDyjDEturHsNsvX6DhdhFg9u5qsa0wHOGydSZphKRqlzBwa0VzBzhp2o2Z7X8GMzLnzT1l
Rcph0bNlcftrIbc7HZGQ6fbbI3rl2mvm3lzrSZ0otK7mwlP3PIxtuu5TbS1eq9OpqpmQcqa1pTQP
Ji1vksSIbdJzamzE08W7ZAUZHO13r+tusjBXd6IHjjAesBvmmtWTf26MYyV8rXpEeny7TWcXtXzs
aIGU07qLg/BMEyRum72ubgyzKYVjhQMLw3aOJWut2PM/one6ZRGlCa505NG0xXWRx5zVTqFSyd6m
GIIswcVQzw0GZ2+lxiQHIEJ4qC9x4uy6KD4AwlTPe+IZn8Ymav68fSvuNFfYKMdUWgixAsvBvD4N
WRP61xP8dcYnfPy5BCAVbCztxWEeiBfky8b1mhbAYDjgGzqQ7p/atPsq4xIuDM535FEtlv+ZIIqf
4ark8ZB7Ix+YkNmFG+JUP6ZLTG61FJyW2j8UtVT8FYy8ALtjRO/0e2xJDtnVShqMJY6juq6E96ar
noR1YU59pPnZxyGR73jAydh0CoRdJ8OOAyF787rndanzz17hoM6P+qDPhbbeWuEvaLTZB35VaDtM
uRJTSDoyJpe4QkgpKoxz9EqmA+1v47bqHzFLEXmKd5/ioW2MKGvyNcUU1oyMJHCGagWWYC5zD6XL
b9mVQot6H5/1itiAOBkgBvc2QUqc5xNbRExBbOLIS/oaP6G54lmvahHLVs3Q4fGxChrIfBOr9FrU
FRxIMjTcQFUBLalk95IFxFsi5MWn7sGc7QCyQLYuxoeI6nvaganhbFuW7L2qct1fGu4L19V2Xjfa
Wqwp9KKEhGEpRH1SiwhZACVi+yZ7cDLIj40A+1pOKUQGx6ApIWQSEEWgh1iV8Kvgz+tFHZBJMp2Y
RPIZ+M7sTJgLqFXVN5MsK816kZk1lgrdSPXxIMvbauQTuWS8YHHXrYT+yhHanAYtAT4KQJxAmrLr
eBjcQgJ9rW1R8qDx2G01Hg7aq7m90ySZuUWWzPOkvb+rGetAcIjxW5Aswuc4Mb8ZGEmvJyoXmsA8
7OVQyoqpEBq5WcePyQey8juzcmMTOq075hG8eR9+CyaqXYK7J3j8OEmhe55fQG1v5n4qrXSjSW8b
fy9pptauc7dsSXYBHyW8SEzUsTQpECBfZx/rq+t1C0sUIlVGKlYpZuT/rENuZQ/fH8OudjRdRP12
TxPPGgamAlM0tGhIj8qcrkEAPhlmCRAEWD8p3zMSRkx56BWE3dJE1PCEcP2nen5Ijq+NigCF5/il
w5aXBKIPIzf8oXT9Uz0j4xkIqy/ccYDorpp8YTiuiHyMDT8wPF3R/bBhFSlBX4R9DmIv/M7r3h6L
7wYe9Wc/KDFDBlFiEcpmEss1qVtOyQ61J8sMLtmQyHInzSCyVEBkOUaaDgVTcf9M+kTG+YRvoqMf
Ovnd4Q7/UeE/+PPG9YgL7LVQIt00z13OBBb6hCW50GRi8OpO2Mrzb7qPWyKAyzgyOKyq+WY+FF24
T0b66p48lS25nbjLj5K6j7VTfvEc8Lv/QoTumsO2mf+v8M8levtSEi8Z/J6HZOpbwLuEs8VsQbeH
R+e7hs4/DD6qxxzMb+fjGhhNCXNJkrBFNrmh/+qULyiHkQC7lFLfx7C+A5z86i7EDmT0NOLyOJAy
culwc5CtLeGm1wjpatIyLEs93FNn3snOYXDuuZ7rg/xifmsZjE62YcB4TGswxv/JlrUJkX+Fpo91
VJzllkR014iyJ6qIfwRS5Rn1W04gmOexUqznS1wZuH6DO1MMloOGm7nSQ5PCTlrh0NBoid3oovP5
ZdRZDBLjpJwkmx0QNHlhg9PshIQAlkCs5gHbYrj+O9b8WXUqmXGIUH5w4bb1Kq0QSHmedvmO5ZhT
HeCdvUGAFYmFEjzjoKPvgXaTp7OJv7YTWdBhQIGSLoil9kQAmbpLtY44Nu5XZVtUpLtDHTYcCzhv
PQuxm58u1rMd7tcmJo8cCOAhH4ZpvrAUozU6aAsFmO3uR1HiF4YjqKMzyd8L00ssxx4QI1G9z8Te
D+M0AoizLz9qermOfFcqflRN4GvyKohaY0germVua3ZlLxsBjdYqizVKnDDSkc+1BboKusYDxW7s
ICDxcEdB58AjATlOFhRNzTowes2Fdmi7dGgJz6nhY9vSqNmwukGdKDgveBOa4EgCFkPlcCRwtXzE
s++ivukOzJMB3QIhLHYqgcTvBoy/vudeJ4FXIH/yFZy5HppDkP5LvulTPtIhzX+jHdFbk8dEqbZz
SS0FDSdNtmXSHw5LdIh/jQelIBDTUmM9XkwvGZAbQV8imagjmdb86hINDCCpNWIoQ6vSZlkkLK9a
fJJFFcd+UzhI3N1HHHHZF9fe1l9+1OIjJZFZ/FnIxvCVXtVeWmw5Dgl+VMZtRHUjlF43KV12Tg2R
9SmNkeOsAQPNDbIpNhQ44aDrBxSOCIINnS7Fgp8j1+jlW+GPXqqRAsQvTLO2QBG9pcG3mmtHuixp
1oxoH5b4RDTuXyiNUbRQuwGiUs7wB1e+ie/wj4ISnB980gf4sJQh646ptOr3Upairujn9fKVfb07
Ky0PQzCPMwd//25oOfR5n5BPzMHyrqt5V65gdiDFBzYE628rsoskW/Xm0HzAgEjzQalC6TDm6DhS
aSw0uvZmCAJ/llaWiZZbaQuWsxVFLlsxZzJL/67bVvP6hv8wJm3yAsV5WlTm539t3bdHqjw9ekn/
ot5S7vXn5iIOe7dUbQVMiNO7eJhoDfVAe7RNnmpABDhnKoQ05kxmYK+/1jJlu16Aa927qYve+92I
qn3vDIKFPbTygM+hJ0xglgvKINXpwZP1zk0h1BLmcL5KEuLh+ucawiemIYDXbIs0o2JHltg4lj4Z
dzGWXMbb/TBo/Z97lDq+7GLKrrbkoddkYhPOnxxgrDGZsAwTHvB2HwLHUg82YU1V0ml8F3NWJV/J
TDQU55zVBq8y4AnhUj3zsWTj7T32mADUkoMw58u0/24Kzgo5vwbvxjXlsxF3YJagngzTrR9LAhjX
PoIt5SS9usPjBHx4uj3g+MY16aX7ZP7fF+2lRkVjwXl470UPADG5ZXgAmyOcNX4icDanC/B/gUBG
UpbQbZFA6a0TvWg3uL7GYs+8liUOMXdJZ7WpPE7MuoSEdrYkycZ45RdJ7vBBnMUtFj5ztwuK/amt
BqtFuDCeO7sJU92e99pi4SkG+sG9yLPkP9UAmHifkIm95YVPm7GeKX5t5s1MkQE92FWPj8J/UXpR
IXfvy/r0bQwKXFOUkgb61N10cddV0J+RvFD1x7qDjPJaPDgc1zFA2wwx/rlXWBhOBKdJyG9ERlTZ
7NkqhHvzRFZH4xMSKQyAWOdm97TzigzBwoaq6UY0RX0GiIQFVlDSA3swUIr+f7SxZLrma4Czrcjn
dkHFlAO+b/nIP/0hU8sxamsBoGSJ9KVK5eB13MXsGh8nFoCUGKw4PyemuZs6E4oVdbLyGJ247Qh2
8yGMFvD9TP3hhDbLKc437+ltVSXUvVJardJKzNibziVU6PP2YW6jQqr1xHk0IOFjjecs9k2k3+E1
1DnIWsx0WaRD3bmCsuyirA==
`protect end_protected
