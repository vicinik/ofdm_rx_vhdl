-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
emnFfF3nLAu8gEO+Urc15ocbA+UcQ0lu26YBAJQCgK/kyxnikSARJPrHyRLA0HrfAX61ag8h2U02
t1R84UMT82XmiA/1Indmi2O8BqTQTJeJQn1tbKzPA9yQfQtepxYHd9ApBWSPWIm84H2DRoOeVjAT
edNbE6I9zTImAsrPlwO1prt2vobgFEaWzIqpr1fyhpeHNV9k5N3BVdKzCqAa9hEQjbknOc7cbnyp
RZX4TjnzqZojZMWnb+GIW4sVKfM5TPXnRrMIIBFQ5Korl+wezuQ5+Sks7fpU0YPoPErI5yOTnLSw
xKsBrP9kY/P3U3NTvY47RmuZwBKVFd3hw6SvBw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7520)
`protect data_block
YriOVj9Fe+PSouMY8zWKwW06H200HIbxPlLM17NJ8rpHtu1TXzNJbDwpPy1gN/B6n48QLi2gu8ET
hjNDKDDkgA9MRNTXgY3sSsh5v4H9NXARhipacfogokrxzQK92x5998Uvpunu/hJxJXf/hHEGle+S
Fs8r+fHzugUZNCOZ9ncBNzwMt1RMwNIuBgVQvHIadQTP8qrhC2HqS9V9u1txnQBSdSHb/XRi8Cyn
iOU9fNAGUXEr0digB2WSXqtL/teiUxa5WrJ8+ytEFHJ5Cds8z9F/19lEl90wZsMCj/GZ98lW3VeV
BJN+NKuiQxUu0f0oFMKx9J5n6OSuS3/VUZirYXGKgBCJwW+XWSNrtD38kXoDEVzhZhF6cybgIo6/
KrtqWRX15N38b/8hTPFtsb3tnaE8FXfymtKGyTHDFpQ1jN5O2URP7MKFHocrY+zMhzb/DFsTa4rx
IMKn0deaZUGZCtKgOKzqKJohXH1YCJ3s1QL8n974YF3UXlPdDO/Y7hWt2TwsbMPJ+MHE2KbsrkAL
7FZyY4wrM6dmSfx68357LXaQTQrEkfZ2RslEudEwYKxJtOlu8HZFwL5ir3B0iObIRjKWwDNKSL85
dvjWDUk7pSx3bPrwnU4swxlVU+WZaeTIc5TXxqogHSQh3VcLLG6Q4b7VSEPQTkF0QNBzNoTcZv4G
8xaX3/zTf9y4mTVQVycOQFeDXqCsnHkCb+oz2lnwhGIf0jCGN6GjqEQjFIMvQxEp0BDwX7544VsG
0VtFbqKIss0EIsEC/XFQpp+fEWNTSyI73iocDRuzTdHJsBtacfbcxpLNnGvzHiLmMYhI+cl/85tK
ZCOzTZXcR5MnaZVZARa8V7jjFJYBDb53DaCRSpOznBJ5FG+BlBbfO5f976JBRJ/0jtX/h14vrViY
WFKSMWgnsrc4xZcMRHIxRycyb+LMvLMV0+Kvflx35vbqPcDLeOH1V4W1jbsbVGluq9W3/HjAT45W
seBF31QbSyX35ozGGYNFnh3c1s2Mk0FOXnhCeYez4sACqEqMQJ5S5YF1nfVLcjJYztsWnXnfhBkc
g59qEJrSdITmXHvUn1W/mTtKRdKoL92WVl+SkA3Ikxh7bbNmSvW4II7BfppsClpq2ySemCgRhjnw
sChglZ/oqxKZhyRRPnx4IP9tp5x/kDSXDfyAg01QXPVcZbkDyg0zKhNvFbXs3RfFrVcCHiIAIEBH
+fM0jtdgOYzmEtNTlpyMcbHj7UzvdsgZykf7Chp02nO2WJgfTo96LzfSdnDKRaffFx4nw/uHHVCN
X70Rywj9P7+fKhIV9bylzDb9RuzekLNoezty4foXVneecIJ26xW2leXnCalv6n/qYsEQFsMIRfan
jGOjyeAJBdCIUAnY/LXVCv5Elw1dUkBpdMrAw7VfbkhILNe4j6y0K8Qbe1042NdH485Z0WkYaelF
+kjhwhMQK/dzeibrWno3MHVJbatHb/CapDrj/v1a5/vX40R1/EGKttLBCTlEMGAUImCGwyHrDuV4
htIOO3f0ODr5pYalxmzo8ZJJqUgDOR3bkdzPZK/oBnX2uDIku3m4bhKbrZdxX8Rky3waQS0R7bQn
nPanUpo0jjwkvU+GXPrBvbdKdd0bvRHn/KN0P427YN+6lhQ/M1+zv3JEIFvEXRwpsv6W89sExI1P
PT72nHUebRlmYPu06YeOt3SPgmfzFBL/wJDJvWVqIxTtbwx8b8vJ/regAFXS8tcD4wdF0y/u3m0r
WoVdTA/+d6UKRI7JN416CKEmlwz+I4IaTxvnmhRDJTQphqBGTdpgUqQZjeovuD9FfExejN8gElW1
7TVQLF6jSEWyYV4Fw1fQyAVVw5gI5GCP3nW1688ZOAoz7d7e38m3UQhMSHen7Qs5939lIqMR4gTp
vTpRFNsjIS6YKutUAlbKfitr8GI9W30toKnqLnjIwjwULVJsuKdNWs8fAbzrbxoNJ46A2keShkq6
KTOOpGkVaGTfXH8cwmS3koABm0ucF5xO7N/GXkG/mlU3tlFD1OH5vuVDkvZYG/AXH6vSFWf4jMWV
xT8VrEnvBXWJClA1ErYL7jycLLMnQ00NUoAY6W+Lvki4LpiRBVdWD/vNVqFmaKwNat9zY0hi08U0
xYMBwvcebQsuZKLV1M5GugB90mesxntKAKw1iIord6FhKOQUI2ehifzTM89ptBYfV+8Swra1vKgc
EvmKZgNF+WuqMHP1rreB1x5x9laBEVxoiEG96mrY3JsX/+xj52NLlcylolY07FabBFX0nWfhz44j
UrHhJWTMAfpcBxR/gQBqSIcxha1H2Kq4al9aQkHfc7t5qzNWaRvwt2SD/PEHR0otVA4Oc/h7rV87
6qReI+/L1RXjfr+yBl03Nup+BEH/xIWWR07OqVL7BrFjsLvvkbqjxmek61PkanrOA/JhDVpVBgvg
7Lfd7tQJZfhbhTWdvYvpBz81CK55uf1H5jxr7SW86j/y9ukHu4s+ZNHwMVOm8KrmHWn1C5NlD5Gx
PxGkHAAs4oQiWFl5lHeci524T6alvVQQGVgv6O/odd2h9kQbCL+77kJpVFPEb3sEfBhk9vmgdsWh
KyUSv0ZCrd5unGjSzCKqGiImtkMtLuZZrWKvRh2jUCV6UTUBvA7P/jpNs6JF1mdfJ/piGWW2iGvd
f5P3cDPiTrDGyB4QKW2lBf2J2Qt0aKC2oKFE+ntWE9+cJxkEceliHFclQ4yIdilOlU0rWs3VbwsM
i059wOuCXTPps1lPW2h2NKttCf1G/yrVG/Yevbu7NNpG/HiJaJyX/leVY1D2dqrTjwLyzAFDAJVG
1xEAGmwA0PgmVjdCHlbQOVclbbLTO1yvYpbvHKD07Nx6kMeyNpCuTIYOmNZrO5RqCb5dR42S4qzD
k5qk3Akxd9BuBQCJgEkylhTO66S9TMBSuZZMJvgsJIzo1Pl+hbDDo/qFfxmtfk7j71SxIcLiIrF9
EngoZ2bfB/nnLSbCxklng2ips+W/NQTsxJmDcrSKH8XsbXWQ0eOwHOJLcvtDgSsMmC8XtapdEAbE
a++E2pGTIIpV54rheq7xvGawm4V8AbDTpyH9BJQ8kbTnpHgCqvuUcsX4yDC09lD1lcNrmODUpMpL
1SPpgJe7Qr4r7aTl3WPz/C6+g15rFkwktmhreV8IxKl+kLw1S7DrnJggCHTu8uJG3vCjl0rm+g/y
pmAGQ/zmIFhKTnkfhY8MtG8Z00qfAnHbqcWIghpFFVvPCUggPTS8pPNawbnozm+BzFBjZUv4+1Bb
ZqtjjJ9qEzEv2MT8iRyVMakrK+8LHRjdOFrY6sN7z5glocvWwbtCeXEHl18rRzz9nbi4Jo3612a+
r64B6yNRRbMKdSAEB3UcLQsroMnvOrrPafc5x1FaC0s4CA+Ey/+Nus16kbrrFFmQQm+lxUtPk0vc
7z/hOM4kOsYrCaUdbo/QqtnaIQgNVBbiIym2pNJluIk05BMHMHclIc7YdW5fr3uuUZnajlurwbzW
Jrhfx2Ea26VyyqbO+LZiXpuHXN/s6kDn5y/6OGpGc7LCyLS6EEB/kFCcrlaXHlgmRieYM37IOG3+
Oa5rupWNlhL3Wv/MTMYK2CT3mKcgnxRlqJh7VlFFN1poOU69+3xLVmHwDkqKrN272v1il2N4wRFI
JSoBMzgB6U1X3tekirADP/WWLgMl4sFhp+Mm3R+oYXdnBMM7i7NN4/gjR2DwmQQuJEmd3JttRSNy
W9YeqBiIh5vUCbiz1ummxPo6tADutHVMTRdV1smXIontFLjzXuC1aA4fxHQWfcNkBVXnhmKlYI2v
tyaVJTf8Rhlm0PKbrmL7ARkQ6taCt3s1mW6Py83eK0Zjw42SsbdLmHsEVDFp6PZiHGFLpP87/c0z
FJ+l4HqWI/DNnilAn+nm/3o+ffNRSH1JKP/sCcwgsezjVSyLa48P9cNldwe8BN3phhOMvTADHdeQ
GBgUI9lx4aXz/TMjpjf9jnvd6Xej/wk9MRq+2PuOsVtd5ApR/TXcWOrS9TfQ0n8emM1jAYx4pi9M
k47iuOxWTVSceolJudkcBGoOZVJhzowH7Ake68/+peP4EhQjBxFnr3522Urv0tJclgo8R7d2Wnny
tJQz9z7654LlsTgMyv93Qi8uAiZ2Qei9etWyrdJPn1Vl8gv8pFV71lnxJKg/NEDfoiF4U4ujTjyq
AWVoGHVQLLSNYiLaDBRN8PsbzFal2ffI++te8n0E7k8xcCKjGoY+y69qEHO3ZaPERn9Gfv9cJRwz
8D0X7Zy41cptZ1SiOdnbDFOkPpVnnZqPlAXwgsPuwaEH4QIXNKoZC2DHy1tUTjr2qEbTMTTmnnxt
vWPnf+tYniEWFLG3RtoOJGD9V8SzQXmv3d5g0bFKTZCWoGaoPbBWHtOf/O9GQTzpEtGd2RhdIF/L
dcmi2CKA0tDA7JoFEXSLFmF9TeJEL9PMpgyUsE9hGMJROBB1y2NZQ88QsVMzNJQg7KSn6d4K2H1K
Ib9VWjeMxFh977mCVEFZ8RTk8LbojmAQNUTV/ecBYqBMzRo1ZgdkoABDAFCj/SKoFTy2N9LqL4i9
3CbWVZxojitNrpwr3Lx+52YwWoH/IaqHF4FhjTB7VAX+Dv8nsTjp4Z5UqeQ79JVHMcfzbhOcqUYU
7GNUXT2B4F95dMd6SizJuwU/Emh7LYe8hbjNqyuIN0aWiff5karOqoaG1VX9SXvfomABKSQxBs5S
DN7hYPo9xXNA8n2qcXWf8+ymdb9SBzCAmyzLSQl6WfLulcB77exnumtJemKRbbbw2+2jTgLA6MrI
LGgCSCaj5OPOZWv0ysIvS7O1v/eaRqepVyeob4IY7+Vgc4cB3FFnew1tHd7T0Okke+Kz+zuQxJlQ
n5LGVizgjXnvvUTYzLFSRMEh4CjkqiS+Y3Vmejy5GZHEkhgzqeoLcCCy94QMfAx373wytpik+Zu3
6PLAxfrM3CMiXZwfoaG2FMG+5R/38etsZ0vnJwJ6Te7dCvisY9fEweVAVTEasZtheoFBaKlyxCgf
AQhLzicVE7STo2ULvW1ZvFYIq0GxGkZl1x4jj5Wr+Z/Dcx9BSNyRnJwxDzf3ctH9CvMMMlRE/Ew5
W5Qv8Et9TXCeUgGjl+TuFp6YAl2ZiMJ+NEbxzDGg+PxSc6cn5FShJXK+LTb2Go0NC0eR9Nk4RoqE
M2BZtro5GUoqMGHsiZ9uS9jx1awPE62fn3+5yNFeASZ72bXfaHZ73azyf6bTHeOde05PNBwhsBV3
bLmZRUpvi8GcDEfA51GlDOfhg2jLpZV/A03A1ajYZBYDIoE3AK+ZIoEdKN/7TpkXXJQa2AEW1HIG
/h+zU1TLYAKcjm4IbuWKdnVwG2vm2AshmbFidDV0nMsRz941jnuNrMNoTf+qmDI4s6eCMPUPyYBa
+XrJP+9/R0uxbUoj47wyvWrTHMRlB/7mQttLGuBX4Jth/76DnKEBYL+4zBjGShWNG3EHfTZay3gr
YoEk5L5wSsyAWDLBW6BOHAsq/UVYT1ESCAoihJAih70OYZoDSIQPuyBXLFnDF0hFIDsRj7zJMfnB
P8zm1kKu9ChjOvz++ZvlK0bMyonlkNPX8XKkfAWvBJXYQeR5a6oMbYM9OEwYymmIubbvX8A4uU2A
xcidd3eDuas3C9vuTDK9OWDUuwhQOsdRsf6ZvmcPvWMOtz2e31yAX9Fk0uxkMw1BYGVSI/JftIjS
FwJn9ULKSaFfcxQx2RRCkFqJ21Ydajuax2oB+l7o48wBMLz5n8KM/CGQGPHEloVcEX/k90gdG1he
D9V4ctrDPqr2gcdbRxEJDPI1opKKEw7iPJj3FqQ60pxBtDMAOEeOGFQmgWVEtkeFRB4PYJ+4GtAZ
2bfQBwOhtQmg33mmTaHhZnrmmcBrDL411Yxhy6xLwc3C2lFE3wqgChZLqsvWcqHHddXeEssIvqbd
omFbJtR2KUwdOqUcItogvUDJpVYwBJ+hJDD+/MhIErFjsr52vCRtjXAVYe17DbEyC4p3GkXCxpYg
VNvGdHRqNYvfvB1/fk1lizjKoff3Usob8L2W4m7VLAAypvSk631vmW5PG0v/6VN7eq7Yjzhuq+04
OQ0DplR8H7pz9WlYwCEhWUQBpWuwP4Bpndg9QZgnZIGDwl+G8Hu0urfEcnnKQd0j1JgABDZSqVT+
eI8EUJWU+nRAg/x+Kmwqpel3hxDWavkJp2LpTOFmlKv6GTJlZfh7LBxGwCyy2dSOXU4MNjCsnvN4
42ZFqm+TAW5WQl2Yb9FRqiKmp3ENuj1LGDYkRZv2+sGwlRB6OtbtdW9iOl0M2JjAci4NEsuSqNuW
5SlMdCaiiUdbMIeFb0YH0yxbMvoW5doabeVhGp+THu3hNlna9JyIgSqi7zTBF+W1lbsWDHGyGNjh
+gOR6aBhHT1l7Uqb7/MVtSRBVJC0PxIU2ZYOZG0wAwMVSlIOP7zPFePYeHYj6CyHCI9sJCPOpF+N
GtrXL0DlSLyzi9CEQJztqzZ2VmTBMhOOFe7SmQ9/QwUEYS9yEq+HKNScfQuXsDtrHwX8BRHkBtVu
ChqQRKyXMAQhzW3ElgyKtu8Oofy+SNVOKRpl1VbFMYDsQHZYCwonsda/JG8E1Oe7wyGu/NnsKvmO
QYVa405qU4jrrsNu02LIGfa9fyuaR4RgHpxqgcaTia5zja4Tq6PAWxnXZMHFbuuUDN/m/BPiLa5c
mf399TD7exsDRXv+tkYqe1n6uVSggkInGLa0BakIwjtNJgUZiSGV6s7Ek7J3VB8pUmmI5GbPjDfs
aVmDpSEucb5L0F2X/AaDIOsEoyA5ti6ivRft3BDaJ5XEE5Uvh8gvtFfCG2V7P9fI0cb5WF1bv0SE
SN/Hkt0nh7szLQB6TeeWMHH7mGIpyE92RAkkRZAYH82DMrJfjTqGYGIzIeKcdKx+s7rokwyL8Uls
x4QKT1Jkj5mqhvWGcGfO5OJPMunL5F/GBIJDAZ45iDVBWOliWB+N6l8WOZbiGKYbHaUDZyVMQVmb
Xl0c5K3WVbmBib7gjV5nk1pK27lpgZy7xXhWeevtPyxgSW4XdPPT9ZlmGIe260UVW2QM1ph+lFht
d1WTxrkKuWR0rj+TlcGmh/MlndEjwwRjEbWASz+dY0jERMEXn7iXTrS95dvCZPjC8i7PlD8JuWFa
SyYwdzKFT4KfDEWgal+Gl4cZbb9j4g3swpYjW3UYYq2yXjnu3Oyd+XwgHtPKSHaVm99RKOXr4AJB
IzlVr+C5lnQiB5eQnPdVWpw1iJ93DkOIRX2DmvXapITt59yt2vI9q9HWcTThC+m/X08VAZ12ylE9
aLS+VpEGWrA20gHiHj7DCONbrnGmzadUHBDZhQJv+JCGKqKixb4b/axBVsc5zvxj3jhhHjO64pld
tcBk5WNfvLGrEXkj6ncKFlA+dmp+BmHuR1KzOgeXMktbWUWjHIbz6yke3I3Ryx5fLlu6Umre3FUD
x6+XgulLMFihABYs7vKrdY4Ic2t9edzfhheMv2G+kGEMkks2cVekNIj/LoVUriZMlhcDrOFyteed
74M+culF1ENuT68cMYyB6qSc7SbA0KUSnOAFlaetACFDl0yMZHdZTNeoq++G1QHJBioyQJhrji4e
miYVoZUyJpUR9iOnRUJBgPkeDyjLgEtTIAhl2D1ceCbnv7xIEAhH2BLraFt+uTqIHH0Udq8jyHRa
m4cuK1eQv++z5Yec5y01wyBvvl80wly3HmHl05gFJ1T/3tPuyemZXsOctyRTOmdYhQl0Vw/z2geH
8g1Ao3qrLRT03tnPyWJFJ3IXC6G0O+p9v1BVL+yp5SVibiwQoSO4K6SFmTPnssAZDd2ea09sFhCn
WSBStPLBzyBiEXPe5hqzPoIKNN+sMtitTD97/aqTVo5SDjeymu2t0ASfoHfVgm5Jo9/2bc7opJLI
9hOy532qGJPCcg2Pk4237K0qM6hGrSe19Xgm9beYUsGVSgJenaK13vs69dXT3Qf9JryKpvdp0+RT
HVhEeYajuuE1b6VEIyoEoKdrM9QAE+Ti2l4NyWVeiwHLVhs0oa/meYe28XFrsQLTaaDw5LaqXwx5
Z/CqsTN6RQRzjdXBYQ17wGJ6gefQj6xn4Gqiuh1sOq3/f32lWBQNidf5x+CuRQXEq5bP6UnW0aqb
ZCsVTUpz77lEC+XHZhkEYXhs97F3bc/ws7JuGgk5yD8H7XneiO9VEDwstuJzlRYQUisSLBELQn+5
NhcO15GX4VFYwFJG1f1xjx9kOFjFtfzPwfcdPJCfb9i+PYv4tOHmu6q1mYkYmZXvVDwe2eZV2kwV
ANKqKJ/OX29uT94iPxLBXCED9WhQcwYU6U3Y0NUWy1RvrJp/fFiopPkRt2plO9iWUoZ4i0njQxgu
OUqA6448nlTjaIQoDnZPOuYofniLRpYpzziVblGaSeGtb9bz0JUCL3PaY5aKSwxHCXIABmDzM1fo
8q8sNsIkII833CSk6cxa0PsA2Kkl0pbEsgdTOiL7QkwZpbyGMLXjfqennxyTwsiy6vvT+v7Tv5c/
KPttvmW0Od4+PynUsMmZ2pe5zDhSE8UEWGWUiuUo9fv8L3CXzu0YD7lQ0tZoZpfyxUOMCeWhesUT
tpgpVtKMmVr3xe7+zSfQzLyJzmdCvJiTwdlg/6OAuKqqzUcgeGfP0RByny1UtM57w2uYNH5bqaeL
04JHgQvR+sxBOi2OnmaysYr5/vAnNB5+9JzCBYjECEhZs5O0KvzlOkXAW188BVsuqXO2m5gasPs+
PTwKbV6w9SWdrS9LYLH4j9S1dMN9CCmeZcwZrA7rEsLObrY85rdSemnsLTQPwwuzByn7WcfJO5BA
Lyy5M+2xzSssl/5XB7KL0wcIFM8976B/clJNbewH6FlzE4a+lC32TR0bgmeasByacz07w1xFuCFZ
Wh/p0+GDFz9BRGNTWE2HShxfxGmKsKqX+SCHLyhufuYQ4E+4ySUgC1ZQ3IDgbWfZu+35RqLZpy9u
H34QTlvgpXW/V4QZv6qgO8PIukojh9Z86Paaj2oLgHuj9DGyfzeYG6uzvaiUrZ9rgadBr/yiJr1s
ARnNzBfuRvCmmH0Z587HhZi+uvd7FPclOuVks2uyuONGFzSoXN1V8DFwbrVcrg/YEtOz4vby/NyC
CsZkGHX5EOKRhBBqydUXVGkq04vjlR5fqIziOP2V4o/00d3TePALt3fYvOOR+Jx+5ltINVMJF0hP
2al5jzFzntmW926p7JnBOT/XiQjULXKdRTDN0MhHREkdf+PD32r9Tr+tDg4TJTtjD8j7L6pli7lS
CmzRnDxz9aLAljj3+o4bN0aGiJlLOhx0PeZ/bohyWhVo+FR5LgNZqNWGW8ysF0T7febn6KYOKBNe
lsPY6dDhRPeNRMv1Kv/6PNWz5ctNV57XrGrXjvGgjAWqoLCvWbYfzIUOQs6KRO/j/aVx8H9TjG1V
OH6lX3Jk2dQjB66N1E3wMuh0Q0ILdr9yIgLeGPO3Na6aE2BHVI9BYAxJaELqbbboxMTdcCAx5HwD
xC5AZENb+n4TKvsT7ffJ1Ihol16UMfr/6WKyvxdrm8HTWcniuGnwi1Ybt2pNpOyELCrEYhMXMmm4
WrqIRlXjM4KhJ12sPCd0xXmJIljgVJx6+MkWw1s1AtfJ+y/7YEep/eiSiH1coCL+KvESdVEFl6UX
pU9xAR/2jmiCC3f4V3/2PRt0yeWI9G7liiW7bKg+rIcMI5atjlS0f1u5Sbk/8z6ZyKd5xSbv3aQ/
JWteQdD05ztTxrDqEvtzZXGCYkRy2AeVN+PfjrOTiXaaDl3WnfV4vDY+APBepKukFPKcb55YND2e
5XIACbtRNnaTR+kDDraecdnoGDtDgEc3vMuTfvUNZa0lt1d0+vSwfOJPkhlDHVhylgX3q67lfoEE
ZuQtFyb5qTOre8M1xGlo/uDT+zTM4UJhqPfpKD9MfRXvckiYekrytNgpCXqnU8D3ekxQTsbiGDK7
MTUqa7O7XajN2sD5IURpJRdoQ8CkItCfr/YrvEt7F3M2mQJdcZjxR+FRr/jAs6X0HTtWvQw=
`protect end_protected
