-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S6p7WqzDpg4yI+DjAx0xDZGLAHdWRwgn7ploNxcrF6g8HeTKPyZrAlOdw6ECDJ+/cr63+6JXYa3e
zIcDGN1otGD34prLv8je5UwhvTeC4Hu5b7jWH84V0x3YnI7yLLjc7sjPGALnCi//GI2Nh7MRk/jM
s7BWXVEKmViWkqoWu+WBuprGYdVWtYCYfq336iG8pzsBPDAA9Gml8PZBTII3rhVJxKi4B6tdo9nl
IsFUAWO6vqA5l+kXw8o/UtYQIMyld5XBpY0bz0I6A6qR5ZO9PsB3CkARb2qHJewdwpp+Aa4W8lyV
ga8fYUVz8hsTtIiDlEELSdlSLqbRopgQDzMCBQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5824)
`protect data_block
MQlXpLWlycDJIhJQ4krxt8Flqzf8cUuoGVoF2lC9MNhZ9WBr5+7L1IhmDkJi2RbKu/3Aa9STCRoM
otkBdewv9Tu1GHkqJEp/bat0+H2GM4U2YhZkg2z2LMbC4ay3oO/gAyqj2LOeNDzRrGS1ZHsIXKex
JL+Yb/nUxbApXtD7mg9GNNgSxMtkRm3RrdHwIz6O1l70Rz5kEtY7UUBraF7yeBjBnAS6Ybjj2w6M
y39mOd56NXlYjoKYBgmeE0JYMGLpStrpNAiunuLNB3HUBZNKAg/KXdd83sKyIRntFbd9ZnM2PDgu
r0k+VOWEDHifgYpNUwKG1Uryc7I1vDgd3fPa1Fe2QNh4HrN4ONFq5GZcVJQllS4mGrreDY0vTGtk
v+5lR/KWxD/blEgrXC/EFHGcrTr0N6g5voOzO+BGyg9ALeThffJDxMn8PufqZu+VpSfEnbeeLxCK
y/62w3oeGX75AAYLPdsobD2zzmKCjNTDp8vguyKTa9uZOpfywbryxF0a8JTi3vZrAt0xGXy3gTaN
5x8Qg/AzqI+oqe/sjUgemZCNSPFp1nW+neaMcYuRcDpqwRbByf1fiHgJ0kPXz/IxA0+DufHQzSDo
2xtgPaVmKVST6PXzn0WYGgVfuRbo1QLNTvJCJya50XtJX2/6oAGw5leCyT8COEHveC+PzFEoWjtA
U9kUCPWVS84znh3lf5/c/n/u6D5o5l8tRZK4USHMRPBpUd9jAGtzNgNbhUZNFgaur9ls1LRx4JvJ
zrwu0YGlRWwemq4aPpKOF4oN+KgJmpRkyidXMnOd1IIlq75RXSQNk1Ccpffo5dTwq3ywZ6SS+CyE
sXLbywstE0gs3t7Ur7lMTwQo3o2AfQamolp+h1BGoOiSAtgspbTQD7TxZI0+wI/5AOzLf1XvWg3T
mK2H4V7GU+aCTQOU1hPnVNCosMjByoxzqnD7/IHK68WBVUMYJvYshexYbACgOrBHiirfb7HUSg04
fRcu/J1pR76gRmwFOTJ1ts7B/FwbV47EZ6X+Zmc6pd4vByWNXGBv6UBlVegSLmTFOIWJ08fEjn1K
elMZ+DMngsTYIcxPFCoypKblQsC8ijSMCnUCwr3/RuAjH0nnjXQUGD+miP6Wj0IC7QvXHVDwlM6o
xGPHpH8apWOQz0RAOcuemGUGgkBVUeDe11HCWHpwk14eyrDXzEnmRotQbpKOV8JWG14l+zQ3lS3r
71e2pqd2p+AdaEbJ4fmhdr4JCzkGhvfo88/Rmb1Jhk9SsSOGixNSZBcpoPOBNPHy3AysoSRJgS2a
6Ou4XEw1hPrzgS7pVGB7ERrTax/8mwsWQa4i0/lQSG2jyH9Z4q6WYdRwnsmi3ueXwAAzNnUIScGN
kvf1vr55R3Npm/ST87muVlzb+DCryQdRZw7mjP+gotxomH8ysi14+HShzbYwky0NUdJ5zOzO7npF
PtDVbOkfnySCY1UieaHakBFJ+0d8hn6cv4+4uqLXF3+OK79cEpmXSUZjH8Z1Bg67H+i61aM1KL0d
hNpuI+wzzbKaT7NMh+O86TLhpVmf9p1NM8s0A4L6gvqB1MfDVmK2pohtMCWapMS+4N7GqWvimOCK
5RbznU1Ub2ywt/rejbJRfgS7Wlwrh6mgJ/A3q9IFXQTJuVlKI+k/toU9lmI3SAHNxdh9lUSxktBD
8gXor0SPRlA5ErzvyCnKSfv5zOM2Rmud6dwh5lWTdEWDcVEQTzNb68cmEszNtPVxhzb7sGL5B7Vz
XLl1HVDnZ1ngpq3Lz38srLTychqxlX2C5NDq41HxvEYIc1vXVZ1ijUmGmPRJ976C5/okDbHWVt3B
Jw9KeIjRrbxtweJlok7rSftILUIR6jL4BF3EP/J11rVsBzC7vNLqxU+WANMLYe/SDr3COVm4tnR7
VeBz+psZOeLQExUH5Uo5DTgWahKcFaJ+VPAvREWrhAL367ruU+ZrdfgyCw3Hk16eALLRqMZIqX8A
OOMt08mlfryNtgke2YBfoArybmpV19Mw5PpFnXiJJpA+rZBr5FHrcb10D6NnrWd1Gfv3OhMBd7Qs
DZ/NyITDEBShgJpkJhHo91TgUL/ALwCTR66JO2I2GbHKHcdTp+FA2wjX9GnU5r2kLkB51PV7dmjB
2sV2r9bZ1zCvgahgKPSX9pxnwTL/eXAyoTaHRZSzHUA0+wmNegM0tyyr82cQoRo9siwtjdM1nLhI
kuc72X5S6k8MPJ76GuhMbC912zsnKzYIUU9HCN58jO8BHUMF0W/m6+iBJWCweRIDvCCnUpiGYAN2
Yo7dw6EGx8XT3FkFYO83T8LG+BfdInfgKZSeld73/t6815PmBBiby3VlZlBbrAFhgmC8JUNjlSFd
+hqTDibTejeQqFKfIvnjU4EcdyJkdPWvP8mFrgaDLH+k4Bhjj9zeeDy8nquSD4CC0skUSn7ATmUV
HXMIoACq0Y63tVqGhG/pEP8WUiRr+M0tcEwh93lE6K+Zbf8idNbwISflQR+oycXJ+9APuNf5KULY
0wXz0Zm48yf0crfNTrwT0PhRB+dpgIE2Oab2tt6yoakADj0afaPAgHHiF/hruzpZn0jwQ0Z2cB/i
FuXSSlBvogDjCu/VW01HzgGRMKroky+pXZcrhmDIMzwLfvsdTnwFmLGW5/N1LMVqpX5kJPUZzX8i
GNfNdRyDZs3DLkl4j1eOHGFxPPlTnE0d23C2iU0CROSKnOUhn/BOiHUdGDtG5S6Sh+W4x19IWofA
UZIyF9kkQsV852YRjkRwp/SwN2ftiz53nuVNMH/+Xhhisw7Yzhd6GvUGt+RlfWXL/l/0TN8ZiXUK
0j6eq5leYuhQ0H+Q+jmAhn45xZiva9vvqXqiCz5HII1RgQ9N8jy9DInYLNEDXGqtpymWgMZSXwHJ
/kcZCUoxKEav2RnPMO42l2H5045CZ7JyeU8BK8ivPgQ115twNMrG3hHWAZyNwd6nXFusb5xPTP4M
covJpwsYM8CoLQ1dAFw3OlRFxquZ2TjwhVvj7HiywU92aK7STdxqFIEieoyFKJ4oWgBoHma65kja
9aA2VhTTPXGAdD0Gm6OAfJO52Vfv+ToOm+LNtUSTNZzCLXefUQRBvqJg/n4+dxnTIvfD3HuyfdDL
Zic8ILKV93Af1CTzBRJZlMlgg3Ukk4aW8BK2vszu0FhOVeJvA0PEgtzKReYqa1urK7hYmOF3wIpF
SIe06wRBCQoL3kgJul77Tl/lYVnTr/ECIdqPvwiuNC3T2T3JvpY1MFWjrbgplGu63DPHlWMWuCf6
wQnnRbrCzrbKjYHChjTbbI8IBZ6s4D/oSZzQXSlZUgChAGhq2cj6cWshGkWXUl1/SYZ24hqG75+M
ittSPQTAWKLFcOY39TWDEMAeLL283eAbMlc8Wz99ESpbIIKNCz228fHv+uWqvCDGtuu6WMXdeeQ7
yrbdRS0C0471qSFF2FezNXfAc8R8KtnhlcvMaMV3x4/QdWMDe3V4BfA/hngvhQojcLLkGIdB63HY
RyXegWlNyJVtBKh+Nk5Qz81r3nYVU3bfVTXMheo0OYn0o844Lkte74pC/PZupPhWR0hJPWKTTVW+
MgOEdtriL08XTn0UHuARXAEF9IzqlRlEKyrNPKS8S8rW4b2PQ5AS3sL81oL3OnpxLLLlnaMseefn
jGn1l95PZJFuERKiepB9v95maJeGvskkW/jXXocwga9JIAXA4RkwDCG9KPTcZjOC0hoEQz2E4Gy8
8kCejG+NqV3Dl+YqhQC4oiBRqzLnvX5mgvm0AkvrMfcMlkR2x60HFwtBQt7lCumy6RI/67OrAupX
+1g6lDr3/GP/5keTGZYi/C9sna4gB8QZ03J5BljiOv9K/g5p7meSiJI1ywgi8cTtw2XaONnhXry5
frL8Cykwfq31wPr1UuO8dRXIWpGParX5TPgqD0W1USEOtGoU6bWTS1AIrEsee1ccCssT9OMhTfps
bGj3VpQxHd1H82CjQB2qME6SbIXJiaRBiz4Mq66YmTwqicrmIKfUmETrra5Ri1bhilcaUIYpkJSs
cbvLmWCiZjI728ZcevImgA9LLoM7Te/jaXUjiZMGSGromF/FhqFm83vesEfRNRFDGatV/T6fsL2b
sDJuNYdu9u+0IrpMVC9u4Bwf9svarZHIZW4HwK3gnoC9Y/f5zJT8BDbh5k0wveAKDbRJJMG5+10s
V3e6Oj/DeJB6egRjvCzamDIdsAqHeSmEl93HS+lsqwM0N/MBDGffZbbg9n5v1Pg8gyeRUw5rlpFt
ol2utLjeo/9DV/RlyJdgLHTGKEw0rK3BpUrA36EmJslAM/9iMugjcWgIraB2G+3au+wIOZlzTRwF
PPWtc1rxCXzjdFiL5izwQzEC+K//CpfyM7roCFiiDPi7eTVVIbvVwSdTrYUP8pnD8pMsWHXElWUp
Z8mlvBtZJQ9qGyabrY6IZGAd21e4mXf0i3Sm9X1chBj5YkCPuVDZ+F3qS3LzfNkak9l6bAqD2keR
V6WT01HChUKoypgK5Q8neNpEoND40TUAVYuobNknihZ5vSYgplq48dBwKSuvwKSEZj4HOpmEzaPw
lU6xcJi7gfTjvmpzaH8qA6YQEEAHDvRx5g+nLg3+5H+HCh3t7JyhxLRFfvwtx+cpafP4Zc8qoZf4
4mVNJV7BuJ7UlzcX7D+TmMZTqZ1EXEbRDs5EBy7yONl8xdhQk+oB6znj2p7bXwVrXPFeNXR6OC+X
2ZJ/z5WSkpC+8Hmedy1cKIe/OWnzShoIF8CQyANn/IGEnlumZik/Es/oTsHebN5ctP1iB8OCgVGP
6i34cj8iZ+QX91kXaMgsVVC/Se3Lgg92X3vzj6ZrF73BhR+BjXYOpAZp1eliqFsW2xLRk3LHVDgw
ozZarrTS4TUI/AqM2aEP9vUV2oeSzshxRr8cid+Ynajr+LGlD5TQT96hI0vpH4ky5X8d4EKtbQnP
VWT7abRIOTxj8GFpMq251sN2xc41R3rjSt5GmUisWn0ketpwdGydn47TbdetPYQYVdj5vDwfYlIq
RzxGNMxqEHl1sD+mn8rvjcCw/b9mM6dRp7uGb7GSCkQtmPbYF2308czWQv5GlOD6ir8fe1WOYhxp
+Wc+uspNkmbqWwMUafNMShHWQmyzocKgUIMvHRqFBQBB1We+5P/8sA8SDCNJREMEkwDsQ6Ubg5Ux
06etbW/rkSrgfFVvjIQsNkYl+JV9diFx+eWju//zi6UJHmEQNXjYHCn0wquY/dkfIqm+YciLPU8Z
feDMMoyrK+HOrk92kmVgVLndceyk6ZowVVADeUOaYJBsewrMNIzqA64KBrvuVt1l7g8JrfBUY+aI
cSreIICPtjkCWQcv7znnTVk1GBfHR8o/SMpUk/1kyfNfwN8CI/I0q8lS+UXgr8ff+iNBeYF2uMpL
y8FsADBAjkKuEIyd9PbMXjJ9CMlf0wJba54RDuINwk589HcXf8lyErANwtW4nMdmIDggirj+bZfR
TFn0rDfj6ttMU/JQ9rG/+OR6v9Ci7Qqt8fa9G8xBE2JHyPpeA5gztvVZPemIjZzn+0p03BgFme5o
P9xUxrneaZgSOxO2lnUZWkSid7ZSqFOqR3XLNaBJr1P8x2nOj8cL+9Nejaf1dypP3/Rdhz+aSB2R
rlOXqGvAliw8Q2KF9kd05e4/TjHEH0esHZXHyQYOt0RFg9jnBOhyvuWAcY0H3+VqckDW7IcLSQdg
Uo9lmnaq3uH5I+rD0lYoiPbrLyKvPwRVO6uD0hxhVmZXRwC7quFDdxL87iAQigD3NCk6iYoSTiBR
q3B26umAkLduHK4QL5GqKCNaMu5ENXqyXuKLixDtzEpZ+JQo1CXV50h2NWfZvrHnww7ID0c1nrKZ
3lXSMQPZXrjFpV3iPiqJVbcomlkNJq2BCyqPnWDVi2z2sj6cYtqDCqKECEHDY+5G+WztksRuAy2O
cOQgyhTWS6skJEJsHT/UnIrLZvsq2gcysN/9Z4iBauZN/udjfVBQ3JmrS4ATb+uZs5Tjxt55l184
ekQTP2XDx1dYHAH2eTHy9TEcC6JTJY+X6J4/DkbB6TtDZIHfFFH6SUIx6GhGl0AYc4rnByngqXYP
lREkqfjTKx4JEiATZvYgfFp1DSvYhb7OPzyMjF0l9j9t9IOXFkujZWsqbOVX+TC2w3CvdgvQFhDD
gX4Ofz0mH317w1hfnqenbYZNV8LBLQg3Pcjffz7TE0D1y61odJ+dXrMvDkMedL2py3Rz0/xays1/
hqqdHc0e7axjC768skWHvwAJTy+HWwdBF7e0XajySez0874nPI/eQllMZA1zTI7rooohpkHo9ZNW
vLe7Xyr4EqrBqBrHKNiONQ6Mbiay4qGvZLYzBTickFAAM++A0tEhSik2+2y0t7yV4jmB6uug4F/J
krcmX1ScL/iKtZl4ntrxR6L1TTqyxDmWB0iM1bG/CChC4MyOtR512tRzQ/C/ZvOVBUvFicdXWR3f
t4kjG/bKbFUD2mAX7mkHiWjK7ATZiEqc0dNeoOho51YA2cjo9qz5Bu8oBxHVPeGZe2t/wN5476Az
vajpKmccA9ddhxhxr4oVt1KnwCdR+95CIE5O0lozDbJbukrrW8p63doBP/ZgOowEUnsw5SKC3f4m
/gEmGrQacTEE7oSirPK/bKpYtQezFtEf+CyvgTIb9Zw2qhG+xMNRZUIyof+q616PBr0n33HBq8u4
LrmzFsq/mCjyoQP12HG65KucT7YUNsFqd9VLOPHT6J8O0D3g/CGl/CTg7ZhWYiMNWgmRidFBebu1
IB+htfLjpbXpg0NpTQUZVD6R2jbr00HyikWawiPP8DI32HVklY55uRiMrtj5mv0LgtlAp56z2x2I
WUK5JUBze4zltb+iJrgXST2X8UdAsVtYUabkoNlqfQH1s5lpETi7Qdfgvf7s27KB9wncctoCAPA4
Idnn8IWDXAVg7s5T9rAUWrNGQVb5FAdrSghmweXz9gBzROinfAYsAak0Tjw4gs242t/CQzD/4lp5
ljHAabxLe/fVcZ+qI1YwWsB44bkjf8GawVhzMuBrs2ypakoNNWzAcMKB8KnhQy3LJ8ahrJ4z8KMe
8RwSwbF7uSIpe0sau/AYDrnpMs9I1AzJYC7uMVXTc4jy8LKwv8G7/mqUgb6jPlAKiB+QXZKygUQ0
CVccWw2fhxYJJSAPNJ3gHaDCbl3ytP3I6PrMrgqli4DvhuSGPeWvuQxJ6u35THycDbdF5WuJN1RA
nsA3h4BrQqKGo5jLpV/SzhbPYAelZEZYwrC30FGh0XTfzpWxm1gyqG2Cn3DtjiqE6TjqhmjO049c
0aO1WMawPpEyIOSxb6pTJwKe/XVGCQnMpFZKqDIoKXiPFoSeXISn6nlmW8D4CEZliCqqZ9Gbt3Ca
Urhk0bS3/2GHNLd75t/BAn3Jnwa8Pcv/xwl8a4YD7n3V/11NWU5S9LZW8XE9Pi551TO+mmnPqZr5
R1i1a79iJbNsgeBp8y6Db7DgvujPgd+5y1yaiaD98MNaHMF3311XJW7Aj59Aez7Nf1VNvW53kHQm
GFkcsc9uBuDi00qQodCdMfMA8yyPBxnYt/NV4LwicGKyWfoXmDM60W/+h6w3FLKbJyT+xAB4X+1N
nKMFCvcnW3WUAzTNiUMbZP192uYsEn+uXpepbXZf9nQHqZ3kGA86BC27qPCMXg+l8iugJjUseOp0
hYFkKaMHt/uOT/xCA421jCaBciGaT5nhEHma9uGZQXjBoPt7WGR4XmjFr6oErt6wUljzaNQaGAto
v7oIhjFb9xRlJg==
`protect end_protected
