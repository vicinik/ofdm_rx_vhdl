��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`�����T;�x��Zg���)U�b����\C�]ȧ�n�ig���uWg����Gb��i>������o"V�SdsR����r�x�����5�%[x�
�e`J��:������D��%�֯qd�����D}`��н6a�_�	�ͯ�m�B�jpG�zy��b:�1v�cn��H���G�#T���n��-:��L�L�;Ha͆{���{~F���pJNG���&�P�>ҿ7�Hefv��po�ڐ1��R����J�䬝|�-�|���/���'O���l/��Tp�i��7Z��Zx-~�P\`J�{*c]��RȾ����%�T��I���՛�BK��W�1A� 	g�ڸ�ISGgEg�؀q��sn�A
��k[۲��4��r�wg<�K'�?[R���E���Pb�1��i(h�W}-C�F2�6��.�(�77�w9��&��(�8
-���Lk��;ފ�f�YaЫB&!��K�X�M~?���V�?T��7��Fv�W@l���*��F� �-d�����ɹBϏ�q$�����Xֳ~�v��������d�6ND�
���>�q�&*�w�5����C���(sW@l�T"�@�٘ᆹ��yb���'��%����rU����2��S��#!4{���&.��31�!��Fb�D������>/7d)��E�Ϻ��Q'�{�ӊ���.#�3��4M�-;Ψ ��f��q02/���r��������T������r���M��2g-��Do�k�lXVrA1c����Ξ����I���۷�md����z���we�zLcnW�%̂�`��1�=|���q;���V;hO3 G���u�mI�[��M�(l[����cV	�uZ���$zB�fP�NR0���
��;>Y�uU�4 ��]`� ��g�?dC��������Y_��Nl��v�����ה�ĵO�SR�[�i
��J�
��B��
�s�۾�����y��� ۴(.ez����K�V�p�T°$�CC2Ɔu�=m�6%�3`���e�
�^eW��+T#�ǝAQ~t[���
�������PL��2����V^�A�����'��|�e_�0~5�k j�F+�����������L����I���5Zs���䙺��ci�(G4���DQ9%o�$��7"i�RN)��=�36�F����j�Z�.Y��I`B��M�Ք�k�=��Oj��W���.����`=ٱ��ɒ��ɿr�����g����s!o����p�l�c��; �w�\f_�˴����} s:�E6�G&P�r�<@���\����TM���ｂ/q�2ع:��W�3�V��/l6c98�J���9L��d�F�2u4����6�U/�P� ���������k�R�ۘ�X���ot,�%غMsdf�~��B��Uϲ�im��&��V	t�h�gX�|�lV2�ՠ%�>*�Y��i,w���<a�w�����Z�_�j.��M�2JG�/�j���҃��?�����[�V9�#}gR�#E�B�A�r/~�����_̂����?cS�U`a^͕���kϜs\�P^�P��H-eo�+q�f^�΃����^뱷��S/�����La]Or6�Z<�%��L�D�'ݵQ���]�72/`:�g���W����ye�E�C$H�������;������q�8���=�B�]�p��L[���#�S�߹�>�;����mD���� �>U6��s�
%��
����D\<�S ���Lqm�1�͡�ON�K�'�1��E_�����.H�.��p�nx�gݵF �/X�f���K �8Z�N�NPʜ���&����l�C���z��/������b��QV2�x<�nEp�l]�T���Z������,�E�
�
� Ea��r�ݛ��ɏ�YX��2��tq���M�A�2���z�����k�G�1S�Z\oPN�"��iBQ&�T�_����Atی.���Gf��]u���:�;)A��8L�7 �n�z��/�g�]iZ�cF,�=0&��Z��~`�l�܅{�j����a�)zl����Z��n��wf�s�z�@�9-�|�y�i�;�Iy0ܹ�"�z��be����wࣳ ϖ�U�=�B�o9��8��Q1!I�
*Z,z��N[n	��:�Ĉ�8�NMJM�(� ɖ�bG ���t�­o.�Y�f):5�[C���n�.)�<��e�U�WJ��Z-s���1!Sd%���=\)h��S�vPf������e&���Q�ƌ�����	�o�@!���X�/��M��F:%��;`o��m��Y�x�b,�_�:����z<�\N�k�t3Y ���Aq��]�4p߆ѥ��T�EJrTk! `	�bD»)���.�>�x7��t�ϵ�\U�v��G�	��
)�������+q��u��r!���P{��mT�v{Tb��&���s��~����g'���z"�nx�d�JF�`&q��8��V$P��V��-���%��c���D��W���'C�[8���U�r����b>��4߉��
o\��g��˧"��j�Ix>S�x��l������ G��%����Pm
�K��f��ȵ�c+�+
d�@O�i��e����G׿a9�#��W��P�'�I� :�P�O�5�Ŀ6�CF]��^�v��&�j��W2W���o���sKf����NT�Ž��a񼨹�y*��@;ܤ5���H`)�����y�(y珪�c�i���#����qS�����ڞ-�2�����İ�Pg��6`/ҥ�B̟�i����3[�R|�*� �go���O�7bf$�\�;����� H����h�[_쉡ǐ(��fF�b�%������.�;�@���y9*�\��<��Q��#Ǩ�W��C>>D�N8�Չ�裬�3�c%�x�%��a(��\5S��H{��Fo)1�Jj�Ls���e���ȰK����P(�{���)��ŷ�iJP$sw+Mo-a?����/��y��gu���E�z_�?�ܨ�W.�{[nej�����<�Fp8c.�q�̱wԊu+��!���&qQ�
��-�tak��ݿ�,㟯����p��f�[u�1�9��BN+w��#�Ch��?I
��^,�Rp�]r|���]�Y��d�X��;�%o�4
F{��� D���yu	��lLa���룇{5�g��=�W,=�%��BXl��ho(ՆP��J|���������.4��ӯ���m��[�n�5��T2��{�����Ĕµ*q�� ^��*y���GL��XSå��"w�Ek��U��`�4��:�������3���v-,Y���Q�o���^�ʅ��r�ђ\D^ �4�'�w�"�g�ҟ9Ny�y_�9����7�L��W)W؃2�h�.�A�F���;��qJ�N$�`�Pb���#�E�A侖��������_��T��}��|#�3$p\���Pe���y��M/i�?�,΃|`r�ʒ@k����A���
w�?*�N�9�.�lu�R&Ã�m;�}>���2A�Sp�	���jgDUps`_N]LN� �zy��Q���3��m�,j8A-*��t��{6�?V|����9C�P~s�)w}i��t��#��&0}� ��ӂ�a�c	9�3��<ܓ�s�2���OE��t��@�#��@�Ts�jA���;�H�`\���k��g`n�Ήǹp֮S��.3�8:�R�߄��N�]��K��Mi�ݓL�D��'��Q���v��Q�����!��Y��K��ֹ��ֽ{y�d�(��Y�wlړ��
4a����}�N&yG�',b����m���bZq��1�'i`��ﯘ��sKw6�{bHX�O,|����ε��ݶ��\	�o$�>�|ז�c��c�t��q�a.��/��p��j�
�_q4ݣ}3�,�[/����^��4�a؇y^�����,��b��Ν4��Dn�gד��x�7X?ac>�b���hN����*� �AT��F t�������^����	'�S֡x��ʦB�M����a^�#��<�x6 N���L���#N�ԟfGCK6��/R1��@%^t��ك�T$`�� ��b�L74Ńaj���o���`
ڔࢼq��<��������x���3Si�Dx}�Q���liW���c���"-ۦH9���ů4J�z7���oO��lxڒ�u��F	�Ԫ��QՕ�^�JY�z]����_z�:|����N\�kf�(]`�U�5��Iqٲ��4���o,�tx�~�F<2��� ����E�T�W��|��՗�6�Ղ���IX�n4:<�1�;�����E`_��rϼ��Ԗ^��[��0FAĐCs�2�D�Ԫb���4���|��+��g���	�׵6�,u@�Єpc�*��伳���U���2�Wm��'zю<(�[Ip?��[���vC5��AC]G /xJ�������W�>�W�bo�2����[<>��2��jG�'s��y]�vh�PknEp�hԎ�w�@�x��ܡLf޷aU���П�݈���+NUl��
?��%�6(������y7��>@�7v_��T ��d���(�YG\캋��4d��fۤ���`�,4��R:��s�;=��v�.Tg�zd�ϳ2���)n�)i��}��^<-r�m5��(��u3��&���dJ�D�z$�����$׺�+ph�G�.dٌ�y��V�r���X�f*���n��=&�m���|�FR
�=�Z�EF���֨��\��7#�ɪ���5?��ٳp1�M����͗����"o^?l��;��{�u��G)K�3���#�S�ǈ����DY��g���1�:�Wa�s1�)_~���M�gk�7L�ڐ��d�,g��,�cޔx�#�:�P�4���MA2_�[ϱ����T��9�^0gB� G%�a��c�c/s0Q�u�r���-A���ox�ϺX�&�]%�c��{jR�;2*I��MX�B�����<��kR�u�����  ��tp0]�����/���j�\���+�y3�փ�Е�<�=����J;\��29�A� ������5�_�*���5�e��3��W.U=j����G9�f��u�Y*}W�&	�~��;]��cFg��	�KIh��[�t�g�oٰ�'�B�zXU]�⫴w��`S��&f��־�vG 26��T�n�?(A�7�S���N�xla1�ȏ����\��C�� �[R���0�f
#���C���Ty/v ʭH#E?�hɀ��V�&���A�LJe���X�--�jh�z��B%�6�h�����)�+��i��g�4�޿mX�@s��6����9� ���́A����S�j\mι�Ә#��<�F/�1Pw����Y���$���ӯ��HˉS
7��yVS�>�ahђ�����i>���5�nrurjn�[|�#��:��x?b-�!����9��;�U�N����Ԝjp� �tFB������RZ��_W�)�a[e��VwĞT�b�4dD���U�H�=��|�����q���z-'�2;.��Cq����J�-�8��)�IdG���؞���F��֢�U������o�]k|�,�?��]�U��U1��H��X|���ǵ�<�U��)���,y9|W	���vnXtn�փU�:Z�>G�D�(�S���>/�*En �P��+�<a.��Go[���r��5c�������=��z�"��5pX�n�� 	:���v�<~V^����u�!�s�f<�KgD����z��Ʃ����/n��òX�# h�IR�5n܇8��^B� �y��mU��[2��������%np�gny��FZ/�b�
����#Ӓ�=<��m�i��W�A�+���2t=������Me����q����.E8�
��J�U1��_c�z�J�wa���z�z��g���
�>�

V@q�kx�
G���ݥ���4Xu=kc�f "��O�r ;PiT�T4���ꚤ>�y�q�L��_�S@G0�y�T��Z��H�l���6 vZ�l�����k���g��ѡ��ɡy�
|�>��!���p}�3���I�@<�C5���ӎ�dd渿z�q_�_)�h4�oKk���=@-��G�{�Ńk��5��h�HF�G�Y�&أm��Ǿ�<�}l�7'tIV-���<IV^Q�e��ϩ�O����A�� ��:��|G����d'h�Usn�Sl�b���H��ulC)�G|�k��W�JEЁZ���Bu5V0��;@;g���e��x�#ǘY���V뇟��?i6�	�ЦR�[����:_�J���oX38
�CÐ���p�H���!G���=���u��6��9ð��ism홚gؼ�}�u���k���T���f��.�X�2���$���2���P
�}���~�_�� [Y�x�I|�D�.ڣ���lUԂ�qMsA��Xa/�$�qD��;��b�1 HC8�6���]�:`N� �6v t�t��7,u���]�������C@c�T=Q�t���=0���O�a�bO��AYBF 4`T~ h��=Qu� �.����~�?���I�@U&,��}�vΈ�T�$�w"���2ز�c�g�*ޔ���aMF��>kuJ��_Ny5&������ġ�t*=��)NVT���Wҧ}�L�;�{3.�d�gɗ�c"�M�������l(^_=(&]���e���[�D���ǿ{��H;�(�M[�Ѱ>��������T� d�=o�j;~B�T�Z�~�\�cYc�dt7�l��|��:�~��W8^2��פ�3ZسCrQZb� ���tV��FTp��?ח�E�N5R-��*���N�w[����Љ��k�<���X� �C��/�*N������?�f0;��ۻ4���pz��c�-
���zb7��ye��i�%�ߥD�N�j�,qgyKfl��h�ݧ��!���*i�>�C*�Y�B�{�f�co��T�y��C����t���L�ְ��^ʕũ2F�����]�"��[��r���/��*��ZEM�h��Y�@"0�1�o6��_���u\I�WS��#�K�8��$͑�cp[=���W�W�O� �a�AR&��޶�����!�l:���
į�'|_���k�5Ap�6:����뚵4v"$��zD��k�})�!G�+�VQ��ye)6�����<��J�f£ɰ�v����t�-��6��vc0[�s���쾆��O�y��p���9�G�����q��+ 4ك(����Ғ���M�[�K��\\Y�vf�{FۼFȝ�w��c��((O�Mp �H�[�@�� @�~ڈy�ƛ�픒\xw)ϙ-�7@���e��>jؤ�z҈?�|�t��"I(R�oYMI�J�l��j�v�+�p��Ĉ�Ǘ�u\�Y�c��')�<s;�򟷳�j��&��N<�8�G�������"g��p�1F�73�]�%�+����?C��Pw픟�򼓢3d�IW'�\r��]�ɫ!�o<�tP��4�^��̅Ӗ���b^����6�C,Q�9��O#����=9��F��0��|z�ˀ�St��a3�x���D���PQ\{�����^�9�k��[��b_�N�@t��a�Tt�1��g�"�R8��TK�\+!����/1�K0�it-�Ε���6�>�M,̙ۥ���QJ�^�L2gc�b,��<�ֶ��N�hB���Wo<��s.\�(��@B��@ M���
Y@��ޱ� �-��%Q?$�����,5��<*���t�PR��{qx�	��� �#�<��<0 !�UU�ԁ,���H-h"�)*Ny576�`�rv��-ٶ�^Q�}BQ������Vɘ�����r&~)�&"�0PW]M�Jl�n_jZ���#W�z[�e1�7�q�Ʊ�.лb�x�V%�T��ް@Y�d����`!c
 �|��Vs������ D�S)cb�;5���ˈi?)�e�etgpu�x��J񽃴��C��T�
L� � �!��tΥ|�ʚz���3�KB���𪠾���y�
oz���yފ�r=SLNUe��,僜�!p~��VMJ,�*�u��*+?I/R��� 6N���ǳ�/.�=�б�jT7��޽'��*��S8��u:�����C�g�_�������w�eĮ�oo�!q!"<uhʰ�
�������1+�>*8�i��M7���sd�S�����f@�9x��g��Fc�?���HD�j���Y6G����V�o���Sf|[u����U���#��@�kF�߄�e2�a��&7i�/J�9/CN����!��	'�l���KwR�ne6�d|�4��T�;��{���cp��-<��}xT��Z8��^ ����Xvu��w�Nr�����ҁ�Qu@�T�����y���񳰁�#�	QMr���]ȫ�)͓@sIUa��۴"D[U�_��r��ICX�i6��s3y{޺�ob�s��B�u��������1Z��1����I6(d⤷5�}g�bQ|I�<�L4�mD���
,��>�}Cn��@,_�'(G�ݿd��#6� DY��5��v�C�	��p@вD�E�(�����g��+����Z�d���򢻐��g��������97/>��R�rF��LyWgL��뽼�خI5t�{F��1�hf#�ܛ��C��:XP�[��Gd�8��m�T�K�+����x|�
|�b<vg���I�������zrN�[Ű������SĶ������kS�������I*�ѽ����)���}\�}mR�Zv�ai���AS���`�(5� y�����kl�G��0��H7f{E��S�5���	�r���7����Qm�I��D���2�)��wS�]�/(�����e�����Ko� �� ��{�°�W�8ڴ�d���cr2���)��"W3(���8Cz?��������r�eb��	�	e��[<�F'��H��<U+���+����w�ף�?	���[8�;��5�_��Wj��[���ɟ�Zj\$�Qx�^(�1ε�齗l[�_�Z����9jG�G��+q'�9��	�>��������1�F����b�=!�|jL�z���t����oэ	YSrq#���S��{.!/g�n��N�M���
�����Y{����z�ƞ�x�s�(i=h/C�?
�Ű�컳���_T���?��kLt�%b���h���3�����\��i'������7��7j�lp/>��ā�#��x����C���::�[���oG��M�K!��xT�=@�ڵ�jY�Y�_�b�r�j\{��j���ȟv`�nIN��HI�gFM��g$�$,���ο�'E���r��,¶��z��Tq��q��������(�o%Ǒt�r��H���q |�%(��������A)���6�6���Ru?��AӒ"(���Qh¤����׫v	5���QyG.���@e~(Jq�Z��C��%�ǖ���`$�	�|s1h��R��#[=�����a/��ݘ"�K���4n�� �6�������	�.�*�
��`F!�����oOw�zo�;��A
�=�07�=֥��
�nl�A��@DGo7@fu��z�?ϑ6�/��m��g�������d�SP������3A�Y�_��ę6��K��R�/]��,I����F%g����T��x%��x�_{d�s�X߰�T"��07���8:�t�ŋ�Qm�C�@�\�%i�@YNڎ>�(:F�yj�޹���*Gk�?d䊮#�����������"�u�B����Z����TmOi-G]ƙi��8����x��!�X�S3�L~2� �M'~Qv�d���%#AI��ޤf�r�S�*��!pʡ�6H�
�{�q�bW��������Hb��t�4����(���íC����sq�l);�_�&pP��.�ױxu��%��H=�y��#*K����J�� ����F障"�iY.X5�詞��Q
w�h-�2�JE��t�gh���g���������3��L�1[U�!)�{�h�,����o|P���#���O���4�j�����o����g�K.��� ��D�4���A6�n�Pү[#�M��G[M�c�a�9�cVg�f)�%�!:L��j{8QO�D�]�-�2�S/t���:3��#�Q~��0GQ�GI��$6b�c���J��'���ɷW��6Ѷ�L�Z���6Ǿ�5��"C4D;�C�(Ê�w���3�1�s[B��������Dtnc�Tx������Z.@$Ȥ�n(ﮰO��mv�/r�@�ɽ'�G�]����#�0{-[�#'��\+x�����t�f��!b�x����~$��ę��%���3FM���k���M�p��.J$ig؎�o.Ï����I�]5����яi�%��-d�a{���^��Ȗas5�Ԟ��+�����o�������a�5!@�v�^�-K���Rt���x���waϒ�b�=8�	*s�"¢��'��=�/Y%fqjr(�*�o��J��d����H���{�`	�|q�7}�̠��G��4i,��Wf[��|$��G=�ܺ��Gj���d��	��}1��UYd컧6#���~���"L�l�>:b�,�1�wf��j�(��kz�DE�h��N^-.�  �#������ r�`��R4-O����������P�TY	�C0�3x?ν��%5��f�''��ܹ��O}u���m���N �x...xU�S��#���@�W��z�I�$�hK��s�Jb�K�e��9�,��Zk��K�1Š�)�p�BŰ���)�MH/޽�1TB�G{
��/�&��ֆ̀�,#������n��>�u%uɌ���U�.��i��Tx�a]��}�j�{gJ�����PR�t�N�	���.6T�a��/��I���_Ҡ� �����p�_8F�.�h����gptt۷�c��f��|U�ΐrŶ�&��tС�����N� �#A���1���@����s�M�8So��S�$cw�.Q3���L�w�B���&�x�~7Ȣ-Vd�{M_8$z+t&2��	;�y��@���>�r�i@��ڦw���8Đ�k�Ŋx�N����J^�!����_QN�{a�
�ꎂ�n	p���%��� �!��g��1��x/
��@<Y*)�:q�u_��bt�Y RĽ A��K�6�	���jٵa�vJB��w�5�*��p4�w�2$�jg~��k�?��|�[u��d��Z�� Ȳ8�'g�'��/m��7��硣g�Ws�vo�o��1h��+�An3�G�����01�=�lK��q�D	��`9ò�C���W;�@_ێ@�h��Mh-wj�yA�aRiP���m*cd�53"�tm��p�w۱9��y��n)�W�v<����@�$}��YT��F$gπ�9���R��%kd��Hp��M��3D��
���<p��"��}T��h��A�C�o�/��?��ܤ�S�
.�h�ob�G׵M.�p�z
T,ƾ��XV�k)��8$���ڳ��%�p��TS*'S��(�&�_�$�?1t�B���?���W�ˆxX�R~eF$ي�/�$9N�v&�+E������Ui����w����ab*;v�����.�[R���\��������J����z�5���Z���m�b�v	�)�-�<�i�_C��ܧ�XOJ��,o�~���ٍ����U����9�|>`������-�s�
qv9�.L�ytl��X$e9Y��oEl"'� ������B2;����땄��e4DOg��V�_��w:?HC��� A