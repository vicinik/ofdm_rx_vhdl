-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
W/jm/kggAOEeHTPTCRS/+aJI2CU12AQEn5mXsJhF1BAgI8uNW/R6IDio7GSZrVtoKsmLFtjoSfmV
doqRXM+6ox17879WQtQEQqp7cr4040jXdGctCuim0LhKXHEoU6dbLFtKnV92isSP9gAqtm9O0EM3
s4gUqZJxHeQlHaIGuwmi7Xo/iAVF4PzLvgWKQEsTq8gcpaRjz4gbtUHlzymobMok8/NaDZEYPvM0
UepP3GEV+L7dlQu8/Py2QUQdbggQAbhQKpAy9DUcq9Qi8fZ1zlsJnb1b3F1WCwWhxn6zpEvb8rK6
EwRXEAuFRZWXvc+Q3EDy2PNZleqtzffjLuu7xg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47136)
`protect data_block
3JTtDuIm/l2gFlP8VUlCcRXJWirNL3zOGOkjyhEjeSyzqmtaTphT67/EbNNe9eAlYtpUTxR3tz6p
oOvxafuX9i/rKfjz33jDl8ojhNUm5oGcWmHdklslF3b1C2v1wxt4uwzd8ZBJb7VWPrDxDGyPjPYZ
XD8RCEA3T2uHGWYLg/HH1X1rmzVX37zF8qy6jyomyRbWil23QL7mciHIXuMRfEjJCE1Qy23fu9wU
mvsxDZs8fmgpEhPUFRYcm4HmSHVr++QZkQLtYVgsVmPqD4zp48rx07knlZqAgcIBQSPDrdh/yVYu
N+ocyTMFQ2UNUBatkXiQQHTnt/Nx5lUIBIEo3zsHykSrBdJAd4l9dk58ZbHddkWLz3y6xnUw+0Rm
L18dou/rknJOpNN65DhV8DVy+aRUuL35GGE7hoCbKPdfN8yVffmdK42bCTFsv0JnrvmPbfFC0Itw
G/ZtNoVmwk9KW1lFks0lIK53lEkFqkCVDYzzON81oW+9/ErWoHpQclFIAmPNu+GciZunlFqJZ+Yl
a1mRbFhJstv6NcsShoVIsDKJscE+4VXZ8DbQBQZI7QW6xqA6YrStryAwTIVCL+fb39P3GkkOZaNd
yc7lcc8wMCO9zbdJ1QgXQrpxuwJi2csoZW+F+icFBb9SdFD8YuCnRFHIJ3xWUdOji8uYJLBLaOs8
ZTeTdsHvleDZpntpdptfuKKFfWKizomoy/81D1xoAkfUl+M6hzpHr+OmuQ8MDu30w79L73JKdzcJ
8zObnvx7Ilg7nUG65PvTzRIkhg+XO4DXC17+hPugDmuWwTaBcFNA+jkvfZPce7EuGm/D9Xp9Mr+O
auYfJorPHKbWM27ix3Xtmwr8T/M+IBGWxag32gK90Kk2JdYtfj9Q4JTA52KzKqLh1C2a7XR2hVAQ
8VuP8BQUuf+QnnBAfP+6H2WwzwpqfWa37hUcp4AgxsCc7ReEq6YbCtzCuC0skLEoBJu9R+c/Q6+U
RxZ68su5I9X4BY8K6vNgN4e2v4WOU3wWWq7/2oSxs9/LwnS0Usg89YjRf53KVVZQDMCpq1Rhveba
Hj+XwZomqKoZxKGcu45NoR2rlbF/Bce/XaiUethtj5wQPfkJuVM4zEausPdInfgLDc473zV7CumA
jligoDZzaUUX9Zeyr9FawjCSlzmYAtmh9uNj35gwVYHELfs1O3jSuyTkQKWXWtzzYRiSqM2C2DkT
y7HJOBq4LX0vbRLjVAlYBejszJGmRzagltfr9JSMuQPzamPRLce9vNs9LIETIxiBrjX042MJPONh
N2VajBXt4EM96Qy4bnYHJXU0lAFLzjZbLsMude21+KyhiC4BBDrnCBROcvZe1GI2z7xT1g3QAwQd
hqnfpU6qnhw+DOuaJX75fVRivP9mjTXE2gbnLHPvVz5yAh+XRkNKj3dOciNQDk/iFe4CpIwKyhRl
zcCO1EIMuVoptzpBrbLovBx/BHN1ClDu2Baed7f/6gFtQDyXQUvvyu8JT0M1CprYe2VVBcRpCvuX
hxZjC8B+ZX2EKNDwv7YMcremze31rWXeRtoMjaLthyot0m342fwskzvRjm4WdZifdVl+ES3AZr37
Nt34chcxIwR+xR83lwNmu7STMxCrObKVYBBF/gfYGni7ObOGLs3lMfzEDkGfYAk9z0NUNbmikV3L
caRI30g0s0krz683JwB85ZYwUH+m0UmN00xQgl/HdwYeMw1VF//ZZB8fPrpfodLNESS8GUIv1v+l
mS4GPLcnpOReAVeqfpj6TlR3VP7pf5DMBFQhsB/GryKeRxmF9zawoHSptkC12dv0rNcGe3Dn8IYc
wOHN2svTE1XduZeAboo4+o9i52FT+TSmkGsW6tm+lKmNVuE5cNqg5RRryuYee4XTPCsMH2QlkFyd
ZJ5Rc8EC3d5tRwf6AU02FdWgKmWJLIV7g7O+7F2Ti5YZVEwBjwPrdin9iejheJTMxSaRC35Z+Okp
Ig4whnqBvFHWh6JS5VQOmOt2DMe+z/5BFYoyzIrtJpFYYionb7qLDHq2xW4Bn3ZNv+yJftilrGXE
Qy/h/pLT5G2ragxKxtt0cG7zWPtsIJVqlWmJRzmiy3B7v3Nz8USNcxIcVQEmzYfC3+NaQWcofQ6f
4C+bRYnOu1ard8ALylsR94XfXmDJRKo7lJFj3v+mMHon37/B1L+1ZmO6sacwGEcMA3I+uGNuzlbU
Vhzwf7uuRBEn7NRsCVA6oVfg2tjGzC3QKStEr5mxhgbylGTDFJX7GH0i6iF2m56ulY0c76RWwncw
0/KzOdn01WW2jtPC1CmIAdqZqrZD4CDViggKi6tjerGpisL/WaLVPfuk0/hg2tIXYL3iB/gz/ENz
DG2YRZHhMxm0131GnzpPb6SF1EM2Adg8JDiNDfTkWjX416jbM23J7sfZkKRfDJwwjWF3HQjfx0f+
UB3pPn8JRK4zQwHcl6HeWY3u6cBBzSsuzfrCu3/nl2+5prPqOlGnNe0PxdJSQpG0TmazS9YBXTS2
Fz149R6c+qdrgK+tZZnA8oda06eJSpoH6Rt3qyjfmXBULwyGWILdxLSYqYOmQ/hT+Zbsm3Pw8CTk
XlE957GOipCtP8XvviN0ElOd9bPDBMGzoA+lX+7URbuKSf3mJe7XmaxVN7LSo2XjllfCtjQDwy4T
bCLiJtrCywH4eBJbzZhm6aOUnkKb9yKgwWkJBWtu7N8sJT3ryK+2GOz8RGiS26IDOTFebA0Ps3wE
FPnP5rk29rA8WEe5RUUGeGcEocMOnsQI6GjQ9zuXbufnkNjtYsMGJMjdd45bA8btKC3vewNQ/pW7
GYrg2Tsd01m/ns5nn690IcBzd1Zy1euCa4FK3x6J8OYTldcIvtts6iQN4gEFdwG5pMP51p92tKb1
AGoD0mc/GvAaDc6wxPlIGKvvkO+pQaSeIuPrHyNxGYBk6gKOh/nO5J6MlFwzCOwjrLWdVWrDTPON
PqCP6/dZdNqiVmQ05dACSAMiOxwfemDOTwjtjZrnypFTv5h7mK97DxC21RIhhvOrzUPnhUySvlFf
OUxWearopxmV+PhSf2yu6SvJEZcKwipEat4PQpnp2td5Zo2xxQE+SpHF5vI82T7CuOdKgUJlY1xS
ZiPTMmBLMaBqLk2C6wEsp8WxglOk1EcaPeR7VbXyEbQSwkUzyNXqn6J9B/t4kRZLC7xHUZkrm2N1
/vbJ/zYme/NIZRDxBwS5we1iOpfwr7KfeXZYEYJp3HtFhVvW5dh/i9kzyOPo6tBLRsLGv/BgTp23
fWu6S0MQso9vymdwppyZztjxlrUbFP384xKsUQApM1clI870QeGqmQErSI0j2tnqPgtIuUg1/jwI
NkgVHSLOdkxQase8QA+RvK0FZB1XXd4xoZhZNqHXJu5c/3ezof3eoDDCaS9QcfDxNnNTj4qRcP8c
OhIq0+6UAStvl2dMgBwfuqUyFSxcskGeykdvN6mskX50Ohmh41jfRJO/PDD3qhGUtpTfsP5crx3r
s9azgTjB5PvPRg57LKrbPDve955nlmmL+xYSeLjttijTseS1XarnqcyLPNyge+PLhESz+7V4cbE+
EzfbOw2F4ytpFbRnuGmCh9hLhMy3k2qu6a95AN7kEE1D1vZBi5z4xTBkF+CvWIWjFHtr+LfN+xDV
mPTwMBoebuBa7E89wSSmlkNPprIsX4mLs9512qAEvELDqnzqWJN0XE7ryTAVxkFQvoM8spPb6XeA
XAPYUNCh99gy7dWOBGEocwx6ZSHQWjMBx3gS1DfxAZiaArE/XGJIXwfPWNGMRzCWf/br95FIjpRl
CEk6uz4LRzss6ZVezInJlRRxjAWuOHhkb4++JSVRq1jNZWVJFk0OReO4Yr/H0jh6WkfVJ60T4FBC
Q4Mh6nSYgP6tujl0hDCePTI1dm7Qg1eWD1M8i+r/gBaOYAcg97s3IKoV6UyYkhYqQQYKzm/VvmNQ
iSKMoXwe+4z+mG33Jm4wu1ye8+aL2qQQoX2nsA8toP7f4BCDaoWn0Jk9mp5CQhXHtIqcbB8RpYH7
mkP91cgU6ZX1+NiwqTS8JxGtynT2jqC42tM9uX8Jknd+1OnfZt8DvjCSjxxweSX56dHnx0dd+feG
bfA89IqM1mPA84bEfWJtR4buZPvOwUS1UtU7+M+aIRSB4vLpCkGCKGxvF3vRbF/X+GvW+1QS/i4y
NtpMv2KasavvalHc+46lkGLt6pm7UOaCvSGVKvYGXzbLzsO1m6DKZICTWG6TDprXwSCp7Y/oYAGj
vAE0MxIi/B9i+IA01pZtylcBBK7jNvdAij3BrFeo7MDNtYD0rVPyHujNV++s5T/66QhgXufWxdRf
hDdZ4tePGahFxwjywYoitK179wMH91o6yI2sMZW+pMag9Ilo/5JY3OB0TaGkKXpuxsI7YwDMWa0a
t2l1RSJ2Y4QGkX68QWLDocDfx+xVS61fAyoenkTtGx3GUW2JmZBjEMWH9k99uDEfTIF3gFK+0CNk
1XCUApS1n/O6EGaPx/r5qol1KrBSf8JAbLNAsH0/w4J7jF8EuzOG8oF0/LdtNKvYvnLSYIibHOmp
agpGmw/l/WcQNWS0bKoe1DEs0vtEY/VgaDIO25YGEHOx0POdz4wUA02mRghtRqmfpYS5z2F76m55
6w1iRlLlO+feEU+kpWQNC8QDGwhDMyirt+XjiVQ+cpMzGAWjw1yhHw7NJhbGftoXA3s6GPkU/Ehd
p1DOUsmji03lgzofj2LrFI/XcyflO9xztx3iCTE9XwNxs0oTe4Lu0OvYZxocpNLT4KTTs/84wA42
EJcpIZOGIRmvQmFBx5QnLtsh6niGnCJXcgGEMu3E8+sJAsig1DHwbbDKFa+2XJsbgTlJZv6ocEsb
eBn0sUjFLgYgnhtuG8seWXmJtFdDLdwN5TX76ePHdedS3sRu0JdwnVRjQCuc73hiw2EgZ2dtWVhH
X6M5yryjfFMg4a77Bgsu4DWQCingIM0r+mw0IMPUGLsFwaZHZd2KFIvxQvBN3bj+z/l+kvvNq+kQ
wyttrsPhQptpripYtr3CARYve55umSbhEaQnWnKym7YxSst+C9d624mrANflDid3kW80DrpVNid5
HKYHIncCo8cGa7E9HeMB29EIkqiAsvX2RJfJRPJl+0RJyVaNFZEg+1c7SPsv7Ld1AQ+Bwb8tRwgI
bwh+3pDx3L9vPbX2XnzUCSEBYl21KKZoxqrSOLJpqNKTj1x7q524OsaZu2gwPIAjMKp62RQTUAUx
8G8u03C+Ww06xhCUr+z5GlbAJlutf3/kQ1PEBRyWSH6IFAmgNNV2Kv3JnS1Z9VaNR4HeObXHORH5
01mxccC3psEvca+CdxvvJHlpKy9ia8754MOv+r7ZPz8XyKk5NAzmi0MA79BYYQLfHgaSznI161xD
MzNFeJWmQATudREPc8L9eOyVeqPhe/ge0nH3p86fc5h0uQyX0S/WyyBSPJ0VS4XPDTSRLMx9G1YT
NSpmDJTd6eyc9Uhau7ixakNpJ5xiMyExYlMzNEXCLrqbFez5sSpEYyJOq0q1RIzdMQlLimIEDJ9S
avQPtNWa+HQcLqCMC40Jc2BxTKlUnZHtjP5LARWkL/jvDRbFdqPNZtR/thRwaBrgtM0lfXmrO/7M
jseFmID2Q/tY8ZlRIqc4usj54uJPfvAkUDTTOlQiCmcG/9P2/HpwZ6k+bsh4Hde7xQIxb+UPSPU0
mCjSUBqgxr3Pz9fTOfKuc2rAjDKAff8sIsdLGlUAzUwj9w8sffiSafOoed3kpAHxQXejactEDB76
uI+Qaxbm89Gpk/zmN8t5HQXpd4Z5KHwCaBY2UlR0u9HLFZXDoPiCp9dUI8EXDl9vUbV6HBsCUX6/
7pKFrHzEQRjmzeOrUoetY4CQbFMSwN5RhM9kfsrs91co5vUQ5/nPYnSyi6WfmSJsAWfEDNtlKy3k
xfP0SOPql1kFTcOeRqDL/b8g8z8sdeCp0C8ZCZI0oAl0oCcCRWn/kBa2+STSOLiMPQX1sZnw/qnG
UnbNL6h1WlzVX/onpezXB/3bYbaBvhlMqAK1Jw/3LtBfA8XY6NiUkO/gZafvvYEkyECWoBIKsU7l
mq8kya355hK9i2LgDQ0KvJReju0bse/s3iPKlUJ677DzBjVEb72HWi/4FQmdBgkgz3htUZDknMhW
/ICuQAVo0BHBWBp9T2gd0+AzNnjkt1qP5yzxiAlr8c8Ioo6o0LM9DeiKX3rJiqCon6G3Buyxg3zK
tFtXepqaEVhDhC6lb+Eboj8FbYDfS8/69JeL3KHP7PHAmHuRwrYP05BxuLnP2stR8zg0hqln8mwp
Vq1cPVm3zQUFlc2HPYSOdDxgJlfqIgAX8yh3pmLJyoJuDSafqhgVEDpnITwCkvvYdig6R3AlriUc
yZ2lfpZTXO4ek7ZPt/zoBxNdDkOFu1DxrvSKqN9HQi6ZM95gY3CfdzEzO8Mgst4hlIVJEM3vqqVU
w5TStTlgyPN4nddoKS6TJZjgCsm7bdtk5eleUpxOdp5zvKOq+0Fsxx0xGinXjq72vswS6h/x/8gU
AjlHyGbtEp9YG877t28SkioRIEwIrnBtBI5eAwkMsKPhKrbIbVSwF6h85OE+//N0AqYgE+j/KcFF
h+HM+7LclZ+Ct9zWwmMrBgfYoK8jV+X6pQ78inEAJEePWAhFqS8ndB12ksnnGp9d0djaZ4svI7iA
gMPevyb2BRUHj+4i1kHyDoUjiKe7XKxE5rSqIXEMFSNvvT+avTG4UG4MBb1esj9qkvlDwcYbTXUQ
e7lDDjCIxWavHqKU79kHwE02ddAq7VrZugGHtJM2K1Z/Es0yjwXjBC9kaKP/PxH6LW7fpLD5SnxZ
OrNMQjKCEmJYx0i9hvNcHk9xQx4ZbZaTdEsYQr4II4yQWyCZOJ2XUPkZdYGSgrP5VQlk4WC0+J27
gJaYWibwJOX3uLes3GVlZwZdG3p4OOlaJbwWzI7oaQj25uNVaouOON8B+Lntm8/wlwyczF6EavtD
0ZSnKNSo62oQdC4ZGdP+0qUxcYU1PWrTTc+AycuOz7piGTVzD93KfoKXhIi1YdfnFvI57S+kheal
oSa7l5YEiEWBhjyvyBlYCe2dsgPDiS7nHw0kAdUN/GBpEB5kMnaHSeS6vIWUhfBHHy0e2iSHs4Pi
VF1S8QrQ0SoV+S3eRU3quV0AIYuu5FHmjbqM9bmecY9L/719Yk7MUNWHWw70Et1Qs2cEoedZ83y2
RYFPDMlNElNy8IYiM13rVYUcBEs2Y3gP7e0HGA3i042K4V/AMWWAYWHs5Tmm9iiTSS/5sGc8cEez
h6N7Aq8qf75y1oS1jSFMRz3iJp4K1AMErpNcnn4T5jguewwbP+oooiM2wMjvcrHt77znfdsjPNaZ
8u3NUpOplx3c4sW50qBKWJHP0Uf5egUVydGf6BRoLp8cEu/XJoz8IFNYET30fTvy+7PlXGvwe6JH
r+immT4LNc/8IN+D2eiIarPzCqsN0qKD3ZziMLAXs6jpg+OuS6rvrYgnWHmi6pepz13PS0+BQXey
IMFo4yMYrSyglzToUciapsd+zayijmUDWeV3GRQAOg5kRAReWse3EA3/nyLAAqC+5ucW198Sp8m/
1DYGXaY3EfM0WJuExxpuCuXossreQs0C1+9gDsQqBa34IepiMITqxLpz+C0KcXb0bvB2bpwdBted
hjQ3kqJwf5HjXV/mCaHDco3Q1TJTl3q712hOMnVHBb6Kz3pcbNLLRGfwFVevef2El97nRmN+PiKr
cYdhTgrR3KagAWGz9kxo30RZ7cil7Zv7OyOBKv2ioMzOStzCLWQ0OHIWkn1qUeQMmqsDubypCh8k
i/U57C+Cka6VIERKmnWvmchQ6zu6b1io4Dn19PC27fUijA7BFGIzzKQuJSRw5wGgAVjnSKnOAxl5
1VUyLeD18UoLqc0Hw/WxZvjAD0yJvBzkiAIz3goUC7SeEYHQe+cYt8OvC8/Fixa/ffD1fUpzuLs2
mKWCS8GOVhjXPk1xgYUk756gEKUy1AQA+L2HwWCDYEgRiqqI+Jd+bTgHOLl3c3Zx4+7ywOH0MgJc
lHz+mk7UemM3LXpRmmM1/eEFGp2A+7KcrnJ7Ts5tPBatV7JA5mHAgHE8XkVWseUMn2MrKvEGNt7I
RRTEKOoIGdvGJICgGZ8DxeoE56WnZ2CgJ4QY9kKvxGoP8ZnhxB8hKyGRyryos8WAEifDJbD7cNJn
zqMbTS1alas2pSV8t2eScfiMMzY8sAlwMlg+1rS4GiPVAhne24A+wc/ANtBvopPr7MmiPZUnB8H9
WxPZz/auIj9tgXp4GF16MQOwyjsULk5rSVqWRcittzkL9tlvPhjdm0qthRvubsdqORBxtVCzjE+G
taed1Rs1LJkegNeN1dTWNG/elMWTnabeTqP89tAXWhyFAvTZ+4vABKCSjf3FM+sDQb3hYZF4GN3J
w9eJqqfJWgj/wPtZpq6Bg2zgXerytL+Iyzqp0MHKtwvDXi7fwA/sp4TiF6zHQzKCPkb1aFtFFUpe
K5nwJexdvRea9IFRxjIGf0rDHlQZX+EDua4pDzAi1EVt+qIphsz4JB7YcWxQiayQILPBnMXKKoYD
zvSy/PeJ9S/W+l/LmiG2LTquxAfGz7Ti9Mf1E7N06+OkYwseh3ArD7LBZuOu7RKx+gMz6BnWTVZ6
nSXpycyZ6gU8it4J7htoVZNnsxngHf9akvQHBAjG9tf2C4dr5Uzyl/VWOOxbcw/wxWGT5za45kBe
71/42dlOK70rKwSUC65DjTqkMnGW1UcrXxXofct/B+XviJh8avy/rt6je7d4mdksVFm0Gs0+WUS/
PUqvZHILkSeeT5FkU8pY2r75eb3+luQtr/Pgd6fgvt3B44sHY8EaC4iepNclLPAxMcU1Top15AM/
PooSQBNBBuTxkhG4uN/s2qtF55HRU86q6QfecAWuS4j1IOnl8q2kc1rQ2GGkqoki/O40ZHkzzS+f
mdDnQc3GWeDuQPGdD9AmjpTsBIRc0cTMTvssLeB6T8J3Y7U4nACahOIqfxiFRDpAXmOh8dD26nHJ
ksF0YRpc03Md395+BKj5v3U69ShgWWYa2np+/hGx3EA9qM971O/Hm8IH6vBpbsqhKQX5IfDrHc2T
W3JQcj8KHfhbEWOYuhpux2nDh2Bt0NO98Z3+hEeMcek5lN3d/yLfPyCNmzSyNXl80y6JZEEd1gnl
37dAZxio6BUglDNliXySAgCFH7rEIS6xAVEgecc3OWhkq0NsPoLhfKVQkk/wGiH1qsHVXQRVW2fI
4ZwUPoYF/7jfhSHF2jkNARjzNXsLKnIPWn987kc1rT1zKjgwZ1nml2yiotJ2pr6gF3zgOh2Wkk4W
4oS4XcOVLHxbnSLQPcqhSCxE8frbwTZB7+OxUMOd1zQRKwrUOG2bJS/XNl0B2oPvuAktvD3uO7Ab
SIQn0eW5TVB8Y8ePMckIIthfaa1ROyh0Gl10atBHxVgP0Ees7apc7FC6kcQLtxH1iHFbSwrfW2v7
ykjjY/jTOIFe0Psz87O3wjjFtB9n/j59HZFCQMiDfUjccp7EQ15sNgrsOwksZ/eeb+lryjUfgi/m
2JoAjWap9/HXoDfgQOD4dSMjOJxe6X+Z/P8wuT+7hJmheM9WIyLACOZXmBaa6q0SKFfitiSdCCyY
wR0EvXhErsR9gzp1gemg29GR8FxihTXQVSWMdtkwAkfms/TMu7aRJW+miAs6Mk8RAMGd11xv10DM
cPVoz+Qzz6OlBUTPTBN2uVVZwH9RTuYTarYZInkacxN1I01ISjE5Pyw+izZYeD3z8cPsKtcgQavo
7/M22Ge6Kil5G6CW5WJmMJ2xQBACibbIdvzJylE5JjihJcSuhCsZXO4lG9N5n8ElkTlUiZqxR0P1
TXkXNnu2dMo71UVmmFpAC7nMticaIt+FjziVaHZMXNvR/fJ90BROnY9hcc6hlFfbyB3DFIGaDxiX
SmmYD2nMC/OFau2vgMy//uBFTQYK7PpK/jmD1OqQjOXGB5r5IfwyCle1lM9+Cuf9sV8G2Sk14zuf
JBpSFExMOU79drrKXVg910BkpCTmgsrIsEMDDyBm28tPJjNRetbpPXh7zWC01TxHlze3D1tcRcFX
A3zCMJmSA4O6FShkHUBLAqXrNVm5yoqqcasHZ4xkT/jZO1DxJUba9YqDTm3UY90VKxjS1THFf023
NFFGd9uoF2tSANTnNjVHWqmAI9yE9DEKFqYnIy385iLpCjiAJGF4HEPWhgbRV4QBZSxBN52Xbs+4
vg5e1QXdkPy+A5hOilLLERBN00P1Jc05xwtZrj0dqGIIbP7j+BK6sLM0awpyvxBrkKRQNv+m7gqH
qPjewiBrzt9XpR9VeTxYh5iZMw3dLg3FvVkr2yWNzM1r0xTY02aMWU4txVlfS9zb71D9ngRs0pwD
pY8bWPSYZxBWNZdutzQU7+QZZ2y6q+WYIcVFhJzr9vsGpMGJyIRMwdyZq7fRfWTk+uyUOj2/BIWk
Rc5IZqMf/41uk4Dgkt0g1jm8Jh7MS0nlgb+ecDbpuaC8qg9dPu02MMsBN6HQVl4vaFpS7ngRxZCL
xJbfEz2wimUbrAgeFu2onsysIXHRUGIlp4pxOGqr+MG/t+EQwZz4fUnZjzorjAr5+wIY0rsD0qbR
QGv/ZuemIXwuGGeFCsl6Rteia0O8816IN4quxNDfSf+xl49wStds6L3SEZRgsMEQOTymbDUsCn3L
vGS8bXaA6owU3xyDot76QUGSztmIORAzO4Mmdl8BamPrgWunxBm1omm5hCYw5LyrfojezOAO/fG5
1ZyLfg7+ZOKswbGHL+XXKe7C0xFPqRmy8ZhU6YBAI1k4U3IfDqhnlkezxSUuMTlbbEhfn0W1fjrF
DDP7wHE632nBlg2WHBDa5Ui9/LGkQUApwv/6UXjTbd1s6TBw+LN1nUbPB1BlXCbzhohgTPq1o56Z
PeQAzPDH9j0W1AIqLxfcIoLgZhBxk45G1gyFV4gRFw6s0vU4xwNX4eDLB5gN9LUbfNIblPCqYbI+
NLiCsSGHZ0sRwlgWE9g1oCo6dENgvvrtyOmcJiLPaoSWyPmVwVJMcxRyvJ1yZZ7KEvBNKsH+233u
/f4z4tvmGWCUe5z7PjbPUuxSS45AbmuV0ABLV179nxcRr+DfjQs4mUk9HBpr8SzreTLHGDxLFpef
Ko9sHrCx0XyK/OzRhohRqEuusQF2T7ti90fCjXOKGrp3tSjvuoMg8RzOF/L5SZ3qpAtfEMTXCH+W
hF59Ob2drlYK6qU6mrVdwM40Mhs0hcBa9Ry/2v1YYjAeKUNVT1TZ3Qa6b3hK3u30K+hRU8nKcrZu
l58vxrmNIzck6Xn/ucfsExESBl9ciOmaXr4gejIaddpNoQ/TuelcKpTYow2FSyXAlh/QQvHYTh4j
jG/LwJ3lqg3Jc3x4ZRhZ9HEiOtLgGQ6bXMMx16S6+9pJRQ1RwaiFO6XAntB1KSwIQKlb9ud/VKp1
eeDLlBhl8YPF8KOngn9JtfFBd6FrfLO4Z9edNDDVYY/lxFkX29Lh5fBUSsC3/voUUDGsvrdR/HFk
xD1wiOSOAIh42nYi0/zfzpyx6jBDyUecmi65CWZkn99oljLDvGAxK/7NrW+CNI0WvKjV6UXM9PhI
PB8+KIrfoozDOylQ+lMNQ/3J69yjNLbL2ONPrC+cd9P8cBaZ6Xu5Pc9Dm3Y9AckanVJ21Zg01s/F
ynl/YAoLbFk3kcZ132O1yLstsBWrje6I38KA115bro8tJ98eMj2/+QzdqNjVRDCPjMp2NXVEYOVQ
B0kvxxRwHDtrkyM7t9UYXnOXVihzHxtp8LPAF8hWPMhQT3/Y5GKikOdhl+5B0UW7Qz8HRsKPxnv0
i3pz8Q2OUw3rmtS9Lig0ljylCGErNBWLPFFZwehnLfSsTEUWNMsp6dfoknydT57CNg5FVRmDYJEm
ITwOYA4ErPzT7cmkHFhZh/QtHWJtuOUkm5HSUSEr8sUW+W7rRbQfMR3aWwXZEk6cyHTcdU8eZKQj
ATyxJ9+/BLDxXQRDq59ds2Yq8QxyTymfO9uI9z3O5fyadKhRpiXL0hjVV3OjypxubdHOZ2uhyyyZ
GXYmMrLyBX9Q+W7VVS1cOZVt6vahzTHS/3OBVZSg860jS/5zFtn5+V91tOpX0cfhrR1R1FXrNtpc
SMSB55v7K1mf7LA8xQjP7JEO9iP8crd+uChoV40kI2jvGMkn/x380Gewfwn7zYGeLkXKlI0+lY2f
GsuK9yNzMzbdUqlvD8Z1NbEXoVmaoOgPbf1tdSgD6WNkqL0u4R903tYM7LutRzAwTmUX+vI2JUg3
KEIFueLtxMCBdjX5gaegO6OdKQ6aLrrN77hq5dGkd5rbWQmy7UwXoxPfa8K/GhGaGSuyzkvlPnpJ
fyDfPtiEze3r6wJzYQXVL28+3iLraRZ12EMmb/0g34FIUytzoIzJEfBqLVEx+N0FVqxcsFNxHuq3
GIOXD1af9ph52tqNO5sdWGsWijKyucal/xfVIoJC3ZYq6PMZh8num9XNaBTc667mQ9efOCf6GtQ4
WYZooLPJ4RceRh9KSLXoRhFjYv1t5hledAAVh40lqGuQMwJDOs2+LpWzSeBwwEx0FzidZpDIlaXY
HdZ+6SrDwwk2/q/SuT7datT+55zCotKsqnG2EpD6qxIflQX6U9o2vIM231WPtC6QdmUjTXSKXop6
L4biDgH7o4h4vOBS/TidYfCmITutajgFnYXvyotcQInkhaOmy+VhRP1G5QLeU68Q/P+HlkmzSMw6
0H1BMK7PvA3XYwyetFAQD9dXwZUiBsw5GM3Fzb9iAvh2hrHGjfAEitNg+wVZ8UB1LQSoe4A8wRti
J7KmoSADQzbhh81njy+WaTPiqZGMkTcIXeQwM5fVAh5WHGSm8Dz2t9XMuv05m4RylkZRDYlPgz55
aZS36Rnu8eXqJFkwvcBKecdRamWj77oZQr8dXERYCBdo7HkU/XEauKN2U6wD8gJ+ZbVo7X8MKPfW
uSaA7JH5yQjpIY2ujM8QLsyN51FygNvpQKzqdVYv/ii0C3DGBvR3+m2+aIWtSadeWM4j1hFwgp60
p5ULl5zD7KeMBjNDUweDm+hTZktqT6llkp3mkQ33Cry8P+RaiWUg2kt/I1CiIk4ZZ7JBhtTvwXl/
kpQNcTV8rOMrsvp6yJsO1Jf3cSMG6pNdVxA9aoI4w/w6laST2T83OKoUXxGPfhU9xKuYxo3Z4RfC
o0FjQh+WKPeIdIVhAYvLI3y69rbFzWPqdIb4OjrztyEYf+Cl8XOphG+GeinV878D0t0Q/j7SeklS
oAS7jA6WXV1lKy0CUuOMbeH7BT/7cZZ0OWa6UR8BFRVpYrJrZWzt+tKJd49e+tfQfxddyZrYHUwH
CWxT+sfFw+Jfzki1+zUj93gB1nd9hP6u0c22+ThmTSELDAWtUgDVphZZdeqsWIHF4/QAh5AiuCAx
ZKLJtz41Yu5i1aRN3r+rjx3thcIyUBoXPsILFoLCaKu5kWfxW2Yn3dLfjvjWik1cL0/wP+KJYsuB
srP01x7rAxbMKGAZmJbIOBHQ46sIbinCb74byl2K90rc0/aUdmK+aBIPCwNHH4znCVOYWTunthQX
wE20KfZbu+VWzWnztCgiaa6OCZ532u22q0SKgCb9zTTCP8JFP4qpCWc/+A/zwk5xlIaU31I0eOAe
P1SPW1uyMX443DOhT7rSlEVyFJOV2IhR/STxk28EUAw/9ifa+97U4gxrHFhtbLO02WRezHYck+yo
5LSPd751JsD3alaCzpQ0E7pw6YkkZ2jqHIiAyJOprwy91vd38WC/5Xe3JtLiuoTmaSP8fxfX8r1x
b/5GhWJka9t6/A1fFDd3P4wU12jS5Msbu1Y2+IAXip8app3Lv0iUc5O2Tem9Bsn1VoUUTow+gZAo
IXqf1H2naPAJ04yYky7QjNK6+NaM4mhoeAjIY7zcA/UFKoubvjfxQqI7XaQ9uuO6HsjJU2uxHuLB
Yey0AKvx0k7sF0aH9RBTw9Sh09baCau5hc59ypE687W7P6XKfVMZy2InBatrMiBxrMrN5MutFUXv
NeBaZfSw3GkkESORyAtTVi4AH0v5lXcITYIbLwh1soZk/bAw7o7sFBt7qUWs31QBkGlSwA98/DiI
4XIFrFBdepTrcMnDIlzbHtAOmGMYCrhlAJe7UJm9sNXy80a/0vosVhyUj5B/8NsfnXD5c0+8gPaV
Bdh5feTRafepjtY0hN64pKfkM3EJsYyFyLYOcswrAlaDU7PBr4xAhLxwv3UmTChE04dyrOHtyaA/
iTOzBIIfz23lf3FIxSX7HCpQYEDkkgca7ttWUNbjRFBg6PBGhUcBv5WwPql1+dspRD6dbqLXTRIb
oSPmZmAbwiIWkcDeB5rPWnQ/sWjASO+IYBCvZY7rjXHtK9p4n4kgR/+ar17n8OoNpCBLDCyCe0vo
yFC9tegfbE5eOtbC1xuVNs0YAyLW0+Sj86MZgE4+C3+nxms3jEe590IFt57OHx/o/e4sFeoUHUMB
DI2q4l+3ajlPcKBKkZaWvjqRHZw+VDB4YIwKvhW30UOoLJ0aEnVFhecy6J8aig5+wO5yBYS2zFqC
pXphqed6JgmRnf0BQ9hrflMsZ+7hOjpWdzqYxQ+8xd4JP8blyy3G1653r6fOA6X9YX3nW8AR9JHa
Tdi8gRtJWdmVePa2qGpTL6xWFuoLUK9Ml32uD1h2+cf8sIxFNdswzZlqmOISQINzh1KMLGB/cCjt
6f1lgfw57QZxcFCsBwimTCFVMpLZ3RbSZxACCEFO3HGsNRZtx7aWzSUsWRVVOvpWajJcfA3pQ6yC
bCd5cMKBYg7UoWD2O3tU+r+rcL0HBE/JK1+a9Mb+cIvV3u65FQMXhi6WXIUraw8mp7219rNDvpsw
lvJsuoivXJrQVVV74QTcfAQx4i53N0S+FcEkcpCOM978S8SOqVp60G0dznpPpPn6SOSXFXAfxHff
aC5hXWU5xkJvv2qkIUimahcKxN6yZMDskm4+LzLL2RpFfh/95VRPYOMZJn+U+9dm8ZWhe1uFXX4L
BsxTBhtVEIMPkY6hcyQqrmvhuWT//Py08RcNBDQNQbMwPaEQuR8FfE46i9sZmihMahPfMPAknhoD
zD8nx8bMT5JlIsQuGe3Kbj2yN5WeUk2tWX5upb0PdMG9ZLqmotFazEBQsLnaciHR61rA9R0XyLfX
pIdhDaBXmP0uUNuqYwOALLaYAb8YKD16nfCsZIPz+C4xnQz+X5RbFWdbofhRhHifEoj9T2KmE8wm
NnBilSnu+Kvn3txz4LxJ6fzu5fk4z+AmovObyxOZgOfPaF/cqrjZoYzc/TwB/+OfkVGc4C7MAaeY
Ugx7piCeEXuTa9UHvQGTENURUmEEQU22fv5w9btCglTnkh726Gx4tmqy8zxh+2P7u00qoCusjCXG
t4Q41OgpUyx2h7DO4ZpdLevqhsTuJaw/f4nPBb1P0tIM/qNKMicr3h1wWDWYl6UrFlrBfZPirY3r
FKxWOwk122ZvIjhdMGMcwWXusP1Fs9B0I1kB4HLCq8BY7JHqyVq3/ZgwYw9qV2+YZts0W3j71rC/
eo5ebFJCvi+JORAzT4xPXRsw2nXHv++YS7Ry3pACY6y1w/KPHNZzMfQMIxZcQqLlXHeitwSFUD99
+3xZoi8q8UvYMlLeUv6Tr18M5SnVie7j68kpAHDDREGRb3T6wSUw4if3DuOXHHZjGvBZsXwCbTDV
NUZ9eK3AolJwuknrDbEVdwILgsfTKKG8yHrqWlCzH0aRKAtamycF6FymCZiEHzcj6RlpvXHK6wC1
c9qVV+ubCT0VsQXlzJteX45SJ0sgwP1XGxlgOns8vzxI/5LoFgW06SKBBKD7u6tsUDDmq2tUUd/a
2Io2QdXGXfSwTdbjgRjIhuEQjjFc6OgN2nlz6+bBocSS2HFhRJYJMuHOp1tZN9uEbzQ00QTGKlAP
40+9KjyZ/K9T1D5flfrFdUzUicJ7n3Jlbqw3rt96hj5bL5+euEjgGcuHaac/oADBWIEgeF92iShq
zBfODHGlLHVjfMenYI0f01uqX+AsTOmC+dUaylJ/n6rWDRtT4q1dXzzwVVJCvkkXtRKM3P/S3S+1
iH96qUGUIGLnUBnYuodycLC2O2imyS9J8txLUBOJtvJtP5bDZarMDNvIs4HtkR+OpE+1HGXR/Xfg
/Z0T0PoHNSP5l0qOTQpc8zp9BOK9WATb8qBOreS4PCzMCpLrWkFAe/JOFSnoSBByiiYichCglmRT
dhFjqYutYi0Nu46IKRqMKrlay0VaszE/peOe4VBylkJSUPHM46PZ82xzK5yHEp7i0iXfvVzXF36W
5cxEx8HKfuu6kBKjStNiBA1v7oKU5Cj2oZ6EAb0lNcpTo65lspMWtxCyzgucxmzHIXKhmVRwlqw3
3YnHPPY7oemSp0Q1/6d2amr/pbTESCP48kZTjz4Cv3Jn3l1TS/iH18bYjrvDndIOS2dZzwt+T4aw
W5544QExmAA9ha/lt0kJqAVN7NW0MUTD6qdIRPknmdxEQmUn2UQjIAbvBgdDrxGiQC+LRDZI534c
nSkfXD4IaYL8YdeQJ859JKcTJmTIbCPUgn3eHwPNifpUe8x3FKd7MgvSsKMxRVxe7Ff4bEsEtImH
g08r1VDkNo7zfAvzCCi1qEEDhKT+qDDSoJF9ZcRi3bR+OMH09zX03+DySoAXIA8p/tDgR3e9ef79
Ux9kNh67K2esoZu5lvj1bMvkjwdvskM+oWgR0u6ZDvaSm4yeLh4PCt5a3UwbEgI1jy3Q2wpw24is
PNH9+bzL8uS//oXZhN+Fe2SvsYps+cIqHVqtH4AoPJgBVf/aWaTsuokPAW6oPZLieQJLF8x/6x5+
rEJZnmg1dsf4ExqzcriOTfxKCrR503RF/QmOeu4Dqs2ahUSzQGWr90G4VOXgSFt6kKBIJk0PJI5o
74Y34zrvv3OE/U7VZOZj62cQRdPTAfSaQjxqzkTPxeo0HFuEOK7F9B8HJ+ZZYNyTVAPwyZJOBeI2
R12VkY2QzRRFQwQSglLqabvaTJLsw/fLwqiNCAIrKPG98Kou2C/n1YQunfePJkFGiZs0qDLgk0vp
dwEMsb7I90dpR8s2guF2IYL5FHJZjZ+3K2J592LbBVR+NZH8lvkrU62nONSSCbMd3FOTuBK5LMs+
96zrKmvCUd7Lg21rBpsS4IR1JcGXfRcUulRfrMWchm3pR0jDQlG7e4cfGiOo2+LH1+Ewu9Oi9Iin
5BBaDl9TyOlZUsSfNjBuHSzZ5A60uFKn24TjErqqWsw1sNi+I/8iVsKOghFjMNnwsPR9YC35Ks6X
Wq7Qk+8/guaocQ1uPx8Bv3pMbwUMxM++tAEsZTDUseJPY9f5B5xjMB2D9x5n9YTZIZiGAAileWo7
Ojv98rtVFx0gU7oP4+5xdganuvbhF68wrLQQVFeDbv90/L5gRBqzLWbKSOnH9hUeegmwFoZjFrVM
Jp/z+wxvTX7Scx/51EO1yHZyooDeLM17m/P8g9wHP+nPvX1fjbkHSjMD2lTV+0Us8uSYUJ7IDtFW
ZxmZoHjcuJ0BlQxZP2UUegfNHt2Hy3unRdgfEC2jPwDUSusramAZGFK+8vD18/nH2+h+VPT652PN
UDlQgXYPYJtvFg7tSNxeOQVJ9JPNX38WqBFV7lLJi8QCpPKNZ4bTVcanbxdaiOPD3ij+Y+Y/YhYg
WLAV0S0yp9VUQYtHJnvDT/FpfaO5cntuXzIk82ZlYXD35cqk9wCNVofr0uHFp/5KXogpL9m75kyn
rZDTN+pn0geO8x3Q1G/c1hnHH2u4YzTF8kV04/BH9Q6uns12u2p/54knMpKCoVVFS0QEoIG6iyLo
JAX76LUELuUY75vQIvgOyU/Ydozt1CDbwzl5zSNW0Ou8EWY4XqSOzzHYPI1PPKzLZamRo2lzrwL/
goPrlwj2EmwYIxhuJ0x4W5uf9iRfShcDhBYGDeamkFMXZ1fipAdHlt3/SBGiS1mDG1nEYWTLZDby
sHKrmbojOMgXABrtzEunvu8HQ2JjbgsAJUnyQHmWfc71a6UoSnm4RZy4ubS/EvNnDb/YFfxmvbRd
7azL/XTFW3Z7e/xjv33uMRXnHXQOQecXrkrdgELAZv0B13Wlp0q/i8wq16H9zMGNLIou+hLYr3Ik
wAG73nyN4MQbxImPj6d33yO8faXgibjWoy+w/NWcaJ6KzZ8wOtk9YVUhs2HI8jeUTLRM8IOPn8sv
qWmqotDqrTf43FABA3hAEYfUpkZW3Au/ugdgaCUGF0hSgguxMma0ssLx4eBoZUUpprqCjExzPYQ+
kBD00dbA0hBJzaQBraXq1V9ZnGPPm9HQuEVbM/GuBvADl2xqtOz9ZqkbxYgdxFax81BQHjHASIcW
ZRv5BroZsyTBut8p4yM/NiMl8qMUhvvJKJtLDDIMYCdfisCaf4/+5wySOKU/WMccQrOzNGzvhzzy
rtBS0z3W8pOsfZ8O2YbD6MFb3TfEcnnT1N+9aKax+FVFKKzWB0I0YfooV5SAof1HOznooLMc+3zx
Jo+ov2dyM+5KESc0JRmRJwqdfp6gxgFZ3GwSxQT4+9fraA7Vb+xDjHVDgZ7NBoS39Yka9WtUwnSV
bSasyxoiubGH/JI7LTw5gunTmYMD43qRfKgPOOtO9DhlZxCFPzOWmI6pCJ57E1YoVvSsHENDP6y+
3J38j+8eRp1JZ2M+YV6fbmyBr9iVUM+WCRdLO+ZxOmem85Xz6HineTjeGFkD3M+B5ZcB0GsXjxQS
kz5AHv1+1k6FDhlUeTBj4P0mn29dklr4d7q4ex1Qia+2F7rfnPSUZnAdVoAO2YQfa0NBbMUZcHhW
iNGN06mw1mmSlpjXt7C80MkM1GBI5DOs32PLCkKi71ixy1/llVyfHUuMUuCG7srjcsUydNWTGS5D
H02LrMG7H4XT6rFfZBbu/JUDryjzPAbktMVuG3q0hB+Dr+QsrpXHpdmKSRbnVCoM+KSWLlLg46AW
b2R957p9+v6W4g1CdHmJsva1U+Z00Bf1wsa4pqOE34PWNrbaXEqxV1nqK/w7RFM5PmDcKJYC2dCk
cEdgX77q6SNZBRwi8pBUJ0d46wKoQos4xxdEYdY0NWggvTnc8UCfZb2OTLvGSRvzHlF8zbRrMBC6
eT9Gg/cSKpqrBlAVKZXcu3UVBZIr/d/1P/1cxoazt2LFSMXUfhzhe42MZzDeHc6qQXSxBNippPd9
vp85Kp/cJjcpsDMlrLZ+YlbtkVYlRhW9Fy0E9YodRlm+MbhQXsOFRjWRthDZTbrRKHrAZYjZD3Mk
oXj5njbO3Cglzwa29Kplv41CV1asXVM3/odUsSM8H/PkoFzgOfBFQN5dYk+zVPIis03n8hVRc1fl
+i8MieV9NmgFDFzG81L2pghnsokmFkhIoBrrfpOvqcfgBSIYeovfKBKsbNB4nb8v3/uPeroA9yRT
PHdsg03iDvoRFJBHuMSuQLkujUMqBkQFUUjJEdYhhPqZfgcS32gxDxsY4RocKjqFc/RpeQNsjKBW
PG5U4k6TRMo98gOAaBuv48vIGS1DHGei54Ruh47rtChFA6ygK+7MQcqN22yUNsskDmBL76nb6EMK
DVzT1wr+l3kJZ4/trvI1nAm48TBYuPANjm46lEqt2HyHyGdE95anPqiHpH/5DOVlF2WgOGtbJbxR
mqldyKzNqLo7KNdSXYMMlfPAO5DvGDMDPTSDsf2ALS1w+yYnCFw4JbWzjL2X6znP74O1XAQ3eos9
pamLhnM69K8QrocuHr+Gw4MFAYzTiT7N2fnMi19jaxOVMZ8gUlDcLJD3T4f40Mvig4nudIWqzGPp
L1I9tsMU3HDpzqzog84HJGUw1sn22sMw3AHE4xc7HJtb3zrjxMGHHYtrBI9I1rZr0YJ99+7zBBNO
t3yyPWHlCrUxatVf6WEdSQ+cmfFvAvns0JKE/i5TEi8h0UY5+RIlstpr/yrb+GXRjnXmfLys9FN9
NEHNvOivnJEJrX98/0TDGfFyj6zShJnD62rt5cKMxj9FByqm4RHxunfEHpdQO5Y+MgWPQ4PUE+mi
Uo3MwjbwVLxJT5ZZQoUWx4+LiLldc4rw2nFb7AnlGuVwbfn/JCYUlIOs7U4Qw68JBspYYNKrEg6F
c+sJ96/PJg47WpxSpidLNb2jmBIC7YvjVkrcRRaR6mkjwqanK7OsvNGBPN7ja6tGN/BObHSupuqZ
ycrIp4Ib4Ib2OmiBKqkVSaZ8azGBEPJVHqNykaRMV/x+dwy/644CwUHPOrIm3ehg8os0PQ+L9HoL
n1mMGFow0zVbFwZ0dvhtQpMlyN2ZWBYGJSmzkm2QJsP8+o6JTef51hUwxla1CjZg6Fmt2TRG++6f
WfOJKJ06Ae1QzdFczP1KQ7QHvnxzSUCpv+wYc+tQI++8wv/otZ6/IOjX1iJ6nU6jzKN0mq5XtW/9
s0rP2fadYDatAhqYonGZUHfr8GVzKMSQJP0JpWh3iR5XJSvzuRnnpHz54vO37Fj2WaVTPYdAUn09
ZXqq0zZTqt8MhCkbj4Gp84Sc4L6kOJKC1rdBVrwhxBWVt9iR/mPfFDF1nYVV7mcW1um/jTry7+dq
+TGiUwzLr/kFPeDU6YMleUOHUBEyRavewoxai7+K+iUHhyEPRHL7VPXLCFjYSbHSiYNse3TDFmx8
J9J3DPpzTABatvUsbIq5sdOu+78iEQSgHp90DMyq8nVPUQNCFCgyiCTKYQb4XxYfqUYuL+ICdhte
DBxZD/8PrKQSyUNLAAscDeQYn15gjzhS28dOYyArD94XU8pwJO2w5R4Lzsj0RofQuJ3mzyqDHax7
N3qE8KtbWK50vBQEOt6QzRlzlpFFHzW0Gj4nNOrZlU8OPOT72TVwF7JXWRK2fROx+Qq8sIgCncap
HMo7yc/RCfpowEMZCcnZbysahuxss5aRtX3BQgC8nUpRjqJS17jrZwhD4dGpQaxGxRpF5pDpgkO8
sW1MBKfdU9HwAmWkXSh9IYqeusd9p0kHt7qetFRgnM+MkvOukzf82p54VTMwxJyIXVYDFBzcN2+V
O+yCA4nErChbeivO4ECr8r4GIdWZfZ4DBBfui911Jwp2DbHTuihL6s7mU5BvptCH/CBFSxHTj9ZA
LfKw3r0IrAod35W0YM5wlMvpVKPSyL93vy9r0xSflgraLjCjXqqpRE3KOiyr49XBtYDoh4HCjcBB
oW4HrhMl1nyp2yjDyVR1lsRNXtQb72i4zwFsZ1XgLJpCTN4/tOiv+gaOCueY4C9ijsyPlH66Euxt
aVnT8BFfJ+HA7RoLQNpwh2ZY7UsMVu771nviTV5WEnaiKPYHCOJko7mACNStffzLo+MtwU6wHEh7
FY1IjeowL3SHHcKiyMh1yyhzzCaTu+s7LEReniZ2cLfe+GYNLWOfeADx1GkWfFWufdus4D2bjvaH
ZcbqUJkUb7RtgniBeYzuHCp+P6ibw/bAiTvz79kcBup8zMIAe9Hl/q1C4vykRRuCSaAwRHTbRj8T
SF9rFURGd5eteJRt9QO0cDaZhAKrl4gh2Olai1pWJpNF1yYdP7YDF8zy46jSCv++R8hM5cfCGmwg
yCsS4d8t/VjXp6Yj5Vg9M9ianvfMuVRHRVzktHGQMCr5N3otibRTXCqFibyKwoqx+RMZ+yeoi5Hx
DEfoGJ2KMR9EN+aRn3VHw2yJuhoyLCOjjJ87aDm3FPAYxC2DRJPzJ9cb4vXn81rhVA+FT7F3eQDh
jLxotgFSnCB3YfgZE8c8rKNasR2fbpSVXNnDDb8pT+cqWHS2+CWAXK3iO/1XCBB4lOy/ipEsk6Dq
u6irJ5EaheeugEEqRnN39wPYCZYByRH2CJGKtlJHmFU9wbhEgDmXwzJ4lhWoneHAdn4smNXI+3L6
eCeRTw2BEOuBBq0kI/ZH5j3YTgESwPek0yd7ov7anEtFy6+sMnJKJkR7fHeFxlD+YSTZpLmBiYRq
F+J/Fb7NdPoaaUm2DSX3Dc2v2rFevM7sdmI2mLV+ETlNNku0lHmnE7Xy9jiGrSwehVWN7dEONJj0
5QXClJDobwN8dtv2hy4FyVjfuiLLuRNSo/f5UZpUMmesGZtFf5iilFaL6jjlYZDhW4xCb5Dja0VX
kCn19jOcOQEO9hHEnzpnZr/GSNoKvVAGPLv5gRL0mnnPhJZ2/IvK47QYxAorc7BMC/E7VD0CYfDh
7fp/Psv1MrwvRlpyg82DDCyIcZihF81g8hqxCPtHvRNHMYWNfjYu/puQ8NFAp6y6Cr8vMEefxI4G
nXZ+PhlGRKSTM8AQ63bGBYXsj0qu5E1nIhMNz11kwvtN71nxxj6XjAUr687W5rXrYLkbt46rxUUt
EhKXYv35d5B2XzoKAydC2aB32atHVNN2NwalXf17YCzPBzWsPchbMIyCmy3l1OpJ+uWYZXIEeCql
DTyQBxbGGYog7LEgYFb4HTfKbOUscaCfhlWTG15dDuDyMCv85p63vHnc6plUzNvuU7ErEXWfaD1/
GsAZRdTel7c7wReBwa/Lv8Yw7D8mAOF9THlKHtlrPcZxhJRxSIg8qDDPnk34LtxukHujP8JSo1us
LDLx3lZvrB9d7ZUNBXZ2ATmH6McLoheZdN8fy4TLBPl0tgFII7w6RZE6kQKGCdrW/gYuq80Tjp0D
Jy6x0yu8Gc9dF1ODKV41LtfA06IxFQJFCPYR+AQwtwb7r+di+X8fn97SYmws9Z5P1+OwiM5ReMFm
XkqrTFQRjdrMbpNPckaLa/g0SluzV5Mi4bBt2e0hY2i10+gEsBPqLuBiZI1Vn4FdKZhdK75XEq1t
7rqdMH4lSzgPLKGkZJDNMMap8iME1gRZ0Sz8QW83/x4BplHfi6srni7SNTv80Rw3RF1Xee0IQDkb
+29ExOmoR4mN9NAga2cdSj7oCUH/mY7rq6WNsJXjLSeXAkbGqxpqceEt8Rrxt0hSWsxPA9cAvzwM
05BAMdU8OtfrXxq1JK7VhG/n9h87hQPUpZrwtwGiTVSLs0b9pJngRqo4CqBYgyHnoK1x+5OUFWLa
5HL1aGNcoIIm3GQ6KuEgZBbDj2I/ZqCBHanJTp0c1ahY4+PeSFWe0jsujxAiN3669n0VxYRA5vH2
0c8IQKWH0845eh2TDVFewZo9r3jsaodSRZktqocrzxub/mDqB7AqSQRYSRplvHzXtdynzYek5no3
kfWQt6B1yYBJyN3hglpkn/2skMrHKRi2amc0ML80IzmbjcFtUGftRXv51MJch7CX2tISk38TfO4M
KYjayi6rSXK5zmb6OfuL08M4c0qmDxv93/yp9xvL329wMeeVUSjWjcFV3n6EuIgrIH3PwygZlAVR
/ucV1GkBLVFRrXMm6eqq4kNg9RTBkr5Fwv1seIE31Zt6ww7rP/ySA64WpCfBS5KSHu55EP59isIu
haUcwJaQRxZj3X26seMtJQhLY5zy9Spp8vTQTbEv1S+BnZS862zfjmJQub3qa3d2tpqZaIq+6B9p
XSHUsV1zNXhHp0Tl68AYPnG/h0l2FsG+0nsY6It4KG+VIMmmJCKGBXh1roNy1t1dZLxMDOXoTbGZ
6Bl83srVEGSdQQo6Gynf16f0M9ArLnmbZml2Cx6vmdPwhxjo5UfDRuAnXySYGdF/0pml3PeBd24w
GTmnzS3Mr4jFpO0tdPLECnYbcJh0JVBhFtjXLLE4tSHebtXD3xVW1w9OQm/BLIClYnnPwAi3GLpn
81UwR+84/lXhu+JQ+vLXVATppp4WOSBAbZ8WtiOiMEFrlTdXgNZepC0XNKEhX9jtOTHq0qYm/h2s
3aJAsOrc28DVVPHqhpWyOpG/ncIaBbvs5FghJo2RsYDfqofjd4bCOQxmT9yx6e3Ce+T9srkIKpZi
S8CHeHMj1iwm/PmS5YC/3hk5sYlQsNOIib4vuQ/f4jB2ndOyYfUpYM4QYb1vAkYvegwU+sHNJBEt
lVecouiUcorPwGr47HJ2SCxTcxEVkrke5w+3LZKVB+GkWClUPRAfM44UPEf4u3yjDBWTMfu0My9z
zFmOSbi1xALkpikXNzPrAuH4zG3QT75S3dytltbs6RLNgme/IDq3mssKBOOoEfd6g13IJjLuvKbS
72o5hUEQ4TMwRcaZN7jKX63MTseKO5ncJb3cA1o07oMId9gf7UBwMTTpWkwMClvl6BaQRMeYY0lR
u6c8ox5LAJ9hS4kkPYsfqwoJWw6L53+aA583glZ+9ekheTrWchhE10sEnlKgRB22hAIIs9ObQX3L
Ce9CJw+kL4KcBcznXflc+vOaG2p8TnCzOYjRIHVHAzyJN6Bhxn0iaNSJ1+jp95ik3WCFafgcsech
HqN9vdxueF/iBDUAnaxlU+aU24phY2TS3O7ceec80Pbyk5kCbhKtCb7QH8aKgSwMxtE0DvpE6axX
jmw9Jsx3+z1EcFpIRHxWBnHp6FqNsi30eJ6s6J+kADnyAtVAsz1/qADfvfJu7kOq+IC6Ts8097S8
f4AAagjGntXhbuQz6SGWtoxyy65bu55K5Ctk52zmDrD53N+t3SZ6FaM8DAhHu9JQibg0FveL2frh
k+vT/2PsSeoOCDAApHQV8aqxs29+ZCbO2BzWQWrak4X+hbF2j+1IwvZsTU5g5Vqq/HtoDykozH0N
KlTAseyOuOWnASUgVONbu+kwbr0z1NOlBhJjZQ+1fs4wTDtXldER+bwnppSyercf6uYuiPWe1kFJ
XthdlnSOTsH6krnIj7D/myY/SenOwi9HUm2J1Izmbn6h6auqYTLbFbUPpalNSGtIbCsHJFw5KeRD
tcUTr0jc/gb7DgvSkmDxmZF2DOOLckQl8r/oKCI/4PvrWeIxptZilX5PNq56U6Q1yxm8Y6yB5RT0
6xGBaQptdnFF8taEf1E84ypeES99bnpYhyoAFy0ShKorSvkaejKe92MztWQiTmQnsfCnyij+gLk7
cwhrL8mc+cS/ja00Gv2ocMzLAhJVOjkpmtMiE8bdA2UwaHoa7OjMUJdzSA+cuZR6HG4MIIOt0mvg
FrgHuYn9vC431F6417NIrF3gwPL7pls+L5wUAW7el24pNZeXrF00iUt32+/6/vei/XCUmsJfuNVP
CAH3XA0Bdy0cuRdtb5LrUUP82SgPLJaCgjzDiNH5WyYou83nWW+9OzkLKrvs70cPo8fS/0LOgyXU
32tRJ6/T9I5KoAis6Y7wormrCsnV5z9AkMgNFq3OvekArz/rEATbr29LkIt8DPgNRy9QiGRT9rUG
Leox7zeQVat4+1EHywc6v79CLaR6+kxhQ7o3uohFvQFXkZ4CL5FMLEW8hGDPfW0b2HckSKV7RAjv
uD7a7XJMg92CGaxVg5ma+LzBANxrvy+y2IhPMSKaGxdP4GYXueics/YNb6Tp5TD8+9XsJWHdY48d
+TCC7laYXLHt7GJAPE2IpKH4e2mXmyLnDzTdHMahJmv4H5SjPQJgcR0d0UjuABK1DgYj0n4njxr8
O9307l/fFLZzOOwMAqc/myI/s578WCuqFpUBFZ4h7rtvYYPDMa2E9vSQbUQopHFn+Sxj94mePTmE
F0oLS0JMwpTUYVDZvJxphVA632a6eY7rJI/dFZHoBc+MLW6miIAGaJvYeJ11tkoiUyxiY+tIkoHc
g+FmGdxj7LteFxPJnRhAIoqH4Q1aaAqvjPxepffLtwZChABRBTjkBHfd8rUVSx4EF4TrYfNRiQC6
XokBrFTmhctwBZP0xEHbbcPtxdNMhHe2S4uPpQEznqKgSjlC+duEaiiFsT64WdLeDsliXzO7dQkR
iF/hxu18CoyB0lULtCAEgXxc2PiqQX9bDNQOMwwqKON5JVknEhJMhVfGETlKst67eLnt6HTD9opb
JyghLwAyKdleFtUTYjzuozhH/zR/eo2NpFYvyyMESbCfOQYqhNlDDqv5c5F2thtYfsc3xZFC11D0
GJckv+ZU4fa8nPntCgwyRELwxzsP+2MKOH1xyqN1vKfQZMm/78JU3Kw7mdlPg40TtR5RCOkQFz6N
V83cYoJJHVkhMfCOqlameS4JB/Igoc1P+T1sM9N1H87boN5bVTu0NbtgBI6E1LLVfJcM7RnliuIS
EVt9v4v1w0B10EDIhO2UQ2OzgYwVxZvXTJybW2M7ybPY3MKrWMzxMTo70HAkE1oeWcaJMzlLuYmW
W6B2AxMc9shMZzFzBwe6KRN3WJzVPQoUBb7j5gBmq21PpNXjBKztW9ffeX+1+EwnCpWq+35ddlWd
LBmrMDNVs4mEqW/AwunfNa1WGIn9CoR2X62DHlQXU/d2Md5cd9llLVeT1yAspdpBxm29RB63MXgb
GUcRDyc5LvQxwfShf1lWQQPw4Aq3C15pS9Z8zEjmyrBVfA9a6reQcXOJ+Bgoi7fqp7bbVc5wmfhk
w4C6LY1ZxT1/GO18/R81CVjrcVUF7Hws+5CZxE/PiDJn0s+ngjMI2UAk7EjwRsUQHMxvvztuBrLV
waQnnt98pv/PWvVfcI2OXNXbjRCZKf+v4EtqFL+f32yyZUHmq02ZHJoFPkKkUPlJobGr0fFF/8gN
c0y+Mch/shAW1E4rLwyZNvUMcA5hnuNDy77+sWpuXVgObcUYv+kZR9smvCW5N6m8W2BV8QFCfJMV
KiSl9dQfECtbPFh/9ypAmZcSyBi/x8nXhYGO4yEzpErh0tVt1XK7NVjc+Si057Ab8B9J9+sM38DW
NCkifmfLfs96HuF4OMtjkkDU9OAEDi8NWoXkCwm/aRsIT40cDDbK6JlFfemCnm1qc4dG3KmCS7z0
nlem683Ux3abgmXRuvvHho773QkraxNiHv3YZexh2Nj7ySYJ3npMGGAMNWH2U9S07MEzGA3JBgsY
7TKYjmsjUwiYxjtbeC+0gmHSijUtB0PM2QuifHuG1b2wcMIzSXMLkNX1vnTaj5a55PZ+YYuyE3jY
DUfNn83XuB1g1D4pQE4bnKL5pB4Omqlf1I7WeZqsAygIZsIw3tAnWglNPwViS7iuGiV8Xj9R3h5D
H/Gu4f9hKc87fSvaM0jW8/y/prpAugiOXcMdO325RSrmvouIduUiNcRg3aGx3Op1jrE+i+bwKq4W
U+jJUqAEwgKn5GHc3m4fMI5cRM0VbPbj+4VsLl1wveSlCvOyOoC679It83+sGN0jYAijMDF5s3X2
8po6/vSoeduOYhyth56V7mOYsxYUKEEQrqS2XD3cSop+BHuBGX70c0KdoN/2rPhWR9vU0Ax5d1W+
61mRGlEtCaAQHbbojvFf3zGheUrZE9Vn92Mz08Kpz1hlPYqYA9jCTAJj4pskm3Y+xEWJTDqQj14c
EsZSBXUJR20dXSonM16bNBAj+majY1cD1JviFKxKYQSPIS1Iz4n/SaVpvbY+LzYRFsx1Oh60AK9w
o1mA93w9kvTp/rKvLfd8OkAjfyC2J1c/+MVstL7OtMPAo9L9BKBcdOLXfsO49L7tTvm6VYEAOBXM
mSzw3P97nYMgufEwz8KsKONEzJia0CoS29RKxrKaMf+h2rFjYnzmOX31nxwhar1skWgiFggxJkRG
OwMiAKHU0oiXPk1nW+Zjt6oYbyCvZnGZ2zA9yX9PTQvQ8FLMMEi+2Z0k1+ye91OTh8KpyB7fkG8e
vOu6WCp7/iHAx3pw+iSPZswZcZXDrwKqf95EhrUnNAhIxL87hn72m54wt1kYqq9VzKhusjVnuBI9
CJnSskmQb7l7Fz3nuZ/7cowfkrSYcMmesXferKWQv2Gu6qWcG0AIxLc63b1Ut1PsHIq+i0GFwLYD
76D9OSsOHrodKxEkyQghC7gNI99RSxZcb2CQr4IDchPR+5SGic84zxwpOTuzIgVqsMYXx7Iw4BHg
+Nb/GBzESJcUr/tbHjWQexlw4V4xguD+hHnbUzkDCw0Bmm+CKq2DonOicpC2+1inu9kRbCIXqPdV
A5kOea2oo+g7HPYbY2PbNITxZTZih3HAZjXt6yowm7wkaSu3yOcI7R92mfxKq2k8iR6cla2q+O+U
Dq/pjXRlIm8JzLXxmvyxrVfOJppgyKUBLLVjr1Qm+cxnCwmnZWM5oF2S1J4EpE4qdLjWLzTxxG8t
ABatlu/cNHtb10WP6PwXq3dDCBIjz74aXXNZxdnfmmZJew1u+AXTiNnpVc7AcyVyzk11588Yg/NQ
d5uZX5VV0wMeCrAfcKT4cBlbkCTwzmQIxXOZJ8MxDOamUrvJVOoHp2GWppXy2nxbozqFAUUrNv1U
v9mLg7tU1HfgC0anaFEe7ZKO8ElGCfAk5DJlWF6kI/vT8gY8zkogFnpfraJ78yj2Hg5rUjLDU7rk
YEChbBRJsyFckIgW/4EftPK9dGjd1vg0VQZ6+NCn65fz+EuxrHv+d7ZMYXrBMtT/DpmUzQ4hhYK1
+C5XUWqzoXZlrQQ3rnGLoGCN2VVlOIfAIfUWzFP/cxZvT2r2V/lZqGVYFclHWkMsEEWf55BYIlWd
eTQ+TEibgWTJK6fEypcq06+hLsBEBrqUc7KFZR6FnS21kzYfxExk/WrGTPY3gwcFC133QTBDsJr0
WcZIdGj86pVCJPzoF9hS8PHYcnXvJ2ydhvLRmcj0EKuiJWB58OX2Y/wo+YifkY7rnsuUKLygx3Lp
Ux8TVOVKQMAcjBqBOOfMpZclUk3FQe+iTe6AwZW4rDZZ51+hwMaCfvgWwTKPsd9EoqZTEnAcECb9
XmaSw323pc7YtK7mQHxZssXhT5b0l5RgFR5TpoU0FmWP39eMHYk0HTew80RnICdvRKv0edC3Xnna
VjvoqvnqeziaIpxFVNb0b3COfLEJUDKhdOt+cXC87eqZFDRZ4oW/O/oGQUFoUufO5w7sWMus/YvD
U5bEebznmgjM+KDi1XgQtDUFv6R/NpI2dXa++VX5qUQG027F7Wvk+N7c+Ho4/qyyUkAwdEJeB1gv
/QmArUFcPn2y7BB+/CdrwCztIAjR9CxhbmqgaED6fEnsYJjAEHZtOnKsB/q75cogMok2pWsDJC8Z
c8L7LcIEqe4iD9BxwGTuY/XI/rCGS42G+dMkHRLB5xRq5v3qN4BPYEi6xv2mbRvEW/wUmVsnVTMD
uPR22/SXE9OWDfs0oG0lCNAHt7TcLWHB22ZlnMMFmK2BrD9Qu3JUJPccRUHIu8OtTBchbyX3qi/u
iKGXBjuppmB1ZsCmn2Yw+Ja81fjRZeC8AeBpEWs80madJcgGFDynl9YdQz3b4So1drQldCAA0vnO
Y7Ly+yNi8H3/HyKKSYC9xug7Ux5Dfx8DPq/HFBK3+XoQog7EXj219jNu2tSUEJ+bCJ+mO+S7wu0Y
1RNZcfasrzTrIS+fMCiXZgD0M9yYtwyfyQqfReL16U1Lab+vlAjz37KZQVXvfZd37QvhHMlFxRvn
Bc0FTmHMyZLiuu4AamIQTYxc9xSnocyjNRCaakxstcMQzdIZe+1d+9P5QJthOluCVgDrJaNS/gUF
7URGOdoo7mEXTexhwmncuX32+EQJH+OghUEB6+rHFcuT2qZYIvEB+BAJI+XPObZeHSvwA11D0YpR
JBOjHtmXGjNA9QPb5WpdvwmtijxDwueZJ9gA1fx8DLZuJSOK8uOixMeTWP+k78UG86m7a6wD9479
GAFfrLTx6Q6f2Ubmt8d3Bj8rb/zTqmEHmy2ZgID2+tou0QZIf/GdeE/nhUK/4KSmA7qhslSvwF43
OJDtSYzYuUJEr04ZZuKCPcDklvsi2eEt5sRgrkLQWxleroZjvqcA+4dmzojiqEsg610kl4CWv7fS
4rE3qQpMZdAh9aS8JJsPqGPDT9mmytyAn41jTPlsWoNJesOheptLTuUnWOYYoF2jiv/L0AAIhPPG
0KOPHKv0MY3ntiV3MBAHqevNDqEZaGvrmHLeoP+sZRcb3WyMvXbEJ+TgMg4glt+ev7/TgUXWiTyB
fc/SXE5b5+Dlx/uLV6eaYmVjPOsqHWS+p7FwKt7PB7r5Lk2b/iiyHwrVTsPC9BZb8gN8hrhdv6xr
TLZXiC9iVQCFiCkNf2BtyTlJkuw2XZYTlS9Ico3kl+ZS5knqkTebSgcw2+C3n8f745VYv82xfGvb
WX+7zeWMgeeJsEQwghpRq8KPDTof/KxJ2puoyeu0LNZw+cpf3iuPTLltLcAAJLOBN5XOxJMjRe8A
o5ZkFtnG3HXOCGYECErNoXLfUwqPMluEfyUmyMQ1aaxVtOSUzlLZYsIErDloucF1fvHhVIqECSH2
nsbP4pUm9B3K21aHal4/SqtsGXdNO4ttKTy50U4Vvdr3a49erzMua/xdCAOxEM/yRhzHwu1F+jit
3kNO93tNSJBFKkmkHvGo5RNtY1BNvRo2e/bD+IL3/+RLxZallAesXoHRq/yrV5VsILqGzsNwvxNY
OUMpyfFvnPE+jl4v8b69o1HXKBJQ5zuQMDQLY8APt60URbd+wSGPW1c1xyrbNVtVAJthHG/wevFc
8xaSiIhUAzRaMS/Yw0RFJZd/AG0bhKy7eDIrR4lP/r3oUbdvoPR06b/XxuvuDrOTTzhFfRw5CvUJ
KEeHuiAxIvaj/LhQEzKtD1O8+UjcvLHrdzCjN3Y1giLJMzV16R+LY50G2veSJLbziG6cU1TjJD2q
pHC7kjV0SAyn28gYNJfbyag5D2VEPcynbBNlpENi9gKuySugs0RpOwgZXUp7AY8xHMRIjyPO0GvJ
bZAYWl+CbAc7FOWd5WKnVoKrjntZn9ltPZIY3yRsQs0botBHC0c0YUgJBcTmCaiUlCcljNF3f6Hd
YF3qnSGm4vGztXPLqi6orOknGfEqpI3wJUVdn8K+JQ7+tlgQ8UBk1ld90Pn8EFEj0uJLIP+RIwds
zlGihNjVZvyaKIQRjjOko0+b6hupMWu5mY45n5xOLtBeIXgGqMIBxgsJ8ECrZh82gh7tlgsi2meJ
vGF9iemt/IYjIwPVc9aneQKex4v8e7uYTON1oWUV0F6VL5TnH+fXiX5J/4x6rBokbxZPMF27RXTN
CwPZQtbF8NsPcyYnKVDonYCEeTze7njyYsNyGGyVu+pTg5vwgnHLzrjEdvQX8qpEk7py0FZtsV9U
qihYUyYINacajAQBE5KVVAGSfCAEW52VdgFPGlrq/PzQPR4Od9gj+09/Ea1SgsLVmV2LVAzGigmd
QDuo4VOdr8VBNz4Tgf64CZvKMI/qWzNj8Etj2iPZqOUwVyCeezhmnlWKyoR/+XaiXFvFnLxHxSNF
nAQv+5xQsVgK6K/VlG2/rQAdWvnoE4iTj/tVXNmLngYyZxNn0M7Pp0Ek96qVXrwUIY4ZkZucumf1
i69pAlMNmFp2523JGXKlpgm6aky6AWgybcNHftp6cggAx97DwkKqeagXBuRK+MsZoqwhH7+ZM+at
EiUsDETyf6fjSoFgPmyXrNQkTYCWlmzXVNj0n5DkX3MZN/8yuEkeIs3/LOQjN40BDwPmp8w2V+UB
oOtdDDsfIRMZMPgR/VwJw0cTIPIC3MEa/zYfffC9fRdpfqwYmESd5k6ImXygZtDAOCirNzUjcxCS
dS4hKeUzFkxeo2bHzKOCPkRKv4QQBKi77mdYLWGpuCXbO0IQ87kBHmoZ35V+zX4A+x5/yuL2H9kf
nHycrhVKF78KC6Qcrla+X7ZMW8QCG5EHJTmvBKicFPcpRxjCf7MmSZyfn7oO6RuOk/+Rpf44aVNl
EvEygol3H9Z4vJJkqvuFh9zsGqox4xRgcZsu6Z8iuerZz5wgWIZM4ZQWEhvkRVp0noXdvXYKOXzb
wVZxj80zomjJiR7H5eOunXxKgDDVXyHbPOz3ulLf9W+ptPEvPJCUL+sEk+EJtlytVxWMQTqLbpsD
Vwi0yxzqB9+Kb1r3NtoDucTZZX+gUvgQDMQXB2nUUFa6NtvsPH8bFFmsKloTYkCJPGqrSw7QENGJ
JFbglZSkPNT2guIaU8eUh4sjauC6jl2FLg8udDFxgOmvPozYDopkvDGrmq748C/3Yym76JMOfMv1
taPrShHFIufu7OOsJhmMzgJI2nS1r1MHBXr+74YANF1QJLPoRdBLMaFBrVy7QaUpDVzVd8ID54OX
s9K+WsI15i+5pfawCX8TRpPvKHiGg1AS+k6bXsQNrzkqWxTgwGmuAbGG5K9J7v08gb+dBzYujH6v
+cmfJx1Ecyg7j2amqh3EhJ3hGYic+ajqDq4zxkW+mEkiCv5lE2piuZyHFqa6ilB2ZwPWl0yBpOW1
s3aHabPjHNOyLwmEajho3xy8BMGRTAC7bx0POyAOoSSjrADX3VlSTzPYWm/jCjjpJhW0JLULUc63
b312h0Po2Hy3FCfqtKzLCJKNXi+et3jF+bXRGJahmR4HuJYMG11ly8kgWeG2gNZRFWuai61AIFN+
1PP2loGOLg3sxlwU1S1RyUbfs1CkH3+2ftc8bi6iPaBdEAhfr2mqhq1naaNlA8OMBIVaCgkguFhg
fIfcPohi4qw5Ooq1w1/lXEO4uH3wK+eSrg1XGt4I+xQ02Wl4/s4nqvqbpZQ2XLfodhB9INFUJxlX
MBFw7Kp7EH249HnsMYLo+t6T2ZTNJnOPtxIH6/p8oM/TBHjPBmm7fUZFD24zgSAJP6TQF5j10Eqa
NmjKdNOmyqTY7dd5HzG9KeYTfHL9JkxlV4p4pSjWR+4q5YQGnWuzUVEVzSR3oFkGRzCZQ7q+511D
PJXzJ4VSTjBkeLozlT/iQ6PzdCGFmJIR0VMc/cHG6nxR4B2aQwtuRT5Yq2DJpgVNkLjCBGCl+0ox
bUOFfefSYwhEUGH1Rm1ksBRy9j5kf+nkKYMasTOi4uve6vCdL9Swq2jNd++aTxcGHpc+Bxt2j0Kx
Ns0jfhXCy7bNYzeOw+BKFJ3rkq8xX9m0gBETXHlKbGRhHOUkh/PWZgrstCJDchiSNdzFneLOow+l
1wzqaKD2z0jeA7+ph6VwZcqdQcRLNJOqFC842QpPExc1i8/eFcizfAAylEfN6Tx/wCGfjhsah+Zc
Qtef87uS87v5VnZyUcp9UrF+60tgZgScCilIXx8KJN+QxmgQQ9MMOm7ePucmas0za6A/8kemr9Mo
zVVt7xwlqSwOTik3Zi/VQlzjfF0cDpl6EmPtgYSvD/Wek00dnVNXzXZ/InlgLkxZnvzWm8UKpBXy
L3AbkwweLVsZfsTUQ0UoATDOx7A4PlJOxx4XYKVu/yUhsTk3cc/6Y8VpiWBsPXybOaFZpSr3efqS
D5wDdp3X68nD1LiFbLH2hVR/QV2wzset9uu8vP17ivqTzQowjDo2CWVKw28ii5i+T/uYZ5B2kiIF
EbKVpr6hh7dUJdQP32tQcN49HSKr6MkVskdAMRYhhQCKf/tx0WCV95CLJDin7FwY7LjDO9v1RRVx
Slk+zcrmqq/d4nKWdarsF13UJ69tHn8FG9fQCsH7SYsMgKV+eBhmmzLWSDEK3a6NHF8TzpfeIBoy
+pBWEn6aqHUiTH9zOToh1YHpJanyh3uLQlyOxfLwwxE7bSwtqnC/o4YG4sSw/Pxl3hh/3yjy+kCE
lrK75BRkx1Xhi4exThICRdp4xi3OxtKmVlRzCCNtbwNF/yJ8XMM0tMhwQJV5QwKfY923Zgi7lvVt
6iWdpghqVJ/66Bsi77gISVajYo0PeWE9Fidr+GPNtztpcyFUUKOJRZ6NhZwq8RX8Vpb1fTlA7/x5
ehORD7AdrJDD5+KdKQG2q02AIMjCl6CBaJ1twEwXXj7Zp4SPisGkgQ8c4QQDpdD8c3Y/azm+kQov
3g27WleqYrucccDKm3yMzEKlrQ9GcSWMVNs5tFXk24CYCj5a3Kt3wvIxtEOo04BCA1hfEH+6oic+
dMTdI3yYK7bAdS7aTVagvgRcEm/RElyw3pELKppNLEihhI40BHR0jg1ifgeOX6mSqs1JznlTGyaW
wftRtDrKUmfzoL2I7fDWKf8zv2tQzpZjd3BbJp849MnmQnMYojZlfC8515IUnZSvtFCZ72pB3XPC
rrRhk8HR96JYD8QdgqV/2xqpY8h/SIsXvL8JpeHJuwgvFIQySnTeYWQvDFOFAck0pWzlGKZkPQUp
EZgQPANoNth+ITQBryDEaNF5m3yloUtgX8K1pCJWOP4ZzKl/ICUMk0E1rslquA0DpOgaOM6jJiqJ
wWd0w2bgKn2N2ubai0snHggotSgVollFVW7NxmTnkmR70qher6ooHK61yigFLu4nB56m5nBIitmS
BAfhk0fB0YYBEtf0SgvOYTa9rtxJsOLvSB/9Fn4Z4696iA7JahYdHjyi0PPCPeht9C0+lAGiirUv
YChGmZhDoStsbG4uMbBV49gjaO/fQKxTX8YaYwDXYdtd+ra9V0x16f0zdzF5r+mXaSLl9SMu6DJk
ifsEoHeI4pEGqDrGldBQlYxmAvA2wY6jzi5uP0rxpYvRSxLQfAtvKm9r9imlk1i2+0Sm5vKI6DqX
nIkB0Zqw8hRE+7GkQBptFCZQQSPNj/bmcL5Lg3nFrGSB39joVCuI265+lWhuIskGFeQvZMjGx4aS
X9TU3g61tol3qlvv6eNGrtHrRNd19cYLS2z69LkPb554DZedqzRPXcvxG2Plo6igco68dBFhqZI6
Na0d72OCd6X+bYAA2DZGYDipkzRDSzVk6bjS27KiWKtOZS32y1GzgQydSQ8kQM61pWpoiWgZ2ZaK
p4uQhc1cDQDLjdsoAolD2Gx3QhHHwwWkU9HU2EvXXvG/mzxqqILXkQP3/43SFR7UKST8PGB1D59m
qFQqCtO3CQxEMMid1c0qjNQlKdZKps+HftGhDmoY+Pkwq+QHUE3m9z0/uedWXRnb/5dY01KVFyse
JIiA62xa35zqEHy2hRkU3YMOv6bvogp1ni2aRS35BBBBRS+1SzYLT/dNq+Nj9+uZ+iv0FgGLRU6s
bArwzOyJPU2jVNv7YQhYxcgboUuaWWHkkP5AblSw/zKZscdHnNA7nI2U8YYqrRO/ggoLpHzO5w3B
ftLcjwl9glAmSvcginhP5zPtD70uwzpOvg6KUyNN1Q4AGzGztxAP9Qg6VyaOu/JIvJu+0Y5DOwHJ
3CDfs/9ZvbVejH25PFf3BS7Zie0IQux73mFq83GZ+e+bE4gXUInbLxph05iRFYo4cNmRoJu/ZMTy
6DBffIRoU1C8waiRsEqAsXzx5pwxnR9HuTYFBg6VflRCCiQ+tr79nwGbZw/MM0OqPS5nMpzOAz3l
P5t18Uiri1kuiPASk/3862Aey4QA/seEwzu1pXnvnjLCkjuNm1uWDML3AZhF7JW6FEd/I+1AJVEH
Ydw/GAVSWclE4xPeytG3vi8QgU5pqQbeBRJB+XdJ5825yjJFfrvxKBHrnoyruHu4Q5xPNcCfNJtg
FBvAgnsx7aX1o4qEvaTM2nrlJjER+aFiZbdWjlECFClUwMEUu0ArxyK8xIPx6X8uzhxo4txNwJMO
DrvE3aJw9djZ2bPh/5eZHoir3DAqCVarL8UmRGUQeL4VJMWjHcU+0A/ScIMlHmXcw2JDIpgx6qxb
RJx2weW5pbJu15OCUBKew6QYST/TT34zOwi2LXtJEYMmiBua1eazBC36najez/6BpsQpSAgL+Lu0
YwpkAi4VHdfhkPpToiS62xjpBfQK2xyXllq3txDQfqpYYQ0QSdN4rX/zxSb937UC/ig1vo4cDvze
V/KNbVqRqC1hYxKu6KYhaGKAgB3ynRXCPL72KY2lWpzt+G5qF4F8HDBkoL4bH0IfDJkJYPLXYjw3
wBbmAaYTQQCm8smhgUxMWqkQx1GT4u0ozmJJEQ/bArUXn7Sos7e5W8YZ2cUSVlf5w/u0W5hf1WGn
lMrNjNLaZwO3aFABRwSij5oc2yBaYVOZyFVq/Tbv3ngLBZt+hhBwlEMcrOnFbTxluLeQNpxCLEto
yC4S5+wQRLXqk+z/kqHaJdnlg4ytm/yDrGwkWBXU3DJiP+0OVh/jJa6ykPAWvZXTdSvjADMmORyV
yLl2wC4QMMqAsE995XeuzUDt3SFMxSFwNeAx1FJCDidA/8pN4vUoZpW96j8EmMNEY9o0PP8BUeOh
PU3VQawgGS+p24gLExu7HALUUjU7GXBiGWPdcG7YFX4y2yA+/oIyghUFc4hraSd0t9cJdyyUgcMO
cluq6Z3FDx7y0gGnAs5Dz3UmNYv248cqlNo4iZTBFFlYPN63cdbBA+r0A5x5Kx4wPfnl9r1ZMVx5
9oKEo6ZbH+FnB7y+er/vBZXJOuAvdadIgVi0E9if/51/3Vw5k5qNK0y65IuXVllGxNslJASGVXvV
8No1aHGfsvOfg0eL4B/gxafDEbAg5mnRPKz+KvEBSUNlfyBPcJPkJ1Z4FAw8+ZelgRQKf0yOZnEL
IDyhRdtOC5ywDWMzSSbS583vxNawu8+NehbLfoK1t1aMSPUdR+EBgJu4+SCAkh07vomvotBc1qFC
COiRCe6xl3jAbVoO8N2pKJbx24yP6jnAUm6ioC1ThP/EfkaL6K51keKD07vx7k7goZGxfp+4ZwIc
O5lKpVJVGwQEcRlu3r+dSoEE4DY1TZ8+NfbzLkoO05n1K4t2x3mcEIfEfZqfjDJXhKxM+9hr31yO
KxD1PDd9ccUWK1ZYCG6uwOF62ePF/8jAfGFvWEMtluPOErVJfiP+G0Gh4ujGc1P8hzF3xuerQiGp
uDI8NTnrxUE+DjOip/JLrTls1zEbUn35JrwXmzGq/88b+27qHtKC1AbaCV5ioSjhqTzEC0scFshV
WhVtBAB+XzA283eDekK+tI4K7rpWbkk6adFFQzeR8aTYkPBqRlpDDHWolMnhcE748shRcAQs+dh2
Qa4fLT7XoFV5yCMiCC8IZFc2Xi+X2aXHcC4JyZl+Oz2tHeJihN58TJ48fppK8oFJDs/hXat4bknv
w51nj9iK0QIBGVIHk8DPPFkqOLCqtusTNO1s0B2jD2QplpaRlEeC3menk9SYiEZVXotvaFyNCjmh
7sJi1LV4OCC83eCgsen2a2Fzc52rhxFctx3oa+sbeYZSvwDxShwfwaB+bY3W1gx6FaT+xluhOEkJ
ksZGwBBQbuNArpRpzZy9uTRzo6xxfiRPQDsPeBVZNrzDdYnpt7nH3sxoQik3eCXmXrGE+jiuZZIo
0PWz4YrFJabrCbYkRdjYNj5dHs879vxaayICttnu/jgbx0fKmUHLlqw55o8hNGwqb1P70DI435Lo
+p3GcaYnhcuN34HqFgbW3fLqcC1mDUK7K53PORFX61Oshjjmz6dpSiRR6bqcSh2Y65gPBWAE/XLP
bTW7hu2rAgclYrkUE8QCPthTYdMaaSfJbHSa/OO9NodMhcySHnnbCRxfiTMY9WrAWOO+npjaiNzo
L6tYBoh8FGTwKah4JiBdhDjxM+Nw5WSIoLD1heVdRBU3iEgVLN7tqW1gXnVecDK9g/wSB2aYTpPM
GmNKCnx4MSOBVoHlp05h4O4eNdpN2nwCOF1Fmy5krOj6tsYbR7wvF0UBuEo6/QwNR6P3oHxCqvTA
Uyewt/yxYDaoWigFBp9jddrnoJzQ5knjTsZiLMlqbTu04MxgIHN8qQC4iSg6+7BpTefEHobk/zsw
3WUCwfp6Y8Ga9t33uOdv4Y1LJIoCoYeGHCwCE4ukmqShx2mpR3dM0mFN6OmOvYwkhoKTLX9s4AZ/
5V+KJa/IATvW32KD9QHTf0ZCKxYAmzQgngKR2ja5kJ5kzNeKXw4vQVIOZK2T+OchCOIkY+hxr0Ep
4wVIpTvX1fCsMdfEPRM/QlB7bfJs2470Nelm4xsYahn5Xt+g+UUGJAJi7E26UJqU7qZqJANAZ6vq
kcDD+49h5fSr3vfSMsL5SbY7hq0HoguF5HnsNrwyShzuw53dxg4F848GN5aGoADiqlXDC3EluLgk
1Exnw3v3R+tFGZkCkRB4HWUMOlWIIQ3H9NwbSmT6M/JJh8HQ6bnDLsGpWbv4XPGLMD/Nac+H5bJJ
KZXzkIAhWiPMubnk6oYhFuveHI2GVmA/vC0J089r271x++hhy+1U/Rjnx8i2QQSK1ADIu4aHQ2Ih
69BzRMjSQYgEngVSIMGY+Z/XAw/DtJPa6VTs6eBH/I90Rpv7H3EzThzo+tDSIL7U8hwDnEwoiLkQ
OuhDEcEX8LdZgkZ3al+9uEn6IqnpjUo2BPj0dm8INDRKCdfmSPXl5sTFpnntE0tJlLXxRaMzqZim
PbC8nH0cFkri6A5BzjJVJ1ONV00U9ZgpoyDvHWjpVUrrTdEvPeqaEYUCKp9tb6+XtL1ZATMH/uLf
jVMvdsa6+5Mrp67qhPAmjI6/0rQeA8exxvYICN+8gafNp2Wm5Yz78xdFaCRGHsL3Voz8Nn13n1uB
dwNHxCD4LSCdJaDR9O0EavI2YzXDCl6gJf13TAotbrQ5p8e33KfdKBEodnLTKyGQuD9di4fvDNs5
bh9jDk7I6z52mqAVtdbK8whCwz77UQ77u4eXJdX6EUzhaG+mZpnYPtij3/V0uBPCOVSh3tREV/sr
e2dZfhbOb7KDsOUSbSprOUX6qNcyTjgTRp5bF8JoFAR+ks/zAMq/jSVILaipzIHkWe+IQvzNFs/g
gPMPxnh1iBWvTthIn6kTn6bNHv+UkCS1tO2AOXzQ5OOF77yFdtsoARAJTJA6RMllvl/sCA5J/uPs
QwrlezldfVZzL/DVTI1U+TEyYPI3Z05AFr1E9rRLd1HTLsXCc48fyJAfzQh+x2ScrwDTW03KegC4
mekdc1CmeCf2Wsp0v3HeQGqUYvL3NdfxRepjxto8cdPtcz1o58cKy9cXMtcoyhk3HRnN8CNFW6j/
2L8hgLMlCulZh1a1XTHq1iaEHJfUWltRcXA2qOmwdjGl62c1qpFIqC4CkFEKT+OUQy0LXoCwm785
d0KVeHqjDUfcHVCCKxDwnXgpMItPXkqZ60wm/vDvZc4tuhZOr5O3kZxx6R1NthxfUYGXUrpnEbCT
ZPbz6wEZ13eV8hte3gOCKEclPtLzZz5cEZ4gQ5v6r25NlcYQ+xcfxoB9jVhALvPjhP8KJBFLmBmQ
nEYNmzMc6pW5JbXxmzUbEfx9seZhG3NDSoLzXzfGS3rcQ1S/SBpW6PNIjf6qqOpskj/MKDJ7M2SP
wjCXpoX6GAeizRYhSkOW/uK6HVPoF0G4JiFv5vxiz5p6XyKJdeNiHezceNx11IZIXHhqHOx/f/yN
TaMBiJ1DFjWz0EOFYalQmUonxJzWJPRmh3iSS+0rQJq8ES3LxlmlvTfE4k2erLXwamTmNVNeUa8t
V7cwWn47hTCEHP602PJuhQCy/q5JKJXCnNfzaX+IEKV7XqUdwiMC9z5Gmb1gOWCenuten8nu6Jr+
hDmpVuDvIorWL+Jf3bUfGG8FzUj3/WWq4SHnrC/S7jk3nXOS+XkOCcf/LsJku+LUh/+4b9uecV8t
NDomh1vvQnpfwwjIZZb3fK8xoc5ptGClUY9vyltOUh/rcYYsgSwX+oWazxURJdFvnEgl1iqqOmx8
IkiCGh6jIb5M3fbKGpLj7Ehf+m1rRqNzQ0XomSaOdjbYO/twwRPzkoQ2smEgA+E+YVGHaTE44FAz
q+TzILJJ9vn+CP3Z2eeGHPbwDmBl7whvzoc8DFmpVnIfz86LjnELTF6HfYfp/4AK3MrgUArGccGC
+7QtpYAy/NdUvw32X3LUJXo1T3JF6BG3WAl/5jgg/8l3KTH97eFb479WBJ/ENPGC06iJ98wUWub5
Javxrup4TC0h5141g79+/5k5b906ouvjyyXzKAZY7H7C3n4CmI6px8Sz8nMeVDF6zO54Uv6HAXoc
WzZKkqyTQGP7ovJcnA5Vfs762EmG9Qo/7JYhXuxN11/Agu+sSYmG0J94Ry8VoETNlmZL5boc4/IE
9uKx+nKqh1vWPtOjYO7pLV4nc+7nGMzjswhpz0pwu05QfcWJ0UaTszysiJ2ArqiDhAyUkhxi4uUU
BaVsIkCVmnWZjR5s6+fuPAd9xwDRVVwxCeTycxk0xKQYqJgHrLUG1aSW1/5BthGIhDIFHAlyU61V
zKXD3X/Jk+phQh3sAG5h1g//A0ry0OF7IkqRwIf3hU29bBtMhBUM79b4ofSArKMHqR0xLdO1qzv8
IxmqwsM4hNmifx8sq35pt7BsmLzg+wv8y8O6eKtsv6N9FF1C/x1aPTeAwu/tfTXzG72czUmI7yWq
ieZJUiHxNBXbbHhQNzHjsZ4hV5OLGgzCCCnsvDK35BjmyNJediMJddOvenHRKH+60LNGL34MRHK4
2QzNj4crYiNJYKcUmSozjW1U1KbtMWnzyHKkDZdO0gokYWSCptZJDQju894vveMDPl6OWsRiLi6Z
vBApaXebToqCV76v2SBuMePYo23hEVYBkTL4NhT5jFmuUcQbQtL1uVyDUHTfPpo3zDF6q9FwsAH4
Fzck3QlJNfzSRJM37Qoangbw+bpphuUuGr1/0r36wn5Hi4CpJaR7ak4rQRYtv8cm2iSfm/iDaDFR
ClYVQFBq0wz/Ea3LzNyQHDc0fSvJlUiZDuT22M/+V6hIpmK6i7YlMSRTzAoNan6Wbv7gEzZVgLVa
jnsdU8bbhFJ9rKlWZIF3dtCNpoAu12CytjnCSdKM2tf3olYHKEcj0Rq0xbLaVevDcUnNsTQUP6Ba
flYcaEHiquXznr5wScf3nVP60L++RJHQjJPsUzDOetIemM6stM2bl8eshT/4kpVrT5A81AQZpige
Ccj3dYd9RXms6Dahqkv9diuDNEZjj9zMEg1EnUcTg5aHoOcHvPBWAAEGb7EGeVDbUfA+8HZVbABi
a7ED9qRBzHQbrqR1wJzSl4V5yQJXMX7HEFYu48CnME11rNLRoysr2Xv5dkhixl5fQn1CYIP4dZ9x
IjDehxPTG1T504olseSKHfrSWG/kXMxbZztF2Vg8PM+KX21FrGnBeZiNnCDkN6Fb84FKjrDHhhcm
dqFvgg8vO1/+l2lbQvDoM0b2nT4aN2jZzkWf49Z+uw5V7OuOOPCfZNeFkL3n7RfCtc6k6v5/FG0d
VFrNT629DkS0FxudhEIxNa14SewP31Sq/ZlM0+9+6EylXTZEDsJ0/FiuuON8/L1tPCa5K6rOxpp1
wWsTYbR8u6/YZChEZ8SIaIs/IR8JuuXfOqMyMmin3DfUF0GeGKfh3UoaLDPMCqEAe9CtltYp7HDk
uXYh52qA96NiM//YBVcDbZhgrNx/irX5aOKCpRXHLwZHq4rSL6F9bdFQA83raAbobYBVQqwY5hNw
hbxem7dmHBQKHw0n3CPJiWFwKXG/zfNho7yMAsg5PeCIsT1gk/9XuLKfSTRoz2ycDY/q3N/I+lao
+syNetMuJeAeMHUq7YKjyR28adzJy2GZABhBth+oL0xr+Dg5mt4lQAbfPOqsx0PUM//Y3UkVjGWY
jfK5YTj1pY2760zBuTbQzcLvL2l9pBxYuxxVNTCF1guVe32sMBG1Hvr3f71TGkJgzS6y476bDMia
uxellpk1E8N1RntuIwukE8l5/fO07ebvIueN54Lqx8FtqkhALdWbUdlu27VoxzJGGiWKJGYCL8EZ
m1OwpwOXmoS/EY1FnQaLAxr0mBfSaTYk+l0vqIav6TjGnt14VCR+Jz69BOzWJxHvWI/HQ4LAlS0+
VGdbzA+/++usCpcgCGxfM4vTe4/yuKfpizsxFHcqQco2L/Co/07O1wUSNamsEDOhaRxiEogfwZjo
P5N5WxzAxXdQJ6ytIGi2z7W561u6LtUS7QP+/q0JBYYep89EmGbx/RiWJEkintqR9XSlrcHTSMLQ
DdLQsH+scLRmVgsZna+yRalM7lBPf0MrRnWSp19Bi9zLM7O7b5iSj+zee4TnPXpbkmoOXUxTM5F2
Arvx38CgtBZZmko0QMkVQPk9U1UCGkj4fbJY2OFLQrZFirNeioUY77NhG4z7i+wmrI0MWX61rIKi
O+fkNqI1jR0p2UFl/hykZZVRcq/+HdJewJ08h+SB2NilIrGOD08Vstr3e0XCkRyfFC5n+yTdPxxu
vsrKpF036BbQIy7H+3u9NhfWlqypNVdgv2hkbFx6qwKm0lr/Irbxx0ATuC3hzAEwrvE0hbK/PjN4
7cup+QCpoZVgmIYNyjjFqiuq3XgdwVml5B4nTC3gv7grVWWRGrE0uTlOn8q9wWhAL5NidLF4i1RK
77AnIBtxpTbHpo9yjD3jNCmZVWZwjWtc1dyCXZx7kJUC8x5p2kjNf1JN8NuML/mB7VeJlNk7wxvo
wMffGQgklewu8NTIGmFyXdLKnZptB5l3zDsFiGoshRKEyfUe8CAB/uOYlpeU8ni8sXVpf5GKbkxQ
Xl7uI2LP0rcIswYlpdjl1WYm98i5lrEjH6Wue9oVMtGiciXvybEXy6P4i/iu7PWEL/GRRWMOMez1
SVVIYNw47Gt3h03gCzFXteWeqEmCUx5Jz5mRvihmzseEwfPnhgBp9hIkK9myDVBV9Pv7T5k9XJWk
FzU+HyaVkSFjPZg4O7SW5j6O4JV8viHBSAO8AYNIN8YXl7AkN/Wvy/FZqoUjWqjjU/BGqS4ucwuA
5iEWNlKXGbTZHqCE5lVTgVVlyEdWP88UHpz9rg6qujmoP8+X+0EBe4Q+hZqndRgOpgnY2lTwH1aC
5Db/dBnafLOm30IPSr+SA/h9R9caI4b4CxoIFsh7gyJNq2nsqX+gFfYKzI7npO6wz5xO+YEgW06s
BZT9X2+ScevhbHOFNpUJars51ZInEKtbRgIP/vIF/8WF1XtpBtUSboiECvIxerCIvQ80HTv0+gt8
wNGELZrAVPz+ORUb4roiSEKBv85qYBw6MN9C5SUXSng8DMuN8DAOlYshATEKsXKdYEz3P0B3fshO
nVq3tzIlVPodxjWmNpZdyXr1X7POxdrMQB4rvP3kmu+0EXspUf4y0SH8rSEUkozppwp6UsF52t1U
7T45vrokHpnQ+lxLqVlwG6b2CZnilSygaYcwgsJI7uvPhUEdJIOKTAW2ospcMmW2ufD26QICFd/x
NGkFVmO5SR35FkqWhNk8b0QFtmw6n6LXqnqlZwKrVXEW+MlpLk1T8syjmjpz37/sTS6HtjfpznlS
N+oEHyfx12b3AQoAOM1FMD5n+MkRaFD68WYVd2OmBPeNNznG88fySSMBM0wld2Twps1tft8sxAZC
MWiXIIDqyHbviOPb+ojrb0Kh9eL9RZODuulPA+j9x4FJo1eXkPE+UsxliTFnX/a75GnL0vcFDTpO
pQ4KVEjt4bjKyVBIeFcrB5G+Hh/iR39Bwr/Nq4kz8ujkYE0MbNVG0dJ5HWLiwAjYLrLWQe3Q2KJJ
q4BMNKs/1BD8SfWb1EPEMQsB9t2JRzwrf5sxMgGEJGm/yY2zTTEAHchnnLdKlgSWC3B8FWBIje2R
abC7krQeAUW+iU8BBcCKGH/k28DXlasgCNRmyDANtrMslTaTREsXNrfEcITRVgYLJ+x1bmH/IwHz
05y2NQQ/q2fdt83e2hAns/lP83tR3HUP9ssK1LMCrM4hU6boUXxqZZLyVvGlk9hApitw+V6jQk0A
m0J7Pkn5ZDp4O+cSNGDpNEvzBDUUZHQwsh7dN0o4cGAi70o9pJJuwkGQ+WTosscD12kRap7K+sFy
yydAlnGGJ8yYrz5O0+krP0twJLfQ2PdaK3a3Nuu8f8M2R2H1DxtF7st3/dIRUUP1T0VqfSjhGbzq
SEttoXUA4Be/ic79W+0FXqveNqVbxYokUmTaJsaHmsJSnQWrnSzq3j/C4voncuKm8wA3xhzMQ95s
x1izwD+qWpVavgujbiU37VAztlBiMwLz07kgddjZRPX9hTKg3z4cmU5pG7XlBLo3n0tUon0dwSEm
Ez0FuhwCNCuOcxdcmuAy9fmulwxX2ga10tv4gbaWvAgyqlSq7yzaSxVpQGx07dnLvbwXzob9qKOa
6awcyS5CGIrdLwudjYOAhptRzvZ3HG1y/rxOOGmcT2pX9uRAld6G613ITo8intEtuMXyMg1VU8Jw
A1u3H0gNQVjHDT9MnrTRI+dCQ8Oj568jM2rw9tmKYH5GSdkXR1UBXjenogpm+Ehiq+DNrhvk+Gl8
7kVjPTaqM8ZZsKhF+vnl0wtmxe/ZXtF0mnYClNzBSQW+TuYEjSKku3RoU9WAvOLD9uc8nPOcmlPf
80RzD12QPyB9w3tqnJ6yWsQClGkXMtMs/tKlwJ56CHYeJIkcRRNqb/nbaShBVjING/qIIVQtOXaL
aChKS0uvRPNjeLBNjNrQxIDEOkZHGCYunZp0Auu9jmEO63QD/vizJQ5BTKBkEklUrwx1P0OefkdG
pCk7q21InrMviFXS7kIxc/zOBBiDAoylCTOME428ucDApmFXfoU3tUEf92PDT+tD8IjU8VzbEfzE
UL6K7rJZJj5/h4oYVYy2sPQ+sMx4oB5qX99I8i9fbBp38TZbkh7pb6pt4i/rde4d4dBIwN5ucAbX
u3LNWoOxbSlgeT26b5CkKA+H0YKH8PjPbvWGYzqcg/XmV/ULTX1IV+OD9BIsrsoD1Wn4Z5TJm9ZA
XNl4x+ScUz23UXOOcIoCeEH1QdMvkU8myTshZVtKRDCySrx23i47JmroNH8eYXeNC1uchQdIcgvw
uSpcyKBJS2p+e73QnhV6Hro7xTinKVDvWiUQnZ5Xnwy7fhMMjxfWX98cRxq2TG1dkucXvp5gl8nD
seHr8Vvc/8zZkU8Kc0N57BpMaAgrTCHhbuncZK7RfXlpQ1TkQ1vOX5aWc7Ojp2Ihdl6wqmu++RIJ
b546eVXzl6EHrO5z1/JsanCE8iVW6KLm7780zWXOb+G0ZwtU5qw8Nw25nBA1+pbiVVxZ9jtu9ba8
w5Wte82ap4W/gWDr97vNJ78BaufWpkS+Jd02gxjtXwV70kbUzOhCSgqIJFBCqGKt5LfXSvhkg3pf
1CKui7uRqk+avAdrTpmIMDus17slk9zjV+E3tZ+zDQOIY/2rZDdaUPISvkEf5SMvliMx2yHnS+Ui
VPilBQZ8p/rp+1HOl1Gb4A8ostdKXirrFzMLmFTWupxECghvuDoozvbwNU67/hureYAFONQ71/sV
kmXHwuOhBRuwyNwBLD1mB1kfOrcm2a2KYZEUAuUv0GMtl1lRsvgSMl5vDOgjg9Gkkgk5lOPSawlU
9kZQoPMtsAN0XSc2uu6/OjUtOALNvzCSqosgxUxyQovFbXwrSpb2lTjSsRoqTolOuuwZPlKRIZyo
7UUj7skOiE+PJclm+l2S2ArBdPvkHOCB9hErgKR0yzdsvKUcVd5gBNFkwjfLs+JvlQjKuefqtstG
LJlKdp4lD15hX0aS9vqFaIuaJh/lMSQfVi+X2+GKNIZ3avKTiIAMvx+Rlna/uoYciV2PD1dWM+/Y
emxOGgj/YjownbzKCfspbOTKB7uAZPu5cV7FLKCG4u5cw8UaRJRDrvUmHwD+KXqZIE3tLohWorTp
dr1oCDp6cZekpEhodDDixfLC+qLX9VeSi9RWBLf5iHVNWCCqZKdeXkdDae36MqOrpY4HKsQ+tOv1
oVpst0Ivpo11uwB7kxn7lzYwAP2WWBPgLIGkSE/cPiUvvpd/GDCUsXwyFKHwbybcz8SxoE1gP1me
QdQpuUYxGCNdJLhp0QzettLyQtqWcGN23lQ7Jqd8pxYWbcQ3LnB9ZBhYOdL3Fc0BrF/9Ame0O/28
tXbbuDXC2iyIFOinzwMnSV9bbxs8XRIiqhZ9MYUPLw8s58NKdf9t28PsuNGkT8kablkU0gw58tK7
atO3Kx2MWTAI8SJc9ZtRsETLxIWF4Fkx853lJfwI6zQ6oe8ycLr7t2ZKCKgnxuSnvudtHRCfoVPB
A63YaZNJ0nUDCiCW5+3wa9Yjm8FopeDAugBzFd9IsRD67E999ux63H3xHpl9HyGkEYAtTl5BDF7h
yndSUnZ0IpDYB7ZeY3AfYJ2LD3SEY842uOfR4tGORQ1NDyc8RSeFaz1u9XWuWjXI5oHpY5Gggeka
2ysIdIg+KGrfH0NTK6Tvc4pNzW5SXiyb/Hy/t093lNCd+ozhlXKtik7pAKEZ3wu2AaU1yUouX3H3
88V7fsGkHNJOdDFLCJDmwBeW0pw8/I7lgCtsDAhSyzITtOeh0KIU6MIgrlEYdggJOdGQchRl91C+
+CilnLkN+eLY6qGI7mZRmVxgTfclKN9ALhWmYaZhDGRWcKik6FqAfoitVn+xmPKoE9iBZsky8jbe
RD44Ql84DA8qClps6/DeYXwU4vIaP+SnHf0jQw8x13dJBC7wJgSeXqSF0fcJnl6IeG6+5s2jVQyP
EEIzoX9XSOkI5nDVkndEzdV9lvqUd6oBPTF6qHWj+FRGSp0HgSLMq/lDKDPHMCyphGOzXcZFsDbO
29SLW4g0KFR4x5ZuKoaNnlb7srTlgeOXOU+7RWpgFxc1+M5CEyrf9VQFVi8BkaainhF7UOML6cRG
9cZ47UGGS3forTtaYBUlhQVe1bEPyni8h5xtBCCBoKPYWLHNr9yU7rf2abNDibUsOEMtVH5YtX2y
HYfqSrV2ue7bgaawCfIzk4AGP0uGPuKArStOM3F4O2bSbGujuGNGmEwz+xa7Zg5G4OLBzvthg4vE
uHUnBMwsSeJlrnwlzC+j8bWp4am6nzDPLctMjkw+mZaIBH0c+pE+Wn9i60seah7v/zm6We4Ncu2V
dsDT9eTv419AuZlXhyFhNxhBZQePh6+/RNRCFoV6Qer7YNwDtZoxI0Yj3L4TULeyBa5bktY1VZs5
rQ+2Ve4RA0MExZ6CFMHj7gE1Bwf4K5b6/57U88xadsTcxWtQKOYrDocpC+FGik/AOx9VEoI1sINE
BOY/WgVa7oQKVDCaaWmLnpxxYHIb01OOB6D8EDn3/e61p35RckMbB/0jeAYgnCfoXdqngj1UOvVl
FYIFw9/adrsGJ+r7NxKRB6j2Q0lVmB+6DaWcU4WbHzT+7PMrQACYfFyK4ic0ShzuagLMbmhALPFH
nB1tW6jX8OcogNim6zNzI6CMqfsjh47k3kRz9bavh+eJNLBUGXlrVsqQawy7ZHLOvD3a26J6XOsj
EnXj9IfrGTTOgO6A6VfD7a8r1podqAlwMCKjQr9aJ/cyPLKdfHOSqktAhOthK7wYrmlBhvT/mBbf
fubQKD0yHnLREnsRerE4Qx+D05WGgGC1WndmfxryoEyEfS9cYC1Fr5wre5edpsdhMWg//Sbx0KND
RCDiHAj7mpGcm51yXRkBYANyvNrHm0oM9jzXoXSt9dCQ6VjFgNgGvz3S7aiWZcwMBmJQsnL++NDX
IcUWVvI/bUd5ATYChczDUuyfga8VF3te6MW5LUZt/9EQu+y0VmKm0k2j1XQfgXi7BwpaGFGpHsQ7
vEVi9rGls+wZ2GY60cZWFfjQ/sbFbDZ58fgTegG6+WaOVOlBMU6GAaeZyp6xiAt2LXZOaQk+QyQp
REA3A2ToiEbtvONyF7rnXpUGa94kNmj7z0LhFk9bOSodBtPP79XvNtCLgM6bVV9CKSw0VobIps/k
Y4rSEKOdx5ufHte6Errk/pPeQAE852PeGt7x9gvAeHZ/OzehZgldb5kLXndlJThXdh/vG330XbNX
1b4OEWOu4XjiFbeIcTTU3d5E4b5msitOii2X9igJLyYGYFDAivXjjl/Dr//zg27ePSyb+z16AAHe
Eul1dj/4lt9XOi8BmjT/zlwd7FAa9igNErrbQaYV8vXbgY5sTq6xHTyniEkcCB9M9kqV5evnd/0f
s8ovND/Ppr+DtEALRNedvUfQVrPDFYHwvC62+dV4NB51FwFe/0KN3jbzfKF4Tdb83rdYZqfahXKP
f+sbahFKy5sYJykJn+CcmvNufhAx09Lqp6SzYmI5AqdsZwnq5ClVq46+fQ0ye3gZyUkQMUG0CKMW
4QCE0wJQ1jj4lO3GgiBVt6bqrhBc+/a20rdxIB9McK5DkG5YJvnp0aCYAuhn5pDdP42ewLXuPahl
QYW9g5DynwcJe00/4mfCoTrML7+Qi2gMFLwRFnA3rd4Z0huVoZ/BHA29U6pv2NJKohKOP7v6n8Dl
+QIBBEwduoIlbw28DEn1C7HizEPP+rCsQrk4oqONLNxT3zZAKVyhdZ0mD0CzU9EoERllF1mctCWQ
1+pLYsS7rzn+i1RulwLbul4ruirXDbjoR4Yg6z96DkgMEmchpKhbRN5QhSzvCSHUxQfigJM5oHgm
1aeRsG+yeJ/awiKeDSxEWVx85F2+LuvtkN2MIAUdcgBkQ7LI6bbMY/fdTttklDsBQQ8R6VBRFj+p
VNsBInMcW6EJnE7hYTyih21lsughz02gYl2FoE7vIggj3W+uPztxwUMZhp62W9Oi/vbrD5HUmzby
zIK8vWNH2ME5yl/mZXhlb21rcAA2G82mNscg85UEP0yZNHUh3ehiGZ/8NkY4rmCZXuVoGu4Vfbfv
LBvOuLvPXPLKeYlOaohrdlsuSZuqqxN0qUc6m8FdNL8fCl11j5sbQQuyVTzjgfqYl9130Y7gK3nu
htasfr036kSnx0hbnUK6fm/GHpl74SrljiKF+ynQ5iO0WnZ2BXupHdsu+Mb/4Npv0PjujKR0SJop
RFarqEVlGRY2XSqfiyqEoKlNlP6ZkmGqz66W2YZfIDMo/GN8p6aQaCKMPH6ILz7/knFTsiH5vu9N
MHUTdLv/yXJywUI6VYBgagaxZOnmn6O8Hzd0PVKS3dZHIqTLREDDYcpljFYF4QcpxASFyVy7l5it
yZ6BsrL1Zaptm9N/GfH+zgrzEsS6ye9W6iPuKie8tbQm3LYxJ7h5Q5P1gscniHggtzwUD4ImC+bf
ArbBs4rG0v0/Un6lUZN+1nllZw9gVcU9yuUcUFfkNdhaUAoljK/4HrkgVBut6OWJO2i/6cJGloV9
6i2LapNBrxjBN2J+gSR/YtzydoBwM43tGfO5zPRqDpQu30Tgu9FUyjOobstLMtirQ3At1qbJ6+4Y
daA0/E7MztZldHz50flunNL3t0JuYJja1zRx2H6dwWwDCjr0sEIw1XW/9XVXkk84WCltKEwlcCZp
XnyTZribZluhPcp91f0iG5UXZbcl6zfwDx51SFKRxxo4rbbtRxSf4IVgtX7AGUt4sQndhfGZ8Dlt
aut5CNLSqX3h+b3pGfkZnNvxD1bQo5fZy0EupuY2C1WFMDmfVq9vHmndgWu6Q1ZJe3dAqAyr7/9G
T9rM9sCG3j19yEKtFlkl7tLOT1ctmg7amYTJbtynvjPsLDuI5QwjVxmnaRPhgmoRZSegqKGioNK1
DQBVDo5+2CFAY3hykHIDWYON6svnjZbKWiTzYPLXXoZdxV8ytXxenE9MMU/FsrFQaE/xqrOjVT0A
kG8MK5ShCPl7x96vgcuaz/qtGoW34vTm3tB2dWUcxOvP+rdgzEVZ7GlV4tz3yzjiDK1s79CYJmtp
Qi5bBBp1O/THCr4cOJDMAB3XEyUXdAFiYPyeaiRiWkF0aV7bhsgK8fVLwyLWy33CmWzq2vBd8OyU
CwCOk8PX5k/glvYUYSQk2VpDvigh9+m/zG0Ay9vV34urgZsvneWZUOW9Yi1v8yjqrY8672GXpBxW
9BdwpAEp8IhPJFMEHrpiPqhrzH5MbPFdfvOnLcXy28G05X49IBeKztKHtOj1pEokJsIZuMwfNhDa
rEieChcrwgm2QXLngUSAR2gua9RnqXrkJRoJonfdocAAnuSF+Q18DjJc/4cW6a8GSKjZnkjhUUx2
/tEoQm32LeIVpbtPv+5pOyU1OsZR9TkOjuBhFF7s3rW7DQkRXNXMgsyD2X+tJGnR11h3QuOqBf54
6Dsf/cFn4z/41aeP1yGoFF7e1V/XTiAMJ5A4SxKyw5qrlzbM053S7EFrScFgZpdaXRw4f3H0+IlC
DzoaGq3B90bNCd4gDnNc/mvWOB+WC1eyPACCXckT59RrvRaxcacrLz04nKOR9GGsD3SC4t20kfBR
8sHOnLIdLbJDBA9191YC0sd96uxponiFW1UI31q8iy8HKP+gg+5f3ZPbizFwxXsjr1XXojO0m9Fp
hUevSlM1BMIoRNNbo4Q97SjP9N5gQFOmfMRTgVPDkJdGdGuTJOUxNfCCzv3rk7psKRMw5RtbcIOk
t4XHOgluXbdNmFnWRZncLg6DJLEwoSAbwPAAi6eaCYSTJe9W66uqHjUDNYNK71+x1zmG7VvgECMd
+vHlYduD9GZVdCjmkiNe+y5XOMITei/FY95cUNm80W3GPtp76FAAseI28GS3kW6fqvB+PNnY9zid
rNmn/L1LyyGxbY7WjJrI/FynmmgpzIK98+DXWyKK8HzEiLtcl4f2tSeCn33oOcP0agEoeLEm9Jsz
qiNrf3uMcRugwCtWse0d10ujHDCU0QXzw7/O62f8/ZQVjk3XOxuEl2+nX6AOE1QjQWVBT6uRo8OS
awaLB4BuZJUGMBwhAYFn76OYMLpTLQgt5grxO4fbjZc4CG1VU2A88n1DHdNApdGiLE7p8PzvjvSq
NPNxZdog0RfEav7lxrgH5XXVLuPK/EB3qzT+35M6RAG3IlbpePZDiE+1AbS8TQ9l0FzHoql6VJIs
6+XlXZSBHT1DB5cfwNi+aaOe9xrfHrCz7T856kLsEOi+LX/2NfMJENZmzxt4/idL0MGfnVWuKQHR
Siw80szRgpVdqV0KR09y4rnfN0OjxYAko2A05O91jEESzbXbtLsmXNZrRQlFa6Ezge5MMwXsgAMk
+5rKwANY5mQ660AtJQQXndkhn/mGNTNcW0R2FbuaLh/n1rdyRwoxyrqf/TurymlPIHNQoE7gVgqk
LttCTVm5xzk/6uV3z6ZHz4MtQE/riCX2by6gmIZsk6GoTkpUKyO3laHoxcmc6b/thJ7oHtwVz9Cc
brQ4dB/vyhwcV5AXbtfCoht2deGBf92ZmAMxG4oZSm4wiAVhqWLYg8uZIMGK14ppztmc6DgMEOWr
TJHbZp5Q1oX/RGtkg0nWcx2lZiqZkY2l9D+ALL798rLrNXPwdggT5QGKxBxfjbDOLYbjJjPtNF0k
3LdfNoSzYdgcU5LKhoNhFeZbbPy96t+S3WNWp7+r7DU+NaS/3TEaqfq4WUfTYK4sPyP4aGg3nTSy
NAnWIMqfvf/x2Y4TEubD4FlkW/QQNDCCK7mC8GutYpDMYDq7RPjl0YLNv23rAtfg99hBpo6gM84H
HQd5B86m+CqLlGtaTgRsXXNBT4xmo0+iwCAuqJPMFcZbr2rp9/vgnOtzvGU3n/v76yGMcNC4clEF
Y2RldbSKZy7SmCrxroq8KU7ly2eMw64Ex5rL4tyPWNpOSoynkBbkanC5vNdmHcazZqnTEV3kYOFu
SWDaf+fMW+Wxa6ovXzY+wNA5A+/rEA9htB/9TempWSKxpfio+Fol1TZOnVMirYCuGdQUZkrYaR1k
EYpWEGhehJR4pt3mdo8MxvqTZodcNRmCgz8QfR0ZxaKiOpg+I6c3cMzOm4SM8wrHXjq6zp3CMq+6
WZ38g3rue2oAPY5ykxfLduL9QjHmG9g9pIEGumom4Qnff9o9CqCx7SCmPADCchTp8KOC3Pcs0C/g
NmmDSwE1GL+m0NSmQxlewtZaHArb8Az9HVhDZelpsg+gaJBTmo3AxGwESsyYnPtePKbpzoLob1Na
nSlK8V3vOTKXuHkaE3Kwbbr+S8n3Nx1i65vI+8AseuSIU7U3O0xPEkdVkM/OCAvFr6VRPC62dO67
KOlO8bUIRVG8OM07bQUm07vksZlTyss0X7eyr7ozqTcFdplp9Y8H/Q69G2CjQAaDneVD2Uv5+5WO
/X310q0KRcNTraQTO88i3Mj7S255WyazVfaVgDpyHqWkZkOS8gc8DUA/mbwJTL/q7Lqemvbm9m7I
72KJzJHcp+wb+2HSkFtvS/ZS41y/EHypQnmoEbvILqfv/78UJC/1tiRv18gkCVdoZanD6FBmSRrU
gGaHFv3zlgTxy2nGqEmTvbDdYKZL/W6rpOMMnhgMv+97EoVrbR2DgdWq0rJ7NQ4kttKa5TNlCnMo
o9ya+U3uPXj/MqeBbh3QFSEzQ/sP04xJfBtNw1bjR1vdkX/DtFUBcqLxZNrc++NNYZGPSb/TxNJl
nJMUzVhwLjxqsM14W6O7XyVUHHZn3tA+nFlbxjEO3UcpxW3thP+KdRXXKcCm0P/5H4a2UVnU10Qq
D5nn6U4OLBUBsweMV12yB5C9VLdpse88v82W424tRWNbb6+qk9i2H2mr2/jXMvngl3WYF/A/w2NP
MzxwPNAAy7rVKug0FntnSS8X8le6H/qKUeSvlqsrULcvcXAz5q4BMirN4cWV4r+pAWXnyYLC7WtZ
98KPPODTjhE/f7ro+Yt/U8FOamq+Q5JN8IxOsWVdAzm/Q7zVaE10Wp+8nnm9ELVtkEnt8i2KlVmh
0lu12HDocb/IGqVZckaDUX6wqE/1I7MEWPS+0s97TDpVj2XNygMqHKxpu5UvmxWegPuzM0Xt3NOg
GvOwnen706CDaMBmoz113c16Djsxw5D+zzoDax/0zhYS3YZ2LIyaHzP1K5BlZKjSip8rNeb3TTpP
q8SwH/I+oo3flfq88QkFrHRN+yZ5ocJGmk59Ztg6pGRm1xM6tsBbwhJquoOYoPzbzjFZIZcxCyxr
MA88/EU+YsEJLjWpmf+rIp267JnITyCd9ASbSL31ie6OB9imUYHbAQfoKQhDwJSZmA7t6Fox5tPQ
OS+sAiMHqrtezEKCLOmGim4jBOxwsiigpb/W7erFhj3yKH7GEAmDGmFotmf9hsEdUmPwm203eG/u
AISE1ea/NIVmjEzqk8BZroHYG6B0i3OmAYtJZrT/BDbeP5RgoNQy2szg3KmK8vkNcsRwtQSqc5bt
4hkh7JcPV2w5/JWGvZHwyEaHA1X9QRb9FMrka02on5kZZ2YpZ8ECdr/+h1kiR8BT6lXNnDOFYoJ2
iEHHRqw9Tgk8Qjt1yXLIsMnCnSrWf/jtxQ/4RIQ1nqnd4aAfOHZ2hvM1pRepo1wLQkTwNfF/CQXm
jv63IrQ5P8Og3hwTGerifxmaK9to0E7Ajsi5QceilkpWiXIUpVX8O+Uw/U0PWmHAI3gHCrQMiQ+s
tAyRGfFwNnwBNTC6cg9EA3khEbqQIiNz6stON2R+5Dr0qAMp7BzvbIbLyfoduB/pP4NBskPMdd95
1sx9bJgipiUo4bDwHULXKA+zVc6eEgWTlXQIgzTphddBDgsj7jxuDP5DUcFh2w4kiTI5LPN6DwW4
JCoWuUr/YEpHKJPDRhQQwFP7LYQENOU2PzA+cg362l65rUlKbgvmeRrVwcumHFoJCUDDbOUwKlZz
REYpc0y6ScB55vXJbCdF7184jZImVNfRV0cjLoaT7Fhch7m4kbI2qvbuv5MCOjppzDdxpsHn6c7N
pbYgrrOsPmSNHAx6XVojch1WGv7QynziqxbkoyE/A/vHGi3fYefQdH6OviqhkBq9AchcI0wNSgHS
0KAfOhjW36kDn9r7ZRENj539t3207aB0WcT+G+SzBIt067psnRku+t+P+NtbJTcv7b/Pke7w7nt7
lQoGBBIdZ5JAk7MbSITUuR1zUK94Wdx8xer+vRmsZh7DXkKr/E2/58/Pm7dYWGmAAkpm81i/aHim
DxTGBJmWdJN8uSX8R4R3JF20u6Ir0b/ryjxqVBtYQwjE8MxJSQEJmbzpjK1RUtVqNSdn+1F+WzMr
MJnEeT1bbLPJnsIE4T7UJNASS3h3sy46WDAFkJp6hviszQBPQsnloCCS8NcbkXhLGtSKyv12nBo6
5sRZZgiaXEI29qKhvY6FEKhCkp9kn2wyL0kwuY7ZLnxc1Qitb8BFFUq4/qzHD6+6i6czIDfhGvvW
iwr75gWiozofm2uSgj4uYCDebWiBa+4hn72FDLWeduLFdTSRKa0q1XRwiEUrdt+UmJLCaNO0Y5DA
ksTu82fjvNDMMxkvvyuQ7e75CRs93lubyApKmRBAywsKPCm3/yY4NNc9/fqFP+3Y5+sibS10Knwn
03LHNfEQb23xZLUd9/1lQAmZgXxSqQxmbWNIhBF7qp5iz261jMGer7fVfUT7TjFvhivgrfwdJMeJ
JqlcQ4tdnTxxwYqb6Zwssd7AVjhjaraKl5tepfHAWi0Wcm4zSTph8AbjeG8UT7SBrF9hTMP03UMv
cu91U6zbfWC3VNxb8fjmq9U3et6mu87yJYtecQagOpNzuCTdEbHZ7jCmyL9okbY/Bu6P7drphG3S
9ZiwOkdQJ64fq3fT0CAwe81ElBPBfdrBCbT4hxS9CKzrhAM1sWw1wzJN6WLxHI8PEc4Zd3e5s/yq
C/AmCnqxJot3jujqR1TdEdDsUOfZ3suAAbU1Cw4eoabBSydqjWXLZ/wP0pLLicZVf2xQQZM8SNq5
ZfP/IYPHgoa+DM+Jxlu5AbaW9F5aDJIf5d1uoFb7iRmU6ysCfSj1XTdxCPz/vlkxQCLSloZQZN+p
l9mqoqy2huKETRYA9gtfFcwtCXIDkYa3d79gjnFpypRq8fQ6GqaBVm31aBHa/40i7ElUuc10JkTG
f/zJ2M7n/rVUhq24BDLWJzP7xmTK848hawNdcA7vPjBeMH0KHAlaSRrk+HzLUKBqGZQRUsM536pj
nBQhGgqxTEOpVEM/41Xj4e9swkAK0fyZHC40IRcrer+W1BsQszYbFZiIUxdKjYYElHtzz3QsGjx0
GW9Y7/vIWs21G6wOlufbXZJapFKXYsK1GWgkTmO53eCmaFCmBDwL6LEMwCtezcweUFqVIr0dhSk6
c6PQIgsf4MPcAlB6/ZsiWmxRSXvZ9jy57EeAbSHPIZsQN6bYPNdVbKEIZS30SfBe82QA4sdEM5Pm
sReoVpH4rVfJu+5bDbFrkwCJYcEsIEcR5NQL3D8CdsTCkckR6tf1tDq+xysAGxOHR0tIwRub6qeV
ROtFN6ednAhH4qmaoU5eRZf/WHbyCk3RpkbP8UDnJ65WoQrDAtBV2hwSKhPyD20ElI3i5X3AvTjJ
RBg73u4NBo9rlTBW8kJK33wXm4jNYICp3VrboCmw3HUoIxZuIRIxs/v5dc/zwYLsoaS2yERvA3DQ
P0aOshH6Ij9ZHWlMhoKb+6UHbX5ACThorRpDYhP38egEzrCbj44LMD3DuO+lZdZG3ZrPRkka2nc1
wSkVYLi5owaX6mSxXIi549TdGyPhHY16TaO6WlOfS6PuGRXDqi6vBFDCt3T7xHkaTPT7/4Lh+SI1
ijulnC17ADU9G05RUwiS9qVT6WMnsmCaYMKG3gfjJIyXaXIQdDYXuoL3GXxxZ6wawW3WERmVwi1u
vokB+VsEneNJbq/IJ1wCkxDOypl5inLDuvUtyp3ua1Ie0eieFHgLpoQWBUVh0K376mtFiRbllfZo
ikB+9qyzKWg1P9uAScXANpS4tlVu+Kvd5LK6PTiERXHw6tefMrNxdvmeWftN93Es72qCZ4/RQS07
93GNQ5cCdH7cIKH7ihFbQGV0D5wFCcv9S2+oyIePyRruPhllDgJ17f1CVkI29dJimeVsQucbsGww
UCMvsnYzj8GZPzeF0ySb4uVVhO/u5C6c5SWu1MLDuAJUmO4iUo5RsKuK1PKXebM0Gh63iolMO29H
MElIN23jKSfONusY7eDUj7tyM4v9eZ4GO42Vg1HRT+XrHJ2KBVKkSTVBM4QNFPO1l8iCq893Z8pX
AsKuxw6dyGX7DHYWINlREapR0vFfK1E79OaySCPz+jPsmFD6qkmFX4Ix6+VC+SYJZZyo68q9fooZ
lQnLnJ4yKJ9e0ACvOANIqMQrwEBZapB8vzkB/z2IIL+zEf8DygkYrRyTqD/5tOLvPyD/UVkFcm9D
06If1mmKqcw32NNRrXdmKMR0TRPsvVKzXTHCkI6zJAtDsQSlhtEyWIZ3WWgLQZz1BAR3JOb6irKC
ysvFZFJysFjHt86CFI7QuHO2BJHz4/V2zRh3T824FslgRMf5bSnkSCWo48haBbUbAZu4eKN/N33s
UrD3mrrcYFxDFGqOxtfJptCKIvUUgzvAxaVkTjlllVSNr4m9ucftIRNZtzk0tnHIc0gw9G8TpLdu
p9D4pmQOsJ24rdDb9ZeLr3STh/jb1bEc85jmWGl/J8Cwr8/kQpbamHoUhnsinvXdk0rjib05eO3r
gTVyJhREwoZ9tznVBfo9IYjznRJzEhAepwjvYMZw2lwI6+WAkXEf9QOkTw3+c6OEHJKi+3oR2V/p
GYEyuHnQewf9YpGVbTHkfdQMROjhJIUoaL6PWPG0SDi4zJs6Da4i33eduS+c2MDcYDZl3vAkaNTR
8w6VfZSvHM0IErdrAXOjsv8kWoSIs63Ql/G/z0rvhBi5YTWBvVvs14jHogms0kC/WqgFzFBP0fb7
6oWNdn+0IjlhQpzI3DLgHpBUZqNCZlGQW9Mn0coXFNxMERdY/AzuG3c+KGZ/XToBrOHKMlay+uba
wtgf98Lk+Uu0uWeAioaBQv7DVi720tYc5EL7XlcODU2hpXUh6N//K4oi/Or8QAAH1h/oIrOzh3dj
Dei4DmNMzW6acPdcIkEInDowZ7bWbYsrOWs7rpgddOzzjMT2s6ult51/PsA4fD6vEnFUDfT4izfN
Z5ZgJANTvRFmHEXaBCnon1FmsS1MKUi/DEQXyQmrRfiZ9Jj8zYggzus12P9bDg6FjMWsAlJABBY/
EZWUeH9c2RL1XKK2W1PsD5lMJf7kgK373lU4bvZejqIBGHrPtdFMrobEAWUVCpqjmwPFqrVO4737
moREAbt2UtnQNOCjTqq0IS/luQFFJobL9KHFyKtaN2ODY4nO6ynDWERpnceZ1p7yvRid3NwDwtv2
kQcZUx/DXInu/EncpL5bS2czcZVT1q4YuBNVyfe8QIRE95DCtZXaOXvF8UIKvjixoe6Pzji9cbxo
1LQ2zCfI/S4fcLkFmum8aELFxrf8bjlU/dFDXnn5duAPIdnhVeXDuvtAYpAa4xJcdvbCVCum0Bqc
GoTyOiDokkLnG3ZT5Cz7ZHBNzqEiSr41D9jW1XeiWQ6ZaEtDH9co2YgdF9sXxLCN+yzDNNcwlqwq
HvgX+5tM+eqoB5UaGTzIrtlDfSJVwnXc15VLP8CnYdU9AvZujODaIs2Wk1T9YjrzVVfanyphLDLe
XF1HJJETlAunwufjH01N/retEZnVgo4FFNvh3zL6LalehGFyC501gDU9ZmVDKYQt1B40LzJbaGX4
nue5P8RaQTHsRoBkhx/2eECIqV2vLxnEpmksdrTFHLIJ+XnKncxDPvQjHIceqNJVQ8xeKPYHpz4v
rsnwW2oKnmSXvHCUbqvO4vKRzZKR4HxssoNBf4vlhm81Pmxy4jbcSnTODpkNAdLZ+aVQzskowQlT
nYukVi938cyQOqxnXVpYnLMjNQ3qUjPI2YKdyV9RsrHGzdPihUzORvpPtOq7OcDMDXwmkGlvjAjU
Cmc1rqB7tPHGUmTPs7dWgoXOwXBIu9RHCIv2nl0UWsqHbLQZKnz3aUxaKlORL7yNT2GB+Qkc4eKx
EIe4sxIIqJJBwsJlZlmJzOUr+tKPjYzXKnZzoynxzZqfB6XW2QI1Lr3RVNs51/A0Jc8R25NYK8kM
V4SgUsaVcKv9H/FaxgqzNWNME6HcCa0yg9qHLb73a2ciuHk0RyongFtkwBbVx7L6DIDfm1OFHWhu
/8XM+txLU62tRq6iswZh3PP2Y+4u/XTPtPsHVkW9v9FNmNJSXX/UEG7VdMkpxAsWnDtTh6nn06dn
mps+SsRSBPZoHBRMr8VzSMqy5N/AJxElaERvl5w9lgUR3w5ezmLi8fda/VR1Xu+OvdYwZAvoHe2u
H3gbrYi5TCi4Tudrcu/FRHec8N3NTDyLh4b8NABf/de6C2AymW5l7gq4a4RWJoUzGVBqe5yPwpsq
SPBrRVIbIqIzYSoWcqP7a3UWXH5exHrEMobDxMsREe3DMef/8b4QEGkLkWbPgtr0eWepZjkbdE0n
UWsTpx7Un9fgGF0IfG4AkO6yIYNrVRWyTczf/8QapzYrFh5zbcZ24lEuou3ukzWhbqlIUhP4r4cO
UM3lFtQw7A8rKOkZzKpb+bIG5oFPAFZOvq8Qzvs92yv4X33XVmqUtcv8Jj9kUMmrXFbUqILQuT3l
0JJ4mzsKvxG1aljNCi/yQfCDCciBajkF+Ikl8VpCJ/eZsSVteZqEdw3NYFE/UzJ5BEno17mSyCzz
2HyNO4NqwBeqe/WTsxMyn7iMtVyY8C6Dq26KHEe9be8s5HGDbMMK4Xm89Y9j8gzuX4EYaoJz6j01
mjFrwa610Yh9g0gMAsAIAEEZ8DV/sYoYuzl+oAXen+G/l5hkiXQvklAkpqj317OMAL9//s/4HID5
X0vxbLNkb19z7NhEbLj8Qb0ns+F5zQuA/3ycV7e/ToCzOy9Zz1xs/UZYLp8Ug7RixlQvifV/+1Am
ty++aa3YaEtzaq9+8/NSA2tceLkNGeSjBdV3PBBDmlFulh10d//u3uAzvXVsVl3pe6oirRZ9tgsR
0I/o3XcLESnAlB9qRDtK/oSrumaOtG7oB6fxUUqMpgWA6Un3eElUc9G0CeGngqz8okWfL19dBmNl
sNHyJLAwSTabXqrSr8+v1yRiyMbU+KEi4OM7KWTYnIJ41M5etdsKavVJob8Z+U5dPqKaQfUSCmcK
T1rHdDZfelzZ+YsA3qA5nl7UNCNtb/EFS+SniJgVd12pmmYLw6MXCSbKpwsMLuNLZzTNOnum3MI6
jLd7UhV6jBW6s6jcLuwp22uMj6mUqJOvlbCXcmQ/x/pOhhoGk46CSNU1+4Z17qxghCnJc9UyPimE
DSFu+33d/PsVaQ8D8M8dzRjIOU9B4Gb+6pjQwK3mXMK/lQr7ZrNzMbZvvODe/3r2bxrpo14C4HfT
h0tR8SQiy9W6F5e/TE+OIMQTE3PI4r7gi1MjbQgTLu3gjjN48/2e57S+uavewQtWzWXPowwPjajr
uCZkhpaG5zq+astrgTTKQCKD5Fo60e0jWBKxfxmDia1DJcY9dKxP7ES+Kg/FFbSPEzU5Y/9tfYTa
qW+izL9yd/KzHYkUI+7YK9a7Tb9PGw0XHk1g68sFsjTshaKr5HjqcFVoVuoMZFw9BGUUkF4iS0av
PuW82eCXgihrWDSgI+aIsaS4Yhx3ONmVgtgffRJ4LmDvgk6AP4nGIG+cLQGpAwP4H3pMD0JStM/u
R3SVz4gr7Xwnx8VqQB1fxXX1looktHoGqVa4z1aaHWVMM7ZzJ6yb3alJFP3EFIa8tzhNtQd2U/uS
gF57HR/W69je0gGCDxYnAZRV3fYbUa/HW76xXASmcpWDBpOS501IMOkinxuroXAoDrmfE1ejXFEu
5NFZ2hijJFPpdzJZVM4J5P+1gEiQv3yMENntLPtB4FKpOJJcpCN+WnCjZEFyDlmp0lxwemeNJi1d
wtEC733IyeqgsJjZA+qMN/9d66EeBbk4Az8OvR5hm3kZfQu8er9BlS8LhWrz9lpcLYrihQFUAeK9
idKUWTy5Ln523MuQ+KQPmzKCLBzhg/4sVaCzsJr7IjPMi2fJdM2C+dJba8e5H0sIWxxw1W7BdK8J
N2GH7NyTgOqLvaXeE8iY1WDoYnF44DN7oC/3sLoIayr02BsafDljAY/h4XdexN3OizI4RSY9btj9
Gur/PQcn0wvE1vngRKroP0e/LI6w8fUYTLAPcI9kgD8m5cjfESXZurdPY8aOccH73txUnVGlN2VZ
JxyMiPuUnwFObCtpZTndlMtuAPEUbCLuMSLFTvWBvmbjy1xeiM9dDSba/BHZL6cAxNjS8Q/uSDPK
s/g6AaUhR7HXNCrmZGwtzFPpfc9P9f/QcaBAskyCFRbNU47P6Mmm4jLhxhOQq87VPg1yStnaKxrW
hyCSiKcslT+bEOAfZ8L0ij/qi5eySFnyYqtnnFdA5LvfLweS/BrA7jVwRFagvHXCqQvvUqBL736r
4KdsaA310jKnHY4UZEnz4oGsJuvHNWlGMCiJpyTBXxQmILTm6iRfZEm0uh//TvKDvS/0sNx1PBXi
L1nPmKbLYaUNWc0ArQGf8jt0iV0EZ933XlyYF4zHIXtfxp89FROh9KKjdZY5DwVroSn5lzexbAzX
ULqpX038CSOksFosa3MPa36AqEdftjXT1OWbEPmv4xgPofH3FkuOFisBIiRHXdiBm5zrwRG5I9r5
WV0P26vLS64LYjNSdk+BvaZtzBokjuyLGy3hoN+mfk2P+nI3PVP138xhmvTrk/3d29N6kD1uNQKY
lWZoKIblA4TLz00KEdbwRnqAwPYya9/STHaSaejWvwQpn/1OeaVBWuCd9xt7HdyKCxkqWc6MaGP1
RicZ4ON8ZT011nH6BkLkEvKfEAwClazdSSLptwaq3pnoxIX/qqwEentLhDvAvNU/TRkNQ67W7x0a
58h4ZTRYqcqrEWcB46MyqIdRdg9CYJwaCPMhVrvljT3VtyXKpLCUmKOHGTmML+fqbq6yDdsaYGuq
mpNPRrmGHlkCBLaipWN7PnL7KZXXYikAXG0j5ABbX8SQf10IeZ2t2ldKIIl/nEOOuWeLJ1dKL4ev
XVUftm6RBo2+FhyszO2uwgqAqObpm/Lr1WkmbHHPvci75cyb3oghqmx5VZzLXtMKhzdsamQN3kMc
ZsMuikLcpuCgDaVmmo3UGNBZv2RulliOEAKluwmyuMqYJT2PllL7yvGcqWLpA+JFvtmRyItAQ5Oj
lHtsJ2lsPEp3hcurkuYmX9sDKCGJXdh5qhxzldWLNNFLgE13j0j/sAJ7+auwzdOjmO8do9+TE6MT
zoParA4odfIgqZagLSoHpE88GLMt+9l7AEKHfTuuIJR3lp258p3gFQ5/jlTP/TxIxAFM3m//kyG2
sc5kmKDUhbdCkz2jMjhf6tGqToZy6iuChYqhPqerrjfaQ5comSYL5E4IbEVeTNpMIVhSPENaFtMc
QjcCMrujYaRm9MaTPlhs00lSwDzyZSiZV/d0Wij5Bw68p+3G4CdyaegN0AdiIGOql07WA/ULqoWr
eRFal3HDZv1ih1i5/IltheCIFx2Alm45BT7YzvYfYROdtcDSanCM1gLMNLjnvT7mnOupSFKciCkG
ywqJDBDM4Qx/U93Gvh8lT0T6U6jHbSMEO/1IYjH2o+yXgW17kn/L6yiaA7YO3+oTU897I2IksWWO
LsWt0Qoy3j0W03GBbYwpZYzzvlLbr892Hspi/314AoSuRR4ZyPOceznl8wFN4Qzg8VINYFdCksGQ
avNYFaz3u2SzES8qYlHLQdnwZLJa7SNQV/DQJAJG7XKHSVR9YX7rSTPfo3GoSh1S2mFTXPlVbaku
/blW0IdWVcj90gu8vXgMKhIW2AQIxwwWTPvSL16aLvoB+RMUx3H6aBJ5hqS0Zj5++siNs5GJQljn
RnuteihTag9PofM8vkpCilkmut2BbTxxkoV/Y82SovmeYrF6SzDYUg3SzKPCcw5L4uOAS4ftV3VG
/OQdcJggAePStwDkURmuN2caxXQcT7/w1zfQ5+MmVLA5xPd/YtKv+Ll1zhZLEl0mDBFkdT159OpZ
qQFft64JJtwLnVQhHD3ePA5icXoihvkyGb6zQUKW/68W/2tAE4razpPMIXSu92z8Rvrnhh8FlbLd
bu8nA5hto+ffFNkIUJTR0oPYcC0MuH2mlxEyFiHt7IUh2yEjgwLcPbMByf5TpmFjUCdidL7Nkg2e
nDPS6tgnrR0zKwyfKYgBlq06rX9nLpoIK3U9uz8fHpiPXKiw/Y3uYprXyX3/hclU+ILu9YUKHouk
/+bAZDW8x5mdod9KQ4h2Jo0n0hPxqj9CVEcogfSwMTXOdI28Wu9ARYOL4+iNZz7NLsGHHOK/8pAA
VGIh4voYqDw5RyaGs/fvL+a+CsneqcF0T3UObNYcjEIqPSFweS/0b0+/aL2rQ99DAMgudIqtiVOr
tjNMs1k4NVX1MR9CFNuINCXXMBzDxD1rpNvYp69js2btOLOEqZPYjiQseHid9DHvSLZLsNkLC6HU
Ff9pGV9Zy5zAoYEGtxIWtsEibue1WqMTUP4YgqLcMHzzwgopjeyZP5NPjgHkA+3iimrmXqZAuSZg
lbZKlZ5vsSJI2bIQ7htrvcFLu+XCXhz/V625EAFjTLg1i48w0LVg/FLeBpf91EW0CwmGi8uZGig5
nOgrM5Dgt8ERvskP3vaL6pVvos/BINHppwPG+W7mkk8tnfjuICV38GHIQF3mMAdaE4oky2gSK+d5
mHRcNTMOZwGWYXKw1sniOVpZYGkjPO+7eBM2tUtDy2XR9SdfCmqFcaCCDOmP861D6F02UR6dTZNm
DT0BIDRUJ/+xRQhMxQtbY1js4Edv0wIlV9d6bpWPimck5PJivoszk/4bg/UvIQng0p7jM3dU5pjC
60LlWZmxFKVgAG1IkdqdTH0fj7EZfKNnJiHz/4IVEDLxshZnoDGIr+ZUt5/hzjx5gFHvkpO+aDOY
Nf9OhLDwPFi9MZvv18+XHdZlUoAwXhyP73N5NWcslYQM6C7aZrKNTRa4UGUkz43qQpUfTpz1Q866
WfCe1ZfZgP/bNXfrcFkzFcAOK8oV+tx7HcBt4X5zLxuhenJVyJ8w05XY2g0ESUsyvBuctoUJTKAg
eJGq+TtM6PDywjTJ4bqqYFge8JdPpDognP6CmIKSFbfMpr873JqQ9B3nJcG8RJn7NjmjapRwkF8b
S1sewGN2sEcwhbYvO3C04PoIo1b/RIt/Ult2rVWJS1iU9F+3wc5g1cQdPPAI6iyDvE56P6H8xUXQ
SfTBWT4YTOrMAdWU91wYI/xn/0OknRgOyBFVgZwWaIMi//M6VSQAjB6Xz5z6/aTOmEjStNbEMSiF
pMu/SlY5TwgIHnEchoZJeV2LijWrhnYnCd524FZy0Rr9kBhsRsFMWR20X3gPGIzvSDsglfVPHSRV
UWeLzeXm/pk1V8AwG2dfya7ORhukYF4SonBw5UJu0lhGqfs1WdYRsYjqxKoyVkTmUyZt/gGl8HyU
3k/Lrd09hlLOHmnysiV5oZaSrq8TCGIM7NnGw1Hu44u+3Xc/Z6rYDDhFAsgt8XvHxGioRUsI
`protect end_protected
