��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i��͌c�iv����'ό1_��A�����G���H��8���ř��'�١�~|V��5/�v�iI��K+Gƾ
!s!&�����r���Y����_#�wBW]LN3�H��'.��j��si+e��E��_�m'��\8���ܺ_�r��
�X�ܾSJWXu�=F|���㪤��"M@�Ɏ�-���1��v"�X�UŽq*����������j��f���/���� ��By��>��A��f��P���i��� ��$�A�qMG�D+1>�$��&�0xq��F�͕!rW�>�9�yCJ�V�n��F9�F������ʉ;3�f{��㫓�~Fy�8v9s������HT��������<��zr���9Te�{�����"�
<�wWq��7��f t�;_ ������8r��O����k�1�x�R�7I��!�!�:'&���>>��#���E=���v��hY��*(��͈U�'�Q��!��)�~t@���Y�D����}ǝ��@D3�Q�m��#�u7�,���t>< �,��5F�se�!���lƑ�.��VOO�������-�ڔE�+6H;��O��#�I��gٜINҔ�+<�Y�'
2��B{�P7(��6��^���߀}*5L�L��팺�ֹ7��rUJ�94��\�5ז�S�o릸�(��"�'h ���A������mS
x�h�)�� Z\�3�3�]ߤкo�.�Gc۵��]����f���Wtκ��9h���O�=��:D6u�S0��⣛�=��wh�s[�ye�ਕ6��0��ai���Y�PIOzn�@3�_�ճo����`f��$�၅co}D,�Q�c�錰��P3�(0N�q�u�����8YR�`�O���+���vxb<������,�',;ܯ
���t�B��l�.�VZ�v�"a,W��l�u=�� E��>�$x]ƙ��/�g���
#T{���d_���9/�#��"���,���F>�{�(ħ�0$̾�:���f?)���-�y��3��n'l�y���`�@��2�  Zk��t�4%��TܪO�W������!?d-B�\�]�%�ݺ��Ez�� 1{�s����]ܷ���#�d�ZD�V�.�rNv�o�`5m]bT�xasө�fV]e��?�T�\DW��"��̵B�h�4F�M���c�;_6糢-�v�E�2�4�����2<��)sX)�_�nlF�� Qd]Z�E����:��Ѓ@�t�=S���,M�w(!c%�Z�4�0W�����?p@GR���g-{L*��=q����3��7���~��BJ���·ڜ����
���cN�Τ�z�����)�c#
ɫ���,Cf������B-bN-�;0��qi�[ H��]�M)��X �j
���k�K^nA���C"D�~4�p����I�9�P �rr%�rC�J�su�pKF~.��C� �:��/jq���e�;nq�S�3����:��E
F#�K��i�U��5��*0#cH'��PgL蘇��]�;���}�B����
���]+ж���t��m�R0�M׭�+�6�췺��T�$�!W9�5�c<˥j�$�������M?+#����)��N[,zF��o�(�|�F=vbx%��h(��^����W<�XT}x�����$%����2L�F�b��Rt�z�'�:��U���hL��6�K[ �eMO��N/���lH�-�T2h��D�D*�.:��0Df���H�W�<��V.^������
���J�����c�N��D�-�D����>@u릨L����	��;�Њ�.*D ���L'QdC��׀����b��H?��zĢ �o� l���G
����{�|�s���d>��~�rЅ1u�O,��'9*u����ȢM���!�a77Я���`Vu�|� ���ٷ��'����V����*ad�&g��	����yA���]�j�G:��-�e��e'�mٸ3���=�#G�+��q�b�?Ì�r�R��L�V���cM��c�b�NOԏA(�@~��+Ж�A���|�ܽ!��Y�w�Wlgs�8@��{����
��ƹg@��Σ�}Xې&�ӽ��A��>�9x2�����￩N��ڥ���0�M-ѩ�Ƚ�op����y(�K��t'_Z���[f�F��z�v&���so�UW�)�@��<=J�����a(#r��.M��*.;q�j�S,4���UJ��NZ��.o*`܌+Ҵ�Р,�?� ٩��pR8yK17O��L�?�5�{��}wP�{?���;!B�����;��M�Ã��%�۳�VSc��6\�q(���v�+��Ԟ�&�6��@�5o����]&v�ETf����0��9������Z�K~��jZ����<k� T���7��U�	���x]�l�,b3��u*��&�&��k/�b�i�@�AU�M�QE/��ܨ�b�<��%+�d���k���JX�Mv�n���҃��կ�t�)��4�עJO��=����oS/t�i��,��I�z�-��T.kr�U��^���AT�1WB!i}p���'"����v�g��LvN��S
�_J�K�s�r�g���r���\{YG���@�lc�p��'�7U���I�]q�{)z��x�]���!� 0l9k;�oJ�l�R��R~4�բ��<?���ɑ�z`�Zgc~�uM�f��F�*P̦�������B0��Y������mWj�L�1aG�'o��1�_R���zІŏX6��c/Yt�Lj���/@T�ɜ�W��*�	")ͬ�C�;*�c�/�!j\��<������y�tcڼ�6�7�9V<ģ��U\Z����&�aoFy�؇�r&�P�N��b�e%�z1��r��ӏ�̒P��2.Hr{J��l~0��xT¢�.؆��>�b��#Wח����*�zĲ�kD-&x�`�,��ˮ�^���bq?ɾ�X䂀.T]܋ɶF�1}F@�)��-�6zI����7��L������A��7G�Xf������Cȥ����ؚ���O����ฝ*1��	�@"�����z2�Ԓ��M�{�>Ӑ۶�W�>&�X���wG$��c��W1ߗ;��8d�oy�M+e	ڼ� sn~��$���{s���9z퉴v�D@��;�����ɽ�9��j~�3���i�%�Op��T���P��#��F?��Q«-Y(:��S�<���n�c�'�+�0
,����C�0]}���Í�$��1�2���y^,��������Z�����@y����iz(�7*m`)_�+%�4�kdi�W��2F��{^ƽ\i;(T������=����0����3I�;1��L�!���>��U�A�'\��&d ��K���tPݵ���}G���+����)����K{[k�N�ēA�C����8�<kD��m�$�&v+��=�����W�F�<��s�`�po�4��=o��eN�6w��p������4Ju6���;��H�$�lc���3Zc�#���@�#Z������_�Ĺ�n6�,󊽕 Q���3�z��Tzں�(��jL��0�*\Y�Ӷ�Z�̚?��$h[�%Ƙ�bp_g���Q �fc��V��.є��h�|�}$BZ�;z���> ���˩D��m춸�+^P�y�9A�-����g���Ǘ��3��4�Y������sHY����EI�Z��͖uh�3e�l�W}p�N��;L�k9�90T�s��k��e_NL���9tg�6�|�Y3�`|d�e�"�*�YO��'^��BI?��x4��u�8E���+����aшX�Q�
��6�k��y�vWV��3�.�#�^IKY�F�c�S�e ���9��\(ˋ� ӵk9��Z�]d0�����Fc�+��]8��6��ca{7�s���A��]zܨ�k�̀i�5�X��׆��!�U3��"��4���Cv�A^4�V�Ѥ{f2����8n�jDnqc��*�;�B�O��>oR%��%_�hݚ��}^X��Pf(mJtr�D^/ﲀْ��V����/�t-��x�������l�I���)��qݶ*%:p��u��'��5;��x��b!���n��$-��o4�!q�m����E�Z�{������6��V˲g���܁ ���X���-V��f�GUg��^?@p �6�����B[��l������מVգ�Rx����KFq���4��7��)'R`���y?~7���L[U���ERZ�������B-�Gi�� Fu�4�Yy��U�5!d�EIdg���DW���Z��W�����BvM"Oyq�C�x,�dɉ�S@Y�"��	c�����պ�.n<14�֌�x	�M;����7u�z� !1!����	z�~�a#��F��U:��1S��|�vg���\�m6��lMS��	wR��q���c�E�x=]��a?��qs�������� ̯�ڸ���6��W)������GE�l�V�1#?���m���&�(���9�b3�/	�@\u�!d����\���T�71����*���MS���q��V[�r�JS�o��km��X͐��#;X_���n�'!LS�Z}S�QE[����@���1C�F5|S�a��Уb�
�5�Y"�U}��}�R�f�h���, ��V��];���*���%sxSA�֌��0i?Y��	�A�:���\x2�I�g��`y�9��f�g�I��axA0xt���/�)s���s��q<h\�; ;� �Tfb�(�S�z%S�+���\�����bZ��<��L�F�hEz/A���+���uZ*E^��f��'��zRM�B�;J`(�t��L�^�3�{,$ٯ�3,	�:�G�+�%����؈{R��̕�q���+h�96��\�d�g��Q&�+�X�5="�\;���� ���Q��m�T�ۉ��6qF��/O��ɤ�Dp�,#ԝ؟b�	����m�s�F��6�&k�0��kx�v3GB��f(D�x����<����KH�eVm����R�>��ݤ2�wY�z��Y<r��l9�\��;�`�{,_v��O��I�g,3A
k^����\�u���X��XX�+Ik��܊Aݏ���{��^���y��${�.#?�����%�%��w� %(�H},֥VŨV�q:��R���q�Z�J�U��`���1��x~
�Ղ}�v�i�6���<��!�]���\R��#�ʣ$�f@pP�A�8KO�[����s���vX��8 ��=�3�L��1קC�p���o�P�XӲc+i�۷*u�J]�b3~�@�L�353�쫚b ���,bĐ������%q}����҆�պЅ٘b�Ap�JN��-(���Z7���F�LC�RMc"���,��,S����b���aA/v��H@b,ܒ���_��x�`<���)v����y�]��w�?.���2�[�%>�u��:��'��?<OW�Vk�Nт�hd�bv����si���Wk��]��"*���G�	8P�Ծ�ں�����n�2غ��p�WcV���)��&l�a�ѳ�-����%@�Fd�`G�e�}[��+[�u�KU��<)���/�h��<۔�'�	��k�J�oۘ|(��݈�Ne�\�I@��L�h���^�>l����ؽ��W�0��geB��{?�h�@d�S+�M�VB"�����x�W��Dl�w�g-�j�x�7,r�6��#ɲ�ʹ}�N�[�U!6�ٍ�~�2�;�&�e}�n�}��mu�a�ƽs��-00*��sjWNfz��%�����X�x��Ql]X��L� @T��
�<zN�&!l��?#�A	��V绨�H��$�$e�����7�.
���)5{
��J5}
�5Լ*M@F�J��N�!�I2jӒkP7��
�_���8<��֥�P}'�0��!^���`/�A��Q�u�~�n�o�T?�r��fxi����"��ٲ���tu'!�m�L�>����Q�>�r
���j�4L��x�Ȇ�m��eŨ1�HMKq���O�y��?�W_��D~�e롡���t��O;L����e��/{8�XC:��)�œ��P�v3_�X��~�P�~ �A�d���hs�C
Dݼ78��x1q[.��M͸���'��� $Tm����#���+�1�c��냻	Fj��*�9u�>�����ғ�-?���K����៰����iC�5X�d-l��?*�~x����[�[��h:�<�P>)$T֙bx�>vD+��(�"� ��>{� �`N ���TL�̵����a|���B��m��OB/i��vv2�}u	%�ܹ���7�ْ��zY�ѝ �/��˪�4Oh���QT�Tm9��R����`�6)A҃��`	��[��]��Kͣ1m]��
�]ʌ{}<=cC��3�'ǭ���Z:D�v����'�U�,+�;�sJs>5�����tG�
���ߛ�`*?}o���2�-�E���Պ�����*�P%Z���7�T���nT�Jf�'N��~�
h̩
�Z�����.R�U�'��x�p|֌:	aJZW|����cN�o�B�ʡ�_-����of?��-�pݣ����Z׏͔L�;�yH�2J
N �&���'��02&ؽ�P>,h�����E
#ڰ���qz�0����ݘ �6����[^=vt2C�R��� ̲���/����Y�3B�؄�=z�4@S x�559���������԰Oƙ��?�V�YY�F;N"�t_��#�N�f4�t�7��v�.�6�������kV_D�"�U/\���!��\�8fNơh$��U�Y�\[��,��Ǹ��/��cٜ/J�j�Q0�5=�	j֐�g����=t�<�i]�!%�<��}Ve���r�۝lc2�ɲ�0X u��w�/|qG]�G3�B'6��ST��Ť�k�g����@�����3�;���j�����-���ץ����$�vWf«}_���Wb��cp�'��jv|~�tj��f��(�2��dҁ(S&$��$=�� <��[?AU�
�i�%
cu�Mf{�5�����1�B���rh�)��;�5Lun��m'ʆb"4��/y�a���O,
I14�!#rT��+hs@���0>F��Ժ������M	'ºW�7����@&y(m͌�|:X&f|s�	���������is/���I�纒��أ���7)�ެ�*^����jgXmx\{Q�%�x�y��n�|��+(\|x�p]m /P��sD!L?i�4&x�A�I)����^m�r~n���"���r�]p� ����G��K�9��h��"5Ήfm�jO�U�e�f*��.DFr(�u���$��Q�,̧�
࠷����Wld��n���aNA,졗����(Ȱ��C;�f&��G\��ꄮF�?�8=vO
}��������P�Z��k�~&����FKq3e�Ӊ8��z�*���g0�g�M�J7�����L�D� h6�XO�Ձ���XN�V2/�r�����,Do�U����6�rƮ;oi�4�.="�&3R��|�����C���Қ*�b�:��x����u�0kC>�Ź_�'��j[Ώ��t9����*�������glH����;��AZ�+���{J����{�� [�9��IX |p�s\���n9�U�H/0���z6�T�M��^�:���v�Մo��hn ����w̸8��%9S���a�� ��:VEǭ�	�Վ���g�}l_I�tԮ��)
�%��xW�?f���a��!:jO��_%��|��h~�����j��[��ڪ�z��HPSm���m�F����t�y��_�3x����[Xd��D>��6 �F���*�YC{��c�\��c\j�dO��xYݭ'Y���.:m�{��y)�-���s<�u��npz��j��v�ᓕ%A��9y��qITxv)�M���A
m)'��96'�[�,6B9��G�pn��6�B(A���,�z��-	�,O�d������I���/k�؁�AS:z�����c6n�~��Rm��-ZR�nJD�O����^ ���e�f���9���uԀ�����_M��m}l������!0��> ��l����4j"(z%W<�*/Ҿ`��;�2� �ڌ�/�yXp����Bm{{qgmբ�n�(�Еf�,�_f9W}�)��/"G��5�@�f�k�դ���Y��&3��_���Ã�.���V��%JƏL�&��9~NpD�j����mg(䕗A����(�}��h�g�®���������2
Ǒ8��I6q6��VG���i�7oV��9�$�.M�5�z�ڣgJq5&u:^b3�3���o,���(ct���� �L�n��2s�ȜP��"9[��$[<�J��r������z�Q��S�8��oH���_+8x��Q��n����=k�+կ��vPd�^r-����*WQ�ӺM�둄��_S��Q��Q���;��K��+�B�aE�S�t$�ّn�T��?��"�;�T��7%���I	+<t�x]��ٖ�}��~
�6e$���n�zߒ�i)�7�d@�u���X� R��Wuf��C���0".Y�!l��O�'W�?���(�^���"{e��9Լ�0��k�z5�:Қ�C�50L�!d,[�Eߗ�w�ԑ����9�G�����a����$��u�Ą�q���,�T{�{��O���AkK�R��Q��K��E�������y q���$�Wc���(�i
�F<���a�P�ӥTaK`���:;S7���'s�Y0*����U=�»�99+���ܩ[Џ�D/[Tp��+�H<V��Xskr��m<C��e�`��t��l �2v02!��P=�J�㿲���fX�!��?����j�}*��3���m��	������a>5^l1Bk�����:|]�m�s�H����=�s#5���m���l�6q�,�*���QrC���k2	5�OfD�ҋ��b\J���i�|����7((#�q\j��[��[�������DRw<�߭�Դf
��U���<F����ו�tC��i�K�[z���,]�c�GK�&j���_
��Or�K��O7����9t��`���@���,aw����m����X�]�{~���yjmcic�?�3h���3t�N���+;;�D4�X��8|�Yǡ���f�����PjxE�R|(jNB_$F�f`d�0
���8���m/��m�+(%&v%�;�����,�"9�=���ݤ9L0%7���˝��[�I�ӶB�������䏄�n��팉�>A��Z�����v<P&��g3C2kY�s����wR�5A�$��7���,�U��SY���URl�e���g.���I�p?;˕"4'� ��������	!]�4�AEЋ7�{SJ��i�+F�sk?�3B�ϼч�[gZ5z���lm̑�oP�@���D�39f6Aa�Zn���y3��\X�~���*4b#;������aG�
bt�q*�Q-��c���^��&gJ[G]=��Iy0;��Wo�3��UNZ�կ�#�^瑱k>�6�1�����'��p���2&0�̜�������5ȸ�c,�*���<H���9?�6�H����,�a�E�B�炋A�%���r�[�����p�>N���d���ߠ�ΠOD��y�~<��������W��M,Ð>Nw���S�OjM�{���%%>D�o1�.')�:w�S���_��r�ߪ�`�W� ��/�dʒBN,���"Q��l�/s���Z]�*�^?'ܹ�w�,���_5�:#���n߉!���ͼ����i"�a����qW���۬��`�t5!�Oz��w�QpK^���Zox�uB��`����|\�7$��q�M��v�6�?��t�v�8�4�c,�V�g�%Am)՚�7!eX��L/ �Fae?*�՘I�0����gL����s�W٘��`#�gr A���bRϦtk|�ѳMn���0GTM�Ǽ�*�Td\��7R���[���D򶿵� �	<:h2т� �N1c)�/�To[��%�����t�[eK� v���#]�c>���S�E����o�#�^�M�������`I�l�>�Y�UW �iQN�EH[��B�8z�ψ��Uiɧ��@�V��^!�l��ZUH�S�=�YO.�`O��^ܦc�(>��{&Р��Գ=q�oi�w�WQ$�r�As��/hj�?�hGK�ՌP�|�@���A�T�]���R@���h��ĭ�`��b�6�W;I{ٹЦ9!X|Ƙ9R�O��q�毺4Q=������IS�++p$Զ���3�+P���S�L$w
��dJ�)��w��_�gL&ТK�q�������a��AC���d�ߛ����V۟�1�h�֏�"��x�5T0�=H�|���en@����B���H�^�Ip�7��(�GnX�����E�?yJ�����/)�0�2��P<Y�'+�] r+�Ld�Z�$��8*.������������!�x�ck���:N�_��k�St��5\N�%�LW@Ä�6���J�ʸ4��;�o��olF��>x���D!&��P�D�Xҿg�M:���W�6��M�v�2&x% %����u�H)4��X�Q�k��0�`O��u=���=��M��� �E��ۀ%m�#.�ujA	�;o66_��a����۫b2֒��P�r�E#gᾬ��3z� �ħ-yx�4P���~^��6��n1��=��Ŭ:zh@�4&�t��lUāw9��=�6b���0�#
���|_�Bb�g}8w&���z��'�!�՘^":�I�,.a�͉��9!e�{�y�̽Ú�P��^�GI?�Qt(��^\���J���X�w6 �l�4��X[���M� ���Y�C�w�^=`��I+���R��5�x���E�R��g���W���E�Y8�G$�kD:�{�:D�uK�V�5]�~E4c���O\D��/�D��9���lR
����BT��o�bϱ�w6���t��7����}�ME1�.�?��>�֔�n���;����7[�L.}з���g�K�S[�  ig;�*A|=B�ǳ�A	u��66N 7l���<��&�4�j�hR% M����Ou;?���n���ݪ5w��u�V5�
a�Ȓ�9�)f��
�4�j&KEy�+�?N��$����BPn�ٜ��-'�ݿ��Y����S������K�����~_k�!3��
"�B�5CuuP�����ka3\��KZ'��|o:������Vnp>>����d��b���(Ki��r�3a��Aww<�t��p� ������]>:]N�*"��%B��Pn���x���9/����LX+KĀ5��s��c���kzvo���OWW���"�.�-�$TH�H�7�sx�� �Ix8̷ɇ��`d9��� f,�����'(�BW~'�ujk�!a\�F�~aˈ���^�n�)�K[.*���F�ꩀrp0M|�h�Z�U<r�P�[F�:=�
uZ��"q.�.B�+jwS�fW���Z<h��W�ICZ�	e]BWb��É�d�c�`9(%)��nC#/H^}`����|tp�=_��v'��x��3�ʝ�pjW�`�=�&Uܪܐ܄iC/�FZr�F�QH�Ɣ++d0����V��0�e�f���X��u?�qg����D:�/��������ҷ�ǿHx�%��� ��q��/�ٵ��`gg |ߖ�ʺUrT_M�I}��xz\=�1R#W�6+�I�p�(��u�X-�0��c%yy�M�Xg���K��}�2�l�-�ཏ�{�u e�w��͆�U2r�(�6Mui
ﲿo��zP�[�z:���y�pH���Կk�����Y�;�ż#��/D�Lއ��bMa�K�`���.)��X��iA��y%XP��I�=���~��4�TR�%�Ԁ��4��Y	�CF�fW�K���v��{(��&qx8H�/��a�XG���_���0���oi)��2�������oj虯S�xɦ�H�T7�\˰^�֯��C.��k�՞�2Ok�Ѥ�%oW���B�U��(I$�C&���xG���i����P���Ql�c�6���P�0�.!h�c�!�˒�k�'�ô����$~�<�o��ޮ�V()h�S˯�*;S�v[|v�!�.�����V:h�g����'�D�Qz��|Ք�@���Y��?7��9�z���)6ZF���il���ʪ�|R������:����j���{��Da����:��n�G.^��� �'��'������E�2�Ҥ�ds��lrC�Z��o[��b�7/V�/O��܈�.Z�Q���a%xZ2��4E<�W�VХ�6YF=����l,��9��hwZ"!���	`.6#~�(�����?�(�^;�S͐�(8�hEH�G��:��H����/��Y�8�I�v~,� k}�X�?��w%(�x ��{�ID'>��И,��=%�{�-�|�L����k| �q��ڠPN�D�a�J�;��D��М?e�3~��2�I{W����9"�?ʞȝ�����\����8&8}�\����X�o<�dK��K��H;_\�������/3�u�o����S�����@�C7�b/8��5I�}\�󼯅s��Y&W �&L��*9�6K���G`1(���F �V7�[ؽZfE+	�=�2v�7y�ZP8�)�vL�s+j�����g�ײ|w��ȝ�t����N���dX��஽�ɬ?ݿ�s���<5m�
qqu���c��"��G�~�DI��:��y;��~��I�jl�pw�k��@��X'���ˑ�����"�}���K��v�9$�x�`%�xgM�C���=$5Q7s�1��C义��µ����b�CqSȮ�U#�-�R ���?�i��o��i�aȗ5��O�+��<�~�&9���"mW�͊�^ȋ_�r;�_���8��h���c5T�����$3���w�~b�(�p�(�Yk�.�e�k՝z@�c��P�D�d!�Y�:���S̪���*��ΣK�u0�N[8�Xq|���s��Hɜ��p�%"����~��KԀ؄�O}N|
A�L�B�.}��rw��8�m9�f+|�gwy���H@��f�ܵ�h`�� �}ج����P��!��4 ����>31�A�|��F
��S��֏|0�@�}��a��R��}Q���C�7/R�f��Rn�qa�������CV��Ջ�oyl6\;+V%�SF��B [�[ၒέ��1[��&��(q�mh-d Z�6oG�G�ijȁzk� c��+F��G��D5���ĥg���y�Aƒ#^���xM�D�(�X ��T ��"�r6�]�>ج��Ⱥ7z/-��a+�ǃ���x'_-?L*}�ۀ-Hc5��/d��F�F���Q&��W�DG#Yc�.���JV��@�����}��E)���mI10./dܥ,�|7�G�B/9p�h�--F����"��cL�+�&ݫ�3��d1o3��{�񘍩���&��W�T��1�h�Βy�O��N�.�[u���G��1Q�����%$3�g�U�pt���c���Q��O�ߩ�Y�P��Z��m�h��RXZ�
	ՙu��㩑
/�"�����Ԑ��CWc��g�q@b�#e^��&��AOPn���(���|�4u._*uKkz�c-�}�9Dl�@?��PD��B�:�q�5����e�����҉��ǒ�I��}�ݱ��@NO�F�iPsa;�'�aT� �F��l��n����4i��h���[[Uq�K1%.�>!"�x���yX�|�_�j�Y��Ĉ-
�OL�q����+�:j��{���C��+"4x6k�}"ɦ,��h��c�?���-�=��~s�.*�u���+��8!܃8���g��'��_�!�@|�c$Tƥs���R�����8�>��a��+�X5L�<��v-~n����^�[X�;a�F;��K�j[QD���Q� 9#~7v���N\l���d����#����p��
�
���,����D���/y�ELl�\��q����v�i[G�:I���2��*z�gJ���Xk����r��`Z�����|A�w|w���pZ��� ��}�x_�)5r𜞮�Yk7�^!��pvRͅ�E{#��Z�<ӿ����	L��[Xl�c�rz�ԭ>�!R_\qsl9�ns�`^�O���;�a�	p�Tà�	,�[8�ǄD����Z0��W��NO2��I�}CIq��aaNd.i�(}R�m,"�"i����h���"��`RTO>�V��\�9M!�l��H#p�&WP����ԓ����D糷>�׿i\��뢴�P��qث�V�X�:��1|�\�̀U��$Һ��$�'y��0�n��ˬ�5�����FvT����_��]�GZ2,�����<A���U����m����/u,x߈�0x��<GiU$�3��-M��ƕ���	�Ћ ?�>0��Or�'
��j�daQ���f�4����M-�u�Y
���D��St�q＊PLh�ͪ���q0f$��8���Ŋ3o��Y矀�g
ռ3�,FNС�����#jb��a�}9�:�<9iB��.e�?_��6R�a��+�G3ҫَr���i|C�;]CW�T�l��n0�Qd�s���yL�:]ӹ�[K��Y��z"��a��w�u�g����u��?��5lW^���{}�v��u2�*�	��IS��������R!�����8R*���A��	���~)��O,�c���C|�]IL�|�@��(�������w2�Dx+F�@b�\x�F[CQ3�Hq���k�E��񃒌�*b�3A���D��XaP=�P��'��z�Y���RDxs�M��t'cv4���I�S�o7\ׅE�­�`���\oc�&	m}�%�ho�����aӚ@�3g
��C,D��W��L1gɇ����_J�*Φ񔢺����=��̔�.P�dUwG
����)�)�3ּ(�W�XF�?ˀg�f%6�V�\C"�ɔ��J-U0!��Lx-�	�*����̊��W��P���I,��?&�>�-i�Fm��:*MF���}K�1v"I��m�#�/�OUs=�P5ύA��oʛyU�F<��(p �X�Br��Z�p���Ѱ���M�.~�t=�o��<���	ɖ�#9B��׹�;v��=�+�<@�<c�?/�ױ��J"��>�a4�����GH�0���<قRw���fVG�~��^Y���K�ys6�"�_!U�|�߶��l'	��l��nKY4Vg��ZO�e�	M�A����'�ϊ
���)�ޠ�F	X\��5��t߹��~YՍx�Rh�Q>�����&�0�+8"�euG}��a!Ҽ:���,�r(���8z���OV�� �A6�J�Dc�km]�2�NcSl&�#E~ޫ!�P�{�rX����ə%�'\_Α��Eq�}=�y��&��3��Y~Y�1S9~���K-��F���*�]�:zߡ]���ز :����E���@�x�E�;1���*���X��#h���%N�Ы%�Q¥+T�}����᎚�%T qUWn�
!yW D���+=��� ��_|��eH� �>6 ��Z~�5-7�� ��lH4s
M��{��d���K3�UB�ͥ�L���[�D��+G��.��E�P��D��΂PB�+�]s�l#�N�7��wqI���͇{'��U.�B�
i�n��D���Hz�<=b�
]������jv�:�����/B�ULW&i���O��F'����QBu��䈕υ(��a�S���\I��۰���1e��O���՘��q�:���ρuƵ�?>z�y��_,Ǡ,|�j�7�M�'���
�	@�z����4���*�zl���sr7C�$~/��!�D4 �R�f0u����x�h�ׯ���]��� �;��r2��4)�B�;�`N0`�|���Yןh���!�n%�}3K �c��H�����2�?�U�<�"���leE�!=`Z��Y,������+d���H	���U٥FB�����bRKM�@ *�ݧP܏�E������9��j�EQ���l�R"��UN��U9��sO��A��;⛢ৌ� 1/.�ރ �%����iH�K�ʻI�mĂ�UP&�k�x4�������œ���������]���Rk����fs�{��nfU�}��a:���fpX�)NW����븪������7Իh��l�I�H���3��ՠ����Ƭ�%г���`!e�`�Ξ�N3DK.%�y�`�E�2�ƌ�c���.��Q�{�Ǯ%���f*��g�5�ҁ^�<o@*�rTv/��y�R�V,�T�)�߱�( h��6��}N�n�t:��6ui�1��_��%l���eZȶ�������^���:�X���t��%h�K5߈O�Y^GV;7�-&�^��ra�Y�1�(�����]����	P��"r�s:�6�J�j!9���s��k�8� \ �V��ě�a���2v��q�m�J�NZ(�z]�T�([Y �Q���t� ;5��c��h��[�W�k�*m���n���X2�UY���MV��7K\�h���s'�<�nL�?)X�9Y��Ў����o���,�㇮!��t���c�ub*P��b'��c� m:�ĝ��UvV���딛�n��{n&A��ŐTN���	�Bh镗��/�)����G�k�(y8�ı�Ѝ�N��A9��<"	�(QSp��G��=���ZF� �$_H�a4K�bOWH;�C�'��Rha���7��}x�>G'�����A��G���
�g$$7�f���P̚��&���	�,�C�{\}<�ndv_P�מy�0���{(5�ʒi��	"[��;<7�f���"�_�z��cXNǤ�UE���	���/�qP҃z8 �s�zS��`/^T��-r8�r�'J�l���.3��w�������X��QMa�y��x�^��ӸuN�9fv����_>S�����v�3�E]�����^Ƣ�ߞ���n�v�@���L���l>�����D&%�}�+]56p;�Ξk�64��<�n��)�P�m��(��Ћw��}����G�6�j�֕pa�YU2~��F�]�+�v��l��KH��Ug�������l��-+�NB!7�n�$�%���#��=�{��P*��`�,��z�R���;RL���b�hӖ���6��2��E��A�E=-T��Y�nw���bF�$��	|4�A��M菆�{�O��מ*�k��I��TN�e�Mu�lw��p�ֽ�L��z!�CY��ڨ��!�P8\�cЈY���Q����C_�]2�+�=� �*mI�s?�����<9,���c�6d�1D ���t�+Ntgd�$��ni�W��^m�`�M��u<��k<�6PF	��݃�ˎ�F;a����NCq��%`U%a�6=o���|�n����I�*��R'C�X{��k��Z5��(U�y��5>�x�@��Y�����͊�L~�#�]���TS��F���i'Ċ�n4�+�tp�aUq���������t��s����AC�@�_2�����})��++�3��Y��6tf���K�L?���p {���^|G+f�PZt}��n�!A�z�q'n[7�6&.��`{%-�3��3t�(dM}�dc�%�^��	�$�q�~�f-���v5�;+M��Ϻ|F�� ������g����CX�^H�/
U�iY}�Oa�87\&�h�^�S�MsF��P	���Щ���q��f*�k}�Eʤ�Oz���ݐ�i�<�vQ�;������>�g��E��V��XL?���2�βq���0@������l�4`���f�"���
%�]�BY-���k�	82z��kv[������P;�Vy�k�1B/��21@�l�M��,::���;��W�V��]�R��Y�z���g�f�����REN���SPl,�L`������y�� 
��l,���=�nQ�Ɖ�:ꭥ!6��Z7��)�/��ll�ړ�S<��C��ek+S���G�+,�k�$�ꍲs����"����<.S���9M��4��b��k�"���V&-2�9�:������!ۭ�uw�������6�;x�,?��&�����itU'�k���6�Ͱ�.�&�KȌԊ{?e���5�9�؊[e�\�&���NJ�q!����Ln�X@$�z5������&z/"�SÇ.%b�?��Ɯ ��5�K��p�0���0��d���p���$Sɟ /0�rM>�a�K�LB��m��������4��D0ku�$�uULc�00{�q�b���Z�̿`�/�j�a7]NpJ�������hS֡�kq|���ҔܐR.le�\Y��4�e�볥�񘞿����+�&�c
�	]�{1*a�=RN��Ǎ���vCe$�̹_��hj���+4�qG��{��u��
�&w�4���-�Î�����<�?�6�P��{@��d�!q������B���3W!u�w14��K�Yf�I��$`���g$�0�ﴥh���m�b�
��r9� �7#NA�N��������r/	�0���lo|08��X�W|)�x��,h�=A�	�h�9�:��>�aW��Nc��;?|�:̋���EV@����>P-�Q�m7+iw3�V��޾�V�
|&[c��r�m�nr���̲oR��6��8���$�1pj�s1��n�3(�)�����'��S8,�P�X:�ܘO�/���O�W�M��^��r͸��Y0��ր�*�,��9o��������ʴ�lp7�f��l"{ޙ���C�S�lȶ/�[�/���*9����7-IV���?}f�۰��;b%
3I��d�"E�+��U��r}HSl� Ԋ����j����n���؟�Jl���D�/
����
�LI��t�!�c��mоB��>m׵��,̃$�÷�?��\��[ߩ �Ņ_���:=�: �B��}��`�G�5*oH��񈨖����B R��<yV�����[~��:�P�����������H���dh)F����]��[y,�	�R�z,
��
A�W�7J��|��B[ l�6joH1����P3*HϨ �K�W�,��@�t�;2Ht���V��R`b��7��A��#�	�y~�I��Х�X�9�'��O<���F����l�uoJ1rG�w3��i0BL�c�!V�Wf%���-ԛ=�@�`�G�I�>���D{L����`�lG�{�We��5����(����
�l���T|+�\�@��9�e������9��xPLd�K���^�y�
�k���˗JA*X(s|�������_�?��
��[�>� V)�Z�-SPKt
��uң ����/�[ߦ��sا�mdd��t�U6�?�[{ӆ�*�)���c7�p�Q��S��V��#�<����nx�������_���s����!+9]�M���˚vE.���e�=�)_v�VG#��e��9�IP��$ق��}��)�$8|):Õ�#�@�g$�-2���6���E��բs0�n_��As����:�&p�N���Fk5�ɑ烙�t$��������Q�1��b�Ġ1�VT(�rB>��ّߝӣ����o�t�CB+�]�X��^��W0�@�=Z]m�0,;���"��"E��Ud�|��Ё��syҁ%��$C^r�D��S��ZN�
�x�wT�Y��<H��Qg����/��U�����E��*�{�Q���%�l�Os(�ʢ�7ܙ���_��\���T����J�XC�- �V��?�(s���k=ru	����(�ͤ����U�R��bJ�qq��UU�����Ѭ��u-r~��,���3j��N�q�@x�5��w���]N)��b����R� �#�oь�ǥpN_��
S�Z�vkH���/kO��g&�@g����]]�ʱ_�襨���(�J8F�=��!o\B���C`y!��{�{�_5�Ŝ��#���Ȓ��POY������ ~�1|mJa�����d�?'�t����r��	�U;�q��H��w��x��IJ!�,�8@�6p��������˔ǿ'�T��p�ՠ���L�'���}�u�"��_�����~��\�48^vX�� ����r^��P�ʾ��uE�I5H�n�	�sOl%���V7�
TT �Z�(�gC%7RZ�"�r�-�b!k�4�~g/o�)!������Ms �_�\����C�H[�����1�y'q��sH�1To'��y!j1�}�C�H9ֵ�ۥ������ =-,}2�r��p���n�)/�U-�D,^�k�O��z�]^L�p�Ï��T�i]8W^��L+ �@�d�1�Q	�Z�s���R��+����\Y�頱��ʷ�̳e�� �]	��h���̶q�͒�<0����s(�����^��!��7|KwT�&��4�R0�Usv�KVh�Ih�T�̲j���{a�W��������f��f�?��*?K�|VP�<�v�Z��_k��_��;+6����#�K"���[�"{�$]�.3m��j���p��d��[�4���<�ŗ8 �$�
�����T��_��Wdyq>N��_|�Ķ���I��Z�Bɀ��O�7w��DiQ�\ф�14*���N_m��{����x�-�K�p��}h|+~���D��d"Y�~F�����7 )�u��G]T{��MJi0�TH��)��s�� L&����e�]��OL��'tsC����m�j���᪊A�@��N�P�Bw��H�%n��]��,/�aI��uA$�Q���b$SQ�)��E�Ӓ@H5����7F�/�7@�bh4)�&�'�_�}aPѽ5�P��#�8��"dD����"g�`��B7���[�����g�"�yB��QI3Ӎ�Ct=l�/8�$�Tc¹�j�O���9�dfu	�h�eW-��|�r��BRR0�X�rCP=WQ3��:��v��v��XI����0x岝U���8�6d͵��#��s���|9{��>������KtLSEm^�����V>�a�x{A
R��J�ի�bO'��5sA�,��p���q�U�c;���J��Z�x�Y��o	b�c0+�����I�{�@�SDл+�� ��p��ܭ��O�R�$�d�ߩqPA�cT��h��|���ܡ�P0!6�������8�V���L�u��-��&Ph���-�s��,:�5�ܢ��OZ�-���|�:���gّϸ*������jX\�;%����'��g�z��y�O��������H0$=����I��<��D�q�ph�s�o����;�|�Y�4���o�Z�/�t��/E��5���Lըj�S��DE�UoóзA �����-��c���UGú��l�N�|���[׌-O�̖U�1`�P��里����X��١M��|�J���������Q����Q~+��*�,��:��"/`[��Ӊ�d�FS'�G���,Uq�������C�wUf�v�>Ġ�z�����9���wa4,���Ak4È/�M���k���@x�����j�6a�?�Әo���S��J�j�
RvK�@��u6��7#��0�;+��۞B�UN�w���;B�}��_�5M��8�Y`�ѰM�3\�Y[���Q�/���D�ʲ��Jf���#�e����%��jث.J�.]'��4��E�Srm�Pвr��e���i.���ֺ{2&�`Z+9�λ�G��#ەDO�T$�	�|��7�oǹj��

�����&�m�*�o�/�n�n���u�i*چ'@�����q��Hx�!���&��hL��ԏ�Į���6ɚ�P1��z������*bL�5�bD	$�`��^��H/0�n�p���iКG�+�C��4�'�|�Ϸq�i�<[�<�o�e1�b3�h��n��� L��4���W�陀�+n=yw��$!��~�[f��UD#n�r�����L�;<\���Tadr����?�	�w�6x��a��� �^�,a<p� ��H�DfV&�b�}ae���F`J�:U���D���ː�JtI�G