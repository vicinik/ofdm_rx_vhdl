��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P���S����OM�̊�Ϧ� ���9�m�4!�PF�?[6l�?Ye0I�'>�������!lݍ���p�^F��ˈy����K��)�KG�1��C�rOe�K%��槂�
��%�OȂp]=>[�f�~v�m�/�a��Tԛʐ�i�_L�`�v�,5�4�U�ß��v_x���fw�]��r�r�P>�QP(������L��Tk�wV���ĕx��D� � ��g�y�6�;���<-G���C�c� �h��_���d�&2Z�;��z�X�'�*�|̺e1�|�b�@'~�T�;[�5��z�!m�j5b�-�x4`"�g�,�I00�I�R8Py
�?�k�dp�s+�s�t܂4�e�&��@ �60�k��7�~;�؂�dÊ�(;s���_�����VDO���;��S׿��.'���1/��x��|Q����0!�ې(���f�֘�l�
M\����x��Յ4����+ ֘��('��S�
���yupi��Z���6T�;��E�b�X�ۥ��D��������^{$�:�Q"5lQ�āF���j�1��u460�w��i�M˽�L5�G�����6A3]gq��M��v�;�d}��p�[���H_��X��c�C~�C��������
����gv�3�c�J���M ��}Dڌ\A��C6�I ��� ��HW�x��GȢ
:�N9���!V�=N���VD��FȀ͜4�&o��Soӕ��$�,A�X9�A_��Ɯ
0��{a/���Ȃ8�8ͪA�X�{�쾧\�y�������z���)X/C�=ri�3''��J��Ԍ��YA��wN��Hw�3Caa*�)�+����|m�*�i:�Ɛ�N�9�x��CC~ WLR[�4ش��-&pݫmt��� ��������;T��z�Q�<p���U\d�~+�t���Ix.�}�����32ټ>��w��a;��� @H�6E4�����(ud!�������K�y|#�+ޔ�
I�2)a$T]�p�R��
} �ЉC�:��0�h�ln��	w�g�[s�|��ی<�yG�ָ�8	��~C�*�<*3�::��Ȭ_6�Nc��sN����`Ca�I�@@�J
dz�
L��$��P)���wځ��7[��+ Z/��p�8oڀ�μ���v�l#3�5P�<���(�E�!�l0��I��!�E�}Y4�����od�����I|�gv�����ҥ���xT	 9�?O��T���*�{�
��k!��3N�T߬�Ma�&7�Y���P�"%u'wNsYMt7i�w
[˖ �5J������t�@�|ܻX���c�Kz�=��a�`r�0 �EM$��U��*�ٷ��X<T.�sD3��2�D%��R�2��(^Wy5�`�&�����=rg��WƩ�H ��{Nʗu<0���"�'D�wѧF.�F*�f�smz�bc8(@��P���~/�i"�R2