��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X VyʐPH:7hCQ/��B�9�8�o!܅�����~8O��"Ve����=
���c̢r2v_j��:��;G�N�|碗Ӷ��������ꢰ���c��������2��&yP}L�1(J�~d���l��&՘���?t��!��\�^[�� �b��֩�Ri��?j�a��'�t
hG��rR��B#��!���o�"�.2�O�ObT={s�l����2a�<�G,�\�MėO��N@��ȭ�	�������a>��~[{�3��<9q�?�iءg��i���������E�/6[#�>Lￇ (d�ta�GW��VA@��I
�i���E �<�u����`�Ҳ:x��,y}����{,U4G}�A��BRfcp������2w�RH��2^���|W��Wk�ߠKc=���LXXY��XUe]��_�&C������w���1�Y�|��ɨ�ڕ��,��p7淎�3��Q d��-.Hip��W���9��R&�$�%��Uik����i�c{��/L�Jb��e^,'A�<��2-Ê�,��_�Hzxs�Vn�1�A?�nĮ�FP	��BAO��K��$�thBC64���T�Qds�;�_���I7�* 1^=K�!���P�������)Gs�t�{7|���up�32�S�t7����O�����rL��6Ԓ��'v�5��]HF�����"RC'⢺s)L��<�z�|��o.Y����ST�/�6Ѯ�\��n2sm�xNq�|�^��r3������X+�]C��u\[�勨��ȅyƎ��(zs�UV!�/���L���2�����|Wh� �T����>E1��+��&�3���)�]�#r�ER�UwV@1�2�)E��%Qܔ��u��ձD���$.(���܌�{".�^�T��V�|�n]Z�>�ܾPӦ<��]�wF��8�%D/�tt����7BI����
�rK�5 Qe�䊤,��W'��)�����~���R{���<�U䰖�6���W�N�D�Hy4�	Fb%w)C�������Rp�GXشQ�B���Q�g__�:���B����W�j�vf$��SĄ���D�r)w�X4+ǭS'U�ͺ��;`Y��9<�+qH5��4Xk��m�VM�����rF#`GR�W�\lJ(u���k���B79����9=J����b�cti@5�~w�id�n��yB��w=TsF�M7=�D���!R�W�)��#���I�ȇ$�}uʶ���L�����sѺ�M���DxO1>q���i�p�bÚ��5���;Bˠ�7	�_�H��vީ5�;RUkT,��f�b6*@=��N���kZ��?K�&�n��t�p|m�u�pj$�������Ȏ�Y/䅼��&�5�/~��A1&� �	\�����ø�F���t��{�����u��R�ɜ�{-�#4S���6�vbR�,3m	�!��V8��/ypvP0S�ʇ݌�T#K[�$2.V$9����G�00SnwE� *�S	��[[u��.->��dƁB,^�C�X��%o�\H"��)FK���Uz2�~�(�x���g_�jD�%�;^��C�y�[K�G����!���XԂs�G�a[Y��S���N�N����������v�;�2�>��Y`�O�֎d���}W�ҽp�,;��K}_b��N~�P?��f�[!͚�=S �e��+r�L�ڶ�+�^c)V+;�RQ�	��	@-XY{y�y(��4�>���w9�3�܏�$�K�=:,�ϋD��<��YZ��Ss(�ظ�]UOi	 oWAE��l�/������i��}��s@��0�9=�)r��5,5��Tra�c���u�D�m�q�,&N�m�m̯/�jYJ��&���m�����B�/��R�e|�p[�k:��,�8����29?{������Rl�}�o�Wُ�����P���
.YҎ�s����Ӝ�M������/�;n���iL���������l6�$;����������e�{���T�ӣ/Or��h�E5���=�p �G>LS��q��V���%ka�<V������j�����0nk�S^�A�*�-zj���q���:v�M�z���,C�i���X&�۔0�����;��(1�t��A_5��o�]�KrU�!�����@*2��&Ą`�Zj�;���E׮V̪=������$}�l�`�P2SS=y㙊7�c�a���i�0�Ė�q��85Y�8Jx���Zÿ��:��KO ۴�(f@-}�)` #��7f�U���g��S�4Y�Xk�,��v}��ń/q沌 !�XT#�����#��V��3l���O���e�L�"{du�pa�[�u��l������3��Z�l�A��S�9�#62Ӫ! =J�S<�lj�bV.�iX�&�=!��՚�@5��a����X���[��'^F<� J3m�@��O&k��?o��x�u9ꑚ����(�v�-��,=~�߈��e�P��Õ(���6̹��εP�
W�(�43�K����`���I*�>�@X���Ň��+�]q�lD�gg0x.i��#
L�L6h/��>p^�� y�d~)S,�3c���b7�g�r~��D��N��"�"?�d��o��'��
��A�ӵ�[�S����$��`:C��1U��}]^�����ű'BQ>:6Ӗ�d�ހ��$Wh��u�x��e��c���ޡbƾ�#�|'�	��E2��>/�@%�A����`șds"/��k�+�b��F�8�����> @ ��&b��� ���A/K�������Q��1g��{��'����J�@f�kV��Q�)(p�ֱ������H�A(ё'�pP2A6<׼'*䓧Ȏ�aI�*����]��ROʸA8��.�&�����^���*\�i'$x��dL�%�����i���"�� �G-mR������%s[��t(��Ų�e�F{�T�UAP^��f#�F��8?��B�� G��	�s����$��"N�"�96�oUD�#�(�� .nx�h�B�}U�����d�t{p6�ۜE�Q;�n���-���t��fV��xE2�H�F�jF��)cZ3]dґ����1x�wUp��hv͒�K�<����/'*��;��&�Z�tXA���8.��yyU;���<����y8��R�z�aV'�� �J��-ӻOCh��z$<Վ����`@d���^��,�[�=/ &g��q �=���a����6<�k���[#SO�c'�={Q
v:��Mĺdƴ�\��� �g�nx���p���޺L�?�%�:��bY�c)!>4��Y����X�������
5$��c{���s;�3��=���V;<Ʈc��/�)�>UH~>����^Ơ#��a��c�Λ*BZeK@c��F���ĕ{a��^�i�zqWF�ϰ�@���hn�����Z�th��+��|G1y���p��_]���؀:�ܵy�Vw#5��L��T��5��1cF��e3���\>�L�𹂫�yPeve�,�%9>4p�[@�J2b�� �̳-���!��~8�y�%�_\$�I�K�<T�WiU�V=8�_�-�B*�,�.FG�Ns;�}��͘��wJ�OM²���fht|XO$_� ��(.�@X�a�����\K���y�Ɂ�wZE��؅Fx;-;�,����]�d�����+Z�� ��s�:b:��{���5w
c~�w�0x��Y�����s��W�K�@t@�6��F!��/��z&/y������`<���M7K��� ��)F�;��_��?>8���t�
�Sc���^��su��!��q������5�&�����/��E�.|;��Q�,
e��9z�3��5���c�9D_��+$1�����) 
��C��-���C`�پ���	˼r��SD����2e�8RyE�>~���9�
��9�}�[�u�r[��k:;J�
�+�[1��OO�z���8n�_�)�\)W�̔7zT�II���/\��{���i�^��v3�6F�2K�� Y�ӎ��y܆�%ޑ�ҺE��:�:h�����T��cФ�TN���u	Gl/����Xᅗ�Sx�6_�þ�M"٥b,���R�Op1.��^|�FJ�q�G�6����s+�X��P.����"����&���I��c� N��6�6CBϰ���-џ��bh�v1_i�&�%PRI��	b���?i��X��wZ�4e�V������N��OHڴ���P���@j��
��'�/�=�%��+p�z�s���I������m{Ʒ�1�uΩ�u�������	�~9!��^��P��â7]U��F`�]%��K���2T���������C��Pu���$��У�E�B�/UԜg���Y�ߑ��t�&��t�D���lYt~ԥ�4�K+% |�t���>�ܸ}���cmL�i�����×pK��.J�����j�aB�=Y�� g����#+j�1>�NM��,Ma���	(��l�F-Ac�L�U���z� <e�;D
x�!��k"�z��'Z�*f����O�S'I�'`����� _��Vn�oߧ�
)�sz�/�t���Hk����0~�ӧ�Ί		���J�m�	4 �dN9E�0�'���Q�9�2��Z���p%�оھ�*�5�]� �1�5�����R�)�3�2�,�pU���/.g��Ӥ����o�Jm��i���{1�ՏȧŦ�c0��i�N#���GM����`(����o�#�@��Mr�o��gGAGC�K0�{�|�"��U@֜�eK��iI�(�{\<� �?t��}��u#M�;��edv���e�.���Kn-e��
��<LO!K0�E��WL��z/ey%�˫�S�Y�*���,��w�G��$f���f'e����@��z`��m�T�����*�y�i����@J��o�W��$ͧ��~�0~W�T�[�i��p�+��������q"�^ ���5絏������\mf���������;�~�˽�ܞ�G�Yi?_h���A&��`^�M��Y�ɸ��Qv�� �`/����=�ꖲN�ϩ��T�Jw�c�bP,�Ʊ�	�/]y�� ���"�R��.��]�];8$4�ESV<V�,��G����2��FK�z�qI�Hި�"äBc��W�G/���nS��cdخhk1����,�p>���"J"�p	�8o^��u��F<%_ʥM�*���O�D���f�[������!��o�+:C���-2�c��rڪ�a�/�͋o�M��G��Z�ia��K%$`c3��b��wz��X j�k&�k�^� ���<�����s���(O
��$�m1��B�i�|����)�xj2{�q
��h@_w\�Yn�q��~ņP�z/�@��b�S�,-���Ƥt�,^�q�D{� �\_�V/�Y��?�>|����F���n��G|;p�������h�,X��\��9g�G@f�����F�`'�P{Z�4)a)�w�q����*���x����&}ڮ��ǐ�6'��͆c�c���O�~T�"0D�!?�#��ۈ��4�:��w�d�R�x�� ��I�xUK�.ҩ;�T�-:��t��'���B����^D��H� K���1oF��2��[
�B��=��ϕ�Avä=o]Ms��J'����5@��%Vzp����(?$8�9~�ぶ���Ylab��5GK�a'��vR���*D6�g��U���V��λ'�(�������Ւk�-��攳� �g��w�͛�̋c�����B�unR����	T��;Lh����i�\��:Tac!՛���'�cc�\��Z����[��@w�ݲ��B���&�Q�=*&�ؔ���U��>��I�@���zg��w�/|*����T�n?��F�qc�,7m���Y��4{/�|3<�ܵ�1��g�{n������c�Z�'��h�v\&e{�`�W��&#�0�������
�/�7����j�y��xC|&�k'�ld�ҿCg�b
F�d�`=:�,��	z��˛x��)Lm����)3��	�ve�^?	���v��#&LI���p\^��q�84�U󍶡�����-���!��[>�sf(��N�(a���*�R�_��i�6�OsD�(����Xj���?Q��P����6��T�I��:9�5!�U40NQ=��B��YBb��u�"]6�1��b<yHz����ҿ� �Ց�8.��1������f�a�����~���ԓ�|A�r�Xrpĸޔ��x����K�-oY�Qi�Ħ)�:�X������I�ᎌ0Ҽ��(�@}�%��|�xK�#<�?�&�m��ÉT�)6� c�jf���\���]a���L��FGdA=��轭��SЍ�9V�"f�Zb��V�0��R���h��3���"g�����x�������c�Y� 2����6K�~dB�m��'�#dY��M�u�y��?w���z�X�&^M�!k�[�\���������7jP	=V�{q��h%23O�\f�Q||MeWPk1��YM_�pO�-�cu��4�\#0O-G+P8�m��$(3|���U~j���)�M)�����"�.G\��5vτT�Yi�J�Uzи-�����c�JD):�OP�h��x����M΍�wW��d�� N�枀�k�t<ř#�{��6���
W�/�� �a��mÚxCW�≄u��%=rf�;"g�Xɸ���Ag�X�)�B�qc!<f��c��}>^��nk�yn���/S�����h��q��/���A����r��W&My�$�r�oQ�尜Zˁ"��-��,�9ף"
�Uh@�Q����
MgK�����9����[����(��|y�s^u�������B� ��6����9 ��f'ל���w�9*���O�(>6�$��מa/aa�ۋ�a��3�$1�qF� N*�����W��T��!�K^o3N_)�kF�뷥�Und� ���N��	v�q]l&V��_u��x�P��ҋ��Ȇ�~)G1�=P�a�A��^������Ț� �KgX��T:����g�D�7Ʈޜ�*xs,�)4���ǆ��ƴ�of�O@�g�s7�'l��3%6�����p�F��41C�|KM�"<%'=D�-==���j�;.�b��e���qY7�=*�!�$N {�`>H�64E@�ݡ�U>�hN�ZEg{�\���*ǥD_��`�享�)�|W��^ӊԺ�t�Д|�rOo�<��P\!dc�D&�#p�(b,ಅ�\���X!��������v�2Xڃ�{W;eOug�Ʌ�(1p���'��'��޸m�&�WG +�~W�A�_PD�����~
����s8�j{^9�7#��z��􅚛E�M���)����::v���R���ٰ�4,Y/��J�O��w=���%�^}�I�lg��rd S���|����~�hw��(� �xV��k�v�>���8(P$��[�E�������(����sئ���a�_f�E�w.M�,ͺ3�o��5u��?�����w���t���0�	E�5�3�]�a򂢍)��^J,���"e����]��h��\AVT1=����]�$�IGt$�+��N9�[-܇(�s �����i	]���5SG<l4�� n���e#�s'Nz��#�����'-�C���@aG;R׏���Y�[at�_���}���}Iݏ �b�����i�˗�l�7y�F���G�P2��;���+P�-���.Ǆ�9��em��'���Ʈ��-�e�����8Ne���`{�� ���bo?�;��\k]�a GI����l�K��:��}�����>�����ݕB�Jᄭ��=��1j�N���3��7MD�͍W�u�9�C���$p���E���!��Vu��l��,/|��g#��F�
S����-${;��/!�OA�����F��q����z���7�<R�:�{�}��a%֎`�Zx�b3�T��� |�rf|���vޜ��yK�3�p�ߗx�[�"pw�g�j�E&LO�n��sN�@�JTMZ�/[�4���D���2m::KF�xhIZ�+7/N���d,�Z����R�pl�`���`�sU���F��3Cf�-x���1�@�̨��誶�%��^<��A�����'��o�+�z<eq}�N^��� ��%6��03��0�~�<+OP6nd�1-P�����)��VҾ���v�-4����o������J(��{�CI��Hw���=׶��u�h�9IfU��E"̎�a��|�Ň��E�1�*\A_���)N�Z��[���*ܑ	�\qQi����@��X��w�bx���r���t<*C�s�������Q��#�䏳l��ߎ��@?P"���6��=����An�f����)�~��:c3`�̌L��p�( �~ L�{W��s
)�k"j��J$���V�$]���1�G��{�c��|:<h��֖�>3P&�YV?t ��1ٲ.rUŰݠ��蹄�QS���0m�O����g�&E�����{z��K��
F�Jc�����Hĥ�OS#C�V[�i���m���t�=����|ig=��}��,��Q ���i�q?dJ�q3MѣbZxd�|N�'^�����:x��g��by232[[>�6��_�f���J����̜b���5Z������3�~��2힎-��"�^%�2�Ʈ�;��C��?��3W�����]��$Q~r��V���a �e�e�k��T��Y��Q��;~� ��d������O�ϢV��̊󉼹�9@�&5����
�tr>O`A(P�Q!�5J/T��K��:��rjeIboo}�+v޻�g}N�Kk�`�:J7�����+-�<ȉˁޗ��j������zDH�� С3Lw�i���#v��xmB �+�Ɍ�>��x��!V����@���3����/��8�����'��%f,��t�����r���ڗ-U����Q�b ��w+B���8Ce���Tm�nD
%��?�@�1p�1��J�BRA��W�kاD`~�TF#`s!��'�g�(�"��f�����-��x�K.!���
_Z�����M��F�iRi�]���^�.���7� �8�t�+�Yӎ�Ob��H�~1S|iuowrh�I�t�n�C9�ؤB�W�>�]VLD �r�Vd��^n�+,1o��^���"�_Q ���ˌ��Ö���B����^��$��b2i�d��J���i�:�{�jg��Z��@B�
�.���h~0����2��ϓ�,�s������y��N$��y�6h��VueU|~����\�U_z�km��_����t°W�)ZE;�O�I�����A��������m�%D(V�M����5��<�po�`�/�*���9�?Lys�㎒�Fp�y�N��׮�`�r�w����Uo
�^�nԱ4�u�v<����Y;���t̀h\�,uz
����qwKC�q����G�S��U*a����;e�! t����5�-m�)�P�)qȁ�q�귆��ax�$Fб_#��0�H���j,Ǖ�5C��(���잂��>Su/��s�ß���Y�ZL[FN|{�pٱF�`�c��V�mǪyq�;h�h� k,x�y��{_��q1�d����}n�эj/b�o����2���M����0xwnF�myf�WcbW�5:�ؿ�:"����(lR9e�����kyZ�p�K(Vǜ\�y�m%���K[�D�����3Z�]P��%Ui�����1�唆����_�I�b�ñ����T̻��&������Y`�1�뒯j��5�!v�vWu��]����;�A�$]I�3�l��������o�e̘	���Vt֩��!���z�pH{\��-{��+@V�dc�u�1z[W���ͤZ�*�c ����%����W�\�"ۄ��yH�Ul��n���bGؘ�F'3�%ur�����z��w��C>y����[�i�_-�S��|>�%�X�U2 �Z������{��gZ���c7 ��J�1��d;�Z��bH}�q'��V㺃�ׄw�Y���q�I��m���%�%�7<�����������҂�܄I���!��.l�h�o�詰hn�؁�jh��#�r�'{��mg/d�1�5@�U�=$� 4Ϣ��u��;���V�>�n��Ӿ���b6B�Ѣ��$D5�_�r�	���WF??yV}��(�*G�X�8��&7>cr��=��FQ�#:^ͤ/e���匷zM�(:�zeu}���}�4˞����f][����(���b�SS08��Sb�kʁL�R�&z��h9P����Ǉ�~bm�b���_�b���1ᵕ�yLbm�#�ӎ��d��q����ƫ����PՈʫL�<;4!8Bd�>���3����(%/bS��X��]��*1�MkϬo����F��x��P�'�ػRY$+�,�,���'F^��sT0��H��$#y�A�W�'f��-�/�׳�����*/�����~M$���O~�b�燩R����H�}���۾�Y4��^ݽX��&�7s�Fv>ؗ�j�F�6�^��~:������^�\D�'�A�r_8�9�=^Akɰ�1��L��M�nw.�B���U%+���/8�ɐ�<מ��	�W�p)��Bv�'�����P(�����9��S�iUQv����"��eP[�i�3�n5�zn�M�z��И)�,|�Mw��bH�u����O$(.F�.�e�$�Yp��׈ND��D����@(n�D������'n��؛�p�C��*�9�0K��ۂ���v�"6ӊ�1��)�P������Yx�����L���0%�D� H�� F�#6۝���0�F���S5<�tW�%J?�wv}�_��RD��e�Q�	~O�G};*�\�+(Jevˑޅ�g�����=c`����s��)��z60 g�L~F�74Vx�#�:�g�wOzǱ�%�v�RY���[+���VO�1j��3�Q�C�X��;��3n"��~t���]��S.3�[�[m��E<'`>�������D����߹�[C���(�5^գ���M�
&אR!��B��\�� ����#1�`��Sd��!{hd0����w��t2�O%`��鎕Q���nF%Ԙ�Ǥ�����=�y�|W���)ߗ��GAG^r�}u�h��&&����^�>k��Q��c�#��O ���:N�W�&1���޴K�O��r�+|w��&I <�W �J伻Y���{V�r��E�6�.��h��dYJ0�ö	��}��}{��)a[h���*�L,Е����Y��~nj�_�"������pmL'we=
`�j��a�
:�U
���gi^������Ʊ"~��@-,��ʢ"Qʦ,�>�����Z�|�*B8���%���t�]S�`'(�"!�% 7�:��$�V��eLr�<aV<��r��+&�S�sl`��XX���Yu�w24��G��"﩮J?��wD���Z#o����p�s�����G����ۉ12�'4���Aڨ抧��V��w��d|Y�� �=w��S�D��\객82��U3�d�Gk�y���ѝ$h�S:7۽�F��`�d_�V��t�"�~��ǘFݤ\i��~�l1�Տ4�@ӄ� 9(|	����4��J�L|,_��D�e�2,����
���2By��	"���N���$оq_��_ ��'QIo�d���S�	#�v ��ڳ�x�Q�M^��Y��sk������m���i�2֗O��m�;� ��'��YEJ@��̺h��E��n6W��%����fP]697�1s�la�Gv�6.YLݹLז|�A���F��p��d'��h�3�&[�A���FIS؁��]�����Q���h��h#�3gX�9ڰs��<���~kA�����N͌��\�U���߼m"1Ͽ�)�]J�'�R��d_�M+�<��T���{R��R����
9=��jb����N�Y�i)���3��l�F�#���9:z{9E�Rh����[�as�9�r*���S�q1%����D��D�U�,F�?���Ԥ��;`�v�N��g�jX|K�Ĕ���MPL/�i8[J���6I�hk' �^�N�I/^������{�����{��a�{�tC*���Z$�Z�a�gV�fwWB<�هk9ռ���������4F�ڋ�4(���[�[�6�ȏ��G���ī:�o�s7�!��3�uA�Q��/��/�Rg*����g�j�� vj,�'�����J���:鸐���b&*Ӎ��G��zxQN��꣧��9�Qy\��͡
�-|X:`��q��/0��,e�j�)|c@	R	��Zn�Xl�p�v��~�ֶ�Xߗ�!ZKg&%�6�Dj@��tjP�m-$`�F�S��m����1= ���^Um`�:��y��FI"w��Ѫ�P����a�)��"D7K���M�'�b��(��D
��]ד��-X�6���.�}2�t/�ӻg
��T����k�| �Q���x6�=#Asr!V0H%��,���,��mQ.6Mb�1АN�K����l��� b�S�J�'�P��[�*ҋX(h�@�s:XL�tP�����sEc��b*8q�5��U����)�3��,��5�?����B�M�����ִ{����E
6b�M��خH�'Bg\�L�T���{I���1����b�*��p�k�b ~����*�-����87k�#���$�wW�������{�&3�\�_F$�v��VG3��"�:_=�����������b�f����?�=s��QM�w��q#�ivD���☰�0짩��0��<,֕<H��LP����a^�ZW���D��*Uw�R�v�����u��}��$B��:'�1��)�r��b�Ș�Q��`Gi}��f���E�5Y�yP7� ԧhϾ
���xt��	H�􎕨r�������S9��tl��!�R�4�k���H=��W2z.T˨Cy�+�Xs���k0􁂏�8)�2����M�r���H���w�*�[�EP�gZln6.����KJ2Je_�p�a0�����gF��9}�rq� ������>�Qvd�^9�dA����E���QɃ����'����N�Ā]j�u�C<\���K�km�JtM!u��Ew[=����y��j�f��W��4���4SY��n���f�"b������l���%���~���e5���
ܟy��!�o�&�Fָ�g�´��8��z��IW�K~E����Th����io"�wEk^Qd\<.|�5�}6�v���ܾA�u�al�F�6�|��t#�Θ1�d��]�vٞm��1���m�+$K�4��]%<u8�ٺ[�:�J�c�le��/�6��0��ly�HNM��:��g9 "5O���~��j���,lWpU�O�K?)b����C�_1J7rW�}��79�+2���n(�=pӺNn\���s��p"5AZ��0O�;*��� �5清KZ�*�1m��LZ���~��Γ�Eλ��X��������Z��'	�2��G�X��w�$��P�Y�!è6�&ȔSSV/���8~l���t�	���3�,�XM3rJ]�T�`��6Ad-|IMb�;A����j�;iN�5��v��˰ݣ-�\�W��)U���'Y�6C����9�E�����E,��=0�?�)}4�,�B'���8u&Bn���K���0��u��R{��j��g��2/��ܮ2H���/|K��a��������p� �ȹ8���p�z�i��8!�r�U��YAQ���k�O�0YN�t�\u�����ԕ�ۑnD|���r��\ �B��t6���F�Ilr9e�	30�`d���F��G5s���V>8�]�9CY�����I{~���_B���Π������>^
�Hl�?!��h�8��Dg�o���.�˙e]�:����A�a^�+�˵4A�y��/�(� a��(�HM��q���wp�мGX������Q�1�iF/r*?3������s3q.��@�5��|~� L�E���q[����x
ə�|S�^Z�2�-#��N�*f1�aJ=v���3JA[:�ޏ��v^C��/�ъ�����ܲ�t&q���ц][��Q�oMYҿ�,��%3�{�-��h̐x����u^ع����$@J��Q�dZ����C������9���W4R��ڛ��lH�-O�s8c��|���+��9o=�ZO��5��B�U�̺��!�9/�f��H<)�v��}��G"�ڐ?ٵ����e��^	����BY�|il��h�Kx�d|�HU�K��,����7<�2}���k����b�,�hEU���f)9V�8`�@-p���N=s�Kd�۷c�u$͒�@s�����Zm;�1k?���:�G;���v袜?�G�$kD�)-N�����K�*1�b�m�ݗ�w�:��Z��ֆ��-d�. W�ʴT�����&���4$T�CS�9��zq�o�Ga����<
M+rHc���Rd����Y_/��`fDd��*�BtD��G&?Iچ�.�<�s�=��pUaP\r�7����1��w���v�t�����>�d��ǰ_�y����EhGJU�:��C�jr�VaP3��
����L�t�`��J9Aj.���U[,iᛡiZ��O'��_-�Qs;��B�j�*Z[��M��Dߧ���+���^]��R�/���gx�z� E�>j(��@=Ĳϴț�Ŏ�U	s� 0#0�;�n� {tT�(,�����O�|f��[i[Ϧ�������>j������w��y�:�	ҥ�I{5��M���2�E7��ow>+,q@�8�o <�
'�=�<�M�a�}�ҿ�"k�-'�ؙ Xo9�8��D�.'�*p}«����-i&��nFN��|b����8^���XD��.ğ�dA~d�>�M��v[������'���~�L���I�uB~��"S�^�M��h\�#��|����Cb�]��3"ƃ�w�Ć�q���e���x/�X�~N�Cd�}�E�]���`%~i_y���n!�b���5�u[�^�h�*쉨��Wx�d<l
�Tɮ%u��K3�J�b�m��Dl�ڒu�8�2���:�XˬV���$�ZXgž�PA��z������Sö�c�$�㡜���N�X����T��~��|��uoDG)���bR�o�V�3r_���+i��V=��Cn�+�@�'�L���;G��&x�JMs��R�~/���c���L�1��\h�d�t����  �}�+�0�W�I'��;[�A͎��|�Fx�[������)��P��M���]��Ö�J0LN�0]>��e�Mq����V���Q�V�~`��iۼi��.�:�\��:�A��y�Oέ��q�QQ���TI5c�*X����XKW��͜�Zr_ǥ���6�Z^گi�i���X>��Lg7���;'�@���o�ʤ�TQ���t��F��΅j�"�bl��ߔ�8���? 6��T�ȮZ�DL����WI��^hIuRV��{N���%uSC���6�S	�����PBj
w�6t����r�8c|�[2x+�Z�1~5]Jy�b�fOZ+��Q�M�, �{*w��4Ve�| ���d�/�f�gd(�֋)"H�6�"/R��]���#w:�'.�?�A�B�[	\(�� 	l���}��sy
4�Q�<W�YE�� �5�s�1G~��怿�R�Z�}�s�[��$4�SDU{�K�r���.�Y�(�[���6٨����S$VL�����珨��d�.�c���{�&���-���.س���->���TMy��2��o���[E$t�� �<Tc
��)��"�)�� �ؤ�P!��L$�8E�m�5!��aR79(�G1n �B_���ȷ��J9���U�t���\��i�j����hQx]��Q�36�yv�XY���4��O�@fЩ����yM�cYްf�>2�`m
Q苉0-*H�����d�(Ѳ\�Rp��X�0@9�Z�ш���Ξ�GJ!��F�_��UR��i�7��[ah�t��7I���#(%ޭ5#T��"�����5ڢ��tgΏ�*[�QrB+r�!T���F䖖��Iԭ��S���貶R�
��SZ�{���Z9����{�ʻ��E��U�̋l��^*/�/wn�G�,L��x a��3�֏9W�S�~@]^(>p��ހ+�&*�ؾ:�R�d,��:κ���C ��'��@g��}us+��6"H��3Ko�{���P����o����) }����=p?�s��d������ǭ��x����3#;��<���̓��P/���D6���R��e��n1g;��,<���}�xq��E�*"��$zZO�w�E/�vh��>�H�sDn>�E�?7X��]���̷�
P�*9|t�4?�
����XZ��}ۜ��e�AF5j�<c�Pкt츯:%:���'���v���L*+���B������u�/�^�kU}�2������A�F���Z͟A���(���Z
���.F������=3�uW��'$�])�ޠj`I�5�v[�d�2=��G�<�f	���V^�����e�����S�WK��(xhi�B�[f1��$h�i8���݌L"V^������J�ƹ�9��#PG,L�����$�2e> �X8l8�:�������-�T)Kȗ�s'i&|���q���R����a�*_�	�iGqk�礐�%|��͋3 X�k�y���̴�RVp�d��Q¬�vx���ƪ�m������]�Yթ�?7W1)���! ���@)���Gh��OS�1�x/X�T���dZ�O�Fpa����!�%!�;gy�N�_���_j��h(7��fELD��
twf_�Jj��n� Ɯ�ʮ|;�mc�[%�?��������*�f�pB�]��4�>����΢���g��$+'��,S�t��W�p�08,r��y�����I���/*N
�q-%=<6 ?�� .*� ��Uy8���Gŵ�NWU��Z�UC�9��7��5ibw>F:���,UG����=#�8�j������4U�����/�Y�Z�޶B�O��t�0�e�TqK�d�mq64� ��#�����U�]�J�	C��iÊ��_i����T���<������m��H�Lo;&���N7�>�����c
"�V��v��ZzE,
�mZ6J׹��&�'�j�*0�VNTKr�~c�9������&夁V��O/nz�S����6�����u4ԍ��andG��Ĩ�T���$]�c�kWCq�'J
NJ�,Qv�F(��5h���*�)W�� �ի:��/W�e�W�~GFb��;�<a� ����D�N=������SExv��95,4 ׽r��lj��h��	A�d�K+���eDkʖ׊��Y���@��1V,��d-?d���i��%7b.P�v2&���5����[�"�� �)\�`�`	*�0�I��#�O��@'�۳|�Z_tWT���6H
��r�YvH0�I?P��8F�N
�Ej����gl�*��	F%$���J�t�c�1≢|ŅX�
�� ah�w
�1����f�I9�~��v�л�m*�}�a�I�Y,�ێ��@���א����%�b��-:̴h�IH�<^�>��k��&�͝@��3��ޜ�My�x��qD�]T����#hz0�U�6�k
�3!%�`L����T/<Ζ����Z��;Bf/bdblx%ú��ܕ��D-�
o�V1[NRH���<`F�,l��gI[�+���|(�XM�IN5��^R�.�@?��Yƛ���ʾ����jO'�6�lC�%�b-�wl㣖^��ګ�G.)l+:h?R8�����=`I�0z�O�.% jb��yd�:HZ8oB���R�:���ЭU徑��3����L�L���_5LM_E��AP_0̝�����nƠ���K|U�R�����3��F�ƿ�C�f�RbI~�sg~#�nH���5)f��}��: �����eƘ��J���)�����-쮠�*��3�̱Wm��oU��vL��f�q����0�Em�y���%E�r֣��<�n�2���#xt���\E��q�K�;�댑w{�."�3ǵS^򎆜z<S�sp��/����N�%������.��/%:��Zˍk%�����Ŏa���`���f��v�瞢�*�mY_�">�đ�My�Q��	�eH2xs �'�O����zf��v�fe51�Y>��c��Ԋ��#�������k#�5<�fl�����r�&@x�H��(�Yk��9����ޚ��c~�x������kʞ=�λ��3�u��a/�/��{���m,	��e�(AsN�FY��)�����@��v_V��M�9��������n�^Z45�I�k(���	mq�P�͝G�^A����6j4$�D-Jp�����&o`13�[��X��',�yTX?��q~�R�.�]�#�*_(z��ܙ,�����x�LC���=��8~f;<.]3��Q� ,� ��&�����m% ���_�Π7�ލ\ ��M&��c!5�7�p�W�i�&9�L@��3 g7��V��&�w!���N!(n���u����t�Xd������&0&�y'�rC�{�M-��#�Y�L�O��=����"|��6�}u+��~"��D�S�O|#6��KC�t�=���P��P�����A� ��	7��o��q��^B�]Ф^Aܟ��\�_���q�Q���� �B�a(Z�D����i��Mo�(��P���<VT&Q��y֓����}�ͣ�����������B`$l�xI���I�9�h��޽~��{p԰��;�K�P��̝���������ƶi!�j'���Ŏ�ٮ|K���p�FvXi޶\�P�E��)P	�N�o�fZ�K������0ը�KL9x3�QE;x�C�Ԟ�6ˇ>�z.3�Y~�ܩ�ndc��GE��Q����m���(n�A9�F�Bq����|j]�	s��b}�x5E����hly�]T�����1��n\R~s6�vR���p�*��6j����!~&,� 	�d����N�����	��`h�W����.\�KdVs���B㛙Hb^���4E�ٱX��VEȣ}:57�4�pr�7���@eO��S��j�_s���D�[��Tڼ����Lm�8unxp��}W�>�,�Ӈ�^���u�$�NӪ�i��D�++j@��?z�����\��A~P|����ғI�c�o�҄�|߸��L�����ǷD�/?�JܟE<e'�\m.��������ŷp(�|":��N��2���:X`�!+���ܘ�u�J�װ3��%L bp߁Zĵd�`�$Fz����wyWOW����坡6��.,�qٶ�;Fz��'���kʂ�����Y}����i3�u(�P�� ��F�/��3�_f9q��ߝ�i�Pb�j����(a���p�op���� A�Ù�v6���x>�<,�������&[���
"Ӌ{s���ħ�!��ެ3�s'�߮߭��M]Xb��&IS^��-��Ϥ^J ��Q�¥-�&�Ѭ���F�vx.&Y���?��W �a�9,�+�H�	��!�g��L���]����~�3��f����5-͝>���n���j>�ҏ]ưw��;]YY7���C�dOW��(tĈl�������%�]�t{e���Y����EF-�5y����B&2b0N�h���u���30�@��?�Jȹ;�A�߭��5 ��aε�\���h�^��g�{�m{�����:ȿ�3�e�(���`�d�[�\���Ej���/�X����X�	F �c�,���׮���u��R�ȒS&3J���N1+YM�jJ�x���W
�z>�"�0��W��a�_G��3���p{�wz �vc�N�ĵ��+�8^MKͦa	�2d!O�a�KT�*��{)+����#�����D��=(Tg��Z����y@��.��*�� ��",T���ԣ�Y��Ҭ�(&ѽ���TpU��۫�K�y���i\��!�F���W��t�F�r}�n����W��ZYԄy��w��S�掷��Gpe�tY{�h~��� 뮐{���?�쌆��8���7��VS�;���I1��������͆D
j4k .�=8h;\˸����-�겈�C�A]~�U3��̵��jT"���/
��sxg�&�EcE<ܽ b�R��6{�-8����v"dС� ~<��&!/�j��2��1�tb�l�c���]�>'BL�^�m��u��^�3ftF�{BC���K�Q�3�CJT����IO� I))k�;1 �:m��g�#����+ؐV� �%��3M�>|D�
C�ց&ZQ���R������J��L��"�x@�"��6�$�n���8cD�P�S9��E:y�u)�]�����7֢F(�@���A8,��F���Q$����gL珎f���Y"T��2c���n�_G�i�@�q�ŒT�&�� f����yđ�.�"r	�f�#�ֵw���}�j�óG,v��b(�b؍؍�?Y�^p2X�O��� ��?H���L�ŏH�:+�V ;�[�����ߎPZ�'  B��t�l���`"���I��ݚ���^4���z��S~~K��,�����Va�72���5r|��T�t�ۃ-�,�cd�=���m�dL�i�t�|���sY&݁("�Gt�<9��]��!���{�m��QFp#u��ȱ�M���)	d�:�7Q��h�;׳�3FQ@B��6Y�}a�����Q˱8K?�߄{1��G3{�Cо�͏,�j��t����V�4+<����݃׃�$|ǚ=����gCd�t����25���ֿ�s؍��,PU����m��d��S�r�������'��	��vg�,d+,��K�脭�lg�f &<9�H��g���2�0Ĳ~���c�\��T�%��b-	J8g�����HQK���$���#�OH��"ǧ�sv��Kg����*�9��48��*�<���1���D7|V��	�c%9u��3���fm�����Y�{JGJ&�G��S��D-A1C��`IV�I���]>�H*Ɯ���G�滚���)5I`DʣH&	������umE��ST����<<��,��d.��x7���@㽽����b{���߇V��!�BLLQ�Z��?�_�6�a�f�J�l%[.$3����+�����wWe���Υf�m�H5Y��g�J��5b��n��Xuz��X�ʼP�N1>��Yn)������o%$|��?0��Ų0�O�1�Ú>�[�O��n���G��ym�~K�ߊau-��52�8��[M�t�XS7?o;&��Ɏ��w��)6�tْc�}|0%�O���GW9�%I(����y[@B��%�Nj�D�AL��� �*#ZF#x��ү����HE�)qqG�+�w"��˅Q��_n�K5�6D%ٜ	̘@�dbbͦ�S���H�(o�*��@��9��̨@C~��2����}j��|�D���l.�� џ��~DN-���fiv��\�
J���u�;S).p^��k�c�E�`��ˁi�E҃_@6T����
N���Ku�����3�Q�ȭ`�e v�t�!��y
��wo�D��/]X*`«�;�F��@P�z�Ϗ�Q�  ꜂�&�bp&n+��k��X��̂��R����ep�u#f	@(�^��ދ]�2� �1��8D�h�?Gyv��çJ�Y�c!��R�꺔�����K�"G\�Ǹ�`b���'Ł�]��=���W�
ꈓu�\������
�V���55�e�q�Ш��hZ��$�Y�kC��Q��;+us�m���Nn��6m�|�u��-g�I��9!�r��#��T��t #ud^<��د����=NW�yݮ���£���b�k���V~�G�v�,Þ
�Z{ ?���f�R���اYOM�ng@&���B�O��M\(���6w&c���_�<�^�"gy���N��S0�|��6xF��$4��.��h<�Y���(H{��d1��I�c�W1Z&)�!����Wo��$�,OU_����P
فC�7��@y�mrN�D�Uo�8K�/��_qƜkaq���
�+%V�a��;g�?[�m
�׈%Z���9����pxTD����[������ ��&��yr����, ��Y�3��3�%1ۉ�!��舿i�l*�=fA]�&�v�h3d+3u �>X��?�M�փt�=�,΋��PT��D����
��AU��CIa���k�� CeӅ�8�.���=�;�VϦ�Ո��G_�#�<��o.R�o��MJ7����(�\�[�`���JgM�������
�[������:���w�c�� ����B��N�l֩��{mץ�W��[�v��ϕA��}jm �j�Z��q������et��T��zc���(����h��f��u��d�����C� �G�	��t�Tn��rЀܫ3���u�C<���	�s�����L=�K�����5xx�
�U�Wj���h��CU�o�� ��o�I�F"���f�#t����:���ɘF��(�{PQ��{�L��IM��V�����<���G�I����~D�Z��Z��H�I�%W�$��Q:	=��Dq�!��±G ��uy��t�i8�(y��1��Ws�Pi]��M@bO�~�=�P�恺G��2}P�p�:��e���t��/�Z�o&dq������f��Ss]J��HI������ׅ�{��#�A����>kj��1_)3�z�l�u��[ᒗb�2�;ϫ���H`�6��t���Q��ױh~��4�(N�jd��:�}J����Uǻ�9\5HV��f��a�(�� ��������&�� D��/�8��KfX��c�����+��<����7�����>���LV���CE�����
$��v���D� )��qO�O%�rH���F��B�5�%�s�h)1�7��������G�1���U�$rV�v�Y%r�[I⹈�K�XcaY���x�qx��Z���dR)x��ܘ����A��֚�6R���hۦ�����^.�S��G:����!�q���i�	K��ʃ��)\g���^Ea�X:�w��8N|=6��4(zz�Hy �2�T)q��D)��)m��0�(t�����>��q�qc�'�OuG�����ac�3f!�Q�R�P�m@��tY%�B� D��u'\��{�mNq�~����U�ִ�8*��;$�c�& �?�)��a��M�؛ �c��y���D�e" KC�1�'%��%�ߚ����d�יպ��N�Ѓ�?�̨��n�U�o�$�">?&F���V�پ`dD�N/����]�6�ߊ��ֲ��3ϕ�(����mn�C���ҩ*�����~�y��m�����4|��b��j(jΒI�F^��K�dM{�lQGBv;��LY,2��dwe�݌�=��oЎ��}6$�\��;�e��0����~W����lq���5��x�&5������NWJB�.�Z��b�N�����F�Ɋ-�F�����nB0�D^�o��q��P6Q�Ӕ�t��D�9���q�g����6���)��X`1ʟ'��{[����q1�T6�[���K�1fFk])�2H���֐`޻��QZ����}V�]��KI~�,����5K�F�� 0�|QY673��O����y7���D�8z��	���x?M]��򙘩"�ٰ��G2F�o��'�7t���i���ou�N�}z�/-��ׅS���0n�~��D������I�
�d l5��nK�i����T��j�tu�/}Eh E/em��0�G1����C0�IK�g��/���Ϋn׉��hbS��<�G��;�.u��^�$�ԳS7�'$�M��]�K�XB]�틆�O7A�::���g4U0b7�v�?���<A=�4ˏ��,������%�{��ɤ,�Yt��1����"��D����ݷ i�lzdS��R�|k�lFT���P��\�B��X�"�#NIt�L��C� �����;W�����0����-)/�`���0A�V�L����8n&�
ܩ�0�@$�=��M��Ot�)��rs�ua�Ty�0������Y��rC�{�-8�^��������+"��?H�l�+�N�����W}l*�6�Պ[h�7'y�;��K+�J�@���E��S��# @d�����͋�;��2�!���U�Zs0��v��ѳ̭N�)Gj� �Q���71���EψFI諎?q1%��$:��q[��������:�(N���g͊�/k��`nN��ͧWi�ZbR`�F|�H���IMANK�t�%n�R�%�9���cy�' ��Z�"к*}��lQ�!��x�הƼTsu���Q����S�k�:�(�[�ԣ8��4%�R�I5�D��?.��ڕ���༳�����g@v�Z|sʧ��Ѩ�C�,�%N��Ǳ�ʔ�%�0�L����˲��w�K�ן�R-����G�����ٛʺB����r��N�T�ze���@��4~�9_�����*�7��q��N�(Y\��N2�t��Ԥrz��Z#V�l(��i��i$�����ܹ�%�m�����G�@]�X������c���u����A�{u�O�n�R11�!�6��׈q��T�
���D8�r��N�)��Ǹ>.��i�j���4c�DG穭q��\�䇗���}Y�D�kb��jO_�e
�JJw�d���?Ycs=l�O�7K�!1ȥ8=[��Ƈ�tғ&O�mA0�OS{4sEurR��(�lk5"��Y	��6�2y�EEv��IE3��I��K_ꡠ��h�ƞ��%���|Ts%p�DI"�uI=\x�|:y�Z��0�ƻ�;������6}f�^*L��"r>==���T�x-�֐���7��<LA�@�m'5҂ZaI&���E]�b�1J̅YU��Kq���yAI"bk��Ɖ���m*��[�CCOJ6���}/bA��k���`?W.^�W��dSiDT\��.�Rz�f�
���}��%��)�~��k�J\���t�֯Ř@H���+a�U������Ώׯ[�pq�p��~�K���I�������B`�i�э�#�y1X���PE-޻���x�v�B��B�EX�Q��в��l�v����v��_�Y'��=�@Հs:��MPP���B+IÌV�x����]���E-܆����<}	Lvk�4a�SXx7��`i�G� �o����$���W��=JG�_�E�e�t�y���� �˴CJ��4�/��� skd$�y�ɾ�0�k��uN��>�T�()ٖc�Y�/"#�]Rf:噇�A�J7o�N����T�
����n'Ǚ����LzM�!O5��DnQF���al��������l6��Pr+�mu�'�XrahΧ��$�b#�혠5�=/���>��|�]�]Q��aVz�xܙ��xb��@ �n���&L�w�[�>t��-�$�:��Jv��$�ˢ����I].x�O8[A�·�-�C�sثWÑ[7.��Jh
��a y�AICX��֏����j"& �� Tv�D����P���_�o�q�2�����k7���R�<�����,;���V��(c&��:"��X
�0��z��7��� ����J��*�����m��Qq( B��f�ݟ�[7k��qF)g?�md|�N b���,��L�~����)�'*���H�r5-|Q��N�ֿ��A����82~�T�����^^���D��Ii����F�ߢÖ�v�X��Q�������vM���axS�����rqv��T�����e4�2���	�+{O�,���ɀ�x;��$��K�	���F_���3���d`�s��
�6V|��=��5�"��Fys��b�~�Ɔ�nI>��\I�	��h�p�aJ��j=�S�$m0%PQu�=*&m.�1N��+�^P8���|�U|(��r}�Zq��GQ��b��G6r��z�ֶ��E�k	K�
P��䝮J�b��f�Vy���<��ͩ�57W���C�O��p����%ct�F��� =��b���z�X���.}3��q��l��{����⵻��k%���wu��"Hc$^��Ѷz�N��'@Y�Ю(C/@�Lñ�@&�A�nnX�D�2^H�AR�CW@'��h��{6��čG����߹~n��B��uf�&�)P&�5� �LAG�z�w�-p�K��&�`h��JMi��D�����S�)�k� ^N&��F���A\Q�6�]&��Xz�h��D@�@����d�Z�����bۺ�^�eF��j�a��(-y,9_����c�OA����iՇ���1���g؈����D�IB+X�(��U�1(z/�3����O9�kC�X�����վzt��2H ��צ��d3��+}k��|x�JNH���($h�>W������ M�6�ɛyI�����g��.h1�J���vCA(U@�ڱƢj[J<��3dbπ?d�0
vp��.ץ;{� ���WF� 3Ps����|�C����d
���i�4��k2^Ü�u㮒�U���U�+r݃@��θ�G��c��ɸ|.�e!Zk������JȨ�/�p0��g��w#�*��(�LƐS��(�J����ĭ�] u�5�����<����1̲Qrl]�ߦ8��]S;g�%�Ȥ��~i��>
:�Y����,����Ӊ�O��yr��wS'�Y}�ԺoL�Xԥ�V=5�J(B�B��ֱ� ���gAt�7��GlȚ^����c�+����N�� <Ag�ﰀ�TH�0}@C���i�(�j���|.�2��as/�JH�
?���a`V��p�O�A��F7a0�#��n�*��ʦ���!2�����_XYI��G�VO�&<�z� �����a�_X�p�B���Ɩ�#(ĢN~�:�W�e�cni"h^T~eĽ܎� �#�Ǡ�V�'���+��*�O�!��m��%x��Xb�g�t�iݱqk~�,����z+�L|Q�b�R�k�<n|�U����_'�E=����z��v6�K�WG{rf������(�4l������=�*�;�~Ͻ�r�]#����<�1��vhI��_�K�,�2���sp�:�q���zTɗ�e��;l�Q�Rb~m4�ƌ�3���U�Nys�^�����%W3a�*Eν�'�R:���f,�k�Y�t�;�l0�d�!|-�%�g� ���+-��V����)	�`ǘ�����i�K�9��+{r/���̖մq��k` qtv�1�ޥ��+͙Q��h�i`��\���������q���aC���E��~���+�8(K���1�ܷʻ��Wn5�A#c�����t��\Y��c�~8����90�UN���B���L��%��*���S3;�۵Q��]ʎ�f_��Q�d2( �S���#����T�?L~~	!�y��j����l)��X��+n&�
���s#�R(H�N�T��t�?f�\:�>N�e5C\W�q�����ҳ�a
�]���΅$b��쨉�);�XJ^MJ,�_��}��?�D�c(<��h馹E��}��T�t��U
$�v|�S�)#��h�~�� ���mR���}.�&����DI5@�+��b���<�:�;#�n�o�~���.���m����2�����w�����]����P��@�`��6��;⊥�d�!�Qt��6(޽\?Q]��x�ϣ�^X�_~��j����c��)�M��N�v��!Z���u�b.�Yq�D���'$�V-�lz�3z��S̮�h�W�W�5��c���O�����J���u�˪��:��C���B7��#�x��c�b��e�^�(ܳ8���@ֹ��͢4�b!�\���»[�l
�L�uձ����vM�7�-�͟�اmH�j�����E�;'������;3�~%݌.��a�d���C���Α��W���q2�ٝ�T�����؛��Wb 3��UDxy�-�I����M{�&��	��Y��yS
�Ncw� ��;�$�#]U��E�-�����{�u�c��5Bm��CA��?|��t��&$�Ō�b�!E&�֒�qh��߳�߹��:7N���V2��Ť`��iRY����6:\(����/��"�v:9�2Y����}����H�~R[��S`	����@�<<�ݳ&!Oz�b%|�ì���9`���*D$eI��M��V� x�	�f�)�5,�j��b$�&�0���w�RW�=�����{��_.6`'h5�%LR�y�^9�@���N�s�i!Ӻ�%=
����-Fe�I�tr���b��!�g��9��V�8�2d3?��_J��ra��J�[����Ñ }��h�;z�!�z;slwy,��]Qqe�'험Oc�o9D'�w�M5M���]&�/JNVB��;o-���	7����qJT��L,������5�޿��N�SH2ڍ��W��J���;�bIL�5���U���aOV�R=�́b��ߟ�1t���`��F��XE��qa�,����ꥳ����I��9�jn�0v�RرW� �J��v|<�o��XC50��wW �jc.}1t��ҫY��iiPM��軅)?�¹�$"����hsi�>�=��av2�U�}�T�A@)��m]gQ��@�{L��M]��r�Zz�P~��R�e.��9 �<�^TD�e����K]��˾a��@��-Z���i+�L���CÂ�)g��p�j�,*�8b��M��� 1�7��a����Kpe��Ȱeׄ�)�ݥ3��_B ��Nd��� �r`d�h�#/:�_D*w]u "[��y�O	�efh��$�T���Zo��ߘc���sCf=���dLy��c~;���f5�:��50)H�{*�j:������جSK��w��]׺uva���oQ>���5��E�a��ߩ��[�AH�v�d�����H~h��M7r2:!d�#�8�#�^+Dq��y�I�q��枖�,��][�?�����IQA��P\(R��K̐K����)[\��$~*���#���Z��G��<�3��S1[ZX7ֈ��z3vڇX!)�T���){��J�q�/��L��%�>��vh�uZ߼�klb6��-;3�C�JF:��U#�ʌ��� F�����&��t�b�D̛P���t!WMb6*�KĦ��=2��_�^��ڲ8Nw���X� �K��}/F�k@x�vA��+e�fU�d�{�����!��H��!''�)�2��s��͛�-J/�:�V�`FF�i��`��km��B�c��*�ͨg�vhS�:@��l�S|���m��0��t]��R���������G^a8V��-p;,e�_nv��������o����brR*�.���2��ˉ�Y�ު[Ϗ�*�F��0D���EI�iGu ���iZuD����^�X�VW9'�fW�,q�-������H�4.��G��:����;ɍo�*������<4��?^g��Gbj8<��l����U-�t��e~���h�� г(�s���,w���@ߏ������8%�����s�ʜ��,%�:8M�'Y��־g�n�Fe��`A�#؁��U�[0S�����\���p;W5���`�m4@��=�}dO6��yIM5��&�&�՛�2�V�j7��s�y����ܠu���NŨ^\0�$)�A+�H����n',�c��ǔ*T��
*��%%P\8��$�,\~i��9�9�4��>41�ӏJ��͝���tr��Ԩl^s�������	،�hR��7 ����j���g��w��e)�f��������s�VWū�I�렀3'����*׊K֕[Hؔ�J���q~��IZ2���Qn�	�2G�rmqdi�}�t�k|N����轓�.m�����b:U]/�t�,�{8�<̴�J�#�B��s �=(:�=ږ����6;LB��EV��$K{��N,k��s]�������m�z:мx���&��"�s�ߺ��o���t�'��Z�3�NY�'�~��{ql`;��iY:����ϙW�‑�A��.+�!5��K��L�S��ˀ� c ��]��^TG�� ʼ��>��ߠ0�e�Q� ���
�hi9�=f��b�:��3ϼ�YW�Ԝ|��ց�U����{��,ݡ�4���]�_�*��VY��SB����,3!���fk��j\��o�>�|:9ة �kO��@
������a��,S�*@/(Ӊ�V�4>�<�h��ϝ��qr���9��y� �ұ��!�4>�T�FA�� c6�ۋ����Vg��h��� G� �M,c��+�`=nx���JQC>g\�sr?��W�hTtBxDO�:�'�u����~4]?�%��Sh�6�ڒO����{}E
�D�v^k�����]��}���^�A�i��ą��Ց �UH�7���'I�-UQbK0���o��M~__��m�ޘ2# ��p�]x�1/��<�&�Hlc|��q��W����[Y���Tm#<,�E�Y��{�!B�0;9H��'����6{s Kԫ�W�G�׷i�x����}bRz�'�̙G_pG{��Ш���K�=����sƦ���a̟� l�ӐH���"C���<�8�"���>�+��p�������E���r�J`��
�-�Sc�w�#�Y����h��}�>�%��&~�2�y�q�}���)0g0%�.��֨$X�ݒo����Ȳ0\}�-W���"��W�:��勹��pQ��:<�#�V=g�|~*-˟|e]$U��|�w�����Z��^P���o��(��*Z��AAn]X��'s��Ӣ�|k ��̔�8r/�|����O�ص�i��A	ԶJ�t5w�2(���� ��G�_��&���� V>�Ot�w�|y�`���W��p$���;�96�T�ٷD3�J������'�f�tp|�0�B��
(��m�b7�;�m02v�E�k� �'�:ߝy�	-t�ncc������j�JǠ-Q�/g7NoG*�:�*·g�fO�ie U���
/� �ɗ����3Hj�MF������a��BĞV�j��-��/��%B�����3-j��gLCZidQ@����h���U���S-
rjz����f�UJ
i.A���m������IK���k�xN�?�2�\'!K
������柷u�� d>`+�j`�4�<7C��!T���s�>�.Yh/:�C�6)����Q�1~�b��'hO4A*Gr0��ݞ��s��b�
#WL	St�{�,z�i�%e��m������� >33H
/�rԥ=�� ��hnz�0�˳5a�����*�h�����#n/r��{�.���߯�0�d�y�c��Y	P��Y�,�Hf���y2sǔ���{�싱\�9Vhv�\X���8��v�*6�-��VI�$O`yB��Q5���Pʡ�)�f��fr�����u{�:��[���u�V��6�a_E��<؝R��A4����:~�5GL�ɽ���I��l�S���V��&Po�=�&+!���	H��6�U�2JQv{:Ɛ��%�mp�����C���>�G�V��(3��N�V���c
?���7���|�C)O浟\劬73Z��w|�TH��Z[�[%>8�I����h$1�Y$̐FC�/��<~EK��)�-��-B�e��w9�v�E���L$wb�~�Ч��-1-�H�&:��)�Ƴ���[*���b����'Wz��ѸXA�1�B�#ZA|���N2?`&�b%�M�~{���g�OO��P��p�2��o���U���P�v�
�z�uz�h&K�:Q6�>#
�Z�P�|��&�X�{Ε�y�����V��Y�=���4I������f�_	�K�ܛ���-��ȉ_��:ЀJO�	���jL�]�� E�Ff��!�FJ1m��[V+a��9�^���VK	����͘��G�"�0x�͈�h�M�VޑI+�K���qCHQM��Us���'>�6��A�FU!WQ���C��ڭ�+�Ҟ� 6�A��0OI��g�L�!T�0Ԉ�"�#�x��3������Ԑyk�0�n&��$^x�c���R�[*�c�u�'F�K� fG�mb>�L�c-p��JP���J�TV��F�6ǵ�ʋ���@����>[f^͜q4���1W�ⶳ�3U���zјf^d�� ��af���/h�Y�����~��MTt]?��@�z��rl)��Y�L��S���OP_U�]u"� �:`�ޅ93��c>R��R��������nӏ��z�M	*���~i��>��#�vNa��UVQ���fr|�K,�V�5,K��~|�>�s�Y��Sd߷\�O�p��6�АZ��%+�ɼ���1^�<{�×��|(��4�J�Gn��ARbU�*{*���)�8���(�\灘��Tq,���d�f���	�u(�7����a#��d����2�R�fd������ޣ_�^��U��#rOAn�'��wh��狅����I����l�X�l��s������;����MZE¾�h�=|�*��	@�:�uO	d,L�ڿڋ��]��9��{�wۅ#k%p�V?U���o%���c??	��L"�A�
@��ϓ�U/.��o�7�i�tw8��UwC6���hGs�ɼl�+��R�$��q r�����rZۀ$M�wɰ�8��1Zt�����h6{[OA��`!�^��V�{�ϊ3b^����/6}�X28k�
q����a!��夦�;|�tб��#P�k�4��_�E��HW���~�N5^\��`��؛����X���S�Z���G���V.8$�<����G�M�^].�Et�0=�Ȅ�����'��n=�CP��q�,Z�R�!fI�N����:�S��a8΋�"�$@:�l��)��=w�D�� ���̕��D�G�Z����E����=p��(�� X�Qj�D��0D���%�_߳�Jb1}���sؐ��WC7!��3 �I��CК�e~>�Rm]���j��A- �/���8�?�*�V%��m\��v���_�.L\�d�m�E��P�^��=ǧ���$�:����O��[3s��p�gH���xB�6h�Ɏ�^~ � UP 0Q5�7�{���G)�JJ��c`+�};�*�]�1L	+�����k��0ʑ����>3x���T��$�m,��W����e�UE:����6?����*����2�f4��6��7-�ݢN�r�Y����Ę�u�:����,�~uY�w� 㒡CK��úP"Q��|�Ǩ�#�(,XH���s&W�A-szG*��}�tC�:j߶����.���q$���\�0b���C��%@h
��Hy�V>s�z�#���(�U���c�$$#p�n�#��[���o�:�x!��/V�LT.�� �ӆ���@Q�����h�)u�Q73'mH(���o�9�#s�Z*�IU*��D[�bn�2�����kd�<��t�����3�w-;���C-y�t
���
�Y�����)��f���7s���R�����ps��K�� �ܩ+�|�TeA�z2:ѧAP��H���=���0M�s�N��W�_�W�|��J�J.�$~�w�j�C	��[m� �&� ��{dj�����2��y���c4c��>N�����*�|�:�U�U���=$Pu)D�����-����^7#g>�[Kd[z0[SM�.6�z"'�D��*��9s7	�j�z��u�Bs|ˍ��o 2nn�P��5(L��Y�y�(mei7���1��)�s��u=i�-��G��7R���C�U
/f��K�L�:]�"_�]�:O-�j�����.�K��cjܴ4���9�n�ZXb�(�CN\k#���mC�Ϻ�fth�Tt`}{���a��}�����w�n�5�/����T��-C�%P����c�+�0k��@��X���B���|����O1�+2U��m�i�t�s��Üfz���?�>�]� W�?��a���#c8x���ir9�ti���{Uh>��pZ��%�Wm�YW2���0�O"�V�鎁R
X�����KYV�@5)-,�k�S��\tܑȯKZ�6?ۖ;�f(K���B�~e�j�����G#@b5?o��kI�Q��*q��?��W�m�+Z�Ī�{��ć�e��o��rI��Fo��`��_XGp��E��	��f��"�kHQ��y����2�Od����
z��'�#?�^
iq(����3�����}�2j�g扳f�*}��$&s���-�D]~q�M�@��Ė+��缙H�R���{;�{�N��E��j�>'�Y�7��"��|���I��\)(s����v(F�bsfV���tTM=f.���)��x H�{y������T#rQ��}�FG�JA����>x��4����q��uz�4�y�L�p7I��a�X�P%X��^��<�ٽ��t;�e���>��|�6�F���KT�&N�k6Qs)'(�5���"}��2ގ�{X(.u�����^AE�Wo��a,+���'�6�j����"�U�4#F7����M��`����\�	6}8�]\���I�l�B&�$�Hح��Mv����Ӈ8x,�/���4�L���(9��?}�/^��ژ9�]D�<l+k\�G�m���
%w�'�H#���P=��|o\R��
2v0���=]f鞡��zp"���X�m����)�(�f�e%���R)zb�����z�4�$Ti��9+�����x'+��mP����
�܂!�C�^��:v����o�Z�4N�B<��<�a��=�2~|�Tb��tץ���\����|O#`R�9玞�	6�Q�N2?-ao	��E*=N/�)�*!qTז#	�����νD��(m��4^U�oD'�g;�ʲ�$�;3.�P<Cqļ���qIY�G���P "�x�8_ǫ2�&9�����:�\���$���'z����^(6V/�����Tf-��Y�هK5,���0�i5@�&HS�g��	}N�������?��x��(���C�K �Ϯ���}�ØRq��i|!�0�ǚ�-��z>ӐPZ+�W�&�Qt�N@��fX�?��IQr�=2vH#n�< ���f]G�����c��V�
6)V�|&�y��ڪ�$�,�fdiv��+�nc�|� _L�nP��7h9��2��/Z]a�r�n�` ���+H��V%i>�5:�y�[z�n#�ͭ�^�[0c���;?�/�:.�Awmf_G��)�d;< m�%{�r	[(Z2OZ���a���tEr6	���sN�6e�����#�5�XIF|}��me0�:�!�������%z���T���n+�,�5{\:���@rT�hl�� �Κ0��rSOu�w�ʌ5ț��ȉ.a������vKo0v��>�-$yM�/��S��)��Lj�ڥ�g঱�{ut��$�$һ>9�����
|o�#�A�}/��*~���N�`(̢[M۳�:F�vX�4�l˹_�^��p�\7�7��0�b�II\�"�0A�PA:���a�g�!���\�Ӻ���\���xPI�jN�K��8�����%�g[������>�l��Qfل[)��^3��4���H���(�'׽Ƴ�2Ag��c�R�
 �����,=MRC��$����Y^����`�]xg�Ճ�6�g>��홫���[(�taeuA0T��)�ۦW%�w�Ժn��K1�@yD�$��*�Xk�scO�u;�L�r�2�ٲg�DJw�K�';�bى�Y�mH�Ɨ[_X�����b���
��G�����]�(���?u������^cj(�����t��Ѿ*�lG^��ꈦ�WV�{"j�s&#�^cM0�d��x��
�ȟW��{��c�#z]��tk��R��{U�*֛W�V�.B_��o�'�Ok�BJ:�k�a������]8HO��O@Dt�h8"��f3ҝ\��B�p��$U߳�I��[��|��H���8��[v��"h[�H�F��s�]��7�����?�7�aKU��P{.����Z��c`��c�/0�D��)2�����֌*��0w��xo~"��i�AS#��>���$���x�o�~�i�RK���2�KE��YZ}}��T�c�ʘ���G��{�'"��ʰ��b@viٕ��Yx�Gwpz@ÓCp϶	�����8G�JI,h�?�'@��u9��Ѕ@6���m(n��}���,��?ܪ ��#L;,*�f���BO�:�
o�:7��JD�7%[�]��ȇ���zj�g)���3���*��0O����v��#P{��iIN"��U��z0���oQ���l"�?c�4r1���w�!P���I���$MdA��G��ouL�a6<�Ū����j��0D^�h�{U ��F�cn�Mҍkv�hd[No�E;fs/�*u���������w[���<����+JۇR��-�k���џ�3@亜�a��b�&�に�j��!�_�]��ө�B�q�P�26rҺ��6��og��=�R~l��":�d�I�05��6N�P!!��dnL����L]3�c<$4 �V��^w��bI�;V���^|�y��\��o���$��&�_b��8*#0D�Z���D`H�~h�s�s���/��3�@�t���@iE[L3�H���;N���nd�1��)�[�#=� ��ۏ�1�˓�Y�;3h��c��ل�����Q^�X`@�K�U�ֈ&	�G�
�Uc%�9�1jA)�G����W�{b�ꭽ�S��w�p��'�<0����DL��_���|=�ݙGYy( �#CdX�-��x�E0����x��b�y�ۇ��$0v8����O���S��3��"X'Q���Ii����"�"����y[�b5��\s��d�?G�E�b�c�}	�mOi?��{���ys��Ɩ	u[��5�rW�1dFtnR���5 D�4	����+n������T���}�W`�+��K��`�l��^��_�r�U�Z��<�v���?6��R��c�f���a�&�s�QDS
��ǀ�]���W}�HP5-�6� wł'�NZ�&�E=B��]7�I���|�S�JR3�fo�&��js�������.�V0dp���|I����s�q��E�l����1�7�6���A�O��7GxK٥�"����7�)��浩���8���KR�Q4�����'ӗ���☩��%I�Ӥa�񘌳�d4R�� &?��%}�2��/"�d�~G����;W�"s����g��*�F��˅����V�{�d亚F�z��P�>h��E��4��*�wg�Q��v�s�!^�HU��x�.	���+6A�Z3x�b�D���3��4;���6m��[6�U�`�i�gd�!�nL�sE�����&��g�3W�&u��Xi �#���r�Aϣ�WT�h��3�6F7�ܓ�`+'����)� �nB�����ʂ�D4,]��#Qe���b��8��`�:�
��V��<^ϡ�V��<J'��Lϔ�J�"G���Xw�IX��H��m󀁹o�Yl�̡ϝ+#�vD�:W�Xl�&;
�I��_��H
�Ho$��*���̷���m�7��~��!I���&E.ϮLR���h]��}$�R�w����| �F���5���������Ťu��NVզ*�f��V�Y��"H�,t@�f����/��S�֡WoԌ�Q��q�%e�nj�:Ƴ���az�������ͣ���d�H������^��A��&A�U��]���֣�װ�q�����������>�����D6sy.��a���-��KQ�����B��m�YAwӤ=���M|����-b��'����R�6M,�6��Ҥ���zeDo���-�<�B= ��3�L����Z.$��9=�O��G�zR)������S�s#�G��<��g4$���BQ��̔��d�����䗌<z�@���.��|d����`�.����՜ͅ�������EbD'��ˑ½�@y����,�dc =�l�9���ZL���4��z�f��E]�վ:O;�o�+7��h��z�W�G	9�Z�s��`v����%��* a7]&z[G�q��"#_¢k�MU����
�|�Z%L�"@ �~���� �`�������(�`�n���A�٘��u*������#Ҳ�#+���	K[�_���
�p��}�И��$
�,�fk�}�o�#p1���`
�ˊ�H�Z˺�ɱ׬jQ��Y�H&h������oy�h-���٦�W��yK˯���'�dьޛB�L��;i�s����E��&|�_��#_���1̻���v���2��<�[��[k氙I�h!�Wz��%����2\Lç3`�2��g_鹒�Lƭ�(0x��sa��6�b��͒�wǤn�n�P��jT��<V��^�s1�#�� )���h)��V�w�7wɋ9#�5����?1���C���e�5�^�c�X�k+�>���@k��������/��MU̽�������Wn�a�d���Fwu_��(�����V��>P�ϧ�����S���p�ɜ=K�ٍm\!�� ��a�J�RO��g��6֧$���g�p�b] d��ub��>��`13
A��rG�_1C"�!��#������:�β�2h"y��uT���	DL9�~�\�P�$I�e�&��x�(����
����
S�*�x�	��2i����_�oLY�#���3�N�|�/��^M��_�*a=��$&��7S�;����ņ�U� e�3si�tx�5{Z����M�qN�����Q3�Y���K��u��f�Aj@���q��m}����5�= �����XeY��┭���� �����1%_t+�Piq���n��imy95�9b�g?�(+�
�l�f����U�,�������'���ƃa!H�x��}��˿��h�[�{����e��.� �VTU����q��9�E,$#h/DO�-�:�.$w�;�{Ɣ���j�û,PW�;�}�@����Ӱ�~	CSSߩh����N���	G��v�:Ie^١�ț��-��hB�.�N:>�����AO$ctxiW�+�ɟ�B��Z���P`�AU���
Äe�R�7C%M ��YY�j.o2��Ƈ�����9�ܬL{��Q��S�BLYR
9>�Z\��2�Jt�e�'D?X�.� �t�px�.�5�_��9��u�[���ʇ�9�:�z�H��3o�o���P���QT�0�a�ċBR��?	��?��08ߎG�T��4ej��їV����P�����~2gW����ۀp�"5�w��&��I�;e��=����'��P��1F���������nW)�=�b��V��DG�4e4R�Y��_�h��d��q>��{wH��V1H���9�gjI-L?��N�
3d.�X��0�F�ԝ=�.�B�3jo��v@�g	ЈNӇc�.O|1��Jh����h�XI�D�W/QˑĬ_)��%�)��<Ȣ �>u� ��ҿ�]z�K����7�(�^�%�UL��,��χ�Ǚr��{';4�8����[;6�T��������o
7Ji�W�{��.�9�☚�c�GFT��q��O��*(¤t���Wi�`p�S͏j���l�z��:�罅I�B�p(XKҩ�z�������RKp��w�5�&���	�oq��}�H��#{V�<�9�rR�O<�� �؀/y�󇃛�D�5$�
�qͱ����uR}<yFd	�j���"�2ߗ��םd'a�����o��?�xL�,o���3mK4��/����m����y� ta���e���Bҗ��kH�r��K~8LzkG$�Yә���||���Ӫ��T��`�4���r��i��z%��3�!��P7�C�yDR�x:��C��u�8g��(B#g��8|=��!�6d���OpE���;�c�������q�S��46��J��S,�ˢ�-�|Q��?@*�|#����]��@�B``*0;��,�޿�L[wx$4��:;6LYޞ�ڲԩ{�Il���	fޤ�qC�b�6�/���5�3!�ϔ*�%.,<�yHcv��F8-��&A��V�PC�����%��2�9S3=��$y�i��_}ss���/�:�6\�(�Y2MbH��:�yGn����y�����c�)ѰB0�-
~��Rq;��B��k��b.3[��#v��Z�1D�4t�q��;U�f�&���� ��AC��/���τg����^�1C�8>�}���g��a�q�e�3�u��,E��a�C?�I3Z̛^��cAsRy+ޗ��L���X|e��{�fzp���*vsv�[B�Sڢ_]`޸��V�+�T�Y(ɍ7�D�9�^�,&.����؎"]�@��"�O�k'�"퐵�_�9�_i���Oc�TQ2��|b��g#%uC��j,�9x��+vZ��ERM>�5G�˯Ƹ��)�h[���|���<����#��G�w]�&/w��oR�6v�?�%Ӆ�ݸ��'(]��H����-XA}��$4_7h��v@�;��}�T!#��h�l"�/ϐM7����,v-='@���5Λ@�i�8F['�H��y������K�Z?�T*���E^k\|�u�E�E���R�K���nm�H��Bb�:��T-�(۽
����K�}hD4i�C���E�Vl��eUM�-)\�z*�{�r�	�eX,X��F �k�~�:0v��G���
_wH !�σ���R��3�ɿ0m�~phv>;W>ɸ�;�	��4�ACJ�=������/�?:� ��Eh�}{�QC�kv0��0x���t��-��h��E'k��[����+ӱ"t�c$.R��C���f7��u
X�ʦ�m�p�X�n�
���!�^�͚T��{H��򁿎";����1��q�;����_�_>Aȉ�|��y5����.�zkb�q�������7�A�j�>TB�ױac�qY��pf�#��<��-c��<-E�% �[���n�|0�vJ�^�y^�M�&��@yM8��b>1l��@K��u�z���e/�'�K$s��Y{P��t�2���ޛusF��I�E��~f���%�������=��(�G������'��g�ë��t�Pk ��q�F�31������#!G�^QQ�xHQ���!�rN����j�V��+����_!7��V>�C�I�e#�D1+g@(�6�f���@�����aA4h�O��ZG���,�N��;f�g�g��ˎmT����3�Y�wH�hd�dy��5F:OZ�6'��c䉛�O
LGX�*��wR&̎fqe�۞�̼�7�-g*�fsP"6� ����o�&���٭T��L/�Bjl�an8"�}H�݂_t�k����@R/{�?���� �1-���M��� 5�`"�G3�s��]�����ˍ����vS��&y�W/���a�z{�G����Kj��x?�$=�������������V�乜���4^]}C���W��ͽ��*��аv����1��x��!6�;�K���5 �-P5~s6����E��͍!(}Ȅ-:�;3_�8Ue��a�&�g���W'�k�c�K���ߌ��U�r�-��Ͼ�^��bQ �>6ź���(bE&Q
C��/)��ELw�.q�ށeI;֚-W������(�IQ_��M~�:
n=�c�Xऀ���i��MSh���S����^Y_�|�>l�8(���!�}�)��MNE��A�xZ��:d,0��6䧈N�1�����_�п�)�w���AA��|!�B^�� ±s� ����UtF���ӳH����ĝ��AD��ST�pˁ���ig0)Χ�A;����|��<�i1�+�W�\`rpkm�^� |#���|�|P�X�jӞ�%g-�X��cŤ\�V ���ߠ��ݫ��n�7����4yErZٶ��{�����?j�:6�Z-�qvJ0�N�\�F�)�<9e7Iɓ�����Gx+X�n�D|A�j+IHE�ש��!����RP�Y_���'�NY��m4l��?����5����f�z���)�E�&KB�kR$נ��+ �A*��`-a/���ꃤ�U�������8zxd��:v��}�����>��TP����Q��%t�J�����Q�/�I�2��!�c�	6�?�z1LD�:iW��}���,7dE&�f� ���2��*�if?���L#�#�'__Hw~�)���i#���x
�e�p�L���j�cRr&�
�0�V	��h�%�?\��=;Qo���g����Е+�4�����3J�T$���)l����@����KF��zi�&�W�. ��N-�ȣToiA�B�N�-?R�v�E�#�U�1v9iD.�[wOº�^���Z���a�:�8k���}��])	m�ŏG�S�@�|�ޡ�>�'u�k�I"���ͅχ���0�-���~�C��=W~Z���5�������V�*���q�ݬ��d�����2�̔g:jEg���e�|3#˅����h���ٚ����P��� o���o�?���>�zF� �n�X�P)������o��^��q�s�%>-����t�����$PШ|7<(~{0c��'�r���a
�`Ѭ߇�k��.'W܍��]+�õ�v+��[�����Z�|��֘1�x9���q�1���{=����q�^��0��k}w�f/>��jM(�<�eX3¸Yw��;B��\��?��I �F�0`��@R�G�+J�:RMl�c�?����p�=Θ;���M��b�9.��G��7�`P�u8�ճ��:C�X�LG1(����
��ϕPi�0$��F Y"��O͗1qQy���KmK��·�-9�N������	9����{8�x���C�W'm�T��n�du�_>3�'uJ���0%N��_mQn��I>�ƶ�D�īJGn�M��\J���7RY�5C�i�c��5�Z�;rc��~��$����U$?\�4?yhiB�����x��<������Ȃ�%��	5��>��6����9^��c~��(��Hځ���t]�X�Ą$�بy��+��3IQ�Wi���fM�<Ȋi�Ω���yc�� ����k{��H	Qo��ǝ��(>�I�_�x@n@��G�bc.�K?>9 #Yf�?Owu����k��}�Yl�*�����6$V��ѳ�#��1#��xKU~*b�f��ѭz"8�齉;X0�Iy˫f�Iԙ�wM�L1��'�8��8�PC����5fP%�-�t�����(I��0��.G��j����e`FJ���=�ĠB[���~�Ȁʰ�1�������4�	�CC�ލ���׬�p����xt?��"���y~Q��/ߴ��R�J	#�O�g]��4����g����[>H3>���#�g�3���yt�_�=�$K�ѳ��<�lp��Z�z�@�_iu%ǐ�
��ָV���o���l}?5��R�3~t�$��j��j���s?!���y&]|!x�Ue�L�W�~tƝD�p���1��^�^�(��YMi�\|Mi�R,��ǣZ���{��*��{@G�%�]�d4�8���v#QYF�Ͳ�����f��	���׾dC�ұ32�îc���6��\P��p�P�ߚ|��q3)�f�tZ<c�ENzss�YH�Ⱥaծ�]�ZI�KN �?��*�` ̤dPF�ӃA��#���?�!k��� ���ۺ��ցб��1Τc�Q���0��Y�q��#�ǵ��Cɔ/w]pw�wR�Xg.��a�����T��)��P��緪w��Ow&c�4��I�e)B�9~S�bf��j]���H!�s�ζO�"�J=�T@%�B������w��8̱�:�6H�[$�h���F�N`�w����F�:�;V�s�/�t��@���}�2���N]��mX����[ܖN����	���������q�d)����|D&	��?z{�����I�����ş�~��0����v쫢
���+܏:{���_�������#�$�9���U�	9���Hcx�
"K;�w�n��_��Ca�L,W�Jb��v�^0{V�`0��99�������-�Ӡ�Ǻ>��S�/���}w�s�&֫�K�d4<oY*�T3J`��O�ͦF\GU��pR?��׊� �@�|�c�5�_�G�6�BG�tWYu��� �LЪg�|�������\n>QԖ������^���y�����`�-�<��	*�F�%)EE�����p5v����Iu?��_I�S�6�� �>MX�hIP����=�6+Ê	���
;��Y^c��;������QQ�ʠ�#�-����?�2$ʪ�
r�$�ٚI�2�����V�`��Q����2Y/��.�oKMI&�u�\RUAQ~��}t-R�ȔЄkR��[n�+��!^�F�@Y'M<��Ն���m���bG�my�iy��4�[OUn,��a֮3���A
,�sLI�qih�3�o^��2L��$FH�W���� ���{�
�i<�mRz"!�[�d.�0��N�%�X[n�R���'���V�� �x��5c�:G��|O�D/��m�����8\:��^�Y|�U��F���$\!���e�@ּ\b>b��W�]�b��Ȕ	��?4o^���L&iJH3ȑ\�<����QN\>��CA��ǎ
����:�}��c��Ū�%<P�m��F��{���6M~��ߏYǌ ��A:(��wt��Ag��6���H[����Br���JM�J˪���������F���Of�HXhW7�"�$��+Ã�0I�9��Č}�wX��F�e��;Tv�S�ȗ!z��˹�������
�eUϤ/#L_P�xr�\'\U�^�Dj�ч��5箾�j�"�?(C�H�P�쨙ǂ4p�!��K�d+�O�����׋`���}���v�� 譀�X��}�On~{0��3'�V* ��Is�������4E����g���lY"S:{�|O���#bmk�-bdG\	����`� A-#��l�m�l��p����_����~��2x���������
���bv2ڻ�c���U��ڞ��xZ؏��7A[�F;�6$�H������.i]�b�B ;G�zLG!����&폻�	����+PgŽsr�nm�m���E>^�z(auQ����=�q��ZG+|T3�B��k��;4Z�<>���f��st|7Ѯ��TP������_�����bov�*Y�R-����]��;��墫��������>m�	�0z�Nb8�m!��<�@�ķ�v)��Y����J#��H��n�v��zڻ������QW��Y�����r�ɽC�{��h@��� ��E������>�1dyjO|n�H�\���y��ښ�/Q���k�U� ��0щ�ީ��]8X�z�վ������5����[G�u(�,���Gܺt.��Y
5(���sı�+��F��L�F�vj(�J�C�B
������^'�@�X�%���M�*!�S��!�����4����+��X�ɷ!�1�C��h8E��Z\1wY�i��ca>�W%ŴW{ku^�X���v�Du�vP�e��$>Js��XPQq48n^~VAd+"-s�Ϛ�IV.wC���%�����	}�m�R�SN��9��J�3Ka��I�H�|U}��N�r���Z�Z�w�t�2�et�����2��o8A�ax��b�g�X]�da���,4���� �=������©#`��p��Ӂ�x�?�D�k�o��9���҉�Q�V�[�y�{��_�
��lFi��̐׺�|���'���z���޲rLgh���p�Dd�.Vrm+Eux�5�Ag$�'n4�j�m�u���� �k:b	&�f���4 �N����`��AD
燔���w��W�{(��H�|�v#?��(@�+��J�k7�R+'�H�I�4^ ��;�g3��5h����M%�9��]P�5�zY/v�P��_�~���oz*B�-��������~kJ�|�N��M��k%� Ǹ�Vܺ�1([��A:�.��%JP"_;^o[��:�}M���(����'1r�h�V=�&�[��9��R�}'M��OR[|�ڭ44��5�w�ÛY@��Gj�	OG+��ÿɟ�y�Fy�N�k^/��]���m��dJ�H9����J�AF��<���k�3�����)��l���jM7��C�3�8�`�	֤�^%ݐ� a��+CT>��x	�).t!��ʗu0p���-�04d��-{+s��$r[T�L���)���"m�s�WFpU.��	��3G���O�"���a��&ց\�yx��D.ƺ؄�}�Y=��P���|����!M��؆�y�n��WMk$��S�}AI����Ǵ����N�? ێ!^ɸf��Q�1-= F#�^�a3���L�,�o�ا���.�'�N�-9yU�!�z`*�0�w�e�O�L���#��ʞ�|aD�y����%!|j�Cv?��E�6A�-��ɍ��tk'��|��Q� k�c��ֿ�1y���;6�'�9�RЉ�,f4~��b	�O�9��-kS���I'z�N*~m=)Z�-X(�uѦ��جM�1��g� ���# y��>A֎	ۀF� c��n�)���-��we�u�U��%�>���L�8��+\���
�0��<y2�~z�`s{��I~�$�U���	��@�pGM�3r����C >���b�'��^�Qqv���S�ș��I>���	��Tp1`�ę�'W��Q����)��r�FM~T�kP�]�u��v||���
{େ*0��%#�v�A"i�����c�#k����ʍ4-�D�
����\=w0��S�lo^��2+(�k��-wr�c���ě�w;�{�w?���q^�%8�{�=�_��ٵ�гjXg�iO���QЦ.f�=y�3�L�I����.|�˙�����$n���_�Y�͖}+;�m�#��]?�k>���]�V�
U��S_�3���C���V�Xk7�
���U~�[����h�g��e��m�
SOh%�U���0�[��Q٘���{`|����i˫�'[�l�|�ab�Q#��x��M�8�?�V.���{��u�sfZ���ŕ�t�)I�:��5i�Ҡu2Y.+љ�E����'*�������8���m��}��%ޗ023��Ӆݬ��>v���+�R ��OG��|�94�C�F*o �Ov���:Ӗ���w��質�"�RC��'����k�;ϯ�ZNHc� `B���V~�{N�qt�%��w���q�2��#��3��K�� ��T�Ƨ�:�x�Oo��+�:ˇw��J45V��ZP������C���1}J0pؓ��8.-�ҕ��v���"jA[��t����{�H�q��i�N�||gL~`p�*f,��F�i���{}�'*xF�Ezȍ�iP�P���F_��e`���;�p(*������AT�9�j��-xs���S-K`_*$��WG��u��h�����;�	v2bӯ�k�؆ �$��%�XII���E��5&��h܁��e��P��N3�A��Z�M4�\��'���.߿�R�nA�R�Fal���͏/>Z.s�i#�z�g~�$㭺|��>����D?��R���#��}���Z���.�?'��yb`�%�9ԆO�`I~�ae�rH���_�1�E�]�g���O�!��Y
i��n񀻴�9�UΊ��05V� �_p���1=��dw�����>���"�9Ò� 
y����=̥ {\��-�}��m{Xq�rj \�=��p����t�.�Oޑ��k9���:����}:Q��t�u7�MvG���@�ؐ#
w� 9/d���ʅ��{S��8�!���s���M�(��n?���K�������O8�91T���I��Z���!�H0�O�i�}Y��k��U����m����%TVV��0t��:����^�F~�G�N����Ȁ��N(�܈[�%�B�v�=�D���X�FU/TF�t����N���Xbl �����q�����H%�קv~q����Ӏ��{`��rؽI�2�DqO�h���9?8v՛��g�Y�C�+=zV�&�&8u7�OB_���Gį�6������]�v��ｪK��̪*�^#3C�.ZC��"���4���#�o���R5-�0G�q�\��@ ["�ݶ�#{(Y�p�E�
��MI�O��X�/���S|ݷ �K�&"�o�LTp2����rCF�Kq� <g� ����4۟B��Y�����D�[��'F`֭%���d!	a9"ح�t�6��8�瀹�wѡ�v�˜1�&������	��(�$=����&^�5{�&Z���*x+���`�37�7��v%�e&��+?��T���R�|�=w=X��vo�Q�]���LI�wU�1Sʌ
<����9�-<;1���R1���"(y׆Z]�~�	Y&�5�?����m�Bо����&6��S��8tv�:u����lmq�@�7Ѵ+��(3`H)n*)��M�l��M�N!��3�y�Ǉ�v��-��"��kSz��8�JӮ�i��Į^����)Y����°��g�n�Y �g�:��^��C�(Q��A��a��g/j(��~�`����1x�F��W��U�uI�2���cr��iPNE[���zt�y�Q������YlH�ַ"�r�J�u+J�3�@BWtH|��h��izf���)jA�V��E��#;���}+�XT02]�κr���@ڷ�?h��%xwe{�'�E���"^,�<�ܓ�l��o���3D�lxذ\�*�D`i���_� !�;H���́?󀮗&|bȵ��������lV$��E�}�s�XލA��F/U�'�DT������E۝������B]��͋�6�h��A��[�R�+��kQ�S��dU�&��^��S��Wv.��Լ\�O��
���Q�LT=V�c���Mqflb�������Y0\��YX<W�i����]}�Ԫ;�8�`��1���ϫ�R1O��ھ)ȢJ��m!xrQ������I��a965�������R#��2C%�?c���>�����iW�L�����d�"�kA5�2��v���<��ª<��`:�3��I��B�;C.p��s���s
����L���R��j(L�R[�L�3=�/���[��n
�TEm�}��}thf
ZK>>1��8�z(�ȅc�6e@бMM,����F���h����@�ܐy�:���y��c��������A����CR��Z-�[�H��%��E���h��0;r�i-��$��v4��5
�������ۂX�����ߞ�,��괵4�hx�}����9�R�]Mb��Kp%}��b��b#����#`�XUWn�0@⢡�r��G!?����F/�3�^���4W@uq�E��΄���j�#�I8f��P�a��Tksh�g�D�M��g���NV�p�$�e�:1�2	���NL����L�A��h��wF�;%�ԆQ�0ZM5�1�B��2���׳ZO�Z�$�+@=�&B��M6��IH��@}{�����l���S���ý��+@Lnҏb\��&����DnG���-�t�N��b�#���L�4��wg�:@�]�E��Wj��KK5oz�f�&��N<?0�t$��!3̦{�qA+8`��
ɑ�?�\`�-sc�b���$�ǅP���ɉ/�'em5͚>Ĵ�<)\0Et�j��~��u�[��K�h��`?�eTn�&��K�<�Mw ��9�W�x<z.��N�Q�]��WP91�Lɜ7�7��T���_�$��u~����ߜ[؏��� �W��4ȴͬ�|?m*n�; �w��O�h���T�&O����WW����y�עL��J�ڻ��n�2��]�I��6�]���7���f�y�����2��!Lawv)|07�cL�4�x�*r�.2,�C��V׺�b�6�A����xֈj��=�̲D6�Z-r�ҳN�	h�nJe
�p��-�*M���L�U�R�y�����ܬK@���A�"�X>9xv�oc�g���2��h|������j�d��pE�;�b���ã<�k�T���u��=��<n�:G)=|�V��p#�U�yI�����p�4�Zb�W�%1 1�1�J��v�dD����g�]�V���29I�H�}^jn���T��~�Y/�YMel�r��Ϥh�p�R������:7�H�+���z�� Z��
��K?<�2 �j���Q��\�k����^*�Y�ڒ�L��՞�b9%,� ��#��?Ͼs[���S�ly��>���ע�����q�̝aɶ͐;�Z�ZH�|O�x`Z�Q7z�Ѹ�ON��CU���ܿP�s�L+ӌ��iv!�t���_9Q�͘�5��#?��3�Z�<����+"{<�;׭j̷Q"&��j:f;��M�����!�U0l��N�n�`i��'e�/bPf�� *b�x㩦�I��b��#���LJ�`?U �ۄ(w�+g�i�룚���#�@BM�:| l��1�f�/�8v^����NBE�^�;��u�.����-�J,�=<���|!���V�}�H���O��H�C����m[U�&�&��C:����@�)u�cL�e�^8K>1���_��>��왎�-�E ��=�;+S=�v�؉u�V���Wr���;���3A�Bʠ[0�xuJ~���$�=[2�l_Pz�y��d7B������A�XCYu�¾�� ��p!���������t�i��4��#��M���?�I���ڻ����4<d���?7@yB�;վ��sb����ޯ��x=��^�~�_�����2Fā������O�O|8�y���_ڠd�t��^A�O@s`�9�s�� Z�EQ��c<��*�sxQ���nbw��U�j(���4�I/�LѧMuN��vS5�?"�������� oD9}�T��j�O�H�����=S&n�S%��H��Kp��Z��*�����g���_�keȴ���NU�g;���i�R�7<��Zuy"S��rJ��,,�Z�B��w�IWP�]&���떖ѥ��Y԰�-KV��$���>��}�`�2X	����o�FW���O����D�"���a�zl^B���9��A�Lc��{�|�l StG����b��o״������7�o>��7����Ub��7��x^8Ƀ9i%��������H�s�l��$!~ح�-B����F�
��64c���?�u��8ig���0����a֧����p�Ozڃ���-o_�HƬ*}f��#�3Vy[F�UZ���Y(t[��"e��ym?�~�Wc؞t������c.LmB�&�"�ͰF�H�gYU�&V�D�y�9�+H"0�|,�Vi���Vd<xa1�N�l6��[j-��Q�G-��{���J�`�96�3ֻ ��"Q�1����e �s���<���d���bm�����;/̗\��|l��BZ�!fZ�,�6ҕ�DX��VUx 
�2e����K�p�i���D6�C1���U�Tv��Z�zR���ܲ*�%�d�)v�3��IOg=���)��P�(&C�>9g�-S������r$��!��N���2@�jr��=�%cAX�o��0���5x����b�1�v� �5�.ߞm�ˑ@ܳ�I�2�����[���$;���YG+�l�M鵺ǎ8h����  \"� 4<������6OQ��ٳ�� �?�`����v:
��/r�������8�J���xC�K(M�f���,�3��Yu9�N�5=*~c:s��j������B�������6����{ {�Nf2V���c�R�W���h�;����b�����&�A���$6�u�������9R�*n�w��������_��s_}�(v�o����b㑖T�3��P�/��[�O�F" aKT����(y��,a[��jT.���մ^����V�~�?�ԃh���NMm��tW��fa��"`&E��<�JS���~B7W�F�37���k�_���c������qA��ە���Kn��J�+�/�jf$��=7x0e|}�A̪m����*_���GďW5�^x(%&!~~(�+|�?ch�8�>�g�3��}�/� �s�!)z���t�	"n��O_�C[��s�&�|��s�S��z_U�x�y3��4���A��
_�<�����ߴX[��q��,��������o������ijq����)��L�li�Wn�{l
�Q� ����y>�C�[`k�9��p��:_��?k8��ʂ�h��EҚ6�����(��9N��]�e����c���M�>ţp0������m�,���qS.�Y���*�Qe��$VAD�`�A�v���w����[*D��[(�@��� �R�������Y��z�vi~��93�,�Ƶ�@0�O�������U�O��7�v1�S���2- lW�JY���<�t�;���+�6����=�E���'��
�3�atG�oB	*M��k3�0�@+�E(�ŀ��,ke/��J\r'��0M�]=yEC���jþЪO��
pb�?Q!�y�����S ��Y� x�J.�����!��o%���l��y��]00s3|ؙJq���O������%/�p��aC^�9!P.���M�����:w=�jG�-T7�x����'}o�pͷ��I��ԗ��\���� �H�pV ���k��z+����&3::ndu�8��X4��ԧ��k(3�
KI��;3��>�y���`�ȴ�r�w72��믒�9���(��k��!9���;S�a���/���va�%�Y[��*���C� �5����v�ؓͨL>�~���c�9Ip�jg���/�@�aHޗr����If2P1��i]
��ũ�FiV�#R���&�T���	Һ��|�G�B\��2�2��r�N����,�������m�����0��cS':#�?SC�r�O*��a�wi�~ń����ic���p�t��)=���4��VP�>S����y���/���c�&�R󶷀Z:��i�7t;�0Y�������`i\�acV볈B�^�{���gRt��轿k�����|lmʳ��f9�0A�^�ӗr�_�$5G)dW9*ȋ�|1�Ů�n����hu�*�m �X�f����e3��E���O9ņ�z��՟�#W�Ʉ<!c�Guy�Q)��	��70��[�L�Q�Z�0�`;z���I\|��@3A鵞����(��m�7���9?$��%Be]K ��4����͎�j���#ٴ�3��5��-�VdY'�P��r��lMhN�3�wqW���;���1���8�v�����
���Z�	�?EW��%�t^�C*����!���G�&�5�Rt���0r\�]X�0A>;�/��VTK�@y$��������q��P@��܏B�����p�]]"��HKݾ+�M����A��a��)�K8����S�6�
.oy_�x��DD��C�ʣԷ����g��pyN�ȶ�a��7�S	�|{	����,��-G��譧J>�Fy�ⷆ��FjA@s"ߍp	%V�5��0Q�1�Y3|���s���u�A%���ż�����&��Р�I�=J|�.ޖH΁�0^��{�+1*64�<��q[��Ը�=��3�F���eٚ<k�h�LF�e�nT��'��.�et9D>��4H��V�z�囂c����<�l>�_TM��/,��Wy.�+�{� L�d�Κ�F�4��V���L�]��@hl�1�o|}�O{+b����|P����⑗�;���Z�U�t������~p���&�f��,�M0�܂��E�����v����t؇���|*��ź��:G�U%��gG!�ӟ��{�'�\�}�A�ݩ��+��@�w,��{�(�3T~���p�+����n�?&`��-ֆH��DY'���#�#��o�c�B(i-�(LUC��XY�	*!"gx��:ӄB>8���Ȩ�y�et�	+h�����]N}Npî�Ҁ �wRߴ�2$	���|!:�
���.>�(xi��[W	�"��Ð�2%����n}S ��2/c��4��jz�Ò��/[�3��C���JYTKW��A�?�� �UT�O���g���Դ����<�>u&�h���/�,�3�9�O9cM�{�lo����6pz"�g�����o�ퟢ8��b3q~
!��9����BC�a_���'�c(ֽ]L��I�N��r�16)�&}Gg��(�z*q�t�����[v��
�G3c�	�X���6��8�#�.=K6�=@�����2������}�Z�ns��(�8r��BL4��-K�����t��= ߔ%�{���6�B^�s����T���EW�\�����*���b&���V'�7��w�ꂶ7hI�����H�Bh�<�8��)|�B3��lsJ+bfV�;���t��1g���J8$wIr�H W�ؗ�v7��9��p�&��jCl���r��*L;L`�R���z��2�˦�e��ЛWh�� a3(�-�I/Bʠđ^�S�� \���Z�^1�dS.�/����X�+) ���:rW(C^�@�N)����
��=z��O�4y�1�o跸-3|-k^K8ʳf��m��zvyEi��.���֦p�(�O*�f�s5J���b�17l�jY�dX����2ch[E\,���� r�/Ȕy�/����]�gvh���( v}���޶�1'�@eMب�V�m���s�uuc �?�#H�?P��ab��<țW���R�?<����) ��N��Y��Η�3���i^(ۺa�ηuQ��aJ��Ek,-n���:��~�3�Π��ڢV�U]Ԡ���-^~a*��UkṞ֠E5��Ѫ�8ϧ���r���xB+�{g����H���?_.���x��=���Y��\ݾ�yD�i���IO��}2	Md����[~PW�T9M��ϓ��e��O�2���p�⮦Q[��{"��}�7	Bb/A �3.N�s��)	�C +��ٶ؆��0�'ʳ~�N�!�A�y��	y��-�,���	u5�p˒�����Q��;pw��c�%�IL�)j�@��������P���Q�8��u��C�a8=Ck�&벂a6m�4�iO����A�Y�G�2�RX���ό�uI�����xj�����Wù['A�@ά��'�Ox|�&3�`�`�'(����j؛;�_u�i�н8�?���c֥���d�����1B/,�(����1���k���I���s4�(�&vq��_/�7D!,x��
|cP�@pg"I�L֨ad����X-IdL���~���?�R�=�(b�PK[v�e�-�h�݁�<�GS$ �?�Ӵ8P�۠R;�0w�������yo�%���D�,��F$��.]𺹇��:k'��ta��*x�b���mCr�b�>Ag��t�ԽmrMJ;��j�u:K���%G8�l<�t�*���=ұ3^�ރ�8�49�Q02�ץ�HO���E=,R���_>Q����O���l0%㘒�;.��1���I'c[�d�	<Z)[u��X����.��C���
̴��%�"U�ȼ4�_.b�P�q)�8�����o&�jӲ��9\/��x�
D[���%��xP�oz3f��7���=��0�u�����7T��O� h���q��-�n����}��=gE����FaI� ����^	��|)	�B1B�F�μ�s ~@ =A�X�����R�x�F���x)�ب��B*S.z�9�)���|0����5ˬX�C(�i�m��6]/�Z�E��K�  �Q����Ճ��pղ)�� �)�j�@%a�-ס��Y��-V�u�NBEG]|����?: �y���-ITE�^�\e'���j{vz7��S6(���t��h�z���9(��-���R��z�)Y*�h����xu4���1K(�Y�H�6o*/2����d�k�:���gB˔����IDP���bOX�v]���F|����<����EۀG>�芬��V�S�C�q��(%mP�H+�󈪈��2Ь0V����=1���,b|�'-r�h��|�FՎO����tT���wT��	۰8�Z@���mO�䊤��'�{����֌�L�����%;F�z�+:џ��JE5��K�>���:�4˷ N[Kg�gx�֎�;��fqq�}-|�bg$�W{_��h���w��tO�D�E��@�V�3&�Q	�6�/�������y��?!��E�*������ş$�v@ɓ�1�cR@l��8A:���2�ub����0����{o���Z��V�$4�,�f1�A��+7��⌆Jk��|�h9��D��bJ�Y�|c�>�xz���9���G#��E0�\@���������5��A�W���m*-F@8������r���c���	Л�����v��EU��q��I�f�9eCM�*ݓ ,k�)4��Q�d�h��"��EP�Ś�w�y������>$dk@��=>�9+�Hc;�	!�ʢd��^	q�0��{�F_�ܬ����+}]12 -a�W��Y_#���#?�X{�P��*{�-WQ��^H�$���mó��v�;ȑ���"����Rz���"��ڟ����a��)�D��}W->i�a�(:�O�v9փB2SL�dw�=yK��l��'�CS2N�;v�08+`������ �ҸE�'�P�v���[�{D�7�2�on��FucOѿ�� ��MVT��[��XI��!�j��	�/�u���4�o�9?b.����0[a���v~�p��
Y��I;��:�Zn$Lp .���\x�h�*i�Sq��P+�Q2HͲ��q��/8���W�H��}�K��a}ôa�%��/��[�q_�D�TK�\�� J�&�b�W��t�!�)qvB����2 V���:B�ܡF�n��+�'�oMP���9��M���,?�}������mӫz�<8xT|[�$K0?�p��m�Ge���9���,8�&��`��Y劺�E��DO��8ׯ�"��?���S�����l�R���2u�Z ��2�-����!�۴ۢzK�6 nm�u��Ց�7�C=/���}�ش m�Sۊ��O5�9 e���=ׅc�&z�(R����t����wj7*�M�
�j�.���������|ҽHM�C�g�Z����3��8�_�c�ϡ�I�����+E�"99=��jD��9�����O}�g)�V ���v��ˀ�R@��R��1M��{�����h�]T�'1�	)C�R �޴�L�6���!�Y��.��E����BW�kx��Y�av�_�ϐ.G�4í"��K�9ޡc�һm�,L�a�Is�s�+� �x�}��E�e�=�d"
���Ӯ)X����H���f��M�O^m/�ln?G�j�3C�	i��6����.q�ba'&��+ߌ��0��_�Ѡ�d;�����ȝ��N���-%)����L]�;2%�7���rP
�=
 S��N+�"��Ȭg|)Oi���]u̜�{���&4�<�"�e�s/6)FZ�9D��1�,��?V#��]x?�����, |m�����j/� ��bzv< � >��09h�b�)Q��Ҳ���S$��#K�H�j��IPя��i�K2�Wֿa�$��Cfɼ���E��_K��atul,;7��`Er�f���5����mR� �����e�Jn�"�}Χ�*��U�)�nV�l�����������s�!�� � \S�|���K�/ɘ�e.�6i��n p��zU=.SS�̷��?U��ԡ@r�)�7��E	R����XeB*ؽ�,�Ǭ�Hɬ��͕X��U�V|��`C81���R{"h�����x"<���>�P|ܶD��C3��c�)��Y=7���_�.�޽����#�=���.Q<l������b;��{/�I��i����lI|b
�9Ŋ�"����[W�M�R� �1;����hP�@K܍�iO,�Xd�A���5�V8C�q5_��Bm^>*t��%�D�/�9A�!���0��4�1"��"�j��zl���юvo�N$�`��l�����k�<��Y[3�Ђ(��2jD���g���up��Y�����+$�;��BX<�f��B��^�?��V��\[4����	��	�U����48�p(�S! ��Y���Mx�|���Oy�e{+Q�'��%��Mp���e�A���z�YLqt�SaAu|��<$.���KO~'�0�����Wc�NO�6T�B�_?�:��K�k�����i�W��hړ	�0����|R�D�G.y�/,�5���=�,É�D&�nk��Sl[��~�s,�g1DC�6��q]�+����X�9L����(�2M�S��C"}����D�[˵/X���9_��m�L7����-�$Kg5�L]5�ڳ�ᙁ������l/���Ҧ�o�C���lhǔ�l}�4�H�`xw�o����*�G�I �^��/ov|ؘbM���`: �|5�dq�A!�Ll���U M�J �|_Lix>�ƖiB"��q�9�oU�(�G���!�珹��ҷV��l���{�>��t��7����֭����3̆%�i�H��d��ō�]�EB�]��3��󤏾KpR��W�p>�9�C�O�X~cU]#3�ڢ�)���Kg��x,�t�\/Q��g���h� Mo+|,f
� ,����=�z��ǪC�|_��+��ϪP�`_��c�5dw}���#p G_��tJ�Ǘ�mLP�_�)n[Omc=���g2��y��C3��&��['J<B�/�r��qf�M� ��Rv���:<
��|Ƿ�z9�Ui�7��d�:��%��п�5�VH�Ƒh�ο�>�E�5F��qk��5r�^��a1��7~oI(����l�X;*mq�(d:,.�SG}9��&�0VH+sK!�D�iwxtR�%!�%_��RU��x 2�7�Y�w~l�N�q�����E�9:4�I��z�_���"Zx�A�K�����UGj�w��%+�lǥ�z��^�\����j�z=�̓J�O������v[Bk݄N9h�A&���V��{� �P79}�y"�OI�5�TQԛn/W+[��)&X=�k���
�y:��Jђӏ�rV4�5�)������M��R�B�cx��Z%݆�;^���0_��ԋނ-ȋo�w�Զ5(V�MP�E�;��}8ߞ*�3V�!]����8�(0�RLe�pb�/��u+�##�Q.��f�d$bXhQ����@����i����iOel�ӟYq�y	���$ԇ>����!��]�B�����]�D��"S�7��(y���S�E���>�V����w�^�/�GP�v[�S��	 ��ͺU�sANhwI��{9���n�ܕ�cA �=W���Q�W�l����	<� ������z��}OZ��P�w��4�l��Ap��~�4wz)�}
@��IבR���8����` �WOYA��*��J?��D9��~�Я<��gèq�0|�gѠ={*�<l �A	���ӟ�v�BA%�����4�V���4T(��)�[�S�=�+܋�%����ەB��ʶ�!5�諠��9w�X �������$�:���%�v �!WFε�#pG���5�-���$�(�ުNMM�9��u�cb(*�c�Bv�H�t����&G��;9��
�o��7v�GD���&�	�{���]��D!z��HY����!�>�<റ~Z��'�m$YGʶoa��%�ao�O�Ov/� �վ;���
��D�/�M�����礪Qd��'�E3�Y2�cjH�)<���$�e���N"��c��^��k�7m⏓�4X��.�����-W�Lw ��h$'��B����8��دSw�.��V����7uu|�%iҒ�O@�������|�g�\��7VY��+���<���_�!�״�Ȧq1�%rXp:�z���*�d�S��*�SZ��2��MJ$7B$kG��Q�Y:�{��*��ʛ�
쇾��M�q�Y���*�g�+.����H��J�����H��rY���Ȕ*�r�N��+�U;����@{-N�XB������<�T��/��P�%L�w&C([�w�N���n��$K4����hx2N-��	�\&�n�O�F���3t�E����LB���o(G��.���BP��(Χ�+��`ℇ���nwͪV8���!��;�@#"��09A�xN��kV�탔���,f��i|�[\�dHe�%�+�x�:E�cTr�6��w�ta"�(�?�A�H#��6M��Ny���]�0�r�����B0Iq�np�!}�,��Ì�+���g�=V?�5�6��s�o�Y2�R߷>Qt�q������	l���������R�ɸ�WJZ���.��� �*<E }���М�J����w�B�J�[�#�JETK��f���=�%/׃�i"o��`���z37���U�D�2��kh�c�q����o��9�˃xc��J��}��~W���̓q�QH��qM|��t6W�$��~�@���}�:b�S<��5���ԥR����Re�	��o-���g�G�m�hߒ5-O�Y��P�~bPԯ$�@��7KX3%9����/	�w���I����Ղ�sW"Ş/y?h���UO�{�{JwtĿ�I*2F韤O�+rq�Rm�Hi����9�u���;���w��_�R��b
�C���is�bi�=��������e��7x�O�Aw�Kz��3U/�:V:�]��4�9<�H�t��J���U>^�>;r�%B�o�AY��Z-�ؔn�3���vb�q�� і���~O��r!���1�>�n�R�(��]l�����_l�/����*�4��=\����O�꣩E�;�>%�O�(}M}���/&�ŊJlw�$��֒wɦ����+�1X�^6n�I�gRrd�j*�g���T�Ih��P��f��� 	#�!"M8ؿ�>��:nw�Kn��L��Q�Z"Bfk�
������O)��/�D@.�Yb�Ɩ��n������a�MR̖��Y��|�)ɭ��#Ѐ���Q���!4��g��֤��j���	�r	�8�F�wݖ%�sv�����ͻ\���!ű3����j����Ɔe9��p�t5��c"
��Y�T��9[?Qh�h:��]���fR�����B�RWs}8�X>��/CAό٪R'��J�FW��:�\=Zc2���d�a��r��t`
�46�֔W��:�EJ]M����"�s��t��ɼob i�
������#I�}�.�ݲ��S{�UC����e���.ðe�?P��Ƅg���	:��Ө@g��Z��<����i����c��屶�ϵl@>�#��#ޓuWo�٤��&�1 �)PQ2= 2L�E�c�=ɀ�/Bi�;�K#Q�zŧC�1�5%����;���wE ��_t��5K'�M2b]��Mc�-��h�GS
�ٹ�e=�#W�������A���_���pd��$-�SL:yqnpĞ�5��t������� o�֑�aU�� ���K�����%o�$�"T\HKR�*\6�C�Śf:��5{}��1�+�2���5�X�Yv���ۧ��
Nu��ʯ�o�a`U�����L/�(���-��ĝ=������[� 6��ޘl`��d#<�
�e;��a�L$��6�H7[s\	�s���?=���EH���b|�ކ��g�wE�K�d50|��bd����c����㐚��9�m�e���Ť�,D�,ߡ���+�ޥk<�D�9݋
�cj����1V[�w�1߮�ј�45����w��ۍ�܍��@4�8Ԡ�D=oϤ��K�Y�ND&��m��{;��m��ً{'�_�.Y�h����>|5\���q�iMm�dAf�Q�O�^+��O���K{u�u����F;p{�k�%:��L�9t�#l��1T랠xY`dx��֘ۆ<mpq7��q�,�����L��ln"ж�=���������U���tt*�M���Ԕ�24����Qͼ]D�G�N�v�/�2-i�2ﲔ�u8Cg��F�ʗk48_���� B��6�8ь��)xך��KuI80x��Q�Ѐn���Q�`0%V��T&������A�\��JL���ao��b
�Ys���yw�v�]L���]���ͷ�V����ݼ�&ڥ��:�X���ɏ �FVQ`��4��D*�J�v\��TX��\��W�����]l(�V ^�"^��y����Q�d�%�ӫS�9q��nSb��V�+�R\SL��(nd��s+>;U�P��N�Ĭ@)�B]�H���^�m�#m~ݔ[�k%�*�5�ƨ����É�A�G�`�`g���{U��0�ېC�d�µ�"�gc-��o�Xxg��?#�rK*���Y�]���b��<����8��4w%��B��
Ίm���O�t������ �g8/w��W����5��O����qF]%�M��"�,+�k k̺�}@]���q~�=ہ�3ACvU$��RLzͬ$j|����7�M���m/a�Z[�\d����GL���+���Kl݄3��J�k&!��p���^��;��Z
.��4��^V����I����eą�dԜ~���bG���+G�y�J��B�$7�������:f}�Ȣ>�����M�׷�ND��h2�1~M��T�:_����ar��)���*l�sVc��dGY����'G �,��9	��nK&�H���� ��D�Ȩ�@d�fܽKl�ˈ���B֦�6�ڢИѱ�4�j�fn4y"%�$�V�0����݁'�����2��\����������a���, ��KJk���ew�1Zx�v�F�q�Ҕ��=(����k$��,=��)G�9�/E�Й��O��6i�r���崭.�� e~���.���12*�����	A�# �v}o��iV�b����'�6���+�}����x�������a���ؓ��Si�ph����K��	�
(�`�O�jB�e�<]���.��)GT�ԋC&��Eic@�O���ꏇ!�q���cTP��qf�G�u}���==�?�i�Ы�a/;{��bl�.N��D*c�'S{x�Tk~��%u����9n��O̃�X���n�@�������]q��$�Ä�{�D<����UY�̐Дi�mF�)�n�͂aMc)XY�pL�"�Զ<Y��u1p��m�Cb�;�y��dѾj  h���Y���x�=�0/�WK<��P{B�uU���0�<u�������:��N�f�a������"���57J̗z�y��>2�D�E,�oM��^�TO1W@x&�������0\��U�?�:y�v�yo@Y����ˠOF^M�8k�� �=W��}�uE^
F�/a�ۄ�W˺L�*J�q��%�@�h'��Z�B�33�"�,Gh���+<!�=�c�� )��mH��- v���!���E�N���
M��e���-8߀�	Ŀ�X!KEz
�����s�g�;��>#��ƂsT�����k�������
���Jf'ʇ����eER���&��I��6���ץ ue���=�He$(3��X��R
��o��X�yd J�}�^���|���lԛ��P�w(�����A������Ѻ�RL���xq"��֙`�r޽4���2ҳ�˝u>���k �4�+]Ƙ?[��$�	6l\� �E�Y�1�j�Z�����Z��0���)��0�+:��)	��w[�G
�>� ^���1���ۂ�v�W����]���I4p�+ş���	k���ԻcvN���zLyz��F?�����א�Ĺrڪ=��C�cl��d0K�)�έ}��x y�8�H��ɸ��5U�s��pj�l�D$~�r�#�e��>�n���*���������)���3��a�c�����P�Z���$�^�}���WIY��"���8�\���O �)I�k��Dao5�^Mj�FqGo�D{u����ɡv���� �C�$���qٜ�ǄC���|��h����<��ȳ�bd�V_U-x��;'��A]x���n���-��ɘm��y�w�u����V��[Z�6M�o�"���s�a���X� �S�
Z���g���/��ʫ���j��G��}����ozq���'�u6��3RC���k�g�t�[i����;L  �%��:���u�ل��g�FKp�is�|Z�Ʈ��ՠ�اT�=�F��m��K�����[�!����O����.��T]��T3�{y�د�-D*���%U��p蔅L[/�m1���H¿/��%�\0�0[�j������|�kNR���G�j?X�_3m~i�c��N�mu*�rV��	}.&�7�q�s���y��na�{�/��9Y�7�kO(p��Q��`u���fra$Itd�R�����Yhs�^�[)<Q��PV������?��A��7�f1C�7���4i�5�}��Z�b��r`s���x\�B��w��������9��@J�f�ߒ3�c
���s�<T� �;wCj'ςX+w�c~r۝�XZ61�̀�jS$-���=Ƒ<���N����K��<�w&yZ��/v��9��m}\�(p�G��
��g�ݺSD�>hG� ����1�,ڍ��j����o�F�/d�Z=��gj8��v����95�vqi�Ϥ��+��_�3z&��h�n!IàG�T���yo/�n�Vs�����d�$"ʱV&#O�$��t�r�ϰU)�A/x��2���R� 1���*�Q�x ����x<��4�5M�ۄf^��]mcH{�ix��1�d�t�\$����βE�DJ�Gz5��U�1f�  "V>7*~,�5�N2��!~;
 �3���-*��?�K��J]�n�X�V��<�a;�e|��>�{֓�B@_lfUa5]�m�ɬ&�O�.	��L����O�0�ܒ��zkZN��(��R)*� ����G9u�TD��n6� �Iԝ�-M���g�9L<����r�_���)���I�W�� 4��l��Q���p]����*�*;�M��c��?3i�����X�3`7C�MI�z���2��p�����6�۔q�rM��k+?%i֩5�gZ&�6vHjd �A)�kwJj��a6�f����bÑ=U������>�Ӈ�����c9��$f�+�U�l����0HZJ�0���Ki0�ϴLS��p�(������	� ��ť��aߌ��O�b�%�37ZD���텳���̤�4�s0}��([�588zx�'+���p��y�:2/LD�����ۤ-���F-�I�K9�9S��Xb�Z�=t�E0�Jc�N)�47S��'n]� s$\{{��(�uK���KQ�U������J�]q7e&O�	̀�ݽh��:E��� <xT
�t8ݠ,����}+=.�͐ٳex8�U�e�S�7����Q�;O�,_�j�6WE�,����Ж����&��|�l.;|�����7!9M75�.�@;:�p� 2�͐�zs�A%���UV�8/���+k�wT��
��m�F����y����!�P|��{��%�HQ�N��'�K���f� ǆ��Iq���|ΓV��$$Nr��b������#ux��_P�b
����,d����,������@x����H�ce�䞊
��VH����Oģ��J̵���9c��,;���(��?��7>�p�2��kj�v���*J��"�ɠf�
���(0E�H��F �}��sdb��F{#�U�<� G�Hx�]̩�r�z~5�e\+3}��d���Y��rs�7o��؏�%yP�o�z��f6u�ҙ%��(5�W�t�4�0g��:�Ц�פ`�7��I�����y$6�W�n��JBA����	̚���T�Ij���n�!�H�
,�l�aC���J/f�l׼�����%��e�]
@����mQ�e����nVj��[��%�4ס�Ţ���ə�
T	�E��$9��!�Ω��!�q���9A_�+�dޣ������(IoybZ~z�4����Ǌ�����(�S� �Ҟ�wZD�����M�j6i�8��k� @�Մ;TA�z�=՚������;�� ��a�ol~Z�="��rZ�� ��"����ݜ��=���'�Q^�~���BX�ꑟP����O�՜壐�Wڈ CƋ����n&�\�99�2�Ld�߹�Q��{Q�XKKzي�;�{k�Pǃa�s	y Z��^Ϳ��G���_�	�Q���k�R�M*ћ�3��� ���m��+�c�Z3� �J[�eǹ�i|�yc{@6������EB`�#�m|�Z7@ހӜ��sf)֧��b�N� ����ާ��l:Jhw2] ǭ�����;c�}@7�u�	v�٣�i�PF��*Pq����Ovє�P�#r3�Pr�k��/q1h��k�fc?�Hu����
�],�)c��Pk$H6�Dci�h�@�$�Ç�����+yj��藨���ڗ��e�V��ͻ0R�u�!E_���H�y��BU�r���Qo����_}���y��B�
�~J���,o�M�V���̰���]!�pl �]!AL�}�e�~����+�M
(��ca�i�2��5~�c#�e���e�I�5�"�^��"�V�̮ي4ڛb�l�`uWD0�HX:?b�h���>ס�_!��MS�֚	$S�*�o��a%��o�6��V	MF�8~K��U�К��H�t�3����{��tzFOrD�S�z1���Q�W��<۷����K[�Q}>FB�����C��	�@��Q��wVG���P�C��נ���g�x��wQ�1�|@g���O8�����j@�VU(��~����:��-M�2΂%�A�[zK�����F�����8���d��2����q
���^�d+��(�3��q[FՅ�šy��:���E*�����á��d���6G���������]zCo��p+i���_4f�0��*EՏ�yh��I@?Byj*�s�E���q�PA�J2��@T_Q�R������\�c���:���n���A2��YF����Ш�\p,ܬU��U�/� �Nv>��
w�f^���L�RM�v(� ɦ�xB�r�`�Qk���aqś�hF-�le�$��䑙Q�-��ւ�����K��?ub��������� ��6m��[U�6��%X�x�������@șE
n�xi1Q��6��6dKE���юв�6��-�Hl\�r��î�G5��)�o'�1$r�rd�EW�3�`�h��7��!�'!C"��S'\�˻�w9�-]�ПP�&�h1�c(���/_���u9���NU��<�w���g��"��G�RL��qUc�L6�M_ن:�O� �����}���
����_��aV�@��ٛ���Np� ӱ٫�t��	�Nj!H�fn%fŠ<�ia2XY)��J���%���0�ҽL������(	��z�s��w��8�T�L�L��=NFv��h#N�I�f�a�����	
\�F{Y'�ꢨOWp��պZ��~{�85��?�vC�uu�:����뻯iZF���[$��V�]���&0)���t���ċ�9.i���|A{2�8�bۄ�θre��4� �����p
�4���X]�0�f˧���9(7��؉N��1����Ǐx&Q5FrU^婼��4�8�x�?���ϻ��~�����d��1ۼD.�
�m�ĕ��^��HIU�jY}o�:/6E}9O�?�I9`d�&SlY�n�x]�!x{���
 .��g@��w�G�?=S7�vz�
{a=iR��ձ��;涋�b�փ���"�����9��A%pX�q�����6�N��-JIL����Zg
�Q��"lI����R��S�^�s��*���(�tDE�-{��
�[�	?��7޺�7x\�U��{�DgkpJl��c���;�]�t�ݜG��!Ku�M��;J�S�| ����^���'��Sr�m8��#�5rRɉ��|;�ie\�\��U��kLlA�il
!��h٥��;���ls�)k�J�`�ǝZ?dO�Z�U�J�¢��S��i�&��h̐"��JM�G���^RG�:�-t�:� ��)�7&����84W���/�/�Æ���(4�,l:�c���c������W6o�`��Thּ���r6m��x�������EI�"���e'�����ga;���-U�.�7������D�����7����Z^����3Jڠ�� ��ńӮt=IaM#� ���S�od�)5$��t���=��+P$|��{�2���O���o��/Z�!����ч�O�bܐ�	q���ۘK�&.t����D"�V�~a�\�^pD���̄��\t��S��K�@�I<@<�@2���K��UM9zB����eb�^Rh�b�χ��-ԗk���`�Z�\T%�F)���T��T�\��"H3v��*��dik���ʌ�ʼ��S,�p��82�5��h��+����w�=���]���������P_ڿ3�ȭ�%E1�}�}� ��5_������_V���O�p0���|
*Te�*)��i�:ՀډS���Y^D>�
/A�o�3A	���2�!\����G�3���Q�*���.�m�DOv������ҿa���aGg@�_�����lyQBi�@�.�l� �M�����WZ+�]�P%T�+ƴ���U�Z��櫚�ޞ)w,#\��h�2�,
��^4�Te����1�T��yv��r��a'���B�%�i�b89��I�F��=����m�jP~���)x�ڂ�	lM��vE=�m���L��p��pK6R�
��������)�g:�T�[���v��H�cy4�l�Ӏ��} ��HR�5����G�ɬ����y��b����y�T.�}W=�cú���gwdו��NVet�����N2?������R�ޜ�oP��u�J������G_�6�EKU~�$���H�	���2���x������Y�pҖ'�/���s���G7�R��$������A���x9������T�Wך��r��QY���dq��f�tk���6�j;+�s�XG'y{�S>V_əH������A]���J���3B���,�x#��y�ίA� �t�N�&��7��m9���j޳}'�b��b�0+34�����#�+Mx�Óo�{�~����_�
k��H�<�!rm0>�!k�҇g�!��#7H����kH�,r�o$d++h�X:�Y:��%%�*�V�MA�Y�u�)�� ��M�+a����t�u=���܃�ƐW��7��r��'�����7�f]Q�8�zצ��ʘ��*� A��c��D|�	\e���ƤūMa�V���K�B~����u���D`fU�Ց�߻�Uc�֮G���(��;�Yfr�3�&��t�)����ە�%�/��REދ�Wȳ�D�t�Y��ޖ?���|\�(��`�S�Dߵʗɧ�6����Ac)�|���J�=���	OT�ŵ���Y&�C��'ƞB�)_m-��0bm�`�Du���6���e�[���e��Cg�-��Tς�6@��T��j�	+L��la����Ǟ�h'��'+sc{1�j��Kw,����VZ(]�5�� AjZ�J
^�233l9�(��S�N��ǭ�W�.f��r��lB��Qk�q�n��%sqiY[5qHwF��ȕgAq\t��y�m��~�L�-�����z5Хf��; ��k���olB�6��:�}Nv�$�s^��/����YŶ'���Z|U�N�;�>��O�2X�����Y�ӷH�g���$O���Wz�'W"(l��y4n,mk���~2r���>����HE{����������)�s�����;Sll�TM��"Q�D����SM��n����L���s�iB0�M9�`��22�=���z8�#n��j�t�����L��~6�N>ȿˮ�p�I�)d{{���6��wt��t�e���J�u�As65�����E_��N�:�0�^�طb��O����6���r<�릈]ݮsӖ=`��Dʐ�c���8��]�6i�-�>sp֝=�Ў�@Х�d��w��+}]��*������Jl����S6O��'���^�ᚥ��ѱ˟��}�᠚�'�D�޻�������qB����<LtN�X^�y���^�f�A_[�\$��O���= �<��&�������U�8�)5�1�Aw�[�Ğx��}�	O	�~������S�Rex��9�I��V�O��؊<�L.����M��	�����Z�&:͉1@���R��q��~��$*o�o�uU�E��*:���G:�(����}Ç__��,�]��C� F�9ʔC���1	����v����)��U�co3ʈ
 ,�����8��Z���;�{�i%P��%��h�ܬ٢�L�,*����fGsP]��N�(R��ފ9�w�Q7�_>�҇�Y�i�$�_de*K^�;��x1Z;@ ��M.�ȩ��� ���p�T�@fDu3���c.-=��Q.~i��V>��h�y���5����U/��42@�&�Dr.?/8gػޮ��H�ߥ�@M"��ƴ�Dw������㓂�-�v�8��}&����T5��[Wo��	��Ԡ@��2n����6a�[L��j�o�H���D-mNe�]ۊA9�U�+����!�4�z���hϗ�'K�!iG1�_���3�nL 5]Ǻ� �Qٿ�a@� t����ąT��+��6��� �<�4�n"�~ϵ��ݹ>�Bd*�P^ZԷ���?t~O�_W�|`�ɸ-�1Á?�?#P���O��A�$�-5���5�p��k�h�)��CE%1�F�n!m���3d�2W���fD��?w��K`f���}e/J�����]-��iG������N��ؿOd"�\,�i�����A�Iy ���[M�Ř�sm8��2r����H)e�,�5�n�{��`W�����][�iR^��\t�ٌ��c(Y?Ē�������P�b"Vи�c��L��L�\�v͘_��G�����]���=�Q�Q��B�4F����O�,�ݛ���+j�C��T���V��y��cd�j��v�2KZ2ȁ�B
�)+�Hr�����\��B'

��=U�L1������Y& {O�)֋A���x���c� �1:����#E�j�D)7�*;I�[��M3�sg�M��v-�S�wDF��4�U8�y盜��$��1K�/�a����Q�;AIs�C��p/G�ɕ~��s�����J]yEA��Kw�wWG3y�6@�ī)�Ǡw%��H�M²wG^�$+���*�;!�Z�m�@1��TG��ghd����АDpE!�;k�5u�4��1;�{��[Om��y��{~K�_z0�w��'+饢������&#���n��
n����t �� ���a�6��9��T`Q�b���+*�Q'}O��4\���kbGIv}�P��4��>e����%�V���
S�
�3��e��(��])m��3ݥ�7Ǧ���f�6EF��-�N�=��qC���wK�d'~��$[���!z`�?(U����ޟ]o�̆ee^%8�&!ca[{VP2�V��!GaazV��P�֓O%m������ai�����Vê0�~=�F����?9E��"���~�y�i����&���#����6�m��7ks�l�����3��w{p��B�����[ͨ��&,�HI���������6����Wdɪw�H~�W)��AP%��<˒̡��Wވh����^��Bh4u�.Ƶ���B;i�0��_��d���(����C>���f��)z"w�x^��f��@�� H��D�l�ugݏ�����׃�6��KO�	>+��NtM�-��s����LN@�ԶT���Mъ���1��5�)��1
(�`ꢌPv�E��8D�cυ	�*u�i��R���s+�+���%�u>|�pM	R�ą��p�h�
H���M�dP3b�3�� �>Q����b�H�u�ڑ���(�L[A�xU�,iշ�?:���ꔍc�Q��뇈��!��V���~)���-��L;|�6�T���-�%��
�W����+g;lgd�޹�'��I�s�4�Ƙ�	�ޜ�*�HkU������sJ`)�ϟ��u�HKZD��v��j<�g?�D� 	)�+�O�WSdR���A���&㰧��]�����UO-�A;�4!���F`�#+��Xq�'����(E4Z�`�g἞���tK?Zl"������
ݿaY����|;�rf��V2�������F��n���:1��w]�V��fk����V�\'�)s�@�?�a�����#�!㟥������ -)���p^��e����j��Ȧ�p�4O���h��� �g���.���m����
\A�Rm%qq�����Lg/]�*]�󙔏!��p��ܖ�Cu���J��J���㋤�:UHP�  p�BI��x�IϤ���=�R(���""������� `��]���S��Gh��V Bf�h���7�-�&�/Gӄ�`x�f�k�8ڱ��Ű$�ZZf�^8v��u�j� gLb�.�3�3@���/�UZk:���k�W(����ؙ����˰�rlJ��.X�xZ���ç�4�aASo�+��G��K6i�� �{�1
To<�'c{k��ݶ���^*��A��-e�V�$��7z�F/W;�;�T�P"�{l�Ƹd�2o��=��;),c�̾GӰ�Ъ̖?4�|[0F6̯O������H�"�2^6*�:"GH����	F��]$�dPX�/j[�p������2��B���d�3󘔗zZ�=T��F(Z�F�H�s�=#�{�T�g�1�i������H�7���PJ�m|?Aᅖ��3|�8!��U��8�"A�+,�����+#�tHʚ�����B�/W5���NR��X}��%�2����@� <�;��nF�+j�C�0-y�`��Ig?�����^� =p��e��8u�7���B.�����GL���Ϳ_���
~�Ni(�i@+�O�-[��,�����q����dq��{@����w��P&7�t�4��h�!�-b��l|/����MtPY��G\�����������2�~��Z��8ɞ�y�|��x�����O�(�tk�#(ȋ�ّ�N[�����W?��}r�@0��2��7�Y#��O�eeƋ���y?�ܟwy��w��
a�����8���Yb`ٓ�f]�i�j������鬤�Q��0X�T��W@�~c�#��[ ��t�9^-�@��Y�E>���F������V���u۔4�O7>�4�J���rl�R��V��3�j����K�o��g�h�6x��k��Z�Fê��VfUQgM	��r�Y9�0���Yl�*�����{zTG���:�dӅ�o1X�p�*���ƣd�%��="m�����>�����4��~`Ȏ�r��fI��˴�x��Z�c����7Ȭ�>X	dƤ}��ׁ�"g�q�}fD.�u�����=k:�y�i�_�}��-mm|�fC��;�
{�M�4(a��H��FЌ���O��]Dx~�J�Z��I&l9�R�%1`e�X�L��QtE�I4��)�h� WxAC�HW���Lsc��;3i��)d+�f�y�9���i2���i���yĊ�71�.���+�ME�}��>������ƹT��a�ؘ�(:Ϳ��U���<sI��>+��O$�:�ܢ5������㙣ƽ���?�RG��e��l�Z%2xݔ��<�G�5$�k�5k��4���:�C��6<@�h���
�hLM�(w�2k����*Y2���`��Jb�����ė�=��8<\=�	R��犋�	;l���_��h�3�R&,��EM�����k�2<*ۧ�8N�#2�6I��o/׽Y��ǉ�����9y�����w�'�d���QQ�6�H��<;����<i�J^����ւ"�����I v�[�U,I���s��� t����U�-*s6�Lnx��:�I�[�1�q��#������J,�ꦸ\$��@35��Ù����5i���;"�����a,����(��9D`��Ex)�E��}
�B#�vL����@��]�u�Fap��'����9�C\��P��WCw�Y�G�AD{�6�����ӥm-/�1N�����g� *SV\�
h�d�����nV+G--�H??�U]S*�fxw`F~�0֨��P��m��uq�F�4׷s�(X�k�-ݧ3�˨�� ��!XZ�Q0���bC��8��	% ��2��Fq7��6��.�Ω�O<%��A%�[��JDڧ��HinY�3��e�^Øl�q��b��ڙp���tc�.���4ң�.^'����Ӱ	�	�=�����iltϕ��,!H]�o��]�F��d'M�>�_XC��bV]��E+Zjf����a
.��y��T�a��#b:���O,���H��*�y�jꄯ@)�Xj�}7\�t	K�S��6�|{�����`DH����w3<�%�9i3xz����c���|�9R���lHޝ�r�wtK^�5��]���^^<� ��:fLh�v�	NL�bcD����6��2���H�ʾ��_���s'��5�Il��(뮀#=M����4�sݤ�l�:����CI���)c�A�wé������D��1,E�S�0�y���¯���T��.*�̝:����hmb��+���%�F�_��M��xZfV)�Be-�A��M|xB��g���� �!��%j�������� �I[ʜ����S��ܯT�Ar3?/؁p���o���}�%���B	I�$���h������K�flc:9��vo԰8��]q���N&��Y�"~{a^Q����(=�J�s)���[�_`�J2���>�A�f��U��v,�zL]M
4N>(OBj�`��5� ��nX�{��\��m1Qm�����Mq��6kb��%r������Ee�k�2,�����P�=�pPO��G3�S��2�~(����B��	��#��`�E6
K´LB�x?�q˶,IK�h��������)0%��c��ﲛ��\Pd�Y����TƬ�u*SETB8>�X#ۈy���(�k�QQH�\�������L2�z� ���C����]�8]�Mj�����EW��}{��x
�J�X9� $Zy������l`�[���q�^�����Q��azP}Bo˳�#��#:*x�D��7g�'�p��Z������a
�\�+��=gr硐.,9�v����:H��@Z{ҥ��a/��Ά�=�l�В�B#݅zp%7�0AT�}z��!~-�*�A׏#���@3�u�c̨y"��;�'�ǔ��E��
�h�@}T�4^�yZ�ӿ��@Mw�c$��|�Tth��9��M2���Q����`Ґksk�8
�VZ{iuH��$����[LN�����;�e�6sl�p���R��q�$���,��Y�(rT���R��<e�nXe�
u�<��w�q@b�s�x(w��l��$P�0c9(�0�U"6G� ӀJ��55�^8�?Q�`	�/O���O=�o(�d������`˃�h��9H!!��o�[-0+��Pr��a���ߘh���w�I�����!��t����j�[Q��LVG`��0A�����&��[�E�A�,7&.Xo�Ѯ�.x��P�%�#/+�v��j�~b�W2ٕ��ց�j�#�b9?��Pn�R�J��G| ���s_�?������k�1��k�'J�=���4u�jl.��y�d[���J�G�N�
/�1g��>*.}񱯥e�Fo�>&�����mӼ�k�gt�/N#9L`ֻ'�{Azo��`C�z\��ڦ����V~�R9�"4�GC&+o;��@^�zT�3M�qI�y�ȩviBoBV~�Lvi@y�����ȑ���Z��ь�d�`idap�a7���}�ևaJ��OӬԇ���v[�����cj�EnU��!�\��+!�1�d�)E�ɼ�����Z�CPY����P?TD���ϩR�cQ%�U��*�=�=��8t�H]��v��c�b��)����Eo�ys�'K�q�;�g�) ��x�1F�ߌ;±���+vD^�*5n-he����
$fP��Zwh=�g�z,�����>U/h���x��e�,2�'��G��D���i�eQ�}���2����}�}Y��n;>�r��j���"�S�nΧUZ����N;f��Peх:ǫ�{��a��[�5ڴҷؽ�Jl��'�} X�H��n7��P���V��[y+����/��X�
����������I�� ,tCm��9�=?��WRm�;�s.��L1�Ȱ|����ذͽx9Q+|l���	���N�S�LoGX�w���̏�#��6��v<B��z���]D��X�!F6�K��8�B���t�Q2���z����/�F)xc3�2RQ[�v��{Bo���\b- �(��s.�e@@DX9�r�;�Y_A�]��v�(R�Ł,�4G&UJ����5 ������b4%�#���GC?�?)wX~fU3�
��Q�&�uE���nʤ@�ʧ�@��2J�͐Aa����&3@��ǫV�W;mH��-e��ќ�o�Z��ٮ���A�J����;�9�۶�����[���׋�{o��z_�?2شU ���4��P&�v �2��~�g��MJ�N�ڵ�4G��)�_�*��I:o0��f��I���������@ ��s�i���� �X��B���[D��R�-�`Dx��FA���l�\S�<���0�z!\�6y�����ҥ��Gw�x���tn`�O���\���p�����%���m��'�^��v�Kԁ�R�y�m��nMc5\>�ك�$N�hA�h�NU�v��T�z��VM��C��{�߃��/��6���c��-My۹��S�!��z��@�v��u�R^�`� �3���Ȟ��S��u�2r��6�Bu:����+��y"ǒ��-Ym��'\ѯ�5W��+m�-�K��ĿoB���1��X-u3R���vkgH������I�ޕ�;����H��R*�y�1���kik5BM�r�e=�F"S�.ڐܻ���+$�vw�##^� 3�Y�w~(�"W����=�_�fi��pT��25����/���7q'n��i(�M'�!q�1�r7��D��,*[�b��yLI���� Uks�� �l��B����M3�b� �Q0^I���@�%��亐Jmg�����s��D����~�=OZZ��]��A����.�E�����=�NUo�+�*��F[�9��S��k�!k��>���T�UY5��$I<CE~sl!��@��m��e���Mf�1�WdE�A����Q�ٱeQS��6U=�)*h�y�Md�&�>�{Ÿ������O����. �V�R�Ѽ�M�7� �֙��_��S(4�:
	�����r{&Ʉt.�A_"Wtn�Y�ba�lX��ץ]��Sʯ��e���v�$�Mqq#��&6�!��*Ǟ5��_p]��({�zg�͑];4�ɹj3Lse@ҀzY���tO������1~�A�z6��6. ��UP���q�T��?8�%��t��ӊ89�"s����f�����b.�ث��!u�����������e3 �<����?'�#���_�󨓓�F�`�����ظ�q�!��f>Π�����BJ�ο��A���r03�>Y�R/���'m
������v+ �}	G��
q�q���L���_F~��s�3�8)2I�|O�= �^��ظ��b�.9��u�
�d��fӞ�n���`�3��<� �拮偄�Õ5"m����`�w#[�����=~�*[��nZ�h��V��{��D;�+�ub~��g�hµ M�=��.�d�:_ T��u��6c
�.�\|�L���jK�{��7���V�t��a:C?�D�����^(�48Y.�D��y���-��f��L���ߔ�jM��G./�f�<WsАf��lT�k53S�2ME���5p�Wp}���?��د����#Fe���n�X��b$���������[%=��h=�ζ��
�m���D(Ò�R؄QxyL}x%Btc��o�2p��1����*�.�>���_}D����1��x7ak� ��z35E5�����qMo���vn���fy����1���=Z���>��T>aNF�- �1��(���1��n@�WB�+ОI-��V��oaE�qd̙�&~͓ �Lז��=�\��[��v:4��F��X� ^�SꤿM��z_E�<��{!��Gސ�����)(߉�>޽��"�T�qq�ι�����P�=7g��� ����v��ь��$�)�6.wH��by�+�o�Ig�s|��m�E�0[+wG��u�=]?D)�������gb�e"���h<]V�ʅ��Y��ˁz�?��ə ��5j�Mve�=��(7����0��;���ԍA�lt睑�b5�D_���pD�M���۩�z!B�V_~��2�C!3sr������_~����q��]���f�(���PNˤ���3�JJ}�������Ov5O��e���6��d��N����'��F6є�a�ㇸ/Es]d�� v��D��I�V>�Q�Q�}���۝�6�$�3�(5�6�HCm�O6�/�;����Ӎ�{R��w��Cu��L�+}�߼W7A������1a��RC����'��)W�D��������#=B(<x�0ߐ/���i��^��e��/5,������|y-��ɯ�"5j<,�0<۲�����t5n	�-�f֣�6�fI�>���X�>l5R�8�og;g���X~�vn_�g4��"�!�aq�eR�r���E��e�0�֒������Ϣ�H*���}�]j~0� n���Uɴ���u51A���O�$�qƝ����Ũ�a��Eԙv=zR����&��_7�V\%N�	_W��mQ�t�s�oc9|��Q��Kzb�'��~�%� �h�sS���������%T[.sZ�R>^�0�nà�pa~E+�n�`ryq�wL^ts�¸�
��㡯��7s���L�ζ�}�uJ;�Kn_ ��� ����?'}*}�_�XF��`40�������;� e�+����]�P ��W{�G5N{�qj�m2�4����,�8>�0��8��զi*9�kM��4��%�rD�"�x�XV���91���K�ׄ�kZٕ"q���<P�Yqi ��o	�����wx��)ct"�~�1Ŀm��(�-y_��5kpE�!�z��.�z F��{�}yHE��'�m�y�6��m,d��bH6u��?e�E��12�j��0�mFh����9��H W��0�i��*�|� ���^�W�q�_]��� &ip-�(���A��#������Зyeǃ\�PE����/s4��Au2�:ily[UQL�En�uQr�˝ہ��}#3�S%^���fr������:�I��qM���3f��MKM<Ь�$MnV��V�v�Y��d�	��˷��*JԊ��%*��Q�8����M,��a#VO
�P8�Q��W����O0��O[�^lGtA�q*�| \�S2X+���,�jg��ş\��:J���oX���(F'���0|��Xnf�T�,�x5��[��ܢ�5bd;{9%U�n'
I�Xq�J?��}+�C����NU�/�����J�o`;sԐ7;3>��E&|���B��p�!<O���I�y��}$Uk�X�|�.�4��ݽ���z�����S+Nݷ;�Y�oݳpW��Ò5��z쳳��?ah� �O6щ�|�U�9�-�gy K?hcc2Bv�W����F��(�������s�s�Θjs1�9΁!��+� �T/y	�Gl��Z����e���zW|
���/o}��!P�R��԰�q<�wҨ�t�%ǞSi��}��`��g�����o���TB�9���y��&��lw���v�R z���d�@�%�:�8��A�:��J���5
`�TsZ9����ae���#c��"86���^�^��Md$��O�\f\z@�KLڥex~o�묅��!pre��h��*�L�(�H��Q���ƿ�:���P���ح�f��Ux@�{E��@�C$W1c��̃��-^@�T��t�&�+N��� 1���1.(6����;�cr2��h�V���)��D�.؈z� Nx�L#wQ�zO��uP��y߁|Q�Vza�FM�;FnF��?�,�A �(������A�	LXj�:u����W �,�~���DC�F�g�U�0������Mc��b��ID���(F?��r�d���ל>kկhc�ҡ�)�n�8�_��ptP-
�M����B��su�� ��I���]�K����`<M��uگ���	B����rA�����n�&��7ؓ���kS�kCN����h9��O�3?�����K������C�L��ց2�7��$nFg��dP�h;��*]!�u�&)��;�ږ����?R�ɶ�C�!�w�71b�H#w�!���3OF�A����ą
@ܭ��+Oۤ����#�N)}��CO�F�w����H��z?Hbi�$d�����ĕ���m�=�8��E`�_\V*X^��$k�(n�H�P~;�E-�D~>�L|2F�޿=jm#��g���p���s����m�p��!��_t�D���ZV�}��9V�Z��[RZph����彺�-��̶R���K<s���rH��?|��P�[�^m��!Ü��Z���U[�ד0�wS�����R�ʟ1.6[���Tqȶ�L4����i?�=�w��'�� (p�����Q���)��R>�^
xsi)���)���v̟U�	2s��(9O�'��1Ư���&��[c�YE&>�_�uy
l,��laK\.�_��X�K-2��i���
�7�2�P)e�{W��Ւ�yh�}Va;x���wK�mm!�Jh��a{S�;r�oc�]q"�w����x��� _���[m�:X�I����:�����tC<`\M);�#�QvQ����\�v��_��� �ps��m5R��U�譟����6���[(ƴ��gz�镂���&�*X>]�<mB��	}�\����2� �a��g.�[3��u*�@NC~��HĹ�����O'<�[�o���Kju<�]`�<E��)��;[����C���ۙ�/���I���2�z��RԱ�� �W�<�F�t/�bճ=rf!�n1^ھ��!� �Y�E����m�����Փ�_"p���th�RĖH��^�.�9��>�`�+�q�}<�~�~y%�sc����nΐ�$�pjW �D�a���<�B�����@���\ �X��&���sX:u0n ��C��/hzW�&���Jy����1F�vPS%Q=�W�"���"K�XӸj�^�E�+�wO=iأ��SDJ�T���^nƌ�n�������
^T�:	�x�r��r��v(�h�˥�d�U���0�D�H���1��T�Ojt5��]��y��wE��a��O{��)����+�#�x�Ll�;7̐9�����~�a;g94%ۍ��	�1B7�C��z��r0F���v��1��NQ2A��v�w�O� z�31���XWv�N��G�s���[�ޥ�8tur�񚧗��f�`)������#�۔k6�f�[�#�V���2�]��f�����r�~��µ 3���� �b6�)��a��z�;�m2��]X��6�F���u�!����0F�[��<�K�˿Q���\�����bd)���Bw����yx�����Yi"~�;�G���1�P�Ѕ�߰rV�n�6G��� -����)I!0.�P`���zM��i7�ܵ�����z���q���t1�~�����Kq�3�08)�PL���P�<&2O���L�>)8#\]���|������^@��L��~0s>tV�iW�T2�#������P�SA �m�	�wISmΆ���W���ͳ[UBb,0�CGUq����۔�,꾱�&�\��
 �5�d�8]h���{�ZZ�Q]A��xF��|����5��h�7OW�)� �W����'�j���!n�J�Z$���2ó���%M��/Ǎ:m��:#����ƀ�_�[��I��nA��l�$4��J�fz��+٧oY�(*:*}���G�`]��ܦ?v�$ʏ߾8��K0��D�\�Oݚ���T%2��F�N��x�"z��*ǾR��D�����%���־��1�$�hk]�J��<�|�U�{Hߛ��A@��M2��(�f@�h2�H����n�/FWf��f� k0=�����I�,�7q�,W����y�[`r�[s��;�(tJj�j�p3��3�>.e�K��%.��Q�;3(q{��nխ�鹹�/��pP3��|)Z�eR��fw$�S��0����1�n@"��m���� ����E�IRU]3-�'N��{�W�� b��ܰ�=���P��"���bf����o f����hC�e,�m��>[nϔ���� Ӣ����I(���G�d�ܛ� H�=Pok�߮�}ǃ�#�L��vբO��Oa�-�r�9�����W�Z�p=F�B��.|���X���QA��/��<J�
 �`���4�)r�������'��'�F��1�`��:�*$�/��	�7s�A\��������!�,��Z��ߦl�q'v�����쳚�Ԥ�3�0Nke��PϪ�pi�� ^1norF:#�R<�W��E�vI�Ք	�M��P6ژ�1���*?gy8�8����:�%�ud��X��Hȯ"Ҁ���$?��*��Ɵ�K1ä�)�ֻ��^�	�r���p�E���R�0	�����J��M��q����ƨ�R�Ӯ��i����m��~��c��G�Q�bţ߫5�,�]���/g����\�����sS��a��|���D����h�>�M
�gk��1��[�vL*�O&,?���ɛA@O��>��-P>=q)5!���߰� ��Y�B㳼�����-9��"��u�L �����k�H?rax��:��xc�a=
J$�������v�A���hf-=a9�b�̐��h4��9�'J}3����r�+�@�������5q����{Or[�8����2�KD�	��_j�!-�<$��G��q���Y2g��N����.f�g勼l�d�!�9G˨*I�4�1ki��m̌O�Kԅ�_E�ceF5���Rm��n�� z�h�GO�"-N{^����]{���MsV��JU��tL��b�w,�� �8�=y��`5��2A�V�?i�};s��']��e6H�m��c,_�*�9tV3%�ȒZo���8�%&Z�U9��_CP��2��(�W�._nT�J��R��1�9RuZ�A�e̭@�]4�{h�я��L�3ah���q0�;�J�P�]~�Z�"�h�^j�;�'D��i6�ęmD*~�nA�+���=��4=�})f��.�2H;�g�"ٌu�	m*������kQI%���.��|{]��c���hဵQI�/��MχU_�0�h<YEV��AJp%�ފ�<S������ [�Ęu�����ߙ�v�꽚����&��n8j�ط	��*DdӇU�l�S\��~���;x�ChZ4�O�?�n��������hVz#���wk<ͬ��d�z��q3���
�'�i�܁������mZLNڑ�2٦H�~���Y7OZ�ǘ�Y��[�gU��	��G�*��o�������x�4H0p[��Xj
�����V�p�.��N�*�e�4�^����lH���<{!ߧ��m��{�+��l���U���[�2}��k�Su~M"�;�l�R_G�)P8�������F��e�,��|�tŇ5�w\ a�_�1 ��h��a$?����0� �ev�Ps`�#Ó����sH T<�	��	v�_D�\�~��х��%M��4�f.g?���!%�b�a�ȹ����U.��ȡ��}Z�Te������,{��v����,p��1�{��g�Ǔ�NCB���QA���_��)�H��4CU����h��2%��Ǖ�b����FfP�jr��x�x�RE������<\�:&�7�5W��)��-��*�7��Gز�6�|(/ou��);�'XL� �O���X�D�B��
���0ưz�K������϶��B��(b��iC//�A�7 v���k�U���.w���L����O)���瑛�刎��[q=��P�6K�P& k�ق:�����I!�}�{�M�X`�B�l��Yt����3M�ŴB[�"�Z��hW.��_^[>��O�Gܘ���c��/�(��qgד�V �]j"�@.�d�8`h<��`ѱ��T��ˤ�U�I�zƙ��!G�`z�fA��3]��)L5M��5�ֆIX��0�z�s���
Z�)�*���d��_���J3�]�7V������u�j�/vl�Y��W��=-�>�η�i����(1���p�5�����A�s+�'�w#H�@�R�I�V�u�!\����)�ܪ�����V�#Zf0���hv"xT�����6��&u1x�BY74Ƈ�nEZM.w�=�ӽ�����6�W�9�#�^.Xh胰P�%ř2��]Xm�i��{�r�pg��%���赟��TKlg�M����4�P�$������z�;�F�A�tOie��w �J�Ŵ���ڸ�U䧡���?{�_Y>� $|m>"V� ��%��x#s��L
�0�A-U�px��ȜX&zs�F=�t�t&{Np�[�>?�'-�jvvFg.^�7>a����(uc��i�Ǎ2��b-~�-K��/��j�R�e��b"�W�n3��~T͎����_]&����\3W膖��?=��Y�S�����n`O�����2���W�:�[�h+��h{=�" ��h�f9��G�]�M}]��*�y�-҅ޟ�W�zل�5�U��^���@�6��4����������$��]�Dă����{�nA��+&�� <$y��c��J�#/d��|���;W�Q�&�����l�Wۮ!E��ێ�CzKn���٦�e���@�ɡ�|�-6��*lJ��u�t�%^�B�n&��34_���8��ye��z�(�l�c�d��IPi���p��V�
(��Wդ��|�7Q=W� D^��7���Xӈb'^'��BtǮ���:0�
��u����	�0�*�Ӛ뼽�Y��*1���_�h�^�z����T�R���_�*���Ee��r���G��~�Ƥ�!y����:NY�t�~{�!���B�=;��z}In�{Ydԫ�}�w��7��G�/��]����dŵ�� ���O>w>�׭���`�A����6��́B�V��A��U��m���~+_�0B���t�&<���:c5��uW��3�"s�-9��0dȬ"�"呈������i����$�o��bb�},�ٌ�=5�Osv�駱$��Q
�� �$��`��F?��|�9� �sy�q4k�'�\�ݔ��7��I�&��V�����ޙʲ�ۡX@�rV��5�*D�SͽNVf��4�6��Lӝ���b�Ǆ��c�H��2���j~�!�e��.uBA=ϛ�-o	]�#W5��8sR�`Qb�/��HD�'EX!�v�w��Y���j�E���þ�"��-;�����ͬ8�<��C�Ɖ��-U��I���oug��
��mz@12�Z��;t3�#I�׉�l5h�R�u�����V��8L�mF�,�Q�s�NS(�����\v�F+`Ep��	)�[�̀�1�,���@hW��n