-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
I1BWErR9mXFwEuTQ4Ty5d5zHgAUoSbc6yzUkJMvz64Ed1wyPQd+uzMStctt5UxoaBb3+GfmbPWmw
V4732za8f7vt4EEPix6ajekcoEuQWav6IRHGU7WYrbSXOr0u8eyqkn6/aYkr7HjdfZzmws+tBw+z
ANFVhQ5wNArcBFe2Iz/Bp5AO3XGmkcFnwn/vhvpy/Wc0HrVJvvJxQCIw5OzGfdxu/eo/HZwituNj
5rtEhwHDVJcciVUJgc2qQoqhsApcP62B9lYdHcEhkadfn4AqPuyWzIxHOvfRpFeN20SFY9S1M9fm
NzzkGbaJ/D8FIReSendcvG8arOKL9KZoVVR2zQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14528)
`protect data_block
JI0cdTr9ZpcZeMQMFtde/xJi8cF7aNLjN6sFOiHs4sbfAQbIfkkMABC6/jTB8TTfNnFf/YF3iYMe
R8hIQ1o3D/2jnXKWA2AqDHDMaL9pnVJ3GWbORNFPi8aWQeJ7RMCI3ByAFqpyXpkAsOlu71Ef3y2q
LrIdNgKi60tGcDM7ipiaLIdzuJnIygiAh/jVljxJrnMBNJqbHT/gOHDUswaBf/DdKBX3PsDs9vQY
wlHvTtMbYPW6Da5c4C4C6W+nXZFdYri5T8Et/ixWKsWtMQ8n9XjWgHTKjgUBNguo/LXHyynU3sFJ
VuB9Hg3x3u1mwqy+wmYEzChmy7m/M/F405fvJIr5kT1seVtdZlrcyEdehZIvf//exDRYM35CjzjE
TJ8rGTCF91NZKfcuW0lk8CI4ksSw8nwJFBZL9VAEMpCIErzGW2ZAZ0XRwAcCZBM1/1c8VQehlwpX
k5fzvx12aro4XijdaSQEFJSfDibmwvjzoAQzJRM4LO+vZHkSvj0AFz9KhO2XhKYltM4K09x85tTo
3JoJYxr14ti81HcG07bfbFktjPv9WG+aXz7Mz6rkZ4FQBAagdeDchXtFVipZ+XHLBSe6SSYfOCXv
LIIZSNP6GPyXJlBiIRbZExf0NwVJ7cknMls0daSXNKigfpfhvrS8ECP10RLhYlL93m2tpU8kikys
Pii6EtbuBgp8kc8K+RSGFaQIGMhBSTRqiS5jQA9dXPpUPVB1Z84REBZnYNMvMBqlFIB3KzcSyKwC
9mfvjouKxpcdztxCX26GUiTLQZx7CLok++43geEPf9XS0IluY3vmGpLWvW5+3iZ1Ynajt5Iw1cIp
ePh95YI5x1PgzgNQR6JrCTQ8lVDOkyB2tQ5T6m3j2BvHsD3xLK9KqA140LMOVfwlJS5LkolDTBgT
PVAKm+B9O3bhsLGEscxxdLuez8Xw8q5FGkW/10sUHpXXZcRPa1mEb9F5fgeGHphGZqwPPKICaoeB
9QhEzgxupPySr35r2MNlPVrQWhxNw2w06rlm8nu/mYMfyQm7AXIiZAKFolwM0JQEvyx5NcD9OcLo
7PgFUk0Ro0OnGQz1irGi8d3HgmTjFDS94JCEQw7rIVmlSoISaTLXSkr1oJbqwqCMibltT/23eBW5
qXchtiAW2ckhehPJsY3F1AvX7ERkUoJzEDig5UMxD142KpU/o/fO8mfcdybJWzQWFt7V6mMYEDIg
p3Z4wH1DrgZNpicUmtuT1J9QjH7pEXKNpJbxwa404Bo+OFq0EAG6XLXYOtOG9h9n2N6FEfTSnu+F
f9r8NCSsf33n/8Y6hAc6fLt4lv9ZFxrklJQ1AO6j5/QdicN1Zf8SGOboL66/eKwT2PnMB3S+3H8s
2B+qqTNqHVtCSCi9xePtxz/WJRoOBE43R6brQR71lkTL9iaKQ8+Uu10fIC3wkJKGUWzPXH8qKx2V
jSBSvIxB8mafVlZGojwAc4DjpXEHabI+I3r+6NZ4q8RpEiYZcL+HTsxsr/2L6M3Bc/FZpbXF/cWV
C8Uwbd6PzqDJLrlgZH8eKLgdxU7sYKLEXuIfCIX3ohp9h6d8+Nkyd2Nw7ujEgJLnbpmVF3O3mOax
uK5++EMFohkPRGB8I2LUVFB+0TRvoHrXPdj1QF7WQzb1R/yTANwoTnSIMOkixCWdCasCc2KstAQt
2geoM/7TsVWqU81D0dN54RldqFc7TYMHgmMlzA6GwecKxVJeczN9UX2e30DygfWuh5EnaEYcITIa
JXPmeB2FDkC1t/03iX/BQU0kPU76v4asDPHQJUXHdXB1Om/S9oFKaI3Kpj4FEwIEt/d7wM41+ytR
x3evX7A9z8b/I0wBaR3TQjKcak1Qq3Z99JYnyJMtDuPKRc8lehon6FTzBZJe/GW6ancX81LcR98u
uytJnQhbraDT4jyJeap8y/K4f0rwxkYzb+YMzYBOjozS0uz3N3psHs+SS1IZIg/4Z3fDTAl8HtLT
xqjwV5zkmfGgNn0HwIog1tniaSVcVcN9suuWETTfy61+iSR+d1N7QKq2YZlI+/+nes0Er9KjgU+K
5DtGcCrI590q1TyGxbPA1q+bsA0X4IzSuMkivf2c/FoxjnjpB+d2J2w8Lg6BakegiZuhAVqDC+Cu
Cx0U5LoDfuziMO21V84k9ORo3JF17/hy0A3PC06OeJGcmjohySiRlIyIlyxqYYRbS9LMcb51pHk3
L7k0qpANimj3RCNCzJSlU1SS7l4oZLji6Wh3/4p0Gj5XntyzV79PKzkwpmHPWUqSEVqaAkwnEULF
t7LYOkMSMUYbxc4SsXytoDNQ9Syesd5jrqPWsqUfRXPW3PcfBmA+jUfF2Le6PutS2+mIHXnIJ++x
P2eNDrYkyvsixEHRJx5MzwiguHGJrqTm7Dua5M0BRLgl91m55C2aUID3uBsTDTNgtiorT5TuaCyp
uw1hVgICF62WIblWvq8PEJC82hPgNct8cw3NXFZYR/tmvgIys85U9mf1oYc9EdH8zCKsEKyTbyHA
pXPnUQs8owuWlsWe4YK1IeaHQ5tqtNEgCx0UtoLdUh0aHR7VAKT88Urx5XFgwS4mA43pFl0g0Ney
MhzBHTddmo5rcccuKJTu4D4iTKx5liEgTWGva6pmHjAluvBD/Jmc25XrvERUZ9C8JuIdZ31ow645
DfUzEfzFy3M5E24BgzhqTrkje1YJjTsJ4lFP9pRKXBhezc93w0cob47Tkou1c9q1X2gJ7zgolls3
IgBmQ99zx8BAfKdAfGgHGCi3L/k+PSfCmNL8IQDw0efp+tdW/k1UciK8r/iUygJsbDPqcwRuMxsd
MTmMJbGNVQ+01X6/szyQCivo99rAaxbsbuKVvFShHMegdUQLjAKInJ3fzaCFhCSVtg2bP9CwdCaz
grls8UVd/Bz4RTPc3LiFv4gByhYL3wPXKjvEKb0w2Rna8pIzApCqT9m7/FUTwI6hsGGWtwo/LvfS
yeGgQWaveCbwUU8DkiGyVNXhrrhDg+uKk47YCcZ4cq7MeWVVz5Y8ZzEMx9PTwhGGoSE6k0WMQK33
UaMaLWhL81zAOqsUg39ZBMGEv8US1dIgpK9YdWKIqzgNe3ZfxsMyMoTWcrQh/zL294BmFBfFQaRe
s5Io4h9llqDWr6Hn1hEI6g7ftawKCX5YIzv4i2BfC5nn8lwhMu5w4msyMhNTg1m2F8B0zekdi8xB
T83ILRDSfjssFpTNb+QMXkEeS0zVNyKXKd81T5dNrE30xpcLi9hHpeXPlAgvb+AFqHreai8Nj4KK
lTz36vUnKYyVuAuuwFHzlqMCONbniaI7RFXYTxcjx9YwtCfnw66lLY4KPixchWQe3YFF8FHhwZsL
ZXwb/ztnbezETS6H7s4Az487fVZbN5LhS3mmhtNgbS4hFatrD5K+ERnSJfd+QE28f3PwnL3u63R8
yoHBFXHuIjSa8HMno84WOCqGBsunBbbZFX7vLQ2TV8nhACFoDmfdnxOjLr227jPtC2DHEyL+ygzA
OPONnkFHFp4ypNSCQDXs2JuWZ82hgak/m8TiiZVAStog2TKvkgaaRL0waDIWra3/wW+Jbsvo3O6D
sd1p/9WIIUmH+omUFp7Ud2TWvxbqTugrSYd0AQDsKzOLQyfbU9b9jxhGv3K+pab+V3hebt+OEnIP
zPucHF9orHc2uOTQ757W2LiHK6z1JVWEiin1BN8dqyRQiCEA6PaOSo3EjC4ps20gVDULqvLtu2jC
8QJyzqgmtbNRh758NQze1cO4X3sCddzZsGdoTcLhwQmrPatSdLulUdQEn/lGIuesJc1wrpYkzeCA
hR4YaamqjOOlFu0FHcI0WCs76RXqEejM1oXbQC0dpvfrxFmV+EHjCfYPzuN7Kmx4D8UUNFtood3b
4wVGVbb5usiuMcGbh/mojSJ+7wodgHaU56CSoVgHD6bEjn3B+k0U/NMlnpKdMG3NFkdk/AKw/JUd
03fGughGVu+wLLI8npl9EZHLP7HSCNfTpyCb0AGTmDKEZqpPs2t/UCMjcOAnQF9Y8sOeni94n66J
/JUmyxf57NIaS2CrMtEvjWTRCyI/Iib4v9GvkXAV97R5gGK058MjrIy4BvWb4oiF4t7HtJwqu0QW
E4x9i59Hw/x01jb0T0MXm+gO7QGfFMtcpxpaHdVe3H4G04ngiBl0mUhb8LRFdMM7vCkFyc57ap0r
rls7yqsRcjbq9PCyVYdpL0w7KM1SCqE/mefaaEAcxIbCM7QpdKk5LDMUIyhAyQu7TUEANK7Nv087
E2/V0Ek4zklZA31vCMnzpcoBvZETz7SeYvvGhVp4sIYIE6nM1NF0TrLVcsemNL3EnWAANcTWTtUW
/34qCAgcwK2QQlgxKNIjdQ+Wxy4HJfBZuvfIYjp5YcVgltGUeKZZIEaxK62a/JwLTD8i+JH1won4
JBunJ2FDr2eYz2p584vrpeblnNwOADopneEE82Dfl5dYLKVxWQhHNLmQCyKcPG6ahesh8eVCsAGj
Q0MNCzoX7XaepWWH7BTZeYL/wawA9icHjknxzLzaby+50QiQkP2IS/NFLNdBqD+IRppsclrMKrb1
ZlTAjVcPVS1gNG8diblP+q8b+9227EAUaH3adUVStk7WoEREPIf8s722Yibg282qg0DutU+9tVNU
4nRP4ZTF6vW0FYLmsONwIQJyJ76VAT7izfDUe3OriXWf3CN1aJwIXUTuIjn6flO5IFh/PpYz+GTA
L+xXg6N8SvVWsqdQv5EA5CqA2rnnWJFBio4rqdWFiYl46/JxHGmKua1dzQJa8uu9vLjGHEMkrVYU
HrBhw/wQuzSQ5ajg0aPZ0tqMD0BzwATPCmUuQ4ewv7JmmNgYeHv9iDUxfbDD2UJir+0V/ogQrrgm
LBcLOU1WeTdaq4AogAA/X2n48/5VQ5NW94WBshRHRRXsD1NxzbsUscf1orkTaVnxvqm0vCcnrXxI
tRxlRGszTGGKdwhXTedsgPIKEPsCHIopHkJhllzHjzam6KucFjreafTFdvjwo5cPDMWqzYi+hoNu
1+6/zS+jvK+O5vAZaxY+SO3P+P3xbbRGxa27tgyCjCBqKdp8F9sfY0sBbyEr9wLensOAynLyL49Y
fbwzaXp9rDnYVilnUCM/s2eALueViFbCWEVUgPe7KQgoHOxDrLskD9YaYmLkHsYD82Q5aNecSI7G
o7Mlq9DyorvekQ7pAucszUqEetmNR+SwmzsVnzY/T9NO7ku2HiwRzIfyZUf+lzDL4GEoli0SCjPr
RRpybBsVAnYQRXMyjBaLurXnyd8QtC52yl4dG8i3wfTEWWa/NWYATm1QxD11QvI34w6WE8Sk100Z
mnY/CHPdwVECC41prxsw+1jnGHyNzbe2yGSAOgwbsPMdlaERBa66Qk2dpxwoG4uhUVEFMAyBmtBl
um2mQdcKLw12hX3o44uw69ZIMhUOve01gWjGc9/S7ZGpdq20wRoJAHCCvicwqHjQyatAgDClHONy
GXvHznmcawxlP7QSxDKHOH69Z1Mf/Adr+AVJAx76e8o84Sc6HT/GCViI9O9VZ8sm8qtbmeBN70P9
3ItslEavJDRP2HBypJuXPMp2BwQkTL2zCe6jYKN9SUO60raa6l/l/edVRlAO5B4+0ksHU5iRL2UC
pOwdo0+NnzY5xgyvYeemR0kLipkUoutdpk7glQPHHpRc05Llm9Bzj/y/FPlHraY2L1JVVES/Qn7c
BgvZyp7EsKzmeORSwj1Axct27FMXW/hUTX9+l4bse/bidys7l45guvVSPlVFHTYPpp8BogGMjmmb
c8LtBGJ1O7WB5GIPvk/XyeHJpZUWeh4abIRwO6/63OcwRtydPhzjWX6N6yYFS9lPGAKa+zZfcdQr
71SFpVM+2psM+rJK8ozsVYpGIEYQVXiihksPyYskY/b3Plmk5ciy9i6vwkep07xPi2jdRpQyJajJ
DCzuQn4ej5MtxwyYyG2eM9Mp3MtED3iEN0KSrlxEylCTNhrTUD8cbH6iPlIdoEb+4zvydnKMaMB6
G03iJAVQqjPukh/3JRUz8VS216bjsl7ksVprlSVCVY3BwSycadDm2pKM+G68BfvQljqPiic0Gz/S
mfX4xBiB/Feex/zQBURMIMswHelwUo/Vn02Uu188G8MMQZT0tidogf3qu9EbBY1iy20a6an5VGq6
+SvyvQMv7+W5Wo0cilQT9FZCUIZali33jMEuxvSm6vhtalGIXZs+r1HV9uskcVKjt5gwcI3660+k
CFydaIcpV8qvcGxnycHjHH7vla9mdPuQnSg8u1SqgGDzgybjgPNyLhqrwdJsEIOyKLcdfz7Jo1eI
/ryE0WARYOIhWOFLhj3qBPQCEGKF90ht3Dl0m78ZyuT+k8BpVg53PfXolIf9juslocTQ4sjVhTT5
2l+gUt3Cy8zRqMqLz3WrN3/pC1rqYjQz8rRyE/kW+q/pZoztyRO/ZPTD8VJkhTn2pjraFUumD/P/
5U1+ef/Br41ETi4uLPWmb1yr4pm3l/hIL4nHKT1BCNennnLyYg594Bf91piOyy87VtqwND/7B5v9
LMjszy6d8tSz6NpLHVEq+FOeZp3jqpBtHUdvTlE+pSN6hg2H6F26cWNXimZi3loLo4TjdKczfipO
X8iMpziSm2/g8IRxryu++dD2eY1bVx2zMNXwaoxH4FEljj9fz1GUIZEQavJd1nJ7H41R/a92xh4T
dh1ZmqmT6V0uGa4gWVQnUsMKRyRdlSTGV0hCr42lBBRxAWRzi4PqOrtwSlV9cU4F9mXpNZ5oniVR
7K0CeKmh8lb4sIb2HGhgyTlDsxFM2GvpOWuqF2XLaRAvbasY0qoXemFmOU/ZJYScjGRA+3HlReDU
MnSt5Yh3AgrtWxmoWKrudmfggbkuD48XRX6uQFqhRLi3cmfGV3ahEmmxuaMESW4hjLnvkN3sX+55
UcCJJvuj5KWo4qNRVO+Mo8Ugi5QC41Cc2csN1q3uMj/oDPdvvHA+4Bm1yU179YcYUdZc5VU+K35o
MWsdzHX5gent8nOAr01N9rpnbAzhiWTaSmWEFKRQFj81ob+c+d64NACDxtZ3yYjleFz7eZ15bN/d
g+x9Df4PeEjxFnlLicUNjvwUVfQnYNc1DaSi7WCldnY5EoPQNyaImgIZt0m6mQt5X2q6SsAXk/Vk
aY3cs9aoKhBJex1O0guHiEYEt3QLG12WzIOnYbPmtc4GNNjDbnNOA920+o3jTSN9osMngoXThdt+
MYNvi2nQEmXh4cmiqW0/SoFqB6Ns4p0y8FaYY50ft4utMSy//gAwXkP4HFnGGFCoDRuPAoLZn4nh
8xQykL0r3pK3iUlJ3ar4dhEgzCwW3WVa1A5pfB75YyJJRMwuoWGqXckZ05oeWGbREE9UjnAedFI3
ikhtNkwrRPTr0Rj68Fuy3nhVuyU4DYPEHjsFaS0l3/tADzHWmnZ1GgeP+8euTetwa5Pf8rKkN2w9
cur88DtyyPkM6nWoU0Np0w+KMYyXePwpv2xPra68TUd0khTzyya1UZ7LPW4gl73GwTwQUNfvLhqc
X3/ZKeqLohfkhL6KSp7Wkhb4GyScFP1CnoRWaASIUY6J9BHcnahs/QotHHDMUiI3ZrFwOigbKuL2
GOgslNYAiYVmegWBsyxaBiDi2I7oT6Q2MXzlsMsR8Q/lfJrTEtTVKMlXXCfqNOEf/WuA0dLqj7AL
rqQGHUVVbzDN8z5d5gSAgAhSuqrmg7aFoZmHJdORZ8PIaZX/nSVA5MDzEkwShvMynWh0exqv8xX3
5XAzNNnqF8djOKUgwYgfOBxPUm48biLBW9vKygzVP2Mv0y8Chnh1tziHhjhWU7K98H1vHBCX7ZaN
Af7ufEcU35XKJgm+ZRqGzbkV7vK47ZU75f5H/6Y0QFxGX5kTGeTYi9Otu1T/icJMVJSGJEiOysxJ
OYfaVE1TGdFiKFzH13vWDPNz/aCqQ2Ds/h1EdSZpRkSvgrnyFd2iPXUNoq+iPs7U5gVvkXYn9rO5
/7h+RQ4FqEM9IhXjDczuVKXeqr0mM6cRPUv57R2vBvxFAtCzhYEr4ay2dF66a0KAEkAYkROym32L
WMNEIG9YIDmG+Hn6Yv6KueXhhingXqDgrKt4VGJeZRCjglhTe33uZTSETYzOhX/SsFX0qpGyrGQI
bDqCI7TLLOTOFY0Mayp1KwX8i3PSyXDg1r/nfuw0eIGiq/5LqJ3qfoqSACOT+uALH2c+v2/ZEtus
PjObMEzvBiEesI97TiERJhe+VyEY91JKc36GF1bWY7kT/C2bcTzQcGofe3MKmfJSHtpFLQ2CQv68
6f6W5WUShGgs5temJOAWdEaPLBXV3SA/7gHFqRSQW3BJw9g2yduob/mRD+rUp4xZI0P6LqVHh3Dv
pg/OC61zisMfncXfQn9ZtIvQ9oZmkp3adsUQW0M0FhuMkvwAg7yyqyEyiDhLGfHfJlj5PzjCc+IG
k5PHFxkK3eJfCRbfOU7qrDbNz9OG+M4E31HuLx5HaDuU9OBdgIgs+9UjnZ0Sgux+UlY0cK0+Hfdt
jvLKrgNXdNA56qOzJ2JfWnnZTNs+3CogrR2qpBjen/3H0nTtGG2nCRVQNclxI60sf2zo5n+CZShE
K0HPxmRHT5HiWnBRGR8KqAh/+qeFcr+9f3FHeAZEo9aAvrrtsWSZ/YjMy3NAbcPzaLETSNMBqVgy
TsInijp6eSvoPQtOfdxinVuQ0nmWLQ/Bw1GuPaP6CAFx24bk81Zdocxg2GcYTMfMRQ1htA8TGHfd
WQ/StkxsIfSTbjWflR1wbA8F7UV+g6nLhUejry44BsLnITE6ONeAKb/DzYYcBoLKkkki2ri0Nw6U
geGE/Ga01nvfENdcr+Vo1IicA8a2BUNoqlgkkrhfvi6iswWuTLIc3W94ThUeOY4Zi+BZUxtxpxa2
yo7ymkphNY/sY9Zhwrk3pF914bxBozZOl6d7x7aK7sXcxDSEE+L9V9a0ojWB6ANO4oCdeGYArBeF
sdxZYZZzzN7Kos0Rpv62QdYS6sRu49Knxsm75XjPdhtCW7PBp+MZLYT5/fZa2RDEQFwhCsYL+cyz
Aq0SUTVSDkl8kjtBsKuzLhH6wWzsMpox9ej7BktqrnaOHUxDqV7Q9Q6LFJAqkeNZR5s18adCqIal
7ef+ZiSsUfeS0ihNtkAjwDBb8+Y1tFJtJ0Y0+v2Km98vU1y53/QWJ5UgAt6wU/D7z3ji/zXwhViD
atGP0+jsAnqzX9XSCKu7aqBxkJxlWSfYb2Cf8bIgVCqvYbJtuhn7S3Xb/vWUvLdpKQaH79DG+mbL
RePMfMPmwD5nwHs5+HR19bSP2BljSNk/OV1egIv481w7H89rNFzEaDzh5lhgDuh1dvoKDuYThU+P
Q+mQOKHe/2Hp2RqSImGRj8fhJdClJo5p0YOh/dEfYvt6RI5gu9Qj85D6wjprXXNWHaY0VlPRPVvS
+z+CAj+20BHmcCvnUmLVG6foZvydJT+4/pDREqoNn7uHSYmmZpGpJPQlgJqzf+R48xh2+Fb+k4KT
wrVWRTASH9WqgfSKcl5N9WRcXQ6aJdrkOHOnFTwSJjn82suknddRzltQaC3XnyBc3lixFxTUGmFz
HVVzTHGMmyc/G8B9LyFCvzyYCuht+IC0L1GGVlnjN5uz8Yb8xo+qYBsfu0OPEDdA6o/8QLq7VHMU
lZHZ8jA0hR76vM8SbNlqyWk1FuvOoB9R5LCd4eDjYrWd+VecEpSrFnyIawFdOVpvPACk8EZcVWIy
p4RlOkbMTeTnfDSVjTHnWBQs1rggNwHJL2OfjUYKwn1a86Nta+fw48IS5tSzw4X9Ysc+qCjKJ2n6
Wum8QCWJBT7ggd9Yd99ZHjezrwi4v7XuUySWy7QWddARYLPodGYDb2Id5axQo+Lmq1fRZvTbVqn/
bA7NOVHOcFsfeUgNWVzS0GOJVJfUt2jPMgL1jm/cGuuick1vRJYwQd60jquR1DYzCSA+ct3+6/lu
6v+antJzrJFUA1ON0pHZZtgGMGAVh0/7O6jygsjlcRP4bcxU9/EDpppXCv3bpFgvO2dUwevLIs4C
EXh7mPo2nnSqvWlWeG3rGD0RQAv9v2axYWlHR67CC6FL2gQRFS1HsByePySaYvfUa1+T1c544YJT
YzZD4hgz95FPI0oBWJXzLXhxBLtf/d9uHpViat0VK4EvDwRmK1O6i9r50FdxbSmgQPrCNuCHwUcN
c/9Qd08fovIFdDD/Om0MWNnRKkqM3azDfemTmv2L+mNahCJWGYjZn7X7rtEj8GWVQAaIIuJgtnXN
SV5N/7pGvBbjsPYsZ0rfgWf06MGlAcCOi7NKKXP8QYvex4LsZdnOCBJ22OpYks8nbzn4hP2qsInG
Z9EXcZDfAModnnLrEf6ikn0lFUTj855Sec703j1U6JIXWNHyO1UZxtjo+eeA4vj2Ma69TNOzrrSZ
+xGFGax36XsxRD3pw1MTrfqlMfuN21RMESLVUVgA7fD8PJM6z+IoHXgFFGMpHXIflaJjBAPSO1bH
Tr9R9Em6hP/1+PjfM62nXiBxLFccuRewqVb00j2JQu0wk/DsAUiB2r3ujISBy2pB3XkUHuqRc05t
taFZN0mnzLVwv/9PqqJuz0I1NnGhCuYS54WDJKovtMzVLHI9XHFTrMpNTIQDs9Aq4LDtYgbXkaVt
KTvnbObw10W743cE7VK4ENIl+I1WPFkEjo+G6gFKu2zYJkp4SRyfJUSsA9cQRuZSnFYNqFTUPEQL
OMrhnaIVEDXDO9nD7m30m1AhrRt0hQfxR5N1vdqr83IrGnMdLij61xKWeKp1FgEOuc2AmIQNB01C
A8hsUL/jUGQqOh9ErTlGnfTyQSa1Q3ZrFgiSca1XLl8PCmWW2FVU/6ujifEVRHauKh3oC/NrLKKV
pT4FjdIEWAu/G76uO3nxfSnhPQyScKafO/GrMeryIda2VXO0O6iw7x8/wwd3qhtLMfbAdpCObr3C
raFi+gN9IowngC8j0ZaeN1db/KBgOlRbYfanRvjSu5Y+a+tl0WFyAp3M4JBgTkbkr1Ua7/wssBXo
ZfbM9WbmNrSzCRlgE6dHgYk/ipMDwk5Ja/yGg8UZqf6FqIYS/Mb9WXosk2j41zKUdJBoLycGqAbP
vGcvSkGCMMgnhlTcRBCzpErCFmBqzOAUqM/XBeAqJepW+eM8DXN1oQp0ThXhMK/V/ZVkUNwKXBdQ
STAUC78f/UQYd4iCkmPUHM1yabhmgzZTNdO1jjHMs4mmIdOovf0Wkp4i2ntSPNMC9PwK/fl66Ey1
sJqa84RDMUaVqpz6HCc6OpTLEeg95A4vfr7cqiXxvk3NQq48DDNnqvWwUFaKSRP43cAA/UCPcDpr
n1OZTmS1dGsXtgS0bpKoosKRe9RgZkUhyy/ZL6Kwx6/AI8Ln5JXzqFxaRuwdim9Ma+bypb4VqZoc
d7ibCOQn8b6Fn1lYyAodGjyloOFYEmudgY2XdRHCYU+jdkpo9kXAcH2TObEo482uJJB0ebfUTMS9
kG+5Mql0MX3L9/pl0/BtI8mU+s89py5R1fq+aVt0ir6wGssjpp5mO5TIKayoyuLMW9QVBnEkAdH4
nZ2eLUumTYjKYFbIevs+WNgBB2oWVfs2Ar4rrk6lQ8uJIwnLLyI1OHA9U07vljg9uatLw0agauvz
kKOS3rnLS28FD9S1u9Xiiw7ExjJ2hxHs2KeE8ko1DkHd9/YkGRQkP4lcljvxFBh0OTcBNIvjzwz8
vx05LHZNe1dhUKwWBfZ7auwQqp8AsvHRrqZYBqZ1VNzbkF0CZqu1L9devU+vZG/VgL2cf9qNJLqR
rGkcRda4yX15+yWtHkdNOh5QHd63onbZ4cAP9bT8wK7dL4ELMyEh1SN1rnb9dMYq+znrWETmITKY
6dhUm0153Myjzl0PT0kk8qbwjwJe7INw/fVFetK1AECaZYxy92Xd0f4qs23WgxK0SLkd9P8nwc9w
lPAkXRFI8vU36IhNqEGdnacXOxemwMOU2zIDMQQPdhvhHgUe4Evk1lbZvFhHqrJSSrrOG6kqy4T1
tEKsLPfcNYKke1NjmH7serQqAgftE1aTkdf0GZa29O7FcmqtKGCPWHdGKMP+Xh4m/TZ4JBD+j2NP
E8w+qQFarpsQHJ1yZPPkTB8OCWoc+PryzD8oxByJrGSDr9PblshsLERiNB4VMjLlPl2me2xsnA84
prbAwxJa8dMzpqVA+5i6f5k1buDDOExkEeKp8VmULDYglH43tM7jBaynA5//PUyZYddsUSfgwtk0
PyJapFlO+RISWQBrJYX3Xu5TxLRi9VAzt2NGxXDkroB2afCmoAMeGxtKl8jAINjc+8UqLmcy9Vl3
PZVqkaqKkEpFrAY6YhP3NQthcPux82xlrVTPLHEBG7Rs2TXQlfNnUy4Hx6Kacook8f/UKBILbJow
k5zlAOtNS9RoqTHS69OFgC5kBJJGzQs00jcD5h2IxEiVmoi0bZukhxz3baeTu53TQzlV59gV8Ehy
HBfukhYNHmj9Sbhk++R2e4DFdVYn45ouNmZFH0V/tsrcOZxdIEqjOlKFQFPPEE4Q/0YAQx5DwWwo
O9AA5UFXuuOBhfZw7olSsYEMOrvx5V+9QxgwUwJ+iLHXj70XBUPPNHI9jrN61JLOGoH3Dxepg/XA
ruFxgqdxYAbF7hYXmdzuoVwwd5J7noAti/QmgdoOA83RbLHs3PmdnODvYWviTSN0EUMFDc51Ue3Y
GRgY7H8O7RKGYFdtZVNpyky9N7bX0A/sklNkRDIglkHg/GMmlAO34nr6SHZajrs2Yq6HmY4ANljI
qCW8dnEL73NTRgC+nhYbAUl/Hlk811bfWndvMWzHcoedVaT0vcVPHQ9Abw9zZ5V0i/+6nhgYn7Ij
froD075CyelKaryN57Z08EBlIB+OEEMpCOUyeg9aIBabYCHmcwCJLvwmxa/Ofk51E2TCtmODq0m9
xmg7vXyjs+RS94Red3E+OL7Hq3CjonBKExF6OFGWXfmqpUik+reQlmCZ15EYbUMvNLd2HJ5HY+/t
lA7WBmyxtKXcfVj9p+WBWNBxC6An5MLrycYON2vV11edAl9do8rnYlzTqNqQRvlT3JZiNKsJ22m9
QoHNfcG8dnOquCEF9cQ5N+lnhwryAKJVIbxG8h+tEjwEWCM99s18NBsQu5FDKEdQJt5SUeYdHViv
AN2H9ic2RClPVMv5VBw+rX5ZC56VNbP6j3rpN74mlHowRo4iXN1gxvCNnrMyJqVVWhu39i+fCY7P
/fDEYiNvm0oJ6ByzmXUwc+jAm97wXhS2PKh0G5ONmu1dwixIqTbshfGsQ6RG0V3nwiw2qkFmKdMl
6wjnEjqYLpK+f4flQqedXgDaslC12n7T420zyQPIzjDJCqJ/SfQACSx/PmdmoWHZg3PlNZY60Xs3
0vC4UipLV8i/TidR1njeMkbBWWgWvwIHKtekGwZAKSeL7HL8WGnXCKVmh2McsV8keAfRO/0axcxd
fc6A+neUHPup4nfi2qN2N6hTlfv8xphkskIKCjWCZVuHINagb5ZxgDtw9d3FZelqZBF29yg94LOj
DjreuOUY/As6FlZdty+x2XWPWYHnxZNHpvXtVM5Qc9U1d/o3pXqI71UMSLkJucMUhW5UwfGzmoYx
/lKN1GXXlOOoYMCJzwHINAQYJBf4LiqCcBSlHs9no8AeHNXcliIqCXHDjhv2oPfYooTmrc8CZo0Y
nQ/VWYkfyPGZUHC1VSE0hJ9qn0cFzFPzVqNmTs6/iQlM9ff3/Nit0KGUEh0VHSgMxVDeswhTWh/w
baBnxrqVJwkC1BxFPabMJDhRRh/ZkVgimlrnIP1xW2UP8JKXB5k3xA9X1nl/WpkkwBkoBTW23iJM
z89uCVqri9s+dGNHNnodHECfSoWfbHNh7ZDMtaO+RkQoh19rt6rE9yVWcAYIO/BT+M8LCF/Q1/ff
2HJkSDdEhLReTDj3HMWv8BeyBLK+2p1oZpsmPuiRkPi6SuZoSqQxQfnWsT73TUQQDqWq5LwWX3eK
KXA5B5cq0Qqz/iqUIT6KjNWiEewPjJa3FLBwavIjpaXIQe1K40eia6UMYORt/1QHQh+wGs4RkqfK
BYv3OWaofnHdoh8dCE11KsD4PGQ/0BWvZjB2K7O5bCiZ/9hLm7tUN58vEDeVfmirJJi1QqmXyYVx
awEYonoS9CDzll2/gITCG9shTQ9/HQ8IR1dL4bXG3b/LnH5GI69B5fG6azusHI9AwPMUiU/muzd3
0rAemfyz3HKrU0369q5OYYV5hdxgjb5KVlkSVhs2lwzssSOBxk1cYkCKy4BtBAdecx/mEL0cn0P1
WneYLrCmGaRVgixhVGq7nspxsKmDL0jkHskoHoM7gbvnZIx77ErrE5ZtPR74XfvWVkBLviruTPtM
PcUJga57Xj1WphyJzaECc3bSmYwDq4JcHf4Y++/F4L2/nH9FUvF0m73zoMEI9aVDnicANWiC5zjp
gaYF6xqCzGXg7WUzpho7B1NUypgC38yOLo5a7r3DoGgvV4hiL8x3Utw6z0tak0E8Z2pj+9MdMxch
CYsFEdNnv+pGZ90PKzMAqZqbYtJhAHew1LRxQo9t9PdPjh1X9e3VVnEIHLOuIvxtKlblY7H03GFA
ZfWBLBkXkVUY6nq9Z2h+wlDv4LEETidHFIWJwaNaWgCa/B5WcoFGKmGj+7kJxdZ+iH4Q1zjPY3Fn
8dLxGpZg9xC4WD2Yu1nZF3QzBDAUXRR2+XVOEWnzTmg0AhDPF6h5ZV7m5iiXhkVCpi15kvuVO39g
LMjTYJBnmqvSzXvQyWktM2A89tvoQ6gZ8JFeQWQUU0lEwgXXVo5rHJYb1CQajUytgXAYKpmiZYl9
IB7YFYt9tgstVfVAAKLI/AEAB6wTM1fKdCqAAYAF3fdbvKTeyVD7vU+21I5WTOYL5K9IoLgKfXNK
R16MEpZ5Di0evxYwl7IQOpLkF0RbYrovAk5yuFu0ahUfEqekVjyGb4RV7T5gd5/zQHS200lK7czJ
+XuyKjw+in68UyZhHBetCv/X5JVGXjIMc6Cn5dsAmJsMF9rfJrIMwe2cwIJw92AWM6gIUzhT4OKX
mCOZ/sKMvqZ8tcuiFzBuv0fgynP7sQy9M+ukMPN4HcnmdOynSljC3W+MnTklBbLKJ6sQ18js+ElN
GpJawfOsfBoaXPEHVXNTatPSiMCVHVPJzKGv7O1HLJ7CAe9J/XbKMH+gq0vQwOuUpKpi93qFJuR8
VAnQYU0KmSoaO4G5Ons4u21VfgLcuNGp6hNfSLzNcdnud/MKgVTtO9BauG5ZYC+0HCr7jAJl2KN1
SYONeadP79A0ee3N/5wovwP/Ly9tci4ArhhZA1HEyCaU0QuyxYEQi82+DLRPWI3FWYA6d52RaYZd
yQzMuYdP5DroXV58DymANGuuZVUVAk2ei7oD8LhrsG7F/PxdQPqttI3rO4FEWskmUaMDVvOeGzrx
pvbLv5UdVdGzF8FfcOjDqH+9xs6PGNTE/4ZXxi9efNbxDet5MQjR2QU849f0v+EzhQLydUfQZrtE
x1WgkY8X+codX6AIm8rLNjQAXMZU/+Pv5w7GFh0+WprViS2nBQOLz/Wq/53R1dO+1JQ1Xl650hF3
1rmS5cceOlfLN55MAIJrD6qWj7S/7AnPLPvSbgbJDYVmdxlsi95I0TjieZ73WFiNwjczM654xEua
hQZG9Kfsu0+cUJ3d4Pa5R40EgbXz3dpByEwSzctnTEYvwuHXzNFIDES+OXhNjo1gcLm4JTBM6Mw4
WyaouaeHMPm88eeTzoXOQPoj/w7OZ1bDsO03XwAGNCnoTdPcsOvrZjj03u7qmCk7qXwh3j3ia8I1
+8Ru7w0ailS5bTqSwAAMVgUIHSPkU9XMsnumqUoujpOMhW8NFmKTu1mTQBqPZbJMaq7bn2+mIpbc
40vfLqSZlEqWcg9AocSYjYUmiTJUTvwMr3Wm5MiBNFKf5J3e+XXMF4yjrn2w+FgAUpekFlFsmDvC
/IFxCbpO5DuaUQpHzT4ziMDma6PpEbZmCYS2A3KRFXqe/zW6vqG0nFX89gfT8vpTEvb+hwZZoG8+
IJm9YhQo2tXcokE9jLPJMggOZw+dyf+PRxFVdi078ADSwzdBm3SriQNJ3iiJX/qMWYsyvyrOWqKV
DzhkH3vlKQlNJgeZ4hLLUhF9bi7VBgSAXaj2nq8d/779n93pMSoFlD51o4sXGC0xbDEB6bdNsmjE
tsQteMEQgrAr0Nal4Hu6skbmhYQBJK14nTSQJy5wAhIg2y3GlxbK0bsZbDjlonB+PpTsZargaZJy
QWnRHRHeBL0NIJbus1pdn3i+Sa+9IZJBjlYPIkGyHzD1nXCQCtW1t7Z7k3PXOg7NHn1LSelz5gYa
FgfRXwEthJwcgkVrQSOB/U4S7rTrVUV7o2rnFZpaJxcJ8RWdQDmCAAyquiyhZRALhSyvmCdw2qHE
wZbbGN78VQR2oeEuH7PeFwe2bFnzxMLKDCqnZfy6WqduAbm+oIfd8gBcp1eOftKM5v7e/PVfl6iw
EArKC2kb8mayJZy/f4Savu+nAB6etCNkPasu0f/Gt0vDs7m0BOABMrUf9EHQUhU/HhFJWwcdmtMt
YYU1hDOU5Q82cD3zTAGOji8CrGPKFvW7AAb7XBWCqJ1hULrSxYscUnP6E7OOsaPS+qERwWwV9W76
VlX9q146HU5vcWxW3VbDXOIHLXXrLh6d5IHZIme4rscKaRsUsppYs6Mnm7t/XYzppV0jeNfY5RFh
ZbhZRTvaA5uBBLZVJYbDrBquc2HCiNVg7s4+sQEUadzSsh98ZlSpLdyRwv064f+mu4fy/D2SPFna
RU9kdPMtmluk/axRJYF5DfhvJ6XBl647koHt3prLvkVVj2MOxm/W12M5RSDkQHb9AipO6x0TMeti
7+Ob6xbdQM7YFuAwYt9CsitjCRKpQrfElo09CKPVmE6iiIsJdBpn/GIMFFqrjhDrela6oVHzcZCc
OfQePWCRpEA3NrJKGXMSbT68XHdjCs7cb0fv/pg/papgUx3VK2P1q3+2LNM5pS+qlkc9DdjsWyUX
Va0Yt+NnxQwMpP52gtuOsrE6Oc/M5USRwgicCqZLVQ8LwfNH2zEQUo6w4YDu0hSM7TnVxhgezlaN
+PbbAkkQkcwlv+aFtGs1NDxweJE8xR3HKRyKBIDaVDe32ecFRSCoaZuVSyM3MPsLw77hPh49kvTt
wF7eHGrGjHj+HegWpmQqL9M6sacNfl+SKNxLJuewVvFJwjJFqh1xMz8QLo58L/v81tK+xP3ybm1+
Tufesk9tK/erl8Y3ppy5XuuSoNXn0bXzhooHu2AytHGn8Qv5NGqsEomkBuaxasHsb7KCTUjbUaVu
EpMDTQfr0bAwNSDifU5Us7nmxHVDUmYNnMMjFBbWgJ+4mofowS801t3jJX68nPZb5CofyDYnAqyG
tBiUeA80kewVNFadcTHrUMrGvCynxebMtXMZeelq2pZYgUJTNqBTeN08QYjZujukqHeZy6x2igko
KBr4+V7t3swYP9MainuuTS9NNdLO34h4LfQgtEZGdbcUUo2vW5Q8a03pnpzMr5kULFm1AJ/pllTt
lJya+LBGNI5/i2JlqSGsoFZ+pq9SlmsN5IfroQ3Jvf9wZ9Cp/ixEX/DYX8Q9CCWB/xtD6IosQnPQ
AsveLl+oZD0tm5pM4VI5IAFa8UEw/qtSvlJv3TO94WpWeZPVYRp9CzVIQwV8Mk4V4bDjFzGeXiFe
KmDNBzgoCUdXXFYooLImtWfJ1JT/G99QQGlkchRp2bfbGu2Vr7/U65Gk7HGmXVA9JKWWTNIEODXb
UmWd/0p1TCKPMfeoDWLCZvnV67fi4CfeOwPL6XzeFvjC/fyAhvTz4y1Nr59FPKSM7iZBmGix2hN3
fige27nIi/7jGKeUBuodTv4N5KUHw6Tt91Inn7966hw0ymLpL/2Ms83vf0U++cTGI4JpdrkI97to
j0yOFlikB19BP0xWu1tDCHQNTc6G5koK+I0IjB3kqTnI47VbVBatoG9A8mC6kY6X7TTl/xrVOBVO
aRXo8M5KgYpgbvsWtxtycusS378fcANmKmoPf2t/rLssZQqgDLJoGSF64KWW7Q7H9FgM4EfCMTFk
SDjZRky87/Ru4qFcXUpb6Mgg9l5OCAl9ehnpUdK2xf/f1LXbIHDpyWA+jxr28D176fhxsLOtrK8F
VwoVTeE0fBdqxHolRXtXPi48H/dQYt3UFMo2B4poeO03WBBQg6D09HytfxHoL1UnfnpfMqFBKokT
oRBESP1Xt8bQ5M268Nbmm+ttmXYjX20P7kULSS3uk35XLTTQtSuxUnw3UlxkAX8VH6wdy0o1d5tq
yjUJaTnu1Vc6h7w5gaRVM7JnIbumyZ8MPiRaOFmOXb19EHrJU6VgHDJvybRDLSL8GUSbsePvij/C
Vg219b5tsHlOxql0fhHj0qp4ssIvOhf9ghPvTNdwt+sEt4cGBBpgKQaVWlbPoywVP7tnNakl3e2m
OEqhqUKbCQobjQ6qR5WuANQpo6xKUPzamTD3LDjcNXwe28qhCVwzEJgUQwd+hsRA7gZL/bA/TqtW
gUu9uukGr13/NSL3VYmZL9NKOyrcDlb5OUITH2jmKvcRh5emAtjDGnSZGXK2t5SsZUVMm8eQQ0LR
l2lfLPyAvhwjU6bKXqiklxUxvE8I9VQF75OZMAQLhrG+5wf8PRJXZcrDuVXXFMRuh0xB299l90J0
HIOUAsaA9pZ7fvbj2D6TIg2xMov+h5TtkaJc0wkbXBsieoUel/ztWD7HTKdDSXTf9B0VZvLofWrW
S0scGARbitGe0jFSUJNgjIXFzbuakR1lJ0wak8NvkJPtLjDXlX7X0u6v/fblIuF0ZwkEtSlndfSp
42FcpSjRwMPlmyX42z26XD0ZPq6VFc3sctuRMe+/e3j4WdFqdRVPiEFo271QqyhstqRXfP3dOMM/
1OPcThyMcftUC8V2x5McqRR8jw22Z0iLeqAKdxHY2VLLnsMeOSvrJfMQqBsPs2Xmgvp8g18vTyfU
YgLiy5YB8uFaGT5dbVgctRC5bZ5W3pLv7asjWYyIuuNnnLOLk/F41xZQjlOoKyJLo56FFyWnl3Vd
tK835Kvdy5ZGnplYkj8Eb5mMX0zaRZTsjiT7BkeiDHxb5qfMvK1czABAce+yaA/4chyxKndf5hIg
AWhVil5VHySX3u2DzyTjp0x99tW1VF28uTU5sX/pExM96/xxidXW4Rlm+jhF2Cs06/W6OhH1xw/z
jx0TIu+I92krJGc0G2aM2Nn2FGgfSDRRsM8gp5PnhO2U5fRlxphoQKTKZ8h44xdhMESwT7lLsZ9R
AAkFJcLWYgIwTAOSykpbZRJ3MY7/5C6vm9aoo733AfAIYtScnO1YfnhK6hjvEdMaUH4=
`protect end_protected
