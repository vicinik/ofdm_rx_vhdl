-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zvKrcXdVThwHdDhTa9EQnhpEyUJ7gEwq9sWczYOUmq3XGEJN5KPb6fKsO7oemmtvHhNoXN4sTTG9
SAZmbOnEm8xy5TXpVbSPdfjHH9rL9UUqiU2MgQ5IqD76d2xoBEpRxnka/FZvGAvD+W8aFnxCaKpj
nj6CfGyUw9IcJcr1UdPBgy0jAvd1RSooV1sZ/00ygLWckfk/XJSoSnX2hQ4JV4X2V5+paLuoEs93
VpgfYxSldgUefv55huUneHKMZzxrQs8ZFBFc5hfao+odIpyViuHPO1evw0UxQVZAAyAChbMdYVDd
7w53MlPXJKdVd52t44RLBZiySgRghhj6CzHT/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
DxGuuPMEF1WN0/j4AtoxkCVdELeoJe2PGLTZsv72ofnGqYMj6fZUjamlZ1BUwYdfxDMLoGPzMpDP
oGPA72mRBfiHnnFFiHE2pMyUiOehihqclqTzQlR6hRq/r+YaN7SXmp8znAJJbGW14JgVEvJVS8Sy
N42Ei+z7DXSOQcOVjAfaaA+OoKEiUmkHBiz0u607hqA9izBZgGWvZ7UhoRKgciUhPN6Ryz/TcOpu
VKLrmR71eVSOA/JWxYuZNFXB6e5J46XBt8gEA/c6q3HdEly2TralgzOUALynAWldjvFNQeGClggE
yvNUH0vv6bnVfRb+HTXJVl1BIG2nEKji2Z8UevdZrv10l/V3nkXPPT4xHruidcvMDTFg8gf+gXju
ppXTu7MYqt3J0HNdvoKepzjothg+24x2kNDal06dB3rK9uXy3N3Zwa1cBWfvV9aUSUhdBW3rzzBz
IH484x+RN2RBr/uyQ8NENbiSxUz2UQn9rS8Wywh/MyGGaRXtSpHlOWhj7aLpNsCKlTssgCA3Fc2O
uxHNubcDNvZC9JKmf97XTTaJnxEBaLg8p0PViQVtDSaa8H+lBzeVsxb3McifQlKHO56Av1hDSqkg
XBHcOaZHxXnzpuJx68dvp1z7ydUD/OyPU6ZY50ScJXi+/8UpYaFMbagyBBHegR9GjE30CIMth7xd
2Xg0EmSLn3Q1Z8F1pJ8DoCXxKlPCVq4dTcMwlMCdQEenYj+16Af1M4GfEGStqUkb0ZOpi65ZtudT
hh4aYgpjluEaHRUoPm5KTkKaTW/DMuzvT1VCnlNJO92/nHM2495YRvl+qExzCodf1bxUrm/cNh8H
0eNRslJFx+kUOkr8MKFFj17PZ7MIP99Fjs466le9rF+SHw0VFzkikZWhyKQhLaJWYVnIr2BciwSi
V1hI31exGUuhg1TPprk/3WPsTV7uElUdEOGz1FgjqEpb/V3fR/GyFu+6YFwe+Q04SDNtRobpkXh9
mnWMxeBa1VGOe+Nmins3/wsnHknTXGV5hOynJwkQo+T2hNqWitCaZ+2OC4amZy0F/o/paBEq3esS
rRvMK8Uc0Uu9FTJXPMTY9xfa7KT+eCcyb/vKO7Eji2eWfo/1/4gWsbyZ3p5p9UalT8EinquDT4I+
4Qg+9TsPKadbNVf7x8VGGKrJYyNExMKvMc6w11vSLiO41xRGBjwWeZowpvYPczqlJoFzQVYTbB0j
EkPOO+bWo1frTRIUfnNosXZLyu3Fb219IuISMYchbgBPZkDDC3idBClu1irwGMGmp1Ez6+O0Z+h+
D4RUOhwQjh2syieZTHjRtrQ0lp46+F89pDuYrf04//lN/ZP6zPggl3B2aOIfBzJ4ghxxdLRAvwH4
hzoY4F776xXDGc9eXo5ogDZEtZqtflNrtkgMPUTu3OMuafcVB5JvWEk0tTrp6/3dXVynYL3RHH+5
B0QM40kJ0UGZPpZY/TTDGVWXTG52cDssaa4o31i248ngaK04MtQk8BieVDVx/57+WWXDc3q+NXCg
YlY/U88RIftiuPdqolwBN4OcDeo/fy13cW2wXOjIxFwDx9qQFSIyQJxP9eJyQE3RuTni/n7tLI9R
MPvDuJoIhflzwMbmTncTMro3qTgGtcsQczy7aKzQsr61abODHhrHTG1EVAEFhMOKDFX0fdI3RMqL
EJhYwUTGEfqLrZwSOnfjxayk0mo7w5Z7BO4NU8HSgoB1K0AM337pejJJBBNYVBOtJg3zog6gTAh3
YgF2Bmp+2dKrJFn2JImN+LTVVr8MfcCDpQTkviyW7TvgKj7HegQqf9rCNQfDCjWBSsUv9FemeaOD
f7tqH49obJkMPsJbDbXWsIxJVLa6WJ/gVDiBs/zEjgsBuZi8HgupMCvQemN9kF8d2MGCvTDUJtxQ
i42L5T49vnaudKIBCl/7WqE4PlWby648DHsrFo89Lhp95AvwmekFUp2kpwqgZyI2kLQS0bczQFpr
EKkoDKbSaVn4+xB0bCsiOiLX7wAhwioE+L5NE1szzXOf0EGxOVfBeLYCx/21UepdNBj585/lgmZX
dEx/G1HQGUjhBdycRqEMewHPnQhVZI74UpMDC564HYQVOBcKBkccqHiAn19PrrqQy7B9otjv54ym
/OAg4kUm95Q+qOO+1zZ/+zt8sKUTgqLcyrjM0SjyE2lit1ycjYesKq2ykAgCsS6GUYhXNq6EjNoY
tNvuyESv6LH+IlmFWSV966z85WGhLAh/Xwopc9str324zdF/xIFpm7cyA1Lsvn4aomQ1hIQYiWqk
VSOr3zjfG9ITDiUki02fsBcpg/iZtTQkuQwmb17gHI4bYvLqzN7GjBHJge54eGGIZesBZ8N5jfHI
A+K3JZT8R7SQCw3Qury805+G3/BdKyKNRgy67Olny1PpncPfM2yWQaZTjL/qtN3vAMeTfskZq22O
RHFioGy2q5LvzsCLHAq4C5LHpx+qKLw+XY/zqbSKEsM1dJ0GG+euE0rCnKPr+cuPrqXrWp5wDreM
/jTzrHJb+34q8vVU02jetiK7aKP3LaYqU0+DJBUWN5iUMxWyHEgBzu/EKdTdnaYDeOZZ2p8lvSJ3
zxrIGoY9c71M2NcWpXx/wyTgOTod8XQew1mrl1yl/qNR7Pi6hpiZfJTAhvNORc0Uffrq3LoYxTlX
BrpAR+21yIZVxohTy0k0/xyr8j1aGFjiBiqDirEopXDZbTBc6krW7AemreS5i/N7kpw6SBU3ivoL
MSDZC7A4NNSRHV5abX2LDVUIiMC6n+li+JsTh48RBeGKWz6+4eSRyRm1yVo6n00/P/FWOKSlgBRy
nMcBGCJrqUA/ttsAWERQYZVZmRQI3CRrvppXXwrszNq5wDQo3VzC383Kb3cN6dYGKLn3Se3dH+QE
+IOxoRVnU1AmDWK7c1lRdPYY2mNu587N6usUUMKC+gI4AiJCGxVOkLcQtf5LaskfUmCaU6JLnFFz
hi9VOdCWNyuLrtus3+ZikV6ooHkIJUO+Nh0FG5Cl+nkyCAxlUctmbO0T6pvkfwyVEdrtSMoOMFMY
2jFD0u/7NDw8Rw9gS4M3pNQjAM1zLJA3D5iplUp/DqVOhlIVQaiMuZZZmbPrHSLi05Gki3jd3Ds4
h7HYiqNUwDuG0YafIlFyoXAwjbltWH5k25G3OX/KhuhF1xLzEn7X8QNsBthKSD6XfX4MSSDO+sEq
oIrFY0BT/0RfR82JkpGf2uJEAtTyjvYvs3XfLcAyY58YLfZ+QjL0OfPhd/kU1DwkCjKm5MzDqC4U
UlPPABZhATZEE6z0sOjvBp8cqSWLQ3lWfrMotAhmBxnWhkAoCodrJLYQFb9067uo4kfxuX38Fj7X
hs9u4gykwZhcD8N9zZCaLHtrfjIcAg/kBRzHvMrfjDDw1xEQ4//fqdlSNIuPtGvCG2Sa4TiXwFCu
3YsEu6p3H+jsaHE0ze/n9757+y0dQFcI8h59uiS4C32sJLFEimD4diXnWqmG8ZOxnp94DeXRrNFH
P6SUQPvglZrQOYwz7Z17IGQDy7izs1hnDMnkSY3+TMkLU2/8Bs81QOhyJCmwzTCRXU4SMIplObWK
nBDY1gzt+7H9ZDSKnxpfV1lEaJp4Nz2oOZmMkPgMlmEG2Ws3PtPUuWBZpp4YGWKg5wlzBDwSMYqr
4MZBsPnMb734d3Mk//2VRP9x2D5msjeewhdplS0tRpylMQQ8sL4Z0G68+fhuKynwI7IhggMmS2u5
eUr1037Vx+T7yCoO6PP1OxHkSaxv1BPBKqYBmwG7qDGe3HWmij6Jj5vSbTmoZHhHHrvwY0xuB/dk
3ICdK3K5g16240u05K309r11z6/ezyApuKQXUwofJ4RAG0lC9PANBEzBGKXDcSXKNUA1bfbuGKi6
T2oSRbw7DrXKX/KCuWVOC1s+YFnS8RpvEY+VSuB/bFnvU5fFnFayV9mwRN3wVwSi04EdZYbaNb/N
H5mM95gpL3pAsDwvI1WZ8/fKiXCjpsL7FbWMpEXbCA75dCbze73ikhQ7EAupAhF//ue5GLiYVFZJ
wTZtFyMf2/1QBkcNuyYi6qenb9OhJMM56soSqsAnHB8J8/kuvr2GiuyrvOFckcfw54HBRRpnWUoa
xexQp2yn0EJ6OH3FBEMH4I0TDiE+Bej7MTetSUVyMlek8mfCCX9vNK24GOTyZyKc5ypQU3zGN9Dd
YrToCZCzhBDk5+lobKMnbp89n0fu2/ROncoVckwqdYpF4yy4NFnHKEFEnOfUz3junOE3NRu/tGbi
smKv2lWATWA4tKUeKptJOxQTvb4L31WPuesRDc/2Z0a2FnQPnwxIf+yQu2RNsjdaGCbnAGQs5Uwf
KTQnI2q85xq5aFe0JGTFyxj9ph0KUUbXPxwSLQ/vviKql1dLgPZyAb5/xUoz7dlIryIjRGr6EsF5
GIb5IyrzwhCXie1M1mAy81e9GXG6ouQTwC/cccXv6J6Q8XRo2BLslmcCCpwlgf8dgpzkbvUWm2GD
0oheJ26eDzXX7HTjzBFUzcRRwoLBfgj8ree/GjtFVkQDvY3mVWVGyzN7P1iCCRxWy5R2DTsXiyIw
lPQ/jpaDeWKSj3LJ6aFyorpBwlDi6KLlR/DUE+MKLHITRjFG/43w/XRb3yau/G1ka2bD0Br+y78t
TEal8MuCZNSnBbkXoEh5Px4WRZVR6qSYk2qzFMlHK412YfSGtDWqK8wftGV574/2ee5StUdR+Zy8
hu2CiBu+G2NfE52Z19EAEJ3jHaGEyBBl6R1z9vp1ix3wqQHxpjsBWm6IrMX55lWdUEaWl/C3Hw9F
JhGFZuJhR8BJ2UVgaNvFavFvdyqjiaMh/Qd2XL27LLCCkqBSVuwpspxVNV9gpzJ/ZC+x6hXkhJAG
E56C3DDHOFzsmfYEuwXFstE9j/SnF/MirXdAMF2vXA3r/JRNJezrIx4t8bmXWKsjG76W7trDbrTh
+clkA4IwIr3uIMnYhQsxZAFARIBFxOdvwVjob//rQEirSxq/zp/LCwXmEt+zUIGG2rU/ba0avbaN
aWZhhYl8XIEi6eMfHm3foTH4c3f4ajf3EP3CbCh4XGHadMcd4bOdEJRi+aBF5Fa5b/UixOcS1A3m
R8B5s4gpaxDq+0nGry3dzmLXGrLbiRYANq6NjkzIDlJOuTl4mhphadWQoqfFNywGZ+H6C+VkO3Ow
ZWa/Jheed/xpR3Fp2QvUEhCiEy6S7Q/uSBH4/iW01mZzkkydPgl1yRdiuPFxJ1c6X+dwGvhcOZA/
eZuhZDGtLESX7KLRypmvcurrJ/LPiNREHElRbRSbtbdSVcDqFb4R5LnVT5/kA/QIe38R1rD9fj5d
zBOgX0AgOsDolyZKVOCBCAAwfjGfu8wKwRoI3VmbiLAIVFU18Vf79N1s0y8ceL6UEt4oxjxGgjLg
pSxc9NizosbD0lcJ5c91Liv6ihQjO5y9lzeYtexzv+mZWJkPKZD6vhQXcje07ClBywQ1w1QSnrPC
8x9RRxzZcST+fh7Mp0sJ+5RxQtqbZofduEQPg267ZidLpeOFLhZflfVPaLrQCI8LbLrHppYmqKwX
5LXXnreGNnEJcvCDvlg3l668qe5xngHtv5E9nCW7L6ihTzG1UUiC6G4e3FjvYMaWNa3b0xeXJ5Dt
oJs+lkBE7ho4EWHL/89s/oN1ObTb3+jT1gpXXid9nKIr9tPurgIbpdMLVC0qVWzPFxw5oPGacJwZ
5z/LsKFvLMf8ko9NSA==
`protect end_protected
