-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
inC37VDS3GYp1HJ2k/8s/IO82SCLF3rJ5dRsB3hnyZ+tkSF05DVp1nVdatExTSH7jg6PKNay3ENH
Vg7yOvE2cmMtU5nSOCwmBQm8qcq21pI7nu4D0ZFMLbR/H/tLF9M3f0sHVmYqUqaWPr/L2o8NW5+G
pjVzuiCwii8lDW8r7e3dBQatL6KG+VaQdWyHrA3i0xkOjKEmEXQI+HHoYaLApQrfFiVEbET64RMe
QWYzh70JaCBvKGu3WTyieVjvrPnpY45keMsq6zvZ0oVP0fu6rvbJAgOeLNd/90VfEZJ9ZvX08Whw
1Ge0/BhUz1tGKvT+FUpVNCJfLZrwRdNMVpQcrQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26880)
`protect data_block
Rb0azX+QYOzuudjyLuFYkRy6roEA+fouAOWmAE7N9ea2pnOEpYeTA0k6kKEVk5rOsOrpkNZARSuc
4OpsHsCLBG2yQeqXmSpegchCn0NRKF+uFLnMlY+nKtskvFGNVwvWDL/OWN//eYhXvcJZpuQPS+c3
d2g2qrVTZPcMNuP++hn4aseoUjjn78TEhsjHNsJTPimmD+N7FhD93bdZtKgCcg/n+/89LQkjMMB3
k7SRzFotILWtk8HAneMAaMiRceJpjv6fDPYEge4nRGG+7NhC8X19knYR8hm7vMLrtgwFCK3dZEAa
bOYz05nLU6PSKbey60EdZ3o58d13z6yNMMDkprWjGawjAhyrgmT2myRe8tkbrB/tG9+AWwSvbjle
lhiNC7MXXxvDUPR1gO6DgCDiwUQENORnz8qutcmPKbYVee5PK/2ugqZ0MWD5+a2mMvloUP1A6PUZ
px/DPOjx66Dc1JNok+8oyDC5kD68JBHMFKPUMvck6rWC55e38u2RG8IbyH8kj6HD3l2FhikCYQIO
ZI17i+CT8SPlxZXAtsFeS5RcpF90xxYWc+FcIapxgewbRAbolGIWqgHoxGkHW/+bN9L1dzUd9QYb
kxvLB3ySFfXoyXxVVMMETXAqISXnzBTUQjRsFA+Ejfyq79GcPxrMpvGQJaSaXsikFyp4BWwfah4M
JtWv/Wz3qbUGuM6WMfGM//odqo8SEXxasW+hf0t/45vwDIhcuSdEZLgVIHFEzJo6sx4xA978iH4l
SZtvWxsQGxFs35DxpDZT7lpUPB5eoB4w1HzUDx4ClKUucAnUR5CYYpgicrCXPKnDlBojekCl1+2t
tBBC3/JbN9XBRV4xofVdNUfcITiz52yjJkc4PO8AX/IeGAvQ4ae4YO4N4yo7tdHvCIetw9ZpWx5l
4GiXX4OheE+6SwamEeBivXAzUFM2kMfvhXm6hSWG/zCRPQ5Plfn8lH8VRbGVXoi0hBLC+wTCf045
+tWKovkL7k4Rmjwu7jKAkgUWSRDhJl1wa6WuDw1grHzXMR8kt0dWX6rvHdHC7RryD/Uk2ffSzXRX
3I/V6Q/iOmttNUZEHUkFRx1BjTdfoeL+SR0XepIN6oj34ZK5bk4P/BFelT2SQxTdTElQTzOaIby3
HTw6DJprqY9hFf8eUMm1OvzCzmjaChKS+TBeUSEe3qLU448Ale/UK2vGYd7OeHgmSvqiWxe964iK
50YoMqBJkp+zKoMOdDorXpuq88rIyll3s2jukpqkbCAh+1EHQwn8n1ncUvAwhNxaKGOYOA0qvjd7
x6q2mLg3LZ9tN/+8c7vcVbeY11HcDfSbYyc7jM1j9suPmQ4xuXTrwCV8eaUEei9bsxUez12Cs/fu
bi9tCyZ/k4kbZnym1ylR8Z7H/xcxu1wo3jrYbYdTehdJq3iTHIyhYG05v96vEymgTWdAAO6oMbzl
0mf62PpTshsroYwlJ/u51Ga5vPywROlGOltGNeXyHbmm74puJ3NvkPWzdXm+sL/Q+ehZjy91J6+b
sCloY5v0CtomE3lebQFR33m40EmyXq1QUoO4M954myGE5I5x0Kxsw5oE5eUmtOYBMNHlp/PBZ/s+
jW4TYNQklhLidOfSiiD8dvaQGVCo1+gYtzrHffPhZ/6ApyAwDbRxedjBScKX4T1rnZjbQh8WXpX0
EiQ4ASfh1ClABTuY6sga8BsLRVbEuBgU/TwUSp6M4i5kG1+PlYH0zXJ18zzyFUBCySar7CtjCk8K
a1/IeCxkERM9fByCPiLya+JM9hx4uE3aNrS4jIWEnGjQ7HBJqbm3B26YQnEjH/LD//uH02koCRQk
JuqbTvynE/RfOWeYhbs7K6ThgnZ0ILB7AZIT4WtRBmOYJLRX0Lg1Gx0k4p8dSCkDcJEsDXmVuOui
WO5YIa/xy4y3q6ampjjLnL3xLTAwDWlY3RdY0klG0FWEgr662AmQ5zWjBAKukJ0BkIIMuHchXaDv
37+6f8ovdmsxiyIoDspyOB4CEf9W8mvmhhHcycqpECdncnAIPrjSjwg+2O5ZDbwZLIrOHir5IU4R
JOMpwJYf3f3Or8hJjCWsuE8BgigN13Unej2lGIAJhbDgWYlKC1bW6JHI+iIfwzt5nrrqrKvGJf7v
z/2yvgtUa6ctPtMRkRFtkeyDDGEamYQ4QHpKLaf034jRrpoZ7Gxa5i246bgeYotvTAaNaJmxAdaT
S0gtPzegBdXd/6YdzhQXKgCVRJpgKLyD8zUKgYvv4i7XUNeqtcVb2+OCtFSXrj9y8AnOoFCIyw5N
DSDFnW8i8SUaz+0oFqjKXSv1UJgIp9lJMuP1Ce5ApqshiyYNiHW1vw72jLQ29P3H+CzCgxnNDall
/WF0AkAIa65KH7gie0FnwdFcxLq66wUQpim5vdQaYI6G4raMsA0WfkZYkxmG8ZrKf/KabiGf3mk4
WSXb2ia3iAQeJFpSu+4rbm99G2EzkgPWW+CQNCCRciadR96K546GHMyShb9M95ai3jdmONhzO7bL
3vDpjBxEuMsOSt/xhtKUaCI/gs0G94Yr+AcFOHT09ZYZ+/yPgEYOqp95ZS3GU8ym/iwo73+HMBAE
a0ff+gRBIFhQGHJJqY1Uk7DYrOJ/nzk+DdwkAuVHchySWPoYDF4+5ge+psPYPYspc0ewTt/QX93W
uGztXnwTIVgxb5bzENkllNR5jv6qH87jVodKzxeQsELNH0goFlV1fR584C97imefP0Ub8at5ewEY
Wqu5yQlJCLtCz3mc085xzoSNKRNcAB0nA2R8ESbOfMZSY0KMv39bBqtRfewiIVwgF6by8WoyKW0c
AhH51i3ghTg8V9xkOqnH+gev86s0GQEwNiRuHVCHUcgebY6yJVnpaoR2aYbI3xmLbv/lROkrRHpk
rva/ogg/ItYOeMP3SmK1U0XsbP63FyMbjNmUdfbQpfKfCDYe0BxZ0ArVeeP8VUQdPQDcDONGJs7g
KgbXMrJF6dfxaTg/gBGTY/bzJd2Jo5b9wiZ5vbSkRQjZ9bn1p4x8mm0gG2zf32HUvvwVkqKPLp3I
LDkBAGYuPrj8N+Oy6xwdrmZ57OwCeT5PCwNDmeJbVz5nD92+c1ny/hL4QfG8QP/8K6hZHIySaPKM
mZLDPFugnlK+REU/YW+VD7LdNL8ti6GmOMagtvTMjtjt7J57AgSxvzukTirPmKdEg7vqy28GzCsv
bsHns+TB/nOM5JOVOR3PR12hNzhiMaOqe3Zr8KL4TRuB309aMlAe0l9G83MEs5IS/zWUu9IWtSRo
eB220q6i1SCUoHA+sU5UBS4NW0e+PCwK0yVdU7NeK70nvfNnXZC6k28m3iBA/sqwQYoQ0zwdQQh2
YR+08MB+/7hKjJ5U+52Q76xEJNNSGjkl6JeHAHCaBbI1ZVYIdkd2TxXNEOdEQT9AFRKcA9I+k9F1
fLovM8e8poXwP4lXcD4IXkNimMRubOyGhm/S8jXvX9nRG1KD5w0eaF/GWUT8uSxQMytbWPehsEmX
/YzhtWd2UXzmU/x6dYsWPmMZETua1fpkl8fke+sfn4zXLaBXf2Ugr7vCHHERaIVdHJw2GwCdgw8+
TCFsyp/2YF3GdMCN8LPDUC7IWGZmTbYgtB4uyoJ2v5ykDijcA//rUMK71bHh2NhLUqy4nzR6IDy+
qYFxcV2ezlArIrupnkA5eGxKiBiXIbcA1QLMQihm7hxTuBAGAj6vAlRy3nk7fYZJE55gc8UzuZsn
pGXmlzzggbKnJ8yT0VLL0U253IlNez2dwD2wudoeZEVVCNFp/8S5PDcufe3dFrAMHnrCly0zOrfW
+7ezigNqMfmxzj5XGJzQXZdgTJZey15TRIE0Wv2W3QqVapT106Bno0uoBMt9zLQp5NQm5/uayfqA
Euu9r1YGdxdjNyFIfl8qQz9hMY/jf+qIh3DDCrCI5lnIkcQu64LA+6/buhVvKt8bhlNMjZN/n9Pc
rwlSg73TFQC/DV8eJMAc9axt7MTtoDx0yeRYLdBHB1LNstHJh8tFlwYIgDWv8FsUL8DhNyZxz1lU
j9//HQwNqnM+8BXAssdme5Dy9ZjaKhDZfwuOmrYSHdwjbWh+7kEMVE/WJo6jz0/dmBsUu1DZ4Wms
4SyG3mahSpwD1EpUaLUbZP2GpwpqbCPnDU2LW2JuxL5rGq7r7fBuzoNxxgKajGEmWaRMxfjdLv+y
XRX6UWcKYO+ggdFRl1gCozKZsVChtVrQAEo4mwBZIgR3dqY9aGCaSGDbVLYQS/JjvFy64EDLAS4u
lOm4BUrA9J6nLP2eG3U6GDKTAK2ON75PV/DS6VvbzAOwi0wghaOY6AwRES2nVhSxOQYVZ99jwvCY
5LaiqApa1TS+v/auG731F23yaLoBx44LcfyYZB5SOrd8gvekBvxfYK1Kw26LUukhfXcoWCratp+7
W0RCkXdcJZYlZ9sdjXW8S5EsEyTFhSZTTNyet0+tYjbk1F8nFw+gB8zYMw2UNzTZ7hYbGWozAr/I
U3vVQo+sfFx1oQKpHP+zd4HygVpilnJ72QZpMRTr5ohcDYMXZZ4k6CiWOnmPNVGbmIK2GBEqMUZw
6WQG7szvTf3o3K/Lmxnp018FX5jyaz1fXU23Kni8BZlICUW5kZ/7eELVUuOM9jhmYHn2loOmR1zC
ZVvn+xYEyPi9igSDk+H6uFZG0R5BB3rl0cl/WE6EjK0BfgOja5T9k11LCTW5U3HYQluZfziOvoiO
iMCIz2pDTNhnH6lXnFcSE0qGnFYLPACnlerYqvFc8byS5hKXUWlGivQcyJUeSwcarsGwWGUY9yvK
VqNcKT463i7wu+RdNPqt3fl5LyuSznCMupJx1OemfHEYMuEHuEU3gOCOiVJhvVH/S6Kmsvhup856
eoIyd2RTPa0u36QKoE8/6xZA0jp2wYv9d/nJ7kJhllisnblIo3pc3CrooYBiBFUZDnLlsmmqFsht
sEE01wuJMmCh4MlDQFeovMSqs8AoFbED8jSTP/NIAShEBFGZj+roj9Mzj/Rlu6YAoHST3MQh1l0f
OnbGNu3MAvw7AjxLVe6aeK0mhY126iWnzp8fpdijY0aiIUNl4ocVN9yVIdyXqY5PAI9PoKS0hWFV
3E60vg5Q4iCijZrWtJ50OvlY6dje8QfTg7aoCQQkHCk7egLTutyJ/CJ3QipGupz0j7DaHP3DL/4g
9yCWK64raM4u63pr8U3FKwSjolQoKHdTjzLpLNUJiVYXqfWIc3HJGdSJRAd9M9ZtH65X7WbWUlsi
WFCLYCCRapKjqu0idBTuacaSTWPTEnfIV1V+JaBFjQVWQ2/TpNoeM5uCeAo9w5m+ijZ0YEun0y87
JzppTem0IhN5+Qnx7SuZysM20uGnn9WXHmboo0lROVu1oG0I+JLWzbYvCidSMfU1VVWXs9qTIPaX
LgRrErfvwVRO8VBAqxlfgZ5Mk1x0Vqzdq4ncL4taWXqTNiPNbnVNnI03lxEQjP54iBD3PzM8Z9h0
4CJM08TfuAE86mLRHZo/8BIWd9owEn5RJP2Df+RgUb6cfrtJ2ZMn2QEJ23QiZbxP+e0C2G9bdiRm
1wGYyP3j+h5xn4MQ8zlwIjIZwMpEPn6TwHJQn6K+uvMDYR6aMepLSf1D63+XO0tp0ao3kXuwoKRB
KAd+Rqs3lJbfoR3kMhW4SIqfWMz6sCfxeT/UDkRYxSj/ulwRb4+A/GgcMp3s9BM5KjxNBK3+flNZ
k9xxSomY1Wq8HsbuQzu2epkrc6YhZKdCzdYgOeVSEL4vBYuE2Oz87l2iz1rbgE4iqTWmFVUQwPXy
T1BX+lntu71CipTQs1vaT+xf46Jx8om0xVdyTXkis7lkIvpQCpOU0+XG8RLyNPdf7GjKbrgQ+BLf
TP5RwAWwx6KRaB1IqRjKxyyRFfIZ/niFmbNoABhaetXyGCRxJTCUIqbLUTrTnNWLv1T5nXbG5w8v
IsOSso2SxTbV3TkE/tRuuBqfWciE6u5G6L7HrLMZ+Wa7gXY8WbekF0k90E0IsQOx988uCS3NFpwH
/09gWTtfIO58NAywqKpW9urIxB0SryM/28eJnne6ZKvrE7/TCfImxTgvqpFjWpm+rtvvnJUbmwx+
1aAFEgtgHdI2y5aYms1+HwqaFwEHaA6pbckIvemMfpqxCk7siOVbx4ucjI0wWg9RkALjRUE1cxCg
j+PDs6f+NDYjtk7LsPrZw5SO9/R3FjchjxKiWEvUSea5G63FE2p3zaEk5VVc3paz03we6Fw4lFi7
KdSdShJvy5XXDfMIf4n+dDpnpG5X9Sdj92ns69Irk+8hKZpyFsSsETB3g1LuuO3vFnn0CPLVbEuv
f5zvT8lgCNfCzWBAmehraZ04LF4SxQc1H7OKeLcWFLUe4SmdeoG3F8E1IZqCfqblHoNMoeFS8x7h
JMPkNZYAosF6JgR2ToaVsgJv3uRKh0mvrVrUooIceinGP53OO2Te+7ywMI1Z7WQZq8xHadYRGFF7
v0iaR7s7t06ymXsenksqRt7mMRNUi2YRWIL8STDjxjW/N+mTWI9sBneb5aeQw0LQsm4mDi+Hxkiv
2bvO46ywP4RnHxSv3/G4boXOvd3vrn9BTYnha7CJmH04pckao4WC5+N87jtkUaHN0K9aXd66hMed
PfbI9wFGUC9vbSqavOPHFGvkTTXHEVc7Do8+5pZK2pRlPOfsM8oUMI66S05abMfVT2YWfohmm7Y8
llcF2JULq8wvVVYb3DeTI9Dz5Skn+jaHEvOO0u/k/6g4z9oVekKqn2okuZwBGYPHk1YiKn6vIfxN
8bkFDoDfHcmJTbRHwZcl1TigwBRI3nxhR1hbpYPa94jik49W8mnykIE1tAdbQ/jPrJc4WogjKrFk
AI/rGFIGc2arHho0kbbQfSEtYYelG/mnx1MVplR3dV2sBpoZgTfD/Zoh4kkjs84ZfDAS5488cQXy
HoZjgNO85eFq/zDoCIG6JlES7hG5yF7aXmg1Su7NgGum3skTm+sMpiWWQhIAqvw19LAQse+vkx0N
k/NFeSR95QPgn9dEIDJr6rF9GWscJ1fUNlzsFo6MuE5Xsk2jPu6uMhOa/rGhfdv0dav5uQYSgkXi
5JI8+gt+OS/cMSXcdQEVKf9+r6vryxAgj1ELFyh4fDfsGXZ/Pk5ludEdOlv3Y3+eXtwb1KJGvb30
xp/O8vDbAZj1Kp4u5fu+srgJ170X7dVu0ygUgY0NVaEdWUrHZ7Kb09ZLATJQRXb7atr12cfP10hf
Ao66iJKKbJ77lqsfAzDNzFHVuu5rpiFTfK6SDTrza7J5lOKCfTmDJixGFkt8L2X9gFKyK9IqRSDr
ku5neuhrDW1WbEyXcyXkBWLhBJN95ryKqkGTDBrvc5HO3+m6iiqIbta1rjOJ/n0Ig9N/1xDLsrD2
CP++C0GYCar0sfxAGIJWNrAxun1J9jRe0TatRl3IBua4TY6eWCVG9W326z6hLOccFjWcIph4Dzug
RXEC72C533OCHryiGX85RQfRLEAP2/bHqOxPGNFtVvukrAJoAzzXE5ME1Exx4S6cZcW2DqM3YjS9
XO31YaTpyZyt3AE8Lf1xydgd9oC0OTk+yctGrfJtqjJgn8F8VxAYbOPU6iWxINqU8GvlbQaBUMCx
YI6jZKkCnOo+wOZ2xHjHEkD6pZfHDU+guPLJ0RoJ0wiUHu1oVKakISSeC+OtcHEWM/AidS5K/8P2
EirlT367sH5A8/SccPDi9Mqwfzp/5VHHkVy4gasoqq8P/+iP0F/sVwe70EZciXPP7NIhdKcjX/0i
dSnTbdyyhIjIUCtrVXUAAVr7SeE6KXZZFbNveDZ1EX9h72brYuTz59EpcqV6JgoVv1H2S4tLc9Vz
EWxgm5wVjAEWgtKNImAMZuWBpRMJLkFyS3KnsXZgjC1AGVXcZjNp6UQzmrfSmC6fAx5egaLIh7FR
q+oEXzElqefU06cAkFRpygh8xSAE56jaSZ7PUMjRpgN7fxf7s1FSkd0lNr9wFL7WDBZMZR2wgbuY
T7ALH5ES15v3WgeFAi0rA1RcAig3tHZcBmBvlz6cSwpHA8ebyPOfSPZTmUXgR1MzrGWRkXQ3SIrn
gpFLtdP7uWco6eaBBwWiHyPzjYobYjhqANmQQ5bc/wbyhW6HsqMr0KfsWewpLyQ3hpONXj72YuTU
JZ2rPYKsF4ThDsB5Hyu2tPvdUCCU3fleb4YvZdnsjKBe8ibDdXixojiIc53HWKTXqXnZ9Y0qubfR
qwdR/YvdErOPTlFJ352pcVpbE99saZqr9YEWg+ZdfGQOMgC+pktv+f7ZnGvuwblksvxtVQy3rckY
lbX9IxP5A8MThT/QFno4cfWKFG496chV5yPtAXL6EKxpDKlX2rntFu8mowxoWtBqFGwBwTUzwwoO
U8m4OV8zJF99c7zhbEzAfqFG5DcUDeNiSmW/u2dL8apMn04ILUIPERhifLOnfUQQvdQgunib+O50
sIhPG7NkEySwQsqBi1WwHhQgKcOtw/lwSsswsChAOVbszxIGNlFmHY8IBTheGl+mW1vo4hf+nmr1
KWImlIZxoucKlMlvBD39ZkyQJcYGPVNKVBsCtjJQo9nzBwYGaokGDt73ZeOuNaCY+2Mlv5t85liJ
fq+0VWfF3nlYSv9j5Z2VHKnA5jbU51EguHpzq0760SOGc+tUxlaYCBIcKk72kuOetEWxKzodZVfQ
+8M1EoYqUShWaEC8qVwDAaZP6cD+KrjTbLny/SQYYNZaXaJ9z3+6jTUlNd61ShBf5CiJS+P7ZDof
FwjxjBau+oFfexxHvtpk7NIPObhQ9K2iN/LqVjr5BWp3pGj8aSt/LPn08yxM5hhtJFYzpS/2YTkt
1s+SIywfVafIgjiRdN9LudxNP3WgB66KlvByokv9Q/WRt5v5yH9WMUEQn00OZunnUhVeAVgzh35A
I7Rg8Tl197eRzez6VbwvsoECMOVGVoUYr+Go1hgxf3MkZWve2tOo05qIxhXxDUyzVaC12jnSvcZG
lY2tGNi7GLiCoDyz6/Mab9BD11wuwZtS831vnN+9aWN7LI8DALq9UQ8sR3xHWZ/khf5bdhre3b0/
8jPpEpaYxdiSxg3K03p5h/INMMxGsMLeDo/T4phzSmpW0TiedLb/h0KQ/upsnYS7Uf/bngDa735S
8pejXFXvgvsDq75AnQpap0Qwir68BVop9MrE+TD9sHUFktWbkt0t6w1XF/S120M1JrFBUdADGWlU
e6G6BuFoYQLsPeoQTBxQaDhOTpTBAuqMvpVeh8nNGKciVTfk0GI8+SUfjOE/xH5FPHAvJ6ARgosn
l7v/NOxeqqyLUn0XUXA98zSIXkoxXQGpDvp2vT+Y/iWczKNfLUAlvLWIqOfvb9duZGF6GV4ondDe
SnzU6xysjQhOGYtnJ9kfc52L0vAskBDwdqElPsqBvfLyVpFUyqo36WjEceBtxLnBMZ7QSObuoAXA
CzXopieKlM2s7ibty4PXIP3T1ldYkF7n6Yb259HUroYXyulhb4q7I+1hw9V+zojzaOitrkhIcvT5
Luhm1/CKNF5pSq0EXCkKJC0hI0lSbl0R/pr8PnXThD5WoyFdxUxTiKyKh+MzKbxX+OOUnB0Cc0rN
9qRJ5cgRE7/sN6R2vl7lE0k6JSCWxAt4NgIcM+GXRnn4z3xlvflfBdQQyjPBVxMybexmtu0TgIhj
88SHQ26VPg8BtuQTCTM7BLDzn1aU3Rc76mWQZLPHYNP1HcB6tBY8NI+kHtqoBRAOyk+E8ejxVLhJ
oUdMV2KZADcsxqbvzJw5ZzMGWsy4RxJotjcdcWH4dNfKd0UZx4qAeyMmRnMDjOLJrzRK62NNUFlp
eUU1FoniuzRvJPODEoQ7ACCGCpqt4q7yoGrXyOqChQqwGFXt1/BhtMvG1uyQqkKYy2rYg5X69mJ3
QeHxXMEuOy8uVQ6Crb7egtJNXTzf48JBSlRuKat/4Mv9pk7mT+Z8HM5PfTAXMsMTALYbckubDdhK
/1w1x8Nxog0ub7WqOyYbfGTyW0F7aMX2UjSQANSsqSCwYPqfc9Sbcu59TKp333YFR1C8qgrb+n7U
MonwudInP0RyeUR2texlEPgg3EnjKQ73b52l9C5EtH0HQgCGLCTEqwFBrlBwlXhmut4lzHY6TzVN
jVOjVMnFAANza4dW3neanl0RX9nKJKcGpKdfx5B01ojLIzJA4aDuPpyjs7MIXQUo8j7QUEugJ/Ye
Jmvo5Fe4pPVqLpqhOf6CVLpZJqBSU6qbS0Qubj/GUW4BrCSdPUgMABLLsCdmY17q2dKBS/FaFVJV
GFdoHokwbb8fFXUTC9kTshVkhRmOTfpJstZQjit7UCR0AW8/ofCZ80z2RMfmSZ8yOSa/gWVfxx2A
jXpunv2wyNx0vLX0Hx6/7kV5JOakZwtzV2jeq7ZpaVmdABnaG9Ntfj8UyGB8i5jkVYHgNnXLwCDk
sJJlLvC9jPUy5TxTp5CzuxbDkoFGiRBM+oKFupapz0cD9+HA1UTRgC7LnawX9pME8qhkrhZph5NB
0dVznNySyigntYMikhyPIxsfotUwL/QwNRIVoV28B5vMi4lvA+RniOVwkqwUA7zVTX0ZZ89RcnxW
e7FS755XVUpnek9LfIfpRaufBYzcoaWre1wUqsYTtz7xTsZSSRTuZn/E8LUrde9LA3pBCRuyL4n+
EoViUmp+Vjo3BiJ+WQqq0sZMKmkrtKLfmVZyF1hO05wJvpAxXrFh+Bo6R3RUYwmOkZxmbWucJEf7
9CEsYZ8CBGAvvjPsZ13UMRljGu9UWmPLP0ofNk9rGhxtsP2K1+O8WSlDZx+HIonAXmuPY/Miv7aL
5+SA0Atf6YjQp/HopVWnmTddKCzIBNLq4x4wZk/YE2gkQMowBbivjwYAdCyFdIcDX0VD9mNZ5AVX
gk0T0GH6EVHvb//Cu1fXYWoI/lx/644CQUk/gq7sOPc8KHYJItqG1QHh1bjlZgkt3wlq4DcUhkEx
WB+/528E0/McWVFF064JBLVMTIShQWiD/qsoFhxkdLtXI7Hutntm3u1dVT+U74NWCFoRu0Vlbk8f
DVlIQZ5PC5p5AM3V7h1EuO5xrTN903kJ7bzNko0Ijuiv3hoeEbNracOWHoLP/V/irZfqwLqTHi5Y
QfWDFS8siVF849ntGJW/gYKlJje6BormRai5WgRWLcDt13yEQRVsB/3Vi8D8jCnd8ZcFX4P+WDs0
ulGnOOwSeY0yPVyCDdm3FTXQuz+ZsLiUPsHz/AKGbimQygX5zV85oOu/EL8fiBXeUzC7nghUg08r
ZZXChPyVpN/00smbzNcwPSqbbzqk0cDMOpH1G/E0m+ze144CjHZYMRPsMujnBQyC7rnrqL5QCP8I
D5dWihTv3UiLo3bPIzSI/fotx8FB3RgWU8K9K8zvKDZSeJnQzJpkzNw05QvOCvnOta403mMr1Mvm
RdaMXFDVklDVZ0kaxWE2jfZT/xJYc21Bi01wDVJqC72hP0UmxKiAmp1M1Vvja80cR34DmIrsQxD5
KRlxkBWMem7GKplwzCyTlEYEDale4/dJpESu0FEns0uwaeYd9coCHTB5bQpow5zj4lNMU/OwRELe
7HegVB29QmR/N2oBgtNlIFQrQyWNt3CS2dHDf8rinpQmUIpGS/PjRjKkJQ0U4lYu2EsOnvFpe7Lb
zhVFwAfUbSlG8qPf5MwJCq6RMKQy0SS43XqT1J6DKeMtH47J5iHU/y8OKT/ptw0Pvf8W1qrF3jTe
2NyfRSb8u/aIL+o5H1yr8lDEf349qGDBxF6bC0p+j8rZ424YtFxrig2Uz6StviFsjwFB/CW0oLzr
0e7gAnpggJYV3nKdnn1FPW5xATfArFSCAp7UTD0Wkx7Qe56pijfMks82KWt21ZdIN+ITAoeJD9a6
L+kWQ3/w/LcL/NwgafjZsGW8ULOCYI9s9iuPx6X/8hWaq4ZWTzDoF6tIDn9lYE49eLR2S0rpTpP2
HiHJnuHSCr2k4nkMXzNnD2SNQou3CtZrOWYWhbvh39xyOPUT3dL/5vlo65rPFu1iDx1kSQBtSkIC
oILW5SeHK9H3Bn6WlD8Vx8RYGrQRFSrkuH5sDhuJQXq7cID0fk9DOU16tOJCggWM4Z54Dge+o77P
au6xk3zcu8xDW/cywnkx8Rf8/XzfVUYHtOXBaV8zITOrXz/MJrUHrsFI6ojp5A1eZ54l4y7P0xCL
ETHyROw1kxIFhNLAVmJeurq9ARFULodpwgtrrh9LlqNQ00TzXItGz1zl6Jwv4xvcCtWMw2zuhEpu
lqSW75Dj/4Pf1n9nz1N9lfjKIClgXBOKdLJgE0a0TWaf665516g3krC7znbPof/k7KdBsRGKPsuO
t31B3UyjWp0Yo6EZruFcT5KqFImR263ttE+OBvpLq8N1x3MFMUu7cqaiQb+Jx/tJSv4rDBg/E4YP
CQBvrjlYd3Ital8/zY1iK5tltp54A1sYCC8XBoeuHmxCW7jGN4iEhtOsrvHk16H/eXJA1hubIR34
hiPP475+uWI/aHVO62lK7YgIafbSiBdRyHr2lRqE2+ciALp22hh08FKAo5LwvZAKqaTvaBlHz2cE
2z59YC/j0OnfUCnww+u4IKXx7/w9rGAWrYZAnXjYei8g1bFovVlsuXJIX/M/ZlXOOTWuJ/HDza1u
eIohnJ4IP9neqwmhiRugZe1CgEyhbotlNX9mHs+Wjt0xpvPBNxVlWE18ecbXo4TpSOhraGC5fHlq
Yz4wy9iZ1e6UfZ+4To6n2071NmiiII+9mS0z16ToK/zIvT291Sokfzgl+IxFMS3v04fLppkEOhxM
FhrisFSPfrGy1AIj2x4Tzoem/Ll94R+15cQ7P8Tik5iChYeJFLYYxXUvEwIs09Ss69ePXVrwX0xS
QNZ5tABp4G2prOgiLGfwedZEBN9AET9aNUjf6YeJBTTV65yF+IWvxqoGd3fMRrumNgEZd9tYOP1n
ujs/6WnJeEvU+srQXeiM49aV1toQO7innQMPr4Imp8o5bgoOeaW7CE3LFPkSaEDr3n8cKKOBVgp6
epsU952TBKxz4R669B7unUDCicYtnx7VPfVbJEEkxYz8hMo+sGTfnjMvnbzGiXjHypvWQmxoPIMO
ncwW6bzm49Wzmx/95KWD7h/Qw2lG4mgF94vNHUH/hcFKeF3+DOhMwVIait6bdWVLJIz7QopYFxUU
V0Dar7kIEZ9E5iBmifQVtQrdEbxOR7rc+JqjvNzl6k+5qTndqAFpgYH5iwzHjDgZNiP2u7KAMfJ8
aN2kP/O7uYlOhk9KorUHJXJqWWRhrHmD1wFbn+B05uqgo84HfMPwW0crEffNjS5XL7BPEvEuuXnT
org5cZuPlwU11K6Xbusz6CPA6qpXhBHFQ6xJDCOXYX/Z9tJir2ZghP13qLhqoOHvJDwRlAabBR+7
bc2Z0v8AnSzpwjq8ySTXU5QADCzsKmUqtIlKNvzQJtQIqGJOenI7cP+YLtpiKduxAFY5k7KvLuVE
GU1VSGapZkom9wfRw2Y48aC+sIJU+Xzv7vEl1YpLtFHXcCQdEyzDDE3XbiSGk2AUI2I0btdbuvgV
4/JNv8OTz8N6C6mt5t+bBFI0ypgeeAAu1gkmElmmr1wVsIGz5M6lg+kfu226Iobz6/ZYIqlziWPT
On9Z+E2lsuJq23OUauXm19IigepN2yCruR9Dxlzi26CeE//Jbb0lTjFUguKJ0X4A81nN34TGF59O
NTtxgtpSeVc3xBxUnFa52AuqMgceqGjE7tFIIoTVLrzUvw1hwkD82Wj7xKMexczll850hTCymPFA
T61zBttmJu+afPZk+K5J1B+aYHilIItbRuyjc6j4ZG7xISc0T+Gu8tkGtFA7GWKyIuQuY3vKe3Zz
yFqTfkA9pyMym1bS+jEbpod7rAoDdXq6utJqCIdde7/wEN7ueUiNo2D1XocZgSRROIMqLbfMtuPy
VGaQoYGBdwlW6nULHAZII7Sj2h8oqLAEUuDJc60eQwqnUoXhzty2dqfyXTN7M5sp84zYKT/vo1V0
D8yrBlHwYgf+fHAun3xTXYlj+/VBOtG1/3mf3WBVwReOwk0g167A5M+eFN4704jnMiQcIFVzioJT
o8hQNLRuvRdqzcDujNCodXDTFKZHhnVInRij/5BA33KwPcXXMYNzwvHp0wGLJFVfgV3k6uynsnD9
GC1tQrOS8qDYjPzThwT48Jiqx5ULO2GlCmi1y6XDrhA4rcCVGtjrL/0+kwEixW9evdzM1q97PRe1
/rVxtaxVM/tOKxzI+4yMiaqNeSb4onGl9wakx7dQpUC69wK4vXRpDey5Gi/gkvJGViKJTuollcHk
vi/lffpfQwBSqYmhwCndDOOuJK1GZVjabyjPjnjmXQCfEZ+/pcF2ME08yXc9P+C4Bf0k82RWMoxt
Xfc1eMnp9iNODhLqitmaD+ZMPLlkymdljwp34YlZwhD6cZKiENUqU+2ZjodozkBsQ4yt+Ia/FmYi
pSI7tM2tCl+/kSyqg7XDTkZEtCIYCS8EA5dxXb7/WL8i0/F9Ei3nmhYLjUvlnZHmKKGyX1yd3rFm
O1HODEZY26/M2Hh5LSEXudhqDXcezYhBGqDXF3gZ9Oj2Fy9G//8nnhv0W72Mswukqlct7oyZty3A
UeqLa0uNCRcdDe69JF6EZGEuhNxQmIq9IUtRRTHtI5VcFZnxDW13g0QEN1ULgvlJUie7Chbrsigt
6ZTGfV73JJC7RoTlfnmglpRRj4qvd4I87KHddurCjLmzov6GOTDp2RnbtYOrDo4OijJYCbqe9xNa
uUqtRkfcp+CuoHJPOP8GATQoEptbLlWBGBl/Aa87qLH3fjrUHIkkHnSGa1vX5ZZOHShzffHUb3We
jP4RXg0mU0d8yp0ZGW9fp0ove5qFQ73Ariz+zTdrn2vlVY4o10kPmrAZRph85XnkfsylUXF/hMTF
Y669GndfaWuj6GDwDZzraXNfQG1Pqhcveq1FUk/AEEX7GySnMd9T953wdIJP6gI2pn7aBQ/yYEXt
BiB/mwyojxN21NV9zccTxDJtfjiwt5mLORU7BLvqoRr7ONedwQczevYNQoito5BCpwTgUtIQmv+p
w8AaKqj1sgaVQ7yLKRQ9MOA+s1O+ohiiH/qUHzbnknqCUivz53unPvVLsZBk0PNbxCAtj6mzQanu
vXUG58RSLpbk1sZV8rBKzZscbcfY5W+iOOTHGRpjUnBSvvBIqx8CrO7TVv/QEdmf7uHrSjB9dmlk
ZguIz2ZCGVpg9iUfGV5kHAUgO+F/qHquczAMKTqiGDiCCIrfJp+hNbmvD83fvyTvhuNiMydrlUqR
zANeIe82SZoIMF/oLaaALai+J+EVz/xr17wqLe4RM6+QGb25QcifVY9I8S3xsFVU/jh/5aw6nK/Y
VzZOHNPitBPFcuD8MN4UhhRFSkurSGPJpy7Ofrbe1QNYVJNWebbQ1bcPqceQjJJa262OFYTSNeCO
y/km2qIl4M5ymlQAUSixRHIVdvHiK/kxogSQrzeZPks26+pUnJEC+FcqAfxrMKXsgOvs6Wh/Jgve
VgweIRDt+JHblmX7vpJOQblXqNtH7uV++l2rf7yrw5Htqy+mdivxIjvWHm7UzXpSpwHBMAW4qji8
Lq+XlW1kbPJChzUWIR+ZZpn3szAxVqHLVCKj7EFmP+DZc6xcjdPf9FDWdN3EGwDl277ySLP3eXwS
2W3+yWBjt5y2izNuoqj/JW5ugC82/ektOu3nxP0rOCCCA6av0TLNUuUenG87CqHrQ7fvJMvpOvGi
XnZ4j15waTdPySAaSFw0/C1qA/lj+f4qeujeewn6vkFlXeczG/0For6jlxA84edAnhxd7mPMUGmg
iHoeRORdOov/oPRSSkIO2niWyIS/DolTvVbLbijmZoHXbgIjW4meY5w+c2ZsG9KfdMsLotCz+Brm
AzD3nyCyx2G9GI8sbe+0K/iQ/zTd8OVcaFYkekU13cnDBp2Yzb3r9PW5u+zk9ToWO5Nv8qjmwPig
HT4/qKXkM6cFmUgmEJU7djaAj7jV+xd4FJ2DbXPK15wQ770b/gh33x6rzqLQw+FpXFUuJve/dmIW
mJMVjJuFA0gn5e8NDzO5TVPrHbvnLFGBwAnNmQiZKYyfGSEDllYKdOn9Et0Zr7Pk1lZnCyB8yGDj
j2z5UY1gACLBYi+fyNjuH2j27BRCOIqRWx9lsBM3a8zVXZwCfanW6/gRh5BFpgxEFcVVqh97g4R/
bkKfzipGyRYmL1JlJFzF/+59Fbec5ml2oBompUW9QWxvA34XY/8n+pdFCvVYYxVdD+KiB9X2Efg2
rB4tOH4XODkspWBpvOr1BGNhgftB66ObY3ppZnUAorxy6TIODZ2z03YNhH7lxxVUSm75mSYaywtQ
cAVUdd5TRinzCt2bFQ7FwHP9B7vZAx1AHLJouyy4RSssFBeMvecD6OAOrhUvi3f3LR5qXaZIJm9J
5sWmJosp5EaP+h6C7CWYswrH6h2ad7LOppOta6ze6sJSZXqUW6gJPQjCDJnYTHn2YIPMyZT+maYT
VLuWCfTx1zGET5OqYRgfwyCEtsFKIoj2K+/s8FlGUHD6jhBbnnOKwrMH9j0h8fVCQeyflFtAx4BK
FEiTq0Tcrb6uZMJb9KESLPhlSDFilQFw2O3x1iiNbocAH2EZDDuILON3DZsQnaRyu4ARQjhEWCQs
CKm6DyK2Gc8GqSwq7+Z05wubgc2hpZK3XHrr/MLkAiSzibJ4/vDtsqZGVb8yUlQ05hggLc0aqDuZ
3U45UX/qcrevq/c1BxIeke/UqPrHPDJP8RVPReuSM9mGyX6nDqpiLDdkCvuztBMG/GMSqdx0H7Gw
yrCE6KAOPYNRdV1OvlJ3CefQuM7utKCWVrpqJPu5CvO/Iz1dZ8lwq2hDjzcG4BtT19rpz2BWfyzh
/dil8pdUqserwDODCBjpU6BghlrBtXFeD8uMoh75oqTbDEcCueVypbe7sEqzDqyWKBipHmbiwNwH
YuHdMqA42rX7cREd92nTBHjEuAq4UI5kgLYS+O2sBfZP+G2y5FaV+zCYeclkV3yNI7AAoDK5AxgQ
2q232N012ruMRiLVfkzFkFjykztAcNMY8YjqzQmSSrrCkOZwr7GeVuHziemW/ANsNkXJ8FueKR5f
OhXZpaE/GmFtoZ6cwXqNN1ztJ+HrwjHf0rPyX+jWXKFl6d0+ltbNiy01ehwLoKElfFuOlfiuk++c
SVFngIeEkG6M5UEv86O4/4SUpFgrtKcQGnk7qztHE1dji4cijA0xEF19p8ztq2fzu9FDt9c0ZD5Z
VkP5loS+8ZEzYZSsN2UoaT/Zdw5CbQ+kk3X3/RnJu5GhIIrVyiLrQ8pCNX9jqvv+l7Pbp47sw2pV
i8K0ju7CMO15Qq5tvT5/UOLZDc5S4xJFbfk3bqJH6pm6fJiefoiP6OJcXTFCyOK9WFk9SpZ7o0F9
GaZ/QnviBBq8lUmKcKBbYrZrfygyCCV425xxdC3q8FJ2s5ddvYFRCHiCGRSHsAgI9RYcRKnMkIdg
jQ/hr8s/4q/0zvsoKXd/uiKh1sPsrNyC9p8zXxgKZihYRJKUkvIiDRhB9Dlao+G6lBW+Bj7LsiD8
2epigkBCkMe8o+LlyK+GXf9Ks5qvfevZWLSTUcnq4Hs8GC4++E15mRqS0bDAC/OW6vT2ewSonGtR
Cax29IL/PX1pQ3cuGm2U4g7eKg2W+o8Fc4X0o1Wcqd+zRj6Wn9BtJK7Q37JBmS07n8gnOgI171uJ
E/KdRrOWaCM9MF6F/i2pPW2eUy2liDXtzHfQQTu0n6gGzRN/Ob8DX1Hh/xy+MLrGIP2y6lfxcTLU
sQVHpIw1j3SbdqjSIQfUssRj9pDtDk8oa5VV/cH3rDaQHGq9AplMgvyo0VbIOkF/ugV3Q9hoDUQ3
oqEfOPdEHRyQjLD5CyFxvrz5SHNzPhTdq+UAAFJQqi4zZUWY3zRZr+WIJGD9JfJg4zxQ3eegiMsS
q8ya/fRXP+BHuU6eYzRHMirZwlXSZ7v+Pas2iuve/r3KLoVemJtvtDYkpeCVrFjKr1Zx+ZBOGI5W
Lt9dndcmR34wqA7lXIen+stFhSItSus7yrgQeOGocE29e3oRZBIJhnwUzhLXI//dHFP1NQZ2Qg8n
ikQHh3jBOKzh61PJxRXgf9AtNd0aMBcj630d1oKX/u3VluhTtzQaA/7Ym6wqtKEwOeT1pdfuHule
1Q0i4n0mwG4/Yf2n5LLpZZcxiIEPqQ421vG8ZJzLxk05+9yC/eRTXj66g5iHld6gnJwiweCpgoHB
ZgQF0NqcXQxGXad/R3Dx+0vtZJixtsXEMddoMDxI4fG7akRVhcOkn/WwnR6oE104gRugHOtIKww1
WcO4U7FWYf8KHiGEInV+bHGYP1HtT9olEgrEEoDGh9N7wwuw6tMTQJARWw9HRBmHFMx21bt9pzTb
OFiEw5mchbSuK4CudFoOGfpAfTCZzVzkTLc1cpCdsnFloFjxwjfrW3VyYUS3DMVMFehe+54q/hlo
dX1M0c1x/10k4TNebIcfUZ/TG+w0iZc8bXY9IMW81SvEd/ZnbvUclWGrEwi0qc/ijgDFPZQnwRMh
m6yBkscA971KZ+oHty4bHfNHiXYpB46gLd6jLONysQ2fJYITvsS1O6duReAFrilcm14832Qb7vvO
80oSLXOM0gKfI3iTuQoAuYZGSAnF6IkfxCgpdTmOr+5mFNe0neI9EL1KDH25wBVJo/K+FIczP+nY
Tl8QE/YzXL+lqV5uPWI1m2VxSlVZUiGOZOs/Bc5dmeIZawI3tRG3bhF3v/ZQgYCj9nFKKrAbVn3o
WQbO2qnq4honLTDsAYTznk55zU9BhiQqibnNtBuREgmza+CKHsJl9UI+NxpGIOIoN9Y8gZdXygQl
x0jpZEFDI3La6hrBC77wI2jhgnumlZeNw+xjXuEVrYfLli7lvkqPNdzKutHXpTuuGZjeMiUIC55J
32bWOuc1yVTZRgipBl0LOxEmKqnja7PV0ICdJ5tB+xlmDWQA1uZ7uJy/X5vuCVZARQFKCFIW4Yk9
Y3IaTNeqXD8z/MX8BFwCviG5L3oPVFnQYjYlo3BQIEDIHjsX94C2gFRBILJMamdDGKoIRva50gAM
/6CsTbJxrqMw+vDGmKO8NrpdeqbyvJw7ICwjTi96Swc0UuKYoaSM8ZyGHWlBDwF6CQyaVUet7h47
CA9/RKtk+okRCtJKKk5ggUmor8GeYF2pk47SA3fM1XBsEBYuPynE0INjl6DiiMoLWYicqmbzedvX
Rtv4EMMtnECCVhW+lQw1AEuZYJOwwWrQTHgqC7N2RVzqQkT+5JOB3qfrVXlIsxtVR3w4iXgEHj+I
WWrMW/hyN3OuScA6vP1Fm1zM2ey71nDmcq9IquIuwtcSo8DUEveqZHkQ/1WgrG/hvJh+HJ7KbKK1
xPk8OcfJRzq2pN8PGaonfPZrdM5c7n8bOeqyPhM7aq0SdYkw/2MmaXQ25B81k0y0AsVlGSuZXJvA
txYFoyoFl/iZjuebCUlI/OwC2jupHfkQ5IKcRgyliDokzFypOtQjvhvOgZLm1wMbvLbTq94u6Fd8
5/jmWwqgS3c+iis0tgAGlVXIY++F01X6Ql1qcJ1fpxlRR4IuTqWgxkKxF1P0ZNiQO4sdl1DMi2Ta
bi2P9geqRuRugFoBmG6GApH788idhMZN5oBWYI7XhV+3FE+dAyRlHp7vOy5uKxaw6SlQsO560Ch6
N+CTJDVoKrbNo2OlXWW/Qv5DPpftoRJQbzzOwVG22cR+CSgw8p0Eo9QsJTIiG/M1if5NFOymvcBJ
fazpW+rxQGboRkLo0YczR3NeZXmheNb9NYGp6/hpvJT2ARgmgxHt6kfVQcamnbuf56tWhE0IHPzc
3QmqGlvQHn5K5xLN+gG89966faYQBGV/hBTaYGHrI2opkxJIilzRqBuY+ZKsaLusJ6MaMep8juC9
DVgd0bbhbuJeIDiaeGE9eu6CJvd3AlabTUn1h6JUPTmOes8YinBWSncwntzph2LZjlSPUru7p4sS
+8xRXWknGFC9Bysn+ioRV0/NCrGx/mjrf2npAekjx3fZkghItk+9tY7Q2U82ym+9EBer+hyLVeoz
fkozSyTjo+hBRPoDFQ2yX7CJ5NXJt1WSumfwYNCOv1C05J770EBqzyDQT29kX8DV7MST1ppyDtzA
nHbZM8vfVnu+mL8YT5cvM5K1LEBkFdqfqina0sc8yJMW1fKLmchoIqqGfh2du0yI6spSV0a8Ldvl
VLjXGkch9vtnNzhyCBFOGPuOrSEgZ1SZoguX68jJxF3ceyd4XWvqgx67NSraC9KPBjE6sbM7CKkY
s/JYnSXlJl1KX0KoSr9fQGtiqlvV0bDB4qwMn6mai72tvLVWdKVcAOBUAljwV2Ketx+MDjrRP3Qq
gu4/qmwEfIHINQF36Dux/FtlqqE3ZwGKWnb0ranc6EYzkR/KlTDz+pBwsgi8OV1x/bQcIOdHZ18t
fGi9FuDaIzl4IT/9EHlqMsUDpnfIVFtDEMTGPlp9Emrxc4s/AwJH85aqK5WOzQPRYCkIUmGTH4Lw
g+WRZWrQXEmAvDwwRxmtDd8qLD8PmOiKUy2sxpjMxP6oKe/R+mNkV5iAMg0IhwhHkBDNC01UfnRJ
C+MsBPAYS/48d30Y4iQualzG6CBeTxJ6CUZ4bVeCEMJWT223DEi79E7kYz2KPa032jXHUAuavouH
0F4kGXf7F6hD5ARB0gff35tna41T0ZxhAB1QgG6F6bFj6GIGOcFu/IVSwTo8NHhYNba/u1M1LEB4
4A/m8XqwapDZRDJe8dI6Cr6eErzId9576lw3RtI1+djOcwljwq5LiYFpsi8rRtySIYFANyl9E2w9
vSc2WDYt2fPNAOaQm3oEIYOWKDmx/Chn5v04JmxpEGrInBLVYkj5SYkNkV5fUwTdwB551wcCuPIv
Ft00dVshOOAXlpUAC/c/y6IyNYGm9q5ToFg+Rvh4QaUyFDAizvHBxSkfMB7tkgUg6+uAono6tY+r
6cBWDGQ/m+2BIRw2DBYk5ek2Y9CcVhNBz3BgDwLWBwKj3QJMKv3c1+qSkLKJ2MoooKHJhYkFIFdf
Jr7ZmYn9livyefsSu+j+Jp4jFU0DlRIXtKX/v7FYso9vdfb+ClkNyfz8/WfBdjEaWsUPrPCfo8tO
Vzn2k1hNufbCZvZvNAnvqbMXbaU6MS1hEEsRwHNSyPKmlb+A+Odgp0idXD532Hvu4aRrHDO4FJsT
asWm5YSUxa9ev61mBlBqUD22a4EiJyA58v98i2iLaLO6wxjLd5AkYqBdVALnawNOHWERx/Y/8CXJ
yWJ+IbBflEr/Axg9Txl1SWtg+n/JAYJgkrbMuvLG5PblgKkkSJSk6tTZhLZ8c6vSime8AjAr5QX6
abOdZ+u9JqLEegRvCJofLbqa1ZZWP/Wtgrfe5I3pdB6jNfYsulVYzZ7ucjpKiFRmXwUiX4/HKAp7
BuzUCKorz2x1upBXtgc8FkAAm8O+4yIr+IWHoC1wgRuL4FzohDnES5Q72uBTkzrg33ojh7Tx8bgm
o79lYuGPDUDD1Sq+I0TmV8t7Bh2U+cZ9LXuG8XKyEHydv5Cvrf917+DkGpAv+2MTYN9XOkUHsTN6
u6zKWdPhAzbw2xdPeUcdkTklT22XJTP6UGPfg07SccJfT9dQ1cM6c6IvfTrprD6sBci78V9tcae5
7orLNT8su6jPmtBla4qfiZCzKWQEJMmXFxPrVDhFoE+ebKwNnmm/pi4AIJa59hH0gMEaxAEW3JsH
OyV6HjiKmAqmlWoQuc4z/A6tOh1EL9PEhCgqebRjX6/ukugiUVuMNTgjppvyKZM92wJfPr7+06JO
Wcx6NW4bL2d6HIL8XLOlQxvwddHtR3Jk2DIdEk7I+/LfeNTv8Std1Chssfbu3NaRmgm77UrmYxRb
A2AVJNaDufsmgxg+YKtiCkxlHM16fUbMFFdkx6uXuhTEZl6msC1SSLuJVw45uaFZVuwLwupXD3E4
dma1I5PJzBhQBwv7QNyqN0OxJA+QvVVDPsDyiCJc1Pr03qk0qi4E2+SLHUT/A9voOvW8WFv6q/iI
M1Ssv3aaWlloX/e0w5JmjI6n0gYPIQJ9T8WsT2OMQ4hp496uCxD1ZdvIglDhtD4bH4wG8PTrwAAg
I+gUzphRTB3hfMzcljiB2LVUjIU7JUft1KkoqzPhDphIsVF3DQ7wqei2XE7r6eOJdU4707WlT8xC
WrXIGCzQvV8oQ520tDZqx233vm7+7pvcVwGJ8jKMHHSI/6x0/RmF4UB96fKoebNlUFHgJGlLhaU4
zLyA4k4tsYzlMwiMlAHgbJthr2yvrw5WFenGhpC7MrurM+MfhFrtlv4vKi8wtGvtAFNivqQn/yNT
lmduN2lRWx7vHvsYF6zQpRKVGDC4FIGOI3YQUALx9AeizQdyIkQwUL1SYxS7Md6q1bSCeGLwyPVT
RTRUDuVfcGUypQG3ud7MhxySLhc8C7iz4HOcUBli284kp3HhtJB1H5tZyqJcZp8XF+kBXSk4xldv
Ik/2+Jg6h7F8A8mQijqMH90SDaRIT3bT08yS/lnr6ls+V/vzpGuwLnOsgosDIqacNyOVknNuhrX/
VdZBjgtNthuGpC3BW7/3Vm2hwhvW7CrfAgbyVnsjbQS+qPpL9feSy06CaZX9EKGj414Ri6h3Oje8
OwgJdEK0rfootb25XJ8KrAqPq0119+x22Sa0/uIok/DDsS5crVBkTkEu/ozFmhSBF/xt2SxqXDqm
dY1gPDC90CyTxPIvVctx+KVL19brXDBwoAPR55nthHI7K9mI/OERVcAbPfBsB1RAUVKHCcNUhMxO
cuozIezYAIBJJTKyYH+qI7HwMPAK8MwJfmfZXv0tKhbpxt1NBRg3x25+X8RhxRc3wzhAQDEv5bFY
/SENx/YmPjgFW0jVYXzx+Oszr1hvy+6uFFrauDycFNfBWsEh2qL6FvG1kwpi4U6ToVzttZXlroiX
6YXwqa4jFVb0OYaKVUUyBfy6MLhQRRkaEClgWJOLqS7POVeHP6+4KKIqDfRP0dUXK9HipPeHVEcY
61/8SLffSwRelyfxuLW3uwGSwR1QmDqMFErf5o8L47fUQGyOCdVU/NH1H9B04BtPeKVxPCkJ3tuC
KtN3CP9ikY1y+gBFmDUljuS1NbcaKVQVDPW1eh6POtecZUSZxQkRy0ClQZIPWA30ScBRknrEnDEO
4X/5MohiCgZco+KjqAe04fQM6c770A0SWolIDP8LV7M0fwrYxP1uzvIECOxVytMHlbuBNOKlYhbe
b553E5bxQnYBeUpwFPBhh1RRviY2VmfE5z7UoivIcK7TP0pZkNLQlvnQToOibKqqlMiklnpybfIs
MzN7ehS5jpJxZB0L194LMBNJDA0BPupcPccNXu5Yw31w+yZjhqzZ9ecG3WJ0qKH7+R3VtpeZLaaf
hywQWcgVNMLXH5nxOi29tLuxB3t1zMNLjIeRz2MMJ/DKaR6YvEx9ihI/HkJ2Ft1VEpOXH3vsECmN
nk2mS/rpTVtrtjKkflor8iCZYXmvqvbFpL+gcnDDZEikD+L5I37XyuGex1GpJ4mCsViHzt+H7IHm
on20j+9DL8RGKql4tkxhSjh7VmeIncs8BaItO43eSEWnI9Rh4IsTFFQjBrOFwNNfNEB2UgxGImT4
99PB6W8DFwU0KQD7QPRUiMALil0WsULzZe6OOiyb46Y+U6qa6RAeDAuEQzw7Sw9yBPKiKbfwLjz4
PY9Nf5XcyKWpMjxK+8aEo7patAh56grfQH/Vqo0B0hZSgCBG+LLPxUSBQqK/1YHiZO0EefKgDnLg
x6VrDSjHl/D2c/M8A5lVMDfQttiHlvWZF/o+R2tGAMaqPSe4fIQf3uuy4NgGbRmrlsNXFMQ8jnUX
1hcld4B7jG3yP/OoSE0zfXgxOJ1RL51NAVoj9JtxmGcqZHwZ/e9429dYtrUnpnbENp1AzBAQihgW
jwZrgs3RflMZVpTgStUtJdocYAILvoG2F6gIvJrMscL+Wxkn7Z/iIWUK6uzK4Ws+AcdKqjJQxV4V
GqHDkImqdtWf7yNcf2lRQuPB195OhKCxE8XnaJmUsJpptIbLd7dnuabnL72qkAW8G9AGerHk72bp
Q0oup1QWc7vXrreMRehiPJfSGEk/vH7r0tZT3Wil9xOt4kW6d8KC67oFhYYjMlS0jm852W6py/dF
PN4pur8qvYoVg6wIizgOxJLMXAmgHLoDRhzKXtpinOUr7xBqHPGm6IkoB1XMcHOwfrbddccCHMCG
sLNvr9d/8NqhqJ2eDev18SQelyVDCdJHjmnaeeP324QwPajWNXasvq2ZqgjOoHVao62DEPUf2Skk
jEZn3EzubOdZf7FdS3n2Lpo+ArMly2VhI7Tm6wYoOD5FP4fTSQDD2DXGXBDUMmT4hTudEtDeMYKD
BL5QSR7v2F7ywCbxGsEXHAw7wXbRZimCs7GO4DipnUxnMRwi2JdHX9md1BLjFg3LNmGbBmO9Ii8V
vNVOqZMUl2lQeQuZp3lfZBXSQCjVK5aTKfnDPMbEmp9B5mgR89kpKE75wn5PQ/YhQ400Eu1IEjJ8
564R+q40Cs+NbpJTCUCg7E72Rmp4wg7CBnzs40ZSz276Y66+nqSx/W7OcO9gb24KYw0wGwglFUyZ
1i9aOpggqoL2z4ZCHLgqe7zt7QoWKjXkA1KdFXx7rVeJzDJG0q8VfGNFcWWKTVfG932NOAOPA8no
iOaUNv0hnUGn4hrqjgGadvjyDbiL3VC3lNEF90SkrRrjA9mqkF6KmbsrFV3hL82KqLqq0Dxg+C/A
7I6P14P4C2m1fOi53o9+f2pKXMygSjDNfO8sVCoY+jJUe1aktUj4GP1dAXfCvRMerUV0DSgFIF4T
rLMtCX92BsmD1off0ebByV3ZalJMlutBMQDgUw4E5rzWAVMHHKYKFSlN8oyl3ugZ7LerGLFpbhzo
QLgBZK2/e86MTbgYe46eQIGg9P8IMajwVOhZ8+6wXPI4KEKp99d4/FwxQj2lOCCEsBw8q8cjRs7U
FC+jQjxtDQ6lvIiXWAk94jiECBp2EE00V6xBlGWV1FjU7GpTeupRKg/Z1NHUC07mFU74OfyTrlKl
g6OSAuzp74GelWWEIZJ9fEwD/IEypEuK4IWjh/etBeX00inyq6HZWbA5/tS3rD3CRsLxfCzz0Zt4
/Outk1aC+ImskXjDNwEcx6Adyz7RRoR2lUF25UgtX53OeMOYy6acQdFseCor8VEkmF1tV/zGNqe5
TtLIM4kesxEAKnCQsc+zIR8zp90OjGR03FxUrvpdHdl9ZfYcFd9SqJtUtfHyeLn9gyh8mWEZIBCc
KmP6jEruTmDq65eTEcesNalWJ45VweePj7B1GIQbUKUPnwUx7tU31JIgTYIEeSxfjjJ3JkLk4ikO
8jFwehfYpPZSlnET62fSvrU46vJYbGHvfuB35nJDhp4J79aGua5W+PwZlXiWp7loosaDDusesYZF
RhQwyCymdK6E9wOEN/V6B9fw4SP5IGp/yZi1mlLMku8Pbg4oGZm+mvqGlt0XH0U4M0fbAhUlFADc
FEHqmkgMQ0u/t81WkvXMdFPqhPYcxgsj0axoLTKE0mZ2bE7V7MFh3X/MWsrMqgHTQArK0qz3AlMC
VuIjfypLEUuuolvZMXP2eAmvWz1uptAMJjYm8RmHS/4/0Aa6RM9mzeTp0ZYWijPWKzFUoryMIc98
AmtrWnoQYcjlKxZs0/TjQQw81Btu1sVyZN0D8RH1XS2klY3gQFzNhzNvojJ1BboyTDfKQjDxX1YP
7YTdwzWakVQBjXwXsZrVt8uwD3GKz5qwsfKJhUA6SXrye+654XY/ocIjr7SnBf1a4R3H6VcoF4mO
v6gEfDXLZQsLpV5PEoSKKSC0QQ0BZ4Lo5eB6Ctk5fpKkxu4r2AqGKzSSkTxL9KpQ3ZF02qUlP+KZ
pN2zf16jLW7irMrE9OxSQ6ABnTnV6/OtATQk64okuohz2VMiA0ubL2VhCiw/ofi1B/xcdODnJn9p
sNjHzPy5VT6pAMrYCD6ovU+3RqXPQi0a/2Eju1iaWmPwvUOL92Gu+v1oO4YxNZ321FAXAFbuVCEd
ZcIFN2UoP6RKA4hl/44+27KNiEPmp7MjgxHh4e0CWWkDbI7Uc0StJR7jj0Q+PVXXyZjNofdEyrdx
K80HQKNLGAtZhipM8dIsy+qeXIU1zkWdmHTOOcTlWa92ifMpLScDjVZD7HuvQDxGjiIyCE+hMiJv
HIC8utudRejFpcwe7rXpEOk29PdRJplbtamQYdk4vyyzkfvR+jCc0trwJmPvk8wU0Ynvc9FGvYR7
4NuOl7o0IgISpuP5WfXscSoDreQTNYf+et+kBpc2rR8SjVeYf2Qn5j5UcQnwSJyHk0H4cNX9PqKe
JRF10t8mWwVtw60ekGmSQ0SAEvhKeRdEiNnaJmpCgkiODUOxMf7qdf1iRiFpccbABr9ZvbWLrw/O
OW7H5RcvE1gzU+UY0CgM9rLn9T0vPg/rYGtWNktj8BiFWyPvD3YeMpJDJiARfF5qn+u+xDyMlNdu
Y4HTn137qt4NYlVyQL6DGAKw4klSUbDPgfYGNRukcg3rtPsM2RuW8kY1Hah1UTJnXE8kGEavDnqx
bEhcLMaSbqG7b8u6CMe4zlEsK9JrZjk4AWpE00hSYJ7J7D3eyGfiXzhiwlrQVNuDBhmLGJtcAV17
N460dJ6eNX3rpQvDAKz/XJ5o/xMI+Sfs28M5Bsq42CPT6Amhe65wW2Gn2cM+ENq4ZJYU4p1or4q4
G4aRlkMgH7ixfic+rOgLW5L7+A7VWAMgRQDqc1fkusnfbqTnqso/gO0FGArJVlwvusNe8RtvvOI3
slT3vd5yRf/3ZTO3sRb3rSKA48uFbHjx9+jUROebtkLQrgQphijMLPNpE82/8shWiCAV1kueHL6o
6hxi6y4M7hf1DpFIh1+4d/rfQg4ckcSQQ3+T+FWqxcSm43BJ+y6CyF6822HNei/c0Auz4zdE/MiQ
edsuEVMbjBBspk+SKxomsIOiKX67hTFFGXDUBtuDx3S93ucsuH+lPpkbmAgmWP137pwqO6eXCjn+
fmkRkmbTNBmtL05Fg0Ax/zT7mCRtGZzKHpfsO5oUSNXQeM14LWcfFDBGZQ7tf31LJU+7x3CU423/
PZZXw7e3ZCzPvsmKXiB+aUqVvQZNfK0q8RetHN8HNBbAOWDjwBcwaOBTIca4D5F1LIrOqL1KjRpI
cXHlPrVxZ8aHEA1bVbgwFQBqSTsAWuMRbhzjtxfWSxEXxue6GhET6kbZcbv4UGLmFXUvRe4FCApY
LE49chODe7Q2LqgVb55B19Hzw7snidyTrYDPJ8/ElvwLBG/RO0OijIXm3cD+qyn7rtpF4lUBLD4X
Vq8MG4JC6SYYzdMur8YAsfBj137hAsgfYA0fLc0FfTSfMCuLHEQmXvtmhxOr7tVNVU7lE4w+uis2
5ZhG6Xw7A5B7ZzdG9OaETUtU0cHeY2DT1P+8lQ6siNDkFDSYIcFPQlFWXngtWMwZpq9qKF6IMIhw
PLoIDmOHX2EvE3ATZ1fj8ACB02MSJVlS7zRCHi7/VcT/nDufYCLaDu9ZAlvX0uEzNuP/FCu+tZRj
fMH6B2VTSsbuiDjvMivsKsYiaU71eIBcXummSTU5FMQVIJMeNghy2oDHg5zs9wMkU+M4leLbbEJ1
bSyeyWG8HsB6kbTtEIC2yVhkxeB+Wb8JwjcAsyZdO/mVCsps0DkebOQSzYnm/kE7WgRiUCn8/Fqh
6vCSnzwUWmLEVTjH682392EAEYbBLzaauI8LU4jZfCZRSY3iO29+bnjk3gq7zFP/wIBiD72dRjiY
vE/ztW7BcwkyqHbW4//J+J2t6k46mIetKim3+VfjL/wOuJFpHDkTP+M+og9rsQvwQBFYL18Q8c0v
a79d3tBSuCaiLEa0TAIac1JNfxo85b9v/I0vrjuXR5uTWIfbN8W0hRhky+PrE3X3JxhJo+l+Z0Lv
ykmj9DVVCNp6lomx4bZdmvZCJOidgcCOzQsYh6QIpzgkGFvsRc0ahzWRRgXb4DEjY9ioWLZLqtaO
AB0F5WNLBVyy5BOz9v/CZhf0pfbh2uysVL/+wnuFezt/1aZ0LA6b/wAj+aweu9Uz4w/aUCL+U5yV
YnBQ0ATKs18uuTGu+bjQtWf+OfWd/8lCX+Afc5BcmU8n/us8x/3YrYrsYzGYXSQuAIYkslyAjtrl
yuOQnNUneHOZvXfvY3/3L/rYXMLylwnjfdgMZ56LXBHbtDS+5k1WLxMphHn92dh9w3O+c7W0qsxC
TI9P8PaNgdyh7V0m8Oq3Ur0wvobH3l/FAx1lEYXUQmVAmPEd0cRtS8i7VFWAqzJhfk1/H3b+rR4N
FrHeWy6ofOaeqjinn3KqimCHUnA6PME7LXG+4DvZ0j/3ooC5gc13/w8CxnCwuz6jXeelFat1fRtq
6v6M79WTJOtOLIT2vQw7Sr4bXk1q+isTrHD1nYYe5h1BdC3cjLEnrbWcd3XIvKaJAN0j2qU8G1UP
UfwVTlEhl+ITHC+ypZxbYG5Klgz30h0GDYtFdQMqQhDQHAnpxpwcdR510URBd6TNjefObVgnxj3X
WlFvIYiEcRXKQVa5Tkj3IJUkGjXI3o8MUY7skf6FChZznbOT6ByqGLhhcXLitcn3F2hyDW88DpgK
+6zwc+80lUWi5sjaoYjxvlKGFxA2n185jyEsa6h2TSTG8GvUmKMnOwbiCEWdiPoV5hYDfzIv/Ig3
f2dUcE3th9HDsGrn7A3ZpyJWWqryXzVem00r3FbIkJ3hQomA0tbmrkJnvyZdNFPJUnPZ/4qbtJuf
y3QQ/TJK8GBhheEhL4iUxzSnfmaoYCbv0DLr7kuueAjEAy/i6IFE+viIDFNYfCs/YPPdsey+LEtu
yTqo1pvLxo957qP61brNXZl3FbfccwCcgfOT6f5qtT+TEY8q1eCPkrsTYOS60or3sWpaDntOxtZP
/6R7UNdDvXkjda0JzWMm0Jq8sSyG4Wa0lJpC0K7CpOXbO0LXyXMKs9V0spvy4qSUba2nmoAxDY+A
fP2aE/uge4LEG6eH23Xa10k7LVpOZcFKZEIhSJvy2S5ua5pRjvI20bKa3AZxH8CEkneQvo5XC7pM
EMJD8Kp1A6kVFff+14U8X2XKhvvmwaSJ1hq39LlF8CMYrHyb4+Csr1aTiR74MqZqZ3yRAF3rbhIX
9NNgCu5Qgz6f/SnMI86AYTA1CcO+Ez9S4d1FZ69vxoM6DQFBqmlbqTGni38GOR6xnDhDvaHn1kTE
M5vdZaVxSFfFbpQNo8Cs+TJrpUA8xf8knAiAdjqARsihhUuutmKN9gKiVe0FFqG5QnkE/40nw4W5
NRmkfI50rMg8KZSM+jJihCAx79NDGrzhXf4K7TgmnrYGJBo4WOPuuzMVx8VxDg6/3VlbJ6gO4baf
LoFebsdGX9MEEoV1krW7Vfg6SmF0WN0SWZjRvrF1lH69CsuY3u/6NnEED0D7lgFVEhK/3dyORXN5
cUZF8JIqHCqRNsU2lVgbT1MQgoOQ+3kZ4LHvtclSJJN7g2f0fhK1hrSP5jBGJxocz5XWWxuWdhqy
NK/HSYMhFBFT2E3fLheoc1sawhEniVww1CYiAdti9E2hKQ3ICebLNXw7qs11/Vc3UZHeBXqu/5mF
7xFNrGUo0YEgQN3exX9FEo32zgLDvngPerR+MmAQUBZ6zOaIX2uGu2iNKTjAHr6zsgVxbXnzm46Q
oD2c5+cW2SEhwKM8F8xzC9NAk7BiZUtY7GomDnK7EJpcG+0kBqoIbsb3Vu5AZXxnCSH6CFITyeGQ
3p1qHe9oOXRu6/SL4nBA+dFTligbyw8qMWOAmOXvC/DuDGELJPVXdtgrSoYuikDAq5AO3d2DKHsR
v+QCzX+Ctp1JEGgHOKf9izSxeZzMZSFKoSKW4Pp8UEqUbgJS/Tqx5nVYbXVQd9M3yWnD7RIVCpl3
lZWTesrcuS9Mbd3Km+AAe4iqWVSLjuRuy85S6IWpV0+BUx6nt3mRt28oFg7cGHZdIwzA5YhCX6AF
kKhjLab4JYI1udAplyiyNei5IcxLsn2+kgFMzHcQ1VCqaxZF6truvVjQdPCix8wEVk2xl1MjUZ2s
IxZVv54rWJEYrNSMJ4eD8rzxgsNgynYUBGd+KO0qDZuLH6efcjUpgwe97gbp9qCVhtP3rQ41Nb8l
h4R0CsAWk2iPf3YXOOeSkmX8m0SNnMi0+DuKS5rlTh2O2ItYxgg3vSJZSzafgi4Fh08sIKH2GMSf
bBYruRDGtoAJapvBYFMB2gAsN7LmWqwK8K3w82QpuyjlAcxYIjE9pKxfOCDHIwiF3InIW9iz1RNG
hu2Tc3IjEQGEaVb23dV+kzcermEvTeKbhcuVGGwui1+2coeTWqMmtgC84Ty41PBQnXem22/hT39c
mJ6wVQAiQuwXTrkNTFHKy3kSdCiTErJv84nlky75pmeuvZWdcQObgXkgkMF+3LaA9YPwLZfbN6Xu
8W+8PVgCJzGOLvAsnMmU3mRTRY5Zre/2ZXM5EsHzM/zUXkhymr+BbDRswU2O9lcrDTigzNL3d+Tp
l/HJjkpTAXt41Cq6u/jL+4kM6Jl0S39nqn8ynRe6qWxSKFTh+BpBQ9jW8M85+jcRXUPZixxAmFC/
CVq+XOOKPBYRMiZAKf/l4fRXtpWTiR8Gp/VSHgy1Y/7r5TiSy7fLJLn/QDO6Mhp2WB61VoacHBgu
DrCVWIQstH01vFPK7whTd2wHQyAxK82y6GOkbnC0DY74pXWBZA4ivXg4QhlpS02OGwVeOpEtORbh
B+d75O2nJYffrIx/TmzUZCfKk/jfD24bn4vSEvROPhfIZ+rk/2AnOfNg2sJuqimmVTbVc7yRHTX9
dVbTKiTBcuSo/wv7AdCXM5A6gujzs4sekdk1iodQ8PcAnjpdwAxuUpO1UGF+lAXBH9o0xeNMdE4y
dyMDGxc88VJV1NgL65ifAuGFZQgi6WuLr/OWiDgPUm9SErUU0YYRuD4ifBDTBWbKqHqiqytGbC6c
/5C7y+t2l7h20L0j0zzY2LEOEq5BLcbTGfWLQZc0YzsJGTn+xFf6WVS93kOYjQirzww0mJQHWkvz
0KOnKI7KWQ5R2uQM1myWWbzRFKF82LC4S8oF3GuCa67IL0ioGdzK086kylMMpJx6DUe03eP1vjxc
j5vWaK40/1597Zxk1pfPdvq9roSCrzaHXS+YFdC+RV0H1vZ0gbmZtSQK9u6/LiaHlivxn+DogKam
CwRKMnaRYolwjOQ6pY/n8oqTO6EusuPt0z9x4Mm3uDYOUnbMSHIX6oU0OuX2Cy4DFPqw2qlr/Pcf
VqEmbO1/BtIB8FtrgiZnj6aU8/0YD3drm1PhBqYwFzYIHITFRDmZFN21mF25bmpF9LvFA50ZzNqh
9T29/H+9cqX2owtQcqsVBwN6QRMEBT+ZKdORtrHH3ImPnoFdYlb4E5qer5GXWgvK+2e4rj1NyDQI
8wLG91N1vMirGKklyMODbhciUVTbRqEa/cYeWmY3y4RWU//M7pmn7s0zPH5Ypd0M3nX3/gR+m68z
N2jQSq5QtuxleBvuZrIbg/rxvMG6hmBmDegiblpYfEtvvdilq1ih1sKYtJBwHQJVUDEf1n8XDVZK
3CHq6OsJ70kqO9QERzMvEBCq+yEEjYHto2o4Hb5CcS+KKtxcPNFwNeUDiNLeOc9VYIo7bidz5u2t
tnPXwPsZCtI4HLGTC1WtdV5S+qnDqc3AagQSctzluDe1TozsRaAYfvykMCxZpi4MOs25M8ZmDJyb
g74eSV/M4+eE5RUAbYqOKX4cDLaMOa4XJrC6zSWn7+BLJjR0Bh6wCjbGjKfEYLS9XFtffnKYAd8B
xzVfn0frbC8jRW0iaUhR48HIbdc1BoopQqDO60C4aOE26qj/VfM5eq0qYHQg4xZiSf4mwoRs1FnE
oqNRxj7Lhn1++70Mm1Mke9vCjFq0EuirWmMufqCOoh0w1aFQO4NdZdkkAMSQypA7n5xc2Y7tcSqv
d8Howxxevsk5GqA1PKEJdcqXgYrqeLPY1Xq7OjMTfXoPJr+fOabnPcdW803Cmx14wCGaNoUSerjG
FHwZYt2L8YWNLOzuoN1yNvYMzk6vSSU7X41xxyDe5OXz7SMGsnR/IaeJyadZtKSTBlzvym9oRKU5
OzWtdCYiu2224XsmXH43cF0Fr6eG8ZbM+DMN3gWjpsplUAfjEzFf4dUXYS5KSWZSr0hGKsWkkuJ4
IT0OrH8Vu+iiGOKMJ6s0obMqiLtdcUID57VxYz99uVO6EoXwXKULWQX/FmFl5pVXhzZnNzGKtrqd
L9PUPnQK697bDcOtSYbp9S/YRGzo2FaDwLvsydkvfmSYfceoNpLX09wecwk9fWR2zpVIAh+MIIxi
/8CnrxlUM3WJdDPAtw9zV418wJdrX/DicyBDu9SNd+QWfoX0AR5Q8PdAkB4fy64YrgTp53yTMFyP
stvjPBJ6E7lqx0Zz0AirVAl1fhdxgKOm04nYxZUFAvwB2Nc+zxazRcpWa+gKDVlnxdOiX61q3Zs7
+fa6HEcyO1cBeceE8r1NFEz9YsrDOpgNWHBNTpan9Ud1vOQ86K51vgEsKFTbKt3hE778SknPNI/c
zB0iRow2Zq/ZWmJy7g+LT1bkwIfj1zCMVGNYL+LNa4YcjYDpGtCdGmvdN+mL7lPMDkJT6IGm7i5V
PTkbtL8568735JyMC7KozDkUklj+39ufvxQfhCEYCC6MPfelJRYNjVR/kyMhJZGWbCZRhomD/vil
J/h/AN9fJE+AWYcb9Vrctp7c2oaR7vDfKkSXlSnss6rsesdNiwOAlmNoZvQKwApy89Vg1Bot96bp
KbbG5wLMrRQ4hqG/e5TTC4v9t6RtdOoHUVYVgNPZ8f6dvQ84vztVbztE8eOLgRnTw1zMgwBUkPGB
zZs54CJ5dzXZE09H4fhspl8akiZloXuLRTadeCo2UE71dyaedg5WWVLowilLujvDV4bQHVJ2TbAY
7WDh/C0kSb0c9RGsJuwth6E5XDg222hCHLvRcjs4A3ojnOied0+uaADSLDrBGgPQkYpGpHxFeojG
XkufIiFt58yCucyU7pN6cP599rLaBxjkikoivsNZAOP43zq2Tw5mAaRlfON+NZovCzOU5iE/xfmW
ggqirbWf3LpyJYmR8LrAhadFuQ/iIGIEaYRehG0jmCnjHNARJGcAPrntV4lCfUFp+hUtFbtpdpId
WT9YV0WUs56T0oEgW0fulX5lceSd9+L74gsCuNnWwZWGyA9HacuJPMpcXJhrtEtBK3klMyUcMkLo
My+fsEuif3/i1fRVsYlQEWuFZqoGOHTFtgeBVSdSLAlzG3b9cxXXb+OV0+eJaUiq8XfeJs6r+/8A
CVMbsbTYFQd8b5uf8Lqk06D0+ZfCMBguaD30pLlHA/BsVc4DTK+kHquKXTCiB537d0FYKcHQWzDM
wnooxJWTrMXBOCqpnncXoFRYkVPrtG1wo5rZM6k/NCFloL0y0NWb57MZdsU3iyG15U0KkmKLApfe
xHE8alHs+1wLFOMtTFGwzpJsDp/uSMAQJyCcRGb9NkEzbPmhkUst3ealTL5lNWsDf0+hGub9HqeG
Nouc1Lp9zIiOdQVBR7JlUyB/24zbnI3qOu39C2mi4cQHH0+xBrzSxPwUZUB524qZCUBHvwNyMDAy
/Yfalol++rSksfC0I3mYpSYXGewF4BkETNDZUt0fhjT8FByMuqKS/mj6wHeS/U8NF3QVkbFlB1ZL
KZhWJJRuTj6U7R5BHUd7eGigGuPB7OuAdB3dGxhMtxIggDNwm0F4x+Z7PGb5viBuOXhm4tzgvs7p
xIwXmJLa7DdR8YfI3YGOjxWtYndB4j5rwFPb40A2pIZ1NrTQQxpMHlsNFseonSorNwHFF/7xDopn
XzuWS8weiCsprNoVV0iTKbUtZ0Ghlt0n25BRtLFv9e02lV/Vm3jCE2Z2/n/U23hkXomN8YX04/E4
3PhYlDxavduZx9YJHerkPyy0nJWTGgWWUS1v5dmWlKgSQ8sr6r4DJWnFNaYcMXnHGSf7TZLrxINQ
w8gpYcn3p3ptQwhoVQKqZou1dxSmcin7o91j5OivsSkoDie9BM4pjuqohTUyPj75f8rccdkmFE0Z
cLJjwSvqlVHdotD2sz/bNvVhJy01lvL7Vx6+AgtmP/uqSJn9E8V7SzSKpxUR5r+rZhe5hUtvNku/
HEkzx3uCEX9FnOF9jYqDIOUAXBAmoLmaVKCUaKrk3SRl4vrnsk7rY0hHSlg9LGZG4ZLenLk1xCHs
Wi0KxmyhazXkGn5eMg7ibO51S4tu9muKbs2XrDoJGc9uMkdB8uWCWZW+6AOrUQ2pU5Gg5tXcuZn9
BONdPOEUCosTi/kpl7clQXBQ9IwojxU8CMG2IVrzr8Vf1NmsRFc6stGDJZFTgOMiBWTX5VS+dr6C
e+IJAv9fWIlT+A6hrLNj9eZr3qT/fKFZiLds1L0ZI2O0ZmGQHurbTiunUOg4RfBUNFsqC0vBMdYJ
c3L812zDTYup5Gm0ICLQd9i2iVt9OIsBvY3z7x3MKKgKMZjRsIN40wB8E9FxcLhnfsEcumnhazHG
BIwncUQBmUrz4Xdjse260n5B1ulIluQQlRspoUYxI5MOZnSDjcaBPT2Gjp99TdP0yKTtAVqZHOL7
Id8rzJKtsMxiN3yOOxBGyAuF9qPLyxiW1I8JwkBuQhAL2CN+4tqD9/dEyTHfIyugLMQbvIt8zbnv
h6JGpbFv8aGng1snjffFwyY96bWeKjIs8LH6YZCO1h7T/BVrZyVzGJuiILQYzt4uklTXpZ0byGSy
BACgc3s+d7T4HQnw4TTj+M7c+OpjDEPjcDTYW9KBl55ocn4awNcGX9YGmTRB1REAp6PWEvOtV98M
qc/ehIa09RORLmM8MtD2k+RIWCioM95bFV++Iuh11q0dn92JugqbzjqXB7BCKDO3umNTBYt/Y4/Z
NRt2z6IjIGe4Q89z1jDjHaNKmFaLiPVHWRn5AIwNczfQqGxRv4qppZAsVKsDGKrDyUteTQM6Vc/j
KoD4AN7IzQ+7bGZW3niAlYg8OLehzOqq5Up/007cpaLQ7327WC/t0NojDfRbfl0txZyXFRzHPMRW
yz1S0vYkU9pC51AsDdNRHsQgFXuCObIi7wh4E+fDamETcgeG8vUf84fm/wrasMldncQpbTEOKd+M
xzQI0f4HWgzXzxtBCzAaZrlqishStEHMsdpXDaaZqN7/tiZ18f0YyUCJdKazpu5lpMExE9reANMI
B+Va1EqHiFh2fHkFtmUxRkXfrt59l04CdI7NJuOtq7exrh6w0QJuyvqorTp/GMXQnD9Fu2wT7xKA
ikYnwS5wcET9g18CpAgV9l/TX5MWI/6yOtQZJ0TncuMedfZhIYkuJqAWEG/NFymOAdTCTK5XiT/0
FEH0xTt/z6E+X2DXQ046mmyjiFhBcXDg+fz39/JOUhbR5SMMjKaERN44IM808LxaDbWqQq2AJ61X
i9NZ85CZZxoh/UxY7EML3Ax7AWw+Nt87WOl71XELQLyMQfwSXh//OthnMwwvzVkDNKQS4kO7N4oh
EI9416HVNGgA66hBfrged2bzDlYdUPhClWIetPshlnGxDcSLdvqP1NPqrCjZwdA+8WwuusobsNg2
CCUlgeP5MCWLk3TlZaC39X9KYf/TtGQSJfGrL0LmBsROn2VkFrl+2Mi9WR0uw8y5B8qS0KCbRHDh
PKOkDsUucG86iACbloaVsqoommKDDu7MePyhnbq4gTuO9kAtvlKvnU49mnvYMNhW7WkAltB5gaVP
Sz6jwo6qa5qfKD5kvmp2HVEkiA74ZQuZzMWn+8Dhea32
`protect end_protected
