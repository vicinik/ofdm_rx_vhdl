-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ic5O73kjIR/FuPwmxXjYbk6JVMGXEz8p7B1tWc99rGoChIUR2MppvY9Fkutsf6X7GoDP/LKtjwmX
dVo6l2i7kMCShb4HR14m9OCgBJKUsF3Jf4fAxf1eDpoY+9Zbxlv20rhvWZ0d4mR25GQEyJMgRNj2
DxeqZ3a48ZtpKXDfps7lN5x/JcxTJHZpidn7AZx/0hFrSa8fAuCggfQhiH/B8uXbIl8aN1TchKq9
ZgvPlSKjfM+tK4ShDaFAmS8PO3R1Ygzhw9tckRswWKjFRtnd3ia/BUHXirck4cs6R5S1KXUu679d
/whnMEBYMCFgw6b+W+Wny3h62p4qv0d7vrAuzQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30528)
`protect data_block
0mBJ5v1XbPf3qZhL9mVSSLmAJtHi1mQZxnxwc3GNkiaBdjZBeSR4u7N4jZ5A/i4rnsLTVOQ46FpQ
zTjzGJopezBejt5GEdBJmfhkMvfAxostc89l0moQVgC6u4B3nt4QC5qQV2Iy/boWIOolLN48I213
WNKnLt/7dXbNsTAiEkzu8exMXiYSAUGF7rf3uJGlCVXqrKpi5fUiyxX0vy4HXGTuumiKLAwNCsQs
ZMBvA+xVegcutGoKgXx64v2h493disqnV+G/X8Du1c05UfiJmYmqvrykTLczIzPPKwohXYobrv+0
A9oqewLLgNBSas+naYUlGO7V7VnuePNTD/bfGNGGeF/DSWNQtpT7Ag45Nvtnvj0bF5UUkV5BJ3vC
7JyTrp74aLcPQJ481zJCZE8o7drwrFc8WXF557iUnFv9rXTl+INcsLCu9vkh3tZ/ExLWjhwIrpwX
/0J4rDcC5l8It37FXM90oj0FPl5z1NbPZrtKwt4An6VZHArFzNJlJUTRdPlyd+ZbRNyO5d6pD9KD
sW8rIzOFyqg5scygWXB+Ir8nNGMxiTFvNVA4ePI3OboN63A2Xd5YSPAQr22aZJKjqtuHc9zC6OeM
780KmXvAZLSq7lXElHS5uCA3E32YTS+oVevxVkLmd+fELAmvYJmGLf4L5mKmMwDDLXsQsoptF5y1
gk720OVVzsefqY1/Z6PqRwvF4dPQZeYhoLq+NXQEW25MxnHECGoYWWKHviDsSGZ0t7wxiYQHYQmC
WiGIH6lfayM/YNcCK8BgZjmyNxcLTVVh4Z3gDy1vm7sF2NMTAQmxeqEhkW+k0fBgJvN93b8Y8oko
JU2gT3SmlgkeLLdkBB4rb7HjEgHH71/oqayhBTttkvoY2ff2eKx5kdlCZ7YnUuwLOOzPot6XsNU5
JSo8YpYvEbhHdjeO6/UVjIlyaxVcDW0N1UzLs3UOLPDxwBCs+5ZSWf89NVFJC2SZUGK8mxmwtIMn
0zoRl/yu6b3o0vbm8iSkdAn5pXBCWXdvmpT6ydWE1SsJTfNXqN2FD57dWBLfh/KN5H4CRmRunFF1
1eXHGiFc6GQB1GAkO0JXxelIzRiUHq0P873JEjpuD64JtfpDsFdBtUBwWnBK0wh0/q3HQBTM2/a+
r8+6bN1UVxDQg1L7GdgeYoyKJF9cpKkAx0T78u49GL5jOHUmqGDVKurWI2cZETxENCcvrfLHCKFX
mXMRll/noD8wCZAk3fWDgHgpThMp1Q+O0ymy5VWzesKy922WBsSncT0cKJctSwpNDWuc+7YQ57p5
ULKe7XtsIJ53C57ZxRANsHw7FbH7zvGwh8CnP6XbGWZSbQPh+TbPoMvPq/Ov+mCL4G0rKi3o+fRP
tScVb0PEj4iTMqAxdYO27ua9pz4lIPiqrxuVrBsuoQr+ozsoUvZ5AcYu8q/dhVa2nrfMe6IM4FXm
eA/VXNNf5gC22fqLKqnhdSc5ezjmID/pp1b7aGRwnSV6T9hKzFcNn/bnwlqUEy73hyAu+fcrkg6u
EOqZk42tXHF8nYWlczuZkFAvXtJhA5Axu7NIk3Qa9ghph3f4kTsNFMCjlhnz46Ju/zWbrzrjtnEC
2lwOm/a1bO+FgaSZvYFjU8CqvZ+0mZ5kXViKKXvSaytMDyD1p6kyVRCJNQ/ZI5ZoWNhp/5W2P1DJ
30RmYKKfGknRSVvR+6Hf/f1JnAUYVnqW+/surslRfLnMPMqoIOUzQxx0+cM8OmWhRYZ2moSqSQOh
LzLwJF4+kbrnekerGKydqrYF3ksF1tzWF6QSb/tMlDvjfZyyBiCVAj8bKJ75Xl71GmAruiD3qTja
AiXhYApFXt4gQTJyvt+2Ohcqau25pz8MkpKpMlqNFB+CnH9HtUzUo2I/hm1BoQ5LHMCYY+G4iiZd
nP7jSiJJDBtK1Ea7WiatMf7pR+GljVKwkln7iDH+2RYqjq5o6Kj6zuVd9beaO04StUGobScCnrvW
iHRfOvzjeq5YJd+3N0sGUrHbM2rKxx8bMmjXS5c2z/4Azn1urYpgC2VEqT45miZNSNk8DRlJFgkE
JMj3tOqXsFVqv2GUEtQU0WvAS6lGysp4CxXAma+tMA6RDH+MHSlOwTUq1GLmEGWk/KbUEwOpxauL
tI5vhgkpLXUMzYho8WTkZWavL0fPBzxXQl4DEkcxlXjWi8S8L1E2ObuR8ysUdPxtzy/tKkWqjS29
PiImwD1yXaeHuHVCQQKZZJvYWkAHHVJ8UIOmzRdCvrE6G4nlEIzxHagdqcwNn704BaLwQ/WTVAtU
ONBTNG6zJphvR6LLz2CBGM45YvCT/a4Gz8oRQLIsIoRTgcpNZ6KH6df67C9bxTnAPHJmXZ/fg4wO
9FYxzSDrEhScjZnqcorOqKU86TTwlZeID25WwoQWv23FII14mZkePwcUajSeAt3zY4IKudsadBO/
5bJBt/gMCs8AsdTbu1eEKioh/S2/Nu7+YjM2BNaSag5xpoluAPAWqeWEGAISxI5ec8redwNXvdjE
5BF+/378HD9Vz93gHdD84tc2EEU9V/WRzBOoaBf4RVBUBqUzgxO0EBO/mNUdfU/W76htw2u77Ity
m0OimCSROIDjkbNumuwL6JABnN3tsTA2koANPVB6rcwMO5ssqNR0WHrT03ekTj74E4uZ8EmHlO/1
yr2vwbg+JcSdPb3ilKur9bx60df7wl1LqW5+y7V8BI5fRHVFW9JyH+X9oWjyJqR0mdgmxkRgK43/
5w31tgtiRjDV1esV/tC5TCg1VdzWxNvQN858xqCg/iLLS7Gi+z0l+klDUB+V2KwffIJ6Wx6l2Wnw
rKVngUe/ljxNP5RjjtbPAzZp6/gC4Vz5SozPmQYcWCEg18QD7Q8SRrV0RhQtVV/bbNBEYpI7LbAz
uWVn9fRB1J+tks0UaXRDlQfoauTJ+s3pS/RaAcfVsaRoAUm/BSytmV1npsy6SYv44EbySl4xnj+M
M5LSwXuk9eKb0dkys/Qy88ahZKzgnViBtJtD4qnTfanHNsfpU68v3mpuk8a3QzjwifZMe0mAr2G2
99DvpXO2eizaV0yu3lpmdlzFt2g2oYiHvrDpb9r7plCRXnTEDSrRXVp9FYfyQbml2Yc0idzLuNLl
ZIleKo4E33b13p/Rbyl+zSn9LR/HI+fU6tK0dfMYe6bCyYt2mQeftj2PHY6FzUVg+dk5FLg5CDK8
JcEWX6h9Lv9KoKIZfPFffhQDTycqNP0iINxTxV7NY6+g9zra+vrloxYfrpuYnLxCQiYgnFG2tQ38
3d5opt5wEO88dJU2QY02q6aNbPe/A4V/6d4KTeI4AybZXkAFKKF6i6sw3rdEQT/3v7BknxKPM3SB
3Ljb1zj37YhYYcqhSTfKuCJBdgOxYjpkgJeipU6eljkHInTOCCtrnMg6amR0d2TT8CbSu48TEJa3
QsYmXI5L5hpO7rRimGupTC9CgT0BqLGyoeIiUnwSTYGLZw/FCejFFQCOROmhm75xYdFDPjbehQ7o
Rc35T/YCOI5SqTIGTVbCtU93OJ/IRA6vyELeMdzPBGx4hpk45SXY0/49hG5jS7NE0t30JA6VT/xq
QhNZX3nbq/ox3FCeRCxOYzA/6EwxrJrdE6IXnHu59LbvbIx6SFJmlkK9MfgqtcQ0XdO6TJT1HNOb
MEqfk0mnh1m1EvX4LIFXjUrwYW50GBlrlm0SB/0HBJtXjSQIXapKh0mJprtmxVJ7Oo0uggHSYVs1
Lvyyu9BgNyGIS96mxvyCg/NmthrEKfGdhTbMGgcAdHvmQ6TwfzzO69sPIYmq8+AWP+5+fL+oL6Sp
7WKZqfge4/jKXEEONFbWc8KYNIRCwc9+5iiVHDTjKgrYdQ3Nlbt7QS1fPdqRUQYlXDbqIbZcs5oJ
IWzNihCc7wuN9M8EYuih+a0wTrVTUaI4o3SCL16QgX+wRm/YtAstGeq8frNxuM46fWjqV5vOdTlR
uAegMFDF9cwLVC5OCs+l0k2RTKbk8DqOh093Std3LD84fbwfmdoEjJia1ZG2mk/k2QbrpZwO2Bas
NYEhaHawWk01B0FOsQkLg/ErmHfGFN9hSN08yP0na9CLaC7UE7kQqwsVWjl4U/012E6lgspj/ojP
Aksyo7zoLcK5VSYDWPTJE0srbSqrgkJ88cNRPHRgRnkM5zZM7yior9MjA3xfChKE703V/5vdRVyW
nsHmtB9hLVP99JcyavJ66nedMI2kQAghVumMXUXLWuhgeLF4GH9edob3i2QhLFjV+pI391FvQqBE
BTWKOtNglVa2B0EQTea575FiUREREQhesPJNroLSSZRdE319c1q7C3DNwZ8xjDgGiONhVMlpoGhk
z3jVLBvEitxIRfrog8c3bipP4kLKm6U8hmbcOMmHsJ7aZIyyR3CfU9SLHTMQSPGU2mBouTo6Rkfa
NWGnik4jrUuXRXalNlN6XmGKQcvoNIJQu2F0Exzdd2o9I8VWVTybAOnC1eYg5HP0qAX8T51B9evo
7odc0xxIcD6lDHnC9vDkgPtDMCaXnrAEkNu2i5GiAE0eBkYz9sT5CioSF0cNH8lLK02Hb0Im++Te
K3UnhTVZ633M0xBN0EmRJ31hcA9nqrhRYUue/FjNAHSBbHToS2cqKS5SwcgSTD9mTEC6FcdEu76O
KwJKfxw/WODIIyxyQdGWUqVrQH8cE4RpvqzbDPTgfGxs37iggT+a+bNedEiRbp2cx7UPFC7cdyuW
yJdz2F7nZVxNL3cbw4WZhpA7C0yI1SixZerWPLfE/qRYRJlgt5nux/frHjAIX9s0JNC6pPmvth2s
EjM5nRjpufoOtmqrHuZb5rnbyamT05HHL/XIqYijJIiyvUbQd//jocf2PVqt6krGuHlH1twEwbM8
F1mwr5nsZwGVAoYh552O5P3WVto+ZD2Wi/ju1+yBzBt0XvSoX3ZcZgCrYEUs0i337s5gzFxRaKbG
awi30lOXG8kpCvDYAHTtoLo95xxAtF5zS2mI4CY/MjdI29gVXjgUPonYe70osQ2lnD0ITwhqZnKI
Smtl8qRzSLMlVIOHY1WjvUD2amiUyD3BlSbQpPOpdCg6oKC+k9lghV6sRo8Tu1SXWhIpW8nZ6/Le
mnvBOfzA1ashcPc6U0Gv/wKIYosbLFyVMYFY8546dKFhIKUK3p0q+Guz466lZ57RbclSoo2he0Tg
a6X/UzkAjhrA6V8VKyFxNUOdsLZmQnknZgtZm5aLO9rMIVBarDWu66dliWo0KcBSvKmUJdWxuyk4
QKwHMXNsyYf128mxpCzmReyoLWKrKb2V1hcc1SC3IjljzYqQKqVgoZpgp2odQhOd0ilzrdFy5FLq
+uU9by/+BeFMZLNxBzp667mh1CKHZBI4zmYhAeDeAOCs4maNcDbplcCZgg7FacwQVohcEl4slAI/
UBUfrZbW/zzzNJ+vkPrInRFlgucRAwC/2khT9UU4d7CENwgLWW9keEPX+s4pdRz4NR1PxJFu6xEX
P4xWfSlIuXwn1Sr9rDMNj5s1BlW5md5cGey+42vY81aGqICXRnduDcdniEvBhVyrpQicbHOkoWPu
GP1Y4tg+QHWaVNWVpCrfIV13w0IpBw2cTFzBmNMOwSwpW5xK9XHu9Y/AdFd0wUZW5L7ultbDGYO0
CWrHIXyQjk7ApB3CdqMj9pXqG85GH0zeOixb7Z7ZZf/TZph6nts98jU7rDnys8xJHMlqj9wBU0Ty
d33T803GsL1LMOQCJ3IeHiDO1HBtTgQBXiS1uuuNKEOj8zQR+u4JxA18GXLpOixSfsVc5EtYwTKd
qcFS/NKO7sK8IeVECAvwxX9k0NSUkUF3i5zhhWlje0wq6ChXO4vzVVVzc+2Uii+OGQscqNh1asRn
cZbBxnoJIVU3bq8O+uD2/8uvYnQS3Pu0iBkGZYWaqiMk9Xlj1DBa2HPGiyhJPPem0lOZrLmiWWRL
Gl4eO0OHf+XK8W7l3QaBW3iixKq3bNXjqDmHXosoy0NwYQYNdwQDi8VfWgWT/u1HsQhCLZNxGiUc
ZcoiuOXJO9tFLaCRTyf8EftPcvuwQNHL+C3ZaLkkoi0MbaJDPlM8mP4106K9j4fIkjQUalJvo8aW
yw99jHLkfJWgvH/0kX/XwSSR7DapnPC845ccSHGaU5fL2PTWSFQqNElGK+YIhRcAtzV4NyhRHVqc
CWoDgdhuF6EAqm40nsYGScaud4r+GgbCBHLRw73E1fQZeMvbSmc4stUCslvbaKxFBezqeWX/pRrK
3rcMcafdjwy12ONj7/o4napUrTBZ8M7apWlmTGwO4HH92qmhHcxF2VdPojRFZb+c7mvm8hg/XbHz
MjqpwyDXlR/i8kBHCVz06suTnzt0ELqm0vH5NRKFaVRJLfpq/ZFml7eca7Bf7qrq/qWALNaEPutS
ijJvj5EoAna6RY491aJpBgaG5LVBgWmTPsFCkdaO42eH02HpCQfhLAbTudsqLQHqjw4dkodQGmC8
R6pFNj8EM967bfycuF2W5Q6OriZBevwOGyF1Y58RvaVFXbJQo/o1o0xAnOBqBUc6/ltiZ8HTj1v9
9G/JwcVtNFZOsBMqR+7s7/Y26v4JcT182/eti0RfXDjo4AdoeB09CoSyBDP8ndhjllXm7jQM02Je
Lvu5Xn3k3wTtdnre3lpOJKpYqiXkreJTFYd86mY0bAnJt4c1eB7w7a3Wc8hmnCWnDuwZY/FnqxVr
J+S4iUFS2s7DBqvjus9YkvnNdrmdeIIuUMyvAdaCYjyk6sb7OMv2Kh4xTiiGlGiJAwOaWN30BuNc
RaERXKABo5zGQCHlXagzBUNGplgCI+qqDIkDeqWGqBcl2/D7+tQFN7dqiqkf5HcKbPu9nAL9NKky
qqwq24ahCsHRC45f3wH0ZE2lTXeoA2q+oxBd8ALuRYTj2PaYzLQkVqeKWVVwJHTptL8zy7Yw7NUM
uL/9x32UdY9XAmAf2sbx15sastzGM4aMkFyRpOepKGfCaxpFK47RKWsBrCDSst27VXbJEN6Hce94
BKmp/W9gGgCxWhW8WR7kbd6GdfSRL/Tk4WGRQz8M+jXmNc7OOFLg5pkbrsJkQOmZ6vGIQANHt0NV
dELNz233zEmtTBDzjzYR30iSX3stqP0n+jaXnVJdnboq3Ip9x9d8adzqOhssxLFAPjEfi7Lz4Ytj
dILuyO1KIbaIzrY2YFEPPHNDfHzjlLs3k/N2qb9z/3nhIR6C7wGx+I4X5aJrPs83IMxeLrJp8+Uk
Fx5IObLRv3qwrK32i/M/DlckOvn+2QDCpEhkXuouHEVFk5P3GtUdjl350DFS3cjAFKr+wSTglDo2
1GmKwmcMEgzMEUxSCQlgaLFqCGbfeJOwVqJXO5xZDFAJWD+sGeWbprsY2ZLJzG1gMSNymDW+SMXa
XvegF1wQ58pVFx9WubD7VJ5de72Mgx+9POqFOVttiNW1gKoF3aPFPC9lof8ceXjVJdi4UyE2l2Ub
XIgILceAxm50EhDf3cvl0XBXTFxF5mi2vLyj4A+PSgXKSMJKoA3h1PBbPbfU5oS3I+GUU6B/fcyr
sKdl7Sa0sus140552DjJAy1LH13nW2lkoZ/AyeV+fDoKgkKOeFuAji+1swZH6H9PEECMXVbP1fO7
MYDZTy7cu35gGbYgfP7FxnoSCG98oGBbfLxIj9VYEbLOMeieDJM8jfi+mW6n1oQ1A66n4mGRuNBq
PWcoaSaquKLJ8gE8DLaGb7YGXbRuwZpqvtZOZnorRN1I6BpSrXfzexC2jYF611wd4+yLfEHCK3do
gmpqfkGx1CCPLmUFCwBCo0BuUnel4nPU+d83PB34tpdbJNAfm8jWZ79ae3pFDszKX/DtPN7Ig6Qa
IoMOaNkncIghR9+DMMMcE5P/HTqEZGi5ZEHnQz3JSbJ5w3zuhSxBjo+93Tgmx8+RSOWegYjQ4vfl
DWOKYQ56sXdYyj5TeP6zS8VSAU9aBaLNCUD6X1/t5lM9xAoUhA9soaPq4E9Q5vLtEJVs3t/dIdXa
w9kMB+zcy/d06kxU28Y9SN/yRxxrUvaZuoDv8uwDiT6gVxITycjLy/4WesK8ehDR6d/CE4+6o96U
hz8UCXr6NSHiYd1hM8yDy2joCjP08et1LvHFzbS8DYSRTC74sFlqY6834WvFyJlc76BPTH5k5yQe
UsTDJnyL8NSs637FCyTOGT0qPxhRnCFkT60OCbqaRsSQhA/7cJ1q2y6WBA4XAL+YunzBxFs51XZC
OFVX9O3wJpWYiGaj/371EcKZfzPKO2metW7NrcaBj/bJA6gYVbjCOIoX9aZzB/onGU1rNhHICslh
j1t9XjeazijY/4S2p4hV+klA0nQp8mdS2hRbIaqIVTYvBBbK32Sduyj/m6RdjEraeoSx9ZnC7vNe
mPkne1MgkCS+x+7ZG8aIoZL9Xv8f1xCaSuPZ3iYPts9ywNZV2REF2hwEb6tOZ1Kq6ZuQKtZRcR5+
sPgYrEAbW/NDaWGfx6YRymadz/Zac8VsXXYd7FIqR2RQDT62m3HlqXvMpigLgJYK4Ea9yzEz1Kuh
+ud5hud0ey0bLbYLoDdcMBQsKwg4yZAa+6Vc7Cf5OHPJUUj5fw8ca4qfRq8j3pJNWO+qrYpWBLgk
vjx8OmENtQJKbQqb6t1MvxJz9xFlIEYjUdRX48tuT1kjTYdNR3c/diwEiX4AOl3OZTn2sWhmz84D
W+YtZgylaEKZPFGxc7ioThbqWg/3ttZUZxjsZt3Ead54MoUBBP+daC1birBkDfl3LfSuYxKrJHVu
u/gR9k30cXINLn1XjgExT0TGWXI0fAmOOJwb7dvzJLDePrY+tkvJoTiIfovxr2KFg0ZF/skICN1h
d/P4e6Fn49MIbTH0GozzgTdckPVwu9yCOBYt3n5gHVvmtrXDY0z8zaNgEEIUALhcF1RaD2QbCOJM
CU7LBsrjiXjzIaWDImwIz34rCxAM0MxDHvjXANYKKETMCtmgcKJZOP5iSyjE+0mq49IfM+ZKYvVV
UPakVqPxFqPtlhXlrtsWOvWcdC3sJJTbbYc2JtXmFe2a4XcFKG/lkHtXEHFuq42zw5Ws+ihcf/jB
qoWYkPRFGAqSMvQt2Cuhx9jbwzVDA/l/Pqwcy40rmzTvV9QpUkRJ9PJxcCivZq5KvyJInHnrtczv
f3wtpEKiQsK0zEZ+gfCFGCJM0j6ywIN2TMDpENQXU2nF7VZ9N77S/9yUGJ5QKYKy0YosLu+D1YNZ
28HShse1zvAN3GAhrFwz81LGvAZFdY9dbXLI9rGIov3/mGuwsUh9yHIoe69Cfgb7nZ2K2mShzSzq
kkyc9ForlVJU2dgJpL7UaimiQw5TdNx5cCkP5VQhhIytcyCiuQGhgrmI05koomdDhtdDzPzl6laF
n8gylVMIqiPaC5ymr/Oqkp2UXecDJtbCJWXw58wHmAEot9b9LWSNgizBYkDY6rgGKDDQrESF7X6c
d8zlYmFViY8t8jSskyvVMdwPgg4PuouKgJMpVWpcvZboIZqj4uJnubHXn9B0H4nbNuB/6y2LOAmx
Lk18HEm1M2yuI/wAHqIWz2g1a7jltqAEfbUCfUM9wukCDPlVZvaLQMvTpyoVc2MopNhGyoVGueJC
98TQJDXFwtiSp7SGjWEKvN/Z/iroYv2HOUIJ47fLSe8m6V5MN1Ng4AxLG70UELXDEnRblw5hhqcb
82zw6YnULz6C/97DnXnHnLY+HztykN23UxT/5/lW3Q/BYGHsLbf66AvoZX+0ua6ufX/kAaC5ltZl
TXGVqFu8nyo7u3ozdWaAqgfONZ4u475z2kVkxlAyNtzqWIXrVAtNj3wirdoP/mA19yeefsvHke6Q
uny4KQ+T4PQIyMgEGqR/c9xi86iXmOkoTOVDYDdsUKYPch1qd4f3TFia+ZX8Sj0d6CZPyDnmxj+h
jE6I4LXPmOssyIVLQjEX7S+abdD04eHEaNRgX2eESEJjp2flFBQYRub6u9yitkj81TyvpaDp8zT8
a2XyGoReAda/XcVEo7iFXzu1dVtlhBrRNaCA5ns1T980EPTlsWkocmSgE7BcfWODwKMGt3QB/ayg
i0cVQPB+PfruQxkgKGsFFMAD+FAmugMr67SF3cPGdfG9m+kPbB7sdfRrFtzUWUezvjIJCAH3avB0
TRco0FSH/tJxbYMvlOtB6z8I7T7Sk5VFs5Nzoc7fxtMBzwtPZxjv7DyDmQcm2lKu7P8p3jo8sJvg
lR4JU5+zWucbIYdjOVLscc1ilWJ73ub1hnsV/TTi5WubRWXN/7eKx8BRS/CwdR5BV+Q+qQxhxcic
knOz41K8U3+OJCoBw7cd513TsoknTVrcB3CTUcaIap/5O0Ih/poaemrwebpqbqhZRSPATFiUoxQC
Wr2UXQccDTuT8PWoLTU0VzvrMoEOT08obK11WcdoD0KlDBV+D3ZrWEMdazzPgjo33ZGZ+HLwCFEn
emIeNuzhLBDpuGCPepoCZMimyU+5GQAoADSk/0h/PU9MHkFI7/wZAxNYBQRGKAgXt5h9WndhQW+U
iGBt767yCATH4FdzWBGZ1YezMkiEP1uRmvzbknHj1I5ACZ9SGqshdrBmfCaufAjz0Ew+hlW29EIJ
DuIQJay+3EeTUCxMn7BXySoqLSl+xAl/n3YhIuinvqQF1DgY3DWqeLdN+qKJ9HvCcoRTi0h8P1ST
pQJwnDPvakNEkewrWc3+4uRAgC93MtBBZ1HjQu/FAaMe9yA4Ti7aTQHzEMi5lFKJXbqUhFfJOIRR
PzB2CebF8KpuLti0nf7rkrL1xnO/wJc9PS6K9IYsiH6r+WkRfVHrYTJ1+vPAfiQxsdDvIfkcDGhV
iz0DDOprj9ueL8hQSUfQO9fDELA4H1DwCAC0+hoSrmEwuh7542dt0MPO0vzqBMuoEyBMMlgLxwSW
jGCTTyLPmQiPhf1OCdGdDqQt3+2FOy/1li8Gx4CXQZc9UWhvcctn4JvepPKtZM+GhsIy+6YIkzT0
e+8yt4550JKo0hvm9UNlG3nuAoo/WBvNgHBnqD9UgqUNzzoJcBgj6ALG+l6DfJIfbVW+5jNuvcbM
DJ+WSiYd35Ndi6uDPEtQ9Ba7/GcY/Py/A6U6es0BwLelLiqXbmyQGgQjUp+fvAdSCI5+3bGZhPNM
IoCT9sz+IyRU9XT3+P4E01G6Tlc+zsn7OzUWZpTHQUu6H2DiE2tlkcGEjREVv1xN+MRE12EGB9oo
zKU5vjXhBW7odASddzJbWrwkXC1dXIrVTn3ITx2adf/ecR7ZVub/oz9wNcmbOjB2DlSPWpZettHe
IWqYRpevidCAbi3b7LOegyPHBv7NggWQbPKchqRi1NYMSP37Rto4QFUuOJg2BgEVhI4cVkyCgwWr
37wTlqAShKHzHSvqP+kq6DEInbjsHUwnSGskw1xlkVxSggzqbu+T1KHn0f8eJGKLdH/ljlofVJM3
JnIVKSjIPgtdhC4RWQ+6JKNaWLNMzaUl2kJkIS9pgNWLNgsj4atKffiS4qb0xo8UhIAh96mF4x0+
zIywYjd0wTlX3rF0+Om6d2IC3l0lxrJ055dpM9DpfcDoPddYPjAkDatDjqBrWdo8pXrZnJS57Gh/
Lji+BvE+eH6IQKchvRQLUINtr0GK6ViIVBNOrgk8uD3XDaIIDoF9ZgzdSvGXIGcb25YZp10FTs2F
7qN1Cc2NFStMGJB732ZWqgrK7+KkI1oK7fEhEyHDOFc+w+38leo5RCLaL18tK7/Y5Ab63Brygrg7
kb/POl2uThE/ts7YbBjcxlcpP5wOInF4Q2Sy46/WfcW9jMx6/2L2fLaTml+M8CEEU/tFZ/MDs+qB
MuOSrQ3f6wmQLoWWgDWp5amR6T27r3FM/gEtSqr1DTCnCERo1DXaZjZWT0sfyGETkk7YpStsXsrU
ZB6IkryZX+rrJ0ZW06xOPaxHvQAbKLoVoeGw4o9y6+QBT7AJMogizpFu+OnbbRhUtfIneHY+oqoD
IGcaak08vTlQZF3wCanHn3cykfi+Nw6EzGxJeFic3gPIbBmtN5XL2/2V2yqTh18ZIOyLQVRPPuQC
t+TVp+XdOHCcmw4cbBmGB6QlWtRF2x/NHphCWQbbXyQTG+alNHcQUyUdPkg52J2G6lxHRZ4Z7LDA
YMY3cyolmKhI03ubOb3ZpxiYS1HMA/OvaV16oKTU2TYnwL3yOe/VHFkg7oSpUIMcMb8xw7zJOg3P
eVQGZvr+VOv1OtfzZrDkKHHDfpVHeQakZu1qFDnqDAbEaWK9fH+XhB+RP7d2i8qP6niX19Ub2gqd
/uhInB4oY4rEbLogfr0lIBjZYhb4ULJs48/TKD1HwwQiR5Y7SwYG4hm9azy+kbXVTsIcMNDriv+v
CoLaQncpsoRJWFmKLYlGl5Wyds8R5kDV6ysJ/JX9xIz8GdEYZ9eWBy9A9GYA/c7iAPmz5weJEye9
8vn38eInxzZ0YdWqxl887UwuwVHt5t9CrMAt35xI/WXzPnTmSMBQ4Ky7cE33rCrDG1mRZ5YgqqT4
+vNIa5bLNOWLS8S42D02+N1R6meMiuLMVkigF7SKb4r76V4zgloJYcT7Opb4719y5VYNovSvn07a
wPBUV/3mhO3M9NH5lOsPbq1wMDNkRckfNmSoYLi4aIe5jxIv8YhvrlwLWUURR355mw0jBWJFDx2s
/5wJoueqglYzJ5WaTFNOo1dfRoVvK/+3bvBMPARH6Jigm29OvjdlB3Ip7Rjuun8IT5F3D/9ji3Rt
g009QiEB6tTlhlhJbi811LmvgI8qr0XaCuyardMKh1mnuo0PNc2crohrmCTzMS0CnFLP2sM8lYtf
pUbArKuZkF5bZUkFoCDucAzO6o6CBs60fyHVFGqwTgXwwTDZryfih9OnrYTDdxtpvv6OHnqSKjmA
rNpwQ5m2ZX/GmvZ1EzqkYAIiO6e206KcUqscCr0y0XM6nvHauHga5jiZuIxqKpYfXPovPM4Yn/QM
aoLywDn3r47PG2aezoyBCP9jd9lGU9aY9lgLeGHHItJAz92x8WDH8kwZ+/sx6p0kJeSlQTuIOVZQ
oz+wpP/Qdpb5gZM5SKjtc4UxLS6xN3xPzJcQlfLtxUwFFVyclBpzVQFbr9V/go9b8FtMB3M2VAta
2bqjFx4SLXNzKiNwNYIVTl0A4HYWFm8xqojohX9Hokkdb6Q14qOSYatbtTCL3FxbR4SkPgjfu0Lr
vHZ7Swjp5qxyaTDAUQ2QVSMWEsMLb52c+sKUCvh8rVDk0fTIyEtvsIKJJFD6vbFu/4E2TkNBuGDe
mONFaaZgiMwEHG8hq1wmZIwWwGi+HsT6PuXwp7rAf2JipOwuVLYbw9zLu34pMD2g409dlTe+SEYi
wlfEd+vQ1NevmMIOepjPPnIyeg9KspjlxWKyPufMQoFAUgx5xbrBKWUc0/juAYjcbdf6f2T+cFvA
yJULBEmOZpa7euFYG4KdCaRTKkrPtkuUgRHU9dTNOoWFlukqI7GRZ+B32hTI0OLVXqVog5QBK1nV
vdydb2/EXRgfXdXqlLhMJIMUK+aR4+mgzDrrggqKfVJg1HEb5/fk7C6BlDIVJEAn5nkhqYW+Hxay
Ua8pTlvGBXEUghREDkALqRp6uYqWFKCfqGN+N39tqLFMWVUy68G5mrftrFcxA1+iiu+DdslDZbSS
xb0nROOGQkxe8Aft0XccKXUIvcXVzbacg7vkLx9vdQO9WazlbZUc2fx1/a/AikRmUfxMR9gKDj39
b6gYml5qapNDmlqrXVtzB2HlbMLoctj3AYlSuCChSp8HyC+qynmpLbWODp0Wx0yQ56c+Mw4Llapi
YSpbFoVsUujKBgDgFxRdfh77YPKopoxfngkeNSqUrxEsfoPLO3dyJ6QliUz6SqgKEtPy6sLvVGnr
CmfX6cyNqKfXnGK0O6Vgp1wgBefJepSFoMj7fkJqbyo+S8Etq1EZyd2Eb1Q6z7N3astEB2UIPqXv
JXiClP1/9rdxHJZC8Ht/+BMFn2nMgwv5Y0I2bnZhB4Rth9ZJV7Fx2wfaQDe29NW9ahWtcKAY+kfK
9JSMJet9uaJDRMvhxO7Kr7hrg0Qkw0Q7WYgvVPKCvFAEUFNsfwALiEpVtXlq7VVxWp8gtfQpbqal
vzwmHmrCq6f05lbQ6M9tdpgSNeip18CdT74OTTz2a9OBbI0zH842UUqs9Yr6M05nwKvoiX92X6Vk
yBCXiLYXmNiqvBN5LFPR+gIR5b5ALl42v9pc5Yd20POKyke75FEbXM1d7rOHgvVhgKETK5tAQDtx
7XoYjJt6IEBG/NuQLwwuaxUtRTiEDGoGUHPbmkyWCTDA+2U/YtXwg/7CIoQp5YXMWC0+2vRZ78Lc
Zp8S1nKRyL0Dz1pdDw4TR0FwwlogU+BdWFIKkXvSEe9x5fiUlyCAqy0CPKjm9Wr5re4JEOAXhy6Z
KH+tUrbdAH9njRaIBhkCqx2OB7gKry+b9s2LJbZI3/8HFalPR1/TliFREtgFAOQDgWFoVBmSJRJR
rTgaMZ79j+/+dtNLuau0Iaj4/EzdAABhPNjpfqLTJqpoSDFt2gB7Vz1gskI5ZTAhR2XwshwmvaCR
iTRYMY3VOQvm02no1KzkF0BkP7y5eD9TIxwEYomAFm+b8l2McscjyXZaF+Iv4mwdg818OAS1/d+/
jBlh7bB4nUNhYBV/v2sMYVXtH9ikCxqA3R/8c2lGXPGlCuK+HMMTUBCzivOSVSI1yavzP3Fua+Fv
PT8aIRvl4ZEwvouj9ec2JWU0Zcf2ErWSyw8x78MhYMqw+RSs5C+pqbJ4Qz0r4NySvROSDlBwNudK
OY7MlcIwdPi0eNEHrxUKGAIF1TL2LTmejEylhfv7OcYtPCs+2O8/4s5PtSHccZMehEzp3yn0AFlJ
fBTdRJ0zypJZb8qnS7u39nMlIputHSk8PyjFYbai6eDmScIMxn9J5PkG4aUMev6iIPm80F9R0OdM
TEm7ES+TRKs6E/fysJbkuBv8n6ueLy++v385eRMsuCX0YwiIZK9ARqMeGTc/bnAhl0u/nQGXScex
M5hMWjt9yaoeW26+Fhko9cCHwWedsqQI6lmMG7V2IEs4bDe/Xmn8VmXmDdNuApm/rxSyxwr1HQsM
bkco05qxACtj/EV+Gwon+xHit0wtnJusO8tFZ3Ey4X3CogvSWeCNJmVMATiTAopIQkum+9BUMF9s
gLsWtGyoJuogNvXoaJUSxURY9bB6/tul5F5pdnqQ0MgfT/FeUjPUTC+axDBufF/QcA9r+AQkbyoY
ApP3hhUU+AE1Q5hSWILcl9/eIdPdIeW6fQ6/lV0iI6JroxMKIvt+vwiHqebndgUlutWPn9cqGuJ9
29BF1D3sVQLBiG0GtzaG3LLLZF89GGR/9PilPITWLT/SJXefA9rehCCSXMiVhfYNBusSrsLs0nnW
GysIrQjO7d4Cyry5NMSluQ9SMhwoL2YaYyIFDzD8NUPcMOFaZgSlDhQZNVuyQV2Ei/UV0JLAteh1
buPPEjyi86/OMvpqDh+ZjZvJDYhFO5Yp1SZtZ2oAY7dgwQQ4exIoyJLFzWUnr1oNQloP+46ZF9hW
SE1AARV5uRg4B9F18vksgR/HQhWjWL8rSgnKEVd9B88tHbfOozWOFfuMWihbFA4tQJtVdUIBGiU0
IsJrrvNmpD3mgES5HWayCHfMfdQbFFX46HI6XmDnMvBQ8yxTyaUk3Zlf7v0k0O/h9JsUSIznwOeU
RSJeaS4nO6qlhz0D4oat24q832MqS3sZKtsUhKMzLqHzkIQHLDwT3hyqp3TXjhkw24QI9Xi4t8ZG
YtrMsqRzImb3LMz8ZWzloyH82OM7tDThQbAPpj9w50SRWH7oVT+IBxLEt0k7oUYN2m1zJSZp9WFF
fsW75EhvBnpnSiaTCRFi2BiHsxEPc76T+oFrmfYiSw3tWDpE9nYQQE579uSoxHy5VCI3YQQMiokj
/KwXbDbFY4s9/JJms+yJR/hLgJ8Wbui1wfwGKeT9r3wfONsHb2cMYFYWsGzn6nei+zSXNLCWV1cv
ccXXewNEbrjHgAJwHtPwJrxbcSDmsV8i9rJKORh8f3MofWCdSi8Z6QlBml75VfZZBkP4B4wzbyJ7
ocetutOj08k91ujeX8zE5KKGIXpai4IL8b+XtJk4cjIf8WNzeCQ+fo5aDAfaqRUqGpUXcn9XVB5f
9joRY9hgn8nDHGg6NAhcE/jiVpIw0QreGGxjllTh/i+GfBkOarUIlUlm/cKABsCyoFki2++GtDLA
1eeJiozVom66vhVcvo+rqeL5+dAl/6YhbDr+YQ7Hp1As7rQXIIo1gqXYYm05yIVzDjKgEIRMj6WD
mqMER9F2HVnEaBbk2eAC7xwOqJWrZBPR/ri08fHEDhbD4mbsW3Va1v3mtgJpHdTaT3k4AhlYt0va
gn3S/EaHHh5UB+JMjoXufOg5UInavah1pM2Rb0Q7lGyYerafnSD564Y0m4g9p/Our0cX6evbL1mU
w8rREbReX6820GSolHqdOyQ0qPdwMXw/tNYi4+lbyAv9S6DaCwCeCV/2yQzG4WiHxX+1lMNPqQZh
MTR7KxzrTXdgipsX9YgD6pv0/NOyRqKoeZZkYZjkvR4274pI8gbizp79O4Y71oqLjohjJr9FeWDY
MLauARVuM3UBMdFikGTO81CgsS8AlcXRhtt4LxmmoDANyU4kiCzgU6UOdbJ1sSmJ5hhrLpcyM4V0
6Iii3W6pf089s/84q7GqGWECuwFsH29LxREHqPnx+wpW6qaOv/oZFMax1a7hRPU43f1JkV7zm0Dw
7L1XccCzaIjNU7vSu0e98VQKAE/Yrchn3Z82yyQ+YaRMVK3VfhxpmQbeXEbEBg+OmHGrLI364xeG
K+NjL9nWPUIt4+lLY0/aHRCBQfKoICwc+IbKZN+aKNbsXRZpipAgQij5DkHzBD3wC0tTPMEvJuY/
m94jlPqk1Fu0GBdlBjRCRBD3qfMAUPkVn5d4/Ci295ZIklvN3KB6vIGpcAFcYsTxA0K3kzVR5/i3
XlPJRPh1bXEczCzH2n23ggvw+ALGoYYgXgA/o3FbxkXw1b2L7KufuHuhvnEpoclh8/yFLedn3Iu2
t6kleEOV6fRkfTYDAEEVAD9kHRWvoHAxxq4QDbkB7A0UNg06dEQisKmAcoJY6PcWW+jQI0b2orVg
v8UYAMhdQcVY2+jHfzHlhU+O/WDnBFbJ/T4+IIhpIEh+CIO04vAakbh3txz4lTdaivSvJLFcP+8Q
Bnfaqmf/R1gVWlXAO+zLxkcDwPY/RnVAXgX0osD/z5KX08JlryRT+r8jMF3nbPl8oegSctcMBLO+
tdtpAW+awK5fgnqSqU7DDz0CyTvQP1WUiUHve13RzETKr0MdRZ3E8xpC76TEzHe70Sq4s5MG3KA/
OFUszpKY5XRGu4PKsU4P7Q8bkesAmq3LIO41C0gfe66wbxxK+8cteAGVyJOPh0solF23yC54Hx6T
Amiv49q8Oj2kb4F2CqaPnKtsU35Sd1KAE8MO3xFMWMugsLIXjej6pFIakxW0DbFxsHBI/0yzHedm
fJp/q3w6GhV4usFV1Ni0BunjCOsAdfoX6TlDz59/A/wkygl3YxkuiDJCZXHVUwNxKhkA5PffacJK
XV4bSgCbklJ+WhIH2CyaT6nBb3qO8ZoatqGWqsduHgymyiPjebjQpteY7hD2re/nAt/czJPUdEEX
uZ4BVAAwXZ3Vi8ibK077TKq0t9hmbSHHT38SVhzajNF/0EIJdiQlcxVXvmy1xvFA6SK2AE0lqLnt
IMGwq0LrrN60DV4cIgKHYYCMZmC9SzWeiVzz5lwBLBT91rufFFvcvSiV8OM3EvKQNChfNyAg45+C
eforgKi4fRLD8yMI3Iz+6oEMDDkUY56rpJA3Z4KftU3VBWYoLTq/aXbJDYzDKfy0JLviHNNyirRf
tpBUNsGZ4BQT1iDX4e8cXVFIHIAkXZxFFAqYQNUtv/ZsR0k2CCJ9YUhMwOKAfuYj/M08Xm7u3hc3
JH4NG1SSnOwhLQ1/IWiswzSc1WJqiixR6buL/B2D+QkV+dRoHmB6Yii6xbVno08OO2gFVVs0iUAw
3R5u4xt0brWUVqomArDvsZMsHa/5j47PkzRemz1UVm0YUK+H9myyZj2p2CFgFRA0nALC59q3VhI1
Fc+6+yUi7iTfxikxtL9y0EElpheVaWzDsrmcp3YcFiYOD93+83jF+y2NY/fw+VAwSNxWp5uXh0cG
JwHlbECyFitmp86ZhU8DybL3/byI317VfNSOKn4mKUL2MPr7mMDClbVHHc3ov4f4VCVzORyJt68L
JxG8IpV8qQQP5k5ysqZDzZnbLcEBfFKiu89JCa9naHTi8EOvpPONy89B1OfSZ6dxhD8QlYD+o+R5
JyL4sLrr0GldkIchSNe7PQ316rk9yRXZYiYn+mEMsbhvxqYznJZaTroLSQr3weDSsWIuaETZSX0i
UqlbjVFJ+wWvCT7MsERHia2oJLIrmZ2+gRyM6fA6luoh1tqqlCCqOUxRNsaJ646LTZdSwdUd7jof
rWxjJ/3UwIMlf7y+ALYdvYSUJaGQuQO+VlnTLI8Y5/p10mtHf6CsF9u1oYTM5wbrkw6cxCw3TbsJ
WCVigNagzm8WPyebyTo3G9AD3Fx83DhqluhTCnB9klEx6llzWd+vz9oN+Epv/JrAfXax6dsaApe5
7bSwI6L9GHkkipMze4yEq3tLkdgsARvjFAayfDH4Wznj2dsUpMLbxQ9oe4vJZLUh1qHL0nvo3XK+
f8iXjZlonIckwiGC5DfO1krqVQdxm6rpTJT05RElgF+nmoFLHmNsGnr6Z+mrRRVAhlNnqj2d5Qo+
uZ9ltBw+mGR4WHPCCpwAsXI/FxQOZZi0f17tdBJu0mhYm2JPGRFQxyze3t+Lau7FVddMrkoVJylh
RL5uQGr7HzWS7PqBXtPTKWq9MuNcDWJ5fgm4la2rDx/7yzWp0KRFhSM/hBLvB/BWe8zSDCTr9SUD
dbIb8cYp2NhihfcsKryW/nC0u2EyoIRZQN1hdwRlDSK8JVkvDgo2Va3K0lryNtd4ArL7v+1tEPWo
v+3p5lGhJe3kmBHRR6E95XjxWXrLgQA/MSAPS3jJQHHtGcP4LP6uhvC3V/qOQoKUfGHPysvSeq33
RovyPhbpgqxS02H6BHYKxZRA9ApvK4DaQ9yV40ZCnN+5ZOkkxFfGyKy56o0NpLRA+1EUsMwGSQjF
geq4Zn/DvVzRyKUDdrvRQoD3hPGUzmomcJOiYLEeuNGd/YWBv/4LzbFe2EPzAwGRlSanA9zBR6BL
WNo08Uy9/P3TesuwHovCjWtz6ru8PxOhQ/egV9SidgbzWcRkQDOBT8afRYa62vSfsB83qFJEHHJZ
LRYPyJpcxIyaAaWDICP3pX0i064SsKjMPJ4kbRHeJ4GUQ4P3vrB9vHN9y4QadRv4VUSJjqROV7uT
67xTngfTQU219fvbjM0I5ez9STRiw3AhwmllC3fwr1DMKEvqEzUYolDgm/IKyyM7l02ev6/sfsDo
uU7LciKkZOG4rvvPXylSirTp5m4JEXyXQWHG8XC13RBOOXzEQNqnMN+tUmppqAYDo1S5kZqIZXp+
5UfhH4ZkKCu+lr5au8rByDnCjf0jZZPYVeOa156msmdmdILaiBzEh1hlijlunBY2qsocdeXgX2Bp
CQ+N8LbjpmhryqYLU4b9TRuVLsgW93yJGk4ZMjsGBzTXXpANoI2Ns+Z70oVEbZFAXJHk58NtI8JF
nV/65mJnWQsV06sLp328gD+smI0DWnApBqjM5Fv35usSGp4THkeALXsmTmn5FPOv88p5ZlJB0cJX
aUrcL3iOy66bvgjwXsw2VKuPM0PdfHDw7A+lwxQu3OUqJV7QK5RWg0ZMSJ6HLUlKm/XEG1ZSTkUR
tISiDQx2+Lo+TwxhdGzZEEAxqGcNdACfTTxtB65zKK308IsA921mD642iCXNCcBgNhgQLGhwiZhm
kbvVqX7BayDhOiXqtUErn/Rfy/qdj/0vp510XsLsmC8W61yNeSymfdWj6fa8eMjL8pePwAdcSBC1
LEg2DvVzmqG5evUKWdM2KbV9Hl1oIRxwMYcYloXgQvYDxNAmfRMaSRauZNBHLcKqxjksN958HeiW
WOdmvgQ8olqB1RR0Y/T8AUAz4Ifmvj/RlG/JiRptAsLeAsdrAcISouoHougK0DnlZNwuLTbqyF61
JQpm5wtXHPETwix7Y95Hb8/fD8ULx8WF7Ex+FIboEQ3ry/hn0i7a2urQ//qBuaADv/X9SZ6Bsqyh
IQ9JzRF4Pva04GmbsPJWi7trf1Q8adrNFvJiPtJ3WLUJ+zuQlotLMktoLtnlgsx1eWtpbuIByWlW
Ebj9a6YYer15vYX2GvqsHLaQZghL8Vu+8E+RvCRQfV03tliwpKgW7j6Jd9hgmHTn+waX+hnVzfgG
9mVog1q0kcLZ/pOZkHsd74z0VReQjtyB644UlCdi6zjqL5YMm5j7yeYFELuXV3Hkopvyoj31sXdw
dPyUjxzB3VLg5of04NITydd/oTD/9hLuqBY4X+zdV7UP2Ojxgt7SHFhqNQw1c61uY7NgLZz+sbpa
s5pNB/eo6bsB5oiaVwczsEs6V+9eP/obmcEZzv+Tn7NXEY6Kl9zxUZUsj0Ia5jUjVxqsIU4ZzSUp
uLYCUgs8irfJp+eq53Hp+2i8h7pKlTv2JeAS8YpeQd7K/XJBjTdr7/tWyGK56ldTGepo6/9pHgb9
5Iu9PXoTPeV8UV764rbim7KuT8YsR/0cUt1QWWf/EWypFAiEYRgMVazyi9nqgHQ3RGponQG6z5wK
ZkVyqknEH5l14hmQf7W04wKJ+XD+VRyV7YFguNUUxDIwVh7MLnEMo4mewllwnQpXogvbcakgj/Ah
nWltPfzgSeKP0tfH9z646SaR9Qz16nzPwNCOCFP0DqdajXgprJSHnyX9PlYfyGIK9TxDZzmo+wFx
2TIHVPOjSDhAlAqOulE8QjtWLIWhtrZIQ39b8PJRnO/C0ulPyO3gkDjQeh3WumM+/rPh1EDAc3bP
1t1WkPn5QU8C/CPnCmkAFH1YrzNVWqQ3+SFS9lQ+E8YSNKFPrZSNChZupGCeNifTp4PUouz2ke6R
HDhoY3MUQ77k4aHQWe6zyRzwMKq9ZiRLuNenl+z6B/mDctid1j2Jo21ZRVGW4Nf5HszdewRvXEIz
m+MNetkCYTGIQUI0t7mDaqAn4Eyq64iRIFsIGnliiekoDMZsPRR6fyHeJ3QVt0oJfYMlvpbJ9wc/
SLhUnOInT3LmAZ9Wkkl/9fGxtaJ8nyyz25Qba3FEaCVhwRZfYxYgOWC7J4biIF5NeMXDCSIsFU99
B8Ep77sduGMMIrfa6JAJuQ6aawfmbEPUDGweSIOUCyvo/356p6zwQ87gaB/ga+NGsb1BOLJO2Rq0
FqWizsY8GfQMCtr5fTq+QEdzi9uiec4zP/7rTJbSNHQU0N0CSoLX16CPCky/qwPof9kldShMd7CX
i5NA/tp1LSyJ4rXn9tn9gdWEWFDNVYyo9RG51+umh7iovseoV3g5LXtrcaAqOXacOirkW//VXUCc
DPAkiwXkTJJW18rY//+7LD2FSMDzuOI2adWzPxxPC9iXNFepxOzxayHX/OnxBkKNXbFFyfKUeCFd
/cMw1erC6NDWg1ce50qRxASnEwXR6pJK/KQXf3iTOqia00uIB6ZoRrxGvPd1/EmEZmh9rRhmHc/A
GFgIjyB6j/Xhw+AfQtNQTm9YO/AIzfCqLglnPx/CQpecORTURAFbptziHt+zh2dElXeG2hp+KKzA
/JNgPo8BHVRYHEG8/x1dK3fQ2KNUDO3Hj0UjTjhgqa6ThjGMUmeJIIQeHLZcggA37as1yvahgJFs
P+qJu1bQOnwTykY006iiJ0UsOPxoYAxJcaiuZZuDRRtoJ8FSRP94wE4Tk4wN/OIUD6+hL0IVJWyF
WvzlcN7W2PEuBJv20QmdKTzIsZ5PVD0ZcIG2Mv00PQB86+4dTQWcNHZcxMdhay0WWxLn1ms2AjU1
jnY63kN+90nqhldaIqjSTxV6DdrzEdHSVvd2NF3x+GK9+fKX/QpFKVrm9kqbV25mxh458ALHEsxd
779kWREV+zFBw0NjSVW54yaAIeLD+ggM9QNy19wkWsSYitvAVSJsVPtfcnIHIB1uygnM0omjk5Ye
IIhhgTwBBo77B8cbFxclK3oUGouY6TZA3IderWyjZAAkcTnpzzH3r0T581+K4F0Y0M3W6Q5sEciq
32fOCF3w1rSUmFya+3hQMgUKbQ8f+gJnhI3P3NhWz9VJAWZMBkKUgRJusI+InjIAY7PPeQTMiAdB
+DOAWSaqdXkar5Bq4TiE+dMLNFdqyAcIkVZHMGM0VJujFurFPAkqDesbOzAmNRXU+gci8lcZ21jO
JmBGV8dIuNPEM2J89otb2YuReeJrwk1UMcTUF17o7VtJm/orkEo0ugWoCRkSXn3I/0zoiw9WfxOa
2r0vRV64Me2I4t6voLKGVRypRDMecI+RtoVolsYY7ex3DpN0lClDrYIqK8kkGMGmW/AyD7bDle+u
02eUSPZgbeDobCSkg4jqSOvBGyPWMIRg8arhK9pQODJofZIn8qZzKOAp8okVIXbNl6cFphweLJna
OQvGZiqY/tdL9HYyWxV5RlWexiaDv8qBdIJxi3ellFLsbKYNNFzgukTnuwBcpXvvjEUrmHLHpmLL
MzpwX1lx+n34IctuwDR9Lodo0J7j43arFTKzIxYxxF9WhSHb2dQHWcIA4XrLHXvxUcTRZipUcLBa
t9igKbGKffj6dFRh3+AAVmodRn8POUjW2cGiPhy8pWoDf3WfpEQYgviIB25gQGqtme6yc3yRt5Jl
MLMAYUqc+2aPwl5U9V5kKXX1RJEwP/L7JCnmntMXgTtL0kJy/betW0V24i/umww9+zL2qKz5B93T
W4EB83yf7V5qoJWEEQJlvEj18mTtmEkOig+HeJcpG5aqE9xlIxT3ir5xPb4kFJDIfgmRtTwk8xzQ
9Uau/IS1ojbAIgNRdFooQeMF9hwP26GQFQX3+n0rDGo2I/Y7a5hM8imhbOpc7IJ4t7aE1yMGpw6A
UgCCJopRnEEAFDX44H/r8YWn+k66ewh7dJvzwmUIJ2f40HEEswA/wdhwmX7TE4opiuxTIYI5j35G
IzLaHRXVDLHS2ZLhiG1E+tnn3uuTR3O6kl0gjQTWPeG2KEwFVsoEyvKQ1/zL22wLcEr7jZ1YWqj0
Vsfv07ezbVS0dyLgR8TOMYlPALD1N7gBsBMaTzR8OdVrC/ffj1KlHXlBg15cp6TobaAJCLQtGnkk
qB8yIJqqSFjfgI9vpAxTt8msjmZ0bKp5TRCVAaod3PN6NNP/DqnpN8OHO2h6R02sIvMd2+/8JpYf
v4HGs2swO0Iwu+iF9E22bHACZiA+0Jym6KSjmII7XsNSNBbQwqbqGIqnBuB3QUDQ54ixjU4jZzbL
EECr84IGbHE8NeedmjCyzMhK3xJqRez5xcBUigRxMZrGXgnNNLrQ0Y2DNaG6GnqxVshuEBPGeVdw
9yHQ9KcJJQLqvvLG+SJNBona7XsHLam7BGOfJ2onaUxY87CN7dWtJYx+q+Pgu5gf8F3e4veQTaCY
Cyd/hQEPKRAqoTnqL1Yx365AApfx2Mfw5ehdYrtIxyjCWFqI0pzeI+D/5x7vKwHBzQZJ7u5e3uUS
fUGmoauGzzwz35VbVnmIUtq3J4Kn+5CNqn0DesUykDYsdZwvJeSd9DiIyanFZoY/snwFU5HV3dPj
5ZSTVDwWdk/xj11AbQaVGOb//6FrXCO4Eu1NuX4EiQePs8HiEx1hd4dg3Wph1C3HO6H88bo+ZpLr
0z2O67P8/MHlQku5tofUMTELj4KIUBKjdx73g6qzZEJXDmuNUPHLApjSVT7/WGV0Ibb69sAUZgmo
opopNS+AF7NZutTMtXOZMR9TehsUjtYK22FeSRX3MtK/S7qyGxx4f4g3HNkeZ2UJiZpKQCZ2qhwS
kh59lpuPU/y3JmoahssXLzUv7sOy21IIkuJ6H9+QNsrl3+QwpdfgL1B0u2bgdyGlxQgVitVTY2Em
zMUkBKQ89av3ZjrLEvSNrOMlW3T+fmFIKKKwngQ6C/x1Xg52jvY35Jp1v4cn1nFKbTKMlmx+ZmkY
VQSuqopZfVeGtba7Rq5w16JrifkY4UKI2o79mazgG/rdTaDRJ+KYZotMhziCPhtS1oglu/FHzucN
6eq8dHGQFcDh8h92K4tDbVsrri7Gb89bhVhuKdGaVnp2ORi0uUvUnv5dAAIK7vytic1ta9LL43zE
KlwWU3yJ4UvbjJSXsfwmQ5qEkgpSo+n2LLkj16aRehuP8UFQ+H1MCvdLGKUqgXRV87AQgCadZIoW
XFHHuP/up+fty0HvE2t+syJisf4h0tS9qWa3rEpDUlP0Rifnpb52ng9Fg4i0uynvDzucG31xhkV+
rVpAgna5ItbZ0f/GtTaYUzxbDo8TOU9osu68s2E08lTFUGVhbStVsBYCl+WkldLr1CC2mWkG5X6s
vQmMuBTMLw/8AVArTAdgn5U7tMtKRLW9bvQeNyJ3ltYFvQ6rbtbgjpwM1EUix0Y8nJxQcAXqtqED
CcQeJ1xyP6RLiDrj2zicqGZHyuItaLLFJf3fdTgkfgGHPqw0VxIKb+DyplubPZaMfYlizkdmqPG9
iTuQ6P9ERqbe7zsNgOz624dyobzN+0CIh5/YvuFh2RfpDwWSr179cAR51hIa8RyGp2PsSw/+7oAo
KyXVUrk5GwkHu2By0jiTi+wONqoR9u+i0VjEWiX12rb7SPqmJRnktwS91Vy5a3VuUfaQsOqs4rtz
O7TV94exyqyrAn+D6Fb6Ol7gWH9liUzhDOE9aBma8mieToyOxOzK5JLwdHm9YZ5mizb2/kJP91/C
V2qmzu7PLCTuy1o5Q1HkkKTxUAselPZA4RGXuk5fMsVjwssrRRgIIowjVk0FyQ9hDzn8J0yNGW3q
/eHKnu12S89pH1SW0MKFTLhXlyOLrcqGKrZGBEVQzpajJfcrn7uZlx9QDy8gJ8anLnqIUfCzw5jx
fVcxghrJs0Ld4+5fOYoA5cCsG34btxSrNe9dVtUo5e4hdLoZKb76cmt4X5FRh20LyTAT/ojLXAD5
ci40i2Xshs70COeMm2StRLH4fS6jsk2nb7uRlbub/HdmX7D4ZctG9pK/gkPaM715kH2tXmC8LIzb
MpAx5Rjn9GV99JdqJxQXjMt80ute1Tf9AtXWw1XI854vUe16J94+nGspgqmbAfQjlP9RkC6LXpkR
MsyO6NBUBj9NPO4C7cKHa15Wkwl9Bu2IfYHgNkRJT/qQMXZwZEL3g2nEVyOrWIiJj85yCdmf8xiQ
ukFRBnq/91Ix5pJiwgocO71YrTdsgBtHfYStEdu3fGpSmnRb9SaEP6QuWjhXM0UENOFQaLfp5bVQ
JnQNVF+d30tk5Ltu6mE0xiedD2hbw9slKughnaKvnIsWBLx9QoFdx8kSYyXg3Hdsks/p4/ZkoRxf
rA/UvDVOLhkG7a4cROfwS40x7RGRBWn0Wj7NUCAfOLX0BO+SRGfxt6hagkLg3r1FVS5vajqMMWzW
T3LfiY9r4uweIseBvQQK3Dtw7fjYB1ZAy1SX4FxTYXPrD3YqSmeec1bLXWuPQezmOO5mrk0VrO4e
ztkuyhP8SzTbFpg+61sLsgK+o+vAiNvTcFKrmB4APbzeegbHbrLLj0INIkYgQqtEKiT5TYN9OlnH
h781tjetnTnwWiDrJef3WsFVJGeYTxRbg3azKo502E1kXuPh6q8Zu1CbWcv8krKWxHVvDB2fFze7
UecZwWVEyQ+9LUjL0Nt2Y+cjZETBaDvIDDbM+FELSmetjhEc+5/kFV+lKHz+GAoaVajpxov9Iwac
JCkRxFTDgJg5tPWN7XzNDuhnkULhgLK9N27UJOMY4xeKUPC0UINhglHuqPXb7Ba2fSVvmEDNIAy3
msw7pumb2DiIhkf2mHRoxdRePNPqMZC2UO7HSRNiaDzcOnX3CDq9Z6brvJvpSP4VuCBjtpYaHl5k
q2X8RXw1+CSOh7fpFlqHbwgArHXwmEoNKMW9jJbNC/F7ge6eY+pj2UqFW4GxV/C2c31UQ0E1xQgq
8V7/jCF26eLKxxubcOLHd/cKxE/9dAeqn5DvNCsYAxL87ip6dMSoyhq5FB5OmDxzhOU6CEeBZHIl
FMLK1gUAYAk4bCCpvRdPQk78wQWZtRmBIZ2pi+KH+m/xkaH1J/BRkgKeFeHH7lSjSnrZ9B9DFZvi
iSee/wa/6BwU4az2k/EahV7KyUFGy6iWvCYUet6ubxsJrGa7pAQzo/1dqW1lsGkCawTLsuJHXYHt
jRE+reW7tXSaOmQzFLSpPbKcEclFMn2Rl/ml4wTKa+fRELwg5sZSFeXxXYX6VglXUNSlUCUDJ7vB
ejde1LONsaiMpJy+cwkzkxozm7RUjuyrkrX+jFNy9uGGfMd0Avn5Fs85A3uZspZ/7i18bUrGOQdF
uF4lTjrFGE94RD551J39q6JGXFhkx4UUVzEYS8z6IKy/VBnRIPCNgT3TX1VgIMQ2BuxaDgEAmshV
W3zaw3q0LoolNBWsp8rqPtV0n1yupWVAlodLY1oe21LN70mPZntxUQw4IHYd9MxKMxJ+LdjWnSxW
jJMC71ZEJ5OhHJZrYMlkEqII1vL8x5Ntss+thXdGqobR/JtAiul4JUFFdH/eLYXxMaSDqRK3gcxb
2FVpRiiOjG8imZiwng6BroaRSihkKwJzNZgRanL4Jax3Q8DW0Qb0P3v0RKBAue4SarCHPeh5QknI
MDGowammRjxoxb0Pob33Me9Mc9bXlvD/AiTTQLOCULO5vRJgpoGDcZkQDI3cMoeNGPYd+mwmuXEb
+Ivbr7ZLl2o3qLzIxt9efUPGmZg29wHaWLMg6vC189crojacZv6x62l5TVtuj0iyZh1qJOfyiw51
GRNw17dsIbzYlCj2g7nhKPbzxvpOw/DCe7REulFJpWzSxYQRmx7kkvYmpKF/b8AfIwdOBI16QHlr
t2xr2UJyTwAloIBDL2TSRUhx8/5tRo0aLfr9fDb/dil9KuvtJ5QpIcg8FOf2X+MjicZ40O5gVa/H
LuVhWaYoa+/V4Mu+TDNzLR6SiYv7x3pvdXbOed7HcmdQcdxwlKPSPJ6cOxUUcHAsGl3ne1b3ygoC
9vJOhBuT0oLiYfrwfu4yT8KxOyXbSXZ7wcoYaaAUUHHgUdCoene4F4Q3C8spUrg5ymeBxVqoqFOo
IPnseOWG4flFCD+wdxLK1PyMpo2NNZayTo9OmgTeZV8KXkGFOWkv4YVVDSA8Z08DaCnzUxAKYwCx
Noh0uTP+NCkX2Cdafz23uCLc69Ao2HOQdDcEbOkP717CapOJ7Yyy65pfnGn2EEBzPvvIplPgr/1b
ESwrmV5LWnU/unLc2YXA0lR54I4xhyzXwQlY6TT9yxs0jXR/P2qCXxXKod24pu5JVJboYiiyVqjy
n1so1TrsO5TpOmXCDG2Uy43DU0Ib4zYNtu3LH8YDTzwKw7imlfPhFJB8i/1YKT5qGCsOOWA3DqWP
oTvzG3EmsoJwhNJAMbGAjsI5wirv98NtBfBzBcEexczsPTUlxAYbEOTB5RbDkqIoo2S3bT8U1WVO
O5S3dYTaqAVAecfP+bOjh/LKFMiQN2RheGxIdseeX+mXS24Aidf09XeUr0KY9m8vUCW29zc6ZSNX
W0HAapUgVeT3PDieDie+SEVTvPUpJjIjhBjydTRo0hQ4s03Nyi4HndJtWlkqZTvmhMetmd5UhKRA
VxvO7O0ItgJ9JrqoqunljZdOakVUL3J1KL01syoSXqiXIamcRSHPQV89kyQ3XYvxd/F1e+LBacI5
MCaVLr4IlGRZ3xevcm67yM3WNAn0s5WG4FyU45Oo9GOsWMYcXmzB4xRH2X6GTXUaOyBSdhHFe7v8
VyYKmZlmCj2hmYEzYvxQ6CXoZQ6GbpYu9q6eP58+o5HhDagw8RxduQ8HJq5A2HN171dezIlPMH+L
E1SxVnm74BOoBavpN4SgugEbVQJCAQcylZMZW8H9h9P79WP466OfBf+S71J9/RJH8TJLdXSMPI0N
0wFgSdrGdnfAaohE9GLkdNvTGXOxQlA0x2JaTFIBNbsfxLHpCXFu9tH0f9jMknzs5IjvVaElGsYV
x7RQi0jjhwtYM6h6lEocY3itEpdECq7kb5ap6yNGKcgMxKE5n5A8c1NJrbT9syFzoUv82muTDtCT
8WYKrXTJInZXPX7pE8PWnIwhq/x8kecRjLG43QjGj5rmnOAm+WtGoO2Il/8m5U+tbnxp19W1Jxy7
w1TMMC4/zSVJpYMDnMgLNO2NIHFF+xIPwuKuigGFLm5a/QJGkSxbJVrQkSWMiPyk3qU/uhTTH5bt
wkMI64CkUQvrNp2VL4oWMncmspndLy9S2LgMVsY6wlIb4O9GwYPYyiQiU/Ay56QLlGr9ccu1TzFe
+HMpCvOuYfdjOu7xDTFUhSqeL4jVlWF53AIHedGEx4YcTq9PhON4A5B1nz5ihxoYc4ywMBeANk+t
Hc76GlGSxmmgl4sDc8/Nt03Sy4hvKC5idc4ociSfIds9Q4FrOg3mB84UqomgSsbXm0lnVlEoUdrz
BnnZEiT+3BnnmIaVpJsbHfm5Zigt1rbXlahLWbQ8iuF/LzBG503lMPTnqgA1I8m6ZtmMdbDIuV15
nl9noVBtUYt0gKbKuBtAG1PcodmQEogM0lA5isPdc6IGt/HPWNFEpoj2VlTifE28E8kca3y04jy1
9hm9CzM+KdLoOYSqy6+6TszeA2A9vzHdxndmsve8SkCIex1ZY38GnRFA42ie8esQm/ZtemvHgUt+
StNFf3qOxYq99ZD6TFHmSUUU2sAPbv9qyVSmygBygIXa3nF0e/1kDim8YNAgXPmQTUxwtuV646gg
8XxwPMz9s62t/3NK7OcO99XN1cGadXY4v43sS3Ak1a6//XFfcGf7UlGeSxWBCWwIE4Wo4E0CIDAa
1d9gcaBauTWJ2hB4O5jpGAgz4LcGpwdaAJvcEPvXfSZkwZDDful36K+oLYXI/q0q0E5J48Ks3uJ4
0Qn5nUdwE9N5T2WCCsLbY5GmcLE71CvZo4Kv45eq6l/qm4Q7QeuMpXEusdijge/b8LZxUjAET1zZ
pWb8QsYs0mwlap07CVlFqLSY8i671fvGo9bTTw33PKJgvkVbltHh+SC8NyB/6PmBL3llB7hECrDd
XYBT32gC/9+h7QL4NcjMqJMvuM3nHpAB+C7JFf06fHFnk4xxlfYm8fnfxQ6qaMJ+DAfera1LjcB4
Iryo5nm7Szvo8UOaJWBlwolmvjOOZi95b9IramctsbXv46a6w/bAThPedYR8jhTZprNfiAVFhrby
9F8SKznvcwJd7X9NXE20rNCTyr/Oi7FzaAHO4vlgotpuGPetn2SEJE6wpbKh3gdup5XuRSbDnH1+
UGYomb70xBWOLVTQsFzUtGLmSdou1NLOxTGGmosCSMG/ZAmpsTXIzLCvLR1hsYmeIurzUaB5I7VG
bXHfSRCmw1fmzr21fiwqrH1SavKKyMF1FMcjIiU39nKktk7uo99zVTfWs7nWXc+SY3cowNmR/V/S
GowLjUEQkN7VZPPjYNCa+D25x6W8QYLvdhCsl/ZkEVBucd0Xdt9czxTqjwziBLWSXNil5NqQcSxI
+jkFywNKVQ9nuDtxQIUSIJeSWMFytQugAn55ENWicecvxW8D5plDk8NntAjKRNxVqYHoR8fKHKjC
5tzGzzQP9f05agFQUlJL0W8H/JpieTPkptMkrR3Aduq1QVMelLp9OofAKkt8PVlkOvJEseDWIR6m
YG6oRN3toabXLFtWQQIfPOUz72dXRee/caAGMXAVlxWRJwI402DlUXi/pn1GUnCwSUK/d1ZJW+1g
BAKADI5PwHta9AUy5Cde20Sg/kIoSPepMqw035WIaZZVNJMTVPlkATfoV1dsteMxYNK486EjXitl
VdBXaEK1cMvORgNBbapS3zvYt1aKBNxtbyxd3FJoDp9jm3xELuQA1oa7FpK9O7G2ot6pW7mQi9Fq
l/sFVVHWGmKccmPtHMD5uITV8XMtNT0QCzcwYsjLp+O+UaIq8AHrevF+mRLGrYbfSKVATqSgDi3i
L29sYr5mPNlD4v737+DtGf84Ycl0V0U1LC6S8O28UMTRJU35PoT8mZ76CmJCHEWFCDsWqwyO8L+n
P2vjjTP5gf+LM0vyMatTx+lE6+E1gIN5rh2LsLovINDIQWekBTmut0BJkOQYoGG4iNwD47lkw5Ra
jnWAqJj01z0YaOJ6ykWMC5AF3ZIsnqVHF4UTKSuqi57mjIBMHsPuRkUFWKdeEHu5GprgW5bU+zAE
xtw+G0GF8QteXnaQNfQ4XtdnXDr0o9qtwDuSeIgtfgJH5IAbMUyhEMcNMZC8lN3vAdgb/qKfKWgI
U1wv82UzUBZxjc9KlpGE3/fMG9i9BygV7llYw/kCb+zQDuAkBqUvZ8CoWg3Hb5QDkgUROn2yTxBz
PwJWd/Dd6msp1in4qA5s5nopGMQMihTmZde0N0tWbSYJf8YF3b6ykIstK3wfsZJBHuQjXg+YkxE2
o1DKPTJXGPDK1QF0E3opiwccNCLSjnq4T50LVp14y8PeiAKouH8HTnDkA6Jl4EWlX7IG4k/o6MsR
dAOmbGoGIRXFvLaRHl0zuLBG4j+3+lpnNJhs7kYLQH5SEO5UCv02zPEcyzDKmM1FFjo3b/vyerCN
VcgjeTjH9KlBdT3+aC4R8hHe8C146KjmcVS1/5hsdNwqLYEGzAhe2f//RUEBSegF0fsnQUEMziln
1bLLr/ZG3exoX4hVjQqwYQ1OAbg+A+Oj+nudzi7lGtTzwbZlOxnEBhndo4IZmFFPtAlaKkymMakM
C0HjJDMvXT5+8/fQuc67hoTDSK587kKzWKjrmkoe9d4DKgfiBoQ8JX6rl0x5EY1q4RSmAUQgnwhc
Eu2jTBIqBd3FzcQCyvaWb/UpFrJG8z/19NYZS2iVMSuZr06Tl2ObRtunJLzfGdlxdzI02mIPgGU/
4Flh/U78KWJfd31Ubug9AwmcBIcsfU2PVsJKquUiavh20ILmEizWp+GoCZGHVJNnnIWaFr984AkT
nCmEEJst93eHv3/1BA4m0XGibSHQpI/nwfPtQgSe4SNQaJCWplkB2IwJ5ezzzECHKsbb7BGMXfAF
NBUSYAoKTovEwdVbOOqBEUO0F0PZ4tLt2uCFQdqT3pFyHnGjDll76sgSiCT9d8L890+DZG8+42nW
49aH1K1qf0sDNzNWpHYu/Bvw17lEfmr4mzuxow0/3TNkBeBbAlkGc+681MUoyYNfp22DfPyiQ6E5
qE13FOS8nh2sHHZQi6va6fFYYgyqQUoa2oY+W0PJq5LNL5s6vNiDu/CcZCiK+wS9L5A2rI1EJ+Pk
84v9b6wWaTQezspFAvQDzB81lLTceA6/iQ1zG/jm0yfiuUDgxeLZ6IjgWKxVaj8DRczn0huPfNXp
7ykGP73Ih4ZojcsdfNWeQcl5AnlUmLeMRA5GNxMoywSvo93nfEupbdNLXzmeKU8f82UYeCgmW02H
smWj6pprAeaUDicL0n1RCwS+7sFd+F8+Uahe3Y2IVGZ//SLaJDjG6kw3HwIJKkp5BO+j0L9DAzsQ
JRIonNDGxPbzgztBwzkpw8J6aUubTGWPN2P9iRs27iFktcHxJiPa0p+NFJXlE6SDMjUeN63jpH+v
9n23BSA3KMCQ4wp400ZcQPI27rRXIkEjXAaLx2zf8/OkhqkgSQCwKkhLXT5mn538RQnzSEneLYzY
uS+8IFnSVLjjg7/pmO1pMIvP4rNfYYNd3+2AfmqPYYIZXQtiLKAA89G327ZkSzRMgyoGW1C6ozMp
6svRj9a8xZoBYhI5mta4zgyxd12hx0t9xrHjZrdhHdTTESF/6i601ysi2PkcB2isPqKZEchc+rRb
nNVglX5Y3jh4c/7bzCfgn0z+5M88SAAeV75QhsHMaaxFl/MsTcv0K8zJ7WiO/c/2UI7/YCI/WPua
x+CpdYBZ0hJD1neMD9FAsBmJkul+wiR3OgYLjOCoWLsS8roI6b+UfEZtOG5ESOGnge+DBrqaZTmf
gu/aS6wm41DXHJawwzaoHmWCOc6ugGMOIiUkiGzw8HElZ/ps4r8BsuYmUw2y3i2CiWCE2SRqbRnB
oVsErcvTVoNTqUci3R2JQbgNE/RIDVki2e594jH66qyCSpSh2BYkqeRPtiiLBPhq5KBsPllHZVOx
l91PJ35yo7n26GnB67603v1o/6NjmQTB+gFU2izEQChG1I4+Krh9Fyye1ufNYXd8nKXDWn6h7pP2
/Y0fIq0Ln4cZFRw74pjQZgrn4OLz0Yafcpg0q3BoDs1wGNc+Cqy9p3gj7oFwb4HsybAiN7neGx8Q
dSjVuPgt/L6I2RtZ7j+3WtP3tECwHfz/Ny2W9HhiIVJ3cKn42WRT+tImtUTuQ9qa0hJQ01qLH+fV
fSj6sZ3XLGhu6werK6HRAby7pr8uP3pcO+9SU6tDHHL/nooBJANLVwKWNpRc3b48rGVlIhHFObGJ
xWX3myXqGv1VeSSdIU8AbGbHy5bvLL8Jadh99Imkl2iVD0gaekHXuaTYwZRnFIcHBoR5Xny5aJ8+
FCM2ee1aFtJbOWWU8ZTAPteSW8wcjQ9IXf/GImDrovqFohcgoCv0ItQegfiGLiqfrZtHEURscZvX
69y1PmJVU3g9Ck3mpT6xVkjoY7xGTJbIizliXraRTTxuzQf0GwvrBr215750tr4SFgjNM2w3ciqY
HjTFUIPvQCQJiymgRi6M4NaYTSEc3rEWJLr/Ilis3MLMrHGA+z2wtaC9Hh/U5e8CZQoa92AcArlO
8RUyP9AJloajtsLcztggysmAlL/lPvOCUWM843uvuWcwfWqnQetpqWKcAJZhwTt6QUfce7ZvKUy5
c9tW4PmJySV0J5tfKJ+yvhYUh9G+JSdR/MQkfppoks+B2S0GzdYIbUAybbWjuVSSoHpri60pDyEA
72j/JKjHH25/zyDFiwQ/aDvtOiVWP7kEKh9x7kz/Kd2Xl5sHR1Hufe6UWCZpWbhWgviYBAxiQgTf
67iExCMAye13lXmTA4xQcqgiB0ABxPl1yvgnuNpOxXimkHCopV+4ZnUUJJJ8+7cLX6vnRh0Rf1++
6OYMYzVGw8pLYfG/eehXsoEwxUQPWV4vbNC+rsI1fIP8gaAmAIjhP0ptlJsU/wOBA4lv033aj9wC
82OEpK3kPCoOacik5UmugEmmqdMwIwmxtKbNEDyshmmrFGXgo19YE7fscGIxEkTfVTRJKBiKHV6S
eCXgmilXWls7uoHJ2qX1WdH6w7PBbOkrXX5bwV6PhhCK1bzmRajJ5sZZzNVRd7sUZEbG+0gTHu2a
+MYJUryohTLncnIDqw27eO+qE33O0QdV8WtAFAEmW+P+eBaYDlriLaiMqY9AorCo1ZNioSI4ZA+a
IHXVZLbkyJhy8kEZmi92Y6AjMTFe5inipdEkJhJED5yoFwbE7ie8T8XIqHESafQ77EOIeRJtBofc
IdNa20El+n0z771I0490sxOQbz/fSClG77ORUmAPXkVTJKFYZfo18qrCEWCdHp0w/bWR0uaY58Mj
ViCyFCntqrfBDpfC5ywLlT5kstNTNwEMYDmJS5s1kxBxsRI4hrzUq1YAB/JA81lymkL1FsFFND7J
YIcMgHL9HkbDLkpSk0nOxikhKWQNfnZOjmk4XALqgkF2uoX9f41a/OaDOf2WEhpqJqG/y94mAH4G
P9DiFk4p1DmE3xxk2w+tucAikdFziYTpixfQNGKyjwniCzC+sGo2X6W04zOdfqdcYdu5a/D7Fk0D
spP0FQB1l7aMbJMqBkodVG8q1VNM8givHJkByZT+y2t3y0inc9fWXVJdZ6+gPUQNpXUKm6vGKzWb
XQbNDdh8pENcLGKNJcho13xhPTygcUFOYyrbV1VA3T0J7O96UBqTdGZzGR+xh2+rTOPlCV8j2qGA
glZin20uvWhTOlOt+xmE3nGPr+PpFMzTqIzOz3m5D2c+12H7PwqIQxqNPPJ/eR0oKTJ1nl0QoBcd
CLNn2roBl4FdR6PRktIPGK6IIcnP+Ysq02jhjjYH1CAWh7pKA0rNV6ksufaV5tEmC+lsIkF3Ju9V
lccHH1Jyy6s/s1B386uCpryvJZZ/Iog9aMy6n+8On4+JRokJW3VDJtsa3KOFZQS8ywnnq4Fqhxn4
4OV7cymV+BUBLa/IZBdPR3PJj3QPmV1tJFw6y3Tfnpl3JtVJp/5OqmKbHjHg4xm3Y46u1rXvfu8g
PzsTkDCoUnhEUiMq4HsPCV7xzSk1db1jaGXfA2bhy1JDAG9gq9PwfQJDilR+q1vlV6qL0roPn8kE
yDpwrrP/ZQhUsx0rn6+d90UZToQVE2+aEDHs3H5ATm/IKVcBC+H6jdAXlIIynV+D0u079Isy13oG
pA1d2F3HPtvWwIXcfIt4jGdyq16CCAcW54dEsaRps+ssdIZym9F9DHb7H4Yl0TVfo7C3gpQS3FyH
i+YqLucaAmrhN3V6Piek4tTFummQ9ICrAr1I0vo6F3l7qrlZDejOn0h6jPKQUp8WEoHajx7tzWfm
mgmaINwH3nWFSDO+hC9EexAqgMrKkBOEBo512Tkg67w2qtP5ZElgbiLsohdG0i20kxsmYyX5XwBP
C0ir1gOIxek+Hnl/Yry2dX7o2Ery3TOJ3NWwvcfqF7wpzO4JZ50s8gJpWinR+eF60MtxmFim03gy
yUxGABXpcNJPlf0LqVhnQoUBr3mOR0M2uYkqB4hZ2I4OLmD6z8LNX2oGLCA/BNGvOnp0vc+lJ5qk
JvfksnD64g7DY+6Do+YMUvexOfAQmhNOStGPDh47RBfw+HKoRcNYWdsYlLOUcLuMR1WzVcz4ccLS
k7K+Do+jMaR1y2GcILVs1Uav/8DVCjvPxE19kn9kUyHf1R6McTGmGmSZy34+DwdCzQXLvB7vlGrn
IHmdndLWi76inVoliq5zRFNpniIBahzkrgPyms0vPd7Mw1xTs7iCbX/Y4Ts16IClb7463KzwLlMx
2rgw4Vz52jKoqEj5UVw1+mJ5xHlvo0ZQvX7Ceq4VErRwgq/A19560Y/2zMtupGdcVjeQOn3wjsl1
hwEMAnUEvOhY1toRVAuXyxZDRKlcfUspjQRfDNDob9FOvJJbDWlYzTjph7IV6qdCcjAigPkufaiZ
UPiHCJdv2ho06a3haCYg1p7JJlSlAnqUq3ADLswcgG0EXj7JvQtQ8aYYYqDiyygm1qRGWOcOiuI8
OHYuGi9jKQ4UXqyVmQdyrvdaAM9A9YT1fKlry4yIiT9oypOiwnMzmpZdUbYjI033TXXjpwSeCkbO
xN7D8QHe3lDodGws7ML6e5weBbLp6H5ubS7+RDLKULWVpLpVGpTjTRGdWWACk3Ij2hKO0ccx7VvR
On/+yaQ/I2S3jx6lBPlnTgOfjpo2G3WvJlS+yK2tEI2Vk9Q35O+8sfVD7kWF8O6A2lMYwcV8erqc
mAhGqdvSe8lV0jT6fisbGq3doB32TEnflNz9ur3GxCYeqdNi9WZfycSzOB+Tu7VEo2FqkBCzg7MT
whu3VQ7+jKmsTthIKQB352yVLsOYOvlgZGZmgfweL0bfxGuZ98oNPsZKFUoRonZdbljooV7aLBzG
dZrvXP2+m1qtPWcKgBmOC1XeBhcEX0JO7aBs8g+hnA2f1wPQ+tDvzrmgWe3BpDnvp+Jkf31HL/uH
cUInjJr1Slhj4FHdMi2f7LiBQvgl14Ahho6v1gX8mtACJCF6EjInpQ5Y5k0vWAYF7BJ54Wjb+Q4M
abXm1pnMOEsezDmM6lmP7H5WGZwtgq6FOdn/I6Mc+rj+4hdbAJ66Qbq6nfUft86ewoBHRnA/UmZJ
837UthFBi8YRfRjWlbWXU31h52G8p21f4LeG82SEmBDU/M+masmXlzs5ZJk3pawOcej0Ct8Qs9nH
WQwLFdT7BOpJzeWR/fq/VWZiBnrx8ZiBM+EPVshDI5Bu0BJe0tf0wysKG9X8m+QsiMqfuxLPvegL
lDjAPB3CvyUemhTwTwidfVy79ByxebryeCKeisXG/GuOvSIWEbvFb2BBJL9qnVMoBm6UmiOem9Xh
FyI4uS62yKyBik3biwL2z1iTH5DtAfv659uxxznP1DvByePFG8jijwKS1MQOUdTGg3qWlXSFCRV6
VyVnW2Tohq6VsmG9CyR0jwz6ZCSUe+Iyqlel5HJ87PF/Xr6cjufb+s4Or6QhkbDABsqo3brsD2/K
kuzPX9xf11XtpMiWNDmABhpQSiMmEKK6slyZAd33RqbUeALCHjHDdOhDQTLS+RezJs9QZU6CJFM2
oFBvxTU9GfmvpBQwGAanCAsxWnEodRlDd2aD0aJ9fq1cfeQgfE7iBMZgVlczElXcoSkdOISvpamN
1EEJJaLDnmUTGHptT3DYa1mJ2Ej+16x7qik8DgnqNkouwlAoK3WCpwFq4Q+dV1uZI37hUMQw70Zm
T2AE7TLHpoJ/aGb29NGiYsGplD5W046ebIKo0P0P+7yef3RydNEoMqJdVdHXKSxf3vpx4Bnf/VOM
ekLVEKVPTELOWhDOfgUgKAlQzplNlgHTVEy8yOThb9DCyPmoJC+CwbwYs+lEil1iCyJl4PSev7Le
Af2/PfaUfh+SSv50SsO+u5i011qStZ1x2F+uFZvtqEz2K0ul8I8Dc7bNtjDN6ZGn5DC6cQKT1/Yh
xm5f5Uq3eKSI/Y9OuQiExYOkuQb2Mv1StZrXGO4aua4LiafefcrSZJ88LW56wItXkKa9TdxZWu2z
VrNNNHzsvgFOtZKmX4Yr3kHvyEC1FY1A3x9gGuO+ZTTwN6dbfHl53htfYRCuuseG76mdxmBzMobi
uX+sz8IxX06TdQvnNs10VzKbKRNNKgnD1YKOs8D+axy20HEp/xI0zngjkmTqA9X6mDsQeaO6Gc+k
rNO9M9NpkxkNRW3bfDYsLRKWtc9zFvoPBt9SoIPrbBpT5CKdr8C4eIuZ5AC+nDMOKEkwFaih3C0e
9hK/bl8ljd6LcN9jepUwyYuvoIDEJYc0i5tnw5wqF2ufdgeRHJqj9x13DJKRRVySuCCrCFI4BHn2
Tk5kvZwCfMS3IfhwSDwDXYT2tO9EJgr3+iAVtr4j6WxdDwIm91fKZmvjG7DksCj9TzrcFfUhkMZn
Vjr2wdRmaZWgL5D4Q1Os3sdnZEIxnfxzt1Z0vrXrJtuAu6h8q6jogmYgNLVkw4XJzVjR1Lkwkcfy
SPHLZpGE/MnvV5KwG1P6LGmIxCBQ25b9XJYyuSZcN7F3zEXLeunyFCqMBymJH8yGnVM3FoB0hun2
knbThkCvKfYtsZ5/c3jEc3HA4htLE7WQ6dyk4PvLh8VQMIYA5jHmXdg4TXafst73tzc5HeTzQxIM
ctimy0sTHRKJNe6ezAcgOJsJmWUO+leLE7QrRAeY05LC4VmVfSb4o49L18iPFng2RYcLiSzdd8cD
lc0rnAcRAZaaO0X8yAJEUa/EItSaQMksKUn03xjeDmtrq33htwJcjyEEKHsI7KYHR+cWvzo3cGOO
Md2SguMmr9BkWNYbHWP217CmeSqG8LK+R+TlIbw5+vZPXOYJiOMHAIGc7Xi94mXTppDUUzc7kyw/
1zeoFF+QxGTVD23K/O+r7I85/rjBavVa6P2KOiFwwcFYMWaSxZKkA/IHkMvWQnYJ1hFQ9jOF0+0q
7Mm0AyycgZELsFGCSPyUlRc7ACe+i2veCPpQON7OHayx0cMbbWROQ3KnccdMMDUppGxCJd8H1MLS
UI69c/ufKHSWgh4IIoDmNOgKC8054uu0eQDzDQ6Pew32nJeI0Hrp+Qboc4DSe/jN5lKQHGrELU/U
blKjd/bKi3DoUmQ6Bhqed7gqBZTbctxhCNQZhdUkKNWpk5y4kcd23jw7AyMoFbz8P6zmn5LCzuCP
OzsOSbzgHhtZGwEqrrMbfnGC/iY7040+J3xE/kDY6B890kZjy9Map7xTUWEW5Z1aCDro7W6SSiZ7
N/ImdU8KapFJ1sTnOxEFuMo/cJZvx5civd7uGcQrlwD4j983MNYoLyCjM48sb4E7NWzgbG/nJZZs
b2yb3jYp+afrluUXLhgZQF+0f44I7jVxJHx0TbAaNNUseGiEC8cIEcazqZz0XFaTmg+GNticldHx
doVuDeltAO5h0K/LxsOsV7WtZ506BOH6Dofm/47aWez9L4UaT0JELMWmNh4oRvJ2JNMSRaNn1f/J
Ljxwr539qbuEmeO6d1S1O0CBxNSaWpsGVecyScpr3oULerG2+Cpy+wFnASeDD3RK7AAFXynLPPah
1RRs1pky9MG13vPHmoSVXi3Lw0c7m52mGjkD7HNN/FQHp/qfXiBL55ostl0ujPy0NTqKg5asKRCp
5UiS4TT79sDYS2p0psn24qZ0gSZTtkA9op71Gcm+SUyiR7BaOa8BMOIzI34ds4fp1Of4aWOXBvuK
UIWsZbaJUPDZ6aRjgFjQWiQrx8DMkEnAe8nzsyqlDZ3PqJFuvK5+megnpeYqn0LIWdi6y3Bi84m1
sSAN3KCs+/Qz/+aaTyOfPyUlhYOPZrPRih3biFcr3YsdhyydFEBKsn/EULliW9ssu36qVKitogHQ
XASwS3YFO9I5fqo58H5qe3hsSzSg+FuhrVqhFcWjwECVwaAjFlkjOEJNTAEd7t/EeXTmc1L+Euw0
/sYRCPtKBicDB4F+pZ6y0H5UahCeCpXO/rpBduB28sfk4N7YwEI3wXPb8twZu9OAiF3N1+kEmFTg
UPv6PfTOZezcxlpL2XiLXB2M8tcJnkE8QlAvWan3jbkgSe74Hv8B0eUr/H8UoRb5g+GoKxWbx3zL
qfeESocVVJKCxcWAdaseE0/fjPDBifhWDXJc1EUxFHPYWEJOCflksCIkREL/97WCBT7gxEXgP1de
3rPEu+3ilymATETMmbkuV6bDKcE3cRJxV2UfS2yZzHGQmtaKAYhBe8NfQwYd5ublFIPR5QLPlTsz
TdzZKcsrW1Qel2M/+s9JtMexPzc6VEp21/x4ibeyJ0socV5BIri/eQKF3Qljs92bzQPgfI5beAFV
2jv9frj1cekHP22l7JtmqD4M3Fi/KFsySeZklVY8HAIciIEzVsmDKVZL9qu/Rdytq1oZXzRHQ/xG
P15/Tph8S/E+JUSk1u0AZnNwUVFU+M2wy+CZGw0DJEw8m4r7KRaDOAgM1xKrr6TqqOburKbmqGRp
WbHYRY36B6ZXHPf2upk+5lM1yd4ohDZzsBRJtNH5pdpxDKf3W6DuBOySGFxO01iVWRJm5yQHgB7d
vEldt+9JKuw/BoAkKokoIEGsIHPmcrj4Hh7UJ2mowQ/AKrLSXz+khnCbRJk6MWVGuS8ntcOf5j5i
nkPc/ktHQopJ8lDOXlO9qfuB+6kheLBgi2jFOmT+CKkdw3dBccHbmoQfvBdluoZ2LSlam0E3Uy1E
x6ZGNLnejTHmVl/dg5UNBeelcXBFXCvOK1qg7Rxwj1Z1sy45JogFReKiDwl6qzbcPXcEFW72GEuN
Fh6Xb59T6LderYT5u6l15r3cWyM58N672B2U0QHqIQ5JcrB50ms/3VJCQvMs+KCwMgJOtJwfC2BE
JIyGBvFcS1DLXf7xyXo1zDAmPglI0z2g9HW4fs3iU8W5Xa4ZH9jzC/6750ICn1UhPWD/ra92OSvj
4rOeEMBx4AffsCIGDB3Rs3HQbz6swwEq5LyZd7KCNA+VjSjit81HtbMmuH84jRhtTOy6JXnbimZg
265e50a6wT8Mx1mcKLbP/+0QMNvGvo06nde/QVBYxaQexOV0tWjV3pGmD8uub8KB0dbdiIr5TWKk
6pYW/dVXy4FBVSbIfRaYfMvmzjBe3rO6Oank0K+Fiqc4iGr8bKRPE+IMKjyTGoJNZieHHHfcfLMN
U7rcIaJBlZQHkr7scequsDYPiHZUHwfjgHR1srf0nW6PzQzKaisGyAyoN3xboe7Li/MItwXAT5w0
gTOSs5i6Vl0xgkDX7OUY8G6u5vSgNEnHV7zh572wJzAviiTfBiG6qcq9TUrJwaicQzIMka2kouvV
Jh6JLgEhcEEXFFbArWswtB3qIlYaCvi1Bn3a8nqHVm9XFVxH+uglsk4O/KRwd0xbz0ZyyhDKDKcp
yAmS61zt6u9UL+Q+RtnaiYhTBtDyRbDioD0BThlZ9ZLG+NT89pEvqgL3fdcIw4BiuQEreFiKj/yB
AYXEqR8nTgWRQQrO9q5Nhrct1zwF6aE3KKNMQD4RP/M4OoO6vpvLQHHk635sabn/ZwP64wsebSy5
muZi+Xgl3QEVV6h5Sj78KzybXamgTRsyZCMzBGosZNzG/R9p9GRcLStz8E2N6hyVbE7geDULusAr
B+d1i0yAHVwRvf7F/JeO8YaIRwogz+xJbn2DVlryLwLlUiUTEB/uumklofLdlC0e9GqR/cNeMnHD
TFRbyq7sye2D26G6gCXZojcYyLWT6QOqulGX62s2jCGTCvFkKb5eVTXCSZVkLN9/ksE3Nr43AOAO
pQY+cR27pMLpEHGspP1dHSWpDMql8HdRyYYi4QBV0yfNSwpxn+7IBRf4R7Q/Y03MsdCQV77AU7iF
aoTt75bB4IYv+tJ5PYtfrjFLGSZruWz1xEKmpPSTj5YIje6jigw8AI6fyWPdKEUvvHjUfKVD/95Y
fATJp+8akPqGTOCXg/IIKW52HdOcGbmFXvmm6Tz/vmv2
`protect end_protected
