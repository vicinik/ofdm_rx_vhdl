-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WyRh0ZvZzr/DNmzMLiSgMPAxYFZbjpGGnrS6az7nc7vsRbTCI/iqUonQG0AvPmEIXrkQJOVEnytn
mIl0FU7PVnNBLjPhdOfKij3bLq4sleF9LuMuLGSIeoUZMZnytfnymw2fCGs2CgbFnmpf18xs4LOr
0o97M/33nPnta2uiT6QblDgOEqh6zearglEFmBh4qjZrpOwzIYiV0tCKYX1MvN7h7KfkiBRcYPtz
SXyGRJUvotz2akAHJla9brNY6LhLzqXT0c8IO+esm3b07RRWitQIhpu/x9vBkL4JIwo/if9CaGfM
1XuMqrsUfDJLl3TRXuDU7mTPtOP9Xqc9rqXMzQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114656)
`protect data_block
n9I/suIAdVibGorUM64KkIwuz8geDu8cMAc5Gu0cTS2jMDKGLc3jpooiOThjynBthkSdicb7tLuy
lV+Sbv9FITmMm+i3JoUpS4S9w0iRfqyulDFAIeVjGKYkm0aASyjqtMOwD+Fom6O9erSCnLGmsWyP
3u2N3RvaZ4NICOLzokeRAhWwopEnclxW8ue+M6pL8S+11PM4xDO1WYL0SeLcAoyrojlTiSeqkeCw
EibG5KiCSZKpY+GWg4mcgwfa1FiyvUAhAOw4OGWwze7MKiS0n7yfPpbQdvWFH4gLlc7U7XHJzDuc
gpDI0ao2spCv1uWqFm8WT92tXSI8NWLJdSprWZuLR1bILouq7zftAtGBYmfYmi8HgKlEQ+YzLQfg
wkjuBVBYqz/V0FDXNVJc2/sBpDiHbStsv13ToIVcfVH4tbU83NOkp0hQW4x30/36IbDHEr1sMPlY
2rk27tUcgqClpSiBPQvobILAb5+ygz960TqYjRZqTOcCJTiNerTLl4trBRg5WyyX0MfMMr95ggwd
VzV+JS5naus1qFDqkbtIarHrPa2EvT8gKTFA+zbHqwwMnjLTB0qwZBw8RdEZgzZ9SvnKlmPTtyNV
NxIm5s5pla2P5ixYX0+SP9HOq/TaNfxebrMSgjOhljxYooppczjr/VRpWIxgBRHUKoLuM3UL/Xfx
P9hMxDDORBBoRRm/4uFSdSjUOQ9f3atn4N4s07HNAN2u5JOggRe+qKgddq3cGZFnYOPYJvCzsWuT
a9GauYrswtC9Mr9mjg7XoQ9ecgCiRrpWa+hoyf0WoDMhSUSEKy1Ky3K+VyEtcTzlZwwwG4ktctOi
SFlkoOikDrzmyXzrdVqm6rWLzwBrwDeAXOYkpaFjCInY5yWQUuy4VYNPahmeU46bYHCEj4f47l1v
6l9RIg7LbxscPrUicbB9gus8RbhjagbU5wU+cs3Oev5BBm4hI9D7Jaxik2yjqRsOTV/hwhcmd2kx
vKT3bRUR5DyWdWMDnAN3nOFRDHnkf/PT/pLj+0zvBvWx4EsxtIzBKU70gCDuxJbIgPEJ/kmPPk+x
hNmLcgw3ygTbwb1Zs6JhNjzxV+m/30De2eQAwmsPlhAzymx4sQ0l1+uZ6uYAv3UR528nmOhejZel
d4MlkT2DNJ7B14Gh2OsLSDMBYKRRYNhHJFTaLjpexI689rM3t8Ntvpo+m+jceFmbZiYDDxp6qfsM
PB/HnYcfbgs99Q7aRcLkY7wE65CB8q/t3usnWiogn4f0KcwMHdLpFP5Eb+ttZKGJYX5VE8ydQbF4
p8AaMfY9f5NsVreKaso1uAGtisnUjQyZb9v6FOUyyKQ7YCBIWMxWeO+lgOYSnD+Hh9jHS8yxFTyG
1+588QJXrbHFiaFVB940FHMEG5G82EfuxOKqKV4qc1x81PEFMW+ggGiOhvrj2Aga5VTqEvGyrmkw
mY5oSG+1xiGGQ5dFJ9Z798VR76J3HPrjOCpOpaYxvDIip1OATYjPat++9uc7qQyfBJ5sfWxJ3AWw
orzWsqfrCjPppbAHWHJDOjJ0S0HOO6hcnPaFtukzLS0xULHlSKfUpteZYH6NlpaaTB69qnvuwVEd
sa/6oAIsjb1mY/YTqZZLPrUK7ThQaD37+0tXnD+u3nMLxwmdhY12lHrfQMHIKiBthAjGhfIaLxtr
4aZWbQlf+VKW7dhXBnWQURIfv/4YVLfFxbuMgdbPexv3xLLTIpKgDb2ADRBD1ZNpl2PiEnGS4swh
Qj76lZdVuDkydInFlFONF+swY5AmzfOBzzpTSScVgCDE5pfim0OsISdUNNvsnQ5cWcTfzstUtrWB
j+rBYgyyNJ/cLCoOcH+0e4r3ipoDTS9vYVv02NXryA98avJ6QNwrtfJZKb2vN8JzydqLg9he4VNL
j3EvQ1NAjDnhVCumFjbObwIghp6cPnPK6NeORjqwtAw1LLtUARCMD7UluMClRFsFX4rWmtdFD7Lv
lbN8Rgaxxk8v1KIr9gMGzpfn/lH8TOQNFUPVAKhgQ3xy56ak5lWWktgD5m4knQ0psiMu0AIUhhpT
hOvozY6U0OC+gTrJ+s1UtbSC1y4BOewZlHx33zDGcxh+lJ3XGyjzpwTiZQnIqOn2w/nw4S5QldTW
3EHT2+wqxwaDQyUCiYP1FOwoLZWQ5n9LaIpN9ScPj2XHZ0+0/BBgaZhw1Z4Jof6Z3z1iHO/HERyi
YH6vwOh1lxGCDLMvoEAQ9if/0EIKqrtXcDDr7H8sVa2VtQNlqEVp1od7VNmaWNCH9YzwqHNe5QzN
T/uRmDDuuER7FxHKkICQZrjTRlhZct6sM1LNCB3IU1Q4MRfKi1RehPveOiFjCYbAra3DQ8N0m2Rl
65TsAhOyq83slnANgfYf/ZKoSeUDTKRykbcF8we6XGhZsINH/mIIm31GxOT6ZT411EdmUFoMHj5R
SV5YEDeButofaTYU/shVpg6ePoNJd2T17ABfzfpqBbmd19UzJuifTjz0x7iqQcdw7EOPQHW3WbeV
WkrgV4Hzt0tYa8Ibm3LcisKwx6bva9ZxuY3FKcKLZCprpvOwUHLPaSQbOz1NCl6c1bESkTuAyo7h
pFhetkIKyJu7EdgJG5pc6C5q4pWMJsvNT7FEExZK+TV4xiu/TPLx+S+eAmak9LXpDT6ey0Va04LJ
hbQHAdTN0cKZVuz2t9wdRQo1uQTJqkO6RJo4CaYd3Ts/X3c2N3u5tsgqnaC98LU7B16SDcynqJpb
w+EFvlN/XBIumhJ0ytkgmnFYawGcsB+4dmBfI4mAKw3l8lLYrxsPsAEcXQb+tlLxaK7iOU/ny90R
1RTak5g89w9f0Mohwnu6we9JGmX1dYxJwbgDVs1KahlfeDbR4YBjX+KL9Bdt+M+Up/OYS8p85zvc
Ylt3jp3/6lrS5M41OfwaOJcCwjE1+jDZjt1hJnialZWBTXxDTKgu2UKMw0zvRVxjJTF5Pwr1Kb+X
IWPJYxp5i4fns/OEih0YVgmNsK0AXwORRtkxy7EmBah9IiQ6/aw+jugeLpOhAsXZvP04p2Q859lw
JYB4ErXuFus8h7E2Tjv6F4DsSYvupP/JonS8EXN79nMLpYhCDKJwpkIofpYwTjjG7jlyBIXiUcoR
w8WNvAO7DU6dKbcCdvuPrYuNK7qZ7a3dTQFJ2PTh8IvWX9+5Y9fD1KMNfod1R811iGOkWea09ACT
1TeHM46NlTxj7Ou2PX5Xw32ouv/oCeOZaGzY9Gtxde4T4WMN1oo4gDfNmKUfasTLn51Kg0lOr/nw
7FjL+/PLnStU+ecGsK0C57uHIKdRKBSpRDDQA+WfGxyUT7WhDSJRmeAWDP8NiA/XKda3i+3KOjPW
OTBbPDCh/y7Yj7daemdexKfEm0+ZJeOb9mp43GBAo0Ixd5rBkU03R4rDNRbYSLDVJ9ciOMOOwVyx
eeeE02Bk++4A8zvAv8tq/tHvgXotkZrTq4vvFOsUJOchgSCLfTKZqCCpK71SK2EOPMMDX5BqU29e
Xlmti8yBTP6drHa7J2Xqp6LxeCa9jvq283NL2gpCcACJK83aVyDbjTSRZcIyW1wIZv21AD2s9m9Y
PRAwN6EyvM+nwdjuPyaSRq3muSrPj5FNrfoWPU0rpaWpxG2KB9QlvtKYgk2rEyEGVxPU2AzGb47n
k8ZPPAr0qHY1qCg68oSJJNe+YSqOXTv1Cxo1Jh9z8NMV0LOthSwlwrVt2CH3pczsYlalz09KTxf3
6gWhKkCQj2DzsBEYIytpP6LWA7A9nrq2tEWtrPEOeeqeCerADn9uy0FID6dN2/HcWMvDT57NYO4x
VE7Ys0WHNGCLGT/0FLv55jJJYxZXmxHDAWvIJkLS2uW7sicmPj7ihEhj1IF3RvPfgiUL6Hzuf/4B
10Xkf8VqUs8HwTcoRL5q/0oeu9IPk8S3yvuBHIZZ1BRIwauI3w++7D8qrSuGZfRI66JISn4cmd3M
8xddhnNe5QQ8cciTHTnz1mgrdksxvfUEl33LeBluJDONHbcOEIRnvb+VGCv2YzUD27lOlHQFkNPC
yc1oFp7pK0K3vnaZbSEkSWJi5KRwjI7U/RFO1aH9Hdr0HjRPtIlqXeycNqCPvGkUvPP5BVaUQf1l
94R13iQE3TFYoxTFlhn/T3FggY4E0T3HJ1KPSrmq/jQtzqMYxod3p0DjKUGigisTQ+al1qKRsu2E
pQFV+RN5wpy6V8ir+SnB0tlIFyAZaYkF7UfcmGPt+zt7mUQ4xyRbFqyjrINRAqupnK7Wm5S67luO
WnbS+5h1Q/tRj8eZI22WwYEp/BAFRUBy8LzdMSm0iv4MSOzPgk11CZcvaI7XG3ojq6MH6MXmVEEb
fZIfN1O2MQVIKT4RkbyLEIrxggczARBqrWaGY+tkD/Y8l4H6PEP6fpmTotihKHzqN632w7feJBlr
YfLofoEbhLWTfimyHNP3aZdNZX/y3GCOxRk44Gd4YnMnIfkwmDRMVcgQYWYUHAmmPFmkgQ8l2wBm
y/UbW8zSO9oF/THoIyqwJVtmC6TzLIIXPV2etvukJHrK6SzAhH65q7HophgRCKXtyhXZF/7KALpl
7A5diVVwlMIbhZvr9W/CKUNaWgINLq6CI0JM0SoyD42ICqdMWP+1pOfWoEPHmOe/vNjwTat7xRVG
6auALYIMi4oy8k05sGFeCpVgpI1nFbhq4nG6oRf0EgPiTf/MeUyVUS/jx9ZDRgGLZacz8X4jQDhj
5WlGIMBgpkQs5F+yN0mGCROmahwcLzd57aHQiQlsLgHCt/ehD6EYX9Sj8uPHx+QWyt1yCKTyOEbM
QrzJnb1BKauJnEnIbkVAQ5AIdFzphY4JxZe6zRvSOrhq7HK7lPkfo1ffYc3XK/qTvJn6okbEnnv0
0emTXlCEZh/NHcn9pgXFEe0NrxDUxg+wobnyqGRE9EkXLLFP4r3l2+b0JWOa2UiO0ro7R/DsR0ln
vj4yRsyA9wXmUukDWHDIoC/n9C8MCYliEr/zmbd9yBMVSyB5yu0djWu9p6M+Xc8oO7MBFzk+L7fx
JODwqyOACR23WgIQjC/TQeM4Kp0gg9Tr1HHDZLdftRSVzGHhjc+IwsKIyMQDhYuYrT4oSfX56gpy
0TrzIT4vZ0/fCJ4QBStYa5qWrofYmdDJFDYiNx9T188L0+rZhHlviAr5Le1J4csPzlF+COj6vjfW
QH7iA+QY2e67s0ylZcq8A5hMGrVRblN4liuEc+3iAG3S8kMLFFDMrRNFqnepIUadWn3Qy20i1I+h
7YQPQDv4eMVZ+uy/9u99T29VKds04zg/NOuyhTzmfd2F2uHKNwTX5lwcF9FknDDtEF69TZze3RcZ
J29MQO+TeEzyh5Qyh5Y9fu/Kv+EXK+tXOxaRkJZHW7/mG+yireQiaf7GJx1GfhOuzT44zloxUYwP
BPVjYze9Z5feV5Ig6mtKP7BQR7eTsx/D+0ES9WkaEnmXP7jpzy2I/glMznHpeOkfJbghED9hVwTZ
SnZMD6dDLK6/Y0iqJ42CLrdjS49XVVq2HieICRALSNKxk1V8s3Z+FaL2wqKbN3ByGxiX2VSyhNoD
8Ep2+7NENSdrbkfMQ+Av9yeqPxd6QvQwHyxpYp9XMMioQx3Q+7ixHn7D9nln7Qwf0b+siV4Pc61W
LksbH6LAaY+47qsT8bcevJFtGzFZCHK4ss8+p+jWNjYMHB0FMkN/84row/jA+3LVajvM/CjHqXRE
UAV4vVvRL5PS8y1kXvLTgX0NRlPCWv0EF9C1OHWVc54vYNKPU88ofKr9lBokJMkiiBewiheqjnTT
y2OU6aMlLkDL4HHLqHa6vO2wwT8TQ4bResDEzv/4cjQwltZ+V76djQ4Q8oZBS+la4skLS8fRyWWs
ACtmslBAsVhXfeIzx5jlLX0tspzm7xg7gN8dZ5scOJVQxOf0KDOSgY+e+uDe9ebsb30RHEweJnyW
+xMU21WufibkvyPObhVL25Ex8eP5yBWA14aRbv/hmuM6/7oeBhw5xINNNpn9UybChLUKHZPA8jR2
EizhBRaGyzbbmCjKvcBIeBe6oestQwS3P+Sah7R/mSCkhlA//cwEZiAMo146tyyGiWNHxNH6XoIP
jfxKJ8y2Zq8JKO5YTXoLXUIpyMen+Q2sPhHprwVMyyHDtsBsuBsTPmMdOvq4jkupno6G8oELIoL9
8zhurwdrEmNNxo0toAWZxZMKrUNcQwWrrHdjsXhslMxDGVz05kvRaJ4qxvWK/Dbzd6cZ2Xtn9EDx
wymUIcQyM/1EtJI7dQUC9byrhIVxuUOdDjHZUARzJeZBOJvmzi+DftRQC+MyZITz9WxExRBrc7L2
5qFORptSONKOU9HHFM9KWaNvRt5THKX3CM6HETXxg43hgCYWDJrgE/MUsaIGb2hosQHZaNjhcmKY
TpMI+FGMdyyDvF7Y+pRu5GpOQ33CLWE6TvEC6SiS6x3TcATP1jK9lMdnvXZZ1mBUt8pfQ76GyYFb
1aKLETXXCAMu0mvxJ6HtwXIm0Oqn2YgFZy31SOsR1g23G7matPnfMUvCVFWT0h6X9bhWzaDn1wJx
q6tosQ5PzguedAOa8cchk1rC4XE8xYTZaBbBKei6KWMrCAsiATVKZjxoKJ/tAF+udH6QRom1aHMf
i/FXMVsbs+Xf34tAQejKfT7Ps6DHMfb/mu4Ns2wJ+ncbV08gpLvMKNDxxbZgBKgNNJan+JdUDr89
HwJpJrg3HFkP8W3NgWEeVqlwioOg/GCHloK5/skNYd0Y1wbYe2AJ9i63GfaWGLFVFPbI5apzknZH
nDO/i8OlFwaAOq6MLAiBHZ9rvam+QkiK1OPTEkIG42arfIsR4H52q1yuiIWg6AdSBhpGcA98F7eX
8S4UH7vBCBp+eLdC5oOZH0Z85YjQ3dqI9q/1A72S2eAxm9hYTjg41z5tjLeM7o9EKI/2ZZcEPw6K
b0fPSfhBs9inrZpEvQ1rTpW2KqD95kKafFAqxkbSYyqKTr3gT6LawbTAzb0EMOP9Enqex5g31gPC
mEv7vbraffUeckmNGJwIwUWyN8y4bz8Ec2fvmYLhl6q7Hnj/Tk3M/g+lE6sjsbnVjRveNXXv9hdF
2/aeMj5kkSiFEy/eO2URYkrcAX7CsXvt0pZo0cdyQp6Y6eiNk7Nz02dB7EcABngHOazlZ3uQfb2u
tdSKTIFTleeD+S2lIPtIZqdmOqOds91MaEZcTwfu8k24vQq7SDhJKH6r+5apnDDHy0LMG3JfPpGw
GLqedirrQdtE33oIIVPLm+TYJvnrlYEY6fIC7FV4t3nALArHlCMWrY6tVvPkj36Ck6h3qXVfucE1
jzYyORzunqnVb8nTaC6eS8kolyuLplwowFyY3OQbOx+1gzhouMh3C1YQa0h1ies18jpymlZbS7T9
igHuhs0qDgYQXkDr19sV6hUDJbG5N/J7Ya8TOF3o46A+VTaXazLU7Vwi/6P7FnnbUwwoKhPb3PNg
bt0NJr4VoAHQyIyOaeGMBoE3F+LOwZNoy0K5K1VjES8ktSs6oplcPCgozJtlURRLXHpghgPbRJMy
lBorY56a044Q5fjRzAS5nnfVLSgGd1qyv75wraqU9yYGY3atJ0Wk/F2Jfn35hIT16Z3NXTC5qcjx
cDGSz9LxDzNAuo1nzBMQMY7Ioi9RpD+je1JfINTFC3IxE/LZas9xaAdFV1cDdmSbsErIFDH3N6BD
bnJGQRFOQSfuAFu/JmsaIvDfAtr6JPoCtDV1Gi5EgcJZS/Ck5eNaq64eSe6Netxo1mlEmCVTXyuG
FsuVfztWXkNqoa9joyTwBV5849B/o89Z3qCWIljqdBotPAHT9rdPqOHJZBU9SfQ8mFQbqd4SopWL
n1NX/kXauyuK7baKrQ8cnsM9R5n5fkljlGKZGAVV9OAboKz6tMpVEHRfFs5TBvpilmlie6LBbYjx
3+bIOX4geOq4BNApLsh1lF2t2j+zTBWiXrNI15IXMa4ywuxBVuYriDfOYMCyO4Pc8TJkDLtONBq8
EgA/k3VpumK7AM997AaIUyptFvL0GczMLvM+dgtAFbNeweVptjA7NMl/GGVC6QR+EZB2CxHgLbow
XXdE004DHNdlnuC1jubtYtwDcI6HDb6XrACmGElrHovw2uueFiM2LZCo1YRVev74IbzEmWPJseNR
3NrP77GQuq5i04k1boOmmK9ubjEVXTyHc26MzCJnhmG7LoeqiyzP28eNnOX6Ulk7dt/CzfZ5El3c
riNzAjbQOgOevbKEy/lLCIcg7whPi7FQBWoocRf9Lawgj7Bkr37tQ+XTBt7JL0BfoX8ny0rTPXxo
l0v+6bgn26x3p8EsUP4iX6OUaiL88zn1cUwEUlYTRYjVh2djhFfCczZiClpKiF9Jtus6Rbrn7YeB
tXEHNlpHXzrowPalAIv3I8Ynsl8I1AofxK1M/DYs49BD9JlMXctye56RrgBWBNpHHmF/spCYB4yw
/gvUSfp/SdHOpCijVqBKVDLBsc2P7g4kunHXHnhRmrbVo/fyFrlZjILgiiMbL/tgeAhj586NIMcJ
Fdj4fZj8VPeMnYbQoQL3qVLnjHcGxSofhF3iDTbKLdT1m29nq7tIc+xsO5W8yNmLaKzlvnEnA0su
dCavXVeb+4R8hT8cFwgASBRwaRC9jk+9BHipsatOctfHyg+y8RJOLXuqg3xg9/olucJytSJjv5Lr
c90sW/IN/+PrqEz77LIBGEp4tAMyKJtFwcX2vwA+MX61Yjj7zwolPF9UY0hGTHMW/PEYdZ36pPuO
YiJROnPUzTBJV7pV1ul6C3fvcWz+zO/sh9k3KTyS4Xjd1CF/5Gy1tp7Yri9VNLuiCBpq3EvmMQmH
bRC0HFSVmiVrVDA5196i66+uc1rvMtuv/3QjUZ+1OCRYgL0M2ElYIGYZR4w7KV6wasVgmcq3RZDc
BvPtPD+MrogJ4it+Z7RIefPM0+IVEZgY+GSRSYC/v1vBOU3SgHbyd5tj2hbzQ/BaxRFL3Un6+1fT
eqQRXwbj5HmV/WXk6zemdcNdShz1iH/fLl30Kr8SUOO9O1RtLWLeIuR85VHx6d4Mj2JHefaLKEsl
rrfrWVo1bC0UUH6KDAy9FzJvlBCfuuB7RUQ4A9FIjhxFf4lwb4H7dJjRdrBaXn4SLDY+DJsnrmZb
7/sVhDOwB+5/mH/+JTkzixsnAVnVwbZDGd6/Pm+LG5WqsFQij5fLBDitS0MGBMg3FNREmVrfaWvJ
ePE6ktFRj1hxGDaRvVWHl74PiWdrFWV9AjoH2WlvdFJqY1OBsztASAnI1MqeslDKomqXqE2K51Ed
wGp1AxpoRlMl9JlpfzS1qaE5+E79ttVGYf+hsWeKxp3F4BKunFkHCKlRNUgA77Lu+gSxZ+6CcE1w
5IstXCYygjLAfKm7M52WajrR5WqRvw89xytFf4W8wUakGRdq7vnd0k4cOs8qyYUIMltqEuZlKXMj
3uYtiL/JUTwWmUk66BApJ/bEluh6BYcfhTomPez4MjGH2yfBCbQ9+d7YFPhpzUxWjxqdhgRRB6KA
YJ5BI385i25akSZinuxfjuPCYI40n5H3DYpWYcs7NvkUkGv6DomIojdQoKImbZg55Np1xyn6iIP0
6kkrDS80SIDQRxqOAVYEmshuDZA9b2vdrkDVePorUjPX1J0l5pE+yRftYrorJTgXYBBk716YM5Vb
Zhw0QFlToasFS45L/ZRnSSVbzEd4JnRGPb3gDYlRn+xtygeHg5jedE79Z7FEogMOJ/SmXf4IVBZs
uoh0ZjQm2arXE4r1eUfFKslXjMm1wHCbNgnpddI+jeWut3z5l8vQ6hBnnieo0OFNJTrMwEQgGNes
TERyk89z7eU/r8STVYsiXDRgviOjdWoCG1ECjqLZSoRf/qRSCxTRFe53t5Can71gd7HRlOq4rN93
XucEdGGDgdAf7XEZScwDgFHPefXucAPZYXdda811TqLM+32I2+wtvcbBU9401R5NMdVQvwTXvkxe
JC+v1CgCnNulKjLMucQpIEZs2YQCLqsHoDgbAtmCgCkfR6q5NA1KTM04X51W+IPFk9WCVfYfJTHI
uR6Z7c6PJ2nesDw1AHS/hHS08/YExyTeeDXQYiZg0OFP5Cz6HNyNDIF/GxS9th6CDH5KAHOuRT08
R0TNztunxnDGDfj8DSwpfy09FHs9RF5fhzSl42qJ1FsN/RmSaJILLG9YdYr7RA5ayC5und8RIbpe
5uQk1b7aWBs7raRV/iq4zA+f1C9qBOtmAWuWsMkj7thcqrzuyNi6XbmoSQXLIt1d2KV6rIfBZ7wQ
XMsybfql/ePMZSMn8T3NIUFcAXsAr1De/f9ZFuSXve3OIaYuiwUuhx2FCO0U63maz9Dw8UvCjURb
ln7yCxXEHfa/FU+E148OYnta+RELI8S9lAMeb0AmbfgaRPYQu+V8XCmkWo+JghFlRawJ0OTOnoKB
73swmk5T1S0StZUwEKKuXriFf7xNuquci2w7lEzcLh6u/ZeIv8hjMrFTG56/XwMEJKO6BSZfIGdP
nu/uZDXBGGD9JBb+fdBpQbK2fKZHzjKsz6bMFOxlZmHIOAm0ScwKwyS3y8kmieDMQL4KDbAmq8KM
kuWvkottWmp2J4CGRYrW/SbXqu0QPAhJHzkmRn9Sx5yiJxecTAF4WIaY1jtrBqzm+BmObROmkEVG
qaas1AXIlGGHx+TNr9cPSyvQPcgam3UGUzlopf77kX36Q7bhaluyG0peSU4hOlKnlR255Sazxraz
yboRdkcTMrsBO67Mn+Qzbig//eaPNknobNZebEUCKH/V4pejlPoBt2tz41P8ycPWEcavMb2Elckx
P43z4BR2cJrQiyx12k/5LNGU2+scS5CBWU6GA+CPXAUBjj3/f+jZkmGA5I0Er88erMC/SngYt2L+
2nsUGni7/iSxpjcOlAvpsgnQAAoX1nf4WdegLbtUFh5aGI+uHqviaTdTpC3grSWSJ0q+t3Kf09Ix
+g1sX1AZ/5apU+5emhOE5WAYsN0mN4spcuuyI1/6BM2pmktLbk0Sbc79oD7xaYXBDPF9xmZhHfYH
oewncpiwB4H8HOGSLLR59i5J7gN+BL15MzvcqGVC6YKzLnzXfU0O+ynUa+et5VkW54gYyiVVHT8+
P0PqTdy8G5ogmFJSovHqQ3ueSYABksCkBb5h+nKdNKYmj0kfmUhL+FniErZafkPiFLHf5NWgz3rt
eaiEVlo7zuS2hsweK6RjV9B3C2f55A+EqvFXeYtTzMdiW6YIMnUi74ZQxymtbvGGcROYztrWGiGv
45wOzfTuryvW7Sn1AeByRl3hfZ+B783x83vQy8isigk734eiZnE1HyhU50ylfQiYUkQJ7yr2a3Ly
2+hTq4hRdPWFOUUMM4z0J8ODWlgV76/1jkqY7ndPh2JJv5MlDiAY2VhmsH8/iZYb0gszpnXfoJNt
wGFdk8WU+X712tFXdHB0vjgfs19DSXvp5WR1AJTA5WdGA9Ydik1/CVsI/PUOhB9mwCjbzRTE14EZ
xsJtB3s0tCzmONlGPDxbBSYoOFNo/8qi39ZIbDQ4obUtG32YHq2hB9aKSxXDLDlaxUkkApjx2Avx
51dxCmGdnB464b+iHRzX9ocQfNT2if3fPAKGnjlceMnMWnWhFVKXbz2qryBEmAQ32EYwa9sXkVsc
YtWCtTv6Si0FKe3r0rhFbCzAx6bxTNkQoNwbcn01k9IZc3N0zb3klGxz6Am2sQ7SfQTEDh597cPD
cYs6q1KYTBjP1CfNqX/z0hErU7Hb3UhusQgO7ZOLlWX/29x4GQ/TQK0J4y6T24uFa4pXBDAjMpmc
UOrK+LrFUFE99viEsIEDgcChRHFBEDCqkczx0E07OZ0e9SmksvKb1A7tj/D4P3ajQmKfdiKrRwsJ
lHcElj3q5i2JZPBNT9EE2lia1B1Fo7rXj06JoLRpAK/leFZccHh1Ac+qo0lkvCgbNEz+ciOnNMIZ
8X6+jb06VuWXI3cKJiCPtnI+QfvX8fq/20v9Wz2pcUNCVK7OtjW2KsO/VyXkLjabwLd7pYWTeGp9
+QNb+HaGnyJuGBv9LyKrr3ARy0AwTHdLfweUbe5c55B3964goBuL6OxtXTBq599HyRxRszb3jNOO
4Wydvc0NA+IHARiBNNwLNP9cWyV0cfEAQWI16LLK6k0EnW46MTROO+pvWCXCA4t2JSomWUEMXICA
oQv5A0ac1tfY9bL7wp8V3l/nXcIwOOIJNnRtM4x9JcZ0dglMD7bojabGICrBWWLGia4EbHCpXqXo
nDiuKyxkIBXQRrHUvU5ieKs0w/R+0mH00Ln7lhusxzNufBvDRuMoIE9Hhf0iOTUHpt+m8CCG/cdV
EzFhV9Hq3D47n6yrLw8N9BbYB505BS6DdwwTWuhOIGuTZI5MiF5y2RMFu92F/IkKSq0IsYDBtj5m
xXeTqjBhzQZXi4QjH+1hweALb2jSDGf9yA5PpKh2ENy1cPfU3sCa1sz8w6v55yKpvgwaYjR582FT
fvxfk1HKw/pqla/rfj7h4kVFB12jNhycxa6ZAOUqakVVWUayCRd/dUY/3mlhVNigetHiF6qCZvEI
UMgZ4AUtvD63hUqBY/kcT4LlpFuz8E13b09hPJj3BoULMunyyTSksDI73YAfy+Vgc8DgcjYzjwjI
sUjxV416sjog8eF/uszi9DM+muedXGUaZw5sBGlHRd03XzyPfYabZYiqZjvx1LJ+y3eVmix7EySW
cvcSvr7h3o5HTIdh7iE2xwJKwM9Of6B4xqGRmNHKe63pfKcRnoqY2NAQlL2DcvqBEWvV6AB5mDqP
ZpOh6a2xOIeyx35LqeT7JvOI8zNqA6v+A/CBkOocApuSLmrJSWSCh+RcWYC1SQsRpoz+iIrI8LeN
w8btaGSB+NocsUNR0kIXmrpoHsc0KYrFSFuupeb6Hz9Wo4MzMNAbAQza5ZtpJ1EbyzvgUJ7w3YXD
zu7/5hieB78EzlgX1pxTQiA6EiFOj78waIRlOY7OKgGgCZ9CYcZ1cPcWLFGQgktUj60h4Rqctyc4
SIZjzdieSFGdgeT+5tV51zGxp93W2Aca/bkXasmJdjk1EDG/GdUdA1x4nYE5q2oXUOCglV6QaWh3
hKultY/+4JPY/pdMFcwBmeUnBvrG6AYIPrj1TVlaaX3SWCzwCRxm9bY+2jEKF8DKloP/4+PB1SCb
P3J76QrHHWyP+l+GsdM2bitgP0n2AdTWp5m/qwxmFIgR7XHnWzATcnFuxXXvmjUPlrwOG2HLYU9N
v4WBxoo/coDgE6uk/OQRVQXiZ4ewYKVYN5Y10Nwv2Sy7bpQ3+aRrpJCe2MRnfRguAhuwxETqd8Mw
yqFC8F+85Vjc2P5vorAVAEDnbLyTv0licGb8i7JKutP4y/bQ+MYe9T4BbNnXvt2fB3qZIfpDu6lh
lxXRo5etW+yClay7RroavnFH7aCTjUyID+owZkNGAj019cDTzvEM89Mfn5tSJH/Uv/T47HgpJxKq
VKzc+Hx4nTe/3vf5hk0Li8uy9htJ1qaOlWYAlB9m6R1wbhRlR2jWWSWbl6VjGWPmyMqtqPgIrHDN
TG/+4AYfeN1htTcQ9HkuZsjttJiPahLYZbicSdpts5t9KIuMSMewNXhXXU+WG4zbQsDZ/U2hyT0i
oraoeAvitGnHmvOq/zdQgD8fBwEHszef+eYMXs95dhFi9PGcAdPfJcjhQzv21f2BYvR5kTvNvVD7
kg+OjOLvynprOD6esqLEVGKcPJQbLE7wjGTiO2bTl8fs/an+Kok/uHuHReBGlADo00M+nXzf/eib
kVqOckXXlRp+po9TwesZwSJHxMCGEOHPr0Art8zBKNnXX/Wz/OvXUPJxRAM4i6aa70JhVKjRqYbV
MToJd5KTrMAuwupp0HP4iB/gnMcR93KSus23koS0jmZz/mY8IBp8QMLXPpwl6SoqcYfoJrWx4opZ
LdQkbEiB9tUlfurI/JWeShtX/gV1bp2qgGhhpyJ+y0A6tbgJwo513I8L8KcmmBSWqtNPwe9Am5is
a3CXRhDzObkldHNm4quAEEc2aAdIHJtPsnqmp0U+4/GLSkZmEnAhz/5lz+w+ljcg94uXv0y/rBPo
WWZ/JIs9hjZwiJuTzU0/O1x6vgIzBQODJrBXMVcPTsPW5CRgXelM+w3gCA+U4wY+a3jsaNmeIFua
UIGIKeERhJJG9KgAeGZfos1/Q5Qv6gv3o9XOkh2zQd8qZw1aJDorYInXxt7rgau3UCyylYo5fm4P
WGo5P8F4MLI654mHrV7wRwaRwFkpCO+ZACKLx6Hhfuz6FPgo2ZsENhwrkR4uHgoIZJ/UbWGUVVlG
5M1W4Vd6UUxYj0+lGtQe1a4yp7jZbbW0ZE73i/+QHUEWg1WVIjaJlRqJ2d35vTXCe4bSo3nkj4HP
L1xstDDo9rqhaAqEd2pXUlzqBV/D78WBubVbRNeOark7+37cM5tq0tZg+OfBzjpXynNevOhIx9Eu
7uy5wDRNAQXIJtnHFskIOfpW4cHqfHkKFsDFFCfdhfJimr+TcfQ52hL2JPsV6Ra/YayJ0E1aqnpD
aWRGZV4I05ahWDdQsUWu3Fc+2bAfpGstOxnqMcJtHstu4tesTA1WZBIIgURWSctyWaRRkoiSPb9z
8E/tLLM6AkV1KWzjS5+WjdCY5BsgPVb/pC96oB4S/g5NX7ATx6rNIWelGetIPIWtgLOu5Vt9/E1R
14HIG78ppLnN7vYzvqDkDh2jd2xNqk95LSf13l7CM9JXX0YuflFa4TCtXWZ2rBiguohv0M1jxPJG
jRz0+F8peEc4Ne5JbEpN/IF60/1YTdjqZ0TR9gx1KHbG5ENoLBJHV2WXKjcsJzwMLIozqxeyov2I
xbXAkNN+HQintlJD4Hga7bgpK7pDDEE0ippE1eMReHu07JrbFJX318ST2eK+pS62P8ZDxZsag2yn
KcQs3En0Viwi6WZnDtL/q54aruIjfAa1WJnLCGw511WafQEf2Xx5aaaqwRep9ya1unmPtShKz2MG
iy6r44eXOxrZie0dJUQydsK8t8R8KLMETPt4FlQvQoKWqjTkkc3eu0l/9TdeasKzN4GHMqdz6+er
j4cpe98sYz5unooY3NK9vH5cQaM0E6nTcSmo/hL0y0tCEZ9rGYLRSH7NBJvUZgF5uyT0jZJbeLcB
5BHzia/VbAxWC4Tl+fINc9Vxjl/oq0WB/l/KRMRAOdE3rnVDQxQchs3mLzOaT+gfv1MxCFx5NnpL
TEdXiLZQwEBBsmz4CTuj/gBeKUco3mProPz68AsWFzf5GJKzsu27hKwjEBlF87bb4WvrPBhtTiE1
CFfUqmKreBv6ApEeqFEhciDTyhkxHlxfLefAZmf82ebqW5G+exVPHhVDAJwfIoWyza3ingxUS+Ni
d0/5sSgUTPCJ5XIKDr8oIvcf8XgMSh6MQlhyygx6fm+QQNiwXY2XH4nmTCq9HeqEjJEKIeOwxXpk
X+FRelA6qY+qn5wRRQ4OKUUgeXV7f/LC1JQyEY8FDvNNy59/nH+8VO70S4FdbHkvlXHLfvWUjfC7
u2PuL3Z9OKLdF20Re+1r7WvOJkO3K0Q5Ar0WL4ah3rt1eh4cuznlWXtTUxIWHoAUY73VE4IWjnEc
snTwep3oQ2d3pVBW+o0T7TNm4sidt8ZzoMnugOVMMlpFgVP4YVH3e25ncu2syP/MmYyxA3V0GSy1
jtkluI9Fm6LMINZik3zUOlUB5P+Iw12ORtEe0c3Fe+y9HIwVEiypftTs1dlS3rLalWSySk4KioQN
gS5dckbC+eOjNXfiAfBu/BDOYsC2Cq68f7PiuIWTCnF/dEfPZ43enk/ugFwLA6ZsaL3+b5krDnUc
S4dONk3LeuV89MTcmpgEKBG6zlF1GroEsggax/Fx7L7q6OhRyStYKA5BlyAkSizB2B7lLb8eMxLF
IBdm5tXTmwa0c/YhYYKN7C0OeTSfTeZZbXaJeJG0SSNtdWfbtNaX4VXPMJE5DSR+tYjdKoYEoSIZ
20kfGpYSAdDbuUiYWcm3UWY0TsnWH+vhX7DhUzvpNnjD7+OFAI0z56jwvTUXUPbxXg085LOHEAyQ
b3v2qnwDujMj0EngX0BgTQw/CltQrO26T+EKDfx8Lpw4R9VodffHIXpeXYoEBX+vzbAJccWlgriQ
zdEQPxXNZfXKtASYiTCRtfyYyD4r1OIbPn6LqxbGn5T2TZpQEOQ/ZqYnR66iM1v/wbbxVfpQUT/x
QAkeKM6HTStG86dUzeDodE12Ce7Kf7PkEaQVGPYL6+e5WyKNf0s/MRRc5sHiwzUiuXNSfskbZBTn
55oVgN8CQp8ndTbN1+nQBXqLn0H49NZ7XLhRvK4bBinUkav8KuoESx756/eid0Y8spNiYU2SSigD
QpeyAXofw17lFW+7pF2xnjWVFv+eLeoTonx9ydCaYdV+SL895M8atLuXsK6hhtkS6SrdSJu6yJat
/6/FqYKMQYRq+XJFknnLHZ6//mHcxYYpkoes5j+/eQwPsZVUlyLSQKE7pEYvYpoY4x2Do/p46wTY
l361ySGWvTPDBYWXGdy0Zum2cor/rfQBPeyJUS/BMWfSgsdeIIyqOUWjHGu1fsVC79dOQ1MNL/Bd
QQo7RYDZVBXTSc6AiZyEsW4i4wNCsIlIBhVaKJlt7XI12FBv1bbeGsu58CUJLWZ8VyGgl4P1fLBT
PpLnFZFq6tR+cY97bgTybVzz+8iDFDUQXy1ZB2aKDM3xPIPL3zNRzJOrq9A9OQh78X+fYYuHgVNF
qdw5sIC9x1zvC1IRXrqESduTIhOIIRirDKBkFx4TnQPSWSqNkiYIBI95zLrVrVH5Z9LXX1oWB4d1
tFputQj3W03Oqj1qQy8uDZHDHmJlZ8LsbhYjSCUjrBGVEzpj8RY6bFOyJFUKiA4c4byIjZMJ+Cok
ViRHqjCeKvs7nbulyKVq3AOmL0T+Ph78Wloxj5Xg53Z4pcXsmgzv1NbhW6kBzcjo/74DCSV52Onq
klm0r4rra1rdGWpIia2TeR3wPZDPl8MPSdr3IqaFYO31EDkrKNlNqzPF1mKM6dlS21tbOAz8pQxq
6ZaBch2b5qD8SCfwWtnHdegqdU0iIzzxeVx4wXKvYsN+N2pkLBOdUwE8jUcOKkMSdDTSc00hf0Pe
suydA93j7fyjb+bk/3fc3ZgmuaIYSvwZpA1sOVkZx5rOEvVS2pMHHytcQ50PNi2vwmet3nkHVADK
Yam3GSSRapAQ4HVLLaMisherrToSRZsuPrdvVQASKvo0plPGQ50hgEs1MAHt2xjZGKQNZswmcjDn
6JOhOYMLIzbBjvHA7dp8AsVIpbH9tU8SHhuqq2iVLuibB/yLuuvuZtbMponnY7HywvZY1iHdnDHY
B4Xeh6bRzGCLcPZm5AXdicSiFg5rlwG7kbKeMFQF5Zj4EdQHXWl19W3AfxA400dfUPf7gwSe/BIJ
qp4ODvGxoLXwE1e5I85IUJV24qibD0O3sw0k4xCu44E2mudurjQkgXkWsYq3t2Crc2yiE9nOgzDT
SF29+XP+yzHeTGGfQBISc8Slj3mvDxWoRcumdTig17MEUZgF5Q44KYyuAMrvmIBatCgCBinSNcxf
MpTZ+o5nIBTEF/6GC+N6CIB+PK54PPWIkz9ru1tyOaj2IKb5TzwfgcstgwWqDXOszZhF+ak3YB6m
hqyJhR+BqU8JAQ3VfN2puuB9vQwfmuJ8/gArQH3ilV3s8R4LTdHQu2VY7I5IpOWCbJjfq95RJ2Cg
QkSsLYnxo+g5C47TvGErKeo6GSY1IoJ3fxweKru1rSnoubrn7X3De745iYrqQX25b9zTA30jaIAh
iSPQTFKsZq+DcFA3OiWVIi2/x40NWIMesFld/oYrqSVfwvu7IYVfj5IPzJanI1rXWhkxv1cNw7m7
gPlRIBdKbSCokVUwHQVsS9Ua6RHKDLTmOlVnCdjEsSNmipfoQNh2uHi4dhOYZu+My/1/CU1b4vRK
Q+EbSrjIqtctj9/lafd/7Ki1h0oN1ZskmHtU8zNEklF4EZiXRqmgLbQyxAwVr5GH31ZGnqlfToOB
irjssZX8f5eNp/oPaK1S1qI8EEkEck1OeKOHzOrnQ/KosDiKGh7hHSUKlGQzLEvjTwTvXqFMFq7I
dgzg0o8nyHjiahi/wRnEMQYYX+a5Px4Zc/7FzGDNmzstr9bQjEr7MsN4lKOIlroXFxhT0lbcNxui
sc+rdPayOzgsTVpBh6WftDdzi9VdM3Z4XCZwGIEAL91GI8Xh1Xol27qQ092H4WBemfqVWm+6fIQM
jdBBnqjwURgwzrX3wcVsQRiOEkBk3Jn014/GLwW7DLn5hQzEp6v5XT8gmOzeqpn3u5V7+qpWN5mJ
mz4y3wGWMSrUagH+ggAjjbNqdd8ASihwCub8RPX0LdZUciGhpJPNK58xT1LxCFnLmCqEGVxVKKGz
BYbjkjDAHztv8Ac8Nv2cMBoj0lsYOwaotGqtIyMYEfiYsybkVFbvSo0+j8Gu+zG/XBeiZ38nTAa3
q8MXcMObr0opR7w4gUcWlkwyGcm2UYfvvw5UgfFSoOF6SyBhWIpyocxgykSFRMzSbKHsW8zAbuJp
r6e2x37NGcnz6is3Bd9irimzr/3fsVKEagOUCwS3B/tO5dhhB3iYqqYJ/3yvUcoUXJpAY3wdjrBd
fDEZEjTPavk69VtqmBYHn6co+pS3ENxlbL0whePobEBGvE7nutatXmcFXiZLGWHEDicR7+mrhlaq
ABwKUHDUPbyA5qLjr/XzjmqVEgQG47UnohJ6xDSjVDj/r/CDqcPiyYV6x+lNZScc5bkh2l7H3pCX
xwbsxOcl4w4CkZLxT948yvq3dU+kpb+flRsDoRaASNJ/N77RbKdNPPXyBdV/wI6r1SmcEHqa9q3/
QA1MZPN+iqRj7/koLhBVR8h1b81QFI6dxkcGDjvfjdapCSoMReOhYRg/5Om300ZRDkHHkfY2f69R
9gZJTSi/n5nY2M28CDkmbQ853W2hqzv5pvmpefwbjtEIAm9jcxtFG8dTNKy1FCJD0F7GyykR8s1m
t8hDPgi3Ejd4GXsONdH/ujcYoEsgTe4Jwr24DaK0Dn+/P9yWQZePNfOw1w/Xh0buu2lp1XxCm/uV
4GwjmN9lW8rpGd2aUJ37Rp1XcZTH+xDGSf7+MTim+rkRVSprxMgxQrTKcG9hoggNzkgG8RSxm0E0
jSm3dhXR4P3hfhRio2VDglmbLK4Q+SXfgQscfubP54q6E8kZhVEkwRCM/x6UuMlUSuajhZ+q6rls
B0c6g6hqKwZltNa/tImm52xwB7HAhxF0iXa4JlzSid61rzGmlV6TyzT98vBlIML6kVTwLWSO1lyn
RbExkSS9gn5VUyUrUH5GJK7gJQlWOZwbJcW+U4g7j3AKgSoKaEdYjgZHRwfwD1PyIOVDyYJEYfed
f/ut5oHVG3CrUqh0j2+zxQyafo+e/d0DBCucmlCbssHWrP84dBB9B576ulxTn1uNVsCphHq5FHPA
z/MCC3u3qoWgdADKriq0TFfVzdE6MYefJAWJZblDRtV1wllNt2ZnnWYioSQwzpqajxV7gQhtYiJf
tfmwIgiOAFOxbj4MmNXcg7oQXOq6Pj/8QobWZUfUhG6Y/xm7Oq9T2LcyIzviejwMgAcasaH876eR
s9cHisCLDenQRAiSzXO8tz0DmOuf62Jer+L7XB3wcaFyZnYJdGEa8qv09oxzOBvL5y9WKt5OFaXf
XyLq4w0L18a/mSYpty1Pw5Q2D1wy7TiGR7WwdUm3ji4iLkqHx+BJcQyOKYUQYBecJ3q7NV60lGni
eT/I4705ayXTliSRNYnKe9oqWgA1c87Dj/FU7Ifbs7/oJZnbMQy5soKbxV03z9w+TW1nx2QF3xZK
T5TYaUqqcJ9RIDDmTV94ip9BfeQWPkL5rE5d+ZpiWsVMVAn2NZ989UqNmCmYyVEUzeg25tRno7dU
0iGmizkNKPZnpxBpfcEDNlg1wSGdveXYfIyViOX59GwKqtjK/a7+MG/ZF+LHz8VFYKJdGdroKcYN
X9JAKKlCQTqPWjI/U2pBinqO1l1L1wn2pu5cs9lQ7qRqoFmtnPrdRYRflPsgSO0BWxzlgQuXZmr5
7vTysA9RUpoHdvKri2IhLgO6gYPzxco8/kLTXQAzVqHUYn95staujBjJnJZyuafcojVrS3TLxjML
BpkGQ7a13I3GZrYkTNF4GR2mWwznN5+7BPSa51z0Kd9sZY2tMAF9sBT+X3dYuL+ryQq4ggPx4MXs
gndsqbfNb4YUwnPIHwNJRyaV9qTsDlHP0rqqd0I6G3kRgwbsXmz3qDQh7PV4W+QT3hoggTdbYLwh
MWgsuNespXDFNQFWpd1fGJq5PtnF80TOrQV/tX5t0cMyf4gZYde7S7gh1E6Wmc8Nxhe2BDPywLJR
uPmZ5yP+zSp1d0Nxly/yF+cREIUt8/yVXrk2la2oLzBvYkcWK2liTVKT1xpFucKSkue9y2dLSBVc
jld1XxxiUylCyxwfZCz6UJdXXU0cXucvTHNpX9bBqoQktwu41+3Q2rLpDrAf0DjLjTl2PWShAhir
XrBYUklTmSRfe1beRh8QTCtlnHkh7ui7cGESVMDNtm9SK8EtBsMA0DevlZbhuZE2ETAfgDaTLcyY
m+EkWP2OuUhlUO+SbofILfueY0rR/KtrItbPLPNzKFZSnaFFi32PeUZTRQNcyqDs1G/cdRA2iTu7
1VXf9+mJhV7miyfhVo2ZOT3CGyD3rom0hUx68C4r+Zl5Y+IEwFdLVoB4WIvjI5qyCSyuQngcP+FK
NzZn61dL5RfyFcnpTqZbRhvoHIIW1bt66/rFsmg3l1xH80JVISsxSEwZ3kLxfk51FGMGiLKaoKm1
7pONHfMmRpI4nlh6Pi9xEOjHlteo4KBeukASkQ1eJeGRHmEqU+p/0VNRsoi1uK+2B0FY3zghXjyM
IeX3Gpke4B0QG5laVBw4W+zEndzBhNgBasSxFQ916C/BUN925MWOwKkv6ngXyh6tLHaDxe/6kmDj
ix7MSQkLKoHz5DmScT5fR3JPNdMQWZZUNp/IcCya8oF44SylT7ow2y4Ej4qen6Rq5UP322uppb3n
K24+YoIycxkDEHiUIT3AeNqY5xm7xXGc+8yl4+68mcQMwClx8qN8TxTvZ+uTecIkWUYHmqA8OSPo
DLPioMu3gjCXQs35QuqqTaktPGqob6AsRus83UiPvDmxwNTqgFhjMOQhaDrbcro2hirXd3HWbuX4
OQgLSzJjPRvHE2uM7co56jUtCAcswk5edU7uiP6GkN6PH3oFEcayfahmZ7SjoVBLIFZzsTP0ZX1L
B2lBAeXJzxvKGBStRZHz/MAPX7WUL0nhTSuHk+M43E8ZvvZT+xMOAJSvokvVthJoaoSuFV8+IIv3
aVXdMs3GZe61Po16LOvqhrwL9hJHrrqkuno8viGO7Y2JCHzHRnDOo4XpG87pVasSooVVOchta8H3
eUjhnUzTE5UPNFuZ7FKYFgJznKN0R2Poxfs+PPLuzb1hbWonMQuudi+OXIC47z7dgQleqrRqFJie
zkcKHHbY54iSzUyesrPCS3IE8FU0IfjIzRalIZofW8KHnYQjQC9aHEpTWGSsVdEFeViX+yPPhFSQ
uX7sIs2nKPIMSTd19xdenky8/FRKRTdqJI/OIWGfnUIJT23lv7tNSlEkRPq65RuMzCHc05TJHg4H
n1JzGuVmm9hhokwl6VBhA0z5W7DsRke8QtFrVDhGsDy0LEQD7WFyF0cME+I03/k1gLpC1AUixh3S
Th2hz2/WiPrWfjn3YKlq5XnFku0oVcKMl3YxjX5OahRV8JOQCAfkUngma/vTZsUSwLe/jn2eCg2v
puKSr01inJIQXeypqrNzdFe8J4w2KhgQz2DDzAjyp069QGTmodS8DFg/06amSM3Xrl6ON0tGgVB/
PIak6rh8vMgv+gqZ89fxBbGsUyBaI5xPEW5+7wshUwdv6yPEkVuPVMfW+bfEURhc6fn0IkY2sMLf
IwxVZvTKtTxv1gJUqYRk0Gku0Kt3af8rfEYAVaZ+Pj5EoZMgTee8znbSfDbbKBqHw7YZnkmyhYxM
JFFADYMN6jA4zBQCx8GMKO2P98zCrYzO9LYLCW6/P0rWH6eE4DazpTAJD4O9x/1p1vhR+sPgZqxI
nupZ10lDWV/L0ZbASvBiPCpEpxUUV0J1GIU241/hG8Gu1wBqhCbU/sMNwa/O/xf8vzJgXG2uvr7l
Ae1mxjDUb6nK/LOW1oe1HrCTOHCH2GFAe2j4bOIkJfUCNnnl9lKY4O/EXUz61udhfOiCHk/SKTZ5
2zMgbeRt1OpNYFMQ66BwNyKKuuTwdvxBRUp+Np3ApD0p/pCDrOfyAm1i8Romly5N/KFMqaDCiiyX
/6EwsC/p+Sj7EBLGpFFDwReodzA6JGP2svOCZHrmGOwJwJDRn5kgk6se31UnaocvDVQFjiI3qOfO
EhvGANrpx2bwgIsTb8Ht8WC6FJBBnLxShxH69lyNauPNdAIZR0ar1ZMcZrsVya4kHUrA2bFzl9MG
GGdDfaF1WSJiwpd1QtUBJRXtsXaFSHsLDfYGA7FGNTqUp6Nj/iNo2fCK3U0PhXa4tK0oh3hsETwM
4xK92JGSXzIqZ77gm5K6tonzXIeOPNN5gYgAIXpFy4oUlX2X5uA+TkXAy33dB5pd8MDxWqDD6ncy
l9hT6kTZycz0PVuVF2xZqbie8kJn8xnBSa/N73OufHKyH5SvWRmWHkscaTjHrSwF4NTvc1Xy8kih
OooV1UFppv6oU18t+nGPbDc0+bfxRUZd3m2B547GFMmmV6Nc0jlQ4hObDm2DUZSDh47EI6DGs03F
+YbhKVU6JaoGKT175xqaboFKZXdQ69bWWetuZ7ClS6M22t1teGrreEkYZn1dUo5OH2kgz4NwBryS
ijSnXjk4VkZKWqX7LHzqBhLHm1rM+q74jiuLUSHiNy6HQcWvkSQISZfGfRDdKHhOYjXopkMtSTTP
US8YtlNXyWatrQam5NQ464vGUIJ2tREwLD47syvNKyH4ONQE0fgJU6mERWoZe3vQczPW16I7cTHT
qOQX+jY1JFjKIVlxV4VQlaDOizsiMj4BstivqPbOTVWzvQrgojTzwJCVT79JJW7s7vKFM19/xDGv
yIWb2R0xRe8+zRIXoeEQWVZgSrlqa+pScB8vX0pMGGQoCbLIRpQyUFsjX2msMckEAGnwl6ALSTwi
RNS9VYvsjLy1uqay/bGozgwZa4peaok3na/bLUgQJ3C1UFSLlmpSunPWOZMwZqw5wENdG79XQj8I
YE+XsJ2+nUu/Z2RATY8toVBVl5YG9s3ohU0G1RLNxS2k+It64s3YkamVq9wf4aCdN4oXAQMbGdit
y/aYqaNRUW1uMsCFVk76jooJGDEETLoYPZ1SHUERJ4QyTMp9ZDZ1HqAJ55HMMCuunzE+oqNNWeKA
YmrcEXKkXzG8qSwRlO0dHGDekCridwW5OoCevA8F31aZf64opK+3BDQA2V4cZCIM663jyyR7WOy0
xOUDX+yUR0gmokm356tZnj9MT9H6zb2bleBcJRPu2LBvs//bgYnLfdtHNydHRU9f3hKidOYfJ5ov
mW3KXUPQn6XBSWj8kLri80XvJV88R5/W2BWIo0Q2h/BjreE41w7Vkk6D+v9s082KvphFSM1ihf/V
GZzeZg99tuOxgGbvV16K6LbPO1ZMoSUhdzR8esDyhLqQ8xIqbfQNhjhLoQJqAAVpFFriOc4M8oHs
xmXTMHYShQBEAZ7av/HoS77KQvf7O+ip5Fopx5TnU7fWGMxGjf4/+J7IfFiGH4wy0nlacSDD7GNA
h/j+6LFrNbfrTvK16E00rySUm7e3OJRaKUQNY1YxPQScaoajs7ybhlh+Oe1VoGD/k0ibxq8b/6RS
6O/WXWrv+TA8q0YdfaOrr4Qun6b1LruF4qX2Ox5O/oJxc3FIiQPDmF4JzwpldOoEK0iBvm15GnA4
HZS6Wwxd0jcVNBnbWrEZ/Zo7J3zU0aKf5SvwiDw166ECKUsZsAk2KhhuPCvDgmWgZb4xW0z1ac7k
K2XeYe2Zwvia6CYizdxKR71fY4KCsJnUWJsl4aKstql6R6fq1YzUNCbY+I7LFrl1Jjj9KIvJghvk
B/Pu5K7KZQnf37k89g5rcc7fFxDL4lhDs6tqy9M+L6HxVZNHlnKU3j5z0sEsYQG8P7NnMvOCGZEB
Y5FBBY+BxL3uyGUbVPaQykRFslpVZ0d5imzgq4G15zEe8Bx2tiwned8ocCqz+EbazjacJIMUR1nc
FKOeWOLwQPRmH0V7w74jbyzxIb6z/iRbnRl4QjO91OJAg3FXMXGtRkMvCpJ4vml72vaY7LKeOcE8
Y0UGKrQU6VB70V3WRxPucd/hcp680bhpXimFsZsf7iDA1Ypu59Ku+njoRklxqp84UU9A4YoiT4kL
EhMR21qn6sKwRWr59xwDVv4wRsn+iSLq49ttvKNzWP42M6KlyHonDXI8yADug3Gv6ygomm0CqWD2
jTk835mkvuQGcObmXKi0TS6DR2S9M2+9mKHzCIEfv3cQxXx/MPkt+FjZdXQ5x0nwxcESiLFFHWyB
MwaH0Rbninhggw26cpKtqNwVE2hRlT2TpTSHjMW/cZjznzlM6l1K7mfYwEr8k+sG0PqoAborZnj/
sR6ml60KSHbYZ5Ubp5yvyGFgHlIE+20dO+u5XrUOMba8htkAlBQA1cjII+DnVsBwqltpXQ2peHNI
nbimdiW4HgVdASPfzAjynxVly2oMJlyQ8BCa+lLxx336LTgQQa+4T0oBFPJ2hrYgFAXf9mdZghje
mjKYJIz+Z9qz52NKztbXNheOQQbZcmbLQ2sLDdh944CZPhhSVQgrsTCXmr2EhLn0izIMwBicZWBk
8Sh/TWlQkxi0YfgNg7hWcOrWC+qeeyOx9zuxMHFYDzl89xXTHgFStOz4/jv+NgOhfWjIyqq+QkTE
vprSqSYMte5rDg+k9JzNyHJmcgOENk7G3+ePXKxi8rwOnhGLwX954mG9ybNSgV79Z1JnxGTXOxRA
hNHnhtkk4hM6ZTxukkn6A8h19Ri0jcj5qBrj1mOs/Uq6gH+4Cmcghs8hPpZvCkPZOcKqRN5AKkwy
SR1c5Eg22RN6iMbUZEo1jH52pt6pf2lBkB6T7Vmn97ZvD8BFMpAbIwtlamB6GxwuERkhxWEMszjQ
QHjDTWjBeega7XaAIqG3XCmNY/5WZ1YmQdpN9g0w5bpbqBAIr3f110rXWWHTdD+CNCp7+cQxhpPN
IMPCSuaiBkRHLOcovGNfbZ5CQliqhEusHHEtrPGzK4t6HGCz+hUUSClj+JlgVKhoRIi2kbFuCP1X
mMgvBbj+oNOXTJR8eHObfgc0O20qVYNLrSBVblXa/ch7I1Epr2rbQOfFswCjMcUGxh7tQoo0nG7I
Mwhev9qoHVj1FQm4Bvraby6Q8lekNadzSFvIshXlD8VcrqICLi5sUrAY7TG7vaKifJNDXbz0TAwB
wfs2da+ojHAjgub+51wi23kj95sxlCiF+0b3YQhF3PFgOL0mcws7PRRBCOjftUsrjmYdga2nrb/m
XeQQhNl3jlIXnCTI+uM4F6wj41dh7fDTRQa2AT90NHQmW5lbe82MKmxs9dZJgT33BzqVYfbdQndi
4PHk9FUMHVGIVq2d5TIrRHIGx7U+KGI7yEaGva+oqXik/UD7BRNAfq+EmokJveGe0PQ0WEDnOxHc
CBdfYINy1EGw5obtisEeY4Jq0qLYGq8XjnhgelhCWmwrbHharuzA0ForQXUcJ513zxbHyYj8RXvF
rTQrsCGfaR6z+kOKwSEVtlGXrnExVABIgQK/AguVL8jLtCuMddgQR6SqRYJANpfKaWn4PzIPZwja
nUKxDkwCDAJrHDFUK2TON4I2fB1/bYviUIb/jdimCAmyLAu8JwFGasQwaxapIO1Md3zvlGQ4wQm/
FBg/0Et9a9iE/IlvzPioBUxaJ/jPTdBP0hhWHmFoz3dYluvf7H0cZkg2fQsUbL3NCSJ2vYi1sUvS
9AG7wbFSEAtiudxqR2DdAJx1dOzfCzWz9/4NbSmiVWGT5roE+NRAS3DDU7epd04yHBJN/ZucUf7u
QrYiUDvFGHxqDLm4koJugM0imZgJ/9lHrfp1hNeO4k8L2V+F8NeNAR/ND3+YEjPbcK6yHNydbxVD
PvUJw/4uw93Lwe2Ri9tYsZfNmk1kkzMwFhe+TjpJBHKAvINgMP612QUVpw8+ZHHz1dAyzXyNNdUM
E7PyIn9A/FThqFKNAVRf6050tsic2jHGevYSUNU7b16IzIk23wHdzvIdLg5JM6A8QaoDExfT3JU0
fMuHTFUnobesR2070Upsvc7KA10Xz/Y6Uq0367xkUxAa/LbVwq1pne7ir/tfia7+Eqncp87il36q
lz8bPu6a3n9e47bl2W73OalyzEtZhRkje5S3kOYjOR3aSXy4df/Kg8ynXNfOVVN6+IhZ6tzt6ZzB
uRva/LM54PHYF0QI+jUp9A4he0oGzv0crwRFZv5ZBjX17cn2i0aTkvLTz6Le+zI8Q12kteNmR9Gk
iwFZKXf+gUQqCEtnOkaiyR8im3qJV3IR3y4Da74kFciCK5NLdRC68Pf3u8Uj7kaAfkyb8QMJgoWm
hBr75nL4hssQXN3sc5j2bsW8ITophpUo78vUJRZY9fyn3z7IaZ+SxsiagpFb3M10Uj4WrcN6QASH
+pmBygSWFlZgUu5DU3HtoXKIT5/kpfZR5vPDJjWd9mM8kwX/4BL6GmW5p+0UM8ynXRnTf+YaF36Z
1WVNurCJcabad1VLxzXo4vSIQl2LfeaaJT1e3g3a6ESMY/1zQJZcHKWWPx1PyHjYLElxMPJu/hWJ
TuB8boxL1rnuHKFXJzQfRGQ5ayil+9BLI8qaKUEZpyXGNKZ862XYuLF2XLGsB1vbxCXlyfeOSRDs
qFH3COW9to+IuS2v4nWYTZSz7qGaiyEJIk4wzfKGm09nhaOcPScFd9UNdzxNFOXM/17yEy8QlUre
1paqtuFwyIDLLa9DEvI5fItZamIiJ9QuDOyq30RXi5ToQJJBvw+sMRkqdKb/7gb++aIApYrg5a9G
uwU3hmUHJ+QUG4faN9Z16vboV+YHxsarHCXGuKe81L636ZpNd6gBv+nFhgjA/XNhwPYTQHk5pUFS
jT0Yp4ATYUQgdbQJov2Ryl7jvnhfVp1IDtio6sSjHhDfTAGwjsObuj5yPegdMJa+7nbyyxYFfRe2
4e4gGaJgYb2x39D46rSFuctFKhzXfvJwmcsKueuOm3yBG/s+1RIrBT9vK39rrXXp1k3ikyYdzgIJ
106njdj0X1WHRsVbQw3uPYvzZMUZw7MEjj4FO6VBVOlEWW8ZZfXiXcdTad3bXfNWWGcURTh8SGh/
XKwolexmH3Bc7LQV2Wf42aR27b0PEQo3aQduboflDTeEtn7DKitzi3+2xT7k5kJ2gOen6tqCVnoW
uH3++asd02+y+jUxe+wX187JIn8TAxGksgKNzPD7q0xsI/8FMrqs8vK31x3zZQDIhvCI2FKZIZeo
UpRKDNu8d633mjI/w3YC0zRF5t4lJ0zIKoTBfiAmPNOfYRJJbae8UDfX25XT8LCXcPXACSdaKaBb
ELljKD3cZI+DEIyB3bFEKyGwMXBiKhH2VnsWcqwHmyef9Eldzj+sb6zNmsLImuf0vUfu6/v2dOwe
qdT+uMMKFJSOfl7ckjOHBkvtdanv8RSpY1SGDDYjHk3MGDlls3CwIGzwo5oyOl/g5NMlHGRv0g6V
shMGnZU+b/CVtsQaEwiuZbbn5UqHeALFSIvYntBpYVCqzE385Z8NMMVeJIbV2jcsdp0bJ6s1P/Ki
IsmwPADeq9zdO4eZjqP2uhujtUsgNU4py6IpClfYIiNQVCtXhJFx59KXHyY1q7IcJpdsfPmW0PXE
iKRyJ3+SqhNzGl+l6Gf6Qn63jwWuCYxF8gCYy1V7631oH8AveUuFit/rwyo4hNAwLFfNTj31N65H
vaSGql3X5aB1NsghSyB9JFXjCKcBY1bxFEcVpO3pgIT3M0/c4ibCC/us/xIQhMPljusWvpgauRBM
H3hfmFywAjOFbUEMklBzHEAIuzQTxyWLeiUiIs3J6FcEO6SvXiYiM7WsRTb/XWCChKCf5iNnmoZy
cIX+xxf9xNIuCWGB3HXtC92WI5cuASQIFfQN2ulXTOpKJFi4shsgs2Vo/7mnyqnjPIdbyUyEyfrd
qwlhxEASnVaZ20qGpN283CLDT1cwJkTJL70N5Om1lV0phHzsqJCCIcRAH8Q0/v1q6tKg8VbqdcUc
2ZCrjVmES3dsJDeLImjW9R+u03WmORy7dIHFL1n3GuFxJc6u3r+FmZIf8uVdLs81NRvxtTj9/TSn
UJEZTgapQCBQZH6XLwrNy2U3WKZDLvZrHgIa1g7cTfYAc57cXj6rMNidOzwCsd9EHn1BnpbkgcuI
ZajdmNdbe2uF6Zz4DR6VOW06QW4fHoBTgxT7/1BGEkylv+jIaDjSq/gItUE3nATq9XZN8To4/B0V
D86EpPeAuN+BwRTb4BvAPOugadhtNJ+JB739z4yLZZLt0t4BXQcJUxH6lAJqTogxEKC+Zqz79sHd
koPCo3QbpKluipex4TvtTRjyi7Y6gEbo6rkh+I9F0WxYl1N9acqttxUSId2pmqhsPHNYMr+27b28
PXFB71sRkEx6HhyRGe/76o/rz4X01ctVj36Ve4hB7mDxerqY3UBcpNxQs7IRgzUBRlKUHhMnisO6
h0f/WMaufd70s0NL3/3DeNylFvzuPzBHWxmbAvBmgvq4dEs73sAXYLmDgrIqcXtTjC+bUKZ4VDQk
1FYHxYngw021kTsZSI6YPhNCGrW85Fr3x1n3VpDCEH7b0aANvkDFsPnuSxg2c9FqnEjUctp4IMPC
HyxrvRdLs8bemoYhRrjmdmvxHCz2bw3Lc5OJK3VHJCKMz/tfNypm4p8zdodskW8np0EF2AzDAe8Z
cTacJPl4OnLRb4v1NhBFv9vGFkCQ8qWrFuQM0QFmzN/sz5l+mpcMHeK1YKF6ydqCuww9cjJ6UxHo
a/H3Y0g+6ipwbG23qVxy75QQL6lvRgcVD0G9SsDGL1fmk6wmIY0T5F93CTbaAmzqw0PclSVcP+en
THAbAF16sl2v2BwQr8IpsB+4scmuaNL/3w3PkWN+9k0ttztKMuNTKT0Z7dJF3nKNpLo1FtxLv0sa
N9MFsO4+4LLk6pcxl4AnBkNycUjQ9VYAZOx4WXmp+MWu2Lw+ZiFa32LQ9RFoydHkMPbvpOOjeVzU
L+nI489PHHjrI/2yR0da83CHf4NYkYWfFTIljgnJ9/fh2O2DwjV4jFEECTrn8y5Wyl+6fTT9ijLm
npypNqpjFBjDN/25pYwAs4efddCNaPrA3YtMGxIAXlEw9qQu3/tYnGbtknuclfoeBBzBRCj1gd8O
TnjK8oQoWUGdx0W6C8Nqr7aX30d0APgoqyVs5zIZeewYSpccWQXuqi5Wn6ITFMj8iTeMT/ka36lH
DzlHUtYiX4YAbMCKUj4mC50360kSlTiZn+tgcvg/K67ujpA4TMCQT/GFzdxjooPD04j6NMGPSD2z
GZrKXr6wczC80qbuhuri6ENKVkuJfWCfQ1icqh5Ewj2QYXTazq2lj9WZABCxivbCMEHzXcyd1ZWb
CXe8NG/VApIJERQV9AIDVVvH5sWDZe1wxB4fH4jlKKNS4cJchI5PZ1hqn3jCfDH0zYqEg3btPk81
31FK5qMCnQmJvQs/QIPBX57RIg3qTORCccABPFnzu4Q0LlHBwgtEOEiUOYXT18QcPTO/HWa41tAE
8TAc038HcwqCgN/TUAzQEUD5CDwGlcb/soPlfTsmGyu4z2emPZ0oa+MtHOxdzrKBNn4/ysRNBGCK
7BrMKQnXR/NOsw3hu/Yspkz02BtBTunnylLk0QQG4vyMH8EbJhw8aISRlp7tEMKxzhW7AQUbV0/g
TLB67m8onbqDP7QewV+v6f70h+aPX5mMj8IP9C/+QYc3ez3nFMPhyxKoSO07UrvvYWk2xvQVm8DL
QFh1PQVsw3Pbi70Sj4g1sku/tStiW5CREMEv/pqDWKiQpyGcm/X3mO6icadOZmVIv3d1WgNorZKk
5clhKj9kGA5W062J7D3j0gQPf2MEJzDvXgX4OGbcNmcdKVn/j+/csyS/YvKdk7FteLk+PPQ4RmwA
sRGxmLbtrM4OWZkhW8Ux8yKn//AwVgYzKCj1BxUKaV1DAwzZdgnLSwutagXqsGTK/iACpOIZwJXA
GPHnKmHWsLCbceB1Iuz/skDYc1trn3JV3HnuIuQcdy7oupZDA7lYCH6fa7NEYn8AQ2K7/soHcXoV
fK4S/MheuN151l5gjsoENDrUEut9NSQM2g2aMDfkE68q3111r7+xFOnGxVzwQsFGP3KTHzoCnNIj
+1mw6Nlvn2Iq9uKJxBYtl3tUDCDgr54DkG/oXU7sQCFZhO3VCanSr88yWuaOxTaHww1KPGjQEmdi
OTWG2KFXFiKPV/7mC+rmsC6XSm3DnqdfCQaGrd+H1R5+1KDvVprRxjtZnf7IrkuEiuJoJm1E3vrv
SdbruLoGgI/WeB0ioKsNXkxUvGVdO2ghYZSCI2KIFBw3ZFU2QhvReTzEeNsASx2U0chu71rQ4BbZ
JWdtkFmuqS09TVgwY66f54QCl3ekRo4NkWEKjNmeSsrJBIzDrbhQluRJwQL+BVz0hUgKbwXeEpmh
UZi2BGv5axTS0OreIjgO+N5orDNCkE8imQYm43K3yuEUd4/2iRTZrm+CYqwKZFQpXch0DiSHuG8h
eXGyCMfs7ZB1QaEiYbbyX1CGsaly2rifFym7nCF0XyXqNM9SJdUWa/G31Ogao41WOChBIXOZnjvD
KI20nKY7b0QbGmSysF7kw5z/u/URtsn1OFLr5W5kxt0p5Z8poq+0zD2RUwnT/zVwManNeO2oKDy/
uXGFfWZKZZpxJ+A4YVZ4Hasvb06HEubCEjwVer9otY+1KSHFYIzN2oBbCE/jYUFUQJZyibk0XxCv
foIYWwWXRN/gh8BM8+GIdNIcJch+GJ5MxinhGaZ9gevlXl+Kqc8zZ0e5q0o3OR4mzd0kW/9UodVD
Bz2Br3a62osSEfGzdtz9HHN8SS1agZvLD3hqqUk2XL36OBTFg/jzbwidhamxKinF7ST7W3TUAD2a
tEiTNSHRFg/YvLjJSuXmE1P/12zLJDFsaCqs7gJ0j/ccB+l6Y4shpQ22KI+xaKfakEEexL2TN7cx
qKE51HF9hdAeu2fJ3cd1BPWvVGRUH+EQ6P6rtlGdkkXKuMy08R+x5lao8W7mj0lHkfC7I/BupCrJ
gi7bIV95D+9eb9weHn0fgLEhxlDs7k6Jm4jpT8ZyGfpF3O6r3BPbw2bQYVNR7xgXIqB5qYnuMmU4
f6qlHvL39ZqyfJ2xZh3eg+1AXL0jJr3KVSLnrnNs5DK/Zbitva3Fs3sGQWb4Gud9XfBAWpWNMnds
SsjZmZ/fRJ5qjwtI5DswKWE1JLbvnDQdqhU9c7MCcu/7Tf6S/25uhQ4WSBzFUmqDYFHFkdC3HkIi
Gt6/DkTK0SOT2A1VTNA1o5sUoRYp3Ja/9YbS7jL5JXquqnKfynpRYCvhzC59Y0cbCZgtDLiOb7O1
39BsJLv/+tdDtRwL6MqXvlgf9FfbbWKSaX0wiCEe9dt2vJSobxSn72rG+Wx5YDJsURyggFiTp3cK
v1dF3Rg1QqsO/IxnpHW+OYW0qI0o+mJTy3Rm1iwzGuFeHg8c0R5PUgb7Hdv+fEatPUTP76guWSs7
SP9dPxoSYGDjvCD3X9SDFhlgaf/zjRy5hOQyNng900RzlfRhqdTrxZFeUr76MYcw/l+Cx2udwAJz
24rHv7wWyaZ+8Cq05CNnbkl/SGsDMiiFqODGujsg3w/8DV8FcgV25tU74Y+8NP6aENRlT/3ULEbT
gg0qGtzp91osJNTCUKxBQ0bqF8mRKbQ822l2ucgrA4gBkPaaW2UAJELZYCj97SoD0ZoRd1n6+lyP
bQzqgBivk59XB3LJREWpVAu7JLl+ZzAVY5CQHMQoBeyEPgFr10YW59D+ry6ZnkAfjlFCcSWHn/3P
4WwVAAiU+1x4UHqFPnLxj2xaiP8V1kjD/6HWUmysPJB9zlTkhCmaQGp+fr7apguOJ0HieB9qIjeu
1rhdOXhGMF1aF5L7fFF4DnRLHmLTAYnQu27FzqmZI5PSrl3Wcgl7PCola3TuT/oBAMwFaGq/tV/V
WvB4cvAB93t6y2NBLvXn+DOpWoBCA1V369rpAHZ1UzMb60hFVzxelcqQrUzrCMRFCyUUygnFt/j3
6EL/0KKhfekuj7urb0qW6cEhwqIeQA4ldCp8xXhZuTC/ZvQtDVUF7fN/gIeZrD+J7A4rFAI7RVSs
pu1p8i+9dQ2+7gpXiWb9J0CXTKb4/NXmMg7k9DyClHdzJuF/OPs8LyoNk/MPyZiXpwTpOaR0SO+c
WzflR3ZW1KA9Ui6KsG4IAMStcBOo/idW8sD96MZqI9R0BKK4ftkziziR7d9cq67ybQt8vmfyzGW2
JX8wlf/9r76Tjr/wl1aU+0A68SUJ2Vw2BWx0geQ6EyGisgBmXa6XTY3kCS49p2I8RNtLGQjR1WXp
h0CVlx5NJcfxMUBA57vrmzESkujm/dxVnBra8MUKPdT/UlJVZ7O0meYpTbIiFP39wBf7DxkLIqSP
NzSF1OBAz1ECUFDcSLiH0cDrjMdNXUtnOSP8BQWp9+hBwQ1sRv2S8XHm4BSLXzJunC3kTxwQU5Vf
PJFey4xaJ9eY9iRZ1ELKLeFTztGLnIBx9VHahT6+4XH0/4+5a9LhKjIklLYdJxj72JfUigU4NHku
yZ7mQOdnS+MYKrRtixWobxA9rh1LzzmPs3XPeuOVF26tYXHBZCcxK/rjjse7+tNIKUsghnUV47Zv
o6y1RjVBiLW28aXfpU6aGjhyIXsBtto959AtnSMngt7/5mukEebXX18YN9yn8Oja7sUNUgb1Ol0F
Y2JwKnqYHF7sBEBvk6MxRcfJAEReCpj1T7nlyDgH/J+lf7ekbmv/NjOC/E8G5plxXxYR3/yYMexj
pXmiijmMU+73WR8cHSBhyzZThC3kp4C114pa9LIX5CZKIAR7vVv1LMmCnjKWMbYYRX5vuILzIhiC
g5ZD2u7tUgDtN42298KKMx6u0JOA2c2zYwbMhqWDZMzkVVH0+fFhlXZ/r6GmNA1/nhz+p+ggJ0un
P/ELID+OKFSc63r5GzViG9Qbt9iRPi1O7qxwj62rrxvBdr3YhWK2liTuReUrwbWxjXgIuauFVky4
RPYItMMAtb2OuxHROEnj1xVCOsAgMjiyk5jyy1BA1uc0/WQqh3kdGesKCRD2ep64wCuieTjzs6e3
LVU97TZc2yBAqDpwJlnusB6hO/qMNGEGy0qEMc8ILu6OH8NRPe3Y6i5DMj1GS3vvHCaD9uXqJZLd
pASbnvWl3l46wSW80ZQ34p7r1wS5g9Ew3m9N3ajan4VmwJJ5Z7DykPEN2tTGezz8ZC6zALdCuTDc
n/QZ4NVzAaYb4bUX0ze+OIY5fjqc6f4gU2UKjGsK8hmb8lNFmMc/rl1eew2UqRCK4os9zS50Uvjc
6GxgmBJNaQpFRFXhlxX/QSERx0igyp/TFq5o6rv/688pKcevuMeVg7JZebXphf5trPZeSA4xMvHR
UGz5SRElCmxaAoZmgoTCTRCkuLJmA5JVDF/Yv1PxPwYMQjm7MUOXwj7uIs6KDbw+n6dY5NHuadlT
QW2STv2Q944IrNWCwpmG23AHSAwrfzZJZcy1YuScnOLy7VxDARId2PT70q816jy88Bl/0GkSLPon
/m533jkbY20Ge6Y84U5SXtPmSecke6HCV6HJ77rYRc862B2n8P9qXf/waQiUzClG6mS32M98Pn/M
UTRT9iL/vvziHkN9MuZALLni7O4OIk0rU9Y1IBb4BvbUprTklk9/WqCCd4sgdcwSx/clf5S1sqKQ
HGJPtHiBccZ7SfRJNb1OLLhB5gAbMJVZYf2fJmpiLPPIWJWSANlmsoheII3H4qehWRwO9/VudBjw
Odq4mnPRsDrnAOcGvylHmYRjqcjAej7MBx24w4aAdls9/qLjw7+SIJDNHQ8+q0zxnmpg9B2IhBu3
njy97saqAuMkxyhEUO/Nz3gYpoLIYgL2Vi4XNm6LU7EETHbb4N7Ktf7Zz9jyUtYSMe8tr/2MFuYY
0jTFLxNZ+Yu+xD4Llmh9xhGE5eAXoVHAJtShVeQ5cXNK/oiKzdXax2HQ/8h7DBPenRzZ2piFbfqt
54KqZD/ZOohM/EvSbrx+mrY4GdxTvTJrGtEgS/7DOhYfJmuztsN56yqVN+k+OULpr+Ody97pzzOm
7hIgp10lPBrfI/u289z07LpLT9KHlDJWU4pNz3obnMmXJ4aCfKmLYJ44/Az4qhaBdQ8ZWfUiS+FR
2ni2vPknWMlH7yZKuF2EkWyHyzutoBTYce0lHi/CyfysQYXX8j1D9dAxpp8YUC4jR1uxUGPWe1yN
kNC2I75FzHaz2B6HLzcR2BHtUn+cUvxP3Js87403nJBB5tJY5P+gkjHXkCkncN+PiAFEu2F/PJYI
dK4ndhWL5iifLr3ZjTcl+yAPdHXFRqDX4wNGAoRbutQ8RyY3hgQTvEiVJvYX2O9+IvF/fP2Lwzqp
q4f2ymOJOQflcEZWuVfwi1SGsmtAHrmvKtHqyM0npacx+e9Ubb1BkuWrMJuEn0FUF0PPJRZy7uxi
AAWa5ASw98gGCIQgW5o+rueBg8Uv48OP9h/sVzAdfX8yqtwVN8XhyWX2+4naNQ+tXmSIzghajUm+
/RC039gNMPydn8aoHRxpKemoELjjtL7tKZFyvfrZk/ob8LdD0GEixp8041siEEOJXb/x7ibnziiu
LVjTPM2QkMM6+ZIajXTPALB4KizImJqhE49NpVyOpdbOna13DWkAkY4PXykMQh/Bu6k4dkUBEYqv
sGWRuWL+CWdA4Pw3TAQQQ0/Oca85hpghdDRgnJs6TwitMFEODXzor3VCZ9KNCWwAZM+97hdOUScS
rBEuISMHgdc8Xk8PspKTx81QMVz4ybNGkY4/Z8SDCeYpTsjxHr+lBziTsUzopN/rSLpe5nUn4jfN
8J9SPW3vCoOqLeElodJI4Zl31OwoyjkS81tCjioKEGn/ooj24Hb4wIDVlcP6iw9HzBS/EexI/DhL
KTOGyLXMF1Q4MkdVXjRH/jm7002lBnC+FDDiTMTBwbiyY5uZVLVYyf04gWz7xMsTj+c8hija6Akq
cvNgDuXmRf4yzA02qprD+GOTxk7RcK/QaMKIP7lSzg6badlj/wBBVnWYhsfFk4fpLvj3+tHqgqFp
vWBwyqt3Ii/quOThSHXqil8Su+gx3Rv14z8BGq61HVscrwBAO8gbZYUR5jYS4I2rJLwpcn3xDH7k
5rbgWRglUFOX33olXgfLBLDjua2s4Dv6LprAoyi7acBMl1MQQ/uAXqB89OuSJsF+o6QurlPnjCZT
V2Riy/lXwOVb4R31DQoS98vggSc6v77HJ/WptUcw5RdlIn7uw545sKWtgFnHDne3vO0rgoMKeDap
uUqsFsEIkv1/WxLQjHU1G6d5e/M00YcWlwUfvOLHs2kNkm0urwOQh1w2xlGzupTxvHHVcc8v8MTj
ozo7G6vyhqiwfFL0OIARsVMR6zGvs9TAG9YHTxtbfSJKViwtGc+4DpfootDiJr6D2u/nn5sX8QRr
S7gPCHsghOXspmiekMOpZxbNM5SQVYVyP+ytHFm1YGhlIui/xdi0Xj6SELxEjkh9gm+lQkagHhSk
6sh8KoRcixg/5aQiOv1CLmPg5I/jduze3hVbtanaVglCbEJV1kKWsz96lWoB4i5ozWAT/FqpIAEr
vTSSjSSwInZMzCfd23uApMQ7n1J+z3X3AQRfIlbTT5W1adIX6bTGLSdbuBX6Gsv6Or2G2UneHFl6
UPp8cW2FxSYqaP4Ts1nptg57wUZb2gVNO7xJL52NRZA8Fn5/LtBt693kbuq+hZ3KSroveQ/7jg8V
L3FmclAGhCuEeShxgSHS6yhGu7KQZKfnYiUsyijr/vMAb8BtiDXYUwjVEr0/pyzvyUaYWFKp4M0K
emVRa6X9rnAVW41K+MOg02ZdgDBMUtWE2muxNq7WQpA6Zm6j/E5wDodZljCy9cE1wJ/NgvSoBPEl
S25QVvYQTJbplBv7ogz11gkOhwTCaBzo/FKYsGbFKIsVuUMIS5If4KfJbTcKYsZaAOE+NZTpJZyS
QXvIi358cLOgCgrXPpQkarC4JG0wtKr9zyEivh1A1Gc7jVFOsR6TcIXzh5BDSTImbLALED/FqZqI
nXvZCG06jXRFKGtUVC0Ldvk03TYGZa2T4xMDpuiEn2fWaKLZauonZMQ9c0niRiEJmpWhWQX7Z2X2
89EXkYTw/IA96l087XValbW8vD2af2NmdQVPMdAdEiPe6Qj2jq0bsiARFJqd1PjYBYItdPgC9Ala
oH2yG/XdcSRti8y7qY5gURdevgQXEddXryLGr3Oo/yfeU31zSbfH1RFbw2gRQaH+7tppFw5qNVWT
wUkbB+bWe05B8TXxTYWbfzXghuwN/Ep8tev0JzlN2u8W5OQhxBnXIaPEU4pUFDXXb/ZcaGkSba+j
y6wtiokJmWS/i+M5LtTB686BfFFM3loImqKD1a42cn0jBdJIrXwTsihHOQPNIP5RpmAY61PIGkYp
1cAxpT0xWZhcQvRT3qBiQNUvr8i6lk4jPkiaShsWROLMrL2O4YhfeP1aYN+kynFdfy+9POPN4dhn
ur1Da1PqcvOJUOVKISKnZ3GiR/lOYQhqZBu3qazzUibVMNKVadifZxvD22loSP4FWKd4vommI1zl
RZ0icZs8vZD7ET7tTdSiXnKxaoE3/h3ALSPQazrJw9lCFRPHPN126tjnJvIB9kXzrn60UQlhqXZn
5Ll9KjMnF4/cX3EQZwQLPTFFIoi4++qYfpiql0isQLLivaKIi4qApASjEQ2+8NuH9Wp4mPuKnbHv
LJ82YCqL/drtW2Dp5oAEC099IVyCeew4Y5dC39V0RNeNZoGmM8Fc7j4Bt6A5bvHh5UGptmRYr30G
eVTKqeycFtmgRqIvdAkJdoqJaEsKh/U4eJN5rrcIkJ07h0w8aPKU225CEN7PCcpUUrCLeQY/+uxt
Xx5WGJObeyxho9lwO8syVfr2cLtGRnSRlK1UQiUpWC1sQaJRdwMgdrAO1EC5RLNa4Diulzr4a6fW
G0lqP+t2q9k+BGROf3eigYCE96zLd0NVSpCP+/FbuQNS8rDtlm6mo1rW9QwXRUsFESzVF5ZEjg8P
ZO13FdS0NLukP0zlKCGj5l6Ne3FyIDNx8k+0e79MNH/3/h3JuPkXdgjBsCw4TU5KDKDVpds6atHg
iENZIjJhEEdIY0oqo7HShGTjrXe/bghHi6V53QnsrLNcAAojFEmrswvjsaHmYI/oxQP9dgrGzEEa
gXx/MpFyUUoa/T7YhFzm5RA2WPVjSVqKGJJQk31ypS8UJWogPifsKk6u4FPbcMgj2Ot5amj+yvrS
BaoIaVzftfy6u+ct673dIvhlkZWQQc9ae2MubnxVZR+zF/aDSoqIhVjjwFxdCC0M/iWWanhYNldu
ZmPcsagapzJA4Os2+ehwpqNJL6cH2R7NgRLBfxBkf+chUYocz7TWYatI2Lkmt6UjOdl/jSE5U0N8
Tp94udit3kcD+cakLPgiQH0mjCrK+p0XqQ1mMvUkNyzA1H9IMiCZF/6vvGhKxrvGFutnD85r8jvu
qV6VWF+etqiGUQ1MiKlsXmc5h2NTGWlPF/vRgxGSVoZk7lmySdfjA7RznqFYTHA8Wl3CYafjFEuc
mDjNqh8J3fdGDLLa/ozXDXWvJLLuMjYvmWhzO6FYgzR+OYPADWKjqNZGl6oiLHDf+NwZDBpDLpJN
xxq0gWwoNahIyUN06zFOxody0hjkWttQPd3NL0VHex82WW58QlqZJbqlmjJrYBvWWS9ER4f3jGge
1Zm/w+y68Cpw7o1yaTUeADOzqXmWLefKtARaqOcXhMzxmGNgvv24RBS0hlibL95lfT9O2LiGL1h1
RBq0Qk+PMqibR/6ynproDUdP2tKPb4Of9F0x2F1/j2XyML3w8sh0eH3xmLJSkyj/DlycChlOEGzQ
41FR+6ZDC6hJYk8Hm36qpgS5gVogVJycCkhRRiShE0K0cNIiGYww2UW9bQFFIyZAatALieX5jkDq
BinrTvAjCGBc8HuQnYYnpgYwWFg9I8cxZj3ohUX823/1EqFv2x6JJ/HBrnwnKpFhfgC6lqBSrFzy
EAyumabxIGR0BGqA0tBfBhlU+/HO16qbtlKTa8/bPZFSFhWYHm6oInZVcT8pSYwRVnvaTQHoNIH4
wQ4oDkCVJgaaYopJJlHXdKNC9L0xgxvDBEpmyFza/wtXzcIOkBVyyFT5F4e/7bRbIoe+cluy/qs0
1vsYj1bMtMUn41SF5EYMPsQQjGeZGpo5GRcB9I9IXNEhf7yL46a8F3IYcQxIkFJqPK2VUaICUOOv
AbBaeq5tQKr5YrRlWUlF/kquG5vEHtQyGadhPl3ldbx4KAigkuEL5LnLFAXLuh5LsM8Ac6Jym9JW
8QPjpTuvd3Iv+w3impWq9c/+t0fYR7/xCvEoBW7gLFq4FuoHA0TpnwCsgz1zplVy+HhSOd1+m82E
DxDM6qMYeGW7pj17ngNmfshRZB8Dm0z+N1BTRJhdNYmFfLvEQFOkEHgJ4pkPgDs9UA6ZgO9S7I/l
z5w4K7G7h4fDGTOELVtVDkVFJ78eMpLc37ziHm5mIBhd1yayEH5wn/JGLIpwl/LuwDDAM3Oykb7v
g5yVqrbpjzbPOp/OTYWMe7T+Gkko5C10deI4ZZbCWqXlMpsYNwB3Wif2bUFrYCw0St9JuwM4a4M6
DYcHQLGUgKgMct0T0pfY3QoAdhnHGyxkmozpTUf9GvOjDY5P3Un6BRAF4DwxB2tog6APxrEEU+5o
JJ4Rp+ukvok3wHHFTVGlxo/3GZmwJd9GjO5AaciYbFb4EzA1ABvtXp2ir8rq2rb5XwU/VJeCs1+6
z2tVdIOpr49QNdorDulB/kumD4QmdElDlWVNcgNGKm5p1MKpBCKRCeSPvXK4jwbroSbGx7BpZ3KK
yWklcPH7uHw8dUJC7uIbAmeVg4OVFaWhTDBDVhr+mCiN7ToQjHqNqsvp0jE7oLEp7SFCIuhcVjqP
E48i0rOvXaWDMsvfWhQslKerOxjDMA5UUppt1Pz3hcJr0QVuUiIE/bGg1ozwxZPxBLxqfOqLIq8g
ndsI6qwRB5xbPhtdMIvQi33wWZtRvEytbQZ3u1/1sv8CNxz4y2zoFH+eFDGAdQpTNoo+Tc3ZKyTw
lpedEzVjjxsn9jFnRdVyCpWSPD0LwAVdDn+bvFqkaEquf18YMMOVwAF4EeFDczW/xBBIi8OrCK9Z
eoSvFGoBQlIPfFgZm3eTts4gY3qF+r7BASjGsVpWltcyR/wLPwgZRvgGZXbv6vbOWzOszLAPLv+y
ZqznIABOl1Ptb0dkUGeB0hzUhiFxrB5SgiClAVPgsxT9SH50li0fLzKxVS56SSKzl38BczyD3rKL
Gmat2zISST8bPS9NO+rlZR6YqZcZodljhaNUY788xIP04wCNAflFNz15FTinCMmpMLVaheRB4z7q
8i6RipYIRcV8h80nMO2n7itLQG32gEvNJNVZBUTsLfCB+N3zn/Tj1vIeICQIjpKeOzFYuZYvxIgr
/vvoO7qIYeWZhFbLWEYnluEUPB8yzA3XF9jmRAxKtQ4DJgEPNGeMNfamB+jh1e4Jpbc0uaw3EQTB
ewvIA7WhhdI6aGcZZ8S19//yiN5c65ITl27s6Bl5Wd1JjP2l81LN57E8ImzzaRFSRN7T+veFkJoi
OVYA7jicH2JzKbsqBHmt6NjfTVizj2H9BD7F1j59BluKZezm3l/PlcexYCyezgUk02EVjDFpQ7pf
Hb2W44rSKC3RsVtW1ppB61t6waP4f9GSPkkyVMU3jcJUtM9DRa9Ue7A1wCAPcl4x271kwq7n4jzf
gkk1qPAZMz+6S/j7nbsxormb68Q+7X1ZcP9cCkf+MpTT3jVlTIVbOE7qNoWHsnFOahfnVqX77/kW
caO+BDeh2It2cbrVQNBdO6uKZ5GTg1FyFBEt5cNC18WjbBy5yTD2X735NXUnmYLfTyzfSB+lya0u
7V4TkCe+JkoS6sgoKS5mTtcX0LhusPsXrQhqo1zoXYwB3j1gRfT3dcpyY1hOMK9uYkYsb6sJIBNw
TDY2EUIBu2sb7WziRqrPfeAW5ZtB0cr/T/cdtqQNP9Lx3OIr7xbfPOKvmsiSheODxyA6LgZ0pL0b
0fRCt6ycLQciJ2BBzCLEpJhBcOhgzo9ooyA8vURGIIbvOxvjLjexG3+ukm0OUgb7avKirXV7ZgrK
2H9G3vs3tQHkSYtC1nhlIakepcmHBT2lF+XHGf2EVEHhGxlAJyNUU8oV0kQt/fuoZ9BHDM9Msef7
3w0XIu8nluopo+SpMw8SIhP6GnY4ZzXYFl/DXPQZe+HgyGcf3Db+TxW0kUnmoQTf5w7Tku5bVDJQ
29wORCsG2hI43AC2RVPhxam6zZ93zVbZV7LU3S9mj7lnvazdUaLdL9cAPa+7PBQQwTEkaCa8TKH6
UoWNtCViKVJsmyJtzCW3/SF4mnkeNWeBhjOjF2XjTtX/2KxDteeag02pqsHjCsNEYfNC6A/ckjyx
lA97rdppBV5ZRRp3WKz+oW5YxiwAOFWPP5g47t0M4Eo5lHxpUdYux91XElOOyzgICA4gn5PsC0s3
/IMc38kTrnMAhdafLVh7DSNyove2/rQj0MXhQprjdPCAXOeFv3vsCJ/lx7jnEuMoZozq6yRanoIt
D4IZIr8mETPtGWbIe7CLcckhUStwWTugEfkP6THP1OYKQduiiIMDJq6BiBLC5dpeQLzgSNIR7mjY
W4Uo5v7DpFNoYLSZMICHnZmQQOxiYETNxlUrtjzbxiD3LwoXN4PE1oMFVl4rFn2eF88R54rXVKkS
evFVX8qdE/xUMh5gA8bPQWg0JPhVneMfYKgPM92LGFI0RD1qH5QOFek5DURph7mSiF/I6B/jPsOm
vWE/0F6/kD8tt1iYLzoUoQcA+Ge58zbNovqJCcchsPrDTVAsXAXgswlsSS1m0JepuPBgQg1WZ8X5
gPPV2Jr9hPUybjSAjXfqdog65magci8QfXeFPuY/LGW9F8d77aL8REXnGKBSQbn4/QcPDgrWae1F
eMma5XRxMFTJ1q8mUtT+dKW73bWcFoDeu5pJPURSI2HkJdD36TRUNJUfs8dhptMrn8TtLFroVLWj
VxibzvGegCjqIw/4CVNdnNgJ7a64u3f/8P630kc6+9HkJD/tQKuTpiiFxPwalQHWJcoeUJlto5iz
IUvctoHfU+ePr02bznpgQBvMajxdw33kTFgYZi1jbE8mbK95F0Ntm5r8vBk7Wpa0Ru0dLeW9ggrO
uhJIn1TEF4y5rYeYjbFC8M3HeRroR7dRTQmuS2DmZTo6c0oVXUgegnXDUv29CEDJmjNDbkjwbRGi
h2Aj+4bb6J3b4YHcglQ/SH3QjwTbutzYJQw7TsSf3A888moUlqXcMqpPsym9hQm2zR2LmXeni2GU
vrx4TCM6YnRHo7+/lklPseYiaaUEjmr8D/jGQQ7zBxz8O55mJDs6j1h+IlJh9MtucyNw/WRToRLB
P5ZsBkfWL0eT3rGsjF1sMbzjWX/MNXojLjUTDEKNTAbdAxMmFxsl5u0QJ0cBJ+yVf1lGZvdgkhzC
3hf4Hk3VbNyKFqjCKacZFJ1I9/EBHRR8TEoGLR74epre0BNlqKw2XzARK2rluXMIX4I3hW27gK5Z
F8efiCL7LQZUAk32i6p9VuV3Zs7gj23e1T5XyTNfeAAgvyELihWjczREmsMOaCbk611zDK3Ke0ao
I3XEbRnIPKFZphHX0fMZHjapDTDSZrCFSWGn3jbRc4x4HFKG9knhXCsOMpGkihXZYis7YwJIJS9z
xPOrlv+yN4X4rWcJnlAhiIWAsvhJ1KzocHM3kDlFVYXLTCJeyOeB4C8r86ntyKvcwiZ+Xo++lyWv
2pfz6Y51p6w0K5f0xi1daOQ5GDVzNBcr6/Gi0P4tuaef1r62WAuNQLqmWTpt42lPvIPBbPL9l95Q
+Rkbgn0PIHtKo0QIrreqmeAuUP3DHG1ifeKeZp5gsoO/sBShO/9gLnPr9zLjxu9hxcXevs3YzKDo
ZYOx6xoEWrl/j4z1HeMatio3bG8rpki9IN5vUolzvkc/e+2d/vmw+ff/iTRgYRoyRm7oD2kENUIa
KnOKFXSQ+4d6R2wfHVL7W3BuVxD4n7hmFJkLkqq+Fht2csdnQiHr5B3oIInol4cGd286CyPlfgjK
Nt0OKuzp7XwXo2f1xL5KsXELwvNnXZrRAj5pbatmV9p3qcf8RMYo0psUzQ20NboLvl1nyYvH9WGl
cxbszOCMcawfi7R8mG9ivCNfGcEEXUiqCMvR74aS1wMfLc2zpT04d64Rf8JFqzkEBJPRXvL3Wauf
gfXFA4hESg0eYw6/hhE4zQ1RWl6sqJwJsvlb0dLIL36S4Kq5ADUGKp6/YL8niMts9LoW+6TOgADQ
iaKHFBgFVGiGXxIowjElqUbv8nC0KutagGGG+y1vmf/lZCfAzDMyxuGqgSX974/MUuCByoGV5cOg
UCP4T4+KwIO25qAHiOxCdxlkl9+wiIVo7nQvBrGH4fztqxPxzl8Q6asuZVZTbj3o9Uc/qRiwlhXQ
dxQ4BOrT8NSs7Wr9h7v86Q15hpDgxPpRGQ8X8/p8rp2HBFqTy3pSb13nL4WYflhXyNn2Q9dL/Vj3
Q8qEFPzKhRCK04St7GY9/emQqhfMdyDfYp0F88+zvZ5Hqvaw4KsjiUcWP6qZjDbFKKBpvc2xl9HU
k9H9Ko2KPzRe9tOGSIcWJov0vU3jS9ZZ4PXL8CV3bDk9FuzdEf2onQxf0ictsMGMKTE/BUUHv78O
Zo2ycUU6KZILP5xclU6i5FaJpmDY6Y5l3oZJGSftzM+v8Nn54PLBFx9HjV96ZVKWC/wZVsevIx7n
tNDXu1Xz1hk3hOXuAgbEeRIBnCdk9JsqAXNFy3wfxU5dOE5HYiVIL8zfQtHYCq1xqa8J0I3QEvvj
VOBcxOq/VovySfMCQZJD/3NzsIr5WZm/5gKP+fw0eJQVwMFp9IG5znzoC0wlNB18Yk/I5gZEm1DL
6jAFo1Vm0Qch/HaNCJmhOUsbc9tzzUugoKwPJPBqvBhPZnEtd2F4R66dxnKuQvetR3rFiDFxUgzp
P/uQA1UUdpd7n0+TcWKsHrSeGkZG50Ff+kNfoB02x/C9bdVyY7SIKO1Yc6UOM+OMwdnCarOqQFdf
j/wjFxT+h07LNCq9/yX9/pPZirp8+x3J+oYeJE3Yy/9j19RndTi4SvVU5nCfcVvKTPpTI63NRbGb
ETPYH4t8nzyjqgyeYLp6cTZhEJnuBESBfZbHGk/KeCjHWHK/xV80ylD/cK/bOMJKPA9/kMTzLW1f
ORlLy4ViSZT75iNaFG852Ia+sxIjEsH/3z2363OUwfbg7YpDQm3NUNPtSmsGDDFvJRe2wO7+RUIr
OLnLkTcM1pqffpEaow5BtovwdUyAUSBayO/kj6otWCKINmzKgdUlSXFJUieCNqlbLJj0kUZzcree
i9YSqlHSDKqlvqUJWgBfm7CCYxWu6lxUoQm7kXJxyLQsJUMw7dxXrk/mKQc4Q4oWQJXfdvKLAbku
58pno3myre6wScdj9Na8kjiRr1toWU596C0KklCSsCT7ZmS90tcRA64auPCfrCOtfnOe28MelSmo
es4ScFK7EFqDh4Y+JxvcwkHSyXmm4gIDfwxkmZ/6vWsjppjoQm0sUudBhHnZiAOEQJ4k9ojMhqKM
D2/hil9Gh/sVYVtb14HO4VJQh4MSiXSbaT2doVYrTN9FrUwCj5be2B783SvC3egCXq5qZyPkbmfc
eeTy2VW3snFWd2Xxrw2rFSO5xOZ2t3KN9mTPDNh83inI+TVddf4TEzpdvLQFrEux5+xp2jxpHjjM
JysMFv+R4SsX0sqX1R1PjBXSREZt78bGnJ+BIPA+6xYhyofSN5QW7JGiPQpwbcgitNwp8anUvCnk
+QhJoviJUtcHvVXpyCBLhhb77wrMnhx+yeL4pFQJNUSYkO3cSHkReIm9ql1Kh+zDr/F6uDLMT2sf
ff9HOOHLlrQ+FFcXk5Pk/jzjo1VwgrOJp8bRJBEJO/AuUoL1pR20rwKQfTWq+JJHgOfOV6FhbW1/
eLIkJaVAzOqt+pZMrqEYEngWgL3Z4sUBYz2A86DoFOy6vqrRzbUNW8wCsrEAbxRgBh5pBKHQmej1
cYk/QlPzUe2m5P6oENyBbkfx+5jCZ0cEBAjB9VmBugCCJHN0bMlapyKvyUcURAMQGgqelD0hx3hy
+mz0IYJi0OTYOfN7nciUZNzJg9ifyqn2vOBQzItTYVoZnNxMRK8/JrQFcK0etydM/6f8vrLltJ1U
1KAOqMcfx0HVRHYzLzKJ0rbI5CNeLxsgyJjJzoz5dT3G5pL6ADwAm6p+DxJLewIE+ZpCu/JHAKdy
f4V0a6wuFo4qPdWtdaKxu/2WxX6PghNvZVlXSsUfzcbYoQ4zleEZzuefcR8M3jFeKcgePsl3p59B
NatOMRbCV1p3WSKhWkblDu6KOwupe3O4JYQzb2TgxOCo18gxJJAxSxryF+Aqu1fQPmzkfnsRg+1R
nkaEjmIfPgiOS78S7wkx50O/xCwQX5jQPnLBzFyDrqHug02fw38tlh68RqW70Bf20EpZoGrb3hD9
49sGGipBQN+sKYr1vdqgAgYdHkjYAc7mIgP0wQv0GSeiZyk3NZ+oqNCP6BD6mjKOwq/6pp/wwrDv
iTtx7NlLIXlnqulJflawd/+Ry1j3tW9dJBcRQ5n6+4atCMb86Il/0Zq9QocYqRCpVZzmwiq0CrIu
3beg+F22WJ4MhkAsA5K1Bv3cwKwC6Gu2XpXuBStKK4Zf5HZ70n5Mp6qyW49HcQ6bK56p3iK8jjQQ
NOXklcEB6zzPcFQbnGXC7vuQzFZdn09/Q8bIXs57NQVK8icChnrhUAD+5rhCgOkbh5Pj7pEwlsS7
PrlBj3ispV+EzmyceWID57AqvnYh33q7lk8j5aEtjCIJMQlNOKQULODwD8tizizknbyYqCOR7Jfw
Toj7JKdiZpjRUk491MaX5VV9Mw2nP15hEp4zlf5bg5VGNecRRkHORi/5BL60rW/EQ/87WEKuFlnj
rcm+UPrOCYW18n3Tr6WcvpeW8IhOtfeKfZ7wL3ScnVHWG24TaPsOT7Thx0TlIMp1WDxsthcLDz8M
/b7f82/Gi/pi6nnzfXWrw3iU4cUiX2GVxNnKFiUBg74QWhruSzPzBJHRDtpIYba+1ATuL763cpVB
WAFcfS5M3w5TYxFF0om11PnaEXfNyj58Adx/OYKEtNcftrrmARaW8ZMg1LDi4DVgtyiql6S0zAYG
f3mYyUxHGJ+gVxIf13nLD36yvEA9CBWrEyMKzbq/mJt9Nbj3Z4vLbPUGB/PW9iCNqveJ/kaws3PW
xAsLdzSt44Ua4KzR984y7GzQ8QWC6gXlg8/svLPgP6HqpIcl5d5rRKtaRCyNPygy2qHKzSNsC96A
W2pvZ3Ev0x16B5Pqelu23wPWr8fZqd1LUn0uCwwaUH8868Tp3m7lrlGeJQsO6Oy2pRUNItCkZQ02
re7PL3L98FqbF7LQ9YIfnQ77bPwhRNlD4qMNaYH9Rjm2wA94fGQvwErJU0KqNy45tuP56uitKDs7
HA5GDyPkTbRuqmS0mQYj1Q7R08/hXrUUQ7Z7i5LK8yBGniVFB/QBJ5FNU/eAGjUJYdup7W/kMrai
udPRE9EO9UIUVhLcWvF2j2SvS5uI8twtRsDhKfRsOxK0gJPAm3TFEJF6mmi0lsHr9tr0/BN6YBFf
C+FR7+ZFGyHMr/8OkCH1eULrnxexNimmkC9Y9Sc8HRkcYWXrbUFtR/cZ4jZB8MExm+HoYCS4Jqz/
QSeeVzp5pOb8C41lRmmOjTnhulIE9Ku8GQ8lyaQ6KzFiBPZ4WE91MVkxCODFjUXuKI7nZR19TA4Z
1RiMvbAevz0fo7OJsYZ+sIdgZ6WXFaBAcxWP+7sSjjgCeZxchwHlYJAWy18RUTK+PIh5SRg7k6TX
EfMMAxG+JTYFmcgsHIFEqDVyQJwALbSLrdKJtK3i7h6y6qEXkEFPfohrKb4qx1v0w2R8n+DR5I4+
FgHVj79I7oHgbBDDYOkS5YUGBDEMlVFLz1FZwOiwRysS+MK1yOTiZufK2UrH7D1dWICyDsKW+4M1
S4BUovHYRJ4wDr7nlxaoFZot9BMkHfpjpfkmRma/x2dCYiI7L1R6lyt2Tzqy1UddpQgA4CIEZRVR
S6p4Vw4EDfKHORfBCg+pnGhuMFtYZZniHOMNVwRVbnGA/cTk8vf0YPWXxf1EwovhG2b4KWos0QZE
hxHRjkQCrtp1vLMWCTozu3ZbA+O/OzidMYLlqLje15MtqT77M/lkUPqmvUVdTJq0422bZMWr2e85
ujGW/FfFTTLsr2PaD8nfKqwikoOJkIhgKWyzWEFdTlPQfSOFgZ8+q/XXbOQ6P7gctp7KoPgSCePK
HP81NKVkBIiGH3YJCbRjh+LGMY2PnGXtIolCGk79NhxBHHNQNh03o1EPqP5EXJdHkVwj8BuyCdgs
EzN8BJ36AR8hnsAaakWEoWOXn2zKi78L5Z94OWNaYZ0rqFs37aHWZs3BP8TvEBGoh0IrUKGM9pAW
K1GUtVW0JQDY9GaO/L4rhMOOryAICKm/Dh+Zh2R3FvegmPIjrRfDyb9jqxW0rk4wHgaocIsf8aTt
1cUK460Y/qb7dGcKBwSRyQgMYQACYgMVJwtfeLiGAJSsl/PzMTj2Y6OLdjJjrg597LzIv7wwMZPI
c+a1/9rmLtOIJ1QkEjPVgjEfaaOMpoqqFKbnl5u/Z7aF0XIA9qQi1u/yNnfRWhe0GMJtWxwL+Wz3
bGDs/DQ7Gm2LR/44copRuJFhWfx40Z9lwU3noZx20BqMDahIVTfcnA3UAp5fb1KMe8t8NszwdN93
J1Ubpl6kwNCsu6tkKGWq2depPd3koFskDxAEr1LsS+wcURdUcHo3ocfNhOr3ljD19BxANnKz6kYG
G/pRIEShnQ7bf7mRjhlRQEvanhITE6aBeGCYdKKJ/sqfI2KsdzAN6esiDG2D1LMDYVqJB/Tw9dcu
lVM5wYl5P3nFH5oipDR79AY8uFbHT4qs2Wj0Jko3IYlmF7yeXOGw5wyPEH6snePKFfyGTtg3ZkAo
ykZWFPG/N1DkaVsVBa8p68smTSODrCkEGU0pVc95yYSoxA7MUGGpZVeY9MSf9SLnueVl7pzTLlt3
G9WJkr/1vEVImsf/h/mBYTMcAT/81QkidqF65PyHgHrHRUDGFWAoNc2g36rXiFmaHe8TGEGOn+Qm
vNV9ZbTszwg0RtiCVnmrkzkbhpNVmbYKteLhAGxwBmYEM66bp5j3SZn940a0gLCk82D48MpqaGrp
7CaEyYBnTIKGFhmDtvm5pvUgnUJY2yHXy96RrnSIMhV8F56yviPpASXNMxFfRwD/qcUfFu03gkre
Z7AM+8OfSh6V92/QJbalLHrUrFg7665rk6tZpS5MsJvFOBOv55qprIvJGoj2YUS4RzkU0sdYzt4f
wZvmyIQ5W4a7/TJOiKC/6XYpNBd39pg3YFiH0oesAonKntFJhcfQiafA9D1voo0DbOuOicGSK5XD
rVFGNC/i3yI8zUiVzSMlESWjmgitvfMM5E7dsow8wvhLWooQkigf4NzzrC2w5FKzML7cTkZWHmh9
AaF3UqrkHLp0srG1aXfmTlQO1Ad/v6i3H0FqwUuXcdHpy1LDR6WpvCqGfHmLKycUGOD25dNwSzdL
2uMDu+mbNZjSFyGohJ6gQ7vYVM8+IiwNPNPcjrnQQw92B2VO2eAxqfmMzYueAuycyHeIn9gXzlkZ
KNbkeNZWhCbuxLj0zq0+/yDTYEDnhoq7DEpS2FGn+W0XOlpNJppxndzu+iuvme/yoX4ZheCT6tHk
J8R7IJ3QdVH6HoZD52Y8xuWsZMQIv7ZLb4XQbS+5UYBa1WF8S5MnB2/nTySBb1BOaFunHQf+YLjt
uvkEp1N5HDjGiTuuObe6fA/J/2FFC0ADY/D8MSUCYi8qWm9923BSuzHMr/jtSTordCQgZmTaDXnZ
0tW2oHCBPv+3mGstXsn3y8Zd88O5oa8XSVIfZBSaxPEKuIeYmgqZ8L7v+CUppWF/NvybVv0T4zw3
aRMhb6pcpelmvM04dysU6D3KIdJgwW03bnPOWeb5DwKlq3ATunNdvs6c5biLgepiIdFZEWQHf3v1
b59/p92tsDFLs9GdApv+ij7x/vKuPoprxL/iCCK4ZRju9ONGFGsG9v509QciYIPSVIY6EcHiod28
Wufouyzsi+9cHIpVO5j+FfBFTe3mNCGK9Me/5m5RNK853KCj2WBYdHMNXx66AAwzkj8S1hf0xm1H
wCqmCUcxTjUHrPosHdtTpCndKYUyYNjNcJuv5XMdXThQG5VpuK5NWPsxG6XERAiVHPxrNjd0jSZw
4SGmdrcnM/fCdvKtcFJfNIL5yBEuPKHq9yrGX2hhjU+7vjEepBwFAUGiAWPn+drD/krS6SNIzhv2
AhKtYnQ2WYKgW+g+pjMmN91sTBVZr+cexk/y+8JgVKep+VDqAbZ8uNNbfP9EQ7+ve5p8XleuaGZX
Btv237VTz13rR4mFJ2xUvTxqRjEbOM1Hita1Pwhn5io+jxknKfSM9S9lJ+rywvXgEhV5uMeRXRaY
G7JGiqntHxeEhkGot+UK5l207JmmzUaH+y/B1HTnDWLMe6ebemf+hvDk3oTUiHtKVrE2HwM5u2+4
1STDEWFmqHMGuv4eaMhqrXkGfIC+PF5rTv8BVLTUzBeiuD3l/oEysMn41Oe9Dgj05UXiAcikYa3L
EQM/Ijz0iyYGyAG8tDreX43W0HCqdN95552rjVxJv9Mzy560RQktzQFqrH8HYwry5E+UeTgzQLGW
+hTymMgw06mhQfblyuomxCT2/NBfk2LGMOhHjxLrF4vNd7+30d5ZWANDFliKVRetOFwFHufC00rP
icUmHdHN1Y9ICIC9c8TKyy5dvGh/jggUJy3yc8+ES7Ryq83D3sWsZOmvR4HOwjnO00fpaKR82lYp
oD63BRTa2gAz6BulGS9X+nC4J/eAn2efJkVetYT/bQ48KH896jBzBWW8uM3poz6sybgW4POjRy4l
gcN6QR5LzhRCdJVQYye3kjs5LFceEdE0JvRoc+HiQkyHW2xy8Xp6fTl5SNoAfPdSrJ0he1s1QfKv
jR3OdmNN6mZOE7tIpzFC/SSwBlI+9mvFvQW0jyQrxSyHZdniz+PjWuoayYL0y3emi51KU8gd4Z3w
ViKt19yTxNgcFeeEQuIx8pfAunHlXpIOjyUlVFs0w8890Z1fJqJ/R3HFrXXn7ZlAbPFLAUn1Krbn
41iRSyKA2OzJTW3tvWl/d1lwVOCDZ87+jOo+sEVy6kt4Z5cl68ci37jLo9MI1FyBVFFLbYxCu0wT
c1Y+ZYJS1blecKKpI0dzTYPMZGBjst5MUPlHTcoZPXp4ZUYViCJghDqux6iMDGIsXLLIi4TIOYKp
hXXoxnDJqwQ+ojTGnS/w2Blnx/CcRsYPfShCDDloRKc2SViwEFfLv02jbjYWcOS99TpyhynNLhbq
rmfxaxVwNXpJQaUQBSFm99GDBgDAkFecb5bbeSMC+7beMWQxjA7BvUpUv3TndBSKrtFAYb/eAIBu
0kA7pDYWGjMZFKFqDbjqSdCzs3b7Wd9Ijv65eRpdGVVfJBxjXGOu5D7RtGusv7VQsUgiAeVVOWjk
ro4amQEmmedCanXDDDo7WwnkjyUg4YkB8IJzJuyZUZMdVv/uoLYkAlk4X823E6xbYftR9CRspByU
2Fk7Mi9heyEPFhxdRV+DDB2/QK7IblywkfNDyXWz+xuPIMronKSmMIVMhUKUc6w75dfXqGOeS/z5
ccFRdELxlPlRW3LNRNNuHFLkN1n5GesjKryK3yfKa/JvxInarTFLbFn9KqoiwBvyk32z0uAV6EGz
L1D7hWSk+LJ9hV3svXvcCIDWSCosHV5RX0iOIYREwhOBKpYi5yqR8PEbyv4qO1ny2HFIaB6HVIH6
2uuiXtlJ+CHPpxwPTU07E/sv5g2zI3pDh98aKGtSZrjdNAU5DZJQ3ZSl2lZ2k2vwT9BXzs7IewSY
EHBPLs4n3YVNJNeWDS4c9XsTs1ve/9fI2DqmhhaTT4q1av5oHu5jP18gK8qGJnfMkrnW+MsK59O1
zCdthvGAxur8fLRoiO8W9iTnMM5SteR9xuiPMdYbKbnsQ9ACy9mK0aLm86mmPekbZCRFeqTn12XW
COjnnIY5oZfJgiZdmwUilu28ggRE9ulpqyegJTlbzQjr2TSMdOTxykGHI6r19UgxaNU0LOeduuwO
dI2/yQj5IfHpBfLvcxngK/kDnfs9p+/KmZrwSH/z/sq9seIntrbSyfCF/G0MoQARo9TVLxwaw+Jr
LnCILqdGKEoH/9bWmnyO83TfcHmAkEoCjp5ahFNtRDYiK2iTyz7GmTLDXcxmiNCiUswTST8n3wJe
LX41kZ/O9R2dPjtvtxM4fNp/sxk4FVivd79nVmHYqjIUFj/tu4sjzzVb2RFttpk+9Ow8RmSmP88X
G9CASuROhQlB56n4t7JAUT/no7uDu11gUVHKJU2nKFVX/6ZLsWlovqn2oxULa1Fp5MB1UXIvI5bF
330eu3hSCoxGD8J3JfWkDE2G8dqbQEhhQaiUx8vg3lx5M4EXjRR4sMq+6MYRmjBxdGGOfmNoVbg7
VM2y1z6tdx0S3SOU09sKP0zg7lmNDfciQtWzq+Gs2qWhiowmynvmrsS9raNIsRCVtAO2k+T80sie
olhSNUmWbxz3ACJhP3s8IEqnslw1IbVwv17S5HmdmWzRXg4NTTvwuIyGQ06BkMYqFFfAV05u3TQC
vgJZKJL2HGxC1qRUhi0M9+Otav+6qVBOwgmry/ZhsS67agbmGr0RqvTtJYUQciWbfaBR6R/2gQu3
GeoNwb/E8VGYrnBs6ICLiR/f0DXu40ysh9Joe2QTt+egns8Y2uCvTutMGE4Lztg4aa4llT0H4A+L
zMMQH44VduRA3NL08VYUNWpl1+ohSY/7kpgjPvhpOWyltHNWbVRW/tfOIaIp8IDWaxYB5ZVpSu6q
kN40hgiSMy3VDi/1JA7QQGvdbrEqUN27jjMOQ/YLITQcmsgBXgKzP3fmGc49j6mdUzRqNYWTQtF0
gK8kTzbGY+wisMmqza75hk1Tq1QVPtxy30eiD02hd9HoU1ffml4d2hqGJM8kB7T+w1uVMjjtPzFc
KOsf15Z1369Vqler4eGYQl2SSlQhZHiAjot+rtr5M1SSA63jQFN6D88/iGIBLpPJkiBv0PnU8yas
rXJJWxUzOUPkKZYZOjMLcHWsHP4MUl3x4ak6YRsZDpSaC1nhcRIjZmqlI68HmEt+GEHLlOKHlun5
2LNTvfLf0lrSaai4xpDNROrq7g2OjOQjNRCSoQ5MD2ZLwO+8iBNG8u5Fb3URz5gKn38IjoSPpbt3
N9Fy8yFZYoNxxP7CnB/DWZpsb7vdG61yAtuGZ8hNwqa/50YjcweY+5WUgje3gIvJj3Wc7GMBucFx
veRFN3bTJLBGar6n9C4un/1EWTDBg+N0y8bHfSkn5UURC/wyjibMpF/mAIBuqB8jzfqkfUMR3zxh
8wXFdXHO6WEVqmlUVcGuH3K0tORSVxb0xe6PIXnKlIg4MZdIJrqncWUtIpZnvNpHBRDAmgTl7Zle
E4/BmKVbvRSu1lo63MmS/0Tkd9spp8nU3CKQkdaZNEyoWXIsXnouUCkNn//EIqcqR4Hsi04tbwqW
mfkwxYBj0HMKQQL3AHWWJVNsEQ1lhi+g4RegJqV+sk05KPQMJDFJExoEFYodQdm2pcns+cRN1C1g
JuUkbP4uxY5JAgqf1SlIAHoeEG2yfRa8xDsf3yvD1cYVB1ZEGi2hhd/eNvG2kz3uM0bDWNIe7oG6
bCJyZrDSS6ss+XakcHHLLYr/sQZM8P5mqNWUHAd8CWVn7prY78xNXTeBW6KfCZkpIH4F39aLOZ4v
qpnkGkZQpB8Rl2Tt06f1jtbZnWpktN35p3+JkanIajICHZ5+VvlqKuEt0IXoZdoM2ZMuNe5BCa4/
QU+ePw6i8Ses3rns5UjW8HMnYXd/y8l379CxZ4L8Op5xIXph6LcQqzrvqmH5Q93SVFfh0uAnx8xt
XJptFBji1iZqyDtqNUP7sfLno7tOItY8Hsrg/3TfD24ebrctQShXzF+DfhQLD2wS0G21QAaQiC02
u9kNrZzstuYAD9WWXuGSPA9eUwGMbX+tvwKxvyhWfGF4HmSVVbZRRbW9ijk/vQukAfsXw5QSGZsz
PPoKwzI75hASkXx+DXaNYSjufKwX2tOFEFi7jDX9t+s/4j7QMCcqY2u9f6R9iKsQp3/Ucm8trOaT
pJmEyYqsTxUkYGdYy4AWcMb0b80k5Z5vGov/sD3C9Tv3EUu385lNOW3Y9BhtbxczkvCgYl9bI+J8
mM/NYbN0hmSs03pI6Ckay1Sc8bzwbqKVHojhHDllW0hiNF8i25/I1HXqtGQOFUI7k91XLvX45iIm
Zf5F4p95bqBHblegdaB7h0wlGbubg08AH5OQuwTHkbOzx6jRuxpJHz5zFjTLSnlB+ut4aELdIyzM
5jO055umbMvasIOx+uHZ+YXnQ+Jv5JYitAy60qiTA/eRzk2Cw/nR+8DdofBWGOR65Q+NMFCmtXnt
xiH/OUiJWKjPjX+vrYQVa1dYvwrT/0evtvZQK086PUN7YoJ3X3iBEpDw4tuuIVjYSuRI2EbfcRSy
Gwgs4VOjVano4bdl9jjn+TRfecrplFcFQi+/asW2Vvcfq6s/Ccf+ZvJxMWMgYi3AAO0Q/FXmDrA1
5tH188ypnNAhObbuozPdPKfW89CiTqfLmuFtYCHZo1PiNRDjM/Ry9Vxy+sBNHkpi4OztDYEBBulx
FX++BVV8K3wmsYC64kzhXSaVTCMqFTNRQRSOK4Q32PWvMMCUn/cDbzQl122tN06uC5imyVqSOqwh
/vjwqbfOwLP2UXUagsjfwEzU/6ay65RNt/6o9uVqBgbOjzrN38tknnH2WlYbQJc6Hk0u/u13Le0P
neyU5wbY2sQx52oqO/Q1YN8dn8WzvMdNWdW0+aDEANLacTGHeC9oy1zvVk21am3bjjxKnDljv8tu
u3bGzckl/FordvqT7P3Z4yDO1Hn1iQY5TmT6uNpL8VCt+zEIGJklrpP0LW8LhqhlLHOMNiNCb/G5
lbWqAXFlX4sm8TpnCOHOoNRg6nmhzAFvCwm5R/VFgt2wep5tKqD7Ar0HT0rNTO0OLlPYwOd8fFzV
Ry8Hza8U1snQzkTtPGqeVzgLhZydlXmnvIXgI0rYif+SuDQjkKWZRhkCj8hQvJFH5r97KO5CWY/7
diyfNMFf+zOo93hQOQ/8IfbeAO9IKuoHNAVfzqu/0Vyy6gF60wd7vODNGHuWmZhfxyHbl/8BvZuF
8j8rflFl+CBVaVldj6IXXnttnHG4vLDdqshDOIgfgG53XguxIdUiHo0haumFNVdogKDEiReGVVCi
5VlZ6nS3ErS9s6fwn+q77cMCqTlRxneLx1jyqb5tVoyZrC1FGY5CW5cgGJFYAWwSTjXwxXgVOQEj
RW042vx3Wu1CL/f1M+O1aQh3zNNV2wAoZG3G7FuB94ZVxDgz/H5XNBO8Rhrzwg/LmMICWiNg+K/y
tmbRcRHkZG1k1xcFupZa9p58dwloe0kymaEsoD8w3n5mCXOjMLsKLotP/DpF8/EEyHz1zWg0xt88
//Q0S0a18SPMzrSdpCH9QjxTXCPf3wQv+vY+nOlLPnB54Lp8Rg/eIsxLUC/+EqwGMKf3kkHPfHmx
agnHWtHw8BO5wi9nBK4Dob3UKkeoQaL7YByjGib3Jp/ylHnVviR2NlDgbKzbtDr0EEuya0zZqWpd
pxTnzHkc4Vm+Z7gu+4Tw5Ulk35CuF+JrmMsY1gxNgqhrXptqXWwTc43XBnsboTTnOQ2pi4Qqw38s
H/2rn0W1d3YYTbgmcW3347K8oaKhKmkx0G+nFITOkhMThQqjeFUvzZmoD4xV32Og/vVDSS//0PFO
vGBpkWfzT30f8TEvIJRMddVEB3ZlSyoi9Xj7w9ZGcAnzdP8XyMSyQ927UUnc3dYoWJ7OcdkjgkW1
pNIMyzrU0u5zFY9/Fg/sMsolCLn6i4GrCu41d/hNMri4WGs8N2zqpAAZanAkpc3WYSw5aXFozrhi
D7nPVo1SZWoQnmp2vfvXIDSF7XHZ82bhiQCIUB6hBHd7D8sWFivOhFUvWcU6GKnsDQsBYjBPdZXc
4rNJudMSnvl3J28hKQlc/TLs/phndSil3RN1zMDFoQqyM8MHNPRKSof0LIzbZ6kEYj/iOeDOYVfb
zjTZLFMhITQIW0Q7CI30wLeahE/QM+kFSHL5DlT67qKF7QoZLGJzv/nwUWNJoljcTvB1kArFYIty
Gjlc+cHudJcvH67B5Aiu9Kv1xDR6GP3KjbNdCMTkzLKshY5JQtxtftABMKX7dlymdME5VYfNH5bC
S1pdEVy78FFWYRBdg1OoWAch0ZeDeNF2XJbzWB+6tdY4oPfR3kz53pVgR1bYVJbxazJHhYbz293L
nr7Mv8rouO7hfv/1dldVmWZYxEtpp6qccKnSUJiEU04rtd7JZBY0/2m9prHDzRdSrWcppDiC/9xx
n36a7DxKx+jF9VOlLGaud/ghqRns4nx/kYcAx4cFLB9jgvqplPJPIHDDdXmTIPBTehYfhA4hkCSW
AZKenjgSuVyuoCd80a4lI6JaVi9BqmZxyvE8ySl/kFs8GlZHCH30erxztg3ecLTtRvTt3EhZ0A5n
ORYX/d8+8YTJBRmV34BzxXJdCITwWEjwNkPms4225XVxsa3SZ6Cofl0OpI1qoSQmyxYaoR3ZwSKN
PnuRU6EILqggga1LLlMHbetqMzVa+cyLU1nMglvGHyfJDehbAaFpVCFdl8MI2wq4Wy+g8qo0rNaY
TaodUwQ1kEV4NHfhBvyGRrnZRewL+CjQs1iRCOk2hh8N5ysl+8/YFhyUrja0CYHrHOVtO4nFJXEc
SsK895EgvCbpgw7ufgyxFr/b0vpG397O/IF0bBYb0skGst5NUW7ksWn5UuW2QEW4uNoH35ZaVhei
LKOZGrhGyZOD0Fei/arPcrkqB452/kubHhbgHVJS5yR6x+6OgivQKO7YMeTEK0Ldb244hVzCWWul
LRYcBGP4D8UI1vFnBxs0bHPTwiWHBCwyDLy0thBTkojOZyPykbDLa+8Z2fuEnrQYUdf69R14fFla
AQaHxitDMr52iBq4NHsgHPmuvPdWCSoG7JkPWsB4YUXK1IiePwtgFg6qTExeWix5VhbMyDVtzpwj
F5bsr/iXXj5xk93T1czhOJ7pF1MKfQGqfxe/40nMFOgxoXfD5Fu+GjvOoyLbHSP9n3Fl2Bj1o8hI
DIsyVOx0LY68bRDsuGFyTNYoKvG29KGbb26d+75uk/BI6PVYQI14YzQ2a2nTBousmdIMRBZaJlsZ
+nEdetUBOeP73UuLP745E0yaYMj7vdV5VSMCIMNaWlJZBIJrWAM/uryZLxxC1BuNYtuQrPBJSsCt
hNy6Mkjp+5VMbVfjG8GJmzQ+yIE8RbeUvKEX0dvgSFGex2ggqgAT1kq9HStNp2YRkgTXia1IyTnD
ALUaIlkdEA0Q0HPKTEP+S6soxXHLIMkpwRXH8j/0re9CGT8hlBZMoDmJCUqVXM+xPEGQFGGHfvgL
Qdf1w1STVezf4YWGLcG888xxEvYDl2WTPUnXNOQTtrKu7/3l7XZJQ8OmK76HBNe2Zq5jV0uYth6C
xpUWJzMV0ejXbSiTw4k9fJiXcxxPG+PDVX6Vj5bYKkjOd3NKLunogyJYS3U/DZD7SYYpxA4RhbOW
NQfdyzxk4LqP+ifAedunM0qy7LXHG7ZkEnYhdh0iop6A4QxNyJoCuJAQfgpqZIvBAIlUDf9zo+D1
83KAaaRRclR5dEYXbUa6S0QitPGq+tFcgRHsTqC7U+cP+HcruB1kMzO3ycgTH1Gf5tJcwz7cpCUA
Xm6RD3ZmDutiosTneRul6E7lFUSoYDLetHL6hukGr8UjGBIlsmekPnaqdIW0HI01SwVdE98YuFZX
AYkLg7NyoisLAW7KHraVBPhmX1vk1W6QCwmzZteJfM38Bw7vTYH8mw1lwYbEDWlyXPbHMLFgHbgW
0PlKh7JTlSerQu7LILNW2WX1ysrh/eq+YVagosMWwW8HYqfbfIryjDFY0mAVC9kR5xsPPBoWJ3/S
RA3ES9gp5esPCwlpRpHFpCFBM3UWyNEkSnK7DBIY1xDMGp+01/hYMLI8KLRDUqKS4nLL55qnq+/K
JsR95ESpMxkVPi4dnY49QH6rFdS9M+Bmkv6+jXRj4iuzq0zQn1luhwnxs5/vSF6uLeQEiK68Yaos
nIlB8lOh5QCp2Qbsz8P8CHn6oZzJsOuKUt2UtW98Qy+Bq1WlScLZ5p1klwZFBO8HufbSSSma46A0
713jREyPm+CXbyEcIZ/pW95qmF2RFpbfPQApLJM3xXFd0qEQ8VI4b1if1V3/2RptqYXu93laIZt7
aXGqyxvb0MKF9PhiHhzrtotR4P7e0zjnc54UrcKjCRkGdRzIYMFDQbTlTNhoxUBr0HvIiTSLJC9X
H5fb2hNSF9bE9HhvCH5VoJBhgf4llOKmubUWpqbH0VKmPaXvsR1zkD0nQQTEDdliJaQxJoWn24P/
p3XcvfuqDDp6zvT+4wFEpei1CGGcqd1LTz2g15asLdyatPHdSiZwaie1RrSCOAbt+YC2Jcv6sF8s
xkVGaZptFZoXLBq6lg8QfSgZD73FDfv+dATGDuVLPCxCJbX9K6uIcUo4BL/IBtVF+oW5f9HFJQ3U
9j4LgBWkxg8uaUtNnv4YqyhqWJdmlZxnfoDJCzbKJbQgXcedW8bYvViOYGa2HFlTLQOKoXeNL/Tm
JhFv0PcUs9tbtn172z/1l1SJD+vol9oukTIgzzKPTg6dP40xkswtZhbIzfAlEn+x2lEWypcbnZzf
wVhRx1gX/qV1bYkXnweRuW+A3GZflylb7WkI8Dbyk63sIuk9ZhPcOoUs+n3lWfxcqQchcTSaoz5z
BoirjVJ1xYr1Z7ttTR6dvI+rGYLS/Wv2XGQOWHc9xyMdI8d3HNlb4cmj1MMFStjKUmWNUyEzQKS8
pgTlw01BbbnMLBewwPbk9d7Ma+Z1Fr9PYitIcrxw/rEuKA6o2n5S7E/X+YUUciFKqOLhJ8f/2B6z
g2RWxcd+5R8EF3Wsyy/Q+46DVrCm842IDHRvYnFafQAiBXGwPFPMCPHJX/zcJQen1onQgQya6vqK
AyBaTS65dHnb9/beM8AiFoAjQM9UI9m0N3cLerPU6b+HM1fRgp4SFyjWSZDxvZn9SG6YiSPutgej
SZFMehJQw+LBWnPylxVOspHe6pAMr738knGY1sFvUpTHB27dqY9rXy0uX1xAI5Pwjbk2vDfTUUSX
QvUQSYQes5ZVRCuJR8dCllREGcEZ3n651qymvgQsKXjbVNWZaLA6DFBHTSuXlVHyS3t+KH8Bj4Fg
jHOY762gcN4QjdfY6iz/RPul6dqudMb/mFhjsJRYXPx//96xCCjyK84Ns3XlNr3Lwg3OQ5LDP6om
rguTpTk46LO54t3W0mGxmW6yAacmMUMaMyNn8XBEH4GnCHLuRBY06ikIZU6HpSOhJYKZBINzhHfF
uZkcmwXN2f72TDol0uZ4uH4iLMd1KJUFWcxZ+bJDtu1F30zkLQgIGsijyAA6oBB0EYSGPPvWClP7
Dyu3wvQCXgQPjgbXP7UuCclQNDLneobq6l6pAlSlloiCayUUMOmp4Pg4qOs2ClTDYTgd0wDsBzFx
uJv5qHwn91kAzu1FM0FHgbjczJUDNEIj/Veg0+gaMLI+UAsWQY+vIgX/s4qZK12wJsTUHAo6CZoc
6fPx1dUARUGnokwDV7wtf66XtgRgJkXI2t/U9ap5TfqtXEOmbyVa0sPZnD3j8/Edxh36N5M869RX
gXq86fkGQJxpt4g9OdBEddaBPwOeGdRavfFATI/UGga9k/YzykhOiKzhzHx4DovQrjFeJI1TwjBS
64eyQbXmXzSVGE0WzpK71FPSACkTKXZwNNo7nTQga5Ot4Gfq+hAzggYO0tS153E9YywAHh1GyiXs
UXvaS3r5W9B6IAfKHqVwG0W1siQC2mjHWSQ+rdizcqS5C15hckZbbbVVsxKUnAL0YJ7YjBtw6B0Y
FZaxNGaTm+dR0nigl6aGq9fdRLWT7yPxJNNvaO2tlBCggaUNhM7JlEnYcyafpHe7q4fKEc3wy5b3
5CqmBENDD83cCXmDZdgerDLqSEK3HltLBoMmPvP3QeyJZfU8D5R3Z+QLgd8DUtyhvRHCIoDsnw/i
47ok9S4asmWZBq0Ybj/XPfw73HHyScxCb29XxWIzaJfxxvAafNE47Cqw+HZ/us2HM9w4m4bZ0UGy
RPnKIA51ktbhVurKVRO6McBHORoUiEtWiHcoo+uGFKkMiCB/C3Vb6mGm+R/z8lhuD0cp97Acuj1J
UksOu1TGseSSOWf/A4Y5GnqhXWIKNirZhs2pJl9rXO109kdtHyM7kFX1vxEGDAnVu3nyHkQOdyPt
s4tgYRUBmy68URi6ny308ImGgAKEvl+ad/ddY5IAi7Z/Y0PaF9jceZVCyyPU2F8Pu8YkckvdbFQC
KigfzK/2QEowYZ81r9grCFfpmhRZ/Rg9oqFT3y84UUDJjFcPupAOFi1p+RfuWP3+LLjQT90WaqHe
58QJohR2DVaL33MXf0TUxGRiEMZB9b+6jMfnVfcu7RkyB6Ryrv251SYUNY9uUn8v5oC2IGnLPKik
Q9sV6RrJBB2KxX+z5pM2voORWd7C6IiyUxor8nUtDY2omw8IqAzW1i1BxqYgFkRXsUomiBDzVT5t
OXH+zH+MeoLLvDL9p88k37QxPOe3otrOnI3huJeQm/Uv7pURqS3vOYQrwnQjgn+aGYepm4idBpqG
43p2okqLmWqVAcvLRtOxDzPgYvUnw8XexRRE0aG7vu5PHjzaVeDlJdsT7Prf5lOzonmm3AHC+Zb7
5CW+MZ/IHNXbeOQzGjzP/HouVE6fzHrUEjQln2B4cKyT1cnH2ztcOSyl2LDgiTxOZKRu0UC5VJM2
/7eSIdt7AyMc7AzNBRhwvemtCaZ2eRVDl/3hYp84ZcJCEGLr7+GnrnVgmq8m7/0gg40QaaPv601W
6E1LEMW/gdnmPfzqamhQc7rLnFr7h56wjXMOYONldlgseiEKbv7/RDCeZ7xa5gUSkC+lmYBAneHW
i/E6oSQBOrXWVUKs6HC6LFNFzKRdkGqmM9lvZ0a3ktPIYuz/LOOVe7LuNwZdGR8SyFwa36UBgu2H
HQRTVxVBoTTe4uzhPDUG/c35T+CYrb95pdw9QaJ8217VNcrfbYQnBioJ410Ci45ufWfzUbNpMFrD
32PmURo0C1ozCOB6PcitSrjhfMuEH5XxmQ6C+01yeYmZfWkvalrkFe2FLi6lXbECJ4yWOMPFeA7L
eiBUjgqV77zIMiw/O2Eku60BMZfqQvQj0dcme9WvQNa0WTQsOM9sbtN9+OVgxRmVOGakQcQMtw51
l6xXEYlR7jOB2GIPz9MnHVLitY/6ST1wGgV+OMHqPjSdEraSJ+Vj7/EGfmltxvp1oe0Bp/PnaBdk
uujOgSOVrAUlWo9051iJ4yFWrNx13/AlMmAXVeTAu4HUm0FWVhlKmc+K70gRgJ//KQn7DrUk7VIr
1hkRI/m8tdXEJVjaudu2hi06mOmOBf25VFTDIetmZFwRO7fovUZ4L2eCNPFQX9n2MNvjwKZq5KKe
laH0i0HaXdH2eYHHBvigOWjo5dxW7a3PNO2vdf5GYMLoKFk9chQRebF/c8QNBpNlM1OZaOqO6z5v
5uOhL365O3syRgmpoiq4q8YY9jlYlWRTz18oT2sf/zQdfqg7R1jH6oH+T3H9dvjmzEND6UyyoyDK
BFctiNe+rOZOPh8iKRQFXax+YxjdRuwD38izHmXZeFlW/hDTaRhm2zroYcE2xkXnW7DgJYjxrbKN
74VabYvuSvwczKNlyRgzACElhrOkSByYMuX4BjwaNP8K/OmpJxZrGtdT3Y0d2MXkr+34z5H8+ftk
5lbN3podK3peaZDiGMKUGFYXzk8A8mhhMu/aq3FDcB0P5G/p69Ln9gTuqf/TXRenKA3r5nMt80hD
mXFvnEOA9jOdams59Eue92SyxZhw4CN4d/15HHi+Er/+xNB02/FBLofVj9GZ1l7f4MI5pG1748kX
ee70C+i4m/l0HAu2byxEVYFa978NxVfGNwzChBbKeXRPjrj/LSg+eSyh25YfJLIfngTVvNcjRG6J
3nSKZU0F5bTfu2p+TM537/XKEV9eWqX4PgFBvCGyNQGohR1zZB8Ugwqb/zANTONS6zqiyXY5cjPx
1UIDhn5VyVcqZfTPWSw4Ezr7Hjjdo0NE8d+3+CVkxLgQUbrh0aVitlteNCvVvcUwCOHprPer4pkO
1Jak4uF70yhpr8Ch9C2k9H0m2uh/mbtV0QtLkOE2sUUcvoTispxuIXvhfeqJRbEd+THdfWHzVLLZ
i4XEfH+crsyC2ljo17Hr41FRMblSjGBe9mArXg8OJzkaD987c78tubuyY9nLnTOPK24jUWfC9KDY
WRA2yM84N45HwqG+55Sa8XodGlToS7TIQWsfnkSvmzy3sdNHL6adQNfwF2Ptqy5VBpgqX74qnThh
/GtWgspor7J3cooGc7aw3CuJjbGW4Ydf9wRTCxFhlXIgI6hTz4J0bTLlQNxQH3PAyDSq507PoNkV
qahkEjUvINL/QAFUJHYh+Zp5voQvWrlXP6EgwrxYGJzi3rdIPRST/3AMcVVQGnhW1tBf3moEb2w9
cAr5tDF6Ys4hVk2/H2PrrA9Qf6A1Ny75hySlHqOd/IaqDNqatpe+mnzZeE/N+rGk6G5bsnWt5Sok
TLhsU8U+tRZMRcTQY87o+pbvuWG3Bz9iOR/iVHABELMUA/Q0KvIhijQYa2fsPglRvSNkd4kjYzsr
eKfy6DAtVmtHhxQa4++GtAzr+dNbHpojvTTBKDb0iXMR8NW9A5cRWa30Aky8gdeid7Juup46ixKt
dmttPqiBLRAbwZVUyI5wg5A6wi1UECuVsyluqxez9zCmJtBGchmMSHYScSXcWxfx7wrzrm4nd33U
8obinSOQh4dYxaB/vntkWNyQzTu3SpLuJMnspaQlysGQCu7emgPVxIntVpWll5hMyatSLeLMB5Se
3Xp7mx54WmeX6yNMhHf3gkpvaE2/jhi/dk15yvBOwD1Dp3FNcKIcvnUm8EVo/Xk0FuS5ROlqXEMP
YzqmaeY4xqhK81qYA2TL8GeYCleon5hWkkvtVGRa8DI8kj8K3P45KVSS7PmAZ7Cz2jmG+Eo4mjo2
NNigcxyv0GPb+DYlOWRhcFKD/N04o1UYFl70144XyunZJlLW1D0B8o5cPtS/qCM7YpjZJECkEWUz
yiPknwkzI1PPDftLMTr4uoe1McIRqgTf1eJj2slfzfl4DCUJ0weTyFVgh/3bRiuhRVNdSNDxl7KG
Y/+11JtTidUhD4IE7RCZpkNKBmpL+SpDkF1ktZ8ORA0mZuHb309Cyyh/HeyAHkOIwHfRxyZ4oe4K
pvuKUISWfUaJ0GXx4umhQTMmOBzg6KyBbSuRuWjfVJGkThMJHySjS3xGyn1CLjrtlXz7Pdqig9Bu
M4dsTy1UxwNlzIGdr88bFDZ83UWD/vLNmv2tc5tXfMlGyr05YQjjVHq8BMxvlnUpOHbHVjGLKGld
KsnKdacv7rO2toyR1BpsE+r3IMxdibf9PP0vZDPVD3laPkGp270l7YKVNqyCaYAr2wZ6O5PBGJ2p
ofHu2EGlayEHc0K/d2xOX42kEwYg5dlUgQHDL96lUygMvY6Z1q3TY/2CBWzhtK0IRgGlukcPLRTQ
yyMvOOOOa9tkr1TDXyGK1URqMV8AyIQNRWJmvKXN/4k/hDMd5Dc3AVH5go00pcGQs5mW3sjCKNN1
mNORZsuPvrxy6zZhOwOhWnLd3ogdrZqF9F82REALxP/HyjObzUgoni/ncrMBiyunlF//WD5fKDM0
Z7lLtISnF8DrYKa3KVYmr4DkXVNtDD7CaFUjZt8cbrZDdUmy82Chb4SlgAKEr/EEmvX+sRxHS/OW
lOKsnOFnaxjFDEXdP6/jhb6O/+CObQcbjd5ntMGFB0z0COfyHZE0gzIlOS3XWa9K7uy/BzzAVjkH
bLmAj2RAZBCuDvGzjuRvupKuhpRzxAFl33F15g50jURT2gMl7NbfSd5Fu1N9MaFFcLYl+W9WqECY
bOjIn5NBgKR+rj3HTeJ8bSooyEux5mTQuXbr7FTpWD9zon6RlzcpfjuiT7prjZ3YRfoBwU0SBi2i
ZkmoFOYYjbHMiW5vWFfX+nnabbPY8tMBCmGO7zQzF1002xwJtycjdms2ihx/VBhaK1ikoqNEHoBW
MLYnSvUPZNbEtWkeCY0+w8wBFsKfr+Y9lL1VnTzptjVbmqLDz2QGUi98xVKSxv8HoIxosCuLbkcf
zmIxyM4JDT3T8e0zofJY/3pA3GN8oBiiq85lNXntzK7BAeyYR9H6IXlrCQCZbGvRGgoqgayjkPnP
T8Y0bPcZWtWlWA9HPJqQkAdRpYjaTaMl1wQ4EdnJRNN3bTFXOaCNRPgqR7AmmCZ3bUqKhJCNq22Z
q8CSF+Cjg6ssa6HzS4ef7XLUnTHCThnz2OE1sTshinizX+pFBtgJcUlCs+TiT0EOVv4iPVe7ZcEY
MkXrDomZJ44UgNwUPOAR3T5gs4y+/7pg1L7aDm1tdIYQKT2steGhUr66Bjdqa1nyXMiJRctPjVfI
4kX5WgkVAuebQrIse+ggfWDPDzEmSS0ehKj4GaveyhGima6iAmXh8ndvbgSD/tE1dkEQcIBkQ2R/
99W7+ZQB8Ph8rogHRBa4DUOVWTLTDdMIVfHi2ATN37cA7Hosm3862xn8HOtGVsKHrJ6ddg5CXziA
k3lgIgCTazHzLdxWjGtQjgFXNDsoAd8YVmYj31jo+YoPH2n3r2p/hjmctPLLbtfI0C8iceoQEkod
Ly5S/pf8oH92PxzzOuaKhujeHIWt40ccyTRrykwZ6V0vYw41LrNxqSs2ru/AYlE9CWL8W3NxBqvO
e9ucETApxJZQdlpUuzEiD39CTsnU+SKjhxH59qitypgkMM5qad7SqLue+XyvH4wrCRy7IJeBwrVs
fGclA7RMR7DWKT0EtmHB/GmEkqxRSykcauINXLG4eSfgMk+eU63c5/gh6TE9AwlodWs+17cxRfCC
XGVtEjEe4bprrWrvaMbmM1G8GYARylSjFOAZpCHNN2+lQWANJ708Rd03CNcnnMyWfi8pUu4PXCR4
TZ13tKPaeIdKSK1ajnDz3zmPr3TnI6JIEP3o9uaB8buXErdHA0jUbbuh9FajYDByQDWIBggjTyRU
HBrusTJ4KmhbLA9zr0Ki0X4/pVqIVtRJ/0HwG9c9EXeOl2GJxAk8DzvK3prWWPcv+liNFCBXnIBu
F2WAyF4+rdNEoRgYiTrLE0gZwapJtWwHg7YeOzLKHYltxDGQeii61pVia/AIFCT4Txt0gJqd3b5q
OTtvTtE8VUKBjXO6r5U2F0uSTBej2xjCuVJ/i8jyt+LzFbWSm946O7/lvGG0pDoQXNGkh/txpY39
LNwgSqrS9sogin5cpOy/c4+l2pXHcJEcLKLWRGoNUapLLh/kMLJIhNTnipyN8OcfvcGrQgdYld7i
r/ZgfAYParSgjAd7MSwIZvLW8yVAlB4rEIPi0zrNoOVFt9jy/ssGrMWwY+b6txMmiYZTsONfLN57
5mhgAFJug2zkwwUiv2byUnmLJR1fBbCMYLFYAcATLigWNHjpcJDkZhzuzDlUdMWwxgCX9mgxLKP/
KuUjxy1bcRe4Clfh8mMMLyP07BkQ+LyvyYO4EnVQGid0C2ahSmM0g58OaI5oIZ7qahxD+DV4sz1S
SBm4hUINUL+oVlOKO9dLOMnbQWuyyLdnEe5jjVHE3JBSQuuH0UlKJzki4lFkIl3JCIhGNRjRq1KC
g/8BtE4QfYiFptL4f/EgiVbxBzVerI6NUhqMYRErxKDPK1jOnr2livmkrjAAm06xLtKoDx1mmsRq
E4lseIwbyBCYKHuPr4+2jI/JfRPva0MelTYp5LyHXinuqH5DHt18p7UW/uLBwa+wzyOWhjk5kf0c
aTGHzyblCzk5uGc6kgtNl3/bmWBsacIJf6WnpSp2HUAYeQ44LRc66tDNfsU2SWkfZcVpta7zWaXf
46RhzgXKK6Y60TvsiiJzKyhgQY9Sd2V+kdA69QTHhTRRH6LD5QthDnpVRj16ds6TeLtjD8ccWqKa
4hpoN9B42yCT/5511QSA/PVwN2nsqDkf5moG1rd1E8nkDF8Pp9yJPJbQ/6s8d8D8qxw1sWt0ffja
oDvyvYQalByREMMfL69VCmlqLwMFqU50y9aaLzkR6brfD5JHyyf9i3kqS4whDczbppFkkHxoqh9K
mz84tKO8ZB5j2h94Llclo+4MelqT1ThviApmmdZqX7n7DY//h288VlvmoJY6c+wQPBoZZUFFZ9xp
BFaTrJju9Rhoy+WW/czIx89IRm8qt2gULH+OqDvAkNDdlcCHv7WXCtB28lqx6E6CIwnbDm8m4H7U
ZsQoRyu6DTV7csTXa37ZRrVWAx8vvZX2Dn2upCUXfy8qKyeb3XU6zfQJgVTFyUGDbOuIuQzNJxKm
nXLy+C/x4AWiWvRLvsr1IHVj9vbjbQkF7RvLhI7G7vMeedHd02o09FnUfJo8ebjzI5pZqrZ7SBGD
7HGPdyaCV3UtjfxD1XBGxk2Ic1NFckr0liCzQrdDMEhJohrjnnI/lxPw6H0mbvTgfP/hsnxWd4ZD
5IT0rDnZp4pTz1ca8phkkBwFDBBdpxRyBg+Am5cdHYG12pgPMskz0jChBX6Sbr8BT7c+9nuftmRj
/+qSQza1JR+3kcr/Agzh/MnyaVnmGk/3ibubowD2MLo4VcD6Gv9jHEQZ/KpucvuX8wOE4ClFNydJ
sDjy7jX15qaHDUM/nO9aCXjCWHxBFHhWxy4Xlb/9B83v3aMbpzkeUs3pCMz8tW3hI5r057OHv1MV
AYt/Ri1sgPC7Xuq8jqnYgcvdd2MUp+xpHOKOqdFibTbQz+qsA6zRg9kZpyaC6TxvL65x7NAs91r8
Z6GIrQ/CRt7MjLM2T41rcw32CorhFFyR6PFlnjrvFzxz0tZo+okf9yK4xLwD+ZaYazc6rSSLdnCa
UX/W0/7pTWHMqw7WhxYiS/HbZUBagAaoDAG4aT3K6qNyGRTZ+EK26XjG3dVLrOtMNhgQahg8/mKy
nRFyu0GJ9GVxe7uTGAJKgE3miRZ4Q0x/SgFj88FNA6gW2OGwKZSo/eb1bgHQwK2wHMYZzDd6HY+A
PkGBha3fhh5KZjLQRTqpv334WBv8ZV5JNYRZSo4glDD+8NFNH+izvaejJrM4qivU0RlgmrCx8TSg
Eb8cF2AdQxnhINpAhoHO4LsmIxwuBKGAFCUIHMUSzQ7rXXwONsQdRChQ8fv+Cf3cZPtbdJJixcnK
fY1E0CGsW+1i9fIjHF1neUhj5QJ/u9rKXH6ZAHGo/22rHdOVHkJ8PIMkt0LRjYOK0YI4I9FuUGar
vcs4ENSHS1mPoiOHUsrDlWnpLkifslPCotg0G6gzttlX21Q4kth3KyDx0NLunIIkUNFAlwvYDU4I
yNVOsKySB+pCs/u8XiHU50Uu5fw4VM7zOac2i0jEcXPIdMNP0pb/LRB/KjX2yyebU27TjHoBmr+J
CGViZxmbILgUXfM/Px5LCILxFwO41zsVgo9h0R6MRyIj9PqJsxK9Cs6rM8kbdohUJ4q/zBFxHhSQ
8IEp011bv/BWv8xWo1FZ8glFsW1xw4x8+1e7kaCltDaqKnsH/aMQFEXLo069oArBu58O/qGpfoBg
3tCyXiJdbzl7z/U/9VTUAUS5Ipc3bP8edvIkFt6aDOeznQsOirgrrjxvybwuaFZUOD8FWI4AtMiv
+G1MuX1zfyf/HpdZ1CsghiHkXfjqcBbrR/YBvk1adwiTCIs88dKWcMMzmOXFvAyweewhcKZYYtkq
QAhnygKI9j6yJaDq3RHALjW8iuoYUtu/L7z7rCKPwnMFFzjBexyvSDQG7RAtdXmSzc++BhJCQwWG
Oh7YnvquYu2ohj6DAfYTK9lTRlbLrJFz9ucg65f8HGVwbu89q+6MilGbdFJRA1hBl4VKUdVgKUjQ
f1nxun2LiP7wAM2EalbgxupV72vHTrJMEZoOHxykprQ9dGOS0CmQe4ekpf4qLq2Sev7/yc+ZUaej
vXSup+NfRvEHdYDBKg9/H2ry06D/WK+OTPztesAqZV9kGm/SvDs0LGcsOIGOpoEqrmr9wJuENqxz
gIhRwBo35jP5zRTKrUGqIyk4hdEKkej5OINHngFFQODNopYeqxrEvfmab4ZzQCI7FoYu6eHGT5bN
F72qKIyXZeGFyCpmeN3bPhwyOJJZHPK4K8cpKyV7bXmlownVk9CjngXkYYOOrx37sbt9JL6m/7z3
y0utIrZbLFgyFBDqQOIs45PWl9W1NZ1ryA/0f8WTl9y50eucSlGR4hui+TFMcFAWqHw47YKAo3az
p8VsfcW+JR9Z+1wl2gy/UjkUlzfNupmfInLQvhhM4n3m2J+i+KjFwxuxzMuCxWO0qu6IK5/aaCNG
RMxU9hJvQVviOrzFymeSSDvhuzmyduOrN7j1SSQmqY9v1mzMlYlNCxbJGlsgkNY2KspMySaLVcel
jteMuibLerCndObz5iRylzzapFHVE2nelgquVADjutAxff1DJdXgJtW9bUacEzM44pf1laERcLQW
fzNzzQtnrCirraeUTXGJeoh3iXeiumV+BBkLy3v/RtofSG4PzLniVn9kEM81/KvWZ7noTGPfT69l
AjlNdq5BAaTNUiocT30yYzz7WmRmqi3/XExpd/l8Rns5dS3/Gn0THuymhf/85PSQjhCMD+18V4qR
c+uYalqmgSP7R8U+4vpiLKxqsgGaV4QauZkFAj/J7P71XwGGmv/PaNNxhw8cV8q81Zc2XGdpWIQw
NwNDw37Nk/D29f7dpLSBQHHkr+2ZpFAxS/4xwuL+JclYxL4SSkFm/V9m+RExcibO5tOwQAX9HnwT
iXtVSfNSsrKn1MzfpGcyhQ1TV+bh/ApIbjfgmpaMFcCO2oXIVdpQf9YUMWxgGAdfkaMwNbZ5xSeR
3Ojfh7qK5Ypbv9tlsZa7yahV94VJVH6pp5of+poCh4jAoiRIwwI7tpcGZVM1OVMWYpWjf4IyFL40
J/OZ2TwxdBwBG4HOULsZp9X0eNupquVhbQ0MLFMWNcTPfQ20wLETtMuPDU04FK1wwxzbF+G14pDM
MZL+aaMyqotkb9Ikvw2/yWKOvZzgd88O1s1C4JRfii7CE0MDg7+8dMP3afIa5swE4IJllCWgva+S
tL+zM8W1+41VKBij0J3TE67gxg9ec8afHaiDYGlcvYjQVRoXVmLxbrc4K4imo1Jx6rFvRqog74U2
Lsz65JVTXyT25KAdxz2UBNUhhMbx32zBTsWCNoJJSMsXVE0CJGTEfGRSTzdMs2WeWfFd7DEeQV1V
+A5ALAwvLbtKYiAg2+YISwJyCGY59gdSHFnslQ0LuF1BQip9wDumUD/JPFUc0/ROKdrry9PoN7ff
KdnNoBiLhLbg1J7QW0oNDIShHZxKXIZ3wMHCCAtzfR+ER9ykbbWbRpKWs6vPseNlIh4FILn+eiH4
fbjq6LYBqlwVDCO0LFKdzOBMQEez5MsUF34UhIat3/pSShzzpMiyOWTBrp/pNG2GzByEygcVD5tT
QLggodmKQ4F8gJIteaN812UVqZPnGrBjsgNAtWl2sTQWmhL4750DVjiDISZPhR9ga29KLu9bJRaj
LbM0ojcCIfg0OaZmcUSHSDxRnnYBsT3fqg3KjxsIT/wgEGKq9CfLr+61fPEHSWrf7O6vsIghLaed
jpVDxNh8neqOGoZieWmHd5F3VTDtn7K2ACAbX+dC5/1rhOVfoKDuhFHjBZ7q8iH0Potu9EC2Zt6u
vQoRdJffAXKJ6AH4+KOfHygEDkR9UUmXhAK8GyuL1/1N4jcQfMqKePYC64mEi4GfSvR9XplTSmWM
w4cmc1WIY9oPozIWQX+Fi4nre1DffBVkQSIwOFWaYHVoZOfiYVvKDB+9WHNXkZDbdHkxRhtSajlm
Im47UQ2qYIjtm7FgIOLhAt8+nCV2XPx9wWujQgf4jqkHx51eT816yBF7dgqUR2isjT5vXi0slr3h
0CMqJdb7Zu12GadHZ3ngRxECEQzrbl2Hv3/UEswdGzOy4KG7trodbbZPqyAXCiUhYsujNpLd5E59
1WW5/qaOcPlm4MVJ5dSvg+U/yiW2HTrQgFKfqmvBDh4AeT2nXtgyBMPkUTtnX0bGQTnNG0IXeui9
iQM1jsgGyBOdMYBJr5UIy/ihKWsvz34mTJMfIH1NMUR4ps8Pikv/gyRCDIuklgXQ/vwQRjGX+df9
rC2bkuLH0NfmaS/Nxv8abK5vDFmOos9JJqF0yTPgK7cyucaZcpheAvN2vCuQ0xRro8kAhdBAbRGP
UOEmUoaxNPMuuj98hBThTkM+w1/zR0tEYASbdr43C6HyC6SnAvtK4Sr3tjMhLzB7B8dGPeOe+BgY
701GqWCqVjoqQTtdNDS52yAlLWqJDC3fWpo2VqlrDYStx27QpLV+rHOXtKm/FZ5XdlKuPrzwoJqG
q/QfyWF3UxXQLUDDSeQDloiKX9b3/QLPsvm7dUI4iwctVAl9yKTkBUc7NCR3M54WN3vlr6/2vIrV
YvZvfNl0GT8L/0VNe+yA7jcX9Dc5dP4p/hc0xZHFDQXkbPXiZCDEeEZ5wDrfC1PMSAzuMjym5ggf
f/yXuqVBQGiwr77jZgdDRit4lIPunm4T6LOw9rluRE8TrtDInk/JBakPdqEOjRWG+STuOQnTk1nI
dtHEnOBS1vu/UQzaS4wbd9Hlg3Nnk+Sf5TCVU21YtvqFfkEPw/vLPE2LVOEgxk+AmRGtEOlTqvFs
Sr3tjh8h3WI/uB+4hGwk9fb9iHbRpS0IJQigbAn2e/IzGLralxIJURUTR/JaoH/eao9epVL6NGwv
ENuEa3K6tFiII0pq1r7Iyokn61nXwsW+winw/GPVQoIv4rKy/pGRkDekDVIBEFwSIeJqJv+DqDLM
uam6YO56QgGTJNFDDX3iD1BU8+yKU4BMaG4cTQ4lJXG9PZJnLy6Xd72BfKdrU2mwNovPD3PIT6Xa
8ZKRA4ax0bfkSC8whI5tJB7EwJakUnTZYu+/p0TawydsgbjTnQao/EostFSXfbK/cOIJZx7SRXD+
e7v3rcUIzeWlOCFG1HIUj774kRWH/gwflFFhbRbsHPNA00dEHW4hLTqZvzqpCDxgng7VAFnilmm/
Gw29Dq6iv9oUEzTbwwuKa+pCy3xfovE2DXZWBHggK+Op7mbZElWFWQFFRESyp1f3cBLsZXPaRpMQ
tv2K2h/kgD0ekwHferFyt13Bu+tju2bWnVwCkI9zITgYALvys0CKHvBXrDwsO1aUD3J8PbaXTC+4
3VbO3jVW874S0rXTKZQjoIXVybTv6C+u5vnAvGhvpEZfvTIGxFw5otMDxNtp5TtCbNkBUG2Gygr1
VHeoxYkuyFBGGjxkNGvstmJgFOgdfTXDHzNk5U9tXsh+4Ki7Pr+mNU4bJ3PofZNY6B1taJNDHlt6
akUoLJVmaEHeNJfdUQcQw91h1niFchRf569a6A32me3q5cpCGsnaRX+g/FQdSB1mtIF3rxr/Hw98
e15eQ+/VSuJwL3i/ENIaISxsmMliKB0xe9z4kjjfnL6K2bIXJX7kcyIOgoEuW/XW4PWN7shcgZJN
x8GusiiQLFuP4qA7LoUIC81ybBy+O9Ql5E2R/UNY5wsztt7YRkAggaSjFeDp/WzUE6R9hA3u7UQx
Zzsn0KHNEHsdQnzo0nQuSRHgq4t5Ytpd8LTXNjsJa0cdY0rYnWr8D5wGYAG6eduff4F9RZ5F9mX3
wh/XZDkb1E2toIpUCWwu3jWagIeeSsJTVyDdcxucxYBf5mIdNhF8yl45qv1wvg1TesTE3E2DScQe
KrNH8xZuv5uFHUGWzU6DjG77Os70clK9VWzBelFOdLXXht5qXYCO1jUzBA68Es4UlYZK1+9DXF0q
oj3NNlb9QdgUvwnzvbB6zUqiz8G153Ro5X4aBePWFAjI35ZDVev+5XQe7z89bOeGh7O+PPOI/Fzm
c2tL2FdK9DYwq16HTY3uGSCaKA6fXQwg6YSA4MaEK5oLyJJDzt1emIwVsVfBnQPma7V9S0mf873r
WQ/TjqvUwtjxRXg7mzvlWObdK/37I6rsddVIbV82oLFDG5ajm/76vptBh8mcw62nHzRiuS29+eDy
Qqmc8tDGeo8NRgVBs+pSPx763JNn/eBx6reFvsrqbH9wFwLHWG63QUD/KVZKCDtBHZeG41SyhcKD
32/nhEkAQlxpDFC4pDTMVq9aQblcVUQkVq1l1EERCal8MulhmcwEtsVv1isva/lPjyawzyaL0OQI
Csli0WyEfjHNJZopuugdwpAgHsr2JNuH7vQ6y471lk1nmGDO6BEq88+DZ0pUzwYhjiH9LFlUcdGe
YZ166vFuaU9NXX4Z8bK3D0ZrcYWoibNCZVYM9maldStQec1+VJQG9p9GIE5PCjCfZ1wX8OZgMAw3
BWS/bPpoDyays6a7DdvMH18r0e0zdspnNai61WeW8bZ9lfmyXRv40INXTEqOoV/RApQ1XIF/zC4I
U2AJI5M0TyD0NTMQVle1yvy+/xFPsMsoOXoV9Msr3a713+S/DSXYcel0lmtHJ/k3/wXc/A1bAXGJ
NSoclnjkyD3kmkrW1JdSqFRT6RqQImMoi6RvR9Ho/PAN6OuZYnXqlMk65YUyqpOraFLr+QwKO2g5
5X07CSEFD7DiZlG1m7htX/67jS6NPGdZtzHGEudAfpkiBYeEws1VSYIPyV2GoP2nO27duBozOzF0
uh2aZ4UqUMj5O6yuAebamK1s53PJu43FkVGl+FhU39pRxLWk3iEJX5WSyX/BxFW14vcy8gPRvwxo
yAmEdi1YWGTEuYpQK6iJJfDSAa+nz2mBOMHYuW6Ln5KfB8cD6XWxY/F4OdHrKAsiKPjHHRSwi3XF
0a8XVa9rNc4vERVREh0zDiDPZllxcAxhvPaxCjMk9p7qsoZ5VBUGAq7SQOxOz5ab6gDv7IR3bYMf
VrlwE6v/aHayrP0Ty1cOkqxnCSYzOKxQ5FgO+nfxIB5oegOw/G7bfha7BgFctSCE2Y9UeSyjxnxj
ht7Hgmc3XiZXYTMpcMv3mhXihpUWsLo5vmx95YcOBJN2Nd3uocYwm1Nhc8npwYq+wfk2W0tyR1CI
8E+QMG8kxgN5uZS8IYCNyLDle9f8RhB1IkKcRIOOSm3WpB6ZJDEJU+6e1QPVhaCd67TKCAOYGqBf
8NaSEYxvUoAKObXT0v2bZQSKOOvhx4PbH7Q2xqBMK9rL3sHqOwLE8pcKLspfKOihz6UYCDBhuI01
Ou8awOxeGpj5MPe0Zrrt6S+ei4CCRHp3rfNA7PvHRLjycsmgBC6Aq4Nh4qOgw7Mq/rAopkI7+t8R
bp+sYJ3hOBAqSVsMqgqGXGKtiz39DAM8TpeLkmdVMUNakVx5sxmH4o1+3Ob3hvKZJOTY7yOrJqS2
Boq+HVQbxDMigJVoX25CF7OreQrSfD6pzLHcc3DHnXrzxpZuxB8UJkm2oUiNIJrG7sm25gZAC2mP
d2WG963qXS+00Ostr/cbhX7E6/y6GtoPs4arQ7GyCWQOdsukW6+vCO0OkSIrHBym2dDiqVHX34DT
Qos/fTsRBc2gjwLOLB7qd+f2wfM3KRfoewHjHZ7i3rPzjvLTVwqr953xyWRx3TqWEHLAYRmJBh95
xmyqD+SMD0yS44R2QbvrL6YxD8mzYPyrsm9vmDHbH2dVUZqwCrvDJqsnIvsnI4sIrveROPWMsavA
Pas10aodiXfCFQrDblecNoFy9+K+TpGSGh9peyJbY+vg2TvExqlq0TantSzp0TebHX6en8sEmtH3
h6OPn0sMT51jnycE1E9s94olej05QFplFtTXOS3g1UqOnXze+HbrZBe/SDgejw2I7Aw3YZy+X9rT
KEZHP0T6M101h/LQ1ucpMRyBRYCi42ZGYKD8sSiPisAacVHnaxPX0XDi670Db8A/+q8GIcrl33QX
SaUxX/JOcA+ij8d8/NXyHy6mWFhyoq+KXJP+aFhcI6xJE9hk3Y3BUy2aw/+BfcxPdgW/qPvxsfVw
ET25miwUr11TCDpC0wrV12Lw50WXrFJ4D4jo5z4W/5GfcJ/xzl1z8uyI06lnGhPgfJO2rr9bD4f0
MXS7Xtrcojf+4xSxzM3shfescRvB8gr3GI/XoEcmEpkbvwGxLt1O742CE29HtO1WYkz1fl2FgXtT
1zaCE6fhJwjBU1kSn8kV0dLuN8N5v+RGv+A+NVFFeWOK43hz+2FL/vN1RLwpdWKy7QQ+Svc3iXgd
pEqvgN1tFehDbTMfujHdCq3ltTVZZZX6jzilj11sYQ6liTO0i4dOkFH+K+AbgL8ieQXyXOy7KZfT
2oqmxyBuFbg6rGluxumNEfxLulbNZdFyPkrzvTpf3JrOd2Ml7xnq5t1vHILqvvGxdfTBvdXY0oYN
j+fOPFWIESNGFAvFbfweTP12e4KdpoNQCBjc/SmYBcJ0eQTNwQpG0IrSLcQRzuY+XJnhPZCvxAkV
wFsVQzfyoS6jPud1dzc3+iabj9xbf2mtKJKFw/EQhmPpPTpMhLuM28juLC0NPCU16cKbC50WSjTW
5AqSwsykm6NK7sGGDSbmN4GX32gasdofiSszR0a1w74eSIsM8XH7ASM7ai1SKI5v/idiiD8eM7o0
zn91ICF/S4UFGLNMNU970KQUopX0+fxuwJfd2HaBV9b5AbOFswuZN1y8h89pdmNxyCcrf91y+kYg
/T1+eZ7dcffQ6H07OUptgisFaZFPm1FLiWeggjN0ceoTh5wSY7LVjAtqMslwG7Ce84zeO9rXZN57
pIyyaVT9W7xAxYdB7B8pPb/DnUj0RsdaeSl4DUyF1JhcRfirt0pnxh4k62g66lTbHIz9jhtZfe9V
euwprNtATrp1OreJXWWnWETJgWVLKXTxYuVu63hFoPVc//XIdFL27At8/uX+qxBj1SfycxKc1BO1
i+cSYoR2F+6qvcGAXbMxVAm+KMKj0cA3e9+GOqV6Eg0vcMRd9cwGF0j56mod08mUQJLxLLp6rMbn
FgbmFf6ogrQ5thoWZ35nxvi2zKcNLonUIuQVWWSmGfrE4/3MoRMgGLmVVH0Z/LAiih1qVWuM9VYr
gBI7nyFPkAl/POzURMc/E6naPsCZubJobLU4E5iNpIWtYhpU/6oKVUIJTaq1yaZZbAwR4N3QHOpS
zo2HiToHLDaB6PJ1xiJ0tGdF5lGHwaxTravK+rrcqIkX20BbRikfAtMAY8R0WFJ8MLvx/SqdOjRN
Yzo2RWZXvX/h6psEpJv8bu5X2QfTr+fREJu2BuETymCNl1CMn771slJOL9bLPjXfOybsQkMUiBlw
ZTP2VfqWGe9U2WNeDHeF1bOxSN6ebLZ5y5RmQ2/kgvQsCdJOfIgKlPxh5psqSDTCcHK6L6JmZwJ9
CVIL9cbxhgg7awcatl9Y4kUfx3DLANLXlOpDFsWplAE5QEnL6OaFtwVSgTJEePN++/2i3BqlZfXz
A0Rj6/lvqZ3YguZFoiUA3bexbGjCLgzN8MyCSdrfvKER0Ea6Qn49liU7QWFG1/gd61ks7XzykPQ4
OCWObUzsSqQDdCWv5nQT3ifbLscpK2twTDstpjvs7gMlAgApoKUaTgyG1MgBM8U81jHh03tnR6tV
1n2fFXU4+0eAfw38P8dKMgTKwuciegi3TOPXrj5+s0DLvBlrwnPxNEG9BlhWFZOTjRMx4efjDN+V
cIRTyOAl6ExeHKlffV6RTztqM9J9wqeDLT7MDi/YfUsyhdAnvnSmqTIsg0sFdmpx7cd5WkIKsn1S
EKF1jB7VKJNBpZSkBQaMuUx7DVILdueXxE4qZP9cjPltVvLHv6dnztP+ip5SefDSeG/wIJ1BVyRQ
0EhHlzWFQsZVor2XCdH7/8stYu+Ec81DVjEVnLArwvcexH12WQ/MZGXw1/wYL4oO+eN12C7pPmLX
LS1BsGLCUFA9Fz9xDWm3VFz7N02qhSqGFvHqIF3/KiTd9SMAPCD8wEIGWSccksCBlIkyfJuXKh6Z
EGC90OQn+BHe869IOLauRY0g1S3wc86atMWUTXJKHq3wZ6xpIxeu9tg/b39mSueP0Z8GaGxljRte
qAYFwAa8MbR8qr7wP6VzDnWW9ShBonzqUci2oKEDTUgGUMIpHQw/wqS7Hgi+qK7LzTi2bj4SI90T
ua40VidRR6WxlJuht0qSCOhEhgRZ6L3CcQrKilebkrvlW+KiboFdL+wGXY39cdMpU7oMNqcb3QuU
BNkkj++eod+b+PesjMKMkmf8uci+mFCQK4DSXDKUgkaWVu/mMXBJHPDAXH7PZ6ya1DiAp5K9VMRv
zndr7d+LHTcXsQyFnXS6OcXYiMdZ57M0R5uSghUmaRaz84IBzqn4EFFuFt07i7AmnBPXxeDgdzJ7
MuNIFygSn/r16unKmFrYq7aYi70KqmgJNy3l7aX1W/Cx4q1ge9QlqAA55Ha2okimrFE0BRC1lFqP
nbbsGhGkMCCG4CH4HoeERJ72Rl4sbIM4HjOCiPXN8Y9t06kxFC//As4LhvC8OUVW4EchXqMCr3Ul
G9ViYqknTyRelT8qrbgOZlRSmuyDYkQH3eM+h8hml8V/zy6Yw22bvxTAxiNCO+LrKIjWEIaywT3y
Z8peWZ9u2qc/XRuVeArXfNGy7Y3N4mx4iNH+Dgqp9jbEg/JnQEKjElfWmg2RV4tOonN49NHj+CXF
ICaN5luPpx6nXZQ8OR2aVNwpJIAiFhMlzRju+By3II46HuJYKw+gfMYF0ScAHJKTaxOHtcjnI+82
3LbG65zDMH/SPdF2rq/D0b5fDa9E8OsAsFhLq/R4CJLIKsYaKs8YfGS9e2hq6VAlj4xhG4tszqIC
tRbaR9xw2uu/zS+siJ7RzM7sNnQCAyMZDXnX7sRx9b9lAOf71aqZc7nUsjapO9AGLKmSisR+CDQx
Q5iqy/7g0OFYONG7p8aR9WTjLrNAJmESqXZK59tOq6WNmxC7RSKD5KMpWSqu+nS9qlOT5jXD5yE9
gmOQ4QFhYk5vl65Sx5/oJhJhTBaRcwVdHnH3Ahu6zYbuQ1eGzsJ8zD+is0SimeC7UrVsVZFXWuo6
KiJQevLBNg/HS0fXZueXCssC+5MJhEKepn4dIiL52l+cfRysl2ikZchQCZjsISsehZB6nBOBcEsI
gyJL8Dh7fDR2dZU20UER1zPYlBw3013iWpcINugSCIbWzmB7Wmz6ZGxtb5ZlZAfmjlPDtUeDi8Ce
afVyRuhPZglVQEB9PZe7b04BYPP7MfNZrIjkZQXx2w9XZnC0U3PKTqbKkPGnf/tL3jUYHim0Y0s5
CNsqP66lde9AAPhN20awWExU+7dxblTNG3L/RpeXKDKxig4jEOWiz9LJ3PaoWdvYuNr7eOa2AwFq
R/Ms6odzDEYv6qzi1ldpx0yTm8zo2xpLUHZj9hlmacqEUI/H6qfzfkxgDNShPcSXjnU6B2/uEsg1
0rF77UgWYhOw4iqj13s/d/rz8q9XadKUGEbziwlXH1MakJr0nXfmNm50lbe+fp3okHWUqFut5riv
WTG19os2bs8GREUu8Pp97icYlOUc0cRRkmg5nEWwCiq2R9+MCes8mpHxytMzQYFIIZSUzcCd29Hg
2GSPlO1qzFmSMIz9ljBP7esxh67FbcC7kBVZon2vqipkpf63Jd4FEkXvLBO8eivLkA7GoDmfqoJr
QqNyQlTDAGI+VaK7oO003Wvx1uUFXiyzsnav3YhMC5OaSxKiqO4frjfih2PhsAJQff+LTCP1eNOA
aWWvCmeALJMdfLFrfipQ31vk+zEe1uPGi8XD0B2mqlmNszUIaKHDNHd9UkWCgu20mBdgJ1lS+S/5
bxEkXllUEFzeNdM33cBqCS9Sgd3lmSwog41q7ceT29EmGDSmEp+lfXr7SNcVN/CcFO5WkUjg4mPl
lfsrucJKV4CRqP2HJYhw1NvBXJ+Au2U0ilUVMgySGFrPePgYffHKUp8u6LRd6KW3piS6Bqi1BuoV
N1z6RnFuo99KdTe3itM0fu2xSyDRcjWjuH/0FHq3DPq61q/aunDiDUzDQ0cQcKQWUUHY0/AFciPV
gDUp1aP7Dexqgn5fyKoSumt6b1RPN3nG0oPq5ozduodGF7xTVqTZy7M2spy1//31FLsf1H7xzUDw
ptjN43P6EVgqj1eLWlqLqg08sk5HcchvXAgDrByfvGZ0IsWIFMKaCWXLK5bvWHnD1XAf/8YIw3rl
hje8pQo5CCjsj6Tgh9K6mISUR0TDZH7BfCk3AuqXydN+CttRoOw1mbXnhPW/4WhbF24RfvECO4uD
6LqrK9JEZjX4mm9xafziAe5iw9Lf0sfA4cwPAjWjJnIFHJUpcVuvNY8hH9bGxnMUcHAPemKwD6tg
yhV9TS/KSj7VdZFQ/RZmLWaEKphmIB0bKwH50Feljg6gaJ3g/+Jv+6faLsY1FtMjbJRRtFULGaob
PWVgrTBjuhCNMW6ELGXy6zMYb8pT/CNo4v+NISAo9aq4pvWwJFdn8ejEoyiU0typq5jc//T70bNu
R8Zcsb1EHmsr/LgIxkPXX6Qr8fg86+aNdTxHHoFoUK6fTN7GOFfEhyAZ5SxOtMfNOWzicSzN7vBC
sHhW7KARK9mD56Gnui7lW5yUv40agF7N1Cb/fF0ccZRSqyFs8RevpVQEOyQR2ERiWjJojiBmt0GR
UHFWBI9Kkvs+3cCAHc2sCh6I+ImV2Utdt3EUDc6/Sd9WxyhwvhG3YApgTaB2KCFGswU15lunCwLl
XUYWADut/QfnXlycKuBGjn7+lYyKUR/VNbSFZzRs5I0EFpuw7UJ8kgZOV+inddMuFJSlUkxg9A89
3NotaPk7Lk/wpDVblVBq79JC1NnoCUYDYAVkzFQUg9/F0BU0yxchSL+YHN5tFI4gR47UkexBsUoP
osYvRII51yCT50Vy1OIH/7fzSPwXuoVeSoAl2AjR/2bs1cS/HfCyLyM8hN5XCrmDPPdz9PEwY1wz
tclvtkaW6vCLUZLTRL2nCWY/QTKKFFs1A7gyXpk5GYeZeq0/kZ9FYBkPSHOP5exF3Y3vDgtyeGu0
HqQgWLVgWxH2wYkkc4mugoTtJ+uhNFmCbTtdbSJHdLneK1VkDtmdmsBZAMBq6cV6hwhW5uBpM+zp
DaCWIzPDlC5Mjo+girQx/991x4hRV/9PWPheSfXtprt3C8D0HErKmqPgcFJmB7b8oGiy3XQrd3KA
1Kzhm94nhoTkTzyOVRrlvLblf0TC4iGzTtvUaahPIOTC36JRr7gw6gHIj8at4JZnhvUnQDm6W/yn
bVC+RtBv8Dwewk4G9Xe3krmRFXHLH5stLIWs2kT9clcF2HExxasQl0y0t6TFbm+dx+0xoWvXN+p1
+D15Yqc3+4krO107RIr1ILuCju1YwIjzLsduupn3OT0VmrR5nQH5I8uAyz6VzK8nr2YvCuKY0G+P
AeBjoxj6O2ASzP9UeSuIo0uOv0R6HoVML/X/yhl6mq2kgu/AeWmrR9TVJZ44n0AAYMFVpTqiqmBW
cTIjj9nNF0JtEEFKWHe49q3uAPBBKvLrYo1wWu2mA2zlYpT9uqPXCSBWCGwNNbKBW/fHHd1mMcfS
qZu9QzLc6158thohPUbKX4tOJPrEc4MPFhi8lzfomphE4aJnNq6fHsDgY3fVmneDs+d3xGSDvJr2
wyPm8zFLY91R5V2utS/k2Nl9FGpOU4mENZsiaGIml8Gib83lL2pIVgqN4uW07SDjewtYw8EVWENH
yovo+IzQ5JuqqyjNmo/MJ6f7WVLPE251n3b8M3HK4Ulw8pZA5wVeJrYV51qHLT9ZwLSXMt7guLAs
qRFQBJj9KYqo8OrrX+lEKTSLjf0vqFg7tMpfzWbYM3qxD+SCZrTQQo5rgkwWIxs2cQFXlX6yWZJA
7O1StJIHABJl0JsG/K6z2cc3jLss1t98vMThk1qJ+sWfaaBozYx/G7V6glpkD7eZ+/3ntundtSHR
jmd5rxO+2R79SojZrjZh5VMUAWs3+ePEwkBqaXqnQXe5FZEPziw1h0yAGAo4vmBrFzfoVvEi7NCU
zOM0D0cbXMM/tM6ALna6aQ4MHC4OeNulK4+/FTrAc0DAc0i4DtFD0HXhLrxjPqKBaQb58QPoj3yo
jvob/XoubZ8BZoEwRHeFX19PPitmu3zIoftE/hu7+69cJOCyFDdrFHMirQ0+8ycfuzncPvcv/S5p
QjKKwuQ3Ec+pJqbjs8dtknoNUSe3ZwR5uk8lsO1pc6O9K1Xfhkb+SmFfyJZ8RSoL9RnRqO2x/zpu
XyE9Tsb7YvZIX6DZhtkKx6HHy2X1fMaJWb3mGI597MfDW9IA5P5utJSBpDhMIlLOi78jZm1Do7pb
pIGn+P+2CWvREpODuQwi+WgLwiwr5AvAWaG4q8U/D2Ao2KMh+0n0azAaDq+bQXcaxFL+2321phZ4
tiEP31az7xZLX8x/JSC+Nm3ofzIE41CCpRWeTCVUiFY7ZubelNLlQa7ZR2asRWrFbmF0tWaCRa2f
vmHVGGN5aYYx6DKAPdJkbPhJrn3QssoSLn5nZ45yTFYf2U0Fyz+V3zqm3gEZg5EeRt6YnWqJvFY4
E0wL2oPd6iBjDe5AYZ7zRG1umaSGGqYpZKgil8tgFijRG+U2wFUvd3iO6kfp4drp5XkW827MQNsm
bHt16kvs+4oN5Vtw19ht3oBlxRpl0AiHr3Eb6pD+shIIUgG1djv5ldsqjc8VfsqpNv4SYTF5ORbm
KcHkyvbc62cYMUr/1W2UXWS7iDoarMvJ6WLPU6hHBLMKsW9JsVE9jE447ehV4f+uR7GCLClFGjxH
TopkdRko3nxdDIhJIQPlHbZrKmX9y0g++fZn2hCg94IJy2HudDYE5TBJIjLWlSz4MMJzA3YHGITs
pMPhlrZ/vLmJ6mzPmEyPGEMyo9L5xNI39fzLFxZO1RcwWpHD6J//ITjpwrr4pYVdjMJs9lSR75UL
nKIzdm2j+fso4bJXwwPz3oSN9R3AKrSaqw6WNvO7PiPUBR142k+PCZ2ueDLxz2q8uJh0zLtdMj5z
VlhlcWG2MTOIQ5cdkagt7NEvGRcLHM00125qpscGg0KLoy98wy7isBhWPb1DMqcLXq2bmqoqLUIU
WS4hxrPEzjwF0HfATFoK9i2ngB1EsLKu9W8olULO12INlO3Nlc9YSIiBo2THgaf6+7IUVXMnRnfy
M3xJx+Rj8a0yweLb0tsGDBsSUn8G6GVE3ukFXmO6R9uuYkVhEjZuyRQSWy1UGXRCYSAD8Uxt4h8U
d1LIF6N7Qr/J2jH2v7mcFObe2A+pt/inca5yR1JgOQt4cMk3W8rPmF3rMSPjEGqHcMxTIivdjwQX
yozqaMY7CwePqCK/AAVtO9ochrVouz/sUFbu6BcLidyZPHkURX1uqQeF5bHbmEWr5sFk+EHwp9/d
OrJygr/wR9/xHaZO4dRWEoA2tTn9Ra9kFcCqC2a+LkElAaTbfVxq60xzZy4fR2D1dZHQJVlzR/7T
MMkQqCQBQHWSkXRF3Yrm3BJH5h+GRPrfUzkQTCPdSXWixIxamk9sBrC/B8roGF6PCV7RgKCFSV15
lG3iMGMNI40EgO0dl2OhY4R2EhGU8NxYBJ9NUiVYxyEeRhibPq67e/usUogjMpCy+LaRWYovbWIa
baaeyZ0A62v9ILNPhO0D7zQ/aBSJko+DTCuHlDHutyzhwTQ8aNK3xwWYEwhuaX0QNg0QJak5VdAM
xU9jpqsUKJ6JOhOB0BAvuspTy1WiZdW+0zfQksaddnsx6L3TIFdKO1jTuqHYKdhxTAkFzUzO3AV9
LdujwuU1tL0EJunQShGfzGiI+PAmyc5XB98eL7tGXzEjVcBrvOYYh0RbP4Mqrp9u5jpaHej+7Q3w
a9NKlierH4pPCeiUMai+FyhSs1AMk95sM5XbYw2PETWmjldRfeI/6yY975LPXfKAcDZIz8tAsNDN
EKngc0jKgOTz2/CXRMGT3GfKG9UnYuHLu1Nc8aNYbV4yImWFzYD/TqA+FkBgWRStnJRFdE+U3QuH
B+Xy9T6XqUfk80o1oGnV6mmGdeNCtFxYQbkfg589rADtBgYcq11++txtKS5iwGRYwOSGl0TeSFr8
dHmoB/dYB+aeeuIi9cVbZFdZAN4m6jDub2tmoMidolr305X8GzhIRAcfuqg+nJh/p5/TKBqjFwZ3
BQXgrNgs8FLslsSy/yL4Fsl4KyMQgtQReNPemvRXlRjAxoiqTsV0p9KH7XjItmx+HpP6x1TmUcpG
jSPNWF3BMUgL3LrCwtFeyWPbOMhQy9Yz07Z1RlYHXBFRpSaoQW7rfeYn/g9t8/dOkck1jdhnB2wN
SOrLfcu/ZXuUfUeQ9dGuSV/YL284+jruV+nxiWxcx04li+WUeuCRkfAG2kCQ3D3RY+IS4NHK3b/P
miFaF4ZVOrF+ASSmvksZD8qnOC3q+mJ/4YMQ7iel9SOoWKFXPn5M1qYBmWUl50+6TxEK49BJgjH5
AAmle2RVy8YrJNVzofQevSo23S1yfaBDjhVvpjz5YvGKyzQrFYsF4fzkRzxEJGAa+btEgnHHbck0
wIpFDpqC40wxaQGRWtESvqRsLPd3bEA/4U9gPzGOnCgVdCauFR9G2oK2Q2ixHJ+zhESghu4duQic
kGiunsatwWpBW8ApDwfM4+PKaZhUs8IX5k7zcsxaNUU0lG+Bl/n0/fzQ0B26S92YYKhWfHfmJ/e7
d1DnWRWJfghDF7T7toWXElaq2QWbNgUVhlvdS6en56JqvOFjV6oimFAH5Sz9bxyHyCi0hippRmdK
cqFxa13K5D2LfENtas+UltwKFc9Nf9bHCAJyuIAcYFkbJu8kOyxx5y3bwxEKAGfVdRFHw2kEDAsO
+9lJZ7pPc4RoTKflovPT9YdgffmNEOflcB/LOUmr4/dH1T/7hLm/vPA+mwsP8Fn8DgxJk97iNcBT
762Nc8ZPbrgdyN0rrwYfpThp/75AxKKpz7iLe8Wv5F80xdUFCsrFg1qAEPnXPjF7Y0n8EFcBP5Xn
RPVw28ePvTVKUso9UuCbqdJUnE5ywVqP6dUykIoP5Du6uHa4bcA2U3rHt5Jks5LajPw5kPQRb5ZF
wXG24GNqUu2cf8dOxGBAyPx94qhk2OzVOBNbJQh0/slomj8MOzdKWpN5k2O2VPlq1PVO9DY8eg1t
NDTHkDwhyB67gM8/VkCxmlMWWVWXuL902m5L6uEJ1SxkB2mvu/LV58pPcOKan/3cGBtkE9RdJo+5
vn5flJyBK6O1BpwnPCSW4gR2hQgKi3/PLhpTHBLVbLxxhSpOwNOVY1YbiGNyRq4BAc/UxRhnpzk/
hxUZJ14dnlCoz7shvsNGnTTC8Hfxtl0m6YyQ4zW3H4UHRDixm5UCLGfxmIT5Gb9lUfUp2KvKZ+ZL
XyP94KbQ2PKoiIAenJ1BvrziX94kuttkF+JE7gv7GPc0GDmpTQZqEBYP5HiGqY6RYEtbHbd1CEDA
9z/6+jQeMnRmKqcTRTzt+4ONzk01JZ1JzMyC+xI75QycnocMLPoO3UIenoZpPqsIYk/DeDeMkjPt
9Z47RquqH7OmW13tYnkcxGoihx6zpQi8m12swtuFs9Ahz6ZpluVVkinT9BQQ1ixhYCvZRVv8vEgw
m4VYkHLgIcQtHVBImvWmJPyxMYLM81hvFzX26nvr9WARnPwABu8UOvn7an7nD6Hn70ScWEl4sQIF
7dgm11MKGQB0E3SjnJBor9a3RMCBHuF+v4ejyqX0CeUTLNre+yrotTzXxRU53S2NAHp40dZfdDzB
KlGQEvDqgwETbVo6ZYqAPH43WrY7lh8WmN/7w5+/AYXKfF/PmpAHE8PZr715aoSdrVp70PZQ+91Q
YJzz7ZxGGfdphY0ZjZcC2ysu973qJNcsFP6fn6KFvG71M82Q8L3zfCswBSNjXvZNLumoyzE1I23e
iuQ7un39aqgPje4PaCHDLN6t014sda/f9cyz90msEAtcnNiVm+YGeUBgY/X7vlnn2DVdpxYPXWXz
e65CsjkU+YMFqVTb0R61tHceVaz8bS3b70qbsAYx6Ldghe1SLNvi40ZEJU9bqUQlRTusfSRJnw7E
SvtSPuni0ozpXz8aINrIlYtponorXAPeE4l7bLASd+7KvZLaXk2v0ccZ+6wxZHoLxR4lUgN/Ogcf
0lrWAJGXJglNK2WWc3qyr+DOVRgkwQfMa/1HnXUTowpInkA+zcUwHR8MZK9e4Sp7M8WwPb2lbVxX
n+FzODPazEetCyJW3UzhVtSWOTc7SKCLN4xYMrF9R2dtUsoBZJTlTB4O/bNR0V9wJk4daMOxhqWq
28ZVRBA82t0T63VHu7AxPShAUJVtaE12SmqlwDxnh+eyMD/A9u3sDchwLmEtijyZwGQiBxiThkRB
7bcH2EqOKTzqMLv32+OtlT5nuOiOdb+d05zr9TPcK3xyoFYTLYKcSi0gs7D8QANQefeXYG7ps/JR
7t5NDGcByYgFzcxd5+GctVr17oHIqYRVEIrsn94IMwKVWcAC4ifqLMOjHIGEKYM4Tk6QxT6jEze9
bBU/R3Vi/Nz0llWOWLxFuUO3qfhsMQjuKinAq5D5kfHOr1FEaYM55VVwIHW8eKPG7zwcm94W2bKh
ar8nMJIeWV7XrW5W+IPiwPbQnRVWMykgBbE2sa3KxKJvDSb+CjDvDKBTQlkRWK9im+Y+5ZiTU7s/
JhFUNsmHNJNpK323rT3WovZwtGYLIyJ0YlzYeAhx9KoChM5qyDwGwFXcxUH9WfS+gzXou34quTHb
yAeEUJSjw2E8AXGbR59QLXQjkIEPn5OmkXo+vWTDHHJmBfpFzLQheUHSNgw/CjDVD0rdgVd46Obl
R3K1VK9UG1Tba3FdzNdfz1Q5zX6jGlf7oPDSbWouILgMPLl+uNDwzSdVZvg2XeMR02WPRmZWIeIo
yB/wFeld2blkpCju8mpbsq6Arr8dGwb1PfHTzHn3L/bv2Uw+vigmiEBBA37E+xlNX1+ipKuk5nhB
IB9Mlxld8Z7+ikv177fAtWlt6T9NG0SIYIxoIqwS9fL7iZQNmbjPQzSiUNxq2DB4Hu9d4HkbVbHU
nRdKbsEPiFcAmrGGxS88/Bdic47+F0Xz9FOpfHuQ5biBI/r/AGb6XYHyZFifQ+MM+6SvzfC1dffV
jKYgBKJ/3+PP2+X/+JPTJGSsRzOAAxhue4NYXLDvN3DhX7UDW7lIoD++4vP+h8Wwg06S6DJ1qT+Q
DLHPUAO/2ZfdC2J+xeX96fZw9zyiPYA+yoFwjRsPg0rmOkYrzKczkJerY+nDIF8izNkrRwREignS
FCdreZZqgYSM6IhlfmHfDyuA0Mrouvd3SxriJVPFR/S2e/Rs48SIl0isBfnmWC6nGVzTexP1rw1A
FLhSOFzDL1sDDv/80+q0D/fMrGdDkQLs3Suo6JF7oWEij+zYhH7yvLMKhilM0I8wtkiNbx/DxMp+
74VEVGEJqVHkh1X6rWiCwLKa94rFKQki2K0I0lSMVBxD2zcXZ+fqH0T9bXB1WQjzEZkNEVfJ9Rso
0IYxNpRedvcQn6sZ6r0qkBDkV2YqbnntTzGxHRbS4KvYTSWBAqhEPpavFsHGavB5l/W1zz4cKliP
WIIO+UbGHfRcDQuLV3eWGZbRXg6QjY6R392eOrtkEGeYIzm86mUmqDSUX870tGao1GbeYVGIiPks
a7xxizpAouKDCdQFYIGl/s1lrxVgHHKxbOlyQDgkKl4O9rhsm8wDSGT52/hXVAI69T/pfBeWxKNN
haCPFAgBzV2TU7jC3omIBDu1bKJYIMd/yP75pBFnQaC0bhxHsVBu+xyr8KN6kWKKSNvRAiZyLN8A
KzqQ/MruER7er2mN1vgL9j5aYEH0XxvzaaIHkXyv+LnhfXB669IPPYFvRPD2UZYrGZr6zSRR7F5X
vjNZ9EYiOTCgxL7t41Hwa2aT79JIN4A5yh+uzt4KjDq1ie4TTiM2S2lGVFOaWA5+isxsNsjX3AQr
KHLfe0wYm75t6aEWfDHq1zioIU/+q2qc+qjTRW1zxyFvbN8idAafmWlhi3/kRY61pZTrJtSKFu1h
/mXX5KL3m1VqyGCQuXDEmm2AfhFUHSdUeqya9usyKpisBYrbTAvdQQtJZ+mk3JYJAHYNA7MINk8X
39UuFAiX+xrybPsd8xTuOUy9FQiKmacXf75eHpFSKV/zvIsJ1gganROv+uVZIWQ18mvsuYmc2iLX
tLh7DnWyU9i80SU2/qPqp8+ZnAmCVyQH+77HC+8REi+TReE3xgBEd7UMKbvhBLqGHTYMAiEXsCKr
Ox+fDTN6j2yusHlukZfYjWYf+jttJk5DccEJUHX22VE8N8skPoNs8V5I6L7+h728GTsWC6IkPzKa
071ijdlNJsrkEuNq8RntjHJr2+P8mlyNn4xCzDk3fDsWpvoOp/i+r8c4fVbDbYphkihQTFHJ0UxA
9/outpAkFl+AbEgkjh4bywdLFTWm/0w1CRgK4dbOrcoNU4TK3BlSA987fuuIUbdysy5u14It8nd5
jH3yC7rOYRQUqphE6JqyF9DzIg2yTFvgkjA+gjO6jSzqKsVEOAUrNWJtF1Or1pFXU76INZfyP5Pk
6wXWehtgYKiDIv3WA7lnZzlkUKJr4vsEnm0Gl/+wSHMJhK0MsiR5WX6QpSOF70lFc2LgxaZMu0Gu
OYXxfFC+GuccrY8Wgf0C+UUWUTdKaz5WU21NTbXMnnrRQsYgIwCI0SUnsRaQa052xflmGshMhnuo
KVpTv9y6jOAjmdQogO0MY0FFlFdXZM43mQc0IScBB/BeN8vMMezQNmetZEe8vUM7VwmIqZDxX5CE
qBqdV6pPEvwSUhzbChkuX23jH2YYeTzQQhwixOuHibKjboK/J24mr+EEZGIbbBsQS6GhkzZ2mH+y
v8htr+bl03SuSqn/elJlfdVkFSgtuASgJnGxcQbsi/RY1jrLVsBKRvZ5Awp0xVhx1YKNOWhF0+zI
5y3feCkI2iQFaZf93xWUaUbEG25UW+u2e5X7PKZoxflBpkJT5HQE9a0V604KLgwFLqC90dsgQwbT
0HWVLF09kr51OLYTX95rRhP0BuXrltTP/dmOjBJSkgZ0g1bgis5dIC095Q1E4oR+iRJ+00tu/gIA
UdfJ24NIDtYgM0PrDcY4fOyFOBtRtQ+EaEUhW32I8Fo+1LUyF19AjNImM2tePMX3RzgO0qGmdbV/
4mWFQU3I9vL2nnY9IMxhYRlOt0/zpGICbW0Tq8vCucrHnH/swR5vWblQhEcdNBaMzgwOmZAl8x2R
Ggi4A7UG/7QsDFuATDcfEl/2SIhXBgmRbTlx7pWLQSVEdIpsWgwqArimCOMDBQzrimDjmr26uxtk
kj6N56LHiC7OU9Fqoo99VSJ8QZ1WEXcGK0AoXf9v093mcaXSVlqhTMepHV5yP6KdIy0rcz886we8
b/1x4p8ZiVW1XgBv3TZgU6HpQVlck/hTJEa5h5uDSUT804SZeKk0w1/RLX2f3y4rHiCBCQE6UCRP
r0pGOsCuHZlaeT5WN92199XjqrxEnK661MYs60exf+hgU1AxReRg0bJ9KPKr+wwe//shhVu218il
wcExWGhm3OlMekFjvSrmaudX0yMh51Z9F9E8ohiJfZNJROBbHl4yauTZgsDWsOHMOWk1rtovMkCC
GP+2JmldA0Fh4GDMfs+OMKTDjYZs7/WL9iKpfARCYPIpno5AHUSVEwjsZOgi/KGXoJZO8m3t0Okd
uvHlrWDR4KDicnP59JWYhTTtTaryuNPTqxS2bh0InlSxgAj1g73gr7QbStsg0g7qkTmvchAVoMwa
UURjdEm+w5Txue65Ml+LSm7D4v6/r2TaNPY+xUibCN2JmQkr2Co59CzATDfF43yztDOx9iymyD4v
WmMgB2J9RrylZOMBKf41H4YBDCGJvSfteN92SzkNwDsObLPm3vfAHg2yOYrDtqKfKX7HKwpVSBvU
rvp0CjsXE1QMlw6pvTqBpDBQHKoygqb3eNwfaGnQ3+8PoCNc4VAdBL0xeTd5YC3mne2g5jUaS72e
6HilPVFHZX/ZbiRCSv1ASzw1cdd5Jp9g1tKIdqBEsA1V9ePgrMtR1y69NOJ8uQGoP2jXrz7BTE6S
18/yXkFZ1PmiNI+osR22ifBAPioAYaxfDO1hjq7NewuVcYiJfjuKtkvFMv29TEWV7yRHTMQnjqj7
jn6I26rJsQkc4fgXDgjYVnf07DowI49odUyWrAkF0LOb7z4Yvjf3Gb2bJPIA/vsmHTV1ZVSMNP9R
+7Zvbgq5J8EA/KKWdNe9+IK4znP+Nro/DW3iaH7bWqIoCbWPa25AcuPPZu3RV2asHL5iJPEB6sbk
90GOFFr9Sq7nstPzE9qBlnp9hxbQNsbdKGoHvLq+YXl2/2ROneIelsGzutJCyCPQSBBso2jC994m
i+eO6wj61wF+CFPSGI4dewkGuspXGWHmFJy80RJIIQ4+tYvyC+qsDEiW5bszoMpW1OzawJqmbC31
/jLN5I5Xn+8qz6zLzKKS4tgB11nAnjg1kmGSurDxXf49sGWfUlc/vSlf7FuK9zDNT2SirEkpkDbi
KfBak1DnESea6hCfp0I/fcVmU97LuDnREJqloA0ncwcDtq8M4BNnn+4/A1yYM6hFDJRVk9efKcsE
pmJ34UKvoIVWpOpzxKbJIbWrJhdJLPedHa3WSHm7WuL0Epe4PMRmaZ0RjRXuGzHHMf60ykep/jTR
/H2PrLdesd0MRuDQ5JIi/RRUyVzkAtf/J5Qt70VkSo4k//l1X7/30n8Q0VWo5EMPzDXl0+kQ6eoU
dKXGZ6nfb0OJ21sxCgEqXLKkVQ5cT5a1i1RjxowWcgOKK2SKdTiqOeFFCyjq9+KBd8fOGYZmVOE7
RmgkdByFplMnfUGhyRSPaD2KmeynsW5tz2QSpHxSJN+B2TrW9dFei/S9mGB1A45yoiWcMysXBghp
Z5J2kAXfoaU/PkkgRiq+g5Tux7n+AYV6FAmyXxhKh49cjt+hnVhfrbuTFnRJ9W5o8HNzY1PN3wnN
Tj/ecFYjAZh+OPCJ0AZwMcKVT+YJEVzADNwPCC63dohKVRLX7f032/DJm6xw2xksQOYb1umI3dZl
yHdJEXTNAtA8xrH9y+3toRFfT07UCSzL09CweA0/MeYt5T3AI26peqXb6j2V3VzgemGTjpNgoOsn
YYxrXaQH6l2QnWkIMRCkMgccr7fKQR4ouLQ0ajgiNj9YVInw2fy1Glg7o1VKBHN0VRgkkLmJ9QzP
fTFiEoZFKyPyK0+mZn5ybT73Y0rvEDzg+hbTX9Y/K36S5L2wnI9LwgQDx79dxq6c0BYJpKVC3VMV
n+RJoP+xBH0Dw9OTnlj0/MC2yzGPq4un7nW7oKT5xPyVasNkQFiW+yqwxTZcx84dTgNghwSaWjKT
SCCV9rP60lLHfASO480zhKzDkHq0w9gl60KuTrmq2sHkqkw1nD8gFhzYbNA7odH5zYtGFhgBfTsq
Wu82oGGFDKSCDpwLrBqae1pViEdlp85fRT8uA2FvZeFZp/7pv2L0RZl5E8dMzqAol48Jz41DCbz9
5jxzv3uyb6ZEYUZwaSQoyq0B5ygZyWCqfPyIJHPn+uh7iDgTX6J9N7eha5KHKkgnsgX+kxXXxI6k
xPXOvG6USfEUcC3DBxf4A/GUfZUpsASo8TYjzLnrgp/qX6Y+PH3dDtmrAbImq3DtOv8b2yWKeohM
X2zNBzbDDAId65V8PJ1TwpsYOHy4bh6eYOAIyHm0kRl0ZELhIWRlCmIzcaYGFSzibwxomHtuqR3A
ygvRFR3We4DYbg07lCbvnhojlXXVLmEX90kKTBbuP3wnyz1XKvPq79TqkkDCpQ8QrljjSfJfN0wx
4sXYAnpLWoqjVaR5OLCJWSV15QoKRJYeQxvHn/c4D5h/Y7K+np8KT7F6h0OpccbY/L+nimlu4N3a
EkjcKa0qCXncx6W8o5WrqvBQmI5GYB3raToPTFG2Pc0FIEMfWH4WV9kIr3DNm29RNhOT+duvl5sQ
ozkUYwohVr0zR+z79xO8FYGOj/Vimpt/fMi60ZOowjWtvhZydH7dvAgvAdfAZ8KS7YhhxGn7rIkI
f9HdJxvYuYomtLPihVxq0/h0Bhkm4ar7iqP6NoDGmYlrFMYlQATz9j517rFp8vwgVEvUW8OReOyK
E0zBtRI5/X8+1RMX3X5ljvIxmelI55enQN1CTwg9vMkm1WL9DE6zpsSmnpZY9Qu2hr+u4zqUgeIU
uTv1164joSN4sccxKFgPf81zaS5tfUj4EvSTcEyuHVgPdhaeOYr7GbZ7uRB4fGcwqrkTqU+tFn/7
SzSLMvPNIJ+hOo1/BRMnyeyYJWbkBzIx/Z8JTIS4CepW+bzzylQgnQxKYFMp34lDCLxYb1Vx8EtT
BkSqf/l06M5m4eTaO0GDZ9mkyNlLCYUky6NCE/O44y2ei4635jKzjpD4J7H6FSsJF0oSCDJLoNPk
vXYrdwfsIM5ir6wQLHYq9qGxppncVIUKYBi3fMkP7hkF1s6kOPa14s0qvcaNr7ikfc+aHOvqakHb
/NvzaO2BIKEynRCLVl9Ea9MGHv7PM+yuXyJ8kbpr3kSAoTz6zM9yqm6vHEODkDizrF96dd5wwp1a
L54HxDl5W60qV2MNwsed0eLla0F3JOrKP4SfwkavXCyTq68Ot5u5tnWuArA2yE2Z/GLJJ0gj/lx1
93X7To2MpsuDgi6st67WkGz/Sw28mEQv6hHW7ldCllwXST+lgWD3IheCFxBLU9zpwDXf2936N0n1
xmnk+ME1gg5yYKYJhsytS4/eFgLKtM1p8Ujbs9945AW4YTQt4MffsNJeJmqcwCktuLxfm1Y0+S/6
ERYf+MaR6NFjDtnxuXKnmPXVuktXTw4oB/1OXYF3gemuDze4PsV35hmlQbHBfg8fhT5cYwsz0iUn
wIeyV/VF3Q6VWxzlMViiESS9yGEMcns1dhYf19B11V2t1tJFIrhTHOxObSKPO5yVNGSSv72sFTMp
TRr+3F8uAN5gqoO/xqMK7pugICHcT7wJL3nQp3U7R4fYpakRLto6J8u0wZTpjEwwzdSneAveAfHf
xHBT4qkhbHrAqi4Om8PrPiD+jIBFMH6N4JTHFnghO7PuXBxEKW7UJ0rS+9/QbageeZa925gXz2i3
b0H6mR2KbNS1epa4vr5GzTAoc0n2zyq0ti3pEN9VIYrqbvthqYFayb3ZABJ7/n+Adl9XBIko14+4
K4f7LdxrHLx+4lNQ65ZcUHPlG2uwCAMPAUOiFwkqsj54XlKISvJiTJAanxXd8b8PMz3UCE4Uuj5k
U/q6Cp5850ocfm51WnQrn+d3A1QtkJrHOHgQ89kpUg6rBCDzSjpvdYuLdJbLAmNHM/J2ISnmVFfn
Be/XmfgSrUqsQ1wlx6f+0xcrXg/YqKrHcjGIoi+ifyXduXTZMqFQ9YJlvJvXnDSgZbV2Z6lji4Dw
1KxxrZLLiy+W4V7PYcVRDXlWssgFCiLRD8+R2mYG0BL/Zr+pgMCUCvQU9XkEUg++0OcOXFNVrh+d
HEXKDZjs9cBP/1RnnrGYF7uMqQUuwn6YXuBXGkED3zaPN2RBpYra6u5Ugr3N2UDZtr3oo7cSxLio
WxkF/wa5kzc9vz2PK0aInMeBIskod3hB/askoQgadDS8ftm8nm7PYSjqC6wcyS8DV4aXBDu8dVZP
Q2l9pjitlEugRHt6+/htqn32Sj/VHoEFSV1381WWUbfuqv5CQJVDy3Gn6KcSoQYRvqkCmIIL6sf0
N0jFCx+UgIXx4sZC0WADMyOmLW8tdnS6ELZMX9HePOiy/ZgE5uQAWEWLXwUHGtvuLhdW84XNytXs
F/bT/bTUDsVv6pfjUfpaTqpyJkO23O0sNEs9Qny2cJ+K/1n6E8K7NcKI9bs6hOEMa8t82ErA2EML
1ALkARiwrYuuF1DTEOpFk1mF3UQQc0GBhH6GrCnCKV/ZPbpTp1SJvGynfyYKw7Q/sgwoFU8N0ZJv
0bhgh1omz15lF0R54t5vZgud2CauBrshDtXFAOaSkWRQq99ojpZXbNHOe5dMhDyUxxuBuzQf1H4v
47TmG7MucWKbo6alf5ucqHCRmQyDTFQ0QlB2NlDEEXUZOV/bOwPCxan31eIOIHAwq1FzYf72S4wq
NIYOl1unQTVe4MrcKMze+ZXh0OqNrkQEOpn527HiTmTeVp9I6Ak58UEoJAE4qDuwL23945ts6tNw
On2EfqLsiHFmbUrgJ+VffuNbkDpU+5T8NYVN1QfYEDVHLdt5h1tGx6RG3HyIxHyeY/WzzrWEuV+M
eaLI+RSGD9XpPzfnnd4CZ6vkzkbJtp1TrImAvmSZDDp350cULHTWg0JHfUy48+6etWjBfFyM7X1g
P8jjtlmzlt24NTI1XNRfNHDlk/dqF6L6ljXcGkE8QI/ntt5jrM2y74EH87hM7oWrWFSx55DPnCzz
aN8NWM9hkFUff7vEAjfGxRqh2DWSBjf5EQ4l/B+Hlm4tttnuxZCjFfzyKwdIA0zR2W1TuY8nchLV
gBOgW5qutHeew6DewBAXvPClpBPEkftpTY434OlFdMEXuyhn7nBzZuJjlKJNHM0HIAVek/NsH7Mi
/HB4dIlKKdc0G1uhj7+KLXFzyso9UzcY6tv/eFY8CLWRyD+ML4ZrbG6jNlYWv2HQe94fnFub89rE
xuqrlg24MQidXctKXlTSu5QrSgJBCZ29lXLJ1aKM2sfSAPz6/A8UyoCPxOKV5woAsXMR2jNZnxBj
vZg2ue9NbACMAPXoQYGUdOAFakoUpdNVqOogrzq5vLa6or9TpA6UDUKOYgajvYltRv4jf4W1G3LX
0m8mDtG50Br2CgSQ0YWNdlrxr5NYtADOpq7K9PMJy9CPwjJKD5qOzt/Ccj7q+6B1yZ8JdMDdGLWm
saTzs5/MItwbc2vpoHrFqwwjVysXRcgKRHI6tYWya30hqVSStIdCnkTes8vtfTx4Az8GgD1AQaa7
f7BdP2zyE1KjoZULcO3XSZElG5FuefFf2DUCpLKIwL1cHEfuz3YKT44TdH4YaPfiY4GicfVAncn/
xysMG+i2uAIsIQocEZiFFIOxr/2hs62Ex+/Nujo0G+cv/xgv0mUbtHFuSnN6kRJLMt9lYJzvA7LA
Z+VSALobGneUcudnVVz6rsqHgQJZiZCIprrwKU0xfbE8efcla2Gk/Wv/qleN7hxe445OX6aRqAxK
rdSzUBPilhsQ3ah6K9kJFKGPEJzGJZiCjI8NSunwwaaaaGf/FmBouMDzj0s5C7vbfuWCHeFp1DTf
2+YtTTIAfaugx/GX0rXeFDr+ZawmVoFLBuro2Q2nqDAS9eyHyqrbS/ne7HqptkxM65/c4luxoZGD
m++Fuwy1h32rx0IdvjNskLgD3wJl0zQRI7L1xWqr9Ws1w8RxdlM1ppv6M8z7ApuQ1HP0CQ0xNmlA
2IS/2h2srQguFZvTdQzFGxH9e1sxEK+4CEnJQMMvUxhfG05XjB8DMSvgfVFkfIfGtWgaRamZGMwo
Zil7OnGA7y4guzwbO3348RYo29qVCucUaWFdyk6QTMhjpybadxYXh8otyopyfHYCRyaPOx9qAoj4
FqVzxqoesMb6WjIuTkXn0g0qxWyCJkUV1lz4ScsYXcGBvjyvr+RRGCZsQ8bTC5gGnvAI8eVAnOaL
fQzyQcfLB9tcTmc5Hg6MK1UM7H7QlJAeWz8BUcPvFAOwuwqqrfXM18xl9cGfUBItfRpXeQbPCYkx
4/wd4Uu5uQLj1JKmhnSEznVIQl/7IO68Ny3LYFXKC1MCMuqMf0hST1sv1KpaHlxxIvB9vSNi35Ic
XX1WMUShn4emWSB7DOwOa8itJLuqpvPA7ThrK66N8sJWIV3iZzM+BuCkJEUK1mBrfKr2A/yuxYxu
Zw8hbrsmbkd6p8rMI2rj8UtMGaUa8xfw+IxS544nNuCaqU+f3Upzjrl6nCfZKw8HTPYb04o+nJbY
JslEHAntjzhP5+XThUSLg9StGKXihaz8NflcKxjZ4cBxCoRhu29+Q29Odn13P5aAY7wTByNLRcMX
77ykLG5riO2qbpir4ENKF4kuZhRyFRgz/9Sn474bz8mn0x7yPoeO0V6cuwamw8o608qlQFfAwlol
CYK4G1KASDhSODuTUhs2qRYR+LZJ4dlc7f2lh0cXDlw7/GTf1lsJFg/bS1d1yjPgWdSPMyx1wslo
sVKYFSxNmsualzWXCUR/R4fK8zZk5dZtTGbv1ILAl++o2S7h1zFlhsLDaEx6FZhmp80BMgHLx8/H
AgdHPwxPR4lS59ZaCX1Cz/fxhBeukNu53GwOrmb/ZPzb/bX1qt4o4adDQaMsGBHCFGBYCV1TZTZU
jscL99klwRN1mT+mf+Zd/BcCCRwNGVu/uXJzGoU6UmP/mw2aq4cwcxqUrtHrjEhqSXF9oMA83MoG
qRJ3l3+cV+RF3hvdjpTOy0jdylUyGE7Nbx/Da/1Go6d2majLfTbX3cVXi/AaiIjiR2tFuK81YPfo
CIuGb9mkHct0mz8ey1nokW5iH6MuM0lRSj/zTH+XdENuOmSrLNBSni580peIcY6E3jg7Ib+ywz3/
R1PFZqHAi4gEPaliYZSs7Ws9kHAugxs/n1VUHrQ6E/w4P9d8AVkQzM+Gapd4+IOzaxm7doDsc2aZ
ytsk5/uLlU2doffhUxHnlO+Y8iqakEuIsIB36THfq+TZa3//T5w/QBh2wURYnd4K3TxQK7yBeYXb
qf7S7sITgZEQyrKy107LsUhsxM8eksQI3w9OUZc6zeC3QNgWobrMzdjnxfjODB7A4iQXKj6Ssi/S
NMRELATZlwUcRTcRPayHCW0cgpzqc52jM+65uxLLwLOBT+z3n+7ffqBxjOD9A1wZQ3VukQHvl0sF
0bml/4erCivjiTMXsqDljYthMRQWBBt8/rSZLAVmchFmYSnA0iXsZsuhTRdgHmeqvgLxOevf3afk
wDW4KKL37cZnA4/F7qAPc16dyn5nvEHt0lASf26g3Ei2EtQuBGwQ//wxNbYXnWr8XOL+my6K5PRS
+JGiOl0IijyRKY1QHoQ/GxRxQ1n9q4anHUU+itrhtRAb+ftkA+ADlMTtQ07AiejA8GKpm8+ZJBx3
TNYRavL7XxwhYYmcwUc/KzLE92qIL9au47Mf79nhm7ccGnYmfD1mKJWC25m5FBksVDek2Qf6rttz
b2nkeR+nBcdX7VSfzAZzY0uWY65MjYLrXfAMUzA2I7J8379KR7AYLcANoa8kIEeAz3Wq4H+dgh7I
1myVD7Fv2GSSqP2AXPDYok+T693onFFa+Dz+fe7WP/tlNG5oeGOrTJNVXnAYlxY9dPebNReJXDAr
tJZKMicJ+LQPclSwipP0Gtr5xbMNrBx5IKnMCaaOx49BUxUVwZXJMQoaYo3j8chipXa+xeZ0xaFQ
uVbJXg9phx0RLrnsmG/I2u0Wogr6NgV0YvTEjeBTkpem0za+U2OMnXUJLWk3WC5QfJTG0hvyB+wz
phXANzm5ftEgQ5mnA2Lb09yqOJRrSvrCBLUsJ4RPotyQbkBTV4IYmMRBVhlqFRyhJItqiwRG1T4a
oNjc1/FR8IRvSAYkpZnN0V/CUm/Ff395c+h1VAK63ppwytCHZdzFEtqRozwLijhcPNMtItfMz8Iz
pmUhE1kOL2iAPioJOb3th8Qtn+KpVyJrL4kcvw2k3bkUvUgxQHxt/V8UaN6C+DkAQ/5tCFkRswBp
GewMHWmJ6TqPgQJh7lxlkwJjvK5Xu7wq3D9I6ey80QvMrciXcnHkwr6DI4TCwP/T0zy5FOHi4AIk
6xNA9q8Iy3wTfr1K92NiqCBo17RT0wPlARHZAGeflsmWOVHlcPjjfj/MSItGb5y6lyufANdRRjtU
VM740SzdjNugPJYv33giRVjzE+YR2Bm9mhpsGxQaiAkDN0AOhovMSRCc6CP2AMnMLjyGAa2n7A63
ua8BlrcfVzXbg83JO19i4S64HS7ri9A5A5a9MGEN0rm2adluAx0Ew+oHslGzIQEVxtNogS/+P0NH
RxmIq8TKdSfkqGVT3tERRBB2hVWPgIkp30rx6g5JSiKWVz5eCu12qQFztL5jx8VLmML13NwtznDj
IOmmQOFAund/U+qcMTEdeu5ypbgubnhw63JsSM3s77uDwBzY5pKUgn8+InxdA1F8Vb93g9+u7Pkw
8EbYOgL3NeRE61BfA84dGsO0Do93AORD+2HztgH+gXj43exIf3LCPWwudnmF1w6pz5zL4byu1Whh
DPALlV8yKAqwr3t1eFDBP+cO+92EZoAZTvxpTXP6DCuBN3pj8GCCePxDGGiosf2QciK3lo4B7Duq
8WyWb0NAg2mDlqK0cFyqq0RpqczhpuY8SF591pCnpifDsYSaIjzW7E/rHEwdvU1xVOqwSA1HcSNZ
0VXtDB7j6c0Nxsf+K5lQVOWFe3RJzFahDu45RPmmPNyR8tSRwV87BVuOyPU3CvvuV5twdiCfn5wZ
Q3fcOGjOSHql/E+hKjNIXfYQNjlSIdnrs8nsqd5l/HsDP3OXegXOWUkOQDxH8uBbSq/DZs2X9teA
Zj34aTo43mg0vlTcUpyf0taQhmTaikHVCks8dH+24Z5edbtClz1m5hVQn7xxW1ztIiXOkcr5NwdV
viAqNZsFaTYDqBv5nYB+KkGPqeBdOdek1OscUXHcHsjTUGqdMN2cqYZMPoHcM+b8IzEB8X7P8Wja
FgZknRveeLZeF7lgPAT7hIVa5/i8X+LDms1zfXmnE2FXGPhc6J5PXi/pXiEgpJ9J8eoH8QX9BkCw
IBQG9sOq06Qrn4wVKlsOELujSTBXffN3IeLadHyCB0pIor6St+zfzder6rQuCM/i/jh2bHwpiwxR
rgMoEVu/o2obpPQwPDHcFjXKNsZ4opmI7rb7lfRGwRYKdlWCv/MLROb2urP12e/v2LzwwCte8+n0
5CWnOO/BpGl6GF14pFg/C7dIkXj23AyPTtLoEPwHJCDJ72H0ZGVCBmqSZXeB45upYYGfrOhLw+1N
7uAXvWvRT95spBE+tCLh8mY8Cdi3lvavRIlkDOFZuwkAbXaL36x8C/y3zXS4qgAF7557SIRPpUvG
Ejt9+/D4LLQS/PzM+Ec6gnDq3XyUHZzxv8BXGiHrB4RY9fu1pbuw5d/H8eXM3pszn4J7Cm2yRtjr
M18k9HKVdxyOthlm6etCA1ujUQ3za5e+vcqZpO+0x3SnsQihsXtRJzuzBbsSCLVpVbP1jkKQFFsN
44CNyWvDg+qhJ0fSLNVdcKBITjTKJN30zhhF92rQTEqBjDGwGeKmrr6ZKoTFSl2N09w+gD41mxNh
NXLRUfGMU4H45kpDO0BDSfSKXvzOVWpMOFuV9lXJ3xODOfThtSfI/bKeyViZ2D9Ow7rdFSwx7lRe
K0uxgDB146u8FEawnwAdc1p9Wr529UgS8D9pcuWe/s2ADkzYx5agU4COiiwfaaQNx9zsCSo2eAqF
eW1FM/Wo+qt6BvEPQazGmsDy2bwnseW6d8AP80jqBydwrJALzHkHTi7WNUtQGZr2/JxItcmz8DWf
TP5AgIR2nkydq7gqgiIlt5YjEwhHu+cuojtiRenup4eWTopgPM694myZlKoePQRTzM9lxnTf+Rpj
ZYoQ5Wx3uUrMiXdeSfpUxXM/VQYQYbgglEWO/MogS1cMJGKZWmLBILjSb41llJyMq6WEaZxW8B8Q
+w3qRV475MWQUYlsh13iaFTKuMO/BqUVeHLCO24a5KGUHIgzKefb24iom7fGaPiHf5dbfPcICcBa
QUywqyODdzA/pZnzcwVbTF4TjJ8KoI6G2UzG2aUbwwgSazoTjHwheIkvGCrtGMPMW82150TixhZp
RYYM7wYaFOpiIhRk9rrPJW6M2gRiPvJfKGhNiMK+aKYhB6WxRyUBpA2ADCQggCZ4o21lSPTYzX1p
wzjEx34sZRGHBJVJg99Q0w0s7YUT3atgLNralgGrFPbkaQ4UUE47rekqjRp5s5moyP3u7K0S22uy
c5MZ8u3TX/11rzk6W4kuVgnm5fRt7obmeVnnKdi6cNQqzed40WoQPRNdnyPGf0hLAPnLSt00NkY4
5WA6ISxsETwr1cFHGB1gAMLerJdh/ApPjI0fxAv2Oxp0LYmLQYNyE3sRR6yCIU+WkHeG5HvLzX+b
6ml9sSpsmX8oxRd4Q5KjEJzHsOe/6jkFxwFnxpRGinJu1XRuuhmMJC6CMyInkc598DuR1D2XgrFn
XpgUr2uzr/utyyvtWAUkcxUUs8ih8IoRbKZ0JECZT0306TU++fEApQjrNtT1Bup112LF76M/5g3Q
pSH3y8oCtneP7MaQOeQn+z3P9FUI6IlQRa44/nzE6kR5fhVNKEJRta3/xFDilPnoebZNrPjrTI3+
Ff4ZApR12h3kiTFgnJXvcouGLvne6y8y3J41SiSmTGFu6nvczvXG89nzU3GbkbL8TYFgCj55rJbX
/LcfEk9Qv81jUlA7uugyhBUHsSfgwojEa3pgr9UsWhpv7tt1vO1zQK/S0tirq543OYsTAKAjYuSI
Mh3eeM9yeNkNxoGno1FclTA3p43JcQ9cMHEz5NzATvIHtc3nMvkn+KFjcsd2fkFMa6sWLQa6RWwV
wJu/yop3/0fRMDUiCyBJTclUkZlUWuaKb5XC9Bp88RqoTSgiNzU0QKNC3Iz2KR5ehTGfMWcmhkYj
P8n4rOv346p8ZsHY/K+fhr68ZDlvVWVc0uqPcnLmxIB60t5XGTZhjvPDtYeuioM/eA+BGEq8z7Bx
LkANNrtu7z+H33EQQ6SLqWUwbbek4eXQYjaG+iNxKrnbRBk0psidFXzO/1mBMMMTS44aBMv+iYeY
+rxz4GaTpEVuktRTigrfyUbfXXNGCEB5tlh6XlrhNQ9VotvEZ95n7sfmwLHpKZynGpZpWGw7DAic
MlVJabWoMcAB1Yqnk8LSg2eX3abyOh0EDdG7iSD7yCMknhLghGc6SNiHC4TGhpbn1Ew94nBJ++KL
hJeFaGs8ocYj56gDsmjfccuzHooJN/s1MLRpvJfKJgoyijEZpe0YR9gJ/or+3aQYur6Eiu+L3EkR
BOe6xBECzibY08zEtuNA6qRNs8e0rrhuZ1SRs2q2Hr6ePTvExWwu7l+D5r9cYvGzpgdOZQyn6Fir
B8oY8UhHfIWAW8tZp2V8JGyPSQztFI941adUWJZ+mEyJW1ofxIVl3rnzMdyeBbNNRc0ZP5lddueE
g95NvBbjufY3OgRH6brP/bG+R2tweBIRfCiLY7jjkGq7d8mvO4hdUqu/Rd582aPxRjiUseINR5L2
dGcJrTOdaS91VtdbjoC+4twPww4snqs2mtCX6cJsYZE7PpJgNzfXui9kE4Zb5m/BTjAc/1IjUXGB
v9PaDuwmsDTmCTLK4M9CoK67MzuDt4KRVRDG7Wqnc8GsOCKQDF84Zaed19vSyY5mV49v1dXZ2k62
4DeSMfgXZzeh4FGiiTvvrbC583sdRUOFyzIDvk6LPtX7ynXofJ9kcz+DJ8jDxFY64cyuRK1akHFw
KkDZq653Nl4c9Xxft6fzC4lc8wJl59IJ2Pt8Za358YZhjMDLuxV0lyqLQUaukM4LJg8q/Vh48xz7
17kc33EBMem6zS4by0KW5Gq+9bNHYRv/ddV4Yteooubi2U3V+UnfvptCd1CJyeaLUwkbRqN6PhHT
loARVflxUS37jBrbVNgIWATIDR6hBnptCftxMqEgRZl6JaJ76mepIwPsZCXBthC+lp0BeEEmujg5
sdMCnEyqEdRB5739IqWtyWaQR21WJ+X7UMiHpkv6270QZVIGaN5ddFLjsM4tGEBGIhtJK2VPrbom
7N2KShIY/P8QH7FEwCoXE4DWi74zAPojdDlZ22rB0PWo8S68hwnU/PpEgS6ExCZo9/CZNhB16/FQ
OcPN7KyyranN06vFE84uU2i3affEWFvQBBqSe+iriEyPMDl96Y7sChJxpQh05uZT12ZZt2/OK0bY
p/CNHW+6nO9cTKrQBd0RC3OEl5n3IweAP6tMfsITJKMCGVIlSP6C32LmfHId16LGlIXCyWlz1TwW
r0IXyQUHPSzdu0FSNKnBB6jxawl/6VqL9OUjaRalNqLyHqCBiyUKbR+S3inqFrZqid1f1hf/SyLp
SVfijRBLzvXQBYu27v/bLDNDLKQFq+/fD8R/GIGvZszRiZ+/slN6i8vb82lNOppNBE8Ob7iZNsqE
w/D59pEz4xltzm6ibNzBFbkif4DeGoDQAt7Zp7QPBIDHOGuuM26zrRd1rtGCN3JmavUCccrLCXO1
FJRbGGnXjbw8APDcXfZ8P3AsrMZKqBMko2m+mBTWX6gwgm+s+UhryyZb4ZVK1yXKnGVbvZkbkELZ
ylG0qO2cpJSC+oIlWYal13+8KwoxOXthTcR6kIZxa6bk9DOtWpfozDzSigzdLufeWYt+2HG6fJ08
mvMPscW6srB7maMdkDBvyMCKj0ZctlLKkMCpgBRJekqHb9XxRSrmM0dx6LADSaHrq5IZvaGgp30T
oLXI3bHWOUv9gTvCN1wDf8dqj1of6ZYeKapbP+4ocCvf6STdsSwSP6Z2a1/Hh8xhodQY+UP65+Iu
zsUvrBUvpUN6XpdSYj+dUKCXVUuJHA3MAjdj7rUjx6nbS+0beCx7Gc370MIi1Cw/kklzEjkWeJ+T
M+EdOuu+wasRoJEmNnnenKZJX6rsUpmLPIs+ImhMxWJSJuuWS+Gt6n4ZoJLMtFFVEQn4dUHHDqIe
5gs1R2dBMYn6ssS5j1c1d4BcmBQRLrVp9jp8dcBw3eUyLe7FIaMbNjjv6fWtyB3VSS57Wl7Kq6mQ
AD94Z413C0myE2n1uz1HUJe2LZLQBh9l+hDeq+vUsVipk4oP0RPv/suchY/nPZNsvJgGT83VEqZo
kh0zbebAtTQFkSuhqHRKslsBSopdpX45lsebJF6hJpH+JNMO2wA3Wv9whgnypHQ8sO4xlllIekJ3
PCf7+bYgdOK1aEbnTrRta7fO79WSiBmbWG4LR01e1w+aUuk412UAc665UQ0ICmi8n+avHcrdj+Sm
jm4b+DvdvD4akeWxQQAKpGWAL7qcE9/RIHHD0XXduHOeRyrmuPvAW1ehU0n0jokNoiw5lChPZ5H4
6Va9cpHnpxXxnCcZtgFlzRad6yIfiLVKMJJosaDjYxYqBH+4OlCuIxe6iqKStCAWjHxYTGFCntbL
/6pSF20IBloVsk2fFryw9NNymYzfXqBWgX5js6/LDLe7ti8BJGA2QMFxHgxqnLaj4QP2MvCSI/Jg
eq2/rY+UPUlEch7vS4W2UzV11V1lgR2ykn8OWvZZdske9M5ST8aTgV6uu8ij1jH+v3wDVZvrEs8t
hO1Nnhry1/+SyIbnS3/pfVkBAaXcXfLrtpKe8HOVI0V4K/UAM+h+FUxttU2QaCewiUaNw1QiZrrx
8eUtoPZ7ffZ7rXGz18B18aBN5Z+1+1IA3AxybRJWA7GIHmbh7fFDhtHhfw3cPP2bmesTqcBW14Vu
4HCddqyvZMdl/dTy6/hj6ZjLqz77kYx2XUjzRR+TPAdfEEkUL62ZCr8MdtWkUQGkkvlxYywpMhFh
8/Dwn82kL0R39ffVMkb2kqpdf/djfpZsqjIhBH9qU3frlVOM88VLtjolR27SmObJxkFSYrijITPR
tw6UOBzb0SIg8JMa6yh10c0Zr/fG8gPLfeAITGZnfUllbDmsChMgrXsOHKqzV8MuJyXOug87w1xh
lNiZbxge0voTn3dI/UNeca/J+Be/pHPPQ/UkVVw/BH6bUC7yST1tcNQchjF97io/RaSgMihZVq6r
ia3eRWbwothdxiJz/rDh1usR05H9P67Td/hrW7zE4dZXkFA+O0ZYCJe+nNCFvZtYbqoVfr368EAl
/hy83PiqdB2bboVYN5n0cKpsdVhJOgfxA9GKjORFyZVmII34rj57zQeha9qmxbgno3lzYrZu5yZ9
d/azI/YzqOb0v+cqUCS34TJBQ/WiE37beI5XBXb3+8iT9TJKegkTk1Lz51p2mAvOfKBAoImmuzfT
SzzYdo5R/GkRv1ymD4AWRRA9/xMc11Kri/B2MWvXzUwI/lZWz4wt2OlidrbMceQbB8hrvOjV79mE
oP6hhSDnvFzunBxBbAlwQix3hipYpGM+uaIvCYfXLCfVaDguOrSlypWDJTwCeCVZ3KK9qdpU5wiL
eGLVa09tMl+lmktFJrebVhusedSFQ5g6CJ7GB9BIalOIh5dKCooE7dgNVKM+lFsDAfH7hh2VWZ9p
zWIt4WF11W6B4a9isJp838oku957/sdBxwtteaB7IqMvZAtyKchkSnyYmQq+eC80lyaD9rqmqZej
6ZDPAmAGOlN7dUKtSttrtG+slbWvYCyYeF9AoO+uaCQFEY574pyQb0PjdPcRXvdESFXVke8yToZ2
WfPVvH1mMZHHvcNk/FihNX2K7FGSJx6BXHMH094WHjPvxY+Avi81YVm3GcosSNZQdnp3D5cegl6t
mNH6AaQXyGYGsi5xE7A+76/fZnRtSM388vX2q94eM7EcL5i8MM1TE1D00Dbw3TNXILIeXOxF7ihT
qmxQFPxv0L7ptpYkTqWfZs/pBsxQxaO88s9VnK+Ur7BmerP/JOkJVAKjHCyxPDtoorYe9XsuYcZW
Obsx8ZBk6AhF5vItHXqjP4njF7uTWTK/ZKpPYiITcOPTeq5RZXuQiYC7iLYqfoTEUxn4m9SMTHXe
Oy7lKOGs5hGKzdGkgizmB3klurxj1O8k7OOYbz0fTxOHV5xst9LIjj/I3PPQ1/JA0QJME1ss12Jr
LNXB5KZfmsJ5kBTh75FIoiC4ndv02dscasRJS5LX5PWhB4UjG25veedwk3w7Q5QEsdkHZlZ5rjdT
JzxUSPabAhHUH2EYTa6xam56TXBr/du1BBpkZu/0nzZqtOJUgKllk7etjgd+VIhf/t4Tpo/Ajl5A
MTZXxR5PVaGyvxpgSeLIStl718XAIVERmcYUnnjBPwHHWaaMGEd+8oPI8oiwYgVMS7pWyL2wQP8r
TYRVu78D7m/tYIMjwRggkeb2OxkXBXeXUQN94EPpPs7hFehqRFPCzCRPGYU29VWAHbTXPe8yrB0c
EmXsgsI3KQaz0/G/gMSVTY4ggrH2zz+A8S6TiQWRNVbbSpjcfCNRgdnjIg+dZPlELE9oGKy8DXkg
TzRPsFdewG0b+ppGOo+w701pg03aHzXMZNEhTyePVMtImRYAD1Em+HueJKEIFBQ8avQayFiMKtf9
SxfEO9U9K+Gz6GY/DWGE3sJU1gwCIdUTNQj0cKAZDMSutowrMfK7x0cRfJTp9SDoDCRGJ0PmJ6G8
rH0UcG5qMp6VbKiOhemRT1wpm2OeL/2GP7GcbGyOGYfTQX19zWXq/YanBDldrnWdWNyGGJSzRE5t
VCAG3K96xxB2u1iVXzLkl66M7HzcEwJ7jy2s+QOy6fBaS4fFB9d0W3n4X51p7msubmFHVBY0BATj
FGxvKv7uGLjnKM2Fwed2Ven9UpA+wqSXDFVIemE7Rvg3mztfLMcbQg03Kpz101lFw6JoV9H53pyo
1fdfaXqzi7gE9tgTghn2IFDZoLW1tXFYFd9iz/VTIiAH5eXnbCHyOfFu57qsuZZsFIBrQzAScD1M
8Lc4bgLosS+Vq8hU0DO7ck0wgrFLHfKOZSx9zjc/nxyVwwUqQ1/1+FfwX10rp3PEzXj7AlkBurkh
TFvay0A8xUw4C7bDBAdSDSDcpHhZuNLxxx6LZr4JMyUcDa5tFzYQcFUgjbtzrkA5opNVsm8bPFHf
aPwfM5AM2suA0ey0IRH5SYsVomtowD824/Qxd32Kl46g6GjC9j/sgwYDhQZcOFSU8plZBCrNdUBK
/JTrJGhXFanlXyz6jtX91KEuLmqhrdAOtGuEGDidi2ZcUC8ryEH+6UnW/yj2eV498ih/rff0fyVo
jLUKMJ7sH1kYRFKVW8l+4zKUN10615I6yWsWZ4/lQea8mHiyiJhLDEokHQI2L0WFlxmYpalJJRBM
3qvAThn3JLR42vzvGGCqWpIe/gfuRJ57RHAtDrEZs7eMFftYS2sgMpWdXnVySt6vxBdX/JwkvPSA
gZcVGzDGqg51z+un38FtT8ZCB0Ct0a7qaMjH01z2rJcNbkN0pWQGiQycqIeLfbzu4cVWlMWHiks7
gjj5W0oEZ8WwfBHZVL8jzltJhtik2XHzMeN/8im0fD4CmR6kusC33nrBsugBIf40P6eE0n9eCtWT
74kQDhkZSHXD6x+wliHRdmaXVlsAjGv0rnBNyPCiEY+9Kn5djWgk9ETpvVMrDdsfbWbJRqPhRcr8
E2/MANL5dDL5coB3m8XrpIqAXi/sLe0/fTvlCwhqvctOIROBQ0pY6J75uhZabshY1Z5aBgLxKncU
KD2PaV+6XJVTOvIGUscuj2+Uy53Pn56ca9VHJrbBIMHNaiGz8CE9K4ZL51XE0/VHmUnAtB1ficKS
F8GTQ5SG1clRzUXiEBolt8lzkvn8rDH5G6WgwtQZQbbdiiSxh5aHy10J2E7YRb19fxUJikwjZR5k
xWdMDznQrgV818FneoTTd4Kcpqd8yy0ppHKhYnoAyocsmXn/hjh9BTf16CjEykSeapdNEMoL8Exz
4Aqt+CSvbLeMm3Jrc6wpD3LFIMrLNI+nfE5G3rmI3O4QvvgZCU0uxjDWuRN0F4s9fz4b2XoJbRgu
/sXmReCWZuLYdlgyl5TNMcs0YcedpF0igJA3CgAdTQrEHaimtdsjJXCpNKL/9JdhamYR/7riQJGn
QMM8V8laX6Ot6ONGVsLQFy9Qk4ZYdiEsBmiNxlQK0NN2gwIQ60Fo28elFM9/4legR6AduEaMDBac
TLEzmh3LZb2POs5MNVvPn7DlNC4e+FhB+3ddo/z2+U+CC+LTEetKAG5LsYcilFCPppCrWAZD7hRA
eX6/umtpHvWE43fjSV+jfrGyK2DSz+54pxhOop78M4luqrxFuBRF1YtcwjFw54AcwFPWtHTUxPgF
8/Pux3sLb8Esy0ZdpMZFrVpRUxacWCos46K6fIy3+RulWitZPJGignTnV6tNfcVkHAiyH5d3uS7e
AHPGSRgvkqqRhSEAKxmgbtChH8huXQDMm9pjQ3w3pH+BSuezeDuf6FnaCvvev+8+IcAIiD4PvBJT
BH+LR9+Shaoubz7dUfnUve1AP6cueVswUZWsG7A3v/jaQo/Vs/5+hpbb9F/YSrQWiKvAcv/xleVh
+tLuH/ApGTGB6TaKBAHDpsOn7oEPrHXPnmm/t0U6EbHvs44nthMLvwRoVbZdEJgCAipNyXYUipGg
vtxNOrlwciz4NN3ME/tbbo3rNjCQSRrWJvJWkkiOG4epWYbGWpjrhnUVP+yTarzxRhuj6BoZYg1w
pcIiYyG+k2XDXL/uIt2cJTghYVsMNAv7irQWwNSmuR3WjoBF5uEEPh8hM7H5xi3No+kQ47jdqQa4
kqK05MUA2HYHhNh412FyaNnCZoyel6juxMBL7hziWMFt2k+TKy8mhQOJy8gaCM5cE1MCHA+kinkb
dLs4pDe0+uqjwvRiXp+K5krGaEX1Judn7Mb6vAsPJdnyrW0hzwj/rBsF7PplyCZvDitjEmweQsUw
CNMd7uOd9h+zCVtkv6LS122fA64ZsAzU6Jy1M2UYDN6Fluwkc9XJhCg1l8KGNEUZpQaWOTW3lB9m
iqmT4VdqooNZJAMGY+GO4wvM47eitAlblZo3nFM9lGp/mCEwWDlGfhst1FGGxWxRjD+RB5sYz7yc
3aaDvEgCGGLijeV3oKakOBGv1zbvlU/cXmh8oJc1htK69Mj5dAnXRMChTu+42Fp7fnLfOv9jv5RA
gAHI0AXasdQJz59HV+0nGC3nqbZ3ajG7lVLpPm4zURFDNUckQrFUg9AoT1I7YLOFQEOcOdgPsyDc
3UsCe5mxiJSjfD5mlNmqzUY7D3YdDbPdUDm37IMBLoyrXj79wykNmD20X52pyoWW3FMNzgI6WTjt
T+hSVACTUNNvmd1EnSTBUQ1wbq6ahBGZyH8pcppYmlqJK/B1izBjg4w8tdzksZoaG0xPYk15BDlX
U/hVwaD2+I6I5XW+oluNKjeBxaLGzIs786tbXAAtlbS99RqvB/l/zdwtuboC7tlO0zT3LDHXuyfI
1m5nPLh/X6NATDl+wuYrGm4JElmnXYMF14dSuWgm5tPyCbBMyfRCJ0JQfWXCKpLigt+5+R9kFwN8
S+HTYQKamkmMa3aELHuGg0vfpQ6KwjWoebojVFfbrzL1cZeocKcMs8+YJg1EU5C6PLbC9Gjy3FAk
aXEPmvvNOaeQ39HxQD7O7KL13cQh2SNsuYckf4ycW8x7R6PWKLawp4SNkZH/vTzLrDoMdLq+8WpF
kMWvaR/wlMkNoX90zTvSyLqrKhN6wBEi4zeEnY2Ai7cDMvEBZ3wVgOArOy7/Fl+gYbk6I9VH1aiv
FMkMqGdTCZoc0ZkX8DXyombdXPmzW8QO6yOd+njt72jurPY5lfQx4dgmgVBIVCOrbWqonWgI8H0C
UckkQg8zgSF4uRkLFGj6ovagijAkudZzduAbGHV+GJMSzErrQciv+Y8qjbmrheiyxmfeGA5bS8H/
LfbXCzAPh/Ryc/i9vXRLUpDPWfqmGGQaI7PpYLYJlcWx305cjY+FVgwsEwhX9hTQynAMHGkdlS44
W3gukyi7/B/PKq0Fgmg8ZT1FKqOlNxXd4o3JSUQbIuTS5RECnKuYtfjYwDAmPOMpbL/4bkK62uko
Ka9LVOFsV29Ptaq8+zea1hYgiDbQtCdZuCjZhJZCknpgT2wRctzE5dUuAkxJvV7dWwuHlHsETwEd
Ezfk/P9mYzEFtTdHRUUK2zd7RjbrMSutdUTJ53ffF+YwhZyiGuiB3fMcFLmH28Z27CLroOjNULvv
3KpByAwzw00qSazc58D4ETebV3zK2F5XJjRhIb48Unq+MHMw8+Kuat0UhVsplpKqiUPihe2lnfjb
/Ykcl8/O7Z/DuVAI8rVjt5jgsV5EBjbt8lkOHNcHMK00M1reqNN85zWaz3JBfTsL6a4zxb7Rf02c
SibhChISU2LZmP3jCBlOWi/Jp+TqWXmwS6BiSuSUTgvH3iT2oK2PsnzAVl5raf7BzztWL8iLCCxF
YrOjTILGkUSZFULAo9TnsbaxliTFqZnn/cptgvVeokAyxKguPzIiCjzPyhLYMdl5we6dhOpmq2aB
4rkU/IfDdwtJkOgmJQ2DJ4AhnFRI7gjfr7QQtGXkGpHQyJxj29FeaRFTggpKsLw4wmAWa+lXufDx
aozo2aqqFfpKgZDe8Up5YM5srvrLXu8j/ACjHZ3ZYRHZHpFbzQBQW9iEF2f6gcFJlM919RkASelO
LbW4Fz8RUNBpqG+QaIyanEhUeClUJLcfJvXcbKF5g8cF/iqM2UgU01lwRISgyTHyTSgZmJkBpyP/
U4Ute2ZCwgwhyR3fzNR0cdx0CGLmhLPdYFlGqKJsyr7ZxOLu+qQ9EM4Uz9wo4jsRu1vR2Hx+m40F
SnrB7nWIlYb7Md9Vr/SoJgcw6OYwtkOZW43xd3nFhLfpt87miF1ljOjFnZ1Qt/BjClAa1X/sm/ur
w+Kzx3mQ2hfw1vcr2bO/wojDx8pS2ntEIHQ1cQGHAPCQuNFcVyRuQmxA6YMABZySqQgQ1ZGyUjtc
uW7rhQfpy3V5pjV5L8Ybknc1osrZXpg/fynoC+kg/GIwNRQwhprvqv7r4vo3kg5v4dGN1z5fD/Ns
170aygNcNHPD3IT0LVibo0deDet60l0M1sMIJNBcX8VgD3LUtsu2waEiGNuJ79W+PWu43v3jbrU0
2mriOQL75OfxGjae7/EDglgT4Y8jEE46gOEtVVOQY+Cj4ixZlD8yo7XK6DlVN0wnEheTEul/54jL
4zSPb0SBNEsDj/11PYqZZYuHK945UB3vDqFnlDSmQWSsNwq58ktRSDzUzq9rkkW+4mi9sITVDCwW
aW4NB2eBxfej6e/ztUwJ4i793ipcAc8HCyQ/T61FuRqYMyhfeFOwX2L4rUssSmnZP4W+VA8JL9X/
yN5J2DooWK0pP5i31rFwX+P9PP3BQHm89kgG4j4FvBOXWKyeBEMdoex41pe6SzDLKNB1CojqbToe
WKguZeSOpnBUkS3UJQ7JEC5CTc6tu994vJVeyOu5QufFghlw4zb0gGEnx8PB2jgoz4CjjV5BRpbQ
biRAdFkuSTxhJFSUXxOLhITe2EKoXCcDE0K8jkxq3dFu71TNy8kL/DRu93VQXuHy0fUUjwptSB/p
m3IJSgg6AieKG6DaQONxki7X2gE1AjItk8YFmImyLqV+hFZTQ8UeqvenSDXcQF+F2ucMXC2I089q
odTAck1Jy+pV7ccD7pwdcFaeUuqLaA2DOMCln3aBYqpgyZ3sh5X0A8hM15gmVmyXtcT/jtteD2Av
KcS7r7VU9MVg3qCqQXFZnvTz+9le/OxxFfLDUt32UzMIS1UJIfEd4SGFaYAWSbXVnVb54AkyLgFz
HKSYRVpRRUw/8W25ZSgyFPvFPMyF7rHDiR3c1t+YgpwiW1BGrASKSUMQtbMczuQbsx0IV9h9witf
GvX+gpw7iVCGSUQ2bOB6lX6gBJ3Qp1gOdfFRYIJBtLYDHzKZz5bajvbHu1Etxb7o43FjzQOsa9b6
RMHZKWY4mlDSG0rU/DiDEbxUE9KrgH2toQ1SImXphUD5ddWploct6jdTcs/We15V0ihgZR1kkiNI
rcLXrD/IQRVqtvz87XZ5ZcT5bA2fuewNRSkbt/PnVToi0HtneTwGJWq3bq6FjNmy9GyXlq0vS+aM
ooxLG/flFdclGx9r02JRZwOlLHWJp9kofDj5eJOUbaf6lWznZ3e3ysS1H9JDV5wEyroYibgOnbG3
P0NExnG9CljxsJdqpb11J7uYcTuWsU5Kkg34tDC2+WefsTtCQD1+9cGDkP0maMtJ20Az649p74Qw
T/SULnBJ5+iba31H8ZXbrgSzvrrOSXFPIn7zEnVQNQg1JwYwYXsmbx28LXKBypksisT7ShIgTj6w
nrmLGevGsaEnx0iB0L/VhC2sAwWaBMui3WjqIYbksLOH/GNOdNvyXVz5SDb9iqmw+blx0fNbFLF8
xWtnc4U+SKkA8Ez+QEyM7qa6qz3p4EW/KUnCCh55O7UKM3NoyYmzjjqs+tIPTN2Bzlqf4xjwa042
zvrO1e0pdPP42t1oP45AWL6oLraQy/7uUsFXtvzM4pWHxCTNzSQbHOoDUhv+tmMdFF2Newu7Fstb
3FX6vFdGdbXGET/LxzOH5TF73IvZMfcVOefFNsiVk7Yfmc46bCn6Uig8kjxeciRpET9JO+MMPsCT
FCbaWB2auFW82KdJNyWSZj2jykUMBW1YuCNIkUB2T1utu62cW2eQWRyb2C5tmEjXcnWbKFP+61tD
xiPayGmp22k47Gh6dk0N6QXU7k4u41BCY1nBb6eCrAQsanHBzp6XfpZ7KrWxuI2V7MrxdqnGdflR
82xzl3l9IAHtJB+dk9ATHywbNWCLLsNIQ2rjOlYvHYz5mnZVCtFwySNOWpDa1VHjZsVjxCNXNuE3
VW+BkfnzCqP+fBc6bEs9oVrAjKZpgb92Y5LTqQuf5FE/HhM5pblce4cowZ7bSQEWxBj7h0G7B9h/
1hfzt9fVHj8KfgdbLoTmA6veyGoqhbNEnW7WZYZvY/vQ9VY5aOXYJU/wDTIxm3qGjNqhMwygVmMb
my/I9Jckn10rJkf/KETcHxRw7WkV/GNeJNjn5R0hc1UiNap2N069NPPKcPgqbap515x8lB7b3svD
gF3JPfDNpfqJghIz1QfsXGkiM7zUH3Bz925xVgNkGxUZDwLlvp+89AfbdnCXGmCmWPuYv3lmAPFF
KX4iVJ2ciBkDNDuS6VUC8VYZEkGrZc9fwn7VMnxrsF6+Dsl3g6c+GT4G4sPPX6heVDmsTB1EYuq3
8fxGs/DObm/1sRougv+3MZInaaPi/sSOuFvtdCrNRcSbkE5G7lhd5tc6cfkibZWhx+0thCpoAsUC
Nk7aA14721PmX9iyTWSi8KDKK9p0LHj9JHLANQig8f2UbNVtSAtvqrmMijSVzYpecSpixUWVn2N4
ZRriwMCJ8kVYAkNlyiVFGEhhQtzishHdteKz4dkmKdaV5ZbmtCqk7TZPte3/JHggf8WyoGCHl1k9
hq+M9pkk5CBHE55EJixb0g4kR/g9RzUHGXvFGuWzK206LwdWq6nRlqmHUZgPfSkdz35M2EZ3AXNS
aFzWXMdXiYhm72LjKkDJNkKnIs1Y13NZIcutmMRYHwNa78z6a+WwW1UxfosYAvW+T+KiwYaYL9fA
JY9TWKzeVZjrwTJnfruW62BDIprKMnKi6I/8V0qmjpgSU+JSFbGQh2e52rv+RWdS9sCV/BfbXqdU
dpRydYp19FBrINVkzna4/pidvOFTSk9fukwZ4YviMDpJsY0MZUUSoj3WlLTD1ey89FYJ88de+Tau
yTgQJj3LdmT42b3/XjB0uCdjbb2APZLjgkbawbMpLB+/JJeS8mmt5JW8KAOTkMLyv3pqEIXnojhI
QeWdx2OXBZAI7kNkUY/vTfphP9bf4SKdqVSbDU1N21AgD8MlzGAzr1MtxzP9Qzxb2TvHN3hcqSIh
kBiXmfhQQK/23b5d5m5c7UKLZ9h7OFcPL2bf3MePO9hti+5goFBiFhRXtQkxEcdbKr8oeukStlvz
CZoEbGaNOJTpEgCmt1xxJlKrh0yKZkFvs232971FGJ7rQcVDymeXrN/J6Ht0n0cAl7AtaGnyr6qF
tFyODG2ewj7vzPhJWhPhpGbicWcyCapga83mumfFqBmgZwwjdhu7Vrd7cU4RVRF2r8ZwggsZkRRZ
V8oU9XsY9YKw0JkUPx1h8MoY178F+P3zBdtcG6QNzSmckzUoz5YJGJOBfwhtXMZ81EawWcxJ+tZw
WCcy337c7HUFbeWr1EiQRYlB3LA9CMIelfHbLZ0l95TiiANPFB0V9MTdAPjyRuEoNmN3fMoiG+e3
jJjjrsiThmwRaSQD24XDw4vilFhnp2kgBDMpmn4248qg6pJXtHJY+OVuoZjxwbxcof7HJIy1i8BA
Vmujw4xHZulalBbmDgLpiDJ0GLHNTTXIZA7Ej8m9wA1S55sMD0dvxpkqFJP+zPgCIrrOScXudkeY
03zZInUKuUDP4XHESdJIqmKHaJ+hX5nhZ4dG9y9T0rgOReVV1lLUsBHR1nqE+x+tWjgM7/An5MP7
Xym/mlZj7DFe1k9WrAxZysMyKbA0hVgQgbcZrDecbsQg3oYY0h+GwsEoQ+wIibkX5bnfCdbPnJ4c
WlA32ka/V/munifJksTflytj2SgTBCbxTgSRukzhzEqbY0PUPljX2cDuri0OkEuXAPrcYZwWgxJD
555WaD6zgRpnu+Gyv0Tw8XRaMVG50IUwUbEeO/iBr4qW6GMgOSeDCm8igep6eTfm16JKA2KG0uRS
ysmzUXCEMJboBMN29BxPO6TQYWch6UllKKgD/zhOmxpar3GClhn4DhWx7NkIBole+JW8Cqz8rBE+
9DSLPvMEsXeP8D2TyEfxA027vn1IWQrAmT2YRivB88adJIphdqn33YSE6kwkm12xhQYPNlIp353H
AtmHycNCiots9vIn3skFAwaHGIBqSEiuMW8NJla5z7S2sOmenKzzcrOB0hYBjr9NDtbbi50y1Ja7
vDTJunGJlFKrMj2bsnQRRO9ksm1FtbEV3ZBDsAnxVT1ERilGtQKR2cYe2zhuet3xylAQ0+lCGaZn
lWqDEKkNy8Fvnh4NkDMytm6eFkRo6Irp8JAm9GIUj8wZgzZc6xy8HPIaykvly3JYRQd/PfEnbv4k
k3QBSTTy6uUFiRWwL+ULt3UmTkyJ8Yp2K3bxBTYL5lfmH83+gaYpRCnFOiBGcZ9iw7cpsA7vFMLb
GZ+bPtLN9UdXAdSWq532CfxeJENLV56etw/40M+txJAomFzv3kYa2yze40e1NzCCnW01kdmbOIqr
tJegivvsukK4SGawG7gknZU92c4RKOCqM/6xTOB3YnU1/Ty3wgfkltScf2M2tvGi4KoQ2r9FJurE
8KkMWO070e2HW0xBfJjPeKs7NUn6su2bOid1SGJnwsPRaYMacIB/3p4pu5y//IKwH7AglSgYS8fR
mythk5CtSgTg6yiJ+k5/lUq6TU4feaecCB9gHhUVBdmCPiEn8c8agc47Q2sOZD8hW8wSLRCmRDiJ
tEjTftso+iYT3qW7BCvJaVwfJqkUNntMxcF95p9rVc46S3dVp6bkxf7SiwNIULalTZRqO4mPo9HT
Sg7Agt2bxmGCHTg7YZS/28vK8+6i1Ozs/WACYMvX6v+ofW2PyOlSR7yip5PyN8d4pzyOidEqebv6
mrfa8t5/Tl15JyeoS23zt4Q2BcrGJpguSTHIN1hiDawCaQM9xRtlYafCa/fYz8C1R1Q9IpPU3XQp
zkHa4mS8kRsDt2/uFfVALh4GQLcEMNigkDGQUNY9p6zqNRYCTbckYNMXzMS/fwwN4Xw52N0BpF+Y
PkgtJyff6xtRsefngycxi3OU0pBkXAheta+LsryPuDvXC2Mk5YSQzHKFcFClR7SGBQ5MnPlJk78g
tVqa5zittNKjwyPgFq6UE5U/kZmfpQRnkspIPJrhQ9H+5OAGWN31bw1mog1YHjY5Y11SSpryMftG
5b30pzcHBgLNVVzduUfbjHy7niUk+cXvlva/vgMWaXs+myfKDXUrGDPg1IZe/rL4VfhAA6ZBScI8
sO26NZsISY7ZDUCYIs3piatEkL9ktrpFj18Ryq++oTBStamiz7SSDwwCsN7SGNuwDOdXoY4cScjf
Ci5j4gCl6PJGlXzFRkSRv5PtZeny4OdR1nK5YNFNP0mI9Q2HaprGJ29GivOVWv/6UhT17Fv0Si4B
GDPOpq3O19wXdC9AXMZn1znRNLQPKniWvl7zetRlsYJ0bqAplPCLaEBR4Ua24yGZw/Sg8qNUKWBt
a6MCEzU0m2kwznVKIlo/lBzIpGTdsRxkPDwb9+VsV+gkz3HleH8AvDbsFQISQVckK0465tmr/4MQ
5g7Zs0VDJvwyWBD27NKqybsMbiymkCyU1RVDrzv5mYLpRiiAi+gkyAOwi9atHYudojlr40WnZVjm
sbxpp/A98ZHaIo0AnhuogApXU2cPStCYH9qG39RTvh/brfd6T2l274jhU8jmfVgPQZMyzHK0/PQS
V1KxQQeZSxiFO7o2nBBkdF4hiNaYzICp0FrnsUWsaVS+Ua2ZQZokeR0w1tFzFp4Im/e4rXBQpdx3
Ij+izEKBie0RcgSSbGhGzuB3tV8u5Qa99dt1OvqxlhYVSO9SURXj7LRtUHpBtIg2i5vvC3ZZepnm
8T55XnrYrWTvDxCzdKR1hj5Jou1ZMRKpFSf8vsFGm7K25m060tg2JdXgigqB8SE5oOAHGMARH8cf
VO2EuhB3mjgV5JcInn1okIhWOYgkPhq9Zp5tGsOB+IO2VJcvNNFLgRgvx2yuMrXMB7saO47F/e7l
pPPtehFqWcZnKthGr02/k0h1eiBUy/0bmMfT6fPyWPIWAq+W4iSek7yNqOkRe2hGx3QctzH4fkE+
glueY3pgp/YMkeKAmCamwDrH5HH6ST0zacIX0ukNsf2f4GK1gLfdcxToMqQvd8uDzwKSUaAL/2jf
BINVkOjgEAjE7PkM701WUsg6sFOqDSZX7CGKBPpHeaIVsE8+nPmi1NIFqVdeAQsVXpfEkrONDCme
LYn1TneXDmcCTCEux8YxFNo9hD/lpChXuataFq6r3Yxttinw57dOwkymUoD9i4yxLGAXHPvYAfY7
/USIivWGqv/BZ3D+NMEvBb2QbmMsLquZSxdESdg7t0txei2g0eagV8WfS11Z33o2hc5Ic811SVLn
6YZshZ16M4QqTBWVVM8177jD59RC9eY6brlgPajcLEV65zXIJkYdASd4X97kmNGebUBxbDwCYu/2
RjSR+QsqzY0G6JhNQEuesOQOlhfoIsXO2ZntT9AXniFHb6r24/f7Nml9MGHOq3WpKCuohfOFwWr5
lL2GOtDvV9QIvIYO7pk2H508DBUEUN1Aq8zhS37eVRg3jdKgihiUZPyzgK/wFv5GL7jTWHZ5MC3q
988Xpo29ANIZG6vXGRKyhJ5idDdBrliYtQjHYk+RjOcqrCBTz7Syz/MTI1ENwH/7pMyKkrXtZLQz
bpaBht+wY5qiY6WmV9XtIyHTWgusLFYafqzp9k+5YRDDnMp52BQ7adrdNTIUgaU4Mo5r1yLJp6rF
/1RGQt1XXHw1MvEErxal6z48fNsRupoAsLYuOfXWq8nrgA0tfo685hvnM+YQ1ZJ6/59sWHlF/oMJ
Dnecfm/xjH1sBQuGtJAWZLc6qwhr5bk/LGFQ12tobM/6npvMjsP9kMLAsi3FeC3Bi/GdouYQYSeJ
hTGAtmMbqRmMMG4QrqBQXju8Cr8kko1RdGbhsk2e5WBPbKJtakfv69pWxDqlvNFir53xjJQqHWDX
N4cTlWGhN0ER9dph8fticshK59M555AItKLihx3fz2U8cATiOqzR7r9BxknU0Od/YjcJ+8rXYE7k
aZPzqiQUCM6FyrOSC6wwwgqBl/tQe4srmbyk0ixd/sTsYEelpniZFrkjyuQDydvrmaChpnFFkzBQ
2aVSJcSMP1EH6ATVd+HcIgBjSKSAPkpkpz75N07efVFJczL3orlPI60iw6Q9dV8tCYFLgHGKAXb0
v4W+CShsefSkDHp7Ep9x4IbhpCAgJeBMgQKvEG8yfSMcccuKeu6Ni0qVe5pc8abaNEWfNPZ/KhkE
6VPU56yeVITckxL/Ytq/6nAwZ4rEXFFui6KSMtzZyTkxDZdtKlmsd/X7ROvfkALQWrbT4VAhY5+C
g5vugUmuFCnH5xJ5LcUbQqDfGxo9C4B/5SBj5J8gJW9+wNplySXM6afUlljd8BAQbbbsggbDTw1q
yPJE/8FpCaEDKxKCJIdhRAe/4TKeldywO8CG+tahA9brTVqZSYGtmXKbaKMcSGLEaVREsIyC+4f8
dFrFcXyNpejKP8NFaXG/3B6pnZ9Jm2AbyYarE6hXUfm1yQuXItK37qjvSvHZXUE/oCHHP+VE+gth
O5ed+VkB7za0YBZm7ZxFw3IAMucYSXamfhOFpL/uJGiB2UDUOsYP7CHhw8Vm8jbZiIvaFaArM8Zh
yL99WKDTDZopL/qvYLix0KtR+4cIW6dbWye+PM4WLXZESj0PXeKHAO59kOB3Db7rF+Lxn5FE2X23
b/HvNnblt9PryuPg9fbgM1CWa40LEwYYFSfmhqd1zmMDcCHCDRWkahj7wsB5y3of2xwpRYum+hWT
tkYVyIaIdNOLn1OUyRiawgQ0MQ84ly593s3cOBzilzee01k34tawBrAG3ypTayFj7KJRQRgCiZC3
lF1dvVRYnRK8QFqw7rVuhPf+JTL9S60r4jP4/Nhnr9mTdLJc80eOIQ7YPKEKtlpmoQGdOaDWV2VU
GjCAzC2X6qURnKnGE6toxmdcXJzo/f/Gb1U6GntgKjpUmTsDo1iX2O+wJqPxr8J9Mayqk8HrzgIO
OKOJxoNX0lS3mw1ydcgJUTjUqyoCLn4iyniDkjKrG8PQLHqbK4oq5dgymH2WpldnjOlLLii0Bp3w
5BRNtxPT3HEeQWHfK45/7l95iFo/Q8CZy4sl4+pIIuO0fhUiwgsfuAH5NqrFchjgie/5QQ8iDvMO
2XWUNUL369Wy+0uekGyswXlIV2SKawaRSj+TVSe5239EdDRiuoT5GecsRmKEv6G4T2fDP7gZfSU+
J7zIs1h3xYRs3xcflANNW+ARCZtqjvu0NOWjdGAKQy68PEMwqNOnpTfqyty9eeteXvWCZkZi7WRn
d9yoJRp1BgHgCVbeZztfY6c46pJz0V2tmhgza5C+KmZgqXWgo2GT2VaFdPbEduymIjDaRj2EtW/O
zGaRKmRnamQViIYLBxx/gNTai3+q0Pg/r4d5PUwNK/rMFIp/58yYt5PUwj/jQCD+/YBziQFSQR4v
dGar9VLsTJqzuLQe5Myat5opqU07ekv+7sXoQi5JEpR1YzQq1zJxD9QLqureNuozuuzfhQQd2lzA
OrKS3c/a2UE0YId9XA9xnbslmmwhmwxNMTPp/lxqcoPOZepYUoxsrwTJtOvKb2PiouwOjgrl7Wad
S1nUqaPJDlIFHA9AUu0eJwY4fiptEZs7DCfsqu5tFPlcHJ7/0SuUylUK7LqegjfLEgJUIELXA2CA
+4BlwsGDPeOI6txuAYaI0LuHOTELgbwmbfhtP/adZSiiFSY32KDoLxFWx5Z8tmmftNOx3xVtb90B
8XDgaaY2mNi/Wu4sVXfzjndUkZDWW2i3kZGwahB5U+l8yTCzb84V2NwMORd9Apet2gdYHie9Tu6c
EBRvOkNLxRAY6Wxzgx6AJmyQis3ghcIhtXy8EPDJ2nFWvOd1E5i8z7TI7riMxjZWs4FrqqNgWx80
yUpwCMncTXcdgbaPMUcKf7/7cJ8PBsRjx0PrV4w+fbg4XMb8Hkr/k0pqGH/x7Zc5B7Dn4eqik0VV
N3vD3QPWf9ciurho1vGwDjT493j/HDFXdzoOYRyg68qyaGHcamwYTgP1YQycdawHv8G5y8PCFGS4
L/wLMDtSI3TV8I5g6951gU3GXMeXYvcLfZ9/K/PSGgcLxJHKnA5LM7bYoBU6kfRBS1kq4EfJGr+X
+lxXJG00nI1Bm6YCG76Ru3A0QG0Z+StEHnSQFMabmmr0kc/t1n+9xCtLJw0bbwnHgZqbEQ23OzqA
ic/qLceoagjMT7C1jgHF1kkab/TIi55fqLa5EKn+dDdg6lVrNgpVa2kdctmBAPhc1ac58XrxpuUR
oizQaxfsIjA+5iLrKF/UDeXtvDq/OiHX/RlB5x51AxwwEc3Sl5F+eg3Ij1Yb47TZecuG/6F2tPZV
I8rKT43+5Ef7gVW4HfFvQmxnQZKXo9MmfTmDHddSodkt86gOfkkRO8NvFOfgqTCNNkDNbmu8TvNp
tdqmAbcCOyjS/fPIClJhBNiIlycQvWy/pBpQzHdMaenDc5SAYdrDZkzjcj/svmID1os6pyeLWxHf
D1zhofPSA/blyVRC+Av+pl7yS/6cBhdmiC3mJxDtQFyDzPIRlB1Z4Ra8/hQ9SWX9Jpr9cigwa2Lq
uBQ3bRTx5gCUXXgd9Xv/4QWfwzdAKWn9n2RXFrm0D16fWF2Gz8Vh1svjKc4tNnbIXZIHV7VpjyT/
4vzuh7yH8ZzjAOnx6cPSDciz/SXemcHGUCMHJ7gDGoBE3KojoKbz555H0HLETPK4zpQHeK57N/u5
5HXiOGiyZDm3+7vrSMIOlI4301yKy4FlBjK2hst9IHhhSiknJWhrluUKHDMaRKG9I2ghmu8Rdl2y
W2uYsDj4azRWSin/L/BS2KzPXqeuGYuQEc1aEf16d7K9tXi4y4TIO8fxwpFEs/+JLZYPsS4JEwPK
g3rtknky+m/byhjYvsHmsL8GVUK1x4Gk3hGZNIIp5RMPORgjqiXaZqJlBjOfYQkpPhvA8b2gcNtj
PH0pl6s7qKDjayQHH5zFs1H1oVoxPAKreiYqVoJDE3OAsORp028yDdssv353DCE8+lnN9o0UXKIg
fiIZNNaYCidX75BRIsQFGjOcBOlL+eU2Xg/429f8CLqOIsZ02RK6aAv2hemsWz4TCZaWJ43Jkawh
kTQ0Olby9/aeE9ozrFZuavwjBMQiH5Ppc0dZ3spDsN+zkGmZFFHwkHXGb0+HV+2WWoqmERxw9meg
WRPUBobUIdDrKbApwZZdoIAIqEmF3XnLniW0lW62mItkm1qaz9SKInB6OUIhgmqAADQrpyb/qsFU
vMHpJnCmgmMglplqKeLtb5GRMUi7YEIkMrQL5+tNOEbwxS4hcKlqxLPFoCThCeHlLexjk6/iVgVx
O74sOn4SuevdjmngOi4L4s+0ZlrLPrO1jDqX0OEDRShwRhAhikrPTyE/OgmRGBQe4x+uyBJvgxT5
6aRCye6Qa2T+K+iWTtiYnEhGihP5K1qRgnUOrIJsH72hXNNS79xHj846AewuB0PXFjLiJ/FW3D1o
ePX/XHrBFyMjClxIM95zG1nuvpjDPbM27uXcaMdVJ7/UScK9caAXnVhw+u/JxHI+SrU3sE1LDabN
rBTHAG4mPfY/UyF886VnwxevGeY+hDVIPAciwZR8EGovuNRH81oNbuHq2HFygCY1/SHA7lkpzWOI
up5mJtpwnKGTvDXN4A6AsHUQ3Iulj0NceeVCvF3hHqu9THvUEj6dnUDzXW3qPD2jyiTQN+bC0qxQ
PNV3NABWmaAkfzlrgFBd6YGGQwCaRzW+QP3phBKj0A2x2unAYbyh18A/7L2MNe0ysSa9+M6YB03k
gGYoO5o9AdRoGE6Jiar0kw0DdCfNIUYELBrj5kZn0epW10mMxwuJBnX9rKST8OIWigB2k9sSQtwR
I14ugd3wAIUMdGgk9Id4FdlxeMfptcaPtpniO4ECYmo3lQr50loljJuSJCQSyrtHqjKHtNZG7Z85
zbLTCKc+bfMUe0hTo1etNXnFVYCaidRyKtYcqU9X0kdFMoG9jzmDJbuK/mEAdjtfabZEMC1RVncz
XqRHFF1tMtY5I+lKC+quF4LreDPxEWWGJrFmTrMMRaLcVOSL35onb8AoN4SKLZoPxhiKgwQdckeT
y8DgDlXREap8psj1L8sZ4HYsFe2kabEv8sd7ISZrL8cZ9GmetT1wP1RrIeNXBgHjFfcfUhRCzeHZ
9Od5NogOyhLI/OdWrzIm426R49pFlLESQVs4FwWG5QiXuOE4dRfwLRxOWGo/laz7NiZ9CpUGwkPg
m86yhxT3idLsetE6YYBk2YtUGFdKJVHQLBZHmOJFoFcPhsKKgAH7Lk/B50hKC32ePRNeaklada7X
dGemJEOX/7PDsS2NqFTsYT9IH8t3WvICFw0Aq1C4brhwjGmYxsexyhIymsQ7mt0iTA2ZPDxEj2Do
j62cNf55vW4IDfNnDUns10L9uSEMJVYjfyT/OeOHiDjICHK6nUU8qwDOgx3lU38UK09DWkC95R/8
sFtDd8cJRgruPWZ7IXaUgAHstM5tWjY/A2xBpvB4T2qhZHQXpHQhAfD4wA4VHlfg/hubw6VzpH3z
Uq2TN+Nml7z4UkThGLLcdFrzZucyE60sB+Duih/pbpSwHYEid6XqAdc/2n2GJ/Sk7PHMFga8Fpft
1jdMs2hXpIHccDLGum6SWDND7piPD6dR1eOXONC3/yJq3Rx/aBmMmJ6fkxToNeM4hC2zVGqeACre
w8Jbsd4AJWDjp8Ao11msuQfwQ2QbJ6roEGyAuvDwBlxpzULe6ya/laql8vYPL77tHFcyYL7uYUXW
He2bj3YkJEq4KFOxCwcnFR57po0j5r+YPTw6Jh+y1I0K5bEda0O/VZGkJsU1kBHKTCpwKStgF8rX
Uqal0hl0R8lsfotzTMW6yKwiHV4W7yJNZGwDeGZ8TVLTSY7KT0ay8KUNUQv94Z94/On2wzIxtq/p
031RexjFxuoapfW1/zJFnQJhh2smkTBZeh3iqUJcQyU9YKNnH4gNqttTUWZcc+ZSE/NpDgPLgipQ
eN7lBxzBf0LiEWK0SjKwNAutX59JDq9YxYYYcLPCdY2G9N1ZrhQXQ+JMkqxDoKyhocln9I5ft2Yk
+5N2yFQKtJiUFaayFgmUH4yaKK9FVZBhIH7C1f7ojr97m7qjLOZC3b3A4UfHSiuOoyVP9fS5Y6DI
ygbRtO5m3Z2vgQB7JGM8PwKVrs1vMkLIVK5iFemLlwC8FE2TwLYQSzAEe2pAG2MPa14FOSs+pe7h
zMyttMhscIFiA8COIelOpHd3tUiXnTeHA5I/l3CR8uGIzkv6UOfYle50EOnrg0CL1Hf5HnJfmelz
HjybV1Q7jq1R1wqd3A2Pn0IUQeKvd5m2AY5zBS4nt2B36V38ZbGcOAOdnIWPkLxu8d4/AsiJ3LhY
5B/S4FpODi4EYgDX7Ri1k5BLeTh6vxnJqnhl4aUvf1SPfs+eISM2QMSopJ78WkMR7zSOWpmL+EEL
AaDAobmer539Mcn3mybHAO+kpLz1ECIFVKGctyUKEWqtDC9FpO8vTMtVVHiisNYxs/4xUBE6b5JL
wQwKpVmAg8sHgiSm6F5qBhcPJLlPSmN9W9akIWMlaG9cDGxSSmJrY48TfLbfC7HsOnzhNBVnIt3V
ENEnMSGjHYac6QgDuQnEY8d5RE4b1YA1sVmxleIdqxZK9SOhcbvE33rMtWv/m5O+/OfC7E7gNx33
J7CQT9fOCzlIDZlhWnPJepyZ3WkcASlllDoqJeFBGMfMEQpSGxz3cRXaJ/DnS5zw5J5gsN2V6gXP
UDXqY7+dbH36FObP1gcXUi8gm66ZHGM3t0v8YIIfpyOIG/AxOfIrTNjoIX1AYmmnmyr843ibrEtg
87TzHaI1OI0+M0vivvRwmAZmT8kcWDqA4BKWUvSv/pLi9BJuAbbgVbsj9tH+FDYSu4B560H4rPrp
yNJwMBIpddG9ZC3rLObqk+mZ4aKJ3mhBoOI5NO0aLNe2Q3+PT9IVnW4fxkb9QXdi8+AepvwFBIAW
THqadbN9yTFfVj6narnJfzczZhh4iODe/3zuR8JA2mJSeR6/Dn1DIyzh8J4lTTZhBIdSx4Nh3P0h
zrkvp9nmCFWctURuVKb2y4yAWmwlzIXd3aVCcynHRW6RD+ht76i3JZGKlaMNg3NgsxQIhFZ+EloV
WyQgfwn7x66PQXKvfQsdDDST6ETH4xNdU3TTT841ntvrQwjvI5t/R/aNrhn1bU/1U8ZPSlVEUrGg
Vp5UbpOWZ2PsQUXK3p8NBlALO/TEb/BuqaRcvUuho+nzXkb5bLBtFYrN8QgnKEYuAddtpyXdM3/V
wZuHNnOK9yj0J22tq2Wds8JktpgZJMDryz0rWF1Jh2FVOTrsYjYDx45GPGyGGId3dWQcePfvqKwW
sFOFaMcZc8UjSyd+MuTtP0JEN7ixf7OY1uQnu2k8DXG7g2FaYAdwC915/7sVDTKRI25VgRm3qflL
tt1jZ7Fgme3x6+KhIa/q6jq7PBLA74zgN//CNrxW6FNtBq7kxtG159FVezF8IHcfVJFL0alA0uEh
DK2oLlk+zKSlmGm7LUMQEAzf23u29mGCNysljKJrI2/qlHnjXjYAJ0KyOwGyIYOOGt2656QnFO7x
QHBYzC5cgFihWG7udFMf2x30YgWTRcaUuGh0+tNC80WMNg35OoJaJb7zN1cj8nCUrD1QnFKT5wkR
ilbwfrVQ/ROaPrQ5In/7hACyipts3aoEhE5F0NPYZyNq6nbmm8tsWq8av1CMnBeFAUNLm94XwRLv
wnGtVuceyabNqfgmD+UA3SVePpvUFm1MZUMC/X+Cz8wHyQcNigb4H30L4F148liBlX1yX9ylHzRn
RbuQiJYLrL5Dx8/Y2saIJDWxfNPPf023Y08j7rgYqVyXXbeAuwLaISQfmf/+UjBAXRXpM5cIM2fF
sOXixCiH21mU6MPscdudcxQ1sE1yhQUuXAnDUQ2InR5HUpdyoC8YNLgz6oS1mcFDCbA3NAo3paie
eS1O6j9lJytygIUNFZkmHbFD1Vp7TnnK23Wk4X/1bf7VhPxuXgRR05GoycfALun6Re/Rxzv84nUt
mGDu8jtxH5aoeaM1WXdBaZRLEdIitALHtwArbsFPTqiX85YXuWFUZ8JgDeHJUxpwJ+qNrRzlR9lo
c7vOrpJeueufp4mbonkDIk+gGyd6EvwThK5WmQJZdGXtKZ4daCPIGdIO9VAR5mN0ypNBBbvKA1m1
rOpbfMU6MpvaliLPyAen79prCsmbpnEvCPsIEcLXpMPRgdXt97bIYCNUrFFXFzUDkb5FoETDUouh
XnrivEMILCak8ldDjLc7apwRt4ogBuua+h+f22UBbdltrGVrgfbq0p9F9EVhX1Pppvr+k7giR+51
AVHcJqwRdTeZ1CoGRwOkLC5fJE8S2w45zaCF3OGoMDX0VAim4yq8prh7kiIAE4900iQgy/zVKoIf
CstllTjcRjWUT/VcWV4j6G9Q2NSLRSRlFFbpecI2s5wrUGCWQ6ta6Ir0DtUu2aJJoShgp6li313a
PQd8wvgJVuYsWxltZsrVpVW148XdsTVZLz8669nrrwTH9bDALl3hIg3uJXVNxq6dxkmfMjwZRAga
U+ZDA+mPMi65Be7/M5+tenIMqy7f+HX7LqL+Vc5mZiK3z3XQULvHukWWF6Sqjs8wWEMEx4L2TaTB
jA6kF/J+imiWSwGaX6k6dRQUYaKYT4EC956AHA6Zy+ZFm1G6tP+t7I9NMNtLfcKMiwJyjv3ynFcQ
sfq1Z7kSgloY303jaJ90YsHX2kL8Akdh4H3W0THT8gLo9b+KMIMZp8SLBBzHPYQfb43A9H/rEuCx
iGDOmbaBQjNdsSrbRRyq+nDOBcHGYdb2E1nDhJldTz79p5hqsB7fv0P0pKjfR0KoA36XvqvxgawH
biQscVzIrktenmbGhhUHke4Hs51g/Q2R0YpBKIT3YlgULFEssTQaWifcM3GpEqEBFmWLXCohyaQQ
l6wBU1brx3+dRua/cisIZuYejiWEvX1cAoorH0jGMUDLePrjIIOJsGWK/tWUoFjc1H26kgBFZhb5
wLm41Vo7zlEewfLz41FtDedBGNq2ZKgq4WaJVKg0SqwVDpVeXy66diJvTJ4TTMd4ESxOiQMEo8jG
ZNMpvTFmrocRnyPORGwjKK3OsVOdirjmSpWz1xCfilbV2fc5IU1/CGINbs0mif1pWZAefcUc6FxJ
t+SXMPlGDnQY/dXbStzdlL2bLt1JQWuO01qFWXFHQhhfxLeAdcMiTLrTW02heNOgpAuQ9YaDdSh4
xvxtMNz1oph9Fvwu1O1Usnh6rFuSEwbx+v6N+TQZKpJAZJ9ycgI/OoeNa9/xZLRZDw0R4aKpUeg/
/9YMUtZL8AxlvALRNftlOsRNeSTvMUM+Ajf0qMClh487MYlAe9ajbsiEBJmpk7DksvNEKrqYPKbP
jzi8reLNKz40aVZPAMSKfwztZrY4QYxHo6xPIXD8nQbxr2BV7VJ+KuO6YoIvcUm4mUm/PeEl7ofM
9+o9LpuG/VxrKLgMBNfBrgyED7zP1OejI0TFKPxShYKjiwH1aJpljKIVXT3GAQtJJb7l5WwIw+5K
EUIxw6dVjyv/D4PijLurkawokapWLPO3ATaxE5hnEyQ1N1+HxaZ39CSMz94b4BfrDcFdM7lmyoiT
Q8y53sccILfyOt+sfGiP80WyL2KoG4oTu+pDgvL5xPXsBPYnKXMOol0gvTsPUX1xBaTXqPriN1LO
1N5ren8dDZT5L8Re33n1OhDSmOHGQ4ZxbmoqrU/wCylwuPxtyRCmYYOFyWF4cBYnwsUTlpB0XbO/
6RUgwD+8GVZlspMq6lGm47Pp3xYQ0jYFJXTpLTCmFwBRvSDzBYyCEimdvIIXWgE1xXKvTfWVTOI5
wuxwD4PUlEdkDJ3BLcfBOffBismT0yiv8ARgmIhlpZAvT0BRiFIOWMyfUFjxIdmjyySXw0ykxprm
P8Up2sr1fo/SwohigkGx4Epthhh7Yorr7BMnp9r6tZxpby4hDnI6/MlEXbtXA5ZZFPG/3kD+J0Wd
2udKV529LO62Jul6lGRuNjSrXMLRCq78wwjMqXWD1ANaJ7fv340oj2VuWJEc25gTCkrgNG9XHB7L
tLYOzyJsM1t0EqKrm8hLFT6Ad19fLaGrN7wJ44PVv5Gs+J4LnfVCWsH6utzRRyFhQinhcRjN5lCd
IeJq5R0eyM/xPJtCTRE0iM8CjJfuMuj/8CnugVBclYvnDFcpf0O7hQYfid/BLpR9mskV0lWTcwFB
boIsG5pPe45afp9rRJ3N5jN8juUqqnMUtrPPF3TVS450sCJSclnwavX2iu+d6U+tD/xhxiXrCmun
oxcb2Uf+99a5CGc5+qDLJ8gtmKU73TfZeiCSIQXDi69KhJ3ricsoworLZ9pa3NmdpmW0Z1JdGiWo
ENmy3k/CO7hHNttUFGxOema/AFJqrEujELCsALnD0oBAUWVh9rX3kdjx4/hME++uSWNA52BaPIWw
HeB4oQWBzAVLPORhrjNxsbdQErjZp1j5aKJ0wCu3JLrJpQrsqphww/CG/7ILFfAoLt6NpgdpwKP1
obHhYPUaymqOADoKNN/3esHFZZM+4pgFdpUnIMWfcB1VliF/x5XzePYACkYH21EDonYolACUrjrN
HXUEZ8eN/Gc6opWn6R/iieq7zTwFGYhtDOz+PwcxdaYHDyy4tbeIyO41kqG0dnUarny7KxtZVWCD
dzrW9b/E2QwAO+gh2j743J/+mtb39RGGGPp8P3kQ6qBy3i98oQ7JVD9MSysZ0if9usk8LVX89rAH
yLZin8mxRV90j2weQZjhY4Lw3iFnAQPOrEhaVrCrV1NTtu8v/u2mJg38zcSiEUpFvG8wpq4nnseE
QBuOcD7IARL5DTqDtQtfCMURZ/35M2LO0ZrAF3IC274WJhgmcuu43JHi2UbXBMZ6Cxk5hD9/qVXI
gifRRtcS7xm6u5jyYUn6ow9uCEPvt1J6I2cU8oAv5LcAPvaFGrRDRpr1tKAEz7bZWunJzf7KhEEN
a3mAWY2sdzrvU46m1cmj1yZceM3IXYzGXzncHgFNKsL6yk1ihOBNzzvgonzZNQVdkNo7HiX8x0dI
XYr81pxnH3iaDR5rIabX1P/+nc6YSANwApVWspO1yKNIYCDAFOVJywTJmx/G/pSIeRiYXJ37XwcB
1o3SACdecv9Q4COeSFGu27qRIqWD/g+c50VWE9FufSywrBIQUs3Jww6eyCIuawf6s28tZ6ih6jkx
C95uEECcXSSh8BiBioenJaTgBsg4/64KjPIEo0pIHP78PLoNLTKo/3dTEOw5l99LrJQkBiD1xAOv
ACYnvm04D2KSA9Bc1sHhdE2XnIssdJkIf0AQC1wyDHIhGBDLh1uH8KtS4ihxvjcTM2iOjUq1oMtt
3go6LGxfXcFxuRPDdWmmN3Z0p6inG8Bu/zfMYO0uSFppcyWskbyUSgXzoYpz0PLXGljE9YhVHTMW
QwtA21arvTANXiVzEmRYg/JoXNY4EjbLSaqDC4f8qwhs3Mdh+EUyPkMWtOsDlXvmT0/MADpqgzgF
ZHNpoHVCuDIZhQeJF1fuZp7h8bHskWP7tn5xmJnJmE6GaRTQPz5UDPftfD0pEzD3MsccuKS/3FiO
GKTO17IqMjT1AnBm+Qupqh4WJ6i367f2S339vd2tPO5AcWu117Su27YiS4b0cqtJ8dFutaiJNXsQ
+x9RbrncPK07m5je8oFizwaeD4APtvITgib1k+IBW6LGAXSrb/WGAwd6r0Mw3AR1MAxb2pvpSHLv
GHeBhbcmJNq+u+BMKb6fkrBV/SDPv/naCugh8pevXw4yYnoJoyYYDdg+IxKIhdU1lVmtFdkRlTJP
1ETPLEkFYog/l+51gUT0lvZJEsol5ApgxXZbsrLTqPF66SbO+oBqAFGeXPaWXOb4213iDkDo3t9e
OS7M/XQrkU5qUfm0gzR2ZGo6O0XWMP2vyWUc/2SFvlwLdFjKbAkxBt+0NDkc782+ZD72RFpIOBLo
bueGnepXKKkPoVIHIYDy6g6Z5BjHxeGV+e86H2y1iKC9M3FxSNBUZwncPASZNgqSnyX4tc11PDz9
zCI8cpe/JrMRz2Ue+1Pl+0Eu07vx4pX9mKZGjUc8W/BnjrYCYalfFE+KuX6kXrnsvsmXTu9d4oO/
CH5mex9brt7xH4Tp2gRp+vfpixpwiskaH0PoC21/im8ppvGf65Pn1WSYKlnUottKKc7v5ZT1jRWw
Jr+xOB5jDG4dQnUXKSRwhnpJo7WePzmY192GLxRr4wWmfZBIgTTbX23U4ifRdqkzyQqkjxT/uThP
VkPpe5teDj81sf8L+lOZhDMelERRZFUYEmpSQaFkByDkr0piBty6JFZyJCVhlJZjAZvKq8nMdJHK
S+ynUUJ26vLNmL+G0BgicM0ls3HyVaCFrCDpPhMGeoudsTUQXT4/hW+KAun+ij43c/rGEZPHa4Ge
WkhhN8OG0RwcYTS6AF3nddQ6XQEsrlY/VivrbIW347TLPcajh3Jq1aVuyQozSNlrwH3ny/lyPHZP
M/ErqjvPHCxDyIOLBLqD2ZSBzrgubWB8/nKcD+tcmRi17MEu5BW3Z7lcb+bbSiaRtgeivMCEEueK
JEisvaAox79EhcqkNqaoFd74L19IgaS7ENP7k60osVD9jmMyOXhx6BhrABROYfsq8sGAWLjgSKGL
gQnElmjTaEZalrhMP0OH9LqTFTuFFbnWLgonVGFBPoDL2z1vV/DBiafLb2ORarhhcyp3HeAXt9cu
c9z5qHUfbgeK5AEMhXBJvYYSWSL+rcudeJ+A4ecx4f9A/ewWRB6Ijbr5b5OWiX6pXks7ny1mz0hT
kb7+kMmVZd/k1dMZJxQFo80dK7KsefHUAENmqAK/zW/wCtvCkybYYm5Be8Z5GKqWxmVz88Pj1ggx
xiZqfVR9AAeQoa5PIoTF/DGhAOaffBPDKFr9K4+rGAUPc8f8gGcoLp9mZrAH1bxaj3ykSDLbJkId
ULBGlKRxUsafry2l3sx78moC51uKV9c+Me4v+kURSAOOPGuda2fOPLY1Kq/33qXx+NfR4Z3Q6SbX
3xxet7IldUdzU7k9a4TIenlNS2uAr0DQc6dYA6Ikun02SWzeMSn23IVExzzl0W9rD5Rm4F45mm5r
29Eh1llPgVTHw94bXi5OiyFteJI+fEOKLGqx0q/eIEagzOG1q/RD8acIj2RmfkM+yvK5IBnY7oYd
B5wOe6IloIqZalUJyo29AMF0eZQhp55hOGPw+b2kfPV3JVgdJ+YOzEV+G37mKMNLg0/LDskkIRLc
Euq5VdcfODh9NA5o6afvMb96i874T4hwTycEZQrGmPhYM+ma76rCY4m23Aqs96gK5DKmkNfnVcuO
czsEuGGXRV16+YYBt6mNhUd7c4O8+tdyXGA3QRehZ1XAwSnsAN/uxjJCTMsHMrq3Dn4IHQZtJRTV
ECju12Nn5Iy5MyBKS/NREwEBT+JW1jRfOnN31CVKMdUSPtBfOH/AfgVf4ZJmEFAxPjb+g3JP+QuN
YJXsUACaJbJQB8ndEqFW42F0vyNc2I7IVIWbHyQybDAHZdcKE4KoCvr2mRUY1QmjJz3fMUvB/RJx
0R4oMWbwKAFbeHmIzDdxZx1uFMcJhAezkWZvbO59srABzyQtvQIU4I3VqStwjYCX/PSKGaePUJQs
swWTJ1ValG+WB9mjuBwIV2Ev7AaqMnBm7/hLLPW9n41ZlY+HrecS7YUUZp5cGjKYk6Ar9XpevFf1
lARmIxBj2KmLabmnjsd3CZl+0r0iGuAi8gDeLVdh2FWxVPsQ4zZljrNKUM7U8/FjNoAniYCA+RtQ
1QKzoWFzFBvwvNol9Fxcmak+pFmv4HAnHItLkbRl/kXMn6ejTgbyq60trbYJ+OBMxfXHv2tKZ2ec
19dlM68mao7SsLkhuPfSDLMnqSK2inn1rJoILHfzOVabvRYjKqYUCohPaIb19UEI5JgMnwU4qe1D
sP09M7cJmzgQPWS33/86Zl1qTHvnrxl6jMiZ6lQ4Si5BBNA2hvm/sIwxr+S+4CwFXjftBKsktX6w
904uq0fWNwknvZnWs4ZdNnd9ObmxJIE/KaQfoYBEGl+0BPMqfcvkGo+Xhg6N8iaKx0nCz1MUTvYP
o4HvR0Ouwv8pBXxrCRVr3yEyYHhgOchdU9vLEKP/OhPqOEuFNHCqvp18dn5NPlQJIvtMWvUyukiA
XFAIgi6A/tjs6ztWJhhseoJy0lCn0O+XimZ6q9KoWfk912izTYvjcpRFVBVsd5rtydajCs4zURI3
YfjZ0D/Qyj+ubp/JClizWt3L2hGC6SU1bs3B+7e8eNS4jILQ0Oz8HKYkhbDNegNFjpEVeS7E3mPK
eFJKT2z85FYHXHusLhskmmkePUcpG2syEWEudaUXSdXyKV7txruKOvfF7xsovdAebT40T7s89LwO
Px8lXZpSv3l/GaXzfeM2yz1yYXC/0TFYBU1ZDypACSRW4p5mTL7lGIPM5Vj5WeG+yzDObhX3f3R8
OB64p3gz1MuvPyggPxo1/XEZE+sK7Kc56WxY90yYf5KGkJjfKs2EMGKMBKT134THGjbrDUvAp1xy
qFU5pAKwEBNxF2FvJvljYa7mmeR3g6JS9oh1tAprYPqA1E3J4Add1TwAgpi2e1cCPEaxHZyoJSEo
LLibizLV8Kf9mhB6rULHHutdZcy17IwSSo/lXE5yTs7Jf9KPA24JcBDf4uws+GzvALw7FTEGu7VD
WbyLyM+JnIbPRjg+8PDr0hRZqhG6AHuKuu/f7VQta0pUZjFn6mv562YeCDlBIlPJM4JaIXIK3UBe
WanXSP6ZZF9B0NV1YFXAmNjKT8y7VCbbYADrivy2G0pUoypjVrDYmFnl9PDaDZfoj1ToPCSTGN3h
pa0khZGXRic2CD8w1WSJK03GnQ360tEm5ScPnxUZvFVcwyWJ6qNd69tv52qFXa+N5sI/SlE2xtZU
0LY68zO0GpobrXSy6sFw3iHJFkhe3Blm16QJdi94z8ZJylBHIswtrizw9wFB9ck4XBmG+v9Bak0N
pH5LDqnziV98JxiSmsIHNag7o/WBo5QDfHifbmBs94A5+gIgomSbtFLbu5Vy1Z9gsbRHcEkQS+GZ
9Lvb7alUyy6ItzE0US+5A3haCmuFrh3UrsATzJmm3fgdd9NAf+U013BQAJE3zn4skuAJDYiFDPwS
RH1kMR01NWIB7D0+4NKEsB/Fe8rbzPE0+GPjn1u5k69PeQqGWepLSol+Faym/omYUAW/pkoVMBHL
bOZSADkGpgwZdR0uNQ3eokujjxaoXYohEvGOQcdbUuRBRoGs5zYA0VMAWsx2xIF6Qc8afWbTiGZX
KdxgAVRzDbmLv3ib6SJsEdrSow/nPjwW+/AiYXj/pRMIeqv42l7RN9eCf5t7AGz9Q78nq03Cxvdm
bD0+9kgElg0gemrpQmYZ1a/dr7H19Xs78cgEiP6f2xWsV/HKfc6ktz0RNWX2VTvsQkaRBXlMdUXt
+ze+wmvXEivsy5iBFGUCbmWyH5VwvM1jOmcUDBGuJMEB9cD1hCOKHq6DgPdi2G2vtRCIrxuNWuNZ
EJihUJzItgV/NG+zWN0jk+PMEwFYDkC+6Wi29cD8eNeVo72+u7DvAk4WlgcteNB1PxnvZImUpkEO
XIRmrA5dPYMlPa1nJhsubCkP2uovVS0IvWguKpeh1G4vNcoqxUYD2Pe6clskzs/h0Pk7T2DtBfnx
MMQKupLI5GWb4ydvG7/H4Pda68GUcqG905v6Tv47AF77we3pOD8bbuK2aKFmcdU57WejT02z4rRs
8mGDdjdr3E4cf5Ri/dUfRx+py3oo4XRSOvzCSc/CfosAS/+RzeO7KXR//W285D7QSwHsW2WUAMgg
GF06Huum3hDmi/ocANkq2yzhozO0eurTzI+YtHdmkBUilFXtRtNPlHSjqvnRYHHyEx202z6xMfWR
1UNUsU5HqCmirgBCs4R1H4OoSGvEsnFSRC9tgIhPyRHyyFbR+pqcsB609htA2uGrClXdhndGYJ/+
mQmJ0BSBcqoCJL9v1S+4hkUqfmiclFh+dutCJ4I6QpNqabT/9bFoj4Da0dioX8vFgbgm22p6lDJa
7e00sXwpw1H6gRu5ZfUCCSVEPxzkUKuMuHuvfeZqLWM3xSAyC6ECewhp18spM/pyzlpocobGaYqO
cOlxFL7Zpk9uS9ioZEg3LzDPf7lJ3v5o3zefZr3OX66uPexzSRqFbQZIb0hSKlOLa8P8DzhEU0yw
5KHmyCRtYQvRo37TuxDAkw/sCKYMsFeLeBRcRDdDFJacZA1dIaQIggvZ7FApjFW21FydWBBR77Z+
ibCncByMLSkhILFRc+7mKqcJO8ee34UYKOdLfQF0erGg4h29cdoXWwhVZRLawFZSyUdq29z8sOPn
6glaCW/822l7lDTlMma0vjBn0QcqmYedN7mFE83KCu2bOuO1mYt/a90IRF6dKHDzwOyBOrYH7L/+
ZXMKaVI1Zroa8ia5J8Z9JsDrtkRUAwJxDPWW9GK8prQi+mZTj2lJ+kIO756PNAgoMD0i1+1p1FsC
n63GoLVkvT380KFnEi2iuTC5SOk7X91t3gg1u0bufuIYISWKo/8lW0/OOd7hDrRFDzE7UuxDVltB
Ms1KPNNyczfFsqbxR9oYMrPB5m1b0goaN+YgRrHnogfeW47EoSscqguRdeyTSywwZa/1myEVqRJZ
5gC4dISt707BhNkvw1OLkcTKxioGJnz5eboHm/IEOWOkvehFTBWCkilx8STPwTZHcOrJ/KH41MHP
zan0MnUtszVFjt2yQSpG6IxS5Ot/BniXs2Nd6smileqCqCJmw7FJ+cZpAcJS79IAfOmZH5dHvynv
cADLZALolnDX3a9v/UDm5yvh7b3KxHoj4qnKG2ff3LPNbyCGnR0AvOTg9fB4oCfxOG/RYUdblBDv
+JZEVG9v3jK8IxRq9UpR96C0dZ875OE2C1T2lKYnubqmqOj9szV4zbIwtvi6nD9oXCNDMyvPiQaW
r8F+aj75r1NtbdgzOQGBVA/xJ8xDptP7pmWG7/+WRKk4J/KGRih69t5vlzeHR8xGFd14t6bG0GI4
ttYQd1GdQJicPkYdz5p5iqeiNbnbetps5Ro06IxRarR3WcZChSE4URX5S2gNKPAOeYX9H0jtLJP1
3nzRo1sy1j9EfdwIgJ1oGlEnuxsOrt9wLvuBfJtWRKfQNy4LH7++5uIEnUJtsx/CZuejGgLUtXgd
2C6X5mLxMZePVdE2utkYcRQy+C+jCj31vYF16uowwZ1DdVT8d3w14/FxwAczRpKC0B7njUn5EfEv
83B+BhtyoUg9ZThix7q7u2V57Qv4JMuBp+CLKt18o2nSP34auL2pwDiUFt5zbT7lMZN19y3HVElL
DP3jvjB5BbeHeAG1fOit01YtDKif54LxSsqdvl1LNV6Mi9F0My/UCK2Uv3qYNEiFn8HPmjgASO5T
hQYDshI1DXkR6+rcaKtsn8kdFfiGzJdt5EiBpp72csRQayiltQo5BOnTDFqeEvtoTebZREQpRvaF
TTmdq1rPEgzkmmCIesmdauJIP53Au1hTI/fhuWG8Kc9z3f4ZR2EugJlVtcRvTH1TUYxi1Q8NpkDW
0U2WKO8u5XeM3rgEosvoGwClWLmjggOsXD3RIpgMWO+57/MVaLqqsIfvsWq72lfVppADa9Y6uIO7
+bhXdIrsD3Ih7pxBC7+7oMQF7cCQTBqAQTpfCIzH/UMUhfOeCMmHmhQKMUbVrfW4Z1SBwJnYWYm4
3RdEY2s/0bxPvTv3brgaKBInuqfONqLU/9ZgNjQG5vEvBCXjLkWAjWgTA1TIFmX2n5iIYUfHuq8W
RUG60ODBjOO0dPX+b5ERpsMC0qN6DfCPg/RCbP8yBCzQAIchccExQeqdUTEE/O/xcXYsY9V6rmWm
PD9pMLaa6zRRcJmipXIXX2uDEWqnOu9Sut038UyWGXaL0Fo9kltu5qQ5daFV+RvvXnIiCxVjnBAF
dCt0duUsbYOVFupMK7skZD/tGTJNGTtmg6mJ4usJXepLSK/v7zUXaBZMUKJCSIrAi+XwnjM72hoR
n+/1JtqKeDJIW8qAm0h/bE7eDh2bLfy6DEZkcVJq7YdidCQnxCBz4b2UMpcuhT9kAOwZc9hfoQ0P
daD5cUMrav2muXHdRLEyzjQDD/Uk1rs1geISGNMpiNmrvDUes5AnRayVuqInqJ5R9TLDhMx4hKJp
Y1igc85Nk2T1ZN6ydUO1+AhvNZvx49bxvfksxkZvnTyMLvrEmeFW/rCe0N+AvLlqDBkRW3Cm4o/K
QIvK50Xfi3MHErCeIOngpf5rJed3ywDC72yLxbQ5Luk4NdwgUXewugzytsGMC/RHESNrR6rtcm2c
iIV8ohokSb71CrFP1LGjVg7V9Sfg8p6Jf5/AMLrjxMzsITb74QOHHDNIWpby9E4QShZ6UlHb3cV8
sfb22W36lvMbg86Oe8EBmPf+07oyOM6Hg3dFVFRumVUd0ekE4u7FKw/uJMVBRGUITQjTRgs1EV6h
ARTciVkZ9Yq/B0iMjEc2gNrv+LJ1zkK3LqPti4Z0jYhBuljvdFY6uDYJXsgkykOBDEX2M9PYLNMx
xgmErTb1JnAN1ABqdrNNqicHXPEuPEIPQmznDA5nRLWD1v5lMVTGOX6xdnq/6GFWvjlwfmAfxxPH
SGWIIAISNgCHaciKZms1JMtfewxvxLXZ6FZHdfAhsqRun7aXNb+8lmg3TBmhdiHK0e+px0m0UVYR
WJNAK/b5Dnase2dwuAWDvHQytBEuuRz9+9oEItj6mlsFU3CCQt+ZieYuyswTE0mek/fbHxYuCyex
9gEsxQ+NmZ3Q08PIQX0NXoM4bzJtGTxVpAikSIL7bGHjflT0aKA3Qz5Zhe8QWvxAGtBgAsXCLzZP
Bq2pzDkAmACBNiRM4rDzLGmiZ7DTxeGmctcr4niqYV+v1CKt4JYAiGDiXZ41qfe8Zor2zTkZk/wH
peE/dOGkBvNL8DfOgEP7YIesYGGI5LbDKXUVnnW57OanCern+bLrAm0hSCe8tiQwwYrOxCXnPIyl
RiyYrXlQXnRC4eX3Cvrx1EaSR6qaXmJ9e2cco8v5qkIEfnOqDKLcIVWXuA4HXpVpHJwAfDREa6oQ
q/x67XWp+0GnSOvln2E/UObpOBYjTuesW36GAgiVn+/mA4uxPuQdz4+IhTd0wCYCkekJZAZtGaL/
7/9lqrf3o3wwqiAgMfkfSTsP8Ij5HOIUMbrA4ghG8K0nMpxtEM1ourqounk57kpZOUPfgKnXsucz
/EEols6FR9lGF1XpHUfYFdIlIZujTftlieFoQl/7pEPDWQc4atAY7uoH06PGKSPxT+tW1+wDPAqL
HxYFbkV0yUY/aBWlfr8/2DIYdRo9oCq7S+TQeXWcT0gqEymPssQ+aFxsk9utk16WKg+G6JbEJFRo
Q9y7Kt//KQpIRh/jdUEpHg8TcCjqBs/n12siXN/dXXbB056IwwMtRODzGe4NgvfEFbalUfVyCJLJ
bre9KDMKpGIbX2x7VSVX9Jel+01kLyPcU21ftzfC6V+paXWt6+jyZn7BZT17pJZdMxDSgZmM3fSR
MU4+F4sm81lweJHRaNmBbLmjbS/MZg/zoowpShh/vyhQFx47X8+kNZPMtlWEenP+pO0Np/OCeyF1
00tax+DavjQB/5GBWUholncJ2S+cuEiCfukPwIvLJzPbVCB8FcI0eHMSbGweh/bRN0AXGWxuLHy6
oYp0v8ZkxR+cSH8NzjrXU5JEdNGF0pBNZxegGIaDPQK3go/7S19clLKi4b6UjzSq8dfk8xEq5JK8
KhCJ0vYtmMRrUBVQ2ltG25aHz3wd8BqWFGhlQhe86PhmdhHkcvx/7KjVl2XI5tMYhcYDTaG/2XNs
/cBe8WJuc6OSM/UyFxJAYbIz3+4kJm5EU8y1iEw+SMKL55DFwI6vApkfx9OJqxl5KtgEfSLAxAL4
pBVbrmlvMA2Z2g2NHczDE1X/Qc/ix1nCwjUsLAFHtzn2UJdbpQAqPB3QlJqS11GtAfG13lGEIPbs
GIkhQdds1humbIwsI59Thxk/1Z2A0FP3JHjZLbCRab57+cJBuBvE2fUKu1UuLWe3Je+evk7Ly8YH
EYoU9uzM/jZN5taTXeMga/SGZ5Zr2QxK7og/JzqEWXvpZwlNgMsUajQDWVSipC80xqsp1X0/OvDs
Sb463SkUPUHG/XerHicivAo2gMagYItVAwqMgJ0OGYJz53WneZOs5BMPyvEuFQ7tjEYnRQwEwJoz
IKsSdd4Jy5Ot+E9X58HhbBOZUGoBW3wBPvRm1WMTOfhDZp5jeElOOcPf6uaL6gE8jzjC4xrc1e5i
nSXF3EZAHABi2E+3gzNOP84fn340HxQHPKCy/FPJlm4rUO1abdN6/b1epdQDRU5dn7qx1mzPHHQN
iOyBzd65QCmrwK94PkTHkzrUGD57YZHTdqKUoV2X6VxU6MDZFPKAO1KiHK+FVmf/G6LpMzr7Xto+
tcGR5YdN39qa2xjQT7JLuqWMNdmCGfFC3i15IrlHQX0Dze+6FI+S+WmeIiSa57d1akGdMPpTqxd5
FW9lmNXqLfjEFdCWr4CcbiGV0N9v/DjDptQ5gCUKssJUf9TMbdDgXwZQJZMBvdA/82h2NPFepVNz
9ets0BQ1X1THQMMeuVmsDUeW0cfCCQUdVEwxvgEKD3UUjBrT2TrJ6qywEORLSn0aHwGhyo3OZ7Vh
bHaT5ktM8hxdakO/O3Rlx4WJBQtAHHLG+2E8XiHmb2MFj32GJENiEqj1Tt9OnkfRVLLnXqwdKewx
sYJx0jIJ2JG20Biy9wmc12itYGJfWTBPnakqP75A+924ePHlN3YvRLZoYuTpmfphBcBbOJGyyRgC
hzcx69RndRZvV/FUuyV/IcInzgJX7/odKThaM2vhc9txGUbd6O5VlNYhqCfvq3Q8njZnEfYC+Mao
VSK67fPctaDEuAnuDJcHZw49luMT6HDOKprikmo0DWdMgT8Hrd4yzGsBMakGeqYak2iX94+5M5jv
8g8M2CpUNZVfrBw9WAJKHHUsPl8SS0/RGgn1KxHZkGULhRwQ7OYkAlgOQ50qNbgguZ4IR5DSLQC3
SsvA2Re1vpFj5utYAVdbYxObBC2czFHU59EfNkuHT4mRHC1DwP4Dp/V2mznMggfvSY+j9joQSWuf
wFd3YZ9sf0BszLjIkh8iSX1e//6vZb1q/IY6aq0hEZRIEl2ezkQpUOpQxLc63iQfE+oOm6bdcz1e
EOoqcLP5WO8vEiD1jO8um0yNXiciE0E2y8uvvpXty1/lTN/buFsBT0X13QJ5jmNOdj2eL0jzaV0X
lqum0OU3k7d9hZfMrlPCBgt66dNVrOtiF5aEVQThzr2Y0obZI1jmoDZS5AGKvS/UPUpPojPu6tHS
xFHw5CEj0FgF8ettQogUlSM57ukQMI3YoAQN6MVhEMiF6kO3ho54QXcogWO1xPqtNzRbYU0p57u6
g6JAlLZkf6c9bJFf+b79oCf7u8foeQF+PbftMsjCJbKS05d7ZOUSD9Rtqk+8SoVU7Wkoi+CTzu9B
tcIiZyjbapHzA49R8yJASKp/2e3efofSu8QmpGzBTmvgihjBSmdPIkMc63FVMDlwUhZBEmgSrySO
fKvMxL1yDw8LwYLzdDE25b4r8JHKPZMKY02btFqhiZIHckeoBNDCOrh5hd22ZjKlHOR1hcXInGTT
l+9Fs8IjqbHbcmJSN5/jjIjuV/W8gC3mWni69ZyYHFX2wpQMa4aeJYaHqcD+Gz9+WIiiRnvOpuPG
7k4vZZfHqa6ZdboBNLLJ8l86iaHwmqzJEfrIHFHDgPsGVwwkW7GhiFQoUfB0xJ29xR62eMBLUPxO
osKvYDDiq3zMOsRFdBMJP8LkM85eqdg0wFUL7Osv+cwRtaHhaT91kf/fZVgInivtJf/RtWXv7GsX
nlv37yaJeTCF0QrUhbARBXa2HdjAAY+m/+Wcn1WLcJb/5c6jJ2H2JBakYddmu3oVJE3+YLt1mWWx
CbTBCsals1dp0s3zlhNfib9PnCvah08zKsqUSbAoEsZL+CiOIVkg1vGgBnwTBxiLI/oWK5RCeHIB
9PT6ziHa5KrpBQI6EzmiI4jKv7pa/L6hlDbzRzNii1bUD3uGdXkTU33mNzpEmDHWuHKeN8rNOS6G
Jvu/Dhii1KqeVq+hwUb9PFvPxunAkES+qoMvHTBgA2dCs7YFomG/wfUMD6FHroYGAy1Ty1l81WXI
VfShLZSlNEtWLITH+4lbx19O+XdMES8WV9W/mmoZE/LWuz7AJQXjG9Gv624XE9UobyqZUQSJQAPl
RHG0Uxy2fOsj0UF9hEcih4ZXKdiEAlN1wIMCU1RFCjTB9VLOz6cvV34V/IjKY4dSQnFV5fwT3WZK
xTqoJCSeJjv5l3ZhtZyZIJ/vpPWXmB41WyOqOht3ZmqBlofBrDHNCWUb9SUWfJur3mfkF5oJx/Lj
LVFP3RVlNPIbszIa9GsHsiH7xq+vgid4IzOQWmFAhHpFxlg0NYreJydk83Tav4XaXuiSEjD2cKw2
e5fi40mkN+Nk33S2adTKZ9u1WNS3NlCgS63qr7ssJhgihXGAWsfZAZlZjtkDkQXgu48tnBV7DGFR
uGruCGEAV4uHwD9BAyvo7fk0t+lZrasahab+fY7X/B25dTwjjsShdN2n4VZ8uVvm63ArS9cVqBJT
3xCE3H7+FAyGfvLHYyeZQLoH4FXHbd3nI/OHAIuSbNxz0WS677aqPZfo2ujTeeMtmRS6RYIsVYuf
pTLHNUMn0TAhKjp7P1G4c2yUlMhC7Gi8RHfe6jTOMugrl51YtL8a4uFBMrd0VkNDokk2Ahrjbt3S
g2XGJiwjAUGhN2Q22dNrOZN12xHi9OBVYzSDSGTSiNPlZjJuYR4o6IwSnipjrnWf50cKrhCDIB6x
Jxm2kSmMMTdHy9esvMCcwyNDkUGTAHtsfkjWhD/UR6mzVHOQxOzCuPDqI1VOnNrKZQWc86bA1NCE
VZs+N2WcfWkQc7CFPAeVm8ExrSWq5e/ronAUSLmA9GMajoR4OZfzpyO2eDYAtKj6f+ziYywud/gQ
JpI3znQ2RMMS8lpnhs3O0HQzDv2FSLFc2Qb/zyeyHDsd0NLzYFqxviYMO3oYS4XXZAZcdBUz9M8s
9vpRKsZoqLEp2vk4VwFisvcr8ZXw5HuCFEHiPAugDYuo7DOY+BR/LNVxWf1k2tdxRVeCRsn7Hp75
uDBMlmn+32YbmQxx58N20htzHzMfjmrEM7ykZVAcNoEyAMsgEtoBP09ruNsjBYkKavTehXg/KhWp
Ur818O7/4OLIh2IwRxLrYsmeDHL2wntBZyNutZOS5xwxAjbqKluM1a2ppfsjmILACYHRmshy3pqg
fzXXMml9xVHwzs9/ui69SrSHTlLTVG1hXkr1QCCDXZVAbQ/5oY3stL+og07/W5MSsBFH5yXeUz+V
LL/2mRQLTHQ81YvYTh/4L0cNqYaIwavUC/hIyIifbbFOb+dcQSfwAuk8uTgh8gcVNxgHqSw0hWUr
EQBymm0A6pF3PqkDr5CsNEcDzO3NdGok1HCG8FQ5yjJeFbxAry6uatz8jKVJijo4xai6tN/gNMNQ
EB1Xm8THYp1Bzcs+YE88i/GTJ0kIvGX3g1to50JY/GcekTF2JRKjVo7XxfHpTLYV9Du1UBa75niK
lTy77wmDPJg411UuJc61PnIsmDo501QwHdy1hEr36/+ZYQYkc2uEwuP4RJUCkjWP1jMfS/eXwzSZ
gXagcqYIvZGsfladU3v9TiJGCseTRvRcI65+YXJRjBDPahkKRLTkNP0oGZuY513CSKiNskKXrvac
f038pRwKsFHuWCryZvF93HuGz/qzoUHXYgIKhOfM8mqt4jrmp5Z1fTw4IudAjy2v4yFZQoqNHd2j
COOjyicO7bpMJgz4ttTDPxFYmzopb0SzYnZ2c8K/2sLWnXt2OScqbM6inurETo3PnLLPR3jkUPvT
Ad7oqgO9bYsmhbaMbEHiG3R2/uEpqX/Xgmrm9ve8hATpnWNAbIB5pvLlfmenhDim1+pheEWuX4W8
1oJDQ5A2lzn+/KbZD9fsG7HcM0jywXSfUN22mKdSFwre0WTrEET+UHtlPrcfhQc7tKA1w/3G0FIl
Rf126mvozw2yLaUO+CKDgvow/FPTz/mLoD+3P0yn09CMC7S1+k0J6zJv0Czzmivrt8rHJStBy3z2
FI2FzP7tIMPRQ/ExojlrBYeXXUM2AwANGL5NMQZlwt5Rq2mbhRHVsk8HTeZtw5G1l9lMA8nqX5I0
FiDMpaAgNR9EnPVBmPEQfiKQm83N/wA9DAvBK0ksd4FLyjqS6ZUOokKAx4Y1hOBXDtcFQCzWN0Me
W7ae5N3jovPhW/h13wsF4n7wQ+puSKGsFFUewtH2J06a3uJNs71hN3v5d3UDdZhQfQ2IxHidGTX0
MEmLC66Ks++HpOcfZHNRUyv00GGkov24FrD+RUdF0+COVX7qr7AXk5Hn7sBmJzc6m3ePq98CbGqI
4Cd3k74ok/eUltRoPra8F2KQw7GqpTXyZUNp2BczO89Runjmi78uOXZm6d72cq6YRXfLSwW7vhDy
KOyjn4le2Ar+cSMvAyS6JBM4dBRmXqkD91hh5WjQNh2jDoQZUo86OYnJu1o480C3sdTSNR0lk0ZJ
f5KzNBPjfF1PoJ0h3jCIx1RQqnMCpVzGKwMBn/B0eMqBkj+LIm3G2pMBWRCFEvORa1xQWpsevcs+
5oVI4TWML9OkjzuPzEnX82ZDLOvNXrTUyf0AGMsOFr8vXW32BJxz1x4p2D5z7c/i8pLhCa7NE+wL
10LJePXLioma555F+sTmPbDoQ+8ZAbyjNf5X5XBjsT9Tq4Ia4VIzt66o0Bl9hC1iB7lDqk4tly5Y
H+iowxidLI/Qw9orX9Lt4p2zpAtZl2gh7+Kf1svOCCh5vERYJDjOwUdvbm0Xo2Ny4O1Icz1oko98
CM+Uipc2DUKCzPU5kb3p45ewJx0fW0XUatt0RcXp25H/9RkliCgq/QFLYCbH3etmedGL6kO/uHIz
KGJY7ToLGEJgEzY4MpPmOjBr7kqU2zSzBnWKXtjCMtunVKxM9y6yoDq9G4kbaOAtyITZf6IbeukL
6IBn2kdCeC9pRfzyqO4yh5NxsKrsabiW0o3fAJFUJiOrh7aI4Vf/9Cp9rdCsXexLiXMXzHQ0HR9l
0mbzJT17QJliYF6HSP8geXD33m/RxPM6Vgep5WdufafEq6oGLRiIT/HEftM8luZDCQhBXHQupR1O
w/Zl1H66fKs7sGYAN1Rp4dYnGWjnKf/hkW8nT5eG2vH+iKQj8Zxw9Z/gZbGxoWh6PJuXA/ALUVtl
ZPXKfreQny3Rlmu0CW57d82443ROfwO2i3caSZVO19GIoQdnbuT2cOVgEN9eRJ/m0p6/Z3usNTtB
UDqOspvM4J80DvB8WydJUCeGV0/yU4UaTK3jF8xlok4GEAHddp/OdCPZJ/R6RnKuTUYvQm1HscuK
OdMv62cj9EyyFTsjT0r5nyOBf2TviobSNrYVlZaleO0A0mWy+o1mV53IBAADAEn7g42kSrxgrRVn
Bd+d7euotxgjArPQKr4FXhnkbyOFXp0U/Ohc5qim72FwI78AsES7ZD7LQYiGyFpcWnQwhftQHHla
HDbvGcU3D140k6d7+sIdAm9JoMmjVio8PztwZatIl03f/sQ1WPHfpsTuOtX2OkFJsgxJ8JrL+5hd
KLXORCrjW56C8kocT0PByVnX7Ahk7noY9ryuQak59NkPGc40UobJ55k1Dx7bWjQ4e4DC9Jo1nZhF
7Ev0EDBhulkUWWQ3KyrRSy8EP64F58ihe8YQmMPtLBnlYKvcQ0+Ct+NMhGhgVSQLH9lXVvlIMuBO
loOKXWg9bNdQgZWcb740f7qJoKnU+MNwhwd7750GPwkSWVN//Ls0CPhz46aWb90QgC8VP8DrfqA4
TlnSIxFij1XK+WLHVL8fVAi/6n7GTVKmkxyb+rmFLH+n0xfZ1SnB1lucdgN/KpPrZp+fySAMjINh
2Oj7kzeTx/cJlMMv9Ws0HqfZLEC1pzi3zJaOZr/WBEKfOH1OT521im5YvU7PnHd/K7AzvVSI/r7X
KMMP05en90NE1gWfeFL7AHyFjA2hPjcFt88Z2snKzPDnUUtnBzEnpMrWZSwd+Y4esRGRGJgpV+rT
MCm6JQHbF01QeoF73dXgSUiepICFTp/g/ZvJe+6RR8aDXd0rn/HrHE8PqUtD9h5fBU03vs7rRzAl
7DaIITsB12vhiox6hxY/b0eo0dLOIE2zzwIwrK6HMa//WQXY8enGlwgzG7NFBgdaEN9OtRXaDzYf
m7CeoIF+o47uQwNnnSWXrTIeZVubGhuTAh5553hsnnvyiZYbzGFYweLcHgD2TFvuQIqwTe2xWEoC
cu7rlkPJfpHMXqHTjAOMjMEKWOnBorTiQTJi6VD9XEaDdOwcnJd0OQc8cAFMdXAOpInZ6pgCNZTJ
oo70g7xTH7IaANZrhe8mPODFfxXtPR/wIpwPVtsRuRKuDWEqIndV/lxLnOklSfkvoyHl/V+9QS/u
3PZys4fMAe2NvR37ukbgElFJr7g2ZC2PzZ7AFpkIZURDzyX4wfu4BYQ7z0w8lK0RR4woC+vs3Dbq
4kLvYPJn68Ix4w7TlsFg0a2EVuFBtnMAMQBZIdoX6xOTh5tJDZGSZZ2V5j4RFvJDfwB/+In2uWyw
dOhJ8xLmG3QNvKrGgWYR157CQBf6kygBkP/m+mR3I67IvnEYqKaF+t3oS4f0SVj9j1QEBJ2jsezj
uMSi6otQPs1+xdKLdg0wu0Dav8mxbVvdOnmMeKDWWCS5HsrG1xnQC8k6nN+N3N7ErlAzcopjYfjM
QfwopJBzOeYLa9KX7jbVSEHzaZ0ZQSmNgHxuUtpHh3YBdXFwiaFqaofkLV8y3O3cmn1lOnlrcogS
nqdK6Y+u+b7as0vUbyUHwm9r/X0FoFrX/WvAYpLLe2V+tCV5cUy4cS6IQRwpuKHOcn9OTJ4UDCZz
bVhIW1Gffg1hcugi6dq73dAKorcVn/PFtQDwzL0r3BnFMEbsi/OFF/SlHXqBwwGC+BZGqP5BJR9S
/r8HM0urIYzu3C8QXk6vA6ZhoRbyx17fdz383Fx5mav4/s7EJHVe6RLOggk9PcQ7VaMTqCiUNafx
7DsPMw1qecMe2DJ8Igs/PS6a/6HlHKxM30dJdalAoA2io6z4BWC+ESBqqQetJCtqlghLMA7b/dHe
74cxO2ZgVCcxyIFNtpI9o25ZNzYtLC8JuqrEJtRYJGoRi8drGOvlMSdc9QjN2Fscj1uLsb1+n0/s
+CsnDI48whiOVjYKoIN61wMdMMUSzK8Y+v1Lr6VYORwpEkpEBLy3hmySFwdLZXJunpQvYQutRhMk
ASSIZQZAi0TbekQMPVSPMxcwexJ45KoMkbB2iWu4j0iTYEKGDH+Ed1o394k8ggNXhA0BvWnfXNNS
tpNCWg54mRJlVqM1Xu3PmVTnNcwc7KbMSrR74wgewEe1iju24fkkbHwE/ZtQjW4iRwAubsE0vqhJ
w/sFp52u/8Bi4ck+owlB9EcBzpKzCC0CgXy4qFLUUrRh9NDLiFPpW55m8jW9K7JfpiVHAWBLaRZP
F3E1Vb45C/R2o5MfY5h5XqKaOXgN8Z29l4hUK3TT+f7RE8aMOVZoa69smjacPp53fa+3EEP/WD83
xCXuF6yoJxsz8RSC3yN+7bF5Zwi4QxQVgu5HWrUDEiWHqEGIqpJmPyogj+bXzQoEFgCdL1polY5r
10TCAIZXeMeS2Gkfd7wfae7q6VzpjWp1skdBrJHGgA9Rhdxg3wM6Wol5+HqDiAQ2UFt+TxJzdjYr
+BMgv7dAIINkw01aTXpDYvCjncRG2cMTZu79azW8/TZrgzpz2nwP28xHcilDf0ezi+bYgc2WoOH+
5xjZP8rJ1VFElApey3kqqjf8nNttJbmTEareGcMn6Poi+sG61cb+t80pSMk7vQBXdS/NqVo1tVkp
pBlFLqZ7B7WreyOTnm9HT8oynP5PkR7E9xhPxnbXjzgJio7lsQLX7ikYhon8MjPNC0fUWtPHCocH
sKKG8YENdHtbUtuHg4wYGZMzXDpP+tehLUy8EBtVBnW6zdaa6NeMNuro3zxtYb2MiZ91Sk/t8Gqn
t4joNieuHIKafzKuBS0uN3gF/zoXtUx95o01+tKCIEH+detQatl+ekiT2zJu5WUwwjdzwiN1ZQsw
xVM9MRIdgYrHUYC8r9TGz7d1LC7z6vN+rM08jXfu+iUi2MfQXINEPN53QKrar+4sEcbeH1lK3t0S
sZhUf56SSLPI50POQ4qN5riIlnsR1UAcqiCEr0pd0YgEmS9QW63BEKm8AG6qhJgqM9uSanayhz9g
N+TNcCb7qf9kN8uLWXwBCCOkPzzUK8pUGwr+FYZ8K1RgtceOa9gxseO0+981pYvX8Cs5D/lA5Z3P
Qg+JBz6I3OLnzn7zrZwYwJr+dCt8f+gn7cBNMJP7psmbRSZys3BFEvYpygyGDWscP2TNaZ+NIqJw
ufJdFk6yY5QPkzT447FQuEEBJMIXg/NTWPIF+MeNP08HknDAfUnU05jJiTkNY05j6gCSzVXE5mUR
Q2NZDzZtfnU09FLDuG1fQl46LdV3NGKFPZ/E/Wm6PhjKYeWBBs+Rth+jMOV6anv5fJub4/ellhnF
vUU0C7RN0e3t3NQ7AOrA+MQ3ed/+TWQuSfB1R/e7EYTydvJLwauCjlIZ7vTl0tEUfIXwgXYol6Fa
GEwdbXGW45CRTAkRoyudOCy9trKzO49P37eYG4I+TUCDepiE4wUHruHRJhOWxy4iOIFeaimMC6eG
n/eeVvXXRLh0iI6U6b98bCVUSn7/ZtORVlTOr/VW1bXnxaEwe3tJB8kq2TnsVk6Yjt+geXM1Osfr
Gm2G6YIgB+sW8ZSCQBhYa5b0/i2pQTJub5IP8ecv8SvLhpV8VrAdebIUi6r04kKELxAaVSq5bSAZ
pzQjuNeGUEpUnC/1VsadIJ5CmH0LkO3qshcO8enpSDalUqsWggTVYtc2kgy9FX8CebaGb6Wvumo9
vgfFLLzQFzzMdVKaqNkXTiDS6jRn+A+vUweACw7Yit7M7rqt+AkPFC0zBIvDVpTflqwaoe24+CRV
x0ZxsKFqqGQRUuhfgMopOeJN9WSQP0SkAPkgiCfUROexYTJGj2IfnHmZpcBBzOxYcnqOJNhnHow9
B87V79Q6e9G19z6JuHwN4pBKIUi+o63yuWu5vEIuoXmLc81eKxJcaveL28gJ7jLiL/Uu6uk4Or3L
If0C1DIGUv+USvuxOzeCNrN0rN8cr0dg7sivFrLwpgKXUWnqyztrUHZc5IZgHVEg6Npmu/Epco87
l2uyYp8H9cZXO4K4rbLC19/o0/aTwDwPbYUw/ftgGMlt0M3DQ5RXufuxmPJCf9vL2pyI/r+837lG
988PEoW2lF89nIJoImh8EqCcpTe0US0kmbW6hSJ+ws9fhIBboMuWloy88+jU/mB9h+cS+UzXAKWF
yVikLTYSFzOFf28pnZQi5m+rbLP+KrBCynnhl3fK0i2SPWJnj+WJqCDiJ1118zf2KllblksHreeM
zFNvTsOi4A35OEnt055h13Hr8Xotj6c3/PfVOpXezSAGGmMWxGc5ekeXtyh3URLPldAa3pImKwo3
YY8U8omKVV9w5R0LWXX1sOUEoseqc+EDyrd62Lyq2JQr8rMJtEo1baxmaJi7VbZKBH6djQqYbASW
WpWcfadsb/QGKkx/RQr+N9EKXeWlxbHFIRUq70tNVcmuTCp56XpLAytg/WUdhVZjWgha5nu4EWDh
Ka+GF9K3VGd8jik81RzTURV2Abf10wvtRemZwjhpKd4rikF59q+Z0f+D2RbrxVhJPBhCre3J8prB
u0X2c8b5F5BPnHLwvT3DNfRhfbkgB2q5SY0LqadHbsi6HrJD1ReRcUmINDiH3peRGjJ9IyoBXEYl
pkj8HMACIN/WSnD2RYM6NCXKcyHMcf3Ffrsm3c5xAhUo7/WqpWPPZCujYmRc9EYvgNjoQbB80BgB
OaiQUw/cUampUoZWsO2inTdtg3QPIz2dfjXIUWhA1oC1GxTqqBdZldoKHtOkVqrNaH6vIU768txF
uqSs6cavKIqejyulpZhJKucPdLxAjLvqRHWVQtYCi5da7AuH2WH9V9rOpe4Iw7i3PX6v4qnqMK68
TxpD4c2BVMD4Wk2eD94C78m3+Qm+4X0l4iykSMX8ESNJRztH5GpS51xw7axR4qbMMMsvHD51fCGy
o7otoheY6E4geT2hTM5IQjSth4vOwV0XExbaOhiUor7RAyhRvUZhuIpJnfuHn4G7AEx/5P/4x5fW
9Z/Xqtfd7Mg2dBvSqb6+G+VwJQWMGMJN5do96YwlXJxE5XfAODKmwckOx2rYxH0nIEBsUelCz860
o5C8OuHIeK5z0RY9UtjHaMF2FC4EAhosxfd1ernE0oUKd/8pLAnSmSykV7igrEBXFFpZXDLRYqkr
+XxbvDKhG+04Nl9oHPRZtXnZyDpQDC1J/pvSH9ZTbfqXmJvnvQjuZycvzDhi+HTAl6IePepVbM7U
9cyEdv769ePN0S68WqHEek+MR3097JsnMdKuGXFnvhfmN3SIEViPpUZzsAjStt4d+RFPwa8p1FO+
GgPidYjvqlY5JxaTu1XaRY9ZslpaRbOKDsFvmmXXIBz1r/Kseqy/hzpsQRWQaif+CnSov9vtd+Jc
g6ksJTm9aqYWuzhWyTj3FGz3Pbo6QDYxrHnT+SFrtUEe+HAGGXo32t0dA7E/OgoHsDad3SOxhTaN
2vuHh2AdvioFQT1WHf3r9iJR19DtGAkJtAmsjoQbsQpraIzMkDrkkaRqz9TZiF/sKA8/DPKRJ8m3
VgxxUl9GlAjnEz9iS3nSqnYRMu/OBqs4P6R4jzXFotqwXJ1ZV8SG2sgbfbCw+TWKZuJxP5JKYbTp
fNjqiM0cdazVRWIZZ7ptFSUARmTl2Ni3HYfSKFkhPQ0XRdxRx9gVPsrTMTCwLRTTMVz+PREJMUpB
o6O748QpTkT7s/NCCdtDp4ab2ZlFFgnTIarVIOJ4E1E6BXlghMTZiFzXzC1JXOO2k1YLI+M0Q74t
iWs5C5hZ6zzBYgGHp3JjYJJXK3afMz3jbCozn4IMUX4h0rM5JGOhzw0mwJqoWT1dn1fte/KQG6ik
gYNmH15QPDjByWh2oGygUQW0CIgjtrmL+0OLqjGcvlBhdDp5L9/XuAAxa4ry/+GrPWEA7vRm7EM7
iGTyKlbNv01ppqbFK38AJxuERkzDUB2znXqlqpLc83tkdgZi4INY7WZ9gB+O6hJU2Sd38VUZ9DWs
EiI0ykbNZ8Rvetxs2950BK4+XXW4hDIfGWwJofyzA0QGERTTlnCpKbK1u07rfULKmOWtCVFm/NC4
FwnYQrNaY1MEkDJkQmiMxduUnFKWL7EzFv0YUwLjfHsaOxFqoK0KOWszJndoZxaDJKKoUSTw7UqN
HtjFtbcOfollUUFPkHNz0xZ/qjAtycEe/gPTtlR9tFBNgsd+6Sa1mARtU+ERi1hp0VqGMvoYwl3t
IdD5SnXVVTHoDhxJgOwq5wWDNLUjJO4a9z3CyW24VTNrzU9V0GmpnM7n/oP0sBDsaMEz2XZB3T/F
YHsNe4FFko991XUPxBm+/6O7z7c2VxD/02QrLzu8KKLOKpXMed8vaR3+kDOR9lkddpVDl7JLpmDq
gwp3QXx0LupXLLmF9swPFi/OQ6z+d+1Upv9D1qi859fH2+Z7GmN7iz44i8y4I0279EsVX61ZwD8f
M6LrvVXGEaIbguYnO4xdkYxUk3ZjxYuE8Y3kpYvGejdTfCQUpWHZ8LszDbTtzOYyjOzsSu4seeT/
Yo8coFej7oYeBXA5Gdj0T9NdOZTUacwH6SiJPVSfC7h1wvR/e9JjkN1ua9y1WUeZrPxsRclYfoUT
F0On4RKip2ZLlXdh0WnUfaqW1afH6xosgjcgLgOTt85Mg5kUw+ocyjoVRojvTdeXAcxgAkLPKaST
gJnbeYCgo26OE5EuoLfGV3wZM72LRQDKTcMnlKmJ2Z/tf5Js/dOH/SBFwipa4yQSmilhOJojDPso
RlXXwiOeoO7dc9gBvRSwkO1Ta3djYmIlHbIRRAvQ52gurXmsiAcU/FZYOEh69n97DZpXu9dsi/gO
n3MX5CwMLS0acwsOmTVLL2F5Nt4SYgsVOeQbhwpeUpN/dbC6cNusRCx8/D4yDh67Y+YGolDYcY+d
g63BNuu2yiHPV+AfeY25gjTiZFRy6nbhxnigXHbbchB6l2AaAGY5OXildu+UtfUkNpab6Y7aYgdH
I4P+vNrj7WJEqPVkNr/ZCW7BxQ9FTsudmLak2y6xNCmhtPCJkoM+sncGU37/chdVAHsXdrf0Yp0v
BVO+GOJGqT55dPLFlCSaX1U0kpitl6hlLp//iDa0G5lWRnP1VeYdf08Ry6AjG9EqUviGD+6YDYYo
Iht2k9WUb81GRNPpUHbcg8F2PbiOaUbexwKK18JbCgJjt0MOM8X5qt4PmbguoUT0Mmtcp7D7w6Fi
AREGc4xzKGRbOLzZyOyXk2hm5z8s0w2Gcu7qsXoCa0DY0T+TfKIrK8GaE84pGN5QFabmEHluQfHi
A8sK8iFNQGqRv22yaUMv/3p4DwJaw+CMDPbnatmlhMeTqH9igsJKt0E8mmLiJJenDGo/36mNoNsf
q1gXHqeqtz7tt5K6JC75vQRBif/Sx3n6s0Jz/uM/V5Ru8j1BWr6rQoazALHI6sthRbWlIbO/8rRS
oa4wC4MRUzBKh83ujffcJu7r9fEBgC7nUqiEqJJ4LEi0ahpd+wXLULHQooTvdseb1I5qzPC4d9lW
Y1LgwYnrU/tPmInAOWrNIg+dDnCTZ8ZkqwmMpCr1vY39vm6HBmfYDE4Z/wlyK8+zSR8lzRtPcN8g
HxcWCyJpEIxIDuwK3B3Eqe/dKRyd/uXhCbTExUJPoGziMuPT+Dtg6iDzV2BpUrp9qaa5kyrm6t+a
inLSsdEMrAR1GkJIVrn33N4Rmu4EDW6J6ypBPqO9ssvS6vbR3Qe3PVbqf5oSTz42kZmPvQkF18bt
rpQOuX4/h8qoSeoI9VYC/MTMsH7ZQrptmzBTVTkO9DDkuoTYfS8/WTMoGCy1XgdakB7GMnfDl3Jl
IVEx7sb+1PvTRjsvX5Px8PBn5tZgD2wGWwEkzIjy/OIQkUoS72uncqVz7b/UsjeDe0bt+FVlZg2m
xtNKMJ499ZKQUAchPszKuwlKHqxlVTgPe0nBqmP5qcrh3Ld4m8ZwAp/d4pkqc6OL3jiio8DCuuy7
/nyf53vks7JmdvjS6C/QxQa4n2mJgvNepT5r1PYBfL7T66CPD9pBi0dPHpcMtI7elOT3GrhWfntq
rg9zVOmHPLpGGk0vV3ZYpoBzMPOeFhkF7RbOIsmfHoynSt3bnOIe2+PY2bHDAo6JJdOMiUqJg8PM
ZEgKa54RmvsC2R7PdrO+dZ2r/dTzIj+7oHF5szIH2JSh8Ui+nVQ0Fa57sScXZSwNfJK28/daIj/L
5PqR+vvPmp207tg98T5Scv+xgpkQc6/WBXbhtTYao1/xgMc5Eq+C7tqCSpMPcbYo2Tv+nqZGkHAU
X7sYZ7lhVG24GK4lbhvpvyCRliU52qjPt3ABQf53tn79NIhutgT9v/j4P62r217zgE1SKmSACaQg
OAMI1CbxnM9mAGuTQLQFjgP4ec/Jk6HGhicodBg6bypWTV1DqA/kT/WC2tHAo1/VKU8RYr5hGTlH
P6qHrVSrqgdFoE6yIB035yDWhQ/N/wE65qc5U79dizyijdgMHMO70l/YPFH8pYPU61xCoQwJUAZu
iDLKg5AdFrTpuCc9jNMn6WLkeIhHUZyYTlWRLucfw6A38eHtOvIf69EH7MS1Jg9Bb/5YkFIPSX6X
WOBbltyW2FWqeUlwzrvAiohRcXCuZFconRxtgmyY1mhhUKdoSmwKFVuTz1uWwTQhqB5atAtsha9p
2j5DIZ4RJSohVIUW4pxD3OTanJIn7ffNLlbA93Wcc3alTvJwv/7/RdSMF+739wIcm8ODol856FgE
fKWq73FM9smFADDtv4B5vGxGTc8Z/TNbCQ+5lu2Vkb3NxVHOMGog/fZTBMBVlSv7pa+Qf/enusqZ
Hs2W7qN5fjIn3llTlZFQcofGdu+UizGitCbwAixHUAQkGqRScIU2edcW7Ggqx4R0ZO6SPsFhbg9x
JdwUrZyG21fhwTXnkWVvptsmdJ5Vm3osvNHHMFRoOqpTiSkEXW2nTHwjGqcg9v/uHcg1goIGAuaO
aHffFIBGhaay7JrC8edbalQOcfRpluMA3wmJV52pfupyimGsmxv/Jh0LzYIhXgGfeW2DcrKwsTL8
Rpt49fNc1NjTxVYvemhwbavV+C8iCEr9bhfDeG5LfAi7lfCMWRqvRIB5t1zRRvbbf3FfET0K8QND
nVlnCQSXgNbilFGXvAogiBSbzTOCa6aKXupN0bI0Zb6lpF0A5M+ofrts5UluKFueJD2ASifsoW2s
TPzEufeoKaMFxUC2lgacCHo3aikRX3yrKhLzyudeUUMo3A4lKZ45U1UrC+Y6psBP4LzD19hqUSLP
f/ZZ57VeMPiE2d5XtJHGOPUQoDkkbFwkSZ0YxdVQRzg4IZ5eeLraPC0y31HBvaimLMf3lZPy5tWr
NK/9i6IFebURVeYkKkI3s4t8FNevl3fuLDg1hTFBv6t3My2wV5Qhz7O3CdQ7v9J9e5NQeuEg5GFo
cVbvrI1c2kX6SXf1hlV8cW6FqPDces0mDOrDHx9a8c1IjmGs2PR/Xlu/9vRw3pjYHchSc6Igk215
I9yI1RpIsFTTEqNzsUkM4v2bgHQYR5jkRwQbv+4MIIsB1nviXi/LJ59QB7PB6PTDjDa8sFdjoem4
9aF3hexzmm3MJ/aynsK+NrsPC9Ldw+DjvtuzY1Ccvp6tj2CHxMCqj2NRDdM8MuiFZ0rI38UKk4cU
lsSM4tQTOYT1nUYIVK6hln4Og2GuWR7RYK0DmkYowq/U8aY0q8auHGUHYAmzgJhXbT4dFKklGkr2
ADhAYTKVMkP2+QT0ckDm7bWELvn7P0OfMneLAQDeGIqfciXS23ekXg9vZcUI7dz1lcDDZRT1fqub
EPmOH1wyZtfd86Fl/qER376uCWEavhVp2/Kt/RnEP7M1sH+kAaKRVLxAhbjgrvbOChZNhNtydhom
Gnp6XRNSVxSIiC+WiT7pq/wxga+4WjaeIVgUwd4YjlJCCBXVKVWKSEK50Dhkie+mDGkyk6Cld3M+
V+qWsZ2oX7aW5OpnVI815DVlsbUkDTKgFklixPb5+bbObIZTLV17xeDtp6ZHFrOO+mKyGibCyxwu
OEqmUMBL0AzHNOxVhRo8nJqY1omNX9ny3KeBwF+SsdBYGfj8tkxEAuJ7ackJSBPiaGfKWXnAzlf/
Dfax4NdALDR/K51EZUYmQM0EVipcu+x78PmrJGYG42equ1uL//jFjQB8d71pAGDHfHSEsx+6KnIC
dJj8hn1Xiysfsg0twhP86QYYqzRZpJYfKztw1981TRU3n6WGv5zsQa6y4sWo8L10LTopgDbyR7mt
HZ8rmHZMQRNapCfDCaY659EstkeWEulyDAKC5o9gRuFHMwScAnT4X0NJ5sf30tUFWo9/KgDxJvmc
vER4TFNkR//vhw3qdeJOrLWUmisvUsvKZ35nRrMub/FYEFtZCzeByhcgYkVp5MDKL+FWIeLX21nw
B6dLKvHFiotcViPA4dp6+r7KrHIK2OLD1Mdi57686wm1piYD8D5HsIbuDup2iET+QiuJ7bOj65f7
oxm14Lp+YZJnVLwqG5U/ez++HpXXgPvYoWxCRRYSQPX4+XTghLpxa6IOYm5dhtzyguMuiDALtLwG
uNvVfiBCRU4Dj58PICkMJBWWGVALdcJumP1k/sgBBBkTzyKRN9hKwPI/DlyUEwvjwFS/+3HS1zNJ
3/OL+SFqXO5FC4LEW1FleA7dIEXQpc4wghQWaNd4x37gWYz65PVnL9k4cY8QtXq7MSQBjMxWJmKl
qAqUU25VJsHN5mAqXuqTWVt7k8gqLMtmgTiC4THFSW4ME0h5AsWIDbWqmPqS1VE68LZjvpAmlOqn
thMMeZVENfoF2AHkxkngEjSIRKHAuquWiZxqlOGnpGKMNz+ofQK16H8ygIC0tWSq4CCDuXu8+DNk
uy6J2jbxt2qg2WRuYyGmC2pdq8c34iBbQS0Jc9YCTsBHpsc589p147HQ412bpPNn+N1Rar45fF8q
KRDq4jd95nre5Pg2J2kWHqVf5SqEdqZ48MGJfEU6/XUKcfLTb1rIZ68CPzuG468DYrKJZ9D8vaS7
SPx6SGK6fIGUCmeKfo7nbXgEKDg9pNMF4mr/TwMr2YXlPYvc6oQBI54AUbY2Qogl0c9gY1oAeRBq
GSbQdaQjgRecZEW/RNykpLLW5WQSDMKOwbq2aO7P9BuE618l9UBLH5U5G8xL/K1w1x8OJhkAl/2n
M4rcVCy5ShnD5Rjc7Bu47XvyC38f7GoXBZxaUEQMbN6Mf2nq0us1g3fXrS2ESBBSMfNZQiXnKPL+
JzcHsxj1GXVITkX2w2tBSh2rPYENVM7CympdUgB6ycS2hdBqLlX/EVHfqd+MvRlKyIukmvIJKvb3
9OzHEvLzoKvzrC+0/L/oiFCL8ReTIGYhRXN+oPCU0H0JeDNYTiJ5sr6WOMa+FV1qmbfDnN20qNDL
Iu1F85OW2lyyVjPI80JQivUPwLIZAVG/lYi9+o4mnh/v1Bdi6IxKmbPsvDnln+pInN6w+OQ95BL3
vrnPQbSaSjLpaUuQb+n0giEDlRhJCmYbSgpOraIQqiJm08x3A0DTpHkW/1HV9YAZTXirB55px4g2
M8laeu2I/kjdQKu3FFcMRG4u6HPfk6mcziC5r29QGCOyBuLplpi/JGZZJaOLlI7A4QsHv2CXdXmp
6vgAj/J3klpdlB882EsEXwUaRVJsAaolL5YZr0+yv3UqE+m2xsTNhqPGW3lIV1orYIrNGyReJEj9
1f+1JF5fNrWwI1OZf7IgO5OU15jfsfcPqHrtzEe0vmvLaLS6/Y8XRUL3luF+62QbxDRWrizb2CO0
j6qmvB+O7PCxsw53j3Rt1wTTdh++0rvLhnnicXrWqLml/dyqTFdq5nCCtAOMmMIoOVSeBMB+P/zp
yHK8IUtaq3kcetGv2HjlmbJiXcSreicIi4TLpuUF3wcHYUBZs/1dryS42cf0W+pSdKMrNmiPWmx/
MIpV6yBWi9PbdkkSuyS4/yKX8FVH0FIUS46jDLs4Ym4FISzN4EO18xy+he3HW4kUanycNDpFTPNB
d8CdiGeSauN4NL72gcmebUcKHTW2Y5sMtzdAGJmOZbYl/1QRORYexEDK7a+4f0Q39z7VdtvL3qwY
84NLEoILBQQG5QM/jbEX12sjrhop//IuChIkS0Hzj0oGHVsKsQeqKcMYyVNUK2QxndNWpwCp+4L0
cKtVFe3QA8L30t9n+769n4j4WJ/rCQ9H0kYlN/crCyopS2jBPS0i7UrsMfaMWb72uNO+c9yscaWw
Q12vFN3TUdfSjEE3X/YVn5sxQJcWSoZOIfUfcxaiCaADHNVPITeYlPVyZDz6rbWdaujSOLwOozoW
4S8cBjA0wIDzeKCkuM10ZeFKIqPriuvSBneh1sxtBWo2EbQqj5OfEf7jR64RBSTnxHW9ZHZX6jsi
923hIxoLnSrabRm6pQ3C3BFsxQyX4qHkSY0qAwXlGstw/xx93lIkasJ0zh/sFQTl3PoE81Z4e7ev
2F1m2LSPSPBBxBbM5E/pJR8r6ZMh0mu6T6DxJr3b1q9kdfib1FYgeONkgmBoI1MsdvDIXrBBRtKp
I27w6jmOUe2YloN0TGmLBNsfllupBeOTaMsvbHlCdFZs8f95OsO8lfCq2hWD+H5GVzSBraiam6kc
8OQjz//Hc0BAgc3C2fS6xcQDwFVJs42OiQgXRnHVBc0EXACoOwmkmu+sel6k6v6peHlVW1iKEhFF
e+/B8PVZ8cJDUqiXw2K1mH8Fh6XTeh61dW8IjClphDaEy6M7vsqRMRZtn/HfQPQwKEjjccKYy9cp
FADXth0eftYckSK6oTb1j7AN+CBKti8nQtAVgWZ8THBiaJCzfHhvRy9Bv2aSW6D8MxmJRGxMw/T9
5rN7jytJn1y2RtaiivEdZ3/7/ZTnKmuOa0sdXFcj3lQFDlQ6VMSTGdQbC7UN7FKTyh1Jhl+sNxfm
7tehDh2NZYBdw+uNcggf/r3/IcMgc/JgvKcrEjkZORymj2F1vo9yGnpFxsoXHPpKnE1YDyRNFQv3
ONJfOEmOPyBXjIWnZZ7O/rThLzY8UNAqIXu5eFZbfsG+etBg0nOaRMl8Fp8rzpKT5iMEoAau7xzJ
IZ5GF5IDVJytR/MPHnh9Iq1czyvLYRy/SPCCRXi7mnEyYYbAuSalgFM6p5THi6vnPxDHaMwyZeEZ
/TAcX/OWmrXDxVFJ+ONcDZCAU0TWEYDu4vcLrtER6Ut5h+TGuWly0vaERPjIVgLfI3OBoVmZkHjl
r14HnZHFan7ZaDf3lCmr0a5EgjMK9/TOCtsGux/keA1H9kPnTNIIV137kAfeQSLhekQsGnpMSA6Z
BsnQ9R9ICmKtLn/BAfxm/UZ8gUD8CGcX0La0uu8g0G7Dt3wKRghrayJoC9LIMldDBkWlRLYb81xd
AQQTZ4D3c1ijU9kTPlcbUf9+vGDyjCGgU0uxXhQO9QgrH1cnJJ6YGxPJ/Ehj7veTAnsZFruBPGXI
nCbhjWqNBx+2fXxBg/BxU/D57N/fye2OUxEVoA5PiF/R/ly/MSLh7qYC9TxDk7HgMc6ctIiQqlHH
ni4kawlMYLzsKYQl3dwKsROn+9DQDhUeIM65jbUZz9e+fVwWKE/vFaqKulS3MSDcIQMcp/rlO4pD
oYrur0IZk9XrO6REzjMgDRWOMrKz264vZImTC21rTjoEP/br5V22ML7sznUDf/OuJCvgTTlYA9DW
7bAB2x7v0sZNbsEVRfTP367C5okY/eGN2Czl+nwEHaAhLqlMXpPcvSeBmMP7JLfJOTDnfupkGgjB
9vdyvBqYk1bT++c/BynslR2uJacLpHyCLBj9WGnv/EdrlUR+TSeATtAyn5nxBBelD17daoT7vHMq
bjw0noqHPw1fYtwC4qiELAY/f47zac7atVODZzgjDLdZL0TnUanfCxchk1qahx/G24e9ry1vvNAy
Q7G39Q0Lt6ZMmgx9XGY4HuEsCtycrcrHE6oQYpg/ypyAKYpgqoSPvuPP0RIYplUeA8aZwv5WmlJb
hW0oaLLQRyKj5bJNvgo2T+dCK2BtwY0HSPNQshegrp6cUDuYae3qdg0Q9ET5EPlsUEjkRzAZRzLs
TYBnsBqgi3gj1ELgDKgyDX99HDkRn+cBAKA6c+GM1KvUHjJfemfhnBON3uwBfFIWrsX7AifaGpdK
p3UwMInFv0qZKNKmm7h2oWQIjprF8B5IGrnZzmwWEREx0XTdBpEHWo5C60eKCq3yiTv10BREad8O
e72kaS9B2q2MhmWnwjmLqY/UjF3Cr7JWbOJWA2ANVZ4HxYDCzAmhKM0VUDDhsNRfgyi9fhoz23yE
+MP26KimdixAH5vW/xLq+xqko0764KhzyFihnB4qbQ7isHIA4DwINUchytr20t/j77I5prjISowa
cm3LJf/GkYf0ZMsbsqSoWoo1toQiwehUMBuiNc3lcY4KjkDRTmW7ZysQk5bTR8zvPOo+Yy6whyuC
f00ey8kOPev/4hncKjnIx/VmXMA7I3iDuROAfZ+AekoEVMqpFG3Hs9O/obesuvRqHtA9f/qGo8S3
mvyc7djjMIvmZ6j0tPvKhuwYZM8a+5kOrA1txO01IJMAo23IB2rDn1HEzb0mVBWOJ/7mCHwp3r+L
oATI6S1Lw88sMA5+TH99GIWph2zdDusIGonBBGX13v6GRi/Fu2Tn+7GUN/Z7C6AfrHdaT1PV/ZKD
yztcFob/tFL+xT0JgPX1AwIpEw8hwSDN494vB9wo8dT6Gm58mrPyP/zpi4eevpVCRLFmQVtKImyp
iXUtprDT5ffNjnJaQEw6ti7HJcOO0nRnHTPFuItqplqzB7c2aiFhdUnQFkkx0kK83vZmK6fJnH6p
5ONMwv8va3VmvjEeO/isFe2F2kIyPRP7xX6RKbCo0b+8HXZ/IwPnGcauf/qftyxxlVFE/14oWiBe
21UEE+eoJwCmBOO6I2WPM6SoZO7lnQ4/PokAOzO5XU2+IVK78AaFhlLCBPtfNNcjpoWQwEUEag6O
gVcKzVHBrD68dv94RiY8JqRcn4ZizVpJAHMDQRCdots6XvxZyVyiKYLW2OLgXstTf1QYNkt/Jr7Z
itl1jyX+iFSuc5symdfUJVwo2Mu0vMq41CT69XKUvh2iEzfJPYDDPjxBUu+uMk2qkAtP5+YG2P2M
+pY8ASzrDuPN5p70a58ZSjJyD/duODTYEvbv6FBA7ZYlBNrUR4FxXTcdeOZxbMAWokc5HhiyHtMv
PRVYw4elf6rCYJ+2wDV6gjtW48ExVOl93xLvdqE8k81gk+ubZmHy72BJ6xIsWJdBX5um1hSuXg+/
ICkK58mabqhck5TjAqdpbwgo9j4TMSxkgTCMjQoFzsAm+M6g/aA6Rx/XGDErAZQSgtU/OGP0z+Fb
0KkRIUP9JIm+WZ522GHRBSSKuMO2LHPGiVkKSkk=
`protect end_protected
