��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*~�)���>w�f�Su����cϑt�ڪ�,t4�E���Ry=�i��f��KNE}�z|h�GH�-����ae�Z)���-�ob��\ * �Z�%P�g wnLF;-ACmA�/6���3��d:�Έ�jo�(��Yu.5j�VT�0�"}�����.+���<R���>��m�����}�W��o Vg�ܯ �i{��3�"��W�uS��%���]�a��Q�;�\�\�*����c����Of��� ��`&�E� �3F�t[�]�<�Q�ڮn�qj$K�G����ߦ$M�ݬڜ�:�j��V��O��#�)�	UGD�}ӿ�s���ϕ��y_��$9]����~G�R����
x�[F�C9g�����"1�d�/�a��C���� t��"������pb�6�͏�J�]0�<E��Y��	@&Bm2-P�x��O���:�ظ�g�a���	^�	+�U�E�,YX�p2 �HXPƖ2�P�;?8z]�.9���q��*�p��b��
q0<o�!C�9L�c���T�,N�����]E��/�l�1+F'���̭5J���1�����~����⵶�Ӏ�����ґ(b��(j�N�[ӉW��Y�2��Ģ�#�0�'޾��:چ�h�o�6	�iNg���%�Y�[�<��U i��<��2���)e&.�t�
�L͋;�jvnR�{�_;�)g0= 6k��K��)��h��]<Ai;2o�H�v4�7o�"�p�!h�SO�z�ح�Ǻ�Kw����˽"L!��	���k�=±%�Զ�`�#��`�ʾ�$���v��I�FY��F�E2�ZKlʵ���`˕"}hA a��)��')Ss���	��fۃĔ� ��I��\�e�3g񓨷��WR�y+���ybv�7o�v�h)+:��Pb(�2��_e�H�`�J��8.�|�Ui��&�"�"��{f��X*j,��a�� ����oKz����J�Phik�L��v�� R�6�'������ܽH�����m皣c;J�OS��N8�s~;&�$ �D�R��Iˆ�傓��,�p���j�9��t��_��3��iJc��%1����]\y�Ds�>�QK@4�}�YD?&�@���h	�qy�����&菋P�	�!26~��{:���G�����?B��g�`h�h�s$"�a��[U�CQ�$)Ȋ��53����g*Rn�-P�j�I`�kr�f�˱���ė�٪�����FMX������v@��	J���H�nu9E�!�9��3zj�\lWky�B�J�6�y`m	`�YD���ה7UV�E��~�n����g�~�z�Z��5;�D|ʯ�ݑ��Q�CǪ>~�.����/9�	��M�z.�E@������:���!BaC\r ��*�S�1�h��Կ�jj�.t)[��;>]�(/�_W�0{a����h������� ����JZI?��>oJE^���)�}����=��!�\͢�:ţ�]M�:gl;E�n�"�٭�}W�O�a|����==ͩ:c�uj��^���e@^�"a.}�##�W�6���.��'7�P���f��̂3`=��#�Cu���<c���j�-<�)I�>c2�" �6�B�-�,y �k}/uy����n�g<�sB��db9�ɘ��&��+�ҭ����̯F]�Y1H�!������
�$�<?+.4$� �$֩#��.�g�B���)y�,w78�/T���X�Bٞd�^��(f��e���M�1�3ǭ�N=��r��M(I�S?B�:�&��_L�W�.��枰=ŵ`�*����8_,������b�Ȱ�t$1��z�����I��[��tYF��K�����2�X:d�,#��c���mZ������<��l�-�H��!�Ƴ�@�a>��aцzl:�<�$�������T���Y�Y	C�H<�+�kh���/c��b���<%�!�>ۿi�#=L�~�h�Ȳ��3�S�,a��,Ԡ��@˰P6>���N��Q��Sv�����],+�O+�~�8D�6]>_8��byTX�����@{���(�ګ�M}n�Լ
_�D׼۳��8�Z������_'�~��h���?�K�w��*�o��㴃$����	n1�s$�w�Wd�g���ե4_V����';����E-Lv�����q��0��y7W���vs朰��I9��=q�Ԁ��2��a�<�t_�t�}�_�.Sϝ�	z�z7Iz.���A>(n
��.��T�R�m�e�����^gb�n>#�x���L�����h���P��v�g �+����N(����8
׋;z�/���g[��sl'�����V,�o�<�.l����D�O�%������BX�+�1�|�=X�9��u��Xd�"O���&A!X�^J�,K�1Y�T������0�5�a�7{��`����!�����j	j|�Ufu0��Y��4Lc��[�$�.]X�~���l:�$_�q9�����*`^׽d�-�+ġ��
r�L�M(U�\����5w�u��jTcw{����a��M+iZ2_$�/ׇ��3�JT�,��߂0a���@�2�#��~�gf��n�®6B�3|�}��&�y2����a:g8.s�dT��m@���e� ��/V&�߶&'��Ǡ&�b�������o��5-���C9� ��H;�Fw)��m�8�,s�O���}2���m�Pх�<�U8OY)>P0�a��%۔����_(|���u�ED��g�����}V%�1�G�&���ډ��	RO����U�ׅ<�;M���y����vqiX;>�+dY�},}Sg��)����݉4R�/vm�dP}����$���,��k�Q�"����/Ae�S2t|RD�ւeƐ�C=�&���k�_���������a����N??,j������:/u��p�(V%� �̂�~�JL�u:��;T�\�U�m�&��)� v�9����9�����UƑ�mG=X����p�V��R��1�" o�������`�,�-��k��mF�h�U!�I��n�H��(��~`�&����>��	�5���p�!�c(AʅNl4��q�?YN�ؗ�jA8�~1L�	`��(��t��wl]��8�q�L�F�D�װ��d�9�P�X��u�(�K��5>��u��ktZ��d����V1�����/��I�mI��S��x��5t��yx6�/�{Z��8�c�߽)��Df�`�A���:RAw�|��d�,q	9������	P`�ZuI�>8R�t�����S�{`+B[E(~��,"E-�����>f��L�x�Q����`5�%w�їeH�b��)`���{�lS,�24V��,�Y�1��p�ƛ�����ʕ/���%_5�wyG��>�t.�`%���o�����M��&��ȱ���ÎA�Hw�t��2�Q=��C� m'&�'�8Df��>��*t4�~uA�*q�L���Uz�gQ
!8��eZ��C��g�_�k��S��o'� *F�����m��D�e�i�Lv���|�L�V{ݶ�Fڒ����5���i趞k���u���!'��x|m d<'8G޿r�ۀ;3r}�_�ם��L�7�G�ͧj1�ғ����b��ⅺqU�*��]�d/x���K	M��� ����bD�uؚMq�f?�?�WV��+�f,��%�,�H��C����'=�KWk��\�<�e*%,��z1J�y�9�Y��.^�L�i^|8�1�cc��۾�Z�h���5n�O�`D��Pia_�~��/�R�g�����R}��D|�ts�%����"9�O�!��ر�0�#�1�2o��ǡ��C�g���� �:��T�T��[<C:��r7~Vx$YTeǵ�M���͗*�(���@l�@Y��p�Z�~v�����zWB���)�����%a@|��p0zMڜ�9��(��!GL;����~s ����g|�6j�]�W��t�!�
ř�|0}[d�fk��ɻ
x�`���r��\.S#ԉ�p2�|){�Y�8�"��0�����:3UW�Z� *qD;sT��9=�WQ�K�iD��� gNT�kq����u��x�n�$�.��q�ªׂ���-E�zWg!	���G��|�7x?����<(p���3�]�`ت��cj%?n�O7d��s{��MF+���A
F�5���\(�'� /������#�,if>�ւ��"��{]����_B�Q�V�^������$\��ڹՂ�㒽!�:�ǩ|�qh�j��0�<���ΈH֩ }o��fPC<�uRD�w�)p�jw�����x'�qw�����C����ßl.�$��MH��L�%WS��	,��jd��]�͇���Q�W!��"�U �ΐ�'�!rk�b$I�=���S�����l�y�R�ƢVP��?U�]�Y�Z ��h3����=2���z�����9c��i�::]��QH1dev��J�k!��7��Q��gJ�2���ڲ��c��9�`��E(�X�)gJ�zTP�}�4_�8�e�y�����&+9[��ҷ�i���[/s���{�nO�b����ϷH���'�� 3@�Tp�^�yf�Ҵ�3f􁟡_��|�Bj��M�&�hh����!�b{��w�k���78NF�?`TYM�;��';��}�s^�.'�?9<q��\騻�1�RX�����Q�{�i��V>N�[6C�j�	j���X�}$3��u���,+��mğ���Tu����{��T�۽���J>����#��H���@��G��M��k�k��5p<I"���6� x��!i�M�YT{���
�	��'�]�K6ú��K�m��
.�1��̲�}�Pi���e�!P��w��X�FS1�ϓ��U�Zũ5=�������T���y���:3�V��r��bG�m��N5��#'Z����ܿA�|#�]b���]��=�O�\}P�ޭ�ϭ;���c��?ls/ml� L��)
�:x(r���l-�����kKOr�2��˭*����8
s�ި�ط@�@�G~��G�%�'9}R*N.��v��w4�*����h(�Kդ�?�=N��8s�4Y���S��4�x͡����Ln��rnxTͷ/�׈�a�ಢ� G��o�q�,�
��Sg �S<\;j�{��=��2��L�_�WE&e=���]r��+Mn:��)��Ir:���DX�}3e�(жi�#'��-1���g�}�
Xn<�sk��K+p�Ow�F�
��`9x<ɔ�F����|$U��hT�]�����,ޙ�.�Ô.ɽ�X]��⣦v�{:�L���%�����
�ל�Q�ڹ��4��W �-(:�ggE�V<O�^�^���5�̷�#��~!L�4��#�T�ސ�-���{`*	��@Þ�����7a�w�
4u�}Wȥ�)\�����`(��B"�
w]��Ps��W���>����)�2�%����Dk�Q�`L}V�s#��U'紉��^C����z��G�\s���pn}���LN��W�V�ʊ.�����.tn����j�f�M*v-!���!9ɫ>
����!�S�~���-ґ���ǨӠ���'LS��\T~����r
!�,�WM��J�Y��+��\D	u��-��ow��.m*�QèY$�Z@�-��3�T��]�9<j�N�!��,�`���>d�xݵ�U�v��23��y���`Uh/kx���	��0M��+��R�'�����lU�3vǞU�N�seo�VAƔ�B~p�w%�/�K��X�S�b�k$(ߪs��j �Z�����e�/��B�"�������Qn��r����2�J�kx~1Y�o��O3'4�Μs+�St.C� �MY�(����ԛ��`zW�i��������S�kec'�Ѓ&l[�`p����#�b2<o�iQ%�r^:v�Y�w3DK�7�P�|޵�d$W��_T�P�Q�j��v<<�
����V(�I�'nγ}Wf
 
	��%�1�`��P��o�����U�z��,���'�Cy�!���h�a��Jª2�A��\2�@=�r��U6y�C�,Gy �5��3��A8s��� O�f�o�a8F�}��@��n���G
n�8�=kdV/����`;T~�O�����o��B�^<����4�`N��A��L���4�L��?r��^1��y(�і,�	t#�,�bwv�	��aن����%Ĵ8ix#@K ����l�L���OUڼ0Wů.�?�	���,Y[�1��*p[.���Q�@r��du���)5�DZ�}��� P�o������(z�@2X�K*f#I�$��� dM�VR�p����,����=���P r����utL=N?@J��C��[%�"IE�<��m>�e����%>��rpv��eJ'� ���|�S�+���$��Q�9sH�v�Ͻ��LNT޶��T�cۊDcd��*גc3�I��[EVb�������Pu�v=T_i�;�4�I%��TΚ/�q��׾8�(�J'��� ���/Xǡ>b�v�kS�"�_*�����օ��)����OL�j������H�;�v��N�~BbA�R.�Fl��	�}��zs��2�t��A��,[n�!<1i��?�:մ�'/��2.|���0l�ۖaخ��(�D�Q��s�L��`���$�ҥ��S�&X �H�r��U�����<�i�[8��U�Ye@�����cQ�?*��r+dstEP>Z<62;*�*#&�H�?�&yf�k��/zfz�O���Fe'hC��:�������������������2�
S����{�a��y�_�P#a�x	ەn|&�_Է%knY^�-��8���;*��ea��Y���˛S��8���
���OLf�6��vHΐ��6������L����G�X�g
M�F�!���[�T� e�P�qXN�i .J���"��O�~A���"߄���E.#�ZR�)�_�T��������ۢ�4g�0��ٱ��½�G��M�ߌJn��M!c%�����ƔC",n>��Pz���@�Ȑ���u2��j(s�rjBJ����e��Wy��X��,f#�Y:�)mV�7Uu�Ť)Q��^�A�Ixo�-9�J����W�Ց�-��>���䌱��j�c���`�I`���� ��`~��@e�^KO2x�꺒b��."XH۳⳻2YQ�:��� ϴ8>��c�Vt�8L��mf�wtW���T~xt�ԗX$8���x���W�oD�~k�@i�D��H$v5��g��r8:*'ʢ�36��*0��]��NB��DHw�{�#�s�/��;�Kj������� ON@�i1*x�q�)x�����Y]K���FT>��=�dO܁���N������ D� �ke�/#�_��`\���ד�k����r��oi��4О�pI~�M��O��Kﳈ�ԑ�*���y���ŵ/�^@7�Y��{=�U�SGdLg��t�9)�o�}~�w�
��{g��@'!�^7����4m,	~c�M*N�����z���jI��Л�����#őa�jC� ��rIi��x�@�C\%��'2l��e���:��\
<\on��ڑ��f�L�h ��rO^��Nn=�|��%�>��w�`��=֫���}�Q!ʁm����ؓ��F�S/ŭ���2���� U�q��N-���=<��i9������&4ށ�����#����TP~�S�,�vz7)I�E�LM�,����\�Rv�䣣oE�#�B�|�!d�ʝhS4�̤"����I����yY�?�X?���6	-�@ːeh���*|��������:K�_�)���i�-��~��P�ؑkK�qi6�7~�Q�1���
�:u�0/�?��r~i�g@'�@����H;I��w�H���Q���k�Q�� �g�����;��y�4EB����n�p��26^
�pQ@P�	�7�����Ag��xǫh�/H��kȖ������-|���W���t���r3
7�w�(�#��R��<�g܍�C��XNک+^�?]���\K�����t/P�Xr;ם�?�/���ȠL��M��1:��a����)�0̋���s=�o�M}-�?��~D 2nJ���(�6*�v}7J��_p�R��N�i|�K�^9ТHC�����$3Z��}�ɡi)��<D'kž+k�_��`(5<�*t�aR�����=Xc�A3K|Kq{�5 ����\�_�<p_�c��B�L������_������u�(g*�.�h1C�W�:�� K3�h�{�>���*w�K��z������M��Ѹ��`z�dN�����@i@y���.�u~���UL������<�\s7����i�e��tZ���[�\:�����9�#9��a?U�ԖD���m-��c!Ю���:��!{ak-^r�)�E��Q��DWoޝ�ԍ¡�H[��D+��4�'	EW/A���#�{NAґ^���8�����0�4[�j�]��,�7���ɰ*���:K�mB�D}�|>�x���	x��	P�$Og
�eQ�:�>�c%�Zu�i�A�|F��NNNMadRڻW�I���v�p����������ue�U#��CsD�{��%��
�;�ďǑ�;&�ޭ�[H�zw�+u��2���O]?m<�� �r� ��e*�ɡ^���n�X��[���Qτ
skOK�Э�����g�p�e�Ҩ�ka�������8��4{��g�K�b(�}��A�M4�#�8SYN��U��ÿ{�fN;�% ���w�����v�)��*�V7Ǒ�a�`%���8�;Z�����ܗ��3�T����IרJ��4��%RA�l��T��i"x돦0�2�u��sV��k8ED�;���PHM~��F4��R�1	K���YWjL�C�l �͐K�偨�@��h=Jx��}�o��Az�A�@�e�6�ܓ.����$(��E�?#�}E�г���!)�U.%@�����='��n�	�p@[��P����,�M��ļ+%;I��Q	���*�W�5,r<����"��h2q�-�7����[��`���%{�)�8?1��������Gf���PT���r�^�+\'L/+��'�#Z)����4/"c�Ge$S!��	z%1�Y���!�s����� �yIr��"@�c �~�B�ӧ���b�Ep�"��<�>��8Ђ���ɋS�.�&phܦ�Mv��?b7sg���SaT�|hEf�@0�1B��JX6����s�j8�����b��֠����U!�9lF�w��\u��т;`�2��lU��q��[y]�q#����au���'��?'(����Z�(�#A����m�"mo�l��L|�qd)?i��e֖ 5T�Al�LZad�l���\#��W��� ���L܈��=�H)�L>'�A_� �G4��d���b/�',��x�|�c�7���Pݹ��B��*c�^�R�'?ʍK����C��~<���: {t}��u�]�m2��忇�`��v�c��sD(R�|��c_��c�o	-%���i6D�e�;��_Jp�W������q�9��]d{]�*	���m%��%LY�No�d�߁u�g/��}%����G���to���@�.�!>ݜ���Q��q4GH��������#"	 E������w�|$
��[8��,��<�E��?���X�1�"!ֽ�7��ݵa	<kN'�x�|�I6���&���x���Ɏ��e�ʶ���F���Y~#nC]����BFnߐ��b�^Qp���a��%��Q&����C��!!���\w��u���L�2�y����5��L9zi2�8!������;0�>ȝ�	h�ý���>�L�� =O���>P�J����a���`:h�2z$�$�ñ��g(����%�N㳿����$����
��������������X��˭Mr[����͵zH�{Ѓ��ԜK�v�<�ŻSV`|�3�FD �@.�� QOM�}�
?�	L/dm�
'�x>䑦x깆�o�T�r؅��[�|�Zh��T���ש�`e���o��,˄�g�p�B�^�V_���W'��R�ש��waÎ}�/�I�s�Ͷ='Y�5�eե�WI3���G� ��Z�2h/��0�\^6SS~P���������Va*��?	~��,N���r3�s��$����B11A �U�k��ի3>X|&i��hճVs5���:S��	�l|�$E���f=�8��~��y�Nu'�����{��n�0؂e�E��!��w�)o�-�K}w��<>��#U&�����O��0DE���n?x�c@c7֙���\���*k���2�ڃD�zL�05�*��QF�7Ђ�_t6�DA$��y$R�-�/}'zըKԝ�20��.։�3`� �B�5�.�G+R��{���H�硗+�Dw٥��i�������ݟ쀜Eu��!�t��HL�bv\����i�ڣ��K?yv��=�{���ϖ	���{}?�n��ߪϢhЙ�,n�W�^a �P>D�i�dCTD����u��d��B�x��Z~Ќv��k�^P������;����8�3K.9�(��aP��`�J	�����{�к;�u��;�}��������!Np��p�� �p��6��ډ �Q��'�^g/%fO��糶��]�o6�;;���Gj��!��� �}�����W��\��p^������LD�Kg_��6U<��]ǇyE��^�;��p�6eY��}�Q��y�i��k������{}T ��ZMT��E�9:N�Un������t�N��R���h[#�#@�o�v�ǲ�ȭ� M����N'�4����*�C�����_�����,˜zVZӚ?m�~���e��,�*�~���a���fД<�h2K��5�$C���21W�&�m�ek�c�b͐Tc�K�ӍaY�v=�ku#Tu�=(�ڋ���g1�G[[ʔl�<�]H�x[U6n�Y쪮���n��`Z0���đ?uJ�̑�f	nW�B1$eYCTܮ���Ozo�̩ڢ]P����cFiQ�����w�lx^�U2��n!�m�]��#�EBT�@��.U��D��
͠E����D������w~G��
Q��6��
�i�HFP1�i$�ǵ[`��\F9#��i�<��y���wÛ�?x-FC��X�5��Z��m���+Z�V弗��o
��_��У�g�Q��ݤ��n�_Ue��'&r� ����@�Z�Oo_#�0���c=�����a�� Vu�uT�÷��|R7����~�]�8$rRâ���y��fnD��㗾�t��YS������\�%�p	R�B��
�є�WF�}�~j/��?�9�`��	�u��>"��8��Зh��J#���G�4~�؞Q�`����ل/,{��V�<�b'��]�� ����GD����C"U�J2_��Pɕ%-H�$�l�6�#�%{�/�u��63',DY?�b5���#�[�(Hd$����9V� �f��.;&4�����%1������^wJ93bx���n@�mO�(ym���M
Bs��+u�k�q����2�\}Na�oiN�@.�
�����+�K�^���� �mȏ� 	���@a�*��A��DP�.m���Ym}:Y�nԌ�,A��mG��'I!�J�յ��_g��"�����Zv�3ԀH�^���Gψ��F��l��g���n�4x�>;! i0����K��(����]0�8��@+��#��ۘ�d�<�c1S��ϙ�� A�a؋+
���R,F �IK�F{��R;��@�$��m������"���=cur��������C5���aб�Q;T��n3����T��l}�
��$���^���݉�6[��:
�H2!�����|�x���#��o�+)