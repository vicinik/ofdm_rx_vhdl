��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�G'?��,���ɎĖ�7�ŉ/�c�tIo��]_��Z�k[���2+��IZC[��\���Y�Q�B�]�[�s��݋@�1^��ukgf௿�۟�SW�ef�_ee��F�Q���U"޼l��+c3xr�VO!�&s�jV�ұ�f{��ߙ�q�����$��(4��%1Q�Y$�p�	M��S�Kf�y$�����a]B�-��B%ӟ��yI0:zSr����2,tJW}�\-�|���b��ٓ	�Ӂ�M�@�e������n4X�w���Ӑ�����{Y��]��@���X��讒�2��/?����=����<��tq`���8�<�Y`���`S����}��mJc2��YG�=�r�f����Y���ov��OC���~ƶ�Y�>�������F����>���,v��D�!��pƿ�b5�7�Ҥ�1aT�j$*�}����R��֭�vY�u��1��T�rOB��,������K�����l��Q4N�W*>�F���o-���F9k/m�V�	��?�M-�x���"���B��Eo�׀H� N�@�yJ�>XC��:F��@����*F�����J�,��#�88�=���x�w�2��l��fСl�5�Q�]��6���s^��ٌ��`�]�4��5���+��+�S"^Q�<�ݐ�k{ffu�"v{c�b`Kɮ6H��ı����2D��R^��[
��B?�.�f��ZG�����'�%U�]�c�$��������$���{jǮ��HRc�ڣ����GU]b���\��P����P���n9(iM��l��H��%'��������fh~yfź��.B���KG�z�P/���>�oHqC�x�Qt�Cb͉��Y|nL���G�� =O*?Ұ�c����̄�;p���-�s�n��y�^��ִ:�1��D��X&@	��Ŝ� �Ԏ�kj�i`������Sݕ� ��pm��;|1�� C�j�VM��3P�����)24q��n�&�S[���Щe{��T�h5�E=��{���
�a$�� �q�l��r_M��{�1Z����P)�Օ���h�Ǻ��mXUr�w��#dƠ!�X��EhM��N�r� �c`�l�,!��fj�>���?aAcA�fВ�e�Q�F�����2�b1�G�䄠N�Hͬ��#iM,����s�*be��W��� ޭ�S��Vq�Ҿr%H:d��>"����T��L�7,0�ҩ���=�� h����À�Z�X>��_�v����@�k>�	b��f�!�W.k/o$�&��K|}BQN�5���ȧ���Q���������J���ݣ��K�$W�)a3�W�Ơ���T���%HR�׆}6]n$�;�-�e����	{�'xi��E�OB���w���6��ER��
��7y����ûU���l[V�x>�"�LJ����g��h�_���[O�>/�3疾M1/��cP�䷓�����GE.|+�긛���_"��:ISh�^�cSos�����C �.���ɍ��/�S�'F(bu�v�%���[;�Ih���yю@�A�Z�:����٩�:X1Dm�K���)^w;�F��X��E�a�:�6y��DAy�^�UI��E�
��b?�:?�.g�EU�݀�%׽U���jE"�'�s�[/�LY������$yAx����Y��^�(���L]*��%�s�UH�T�q~-B���<�y	U;`�R��b�t-��Ɵ���S�������w�iĭ�V�<��氀m�yA�11.���'���`0�h�	��j9�?��D�'*F����LoWW>7�������|�73���g����-�IK.V6|�����z�6[F4ِ!�ϔ�O��Y��l��It��3�s)��.7��K/�c���~�ƻ�: ����e���"E]��k�f�H��zV���[u>;Az$@}5��h��^WnPV�n6/i�/���:�"��kw��1m*�5�y!s�����&�vzW�,1A���JᎻ(���G���W�Z���n�ɮ��$n6�^�fMK�(]5��w2*};` $Cߏ;s5�Ea�O�cG����a9��B#�+M5�5��fXy�2Zev��#>�[G*�}�{&�zP� ��Y��q�d,�a�`��X��[�z$���nmsY�[C���KZa|6}�k�'&M��1������tۏ$3^�B���醨ͺ�b�v��?��-f ��X9
,:� W��@6XT�!a����tـ�J�矵YP�b5/��,?@�ׄM�K�sMb[;��������^��B����6�r,%�P�nS�y��'-��(��I2⌺0��n�נ�0FY\H�>���3���z��~���1 �@�o��=KС9=t*A2��-V3���m�y���,�T*@��M���n��L�AX||��q�e�����V�=���d-Y8�Bh�˞Ff}�Y!:�E�GIibW����0�J���^�QhjU���M8E�ç)և#��5�z!���}�1j[ˑ�e�y�H����c֊?2�HE{#�35��Á���g��	�����ip�+T�#�rt��x��Ǟ������m�72����	�C���^�T�H�``��]a�7��(�4�$����ں��9�c �Pk����vBp?��#�T�Q�9���;��%H�l����{�c��6��f�����R6*��Z�hE����-V���q����܉���f@����]��Y��
�J���j��B��S��|Uz�3l�;p_E�O�}#��W�E�5?8���MMG��̸�!"�Z���wB߮���/&�ֶ��^`�|�ʖ� <�b�	܁����p�r�,g�����(����iZ��D�9qk��w������K}�B<��Y�]S���N��?$�M�*�����\����c,���n��*�p�:��d�c���ϓ~���\���P�Ĩy.�$0iϢP��&qf?�VH�g`�����I�B�x�?�s�F���b^�&MLs����cx&�  ��	t�r�RҰ̓A
Û-� �ǚ9d�S
�� �ߦ�2���Rx�fJ�>��	i�`�hf��ad�Ǆ�����(�Dk����cw�=@���+;ի���:���ƕ�gd9�ud0
k�90T���%�\Һ!ˮ�P��;��*/J��~��z�BQ���y�t�B�;�`Ů*pV@�����#	D�{��Q�E{��j��\R>�"B��
�;6� R�/��%xN����#�l�d�YAw�����@�<z�;y$}n$:v���׿2��ݎ��_��G��e2����	r�@�C۸(��}�x3��N]�mO�֌�;J� ���^��� �cC�4�_&`���+ߓ�ȫ��I9���qߺL0�~������M9��������6T�R@��N/����I���]�o�8Hfq]Pqyq}��9B��>�{[�B�3�� ��j��_�(RK��k��C#�5�wwc��;��!j���*����<��2�D�n�5�!��9�#��!:����M�;<#�:�n?�� ��������O��x�hr�Ñ6r*&c#*�ٖT��$y�_������Zu<WJ,�g~�xT��+��`6��$0�c�h��Q�3l�F0'QeL_��=���g�@��5�.�8�X��A�O���B)"�y�4r �we.v�� �O�Y�Mþ�7��[$F��P��a��E E!�\�%�)��X�<��d����lw��{[�dl�N)�Ȣ���)O~�P�R��,�V������`��E{Ұ�r����A`����!�����d;�3N+.J�[�dG� ���m�}�p(�U$�E]Ĉ�ǟ�������SAYY%������W ���([*_�z��7���1'��8��[���Z��0��;�3x��ٷ��(��U��tj�Uc���V�ut6	�f��H��%�u�#��$$�w+_�V�Ed]7�[��Y�|� b�Z����|�����|NnV����#����f��
6���}�0�:�s��y�c��/c�ϔ�{��fo7�.�/7��0n��J�'�Ӏzi	X��C�9u��=p���k��z�[k����K�Qus��`�yh���:�����Z���Q�xυ��٠�Vb�ǿ-c~hK�D���ћ�nw�p{O��S�
��.:��)�5=�#�m�>���n$fU˿o1�i���w�a��R����Γ���CeQE�!Z̩ɺ��=�t��9�̬��?d�X*o3����7C�W2��������7�;ި[�Ǔſ!���S� �D�����O�>1�"H��{Yt:�",�nP�o�v���L�U��k��UjW��0�Z���"�Je9M��r_�i<��Z�Аt���������=�ת;N�`c}���=p����2�^$	�
����� Z\��Ljj�5ӡ��:���6
U��
����y��b��Ce�� ͠qgʋ��0	����cW��	Y2��%ڜ�fX����ؔ={�ȭ)j������*�0�����q�i�M��_c���P����7����$��j3�$�B6���+��X���S8
r2z���U`��Aw��֝�p����Ŵ��~и��wo����@J�&���TSd6[8��ʋ���`��GX�\$b:r��(�1���<�����V��<烠�K�4���ʂ���� 8iY�[�@J�x�+Ą5��Z]Uj�q�Q�6L\�x"�9����ݤ��\�[�Y�)#�e��/���u˗̲���,���a�=�͆��fSE��3QDa?/�0����$�i�� ���k�+^�=���ѕ���H���8$��#�v<�G�C�9���U�h,�9R&�|X�]z�v8�1�w���q���T���#u�X!�����!�����W�2�uYo���Y���g�yf���n�̍LU!)p�\�V�b꽦{*������|�%^d�]��+
��p��#FM7���KS{HB����7�^%��~�]5��.���C����:
�I���@���4
j��K{�ym�CX>�<��aF�z�L�u��0o�FYmb^e7M7�����<RBe l"p�4/&�}��Ñ��Q�I�G	�pT~�$�2d�q��]���0�V����D\C�s�^�7EL�i�5!ť��f���
�Js��7`���4W^�瓒V݋�F�0�4��=�?��zt��(�L{��0fb�HXM+b�� ����t|SO�(�넖�cMs�)�/��4@k�f���ֽ��K;�Y�Cid�-����B 怬G�;5B���♿	�MKV������s�r��-��l$NL"��y<����U+T���!�y&'s������\i�W���|�	KP; -��t�.7m��TQ��L�[�6�l�xI���S��ؚWv��w�+����B��gAx�a����.9�T���iUW��4?�[V��-�=��"mJN�X��v�T�Z�>���ZuO}n�E(n�S��24�� ���03A����h���*�`$��sz�	��G�l��M��֖�G���K͍V-rdL�d5s�h����N�l�`��Y�Grz�4\��FRe+f���ɼุ�]
HW|=s�j�_Z�E�R����Q��G��lEq"�;��jz� "V�{䯵K�a�}�����
5	�Ma�g+h�h�S�5�Q�DNZ[3��q�m#	��I�A� 6Y����@u�{��F�G��A�x���xE ���
ZL����:�g8��(�D��=���I�����߿I��|b=l�mר��gz�)�d�'�N�X��咰�������s��0�[g�Pkl�3<	�Kovt��V1 /K>%K�O� Zd������L(k��	��i��o�.D��	�5M�Ys(iL��������·���PN�鿭%��ϡ,��һ��ާ��A��&o��N~nUw�]��8U�Ʀ	/~��(�V\���Zr��C�,�6�+�dv�}(���LNpW����h�ϱ�ڂ=��*��0Y��p�1�i�4����~Gh�ښ�o�w�Q(�������2�l܇�S�d��s�Y�yC��㣞T��w����-m<�?��I1�U����>������{�V%2%2UB)��y�`������km:��r*�)��S�������k[��Ȏe^��n"*4�� �В]�yK���f�����b4uo��87�_P�v�u;rn��*���i~������!�r��hF�3W�����t]��K��pa�ȀM�I�<Dk�ئ^�*%���v�s<��|ٔ��ѩ�sC�C*�_g��ӑ��P�GX{�m���,���ۘx9��;��,���S��d�|�S�B��ŃO�]������+
��o�ೈ7J������F�k3L"]���\�X�K�gڒ{�ߤ=��J����|(��N"Ř��|��@fw=)죪^X�N5O)� 繎���q�t������썧Z��+��z7<�#8��]g�JU80kR� ���s2��諫5��.��{�����ٔ���� �!5�:�[<qǫ=��4��+��i�C�y'tG-�M��+�"E(�*)\Z3��@g�!��|��֨Bͷ�y��eJ�ׂ���-����v�\�,|�����}��R�<N��
O�������E;�a��n���_?�ӗۅ��N-��b�.��g�-��tHg"��I�hkkYp�i�6�"w2����uO����#e=��������t��Soށ��?ҵh��(�b"��N���E�6w��Z=�������i���g��:�&�H$YX�h`�{�B P��N�v_�����=]Z��E'���>���Z�{��C�{0�	uˍB�w]%o�@�+-��D�����?Ξ�]���CD�4�5�
��r��l�rtiq�|W��oO��4�3�F��gk5Kc�`��F57�j<B	9���oC��4Bq�g�b��xu��c#�]���rE�lz��8#�d)%H��u�_]�`��c�G��R�Qc�Y�n��O��Z������")D�?
���G\�e[B<���;�C^�-1yK��x,�� �Q�����c���X���~G�-���a9R������;@	:@���\���+��X�J*o1��j��D�����e'[nA��A�W��!���N�~�/͉zOI ���<ķ¨�]ҺU����6�P��j�=�9�@���n|q����~������͠��R�X�v���d���}Avj�]=M,π�h���*�������l�;�Wx)�}X�*��I�I+����2�߆��d�����D�f;��u���)�dY�����<�忹��Y�P%�D��G���1���*��E��߱Z){�K����AR
`�Z���w�V��H�8E���\����B��
zs��w����*�~q��%Z�8�{f�I:Dh!��$�j�l>j7����t:z)y��S��5�q�3��ZC�}'�ToK��k	F�\k}p-��a��u5եт�)j��F�)�������1���!��$i�ۙz������Q�$�
���6��m�U&$�*`���~�Lk�N4���$�����I8�G����8w��^��69��?�?G��:�P��[Ke*$P��>1n;d}��`d�S���ğe�^�o�2�J��I���³���#��/�@v�S�u��)�>?��D��l�cO���%�2Dh�/�"�Lv6F�R�r��C��x��elFXؿ���Bn���1A�m�5�X�ohʹ���芬�)���Dy,W�i�GR�s\��1���c~�w��W��ɗ�rp,+ch����y�'ae�0Y�����5o!A�����6�F��#+���-���ѫ��\�Y�j�� &+H�v���Z�V�ٓr��(�kV[L��~6l�8Y�U���P�>^d�Q�دY��Ǚ] #�JB��,$
�tμ;4*���������� �f���B�*���I̷��V����r������t;�#���F5�1���=�p"-�]a�k*)8�&��w���|A�'M~+��@�����V\ZC�8X5J5�K��+km`�G츔����΂����g�9��R��0��c8�p�'V;r*=��B�>ޓ3�(|�m��~�<h�??���++�UE�	�d6� �1e��x��u\�3���K�yd�β'���[�E�E �]������azW�]H���)��쿄Dv�2�m��w�lhvf�Fĳ����|怚z"]�`W�,5SQ��z"�t#�ҮUh�,�W�PA�yVxX	�s���M����-uы�=���Y��W[ ��������M����F4���#� T�"Fպ�Y�jN����2s��(�:Q"���i�6��Q�t�w��%
^W��aY�n�y�p�����a�Ye��,"�%7�<� ��c�5��y�t��!���u��g��b%���Vꊄ[��e��N&Z2$��&dBc���%�)�wQ����Q5Be�{3QF��5�ɗ��Hpܓ$�/#I٪��<�v&�}Z�DϹ&��������̣���8�	�c�)v��0�<5!;�I��(���/��*S�@%��h��,�k9��C�}��I����D��e6TwU/��񄎯B��S�}l ��c�ظ����\�e+7s�����X�[t���⸽�'�?}���W	���o�1�S-ѧD)r_\����e�e��Lf؛��Yas�ȡ�mc��؇��$)�lg�K�-��:<-�z����$�I�K�V��7�?���)���i��:+�V@Z0T̿�-Q<N�'2��ٔi��ܞ�El�y,��������O�Ί|ƴ��K�j���9���J�Sp�?��[���D���"��2�ІJZs�}�B��!���0�X�*��I��A�U!O ���{�y2�c2d�'h�y��6A�(c��rC���M5o/j�ឫ4����'6)��w<�%�0��I�`d�>B�_�2-��G��n�����F&25��_s�B���iw
J�~��oC�ҌM�f���>P�s=x��)�+bK�옵0�,��D��i�W�tw��ԁ�G�-�9���\��"�y���-�LO6'��m��)�t[=	7I�����s�����N1^�ΒΛ��S�Y�e���K�3tb�覧�N�1�� ?Ys�{�B���qB�)ר�3�p/%�}���/Ks���A���j�o�Ð�e��)��*͞���TVI˗��
O����E���~��La0��s�(���ȸ��,RE��;�����G�b�9ن�vه�]�H���k�N�$���)�B��ҋ�Z��D�i�CRv��]��������ML�+�{����E3��WI�ފ�|*��2 ����E��#،���R$�ҽ��m�����:*�d���qa 7z)�+C!�n��C�CL"B	�u�&7�c=#ȯ0{<-��l�"ҡ ��
7.Z�5(p?�X�X���6_M���w�3��&���6�H�l��2
���ŷ2b�
O����� �v'�906�����y�d��&�E����є���$ o������	��&H;(:�v�$�pdr���1EvOwEb+�WV;��T�j��R#�M���S�\����N_��G�W��Q�o_�;c6��	�8��Q>P6O���R#�� �N���x�&?�Yl'w��L���>dC�B���	W���#҉���Q�L��v<�|Z����'��~��DۨFT��x�&����8�u��*��(v΀�f����x-
��fz��ܕd�$�}����+��n���*^�d���!,��4�H9���(�b�S�9���F��B���0�ص�qu�����>�c�F�o���E2����y~Ey����G"ѹ.�<l"Y-d�LM��jY���R!�$���*���AN��"�Կ��Jŕm�E��%���S��6Ԯ���#��_��ڪ<�q`PC-SX֜&�Y���G�m폢��&�J� ��S��Q9���[�{�KV�c5�l?��\~����6[��n�oI�&����?�d�4Y=3�q�m�+��7�������?�O�)a9ZQ3qHz,(GH����[��Sʐ�&������9j���c}�9(ݠ$�_���mJ;�rq����ϯ��J�3T��>s�|���Y|͓x�*�f� ��a[U��l=����pE�����3�nH�l^f�:B�.���ߙl=��wu�?����s��KU�2;ؑ�\qb^����n��W�dO\*��h�l�E��>."�C��\0;�2��p�#
��鳓���&�i���*�x
=Rie"�;�u�7�2sP�!ӉjZ�(�\�«��>�흒��	v�\��dY!��o1+}�n~|aV�M����f�L/6�Wqj�;n��
)�%�y]� ��q�d{r;��=�Kp�00��	�i�Ȱ��"t�Vg)�*n�����J�U���B��9��:��>�j>��t�h��_*�m�`��ٜ-1~��%���=�)�" ��|:�� �l�����.@*!�;'�:��jxO���/{Vx�R��d#]��:K򨘬�#GI+��a����Q[D��w'�f]���������d{u�`�pl�s���W��;>��W����A����I��+�x��~:�A[�,\��9e�u��tTt�С"2��'t+��cZ��?��	�0�;A���=�"}���M>�����-N���[�[E�W8!{�-�H�_GhcW�#S���o��a�Y����-B�]u��֚AT݀<3�i�1'��i�T�"��y�ia��L��ⲵ^m�u2����r&i4����Wl�T�F`g-�Z,�yy���W�����~.ۋJ)k��_���d���7u��X�,%���P�hR<0�2Wh2lh��.��yj�(7�M�ߣ�V�b�����@ڪiBn��'1���k̲!��U>����!I�H&�Z|>���1��h	- �s�Z�^�J�x�� '5_� �oH�����2�$ew'L�"/��:'NBdd��!��ί����Y��T"P=�t��mֿ�V�=�WM6����]�����M�}ڙ�V��{��U�<"�9d�8р֑n�v#�,K�ӫ�ȣ�F����ӭ��շ�:ph�pu�M�>�1��IY:fq��Dl@�	��;�݋Qg\k�q�ޥ�����K��sM/*�&����D��ߜ�Sۥ$/M�T�u�o�r3�*�)�d�y�Oe(ڣ�t������;�࢕_�V.8ђ���E�rů�rU����F]b�@�@����JT#M3�!�S����+� ��q8��BOo?�j��GO3���X/�{�R�i�O5��R��S���}ʌ��6C`K(�x|P��.���jN���G��W���}(�(�|��h��Բ(�ފ��i8�����3�#��1�B����E��vPO���Ք��H�z���],/||�e��$�C�｛E�e���W��ڊ��u���� k�/����`B�DUHg'�oZ"�SXR<E(w��OӔ��w
�)�Ұ����[T�Ѽ��{,���r2�?��'�8����;*@2Qm��"�ΰ���N���uL
�5d?�-&@�P�J��Q��@���sĞ��?Z5 ���}�-z�+x������Tf8(H ���)���1�F���(�>�D��HH(��8I g0<�Q8�t�"�����T���:Ͱj�$���~,������ӛ�:ٻ��ˊs�x��^���It_F�t/[J��a�,f�R�(1��,��)WJ>���n�e1K3[Ѿ3tu�X%�f̪�nV�+z|[�$����������	��@�`�W��d���Ĝ��d�I�t��׳���ߞ�p�(��5�z��)s޳�i��J&$yE�_�TI[7і<�AB�����@�J>�L��ɔO@�����n~���(�[�(�T<QeEw֯����J�r�:3o���*n�*�A����%��7�Y`�;R�d��^u0�e2%�H��UjO�����"�����*��%������K}���v`w���ؚ����PZK�
opr��ה����j����	��/\4/omO��"��v�rD�e?}/�i�V;�+W�*۰���cp����ӿ���9|.���3=�w��9�)��?^��4h�B��Ncsm�6Q�G��^VSfL����ַ����p�\8�ݨ��������	r�!��@��4ߗ(ʻ�﫚f��oxuP�D��)��׵7^��_����3I��٢���8!��X����4"z�3}D��	!�2��"��7&���/_<T& �):J�"V��|��|���Qy&��I�����{����^�$�82�"0#�ۖU��+�"I��2�<;20@��6�N��t���?F�'�ѣ/��1x}lb*f*-��>����@+����?�cU��Xcmx� ���e�X�)�_��� �^���j@��ZR�$ }�Z��q�