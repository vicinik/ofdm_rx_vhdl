-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
I0E6+H6l+RxDFwkfUrlCaJppFi32ES7WXHraw2qRKYqt6V5R9FgLpZtu5uu553h3mkA7PCqqRyON
um7DOVaJBJsaX0jOqI0ukSI8vkDRX6qmdcyPEkDl5Mq8rOqg4Q2si3Sy9CEFWLR2/ah92SLHMJJS
Js3CH4Dekr36Y183yLMcspuldo2bMFL+wpnjYwxGUmIEfqrKRuq9W7/zVcfjVQLj9o1Ab2KKU1VG
/WgnMbiPl3mWySandJgAe6MfCtwogW0RSqLGixBp+GFnQ+2Sl9TR+zmWMG91MI/2Nv2zsXBS+vMJ
suSzMVa48FYNfw6spuYG8CpBr2JCGSBSi0xU+g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10752)
`protect data_block
mqWVItRxfCcCzM2dRzxNhpjctBjzNfeEOMgkBioxiFwkgQwQgP47BUftlT/bnfHtRSAiXcwRNcUI
jZfx5DBZh7HjSXfCIWPjIUKno+OBvsJ21Y8uKEa1V7SUTcjwK3lNAS9VbGyzxGenpZU+GM1eqZfZ
3fZCc7JsHwMis9qhJiYoQ+EWj29P3FhzSb34cAW1QXQ7y1+mMPg+BT95n2+5hTNQ9IkPUfQEyqV6
Z+FLEpZNuhqVAHCmcjeHBkFzze2HzbaKmSVKtpWrbrBPxHNiHv5ozAUyD17SKX0k8VnDuKgRAoj3
bLYdvs99RrMgs0Whxoug/U4ddopXOsd0IfIY5qoaw9d6M5SNsVDmtMDSWORKP10+2W+E4PpiKv8z
XG8O/ZPlnZpuUJWtvculbW4O8iiJQ6Mvi5Wv6OIfOYxsHgfX40GSffulOgU60GMzeWgS3T+/4j9w
Hnc2PrrvXBNARiYUvl3xwkgyEtyekw1PvGrNGvGExcIkE+HCaafxYseCDlUu5hO+WRgaLfLvEQ0r
kMp/06RGLrolcw/fvw+pfGqUz0CY/1Zj0CC8nOZbEUZu2blsBc5o/cCgLL8RIltq33sAH8xX3XIZ
COr37jAWF+iy7EkZb2cXG7JuP3bACyhSqL5FSCNzsiZJSsUwjDQgUWVamXdmxDQQQUfF7uzC8BaS
lgR12i/9euA8Je+l+t09vZeFBm9jaSkcjDv15taLBUXi0GOY4AuCj/dd+o/kdiyRp6fnia04768b
y1zANkqXPxF23hnXD4cFsGvRoLdWL/bRB99hsL8YvzUR7jrVtL7RzFB/E3TA4ml0/RL+6BJirJLv
V/nfE8jjTP975o+66eodrdRJPjjxU2Tu1rl+HqsG4Tz0ZGFfCEXRrQgjZ/7+FoFh8S6VIXn4L2ta
27Kr/rnvBnI/jZl0+Gc5B3URR7PO//PczRNbt3j8OkfDMX0E3pGDD595RqmuLeihsaJRm8OEGDV6
FLdm7ofbZCVWeYIegJUSHIwbaP7FQCn38pSy2y8JaeC80ndj4uDYYHIyLqRf0GPPUchO29qt92FT
vI+az51MTLx3HAalP3twjZ8ZVoJRAaVlKK2lFwwhtMa8otjfyKMp3mw9WHO8MwRnW54GDxmGG48n
Fp485LV67j4krJDa45dKM/zotfOvw4PKzKwWedrk/6i2TlhQqdSVwVQ8Swsw1vNQcNZ/F6Rrk2w0
m8ugT7K48DN48UlZJZqCk5+B+B74ss/nQKTK1GQ9A/2R5mvL+G2/M23kGhWGbj6Olv64RtJFuJV4
q9hSXWhmuJROCdYd72z+HRJ9WSAfgcdJIK95dXZzZSEXMb/2F4zdbVKW6no6GpV0a/9rzoQ8Ko+F
x8mJVj/yWtdqpFVj3XA7rKYY8V9zNVohIZbUALhX4exTlW2DAJIB9DCoFVV06uYF8wi7pn5RdH7n
ztwomEmJN2bRjvSIthZzRxvXocIywd6ADvT+wWcJ6k1SNWbEVuM5Ybe4rlA2+qc5eLyP9aCHscpI
abZcreyq/bkZe3YjoLeV1QhjvwgLZKV0dAVYTbSi78gyLGRt6bdco9FCMwSZQERp5Qy5G2d48BJF
dqjT6dOTcgQRxn3xSwIY/sJVEwBE8gq8BhvcVpHyFD6/NFcv+Stz8YqSGw3X2CdrtULefr0lfXsO
Jbk7Vjn2FLqxcDgSGByK7/vNJhcbAIcXMkeNCvY5mASrtgLfNDMBEGgG++vEI20NC89nPeaq6t7F
xMQNwi5q2E0TvZyOJfnn0O2tWIe1uoop52Frf/MSROolm12gzdm2Pj9B46j5sZCUjNrJTRc++tPP
ldAt+1/ag6ULX8NRilXf2Un6QaxNmDhCiODax5MPnG/ayj94G76qEcZM3TsJ5g2o1APqx6He1SR8
nXhF2EeeQYy38PDMHKpvFkASZdQA7J4lXB3RcChsnobn0RYR2gU80Q+3JiZUzypmhY1M0JGYmG1r
t97PrQU97k3jRWSI5EEOwqzmkuNzg/DWrDCsCgF2Op231e4mlv+jEYzY6H5jTNtH3lg9WfGrU+5s
TcNu+7n3MOIdRlnjmJTZnVCd1XUFQ4dzGbriqujP1yUStaU1b3LbuHv01tu4FDxubjHrUtaP3+WX
2mfxaLRV1uQlKORCG4oh/1Dp7LXgQIbMkiOIhUskRJFR2GT4wy9Av8HKEGByq4WDmDZ8t4x+8OR/
2yQSKx0jIL1IoN50gFttQ0lABVjRSF5ksYuaisNb6THiyrTCdRwwhr65ucMf5VSgOPkEgklaJJdR
TJWAkiREX4bwniXy1YEeMAdFFiPhx/HCn4wtO1GCZ+9YbjHi+qt5uclAD++uZ6Le1RoCr9KWjh1k
JXpu2PTjaJnkQLjKHBhM5BgC1rHcbKVqcPtRoAMrHWtyNxChO69Hk662/OFFl1fmjJpTdypZCOQ+
mNMGxUUF531eLZJIfIWfCaRslQD9gEWMeIyyPgDyZ8xDbXkFoVc3fgPrJg/bNY1wKbwHGSQxNxWX
xorw0plAQ3LbIlLhibmEqrVqBwC2uU32R44mzdZM2HL4cf2buz+CdN8kd2PHLp7IQ0k7fEXnIHOn
fP3tR/9iH6UQFG/RmDCwEW0DyI+j9LlNjbm62Bv5ezsVBodCqguyLKFT3SagsS8eyS5DJJofNUCO
IjuLOZwHn35lyb6aYDvsr0AS7TMOCBalA0elrjbdYrfT4v7x9cwkAf/tp6hk9iULfmDzCgbwYUHK
yKiv8Jp2htiItYkNiPKvWtdBRfJSiQuXHolpuZLyCN3rk+hmbbRMFbbtFkdTswTlQFCZOEqcHDG8
Owv++DJS/m9UO0EDwe3tY2i+FdGqQuHCvuBWYU0NqFQqLt82WM6tLWVwNXM05jZ+MZ/Nl/ibL+Fw
WeQ/2RWf2iE+IXg8jfhfR62Dycnh/KfWb8MzuX3tGQuHroemCzkbSxjo6ozOFLmwtTLkA9MTpSyv
qZ8xvKKIZQPMkpKMO4iyy7UsEIvUvbB6V3055GpSyy2SfiekDax3Z0vjDUIGKIgqjkixmAIavgPO
r5JkxMQCfX2SmQoJsY7GCQdpj75yY5aBdknx+giyEh4aXlXgeeRmBQ8xD02ZjTQw92tHgCDJZsH4
KYPr3MCbYh09Wscj8IZQNTSnELY8aebCVlMD/XT3R/D0R/xPm/yu0OOBFTJAgn2Zq29zJVC7xqOl
Legah7ApE5iJx96cFzh/3/3GPCn+4oCHaRUPYaPN6tjavvFU2LA5k+b0sR/nZeDccroB1kT/jh5G
JT+T3g70h5hyZBGABgSYTBJrgS+faQ+0kjMdKOdH8/YE577PXsWCzGtJ06FATWu/oAzd5gS41hyC
y0AX+fONMRDlnFUQ+G5bFsrHIGnZ0oSRkceH7NlUelO9zcR3g6+Nm3bw3yddXZ9xc97GN+NdYTJu
d3kuNL7IJuk/058FtQwXpyyYxQZGuTMvUvbOC7QYX0W1ZXOTXrhuw4ZSq2Y82ZXrJnRLSaxzPHRA
HtUdFvfWJqq1c9koMx0vKkc5sfOuMCueuNOctyBGLPkjPxpXkP3IvwY+PjF+gcegcp+En3iEzM5K
Ci0Ma8NKVnSOBqG2VT4JdK1hm832gUN3A0GO6/Kluc4JYJBDu95t/JwHpqS8ngepVbWJLDJ6xrR/
BwQwvT9qatLHrRlUxVpEs+jV0BAbCTOlrStKumdnJV+sx/tJvCKCNCGZw2Y3B0P/6yS1y7KPAeuA
yevLKWMBxzbjPSjyqi/4Vr8mcY0fxvSJSYywnuw/xMNSuvTTZlFDU/95I66taK9Fr9iEcS0pxRaS
AmjsD0sZ/cTOofbh/itn8VgfjoFsB8UDE2tvnQOGKfgO9fM0rMN0QNzILP3O69yiY6JwFks7LbcZ
URB1Mi3FfyT9skBPxffd9mVNgzbkzwHWDkMsI0OSY64Xh0ldQ2Mc/peOk55Wb1V2mXMC68XFDOfQ
89EmYl3mOIizSVprTpLTbY52PZ1jFaOnYwG5nNKIGJI36lhPcCeQtA1H8pS9S8GM+UL3g79AfMRO
P7cs17w6boARVTiC+ohSgRLU9w4+FbwGXXaVeq2XOjz7q4GBsHdzvKLJExo1c5TCOy9RkGf2foRt
KTKj4+mG+v6Q729XKXJxqlLpaM85+sKZeYz3eGMvgHn+7jeKF0RfP4O8tfr151e5ZONSF1qYenmi
jb/zXptt/QnGtDBdTu4H4p8evkclXgmEle+lbkhrZnQe1/l+goyh2/ZaSVpDOTdRTHa8XC7oTtoe
3yB4jmj6ekKIFT4jjFf5sK/mYL6uLa9eRaasbGYylaRiZHfW8jjsdZKkzzoyCMwBUwFxyx+E3ksn
e2Ybj8CLXVtkA/J3Wx5ptE5KvP04a3JryjDtAEOuUuo6350ykB+/fjmogL7zf4nBHGjNQ2C3PCWN
9CHUCP2s+8EgvTI9oiaRnWh2BlVV/vNJIpV2x1kxbo+fdPAx5dacX5ZSVcZAQjWRiUqIVT2AglT6
7fNq/B8OB9+Bo8EA30g9T/Mn6HHuNOZQhOu1z97hMdskZoAUdPzd0bVjoiW7/ZRAZ2CJRFNyE//N
b+3D1qoBvvcE+D8x1bpOOqNJlwjkh8n3pXE7VjSmjspNBqm8SHjX2LobQjv7vwMPOSDX0g6CYjbC
y/y6kY5CZF3mtUcsH8YwugYvo5WAyaHyHq0mRontnBl6MJwoA0rao/Hydzh9+sBHN2YztZELLSw9
UwqI7rk2Hcn71cq4IPgsm5M+pdYQr3c6XsFK3jwUoyoGE/IUdJxhMafJPijwnEwBK1t4IsSdugoM
UuNO6vnNHJbGPAXtNqG62zX3Ms5arfMTCGhXyW4FMEfkdje80UEOTZKJtSZK+luWPdXCH6/IG4HH
gmw5giqGVRPlM3HsU5i+uByVdnn0NSieGzyRRaCGUpcojnXC2Op+CADbZdobJxNyS17KgeTP+BgN
VGLmx0zwH2swGcsneKfFuRP8IaaYNIO5yGHSzZzsZAockvBPUPLQNSGwA/blbn6qWa69NhIGfFWg
pqA0ljOaj3oKT72qs2hiH2nNcfW4dyFLjiHC9Plo7F4y05gbTLI7FyKGoDW5vZGME8ZKG7AfyGtH
MO4Z51vhlnpOlUnnQWGGFR1ED+I5OJ7E6nJp09OLwmKGuizFaT/Ezl6K8EUo4em3LaH4MAmimUgX
D2tKEiio43Cidhn1O1aTNdAjV6xMB6MpNqrZrevWLdB0asw2cE6Kh/UMT3EINyYbnWc59FEsF8vZ
LvzzPyv0gdTN8z/3L09VSU4QbVI8J7CM32fFMzN/882n8HKq0EyJJX1bEzMKPalmG5n8yJYs8lOc
NFw7jShsPHSv+Ykl57IC3lCvosBDlRl/IAy+/PQxyxHTvgOtIyd23h9jnAPZDzm8WnuZRPOL3C94
xcc3j+HGMmAwzcEZzqmEv+TErrUCM8lHf8YboOl6F/VaO4D0PaLajo0Smr0KzP2U0OArNRUvyz1+
3xKWoy0Na8/V928JBhFlh3uodsV3gyDsULYEWCUUJggWcIMHZa8Ax93Fy5d4ZhlEvoqRg1plzfp9
48NNTMhLm2pmSzrRN33lcvtoMV0Fyh5GyFmD/13hA608Xw384PLca21F79Rv88Mp0BITDQhKIjRx
CeFy1fNU85JJXEOeSYBTXn9R/BUcvYjCzeJbXg+0IIjptSxYg7GQ7yHCU1qb9q9VlM4eQfwXdDZQ
myGSN0QM9KuVQtVdBsYGpWL9wtp4PDnCrjyfKRpPDuHBAQkCMUoG3SUNywsnbwJB7P5qPzjfQjcq
qkZ/Z+gKcC2bHDsNkGFMFSSf53NzZnf4jy5hcm7Q/fJIZJ5BxCd+Pbyqw1HJOTLa8JuLGTDp3yZY
lnx34s39BiQIT/rPR4Mq24k07yKmb0r9CPrQVVD5EYCRGBv1Ve7XUuo3YysNn1gXQ8RemmVltTdB
2dywHNpLTbxvbaFMK+HOcKo3qyH+atZBvRKl5CNBxZacHzOJ3zSyhlIsOXjAadJSMXHgrrPB2bNA
NvIybRxDmowik0yvCcctZ1ZAwS0etGY/UCskVdxXYTu6LcPiKy1YUh7uSZvCv29O3rASgFDF8W3w
wQby3EFlCwYHtVhV1yvDkWLoWhzsj52KMBKRzQbyRV+sUIKso/d7zRgKWjnxf0Pd2gSOqPBuXWoF
Ve5oJFnebaze4KHqklA1mwUYevZcVc7Z0Fj0xB4S2X/z8Qr0efmodKoJ03UtRYQSAVhJ/aNU2Oe3
ARZ21ErWHRWgp1xqMm/gyybKgYV7J9EJQ1JZkERnqx9Ej6G4xItg1AY1FbDUPFy880lg60N/Zvvq
d1tHlyf8BMr/jLdKnYAbCE+t+ze3oFka7vEt2aNo+B+F3Ub9Z+jGTneTnKzDgb+f0pre51i+4KPv
+rrtFVK52gIaE5+IoWmjkAhhK9VpiCG8Y8zQroEeXC1s/G5W5mqD6uCZrWc7k5vS/r2VezPQ4hW6
gYKMmljgwrBXfQfrAmz0UwzF8Ib45iNiVchYlIOhOmAlJ0zwF5p1mQuABBQDh3hTXKM9tXNvKBpd
M90jECSsRkrvUTTe25yLd2p3sN3CEeB4IeMqk8YKQOwRn4TQCaC45zqGiuiwm5eAdfjLkQK+N5XU
yTjeMtCkY5HTpMz3QJBDqQq+bnl1aG6YnQ/YD/mNubDgB2D4iIMPgfvfHrQIbvAPG+WujJgOKC5m
lsna5xBMSAcUN4pWdrWaeQqIGi7n4tfz0o9XmK7bpCdLb5lD+SqEaDf4v1g5vcDi40HvCjObYK5T
KcdH84jxusu/DuFwNExdwRqhUPxs794XW6KbxepW8TXKf1Y+JA2Ugslu6Z8NJjeuZ39qWd0KLY8Q
IivNQriUpWlFK3hBiw+V9Ez8Iyi2cmuyovcLNegGSRNVI+5EzM0JCCE4aNw43OS/X6SbistZcwZB
19XevyNe0UmKiz1WSaFmLVCUlIWtGwtb3VyYP7ex70lBjcMCA8zpuGysb/exv50xpQwG84J7vsRg
XpXcPuZ9Tk1TWiPeX5tOSafboYhmtMHHTKDFtE6i8j2yxfnVipdFGRGeyZ/EdD9ulZ+m4MRyC9NG
CpjOvk9j1Yw0VhpsR9Q6VLIFA2Sz0FzEy6YXBm0hS4wDrZi3p1QlSt9XgtX0C74K/eNMuEQ7Mp40
n3tbjjac6DEPkYSqyjM5rtr5/7kNCZQHbjuF1sXpuFWSqVLSK4XjEwcCJl82Ada15bX1ANN3n4//
ZhoEXfipQB+WysvfmlZ9B53qYHNUEEcWfClN6GOizSmGAPHIlNHbu0vnXspIZEJDEVzin5Rep06Y
uQaDuDSFoshM1kkbJHD2ABnmmJMGGdPJXZXojt4WBNtxM3BL2cj4h6klz0sY+Mx81fbOZm/w0gHN
BMMmqadjk9SQrsEcVOak5VZJBrwSfLoDTEflG+hdEVh188HJJoS5ER6WE5mJ777cy0qyubMhnzLy
3KYNtc5I2eItqHQhODgFG08ZHqMAL1huF1SeqQ5YbD1WUdv+5mtt9zhgXOsaqQmk3xXkYA7cLtys
9e2DCOiAoiPH21Td1Bxh8g78UA7xLQU7l6WcsegVkP/HfW6aM8fR1IPvIQ3aQ2mpo8P245QFJU3r
J7468MJc8D/a21ZOo0Vv6MdAS52uRw8qzvU3sDD4MMCtGEuFbqewYHdkc+AIUu+X4+bosLurGOKJ
lzAAUSvp+wE3IzQVk5IP5ewk7eJAvrarrQ5rVFuJ7Nj+DUCYfyui/FoEN8XgeYhe8nOVYh87/nzP
79KLSNQIbvkeheHy6z8u0iRST/hiOsFv/mX65uvhiknIKJDSDfdOvppA9oYFM5U+JfqnJf8kvY0+
1iuNDFOsdL07jJBSy0SeuD04G97ZNN/8/qgiG8/Vyq8B/9HU1WiUoFpfN9Yqcp/PzncTTIxPmWdI
EOEw6LhLWgOzZy1LBgR2FnXC1eL+RqNCRIx4VIwjYaptjbMAzw2jNasAIJ92RjaXjy3sm4a3SuKv
+2xmixCuExlU0LmEQrBpK09dSnzHhAUjCREPJBNi8/1clVbWGz5kpbT5D4q9uQPqdgkirwDmu8q7
RU+r+fV73Wa87blkw5eAmLBJ7TDp4u8X+NXnpSldDDI6aQo6v8bbLqGU+HOFkycoP2AU1FLeJccB
ejndUc23lpkwigTEHK7ecA85sgiZ1ccw/+29NzKDqDFrT6wm82z0dkRlhID7i5bbUzs0wjaNNtIi
tGqq9r0sOL8t4O5T0H+fQb+vaIZD0bNgAZC1r+ziHffJ4WHvJk4pRucMdSYaB58oEwbxHzjbfpL7
iUmTKU52I/uLsvT3sZ930D5rIRXuE0Do6iRt7Fj8WXDf+VignIencBKTAihykxJvN+9knM3s4PAc
Fx2zNwZigO8VhBt3GbnmwiXMOs3gi2RWZmPX7TZRwDSlvSUwW+7U9YydV4VyL3hFLTN/+2a1kXHh
Fk0p6DxU2XK9uqaPIIGA3R4QJ8gPE16H4ese/KP0J6d4a2nt1pEHxM25PL9BbOMcuHbkzi0r8dmS
VIsTavjA/Rap+Q1X1oZKNb3W+V8FrkZufN255p/3l4v5mPObu/jViTb2vAk3rngc6Yt6J3fQNy2j
Cylyi2Ro8AGPIaqV7SZfaoZol6EE5LkPdpisgEvPBWm53bgLEZQcZG7NrxtWMO2ywYiGpaWGhZwt
7M3/gNtnxljO1NBuAqqlAxvG6ykOjtM0z4XZfA9VzDWos6wddKGWt8nUw+KChS5FyuuhMiVvriJS
vJtqKocDXitSPApdMCPUrzTW85Z6oOykyrye6B1J+Ykm5o5m6PZ3aELskpIWOKIrH+Gvb/7UNyIA
ZPuIelT31YkjSYIeWpVpDTJ7v/swMcil1DF+avTJyknc0nTrJyNdxqkelYsbgrsL2YW7EAZJkoDd
gd9/d9x7NM5eD3dAO1qG6E0pUbatdmJEB8el08kgS9Nf0z75y1kTnznzI2ClNwkVkX5nRwgeqWKF
G5lpYtosR6/HQMUHEbSoTtv8m/O4+mSFEJWUumjsO0jhdeCZguJm+esXJ9WkSeFsvigGxf45pWtb
8lOEp5WhZxOp02wtj6Ejpp0EQiT+QSXNKyj8IGbFCNX++htjdUTwif36lN06e1zs7gqp1RHFNTh6
HTXp1jWcB5EPRNLuRbTnaOikfzrdNgeMi5KoFX+HLSRO+5WgnQeWg5GUl77LwVEoviWMquxBrYPM
Fsor/thPK6nQMJkdnF4CQoZnyVZw0r/YNluLdsSKS1p69+mK+gtYf56oxhkDsaXlGnxbjL7KmegN
dmWws2FKoNePI4Ypo2ZuzWY2JFN0t8CR6FU3zw+3R/Rznm07gLmz4DvAnWTTjlpDajMu+UOILNLq
PdLUYoJzIi2MXHixfaJEhKsF1S4YeAThKpOVnHDiNeoQd8yQP9RjHQwSLQDiqR9jOxJBWuss/pff
J/nKzAAR7+RO9Cjrf7qvCVCCqeoMZ4TXOcczFD6cECz0kDWWIn8mtosYmz/SslVaNmoNq2gxLWXg
/4tTPQA1wqCoG1LqC+9nRAFm3fJ+bae63RutAJKSstdxfctCvPDl9j5MUTsy8iXnx8KQaY4ysuM2
MhfWGExc34ElEVejlrVGtxQXYB73BxyHtBPRNBmXBNYSI3Aq5k6ioly6su7BJTHVGKbbYQ73VOwN
IysFoEPGfAm/vf4kFNvqDUh6J0JWvCpZ8H9joDPhZHXuZ/Mx3sTztphRj2JwrqYT1thKs0zI8UEg
7IHXDme2gBRS5XXlOHwEptdRXjMDHjMKi0ZzD4cWMu8GzB0ihKgaSgDitk+dGHmGcw4l65+zTyQD
6JnQMyaMxlPanMlCA7GsW0FBAmKjnWJpIhiCNOssHLn9AF/s8b4IiQrLvsolg9Iu4oxgX1ExMcMW
zYfw4LMwk+ATrHfK+rONd1lY56RZU22O6FvHkre+2a+mhrgMsjaK4sq+J+8GoiKQyZJTJ1N9pG3K
gOVaMN2eKkecVcHjUYF2kA8wCDIcWmaGDdbsCJUWfv9j4YP7fTmxadDEnFgCKkHK6PoXeOhS5QzB
Kjqf+m+NhSu4x5Ry7zzeL0Z86j9s0Bqj7ZfL+rZ3u+AD0vMRxdmvgyaNgX/ZQpx9DMO//Jlg9NQN
yo8SPRYNUaH86L/kyMJC7Od54cH1rasYIwwOFixu/tHn7qGadCGip+FvGbILfah6zF2JFR3CXV/k
apgBkhHzqBI22+RsV6x19Xt4Ob9xCRcMy9Ecg0z3E4GFbDFWrx8WRwTGhtdw+PUk3/UV3j/UqBYN
cTKool18/9lsY014/SwaCUIfOHgKMuWqZ2iU/2OnjLrrfIWdvMbWjj4/wW4J3rQeqj3buQKUgX7+
CDSmbj6DT0waNwdMkhSlXAIo0LoUYcBNDrrkfL3w0ss6K3DVPO8a8sZGszmHaTKf6+O/Mo/VdHRF
YL7ls2c+9vuQ0amIjFaIZ9SOARv6HEYBNQqijFdTPBfMtlzwK3zytXoAmR5UwKvF8dOlg3DJ3Xoi
Z5Rf3e+5mVBNMHZtE9nLNhY4o1HI+GHDw5/B36yf/URl0IF5fgXBglVrAncliE/BPGRy81R+PRgq
DfSpsCDiRW90Dh6yLhpAcIpnDw1iexwCeCgH7+g2khr2ug3gKF/uIiS3aKayzyTuk0k/jCoX/7aw
2jZy9VOgUCtra89uylfVqm6gXD5uqwf2sg/uZwGFckKKB3JZUjKp5nfcHaWJjj74aUHPtT48Inpc
rhACz8XSvaZsx7E4f7F5UVAmUEUX1fujkBd2ykuSt/X9+ZnyJfa6vRzKxM5PikHZYtno0JPI7TvC
wnqsyJqVSRzbk7x1eF82n+PzXPkDTbF9qTuZo1KEc0sq3+OkVhH+4MW2GqJbdcIW7Goq6SBuATHf
psX4Nmgph79d6KFthPpqGRLISV54T5wLMLbR21L/dXiU8o1oba1wjw+yfR+1ULxZtuGH4dGqOnl9
oQFnyopKERc+RlF/gRtEynG7GhfLaqzw0J5PcGaF1LuDbT1PQB+YIRbf0JKRnr9HDjYOxfKVt6Ek
Yl75UZUr/TAwTSZ7JQff42fKHBkll/emk77sngKFDlEvB/IZDGwLTy9HUpt+rqKM/YeAh9DbVfkC
+6xevlRtueEOVF716IG02dlTof76cR90FiZYVEbVin67uSp3UycGC50Iem6aNJIYPS7hRLYCUuCp
wZXXZj06jBrr9DcHJerMzHJfNB+DLrkfLiqwsWZiC9GxJr4NImu2Z0g4+pFo7Tm69kNF1z6NCQY8
nztTTXyho01azUnnrEmdIDm8iqBkj5Idh/zdUl29MdrtAV2uMu3NnlI7u6FJ8ooRmat6qQKJDrb9
LWJMGmefsjVNk63D4Lt3qVF5cKr06lU1/daXYeW85YGdJFGghzOf54hSp9gCR0X6XrDdIvKYYsCZ
zqBhoTIoOUY1Y7pou1MFrzM+ydKFT6G4ICH+nFa6ZgOFpVMVPMgw6aRkpIiT5pkc0CDZouBcvA3m
72ZihKB9EDzPbAQldC/b62oaufTSLt3G3ve4wnZyKvxTRdZGRs60tWPtOqTisKDIataEWbtRgPzQ
P3nwOsAnNxoUH0Tqa5tSQOy3Seg5WXShEKUF+IMBtco9XEVeZanu33okTF/Qke1+BWvFo2ZJgr9A
OA6yRXfe/UdkD7NXeM2AuDTp0oP9APj+PMf6lH70Z6YcbMs4jUazaWFYmmtyx8P3Ovt5xfCkBEfo
p+cFeMSvDjiMfS6QZJ5Rh2ISbmtgIyBELx4vjaVQV08HlIY/gzYiRMuK+aVg4LFMvySbM0/zu0Ph
EhQGrWHuUHfFmjAglJPJTCBru1sOfCbLU0c2TGKicbsFHod5YB1tTpD48Jd9i1CRRLQXZ8Hjq28U
xHG3pBrizEGKQnoZacbh+vHlcB8jwG51avVWiPxhtPvN/7xXiOFFatEBQs7GlSZRdE7yS1wfu+wl
uKTdUCEofD7Q7+Guw2BLL5CuhQ+kW9KV+gbWgVGyKmsbXR1OV492eOgaz2Lc6n2WMzFgHauOIT1h
toUJo2GwuZfHNHLP2q9oDWQe1qKHJFrHQQReSS1oQEsXgaSDGwgP60aQBrS2CpRpLJggwktuqYKu
j8WaLiwCYBmenn/pX57u8gRg3/tvCxL3mX1JTyIHVauKOIWxISHHLFcGSO50NswwzohPhBYRISgt
giJc+SIK2oNtlBAIIMmDBVsX0KPDnBxE9dkoZgCgWcgzWwEkpzcwFzb3i/orYpswhkAVIiuPgDDb
Z1LUAlbexNsXfR/AQ97fmE78mz1TteBS3POUQ0Dd27LA0tdP/8CL3RMwTPRl57DtvPmh8hlucDqm
TstAyC6Rgyd96oXRu9TqavyjEGeztHi5/eTSKdTNVQIR5sLtsO9zGCxvvSx8WhFo91v2EHucjR7O
xIh+LifS8ffSjPkhRh9EjutdDOM8MuPIqF23ZwjRhgXI22R1MNspr8IRe65RCTSeI/Z0HblXEVNV
mo9T3HP5uexW+3AL0peeqjFkhGTmdzt3AlB5LRJZsRgKS2yd3bZB/NQu8bw1wrxcZTtDEqqMFWn0
j7ztbU/fhLP1OMboe+eSb4LA7zshUZ4GHF9UD7iwzf8F4EQOEDOD+WbyNU+c2cZ/oaBtzQXu97eb
KYVbFwgd4l8mFAoiWCKdqWW9tbE9iL1/xrnIwknEs7QSxTjouE9XpLfaNtOkg+8EhiXNz6PJIPIl
QpgZqOhbw4P4yyUK7bj2u+cVfYrLbsMxmADCCb+QOZaAFJ2nD/i2slF/lcMHG9wAEWyjXch7RH6a
FHjjPdFSoLjGg+ocFPzl2QJnXuHwtCqhq3Fuy97XiOWYXyDnSezZwhKA3wWqswO1ZOV+iykwFBJ3
L/XLRnp8jTC2krfCwtALTQGrKrCjrwIUpZaVDE4tEbobB0GFOy+xRi9WX3IxishBehoYnlkHuhEZ
q0JVwmEurKRR2IfNBsuQni7oN0RARb46WrBj+PXmjiBAZf0lzk1P3wbaTFf7PldbPuGp0+LWVTPq
CIM/AYsT9lo//bEI0hdF/kXWFPlfnRAiWuJP4hcA+0edolVQgUap6kEdUPf5wyrnTEA5/wdvZBpf
LDw2zlx7n+mvHrRZSUnjqknUaT6s+wWBEbTcEfC9ziTnfnXNiFVpmUz7US2cbYaPvMXK0ZLmU4DD
DqofnemE4qM0cxenKD5hg0vWMgviTvGLOvSwqGk3bYqHLmT2OhU86btijnvycHZ5cVzScWIXNPUy
vYgD4bSduI1/PShyVnQe4IlvoopcFVUV/Pu9uuXEUVUz/0+JZlAS21O86xwCmVJVhqfDO4TW+eC6
YwcTx/6G0zBMczPP077rs4u+wc+Mx1a+su57n8Zgm4HTmRrrt068/WPkKtC4Vz9W0nu9DThVx9ZK
quX0vvjSmivp0StO7Kc4R9cb+4mZ85BMD977EC3O52eEjSKd8WDoZuQbvR7CWDl+oVCw/x1ZoWHP
J4ZZHW8rZxd0tFnl/pce9DNKYI6Ll2xTNdyq0CQb/yjW0gOuGSF12DcpVWKBwYmIlMdzW5hsWPbY
VgjlnAfPiMTb6Wd2sepBNkt82grsgo6XZ7yRAogQcjA7E/L4ddlnl1G50FkGR7FFEIEZmS0OXOJt
xY1AFnOP5KP6fQxwezHHhLsLQrk//4mCfdbv1r+0XmEeQ0xRQO6VDh+NzfkX8RtDszFE6CdwLkMC
Fs2Cm7qorYo0CCffyJuhemy3uQI3UOwwE1wkBnmZzZ6OElD4+sexH/sacY3lUugx9Nf09F1/SlJ7
pzRE+PEJ2nKwRXitTQO2b8XjRMsorTl0gGw7mKCbmw72ik4JKMRyUWo0ZXDhBHR/0BFRrwMLt0ez
qQLTyR+9EjUSBfrO8rvoVXzZ04piEbU5Z+vCeqteqrg2YNLv0XjW0V0KARnMa4joS77/2KgoFg6e
WuXroYnfyREeG/3IO0tkVAE5BnX9kEezOBFSZ//QZy4sFbqQmxXlIpZW+QH0xwxRPSTWj/svWBba
POrUo9leZZYA6ilGCssZonZUU6hWWho1y4j4Wzhc2ugopFl6ry5x1bvQvoLripB0dem2zWPlC57Q
7nde+VDbAE9SWXc5PkZHxi8+g5PHHCj3m9Ht6aRVTCm7lNAQIOlpZEpr/qsVbpIDRL0hEBB/Pn9O
GKc9HZ3gNJ0pH9UBpFyyNdlWIuPU0Hl3hyXbGqZGlhkD5f405c8z5BK8lSs9fEr32F2+l0130QOO
qdt8EHrGqF3jnnDHB8xgEplL44SWVdd3kQfCoTbspEzpNxhqipc2oU8nTaMIVeBtOh2g/p4Z82q9
qoKGx3ToKSXX6EpV+xCJhXDvwESNA0KyGfAeEt17UFHbr/uq
`protect end_protected
