��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_do�q��+�����T3M���ZC����	!�*]'_��0L��A�vT9����<Hov����Xj>[�=���u�s���!�Y�}>�i�	7�&��jْz!-����}f��*<-$F����I|�hQq&A��&��D��1u�wUM6:'��g��ڊ��fC��D��K6��� fvv.����7w�nE*�b����l��]�gI���)�nԌL�
ʚ�Gː�.�!)��#Ͽ$#�2�8��$e?%���g�i����W�ҫH����ƭ2�N|������I"�
fT�n�ltX%ɖ��^^��b�ܒ2Q�^9��ϒ-$��ڣHɸv�GI���K/�-?kUgHNZpw��3��k��#oRl��*VGW�޽,����A�C2vTG:Ɨmk ~�Ү;^�=ȑ]��y)�s�t��S{�C7v�M�χ�D}t {����S?^��_�ӵ;���*"����h�Z��|\�c5���7�C�&��V�n/^�+W��2F�Ʒ���H��/9V�ƀE���ݬ�w%!�N���ٰM�`? ��ey�hHv@�>T�Aq/%��ck�߇�Z�
8�(�i�r@�i&�����@���Z�5���Z�Z���!;���K6�ПDҼ��������;(-��Oy��+1R:���U�,@�h:YP�jn�.�S����T�Ͱ��*��&t�V|}��Ѳ���F3��d��>�@J��rrrr�O���l�M0H�5�]n��ci2����c\	-�h�B��&��d��^��ݹd��1rR�a�n27��Q9,��I_�$��L�w$�29����S}9�2Nm��%(u?[�8���Oi6j�?y�����θ�b�ΕMh:*Q�ә=�e�b}�?[���i�ȕQ��*�a��?	���7gk�k~ƈ�t[��jA��U.�����)�ML	w�C�������']ќ�=�M����x�}uC��x��	!��������(����Ə�G=��F��K11��[�&Y�ŝ���;�4�[0��t�`�+���I��٭P��ë5����c��ی���dV�K����
.[!X��^��r�h���),E�I�gѭ�,Vy)���K�,9g��&J���v�y��5`<���� 3�n��|�f�[�@����&�$2Qf���~��|�D|7wGUMK�;=�����S*�6�����d��]�svUo�����ʎ���+�	WIO��a���������EbM\U�wC��{'����𛻨W-jD������LqR�6����7'���I*�8pG_5��(�_PH!�v��W�Vӏ0F,$[��*�LQܖ˲2����!�e�ˣ>E�Xiԩ���Z)�	"2�	ֶ�fs'��A5:� p=�ޒ	a�^K��/s�N� r؍|��~Hz&�+5�rP��"&*g
�2l����8�ź�i��<?��d�j����ۿ�s�Ƃ~KT��|�*��/��$�=Kd�z\s�:��8��5����Ž�q�d����eIӟy��tMl��G')�{;����=T�J�\��2��ߟ0س�h<���A��Y:��yS��_xl @��֏���7R̚�rz]�e�c��P�U�yx����ۛ%m�V AK�l�ةE��S�3o.�:��t-϶�9�X=�H�"����w�/q�e�2��NQ8�n�����D����0�QZ�o��L�t¤�Ȟ�;�'����}�ZO�d.][1'm�W#Nz0t�?(��^�7�v�˼Ħiܥ�̣��G�]ͫ��L�󃂒�_/sO�^�?�������A���K�8� �H�K��y!�݊�J�2iTd�8�#���s��_nG�n-��i;������yZV�z��>L?�փ*�1�!���8���3l����F�䎾຾C^�?DD�6��D<�D���&�B��q�O�V��'F��q@�҃ώ,G������+5��]��{Lp���=����`g�kE���>8�d�J�S���U���}�}��>ts���Y�pV�|d��;L� p�{/�h8��s.k�[���%�{�!�Ո����-ڧ�i����m��G�/�N=�;9�.)߿�n�Q����[�si[����� �~2��vnޢSJ�X@o�"����#¤�?Ӌ�P|�dHBO��������F����� ��E|X�P�5&,����w�@ch�Q	��(?�W��-%���C%�?؛�����l����n<L��?u�H��� ���ck�|�HG��ه�M�0�A	�kT�Ԫ�OM'� ��q0�kv~�>���:��gW=���Y�+$5���#��2��]�OZ-�������ְ'���[_=��&���3@@�]����U'��ߺ�� �Oc=:X������T��E�h	��ϬG��o�;3��,�0_��9N�����mx��T�:�g<H+_�^0���1ث>',��,�F1cIM�l6���҇^p���,�M*t�{�D�?�g��לt�`�SDŰ�zi��q�i�%��!�fzr��z�c^�Ļ��>f��M�ڷ�tqU;��$�xܸI�P
��n,p�	w������T0�!�����&�T1�[�vP}�m��0f�u���6��9��<��[��y5,k��8qFp%��~�aj=1���2����ՔĲߺ��I�z��y��\�D��8���`/�iZ{���Tm���%R�����j����֡�s��5vD���"���1���n�A�(����e�<�62>3+�%��u�6�Q��C�6�J�7��������5׆J
^qy�rDvH2�a��l�t�XVJ-\�΀Ʊ��l❴g�"�w�JsA�FY�@{>��s�P���k�~�ǐ� re/19�k�5�X�N�hG�G�z��0�U=�;�ӟKw����o1<�_������&��P =�?���7�����M��˳4P�+t�H�'D�O�S��u����!�Q�9q�;&�9F=�-���3"ǋZ�K�&)�SV�;���,��3���$ʗVI�O���v�31I�*���d��w�m�mR���d(���M^�_pr�%m]�d�UNr�j��ɸ3)�����
�7P��$k����an���S��R�wUDѼr�T|���̎Il��G�	p#\����˽�?J_��E���P�V���?!8�i�b�
�YH��4#u]F�Fy�s|p>�5�SdEN���%^W���p"#�� �o_�f��M�����+�cDl�8�r�ll��~�df���:�+�vp�.�(r�p�� �1>��3��T�Q�o��_
®
W�f�jqWx.��8���C.0��wi���/�o�W��yS�"~o�~�Ly]��zO�y+��P��Խ�!��#��TK�ӽb��&;��J\����٦�$���Pr�PD4�d���R����dPW,����r�N�c<��.�:�NN�Jt���Cw�nf�;�8j�G3�5I���|F���� (V���ޖ=�z��������h�7�t$��}�^x�BC9i����g*�Qw��!��֦�)oi�H��A7_T�nCk	_3���J�b�=X�z�𘶶�m,Q���R�i�AqE�@{�א�撩�&3��;��a��V���	�q�&ur4Y$��2w����,�5)ZD^��5�ߕ��t�k!b�δl�$���t3�P5����Hu�Q���}e�]����#N�1!���� ���G��Op7$.F�^�8%�d�k�� O��r!)�k�/����%��\>���
��hB�5��b��4���]�Ă1&e�Y'њ��!�����:X���~����D�o[.�.
#�t�t�w�9Q�!��aOc/���]�`8�&��t�z
����"�P���܊8.yT�3�?^$T���B�380�_Ƈ 84'�V�k�e�Sf�TH
m�l�S��WQ�ՂJA�VjGԨ�I.���l���O�Bȏ�L�@I@��O�Gj7Wׄi8�?�S����m�R,���|��`�Q�O'N�BIT��;��'�㳖���hmĆ�s.��G$��1oф=���aB�\�g�����;��P�8�hl��*�7o�E����A�݀1-�T�H�,�6�ߢO�*@&,)��C���P����n�V7S:��S����Y�	ì83����f�a$�b8�V�ZTpo��Q7�G�"�A�p���