��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���,�Ô���h�Mk;wjj����=j�ˣgJ$�_����^C��j0|���.�
����!�f*�k�ׇ�B��������@�C�Z5E*�V#�q�m�}x�[Ǜe��35ft����7Yqx�����}-�/\8-byޓ}ڦ[���X���!�j�v�����,���Ϙm���76��t��̻h��jƯ1�s�wa&�m�|!8(��`��$-6�PG�^��x�oק��Z�g�4]/r��b8.���G�6��
9u߬S&��\��wd����쳖f�,Nw�s��qU�����y�V}*k.��]62�pYP�!�N,L�V9�������L��e�CB�;���'Y췎��rL�:�`4$��o�A��jR_��s���f��[}�%���$�!��l���_�����`Y�Uq 9�j��t�c3�m�E=�ԱY��͵�s5:��K��v�An��B��;7�Q�2��q�.����{�|�X[��<1ZCI(�od�K��q�ٵu���ד�t����2c;;��쑩of	j�>t���g���"�|=d���`�Y�E%�!؟?����d��?
�[L�=��Y�I�H��b��O?�%�+�d2/�=��u�{rХ�� �5�(��w�v�cw��G��,��f���>�L<��k���)U�'��yLn1^���_v����b�h\��tѓ�x��\
A����Q�OTbM��@�Ah����TE��L�,��3SK���J�A-�����f��܆a*o�b�@>�[���v�bI��RUo��v�k<C���&ާh�l���>�-t�9\M����zr��(��x*�3��r�쒞�����ޮ��\�}K��."�g��%F��Uh���<���rL�'u��'���x:`���">��n`��@Zm�=�&��:�o�^�d4��o;��q��ӄ��~�����
�j~�;J)�lI�͗s|���WMO�c�-gO�7J��&7�� rkݼ��%��)|�l��*�����h��W�G�1[t��xB��VH Xi��t�<�?�J�mR�k|���Bf�Q��nD���޴�o�O,SQ�P��N��n�Bt�?�7nÑ�U�������4�Bz]w݃Y5�����L�f׬H ��+��٪���B��8���� g�4�����KR�G'ul�z�J8(*!�U!��֟k6��	w��QP(+�����~�CZ��;*j�ꟋI2�Y���G��M�ĻC&W��K�d&�VmK��T{T���Y�P�UcH�Y�qcԋY��ء>PwM���#���`WS��$^u~���hk3H�ށ3�)A�x��Fz@zR�a����4
r%~���L�;�>��Ge�#�Ӌ�&�'��<��:3�v����*���0^�>�t�Z��BA�!����Y��Q��2�I����ADC.E�6�\ri�}�&p졫cVyuD1%<lP��i6���m��9E��;R�g��,ˢI=y5!35g���L4��aQo�ʡFX�N�#�@���%׷4ʃJ�)�^�c�su��n�2��Z��M�튧�HL��`ag��W4�>WB-� U�ۻ��0��.��ޕZ*�bBy�ۈ���������Y�4yv��L.�*b�و����e E�Y���i��]�d����?O���>�Kn�C�ch\�(�c-�a�2�/F�G7��fFk�p0е��?����msD�(��] u@�ܙyR��ZV�4v����e��s�kr6��z0�[���GzW�R���q��7��g�&&�_�m����vf�����.�3�jh�)��N�X3@@�B�n��y	8�Q9��%@]{W��o%q\��:@buR��s�i��!E����8M;��T:3�_Hõ�<���'p��ÖG�4#�c.=ݍ@N�]*�{pm�܁|�Ay��Xqgͨ州��iA$�����~�q����*�����牡v6g�ˬHxc�*��N��c���
�oa��鄎c���ڹh��#�ZJ"��3�dR=�d�fB7��5y��Q�g/r1z�,1h'�B�$"s�t��mfV-��g�|��r�yN�ªz����\	����xN�*�zƥ17p.](a28�X�د�!=AY ������Yͮp�M���r�Wo�点�i0�����i�o��z:���*Aߖé1�izu҉C�%ʗ
�`��8�Qю��|e�{j�@������Z�^Q�;���
E+��"�^�ȭ�_𬦵����͓P�<k�.ԚG㌠��K�ɒ|��X����`nV;⤨Jܻ�J=��i��.[�����H�����!�X_��?�I	�G;T�E�\U%�Rnz�$�
x^ @�W_��x˶��Kq^-=�nѾ��1_�ޡ����Vx��c��o�C���/�>��Xg0 ��3��rm)�'���/��P��*�@.����xH_���E�S��{RIei�H�g	��HR;�X�fA����گ�@p���GA��`�|f�����}D���kW[p����>%|�4K3��%�td���7?ͦ���9��UZ��?��j�EfQw(V�����έ�&�7�c�T���"ߐ��J;�.Z�"� ��{�&Ɋ���|�����U)Z��'s��L�7�w{>�,r��J�a1�