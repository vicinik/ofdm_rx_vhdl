// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.0std
// ALTERA_TIMESTAMP:Wed Apr 25 14:17:26 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eJsNR8PIWZg5kQ49RG4w0FwInOtGauqTcF3RJ367o3hoyyjKnbqqxgsWX/xIepqe
KLiNAHMV8pxtyR7pfTgtbABL7Z/v0+tGNRukF1vBpt5hgr8xzBeHajT/dJtr0Q63
E1VFG0lHajIiKs2ljkXRCVCNdmUaRO7WMeH8G7TgmEI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11200)
+QfT1eVu+BgiAW1UMrNvfBJk3WJzE+RcnOjxL0wuMgCW55cDaWZT/O8PsF6mjTFT
X4VGQqexj3oY4SO7UDHX0Ynqzu5jmiMfJtWmKjZejUQ3xZEuqo9MkPLBjgdYpPKi
L21jFx8U/pd3p3tQZ3vQFQwLngzB5dQ85EIn7m2SzKlCkKRYgbvOtT25A7z6XGKo
+4SQAgguAMWzVPIGw6Eq0VOjKvztYk62UQN2wBzG2xbLYyfuO4gESIZz4a0Wi79x
NVTnBDz+/aGnTypVceIYIyzzEavWuNOfYe5NmhyMnCmdH2SjM5hyGI7agW9ZVBtJ
6+Sjufk9in6W3iYbpz7WdPgGPubK2BzjpXcgI9lmUYAQRafbKlpAwHi08akfOwA5
/fFPAFkC6aBULmllej9mXTExKcQ+ofz2iLEIvoONeKpCy41N1GqKPWeY8Y8slWzD
iyAY68OEN2KGCuu365V0rYTU2JAN++VL5jQpX/NytkFq0BD4gae4Vn5nvBUO3Ha/
WaKYg3rD2lhsSSGduGMdzfqLo/W59xgrurVMq3+NDxYysOfj2srJOnSgcMmZixaF
rxJYZ04XNd/+uzrO89A74+UgYUefIms/nOeGS5elgUejBU48CrfxHx09sBFLSbNv
uynvtZj9UklZy3ooKttx9BJyeSmr0RfpMcewerhRbnYLpHJOP2q7OAi+J1nQu1DX
MvXyQa5QVPes96q9qflYOaofPG8npUg6FJFsCIxOjboCKccFoO4EB+u5TpnNIISw
S4SQqzhtnJIMcdpQBG1Pcjn5q83GWg51mesoJiJRxkj2AQYaNSGmZqDqrKnmgK6Q
3nzAU+JpOsaapDKCFTcfol21rM28R/WtTjZZewrb4Wvbn2/8rnYHmSbmO7Ncbbk+
u0qON75+XiYeQtii2/g+KGuwBsEsIzzDsN99sUFk+Xf5bADPqHR2XRRVm69Veqml
35tmr3dkzIQCvUUfLADqLFAItZtjzK3Hm9+/j8pFsf7cJ3bqSeirSKvGQB62Qy1w
fw+btM4L7u8ZLhgVN8pUwQAroFzdBYcZiIUB2TDoltcf9G1v8tvfO/tv+3bmDPa5
o9gKq2mAZyjV6dLNTt5FPBXh9hr54p1ZaDSq3Fl3IfahAHB0ZoItKaIyjRpb2y2J
BxLhrLgJEeeiyylpIwpmIQzmVL+ytxr6rZvi9d2tKZ2PL2kSqlbDDhobr2uxglvH
asL3JC6oqu9LhszMPCPCN8B675gnW3VN7mXENj61MJNDaGyuf4LDar9DpJOf1xEf
e0Ixe64a8YeSWzMhbP3DQ8ZqzHXpYGzHAzkcOwLNrSRQs2/DkW/+hqqFslpkh999
/eBjcgKg7r53s8BfIBMj/PeB9+etrnhjNpNTAp4ipyTNFDC5Np9JAo5HX72xorRi
ZqyVCVNqP34NVL22P8O0WYRhOthedU3vmJ9x1buBqlOl2Y1lgpiaumOA2VcT+d12
09/Md2GSK84TN6rz70PoiFV5SQUOhxBglXJ3Cv7AgpYMPtBJ/EduiVlRQhbLxAPO
0LnAgkYE+6+1zGnXjWdZZ9f8Itd32Ugkv3z4Kg5PovmZyLYxZPg0XHNJGavgJOVw
LMA6gyuu+Qjm0KGFEQGiuouPSBCCGjK55WW2QQ4QWoqqgS7r+jWpa9SAWvrYsfT8
yJXR4ih/XmwhW9sVLaYlvskIynM2+YFY1D4HChGzf2lRPq7BXEhqXZ23u2uaz0XS
q+b6NYqHXCe/RPgxRxqd3q5NXYbPiyYHxiI7DL6U3UKc4k5UgFQo/1+CGsnXYlKM
AN/9WF6yfTxQf0zquY34ihAJ9W9HH1xpS7i3Rqo3MCFNY+y1EsFlUsuqOadGC0t4
IB0QTGvsEmqmqaRbjrn5D5dVGHJ3oL39nyJIEd6JRqfb4yPuaY9W8ec+Ax0lvqE5
3I86x9ZC4aC5mzHl+hWUuPuvfuQhXc2x8a8Fh3SVuyuweZ4RvbDKsoACm2HrKzJK
BCIDf5xKRmUcF+ufxTm/FSpPLdGhXFRpaLk2CtDTOudFu962nkwK5HQix3zVtvz+
OQi+YQN/6qux4DfoBcSCL6cd/pzzoEi/qub4KNB7Eldc1AK5xpvDRTrlQgAlj3q1
PdLcKqt2tOnmYQJxo/abNhxEq23jK3RHxVF9rPqHEq4kGNBIkBJFnmD+fYecIlp3
Ar2Xpo2Moqk28osb4r5ThV0xakKczd9F6IWWX+u86iZmkbg1FN9TQrIa1PMg9ugg
sGX0n5Gi5r1zx3/rawwUidJc5/vvPZi46URDJvwNrtJP86HKGGrgDZiOOs9Q+8Jd
iTKlXZ4lx+Yv373c9IGyEcVfpapXrK76oJsr9QTeXEtWlGgHTGkj2WRSZUMVKEHB
gIbRko8kyqzqTaAdjvq6pPi551SNkCZ77mu2AUshbBIUtFKe0oqRieosNgMPmYBM
KKsDRnevY6o5qYoYU59apqs/J7INdD1qqPgvKJ0Y/EwqN9OIhuUBSqm9g6d50jw3
ckJMJQGyKDf8QxC1JRUnEJQjWiIlnJWtWQnTRy2qpioLDIScqpRWWXrr1fwZw9ze
KL3OQ8ng5zwiZbVtHBNHyK8Yptc1jVbxwvos5Yb5vVsLRcPRfBXozq4Wk2bNGTrx
chqdU1+11KCDvcXz88CrG5wx6BNC2hN57oQP5cb2uYEOCJn+h36v6+/1Dv3A75HC
WWT8WQSnPY1u7Kl+GD8tlbeKr/t5rjBh+2p16g6+tK4N0l7+C5A7IzzJI44hfmUq
XW3Y7gW8Sfv3/NBqHPaC2bJzFtyUKQtgr3pzvjaT5FmyL4q6k9+UZQALECAxSW7U
RoYklupoWBUdnPmc66U0fIs/OT7XuttP2uLXox6dnZNCZZ10llWOSzABboEPB7wa
GxZVfJ2Yeb+GapOkSaF1s6I4VhuRX3YBCArO9C9cOmun47Rgq9oyAr5i2Ae5fCr9
q+a4ogXCFPd6mCPm1mEmNpjhMgfZJRuSnZyNp8rruzLPbdRCp3QH99++57uJleN5
O3fIH72SMksEB9T24RrNLi3IzNi8yALHTb8m6Y8PB/oOIbmf81weLkgGMYQs3KhX
FbKN88RzFxUUf94AChwX+KT2va/f/FzY+Aq8sPdgoeNeeU4pkPZwUr7MW3DNnTYV
VLWocTmqCnQSbISJz6hjBH8a2BYozHePIj6s9WHsWNOQ+XHZr5Ky+3z3e6sJ+CpP
eDjGq+5RffHgxGLd8wBI9onb/TCfARtKcRGuT+7IhZRJkXBZV9hYGuOEQxwC0X+n
uTDcqdtvAxKiNg2dequZJriaUfcDhLhqiLAyjQ1OhqJru84iCXAviBikRxyoMzpd
DVAPzj5D3Oy/kuG9rlB7+s81hCoyVh6MlWELG/WoLn+olpnZbksb3fJwzaLbo86Z
jQVGkjBsruCrPHRR3Z2UgWpAmBn2jUz8gxd4qv/laXSVkfkxrEAzZvv3mTJfmthU
GVRdH+ekIDc5WJes6QEDcH0SFf17GvTP1hCiehKsg/bDtfxn//NIuFsqlzv+BaG9
eDHwp1zGBSqamCBBo1h5voIyuuGawPoBiC/W3JhaUkjK3WlRdM2jihZK0T/3Ys5N
F5iqv+9p+7NTVqaV8A23Yhjc4v75L5NXbCQgxkFKXvZ4BsRg598HCypB2dXtX0zs
NZinO7Kp8zIK/McQFfWR9ZYbx3LT0W6Raniz8q5jfWS39kH1aeYHJA0RfM6KTggI
dcM+zu6ID9v8mS85N7VHOfgpUt02XgNRnWjum3mQz7k21eRiAnoDtIB6TQDC3lP1
3ACf45YkJrMUhG9H0fx/wsxBK5Hu7fm5UvSQaryDQjQSt/GEyDqkqM6g9t8WSkR1
S+hkn9OPU1zGAXSQq/LkuMWJuSrmLVwNYwaHAZGsx674g7Kf6YDEfvsZpG2Tdv3N
fMgheGYxN14XBoUz3zo7sn32LBFRnB4h8QyFhb6Yx7oEdkFP15XzWnI/ItSgGdtQ
yBIgHLj/XEaOjD9EPC9w3zcC+MgNmvmVhaYPuaCof8LgM9H6WFAcdFdZ2mtHCpYB
N+tRbQs+5jhVTWeSHH6mvXxbg6szPN6vr8ZHSGkeTCnIA4cOkBgsJm+zMmMXRFws
rQqrwZ/zxS4LVxliks95xXxOawnYZkHrTyMREdcceKEqFMyxAbgt0GWkHH930JcU
XrAGeuG9aa2GY40xpg69i9jJ706NIAOPU1IacLTqxGISOg516fOSQXu0gOC1N9Wp
iYpt1yhngfx+ZpouRDpSqpWipORE+zXkt9SSRm6BKyRvD0oCYn44QBQsURe2gfUg
zGdnbEo9aReTJMdr55Mr0sTxMYjqLI3eSPMULYOA0m+isglM5ak9XcnxcbKAdxPH
G07KGSdB0/vPpBs8pph1+tF6hnJ21+eYxNpfiFyjQVLGtV5UJldnoauPwUIXK6A2
mbrO38xmoCZrwotuwjAUmjD7xlrpkfGJM6R5jIJ+XanoW2G6AzlE0mS5DJmqbzhc
VIS+94x30JK1/vUB4NV/Uo11LqO9+BNSMMkYPEwfkY3wb6bK4e4BxZlFvN081DwF
YKTkgN90SmwaO7wjf1XwN+J2Hye7w+EROXClwHKp6MW2AwptPm1zCU337FOVPA/e
WIGuzYtcNuydRn3xgNaP8Ffg9/JMctPrzuxZLZ9D7amnzw5474Xz24r9FRPin9Yb
gOn37ztt3Qf5pAMx89vn6QhnP4vPOgYcKGGVZe/4My8+UocooD44tSHPW2+Do+sB
dOWAGMEaCcGVEiaeQmGufrx85GcF2RckHE+rtSLgeqjdB78BD5pjIvAK1BmzjdqR
EMXtxrNiuGe9+9vdlJpcvZdDWS45JD+EmrqqIAbHAA5aznhKn1ZVanuLWCQ1XDd1
v5k5FgX+yjLe0v6N7yYyMvOrnSPxGQK9166CykjWLHmtmPfTWPZLEZLx7AmkAyC0
RbkWgyDMN5QS9o76jLGk43U3VikeaoFdhCkJRWeKMAf0iZxKndFzPHghShSf+jbo
nb5URvbnVWb6pYF72aeCe1Ext6Nehyo2jwl60XS+F8tPJsYnSJfmmWNGCnbF8wME
F6pCz5mXw9gGwCsYtybWMek9Pen2VjSM+yPjTT9Z6TUm234MD9zSAelKd3LqoiBg
J9HLLUEXc6i7J2WggXgdktxgyIW8cEMu/EuqbtOY4Bl0BQxYaKlppcWdkmKxYnGn
6IEzDyWRenwML8RCWE9I8YCiI2ngLU01JRpUrO5a7i+u+oei1c+XQVdLQZ8oJ1Tj
wwS4SahTMRaPKueDb60cysn8xxK37agUB8CYMJbBA8og+jIToGEU7qvSOEOMGnJl
SLWa/3cylcjeoiIZ1qAvVSxfJBx39Cnr7Wp7Y0ftADKP+HwFKhjYmKnW2c6/xbgO
hUGHJNbYaKKBha/aBHtIVHs19B4eNHTvy6k6yNK+Ffku2W1wt8drHB8lRacsq/yP
wTf8UwYOYGo8wdthiJxWs5rl8OaIsSymro2zfBxcRRvdu07f/piu5h/fprmLErNs
qLESt98Wyt/kTKUbxxeFLe+U87IaIkR95sEgk3MnA/Eq1F32CGAMKZIf8JPzFGoC
EhqqJPDaE/HoV7gtZ3wSh7neaCShv0ynzj/+6wKg6k5ynzTJY6OniorHaGXHJJWz
rmGC+ge7QIGc6hUjGfuXmhPO1GzvMDKU15uq31M14UbBNleE81qJABJPt+ymO8wK
zkLKsaCLwJud/BGiEh9qcYL5z3Uy5hTAJwZjzqFxQnZVza4GeG8fmmB/IWDuokrQ
mSmMjdjkU46BkzUh7GqZ0ihHoR+wEFVRbrAklJLNNA6Fm4q9VGUX7/mgo0bCfOOF
WBiLpijD5avretGt/VM373lLZSRJeyXTaVaex3fzZrK1eqwQbhYN7t4zuVMR+7qN
VF1kamL5zL4zt+m8nJRNf8fGc7mT0+0fR9NAy9W0vk3EbYYTLIh/4Yee03EAPkwv
a+QU66LANvTWJrLoS8ZoXH2YgIEBOlB9FKUCCA8S8btqE5+d4GGiMg0G5ijrv67M
sVa3GJYlWSOoMZi6+4WSq0j5VROXsPapYBYAyGv5kD6d1O956EWLyTupTUxLusd2
DtKjot9OE0rgB94f22JK3fxxnGUzjv725CMYWBTyNcDxHkx/c/Qho+nODraQOWLv
jH/Uegz54FROnAKLcyvVoLc0SS/pPuMQkbcSQcnSAR/ox/OYsMUxM0iqirgzyg6U
ObWXx9IdzrXVwxpFCefs0tQ6xGum1bsthn0xYFkO9C6hsZc9uFHrUFQz3U0J0VA1
9vID/HwlQhH/Do80pr49bkQ3mXG9UOjlWyPLUEkfTe5OfoK1xLgHV29iy0xn/4Gi
iXC2wm41AdTraqhdYpyUuoGttOz6dj4RE66rIUqvSGWLBFP49hJyk+WAoxJRqIjQ
Dcm4e6ldCnj4bviAN/H562e2OzLSBBz1Ro3sAvwIk7LkXHEc1N1OEh/MX5XIMDkK
ZgpHLLr3Gwj0sDPwIIhnwFVniYO7TZ+QNh9+QTdFlom+SJXApD7MbfYKcjMbceWK
7ql0d3DkWFpQp7DQXR/lP7HZqBPax2+yxaB3zYTCHA7bHfnqC3sCgOjPHilZ5RfG
sKvmhhQGG2Bwd9TMLvOVvZlRRUiDgB5tIow0MDwGiofyI/0whnRT4kyTaiTaiE/O
XpToSW1/u5iDeVWcoC2V5dIZHS0NgsHDZ1IC+aI235VSPQAFACe+0oCPU/IMxZe1
QXajBSxE5Rrq3SorJS33SPx8a0TjjZc/vve6dOSEM9LUQQ5T4uT3RFsxz2UjrTzu
Xqsww7RpO94lYBHoS4lLhmIeRHpQNAeAHWJbiH2imE1FdA7BmU7NgqWZ9CFCjEFV
P94qecdxiWhBIBbpizsrPUJC80wGVfSKi9DvMqWGjEEDSZvxLih5nIwBNqVcP6fg
eQ0hPiDhp23qtj6CvOrZ79dVRNxf+a0VXbsJI36YNBIsdJCUT3XETjH0ewRyQyOJ
UjSppB5b9j1TgrquC6fFODDoGdJWBoU1w3StayzZpPcnuCL78iX1T7u8xECuFWQ7
lSeaUEcide/Myf9mUkroOt9ZF+aNAXDIcpl0klCSSoLMAfd+QDvQMQajveAP4l65
BENU3F7UfbH5XG4Trm13YIFxwdZR3H0gIbNms/yLKJiiHuUtjqa/oLMsLjirYBpE
SIjGy1hg1RguN4+Dae9KpisbV8aqqx3qUXwCQSJIn3Ynm0Wv7PF6tpf8I+EtApnC
XwMBbx92DM327eLhFFPJFb3W23iphCsxqN7S+F5sOkJ+LgumRQYYQLuLCMpXzQzb
8892rJRYB4gJiunFnykERegZ21YDI/Oe9n5CbzEFtmF9fXTbGPPaJvLdyzs4hXXG
yOihFXJxobxnnLzidTQ2A3WM8KJlUd/wf01tRwvbNUpdzvS8z46Y/8fu6oVjMGa3
wrAp+LuJ43jfFw5nnbPhIMSao0oEQoxeSFLXKjKFPNaT84GiABGqLWaSSfi0QFGn
+nYqbYcmxk2gpR+3/II1JQA4QNQyyyLU2OfbmziI3xkfFwYYkJAwCKlsnHExYDG9
zL4uvPFxQzhP20e1b9W3sAX4M5jrJUVP/U6gFYttGohla5AwDOgBMX3oQMHdTXe4
GNUfyR9VfvzGC6yq1wTsYf3nKMDqlxmdxn/dL32lwa3v+18qaONhYZUquGyaVyIh
D34ko9e1X2APTVLCSc6dI21nuvCm3vzdkqjO0q71+3pYs3dPr0LhWG3TsULmurWz
r7S8g3yE3BccGCTzW02le7v9M48+XGgdC7haMb795DohjDqoFWH04IGXQZUtYbWl
IrksoW2vLOt/hGxg55GHMmEwwa9ZPo4IqTHOevQH9kgRu4rYd3tlbfVXt5SKVdC3
f0KlbbngpHJzl8vZf9kASt2E3euJsAX8g8FqDTgagiwCoLUQOH93bQYYqMzG+6pJ
L/sWaYOkkrMysIDNNs7Nsv2Ai2qryNbr6MNWgwlp9f1zCdkfrs12in0ckuF/zFC+
BFMRtK7svnaxeTSk6OkWPudmgKE+muUCKEbMhxND3rNa3CM/NEeQiC5sU2/rhwk6
myl7+nqmFn/nj677Rga5rvHw067qbJWMee5RLJYIxwKUg0d0p6AyOmdrimjAqNMU
vJV0fMn0laGJX72/qiZ7yizplP8rx1tkk4LhvN1+TaO4oSuSEDLqSCux+YShi3QC
G5YQCxu/5dywwxfFoasK9eoff/d25mJVs2ijaVa50Ln09SBm80zKO/bZ2bdvkjNM
OujkQ7cizN990aMhDF08GO6pf4k4UaAyY/shOYBAhwtK8Ztbi1l1pCrtK8+A58cM
9vQi2qk+YuUTB69HNPspkI4T/6eRT9D9B/m9zEzfbrZsnKtW8swas+iKJiL0QdVF
CiiSXF2xt2nUSM2rhP5HgWz+ojIrsO5IPrGgJptGfexNX4iuiqmdiY8RYHkDNYXp
fRMVLMZi8KgoqFKiJLkztkja3KdiR4Vz7LUQsO3pRtOsotNUsP2Yf7EyeP35xXBn
z/EkKRxwvKmavU23PC8qXGfvdH1lB2wl7Rq3R0KpUz6j+662zfOmS2D8sWfIstld
1fvU4XqSLZDc32hWGM7jO7pyAC0XXfAPXhVtt+fmNY8pTOwYXm1+Uj2pRhp2h8i9
i0LcapnG6noDWJ+HJNVin2xAZpiq7wLpah/Ux8lxa2OLM5cnKpVeeHwfV4sscNGn
aEJfZGFo3k6LK9TK40t4n0HXb+PqGH72a35H0kiIOv8EDoz26HGUKv0PEwtL2/Jp
jpGPyhlwcsQS2kU3KbU5aIqrmv5M7z8BcrXxgrvRcJ5H4cYSQ5oh6+6+wHOznmVk
5KM8Hx8JyP6Rwh9a2UfwaQP8o6vm59CfCFTRn0mE4RKjfvYRqrpmwU7pQ+sBnumo
/IC/nw5BAZdt53iTTNEIxLmP1kKnQ0RgbBOTZdXFhN2IseaWs24R+74d86801jgl
wpZgsxWRFGInJYD015m7cR5qGlk7LAQO5QO9z0QOoxieqZoLP+71IeLguwPO+Ql7
YEhzkJEULf8AOnig5IXcgFxGQKHYdZjVNHR1/p3WmXaIg9jUZVnMyUdloOAPudgg
eMukOP3bzqMFo83Hh3UEoZ+9s/xv4sbl7MgM+6YuLG07QehFIqmB+j1Z2baZEUtI
6RXZVbqmXsI5gj7GLM4VwqhqBe25JZuCrWzHR1RQaG2fo8IFFCC9mvnlyXx8eZF7
yrffMmWSw219keNUBbdGatEDBGgQ5IzKkQff84qZDZngclWwV8tdiPDVYulp8jM2
yS6IhL4Gilya1BEX1kIEL7O+7NJ+M43gTISnt95QXGb+4OlIZp4U5zUrGLjPY49g
dZMRSMahdXOiuiZX19XYLlrEcJ4a7zGi50dm6Fzwbb6Wy3ZekSM5bViq925KZfyM
vAtHveetApIpG9JeRhlZEUXGD5P38sL9HvXh4xCmeAC0ucajSiNtLh7r8dn+O/no
AXvSEWrdB337ghLzuu3wn2UvVs3mpJaIcIHQ+MY9FoVUnHf9JrZZ/EAhcGXugaJA
Kc6I2EecWu4SpDbDAJI6cXiejIS8RpMp7EwOhK4Gw0yZpVbdWQmdhcRfIiC+7guS
IpHxcjG9chvDqDbIQV/BexOW3A00vs7pl4zPJ35Con7FZESgoqUabnrKn8zImz+G
9NejmVIIsINl8PI71E8Id9xqJEf+7atqu16NermZhcnLxR/tS9p40oa6S2Uu500W
GEC7kYzL/t3w0CuHOTPK27YnzDtG5+Mur7Bv2P8W+kJOzbzhwAYNm76H2BKjok4T
HRq5LHHc+i44ylBrtxcs3EOwycal9uLgVZ+h8iWug3stkit3t0EZa/1CZ3Juq0yj
rklSqDjoEjdOYcDDWyFODQPie+3r+GbqTGtFCNMOtk6EJjcFvDhF0Df31XmQjpOi
UTBLIVBYnD61MPl8hgTQyPdmVvjw+qG8j5JrnOS7Kn3CzU3/2NN4C1/kdD7u3TV0
jTFLLiALNpI3slXEfiMxgO9WDocYJlsfB6h4Ghrx+XCUeu7EwSzDufnYbNnvvdJw
vxz1VP5Eg9IQp5idzHqJqWOGMQDS2C5971DXRdd21cM9SOh7Ge+9aI3pS1ZooEg5
3YlXa2jAjtx1fGRSk3h4gXs8g+Xrg69AeyxvU9xjF39leYw5zziSKhDRA84Oo+pK
wsJszu3xKj+gd2On++6r3WYXBDrd7jUkWXq8zYav1C9xkPQumfQPlTsHW4QIrOCx
15Da5ZfvYxr/eyOOk7hH4Bk/4Vjl9qB1K3s6V+l++3vazXBdVU+FMHPOluADWkTv
MywTAUj1u4qxqTfzqzodlu+C6gbUNhUaVpPcIhCOGF062eG0pGl0z25GgwjDGCkr
hSa/YbTsSY8yfCtRq5zL1DaTDx/H1nCk4vEulkFAzO3iiuuOjMu+QMDytQVMKrup
5Ed+sgzykr57h4Xx0CfYWcTK1HUfgSdbM85g4vbxIBS7K2576rKXso9V1bZr179F
gU+1UJUfYFhiHxCb1qtEbCN/GI1q00sb3x1iK6U2XMSausqyppv4PRZnTGM7dvkL
6aJLY1HqotngX0nWCLnj4Fu0q+hF1mZZ9/OEeSuf3/Yq0+hIHoRYasbEWhwbxw13
JWCV2PQ2ftObssZ9ptI4BSQLbIJ62vaHmapA1PWwgyRBLeVtbFdUcHBlgfzNVrNg
pLru/bso5GV0xiMuSSpid0n1szGnAH6Z5SqOScPRYJ4skF2OPuAyj3EGXxoz3ok5
bxyStCZUNSa0bKr35WdPLt8LsGGiTt3jcw0HIdwLQZ/5UexNhM02yKaL3tQeATWx
UtQmgvrGngazloIRlQk+JX6zXgKnsndntrxyNOyuQmbu0zPibctbVXNYXgp+8+fl
XocoSoUdbSa1+j+KfrSqqFQquWoDJ/qpjzWx71lpFrbhlGcX3zw6OWIOvy0+3bU8
KBvt2RyHMiYQBPvUB+YtBrSVspp9h3FF5dPjxyzI3yPdl/6vYWrU1wGovXBiI9sm
9g/XZ+k8tmQV/zA5ajR6Ovi44stVtBG2HJaIlgIQD9pLZdFyV/tkkqpODzsCrIE/
dYi18YgCekhOGUNGrWrABwN6C9PlrV9aayFYU0IkEheQPSqjkBWMjZArVBY+Q7iY
cPqMtEKT4IgRnVGtRazDwbHJ8aL5zXACKboDlngkRa5+1AWkRf2cWQbQsBCYYmUp
3Tt0FOYLM+X4D2ICSOAVYDZiaR857YqPs0SQ/VIeEB4uxERjBbt8Pfj1vMJz7qlh
+Z/LzN0jizxyZTgJlaD5VGw+Yzjti7KouKSAvEgEytnlN/hEeP0PA4Hn0zMClViw
rX9/ONkA1HR+bPhRPXNHdKhqdaGWmlpJfdRTnBo7h8SsKF1iK/THNWcrJrB4k6Pz
9n2IaWt3j6lWJKDNChFk43pH7ZvAJoj33LXwVtK5pciFrXVG9A9IlRXit1B5il2d
bMYyCAWFjjMKHdCaA0lQzDvVl9bKsfeNTmS29FPcNN39CnO6NfVGU5PQYMbdoNGT
q7y+NflnoMitb6ntaKxifFETcumY1KUI0yo+o0DOxw5IGvLp+XedKq66VqunEX8q
4C4MzNb3e7BsMBq5Q7q3bObEovWsaJa6MJWz5OG8ESPv3BVWWoBsX1kQoKPFRgnO
yVvHGyOACmvXX2vUMKwLyynQSpufwF5lAxMYnxqhbmUXu/dDmkZxf7jz0rLbOzo4
FOll/Cn562Z5p8zlb6nE1G8RlauZPd1bXBVJVh2PBrNhZnPobMn4rrLZtzQAeefN
6IlKJu92bNykSLPaPNHU1Q9Y0+idL7xojahFPj9VLRB35zS9ffHXs4Hk+uwa/25M
OEjo0vrAx7DUE1jl5K57/8g+n5FMwokkomoZbp018ql59f2hHt1UjyBtJhHskm8N
JozMO25MDJ+oZJNJzUiVohzOXq1FGUAOFq6QvvkPDv0D4x7y5S6OMw2UcKA7sh1V
Ty1GM43PUrVEW2JOxsnPownyiV2oHHuE99Ije8HRjVMpfChPa3cqxzjpcDO+WfqM
wAXjjgwHbYm3O3e97bCi8QtDLY0/xBQr0QxkIyjfmJZItELqAQ7U7ALDVqR6WmsM
8ITBvQnv5Y1UGbPCNsnBmOGb4KT+rNk6YMmCG3jUfljcYFVULc0R7ORoiUZpes00
QggOJUTt8ivSDu5QIaUfb5TFY3mxyPI/ziI7jiM3swzspxxiujp/+/99HeUtCe9/
e8bLcJUN3a5T/sf27wNQN2BKM8ePeNZsU9D2wago7iH85DOAEvpDswFFOviFBD3D
IvwI6AoLBc6bgnE+Pfrg/IGYt5Ra1BuMHBHNPv2qLkdDMqLPlhwsQuo1LkgLMNHf
EA+hnVVig/0xarezcmWyl58hXbWDMx45ae1NQ3bpiurnPaf000hJD13/ESZaLOmI
yfd8YgdrYcZYBZXXhHlBbiWysLYsg2B0Nm07b/g3YJkUTZk0BoH64QXoUhxEqKBO
eVaAFT9/B8RaXBLCEozlDjkqUYLJkaFN5Xl+KbHDN08YkIQuZcLvq5x96KHJ8VJz
e+hjJWy9FSFBfsSf3dxqYUdtVUxXw7qHD+1QVg2h1W+meTpE9irAzN+Hy3a3z1/1
bo+f2c9ArEOPIb48zfsKbBgNjqcAXIsO/VEkzObRMCzvKIoE08UESQwRxQLDDBOy
2NYgP5WCuE4APrAvLeeIQa+JUaiZiSzxAVDv7/zQ4bz7hEsJ0WXvWJ5ZjSUfJ5KX
zwDrdsUtOs9RSukDdlaJC206DxrXtRtnWkRXxspt+7p701BFst9uPlWrfVbiLFcb
LH1u0cnVh8USqsinhqPyvYtK54GEyrLMBqJAXXmAxYObKMzUnQ4N7Vbra+Ns16PU
4Klkcj0fj6MxA7RF5GY5M47aMsUU8es1Jvy9AP7hzZYAXzutpjttmstLvFoAobRz
PEx4KJ/ry/1qfaLGPLrTamT7gnMve5K+tSr+le+m5WfBjCcICUbNCsfz2P0c2gEa
//k308LcEpNZQBLImO9tiOhNZ0/FsTuSU25TEnnSqdYrnQE6qSaS2dDhJSdoPNyK
t+33pIR49NZSCadi1/JVtSQGYP4aqL7sZkT3R3pKMqdVSSUYctRB8+l4v/e08Bn+
uEuxhKdug7YItcFTdzpaOUr/CjAU47TO4mkuTFAac10Aogo99PFBf4E5fe78Vl0D
lXX0qO48EwYWVpR3UsaKyPJz+LEUml7SJz6jeDIJI/YewiUSmOdbjpnwuXMQ4qcl
qCmrWzXkM4nT2/Zf1+nnKwdAdznPItoeUyLG3jqISkLF6/0gaTa+NnTgabWJIo6w
d21QoJTKpvBy6pAho7X8SuQq7MjRFmGZd4BfXaIUzny0F3+U4cLLGisBIxsPEJs8
bnrwlHsRoO0n4rgQd6xhtcC4BaQ1xYLAHSvzl48mED+Av7RP95uhoA6kiygOGn2x
JZAw/gqIeXYh+pX2piiCMj3OjAwvrz0ipCV+TnkdryxR+rP8QwrvO/I6ako/h+bv
+i/nNeYqrCkr3drocygtsjqVnMca34AVLJ3IJ6cTjh7WXKGOi34x53aTkSeKha0/
StrdeKiCw7iQIAQAMghs3RAcZ3Re3gO29JIdSy9TKT/o9Mgg9S+pJft52FcXflLb
/SNtVNkKDDb90+OQzmMzc/WN9CMBLpdgYAGFMD/NYAJyb8gkCQ1EBokFmG+LNrf4
82RR0TkHC5FyVcS+1tutIqa81K6qETpZoHzCRFKEfvdPlFI5ApPUf8+QuBO/dv63
j2hNZPO/atsZGAOnruFYPfhNmukVJ8Az4ugUp4YgJCZAiB/b5smmmu+pshC1jcpd
Yu+2ObwdGkd+F+j8V2YRskbKfxR5ERqsoRQ5vtv4q2F8eBnknWGwrH0g/yeI3o56
lZuT0av0UIjgV1tUuOgkolmM+lN4MRGUZMSrMj+0hYl03hmT+dkO1NUkjPj10f66
6Z9s36yceVb0w+SRqV0HlDVlsEjkQnuFW73AJobH/r9ZMYpgi/F9/7C7TGD5e/W7
AXcXECW9A+BL/d3egJ4KrPKcYfUDGDbsLrFCe4bdBNLCBxFxwcJeMIgmepk3GN+O
8f3UK82uH3XEXJC1Wrx2csCgqTapaYBROWj+xe5sGiIBo/C65yqGTf2MmKMeKs+X
xVHd4Vm+HR4dLKT5QG2PmyQRYsCv4Z8V/N/MixDu1aNT+4Z+dnieiPnh/gx8cTbd
JxVLCXa6jSUttz0iSKiUZbegwqRCtXzB2T8LarNDh9Lt29EzPsZ5DnlUY4jbjGY7
YhzRQ98ynu/l/U/2S2eAKQuwqbcFxAh81kYRAPyjuFAKN33iUo8l4D2dAnvgeCdP
QI1BdqhjL3CHAdFq/BLBDy/4zEd1TMqL3gDwnTyi0QylMU6hhHgkoT9Jf3tqXYcK
AXGO9YGH4xhXOajZmBKK/JkNmVmluHcOxHiCd1AgJaCtPd1hZ3RQURRp6HNAkcqu
veoGjPLkvxW9m3lMwNLaaAIZWtEnh1Tlakj8fEHSpRdVRMqeaDMYGBFy8lmTYyzq
Fda1zSvt21gUWTJyIVX5mFCU5RdJ7Sd0itWWOX7ctgrWarzSjEk8h5NrKEjdWRPA
8oc455hwt5vgWWINrTkDm/ximdZHIl1N1ZL3aZjuqJwU2vKvs9j7BtiHiLjtbeL8
ncrhp26gIThvroc9EwWHBxZi0v02jNisDzehZVupZUQMRHqGWL22lbuYrmfekPVz
ew5nbbMhqBjxno5bwNnp3SOaEe6DKhJVVAijTVRkYWKRVSiLOwa+vwacd+YghyAE
ISQP1dZ+RXuBlchQ9VCggNjXTU18zQHSr1BmOqz+V5jAleHWRnondAVCm5TUFNGr
gCdhO9aFTiCg595Qd5sVOnYopKrnIjBQH+ALli3SBYRGZotsCxXDXq1VilhNmEL+
TTZGyiay3c84GNpIBzSATA==
`pragma protect end_protected
