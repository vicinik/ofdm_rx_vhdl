��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�G'?��,�b�*i!��f]��
�^��መ�����W��y�?�x풟I�p���j�ؕ,;Si�o�Y?�q�"tG}H?�S,��Z�fz�Km����6��-��o�yրw�y� D����a��vs��68PqzZ�I�"�"Zq��G�("��B��G/�[v�i���PurX���q���An�4���A�POOH�����f�*S�ڞx��'�%��>����}pB������*���h}����l�"�Ǹ���3u��s�߀�ye`��Q�J����"��>i���s�T�n���7���U���(�
�ؽx��
�����i-����͙_������%em�1�@����MM�9Ԋu��HV�O�u��6��f�(� '3��#�9'g�>�7零H�e�A�8�/����� ���x0,�Bk���6<)�-�1j6އ�s6"�8VlFZX��T���x�_��`U&)͉-"m����H�baK��&���h��lP�l�`�38�e�Uo�\W������n�A��1�Rb�7Xe�۽C-�w� ���j�ۮK���]Kq@�y��LfR2�&���V��k��^����~.�JA�u���
����,1�����7֒ĸ�{�lA���7���4��E�£�w���>�g�EqCIu"�r��|-g�q�1����~��4� -V�x��3OB"x�U}�^�� �CCX*�	PFD��%W� \Z��B���n������XŐ�P�S�貨#)$g��-�ɔ���8e<Oi[c��Fk��ߔ��T����uRa�w��ÀAk,It-]���|��
��"��^t�V�����Y.���\�xI\A�W�M�+�`9��ƫ�vz��ۭ��6W����Gw"�OA�FɁv��_�a��	�3t��e�ǆ�S����`�S��c<��O��}Fܜ�M�,;��8����LQ�j0�@���]>]������=~���ߨ�?�f������/A";�=D�rn���K�>S#�h^9ɴz��#ڹC�T/�� �Wªf���e?\5P�,�
���{�PL}X$��>�o�c%��vd�
Ddy�������^�Y�8�8�k@H���ƥ pB=8�˦n� �Z�7�k�)�����4������MI=��J�Sx�ȸbY7�W!�s��877��>�ʹ�����O�����0�[7�S�<�XF��In�ޔҤjS��=[��3(�/��;Z���b�	��Yh,��{�3��
8�ׇE��'1h�`�qz��n�A-�߭��C��*ܲ�_�]�G��Yhsm��RW�x|6z���tR���siAf��Gޘ�܅Jg����5JQ������?hm<Y�(�Є1��:��
�wv��҈P�G�@b�y��>cV[]� ���*�OV�"�\���PO�u�+d�N:�ֿg��&���}�����s�)p��l{$-9^�R��b��;"�dS��X<��7mwj�L��G�dt�6�~���)-�"ɿ��Z���$��>!S>�x;��������	�&븰�;�N�/�N���9b�I�?��0��)>�(��("T*�*��Z��C+Y�s��u^����yL�"+��GSV��Ŗ�L�:z�� ��EHMT]�Г���ES�l�+��z�wk�ŖZ�c�� w+0�#	b.���	w���'>+82}����-};��/���ԲY�R�0��T4�ej�h�Y�~��Fg�{���R�c?�Ru�B5�G�~]����ć�Efh�=(����-f(H;4�+</O�K��`R��`�2�M��rW���/3�v|�P6�¶�4/f���jF8���t���&��I�ǻ�.��#x9�= A�#R	zT��'�S�i�S���͸��{F�I��Ȳ~𼑉�I�3
�8֓_S�Mpr�%�2��L-�ҍ'ǝo+�5g��7ڋ%�kcg�|L�Dz���د(t������¶<	��!}��Zb[���"̀�Ok�q_a�����l@M0�^����&S0"���E(�hZ�����D$W�<R���Q���d�ǈ�7�"h̸a�%Q�h&-Q�6#P���ND���^�׽1k������H"��WFQ�����H>����xn=�KE�X�y�����;8�I�IxO8�_$M��f�S����-�Z�?[�%Aq�.%�VP��UpdC�cu�2���X�cltk��ݶ�E#|�Bn��-�jz��ݙ�~d�&���|}Q�������R�֦j��w�ΐ�4���C�˥�m�-�3�i�������y��T�g �[��q�)U����q.�bltUl��0*|�)ѐ�L���Zy���/S��׼���g��5�W� �^������ �D1��n��;�[�1>�8_o;Y��P�0',��h�޻�Sw͆E�*���8�����{�(�Yi��H��ܛ�5G ��C<����
�����������%48�:�m���%�g�4�go<i�f�����d��@���0� m��2q"�Ǻb)��m��K���?&��X�ã=S^Lv�ʷp����h�� �b~7��Ki���e^��tR��s�w��t/;t,��t(<$#��KK��?G�=���F��]J��'j�v����V7�X��H9u���H�s%\}Oغ�t���c��~JFʇ�fp�7(�ʥ�J* ���q�a��-�~�}#cٺ�1~��Q���AM2��W$ڷ�� �c�����j������Í�<�sE��6��?�p�4�Sm���=�
׍�\𳑰��y����6d"=�VJi�I���`�s\� ��"���h���������C؛��x�f�;�o�5�io��|F,��=��>�ۇ܌�;Ⱦ���&�%h�Q�7{xar$�5�����C���8F����.��GX�I��NNR��A��
�xd9ѯ�g�wH�~D���tyFg��U7�R3τ������,�E3�;�[���K$���u@~%6m��D����
�2����}�qI��bd#������>_"�g���H��hy$v�z-D��Q��NT���'?#���{�p�薔��d%I��!�[���;\(��e�#L6��� ��m�<S�)�_Xf�N�mN���w��ֵll��@��Tn�Q捳�4u&ĖA�w�����*��0b{��cP-k��=b6O+�|T�� 0�c��d����7D+������~��>�x�9�}ouYn}��P��y�>1ӣ�$�^�A�9l�Y��l�b74�!A��8�}�X�̶YwEk�9���|q�'A�}>C�����|��HvT-܀�y�V���+�S�>n�/2e�G�k��{�?_�bip��Α�]����?Ŧ�"�JIҌVw��TdY��,C��2b�b��D���W����AQ|��Q��"���m�:6�	W�����f����D���c��5�E�wmR�Z:0�9`jiI@���"�;d/�y�fA]�ƚ�����>Z_a�>�Ju�����JU�ׂFh���=�bĉwV�yxd��w �ݭN=gI���%�	�� 5��Џ2�@y���X�h��/'y�j:;�$#];zj�Yp?�, �(��.;������݇�Dޝ8y��@'���51���
��ݎ�;,As�"�`Y����W�4��*e��Nd�zS�]	W�!�	��{�]/N�%��_�j��y�_*�Z/�
������2�C�߃�bm}�a��8�k���U��)���F�!q�_� |Ɗ&������~��q�[j}��tUNSh��s����r�һ!�5�A�$�u����(o�#6��#� a;es���q*���E,+V@�)y1Y��U��Ϻ�j
<C�ñ(�q��V������� (JR�r��~,�{�YNS��Wo8�=�z�?�՝z;�����6�
���s�7��v��,��a����Sd�9�AD�y�q��O���7�hi>�ߖ����f4�?-WŹηmZ��Z�[$�Ig��ڮ���Z
�]Ѕ$�ҟ*ڿ&��g~�%�����n�x0���=	�p���s��=��~fӅH8qJ��"�4�UW�i43-�f��s)]0v8��A���uĤ� ��b�+�����Q7PH�Mp��}�f�F�u�ڶZOG�6�L�bs�@��#��{~EAܔ}\Eф�[2mrT��s�ͻ(E&#���Q��V8c:-j�ܿqT��]*Q�<9f�l����>��!̭q���\���̡	��t�Q����G��_��&��Ǿ�y��pB�>�@͖*�!=)�7|�O�5�U_�C}Xx����`�~����R���$0��LDq���H*��g�nC�mu~����k E�_8��>�		���~s���kzAJͨAԨ�e�����"_�pX��K�j�%�%�-������|��>.�hcX�^P�_֙d�0Q2�"{�ĨNt��"A�$�
έi���$ެo+�%\3��Y,���H�z�W�k����.J�x�����L�t�/���Lji[���d8(:�X�LQ8�<2��C��a"/%^�5��X0���C/"�oP|�~p5�_�,$p���P�߷�f�̈��n$@��@Z��h���jU���uOf����)�l4p%Ɏu'��}�UVIC��Ê�Q�ԧ*_��Z%O�2�0�[^͜�Œ`���3�[��	Ս���U8�I���ői"���V�.�s=���,Zu��X�[��V@�ۃ��(�z":��J�S)]�J����w����*ڮ�
�	8^4��s-6��w�
6O:�t��y�}PcZ.�� F�<������ĵ�PU�%O[���瞕���8��
v���EU<��t�9�@a�ɭ��C|0�[*n����g^6
�T�|O������y���	Op�̉����փ��t�u�����7"@���W�&D�-g�����b#�$f9y�Ui��_��b}���x!�[�3ƈ7-�H=}���L����"�,z ,��.x��ߒ������$��_kF��P������:�={����4�/7��?��9����p�G���<k�[w#�z;`o0���4�ړ���ҭ�R0d�poc	����+U�{2觽��>m1~kf�S!�ɖ�?y�8�N���[Gw�2�M@ ��i��-ѼVX���M�UM��<��N*Iq�	Q�����[H�f��I7�����А1� ��0��c�i��0����WL�Y��\d���f��6O��Ho�`�C��,tN��h�c8ڷ��Q�\H��?��̃��,RQ
4 �E���7�y!Ri0q�рA�O�1�ԍ�~f3���3X�d2�=E7�KD�ߩ��4� �][�d�f,2R�R��HPM����T���&di_�/7c�m�Ye��R+_~>����5T<��Y}(5��G��wtgc+����B0
�ˑPO;����!��'�)�Rz�<�Rv�}��M%�l��?ӱ�� ��r��?T��i�"�$�24"I�9����9KN��h��f���d��>UQ&�K�2��A+�b�����H��$z�{o��XB�@��ݽ��v�*B��[��[e�yrsm��ۅmr�T�˘:�e[���5��Kޅ0f��쏜�K�KQ�u�g�'�D�������%�����y���EǅY�����z.�o-��`���x�Ҏ"#����:B�f-Y4n��@S��X��*�%x)[K�g*���X�[8����wHX�n"!^��5�����tѐ�3L-�ƅeZdv}vKU�c������Ӯ��l1�e�D�oII��J��f]����B���P���-�=�����y�H�CM���v�oݪ�� ���m�e�Qx1cx��b���q�Oy�t~U�:l(:%�V�{Ș��נ��)�P
:��Vlt�Y�ڏ��0���p#K%�����Dh1CM�#9P���>D`��P���a��q��|��c����XQ���N*��(n���?{(���FQP�3�`���17 �V_�̬���͝�:� �tjttk9A������R(����[��ӱ�G�B�]U�r�����pZ��v.rn&�y��_�4��k�z���\��h�\T-�U_����>�����a!H�Ux��f���Ƿl���Z���]3O�L2�^s8�N��>>M��Z:���O�t�B�:�&�K^�&B�>��d��`^h]\���Dwȇ�b���5!�Ϗ���~�G,%�Dy��M��1,��Sϧ�}��w�UU�փ������`�w�嚦B��;A1(
�:�/�f��X�>h"U�KÞ�J��r��)��V_�Y>�ew��y�
N/m��vG�.�'@$]�$����֞�u\?�Zt�p�1ޣ�;���{�͞ �*��	�6b��0��%_�A����H��f@"G���nl�*�g(8�$�p+Ut�g_��}גZ��̚wйe��y����A�
����蒾�,4�-L�"ۦ���
DY��㹫������(L�cK�Δ�|>C0K��51Ǔ1������C�C��9M��P��^��q����]����T�I��TN��Wk��|�uM�h��Jc`�y��s�}��H�ī���^h�&��pW6
�:�a�S͆�~�7!�F�o�qA�$9�С�E��y��-%��Ƶm�|ֻErn�r80]i�@����^��",���z�o(n�W �K�&V����C����bH�x3�7���pk
�s��tvB�d��l�W}r`�s���#0$q�k@�"��dC�p����d�#gW�	*X��OC���lL�-�<�E�#��-f�wl�k�v�0K�DX��fI�\:�	�� �U� �VQ�ûE��-\mD!��d����;@J������D+��\�_#��ӒO��,��Z�S����"�]�[�!�a�R%��O'�9��f��1vd3n���B��U��h����&D��Ta���C =�Iǆ�����qK�n:�f��`�~��D`�Rm�(�)��(O.���_\��:��~�[�!gO�obo�'{O�/����1�n|yH�ɬRK6��/t�l�z�
&�.0a_?��� �h�[#4+�r������A� �� ��#x��n��O��"�V����EGmv'�*����g/S�,׃?�G^�Z�V��y��{���	_{�{5���,�^��ފ=�����!:�����.��)�-9zD��)�c�)!�S��F���g<�k���(�sPޖc�5��b�^]�6�GBl�X�ȳ�o�M_ᠩ�Dk��Wi�ŨҌ����5�~��@�`�*�vҊ*����\���k*N��3��(��^�6�Q�
Q%��#D�U�<��ܓ/؉�����,��B�Kك��i���M�,�0@���� x7��dX���n�h��vvB���˲�a�(���<n���<�|� ��U5T
u�a���#ˇ�ѯn)v������ ����⯡?�Xy�������|9M���=��s����t�ص�@km�'��	NZ�N�x��gu`I�S.��T��zs��e��Hv��{�DH�������	�r�^��-���5��b�w�N�%��ņ&�yM��-�+�p�Y��+��ۚ��tS���:ੰ0���(�5�m}	!;����p7�g���E�yTs�J�o5^�X��n9v'� ��/b�;�i�W_����F��;D�q�}W��?nO"緯��YZ`'����O�0e>���u��>�s���-ǁ���0�j9\^��кb���w D���� 0��|eadW��Bu6[r0����6II�岓�Wi�o̬
���=�8�$�U��`{C���"�ծ/����e�f��w�>^FΘ�b�����xo,Bȿ^><��?��Pi��l���sw����	�+#��� ����D����Ʌ�'(�U�<�B�Y$�4<�)Wi��I.:�$���=v�+8ĴE�_�a�d��_v��#9g�ԁZ�h��U7�XL d[E�QAp�	4�wQ���K4o���nǠbj�,�~�9}�@��=�+(]�戝