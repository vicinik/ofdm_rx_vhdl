��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7�����������	$��BR/�`�f����=|o�hN�<Q��^0Fx{!o �<v��	 �[���y1�E�Tڅ7I'��7�'^#��́��y�'�a�� O�KEʇ�m����@��=P%#3��(M8���p'����U*9�����J��Zm�;�}j8X)��Ӗ]?yMm����mN.������j��p�]�H��%Xg5Ԥ*�X���9y�J���\���7{�f���]V���^+�F��6��?k	5�H��9�<���w�at��a�oA[3�r�QA���R'�`R�^�鷃07���)ص2����d�\�跮�:�˄�	
�bqMBܭ D�"V}5y5�"9�|,�K�T�҇�'�.# O�&N`�]�סO"�xN%�������(ԩ�5���5�M��ԴxR70��iG̉n�p�U��}�O����,��!S��\ ���|~�Nl�1k2���뺷@ja���7~�&���t.�,X�]μL�Fe��:A���NI��K������O_���*Y�#��N)�����R�*�vDh�#���d��\��1g����%�'�?���%���T�|�
�Ef!,k�J�	�m�-���
ue��e� Ѱ
΅�옐��+�k�W}]�eC�~��
a1߁���N´w�1�@���9��#|�>H�t�QU�bX���5>:�N4L�R�;��xH�����6 ����0�fv�qWn�|��rò9t$l�%��³8�0&��`�"PM��-[_�a�5ѷ,��[他���\>݅/�4h$��
�;�W�m�A���2��aD�q��A*&��W��)�^�T���\a�8]��F��[!�s��lFZxy8����7�6}�
��:��7��b9<�A#a3��XYu��������{+�C�~�^�Y����[�y�ޚ/W�"��_KI�#��̐f�[<��F�<d�H�q����u@�/\�ΐ?�DK:ն��펬�6ܛqf,�Wazh3�/�m���X(�������na�D��vψ	<��n�����I�����u���L�7T��!��G�K�ӽ3 �)���ބ-�*�y�9��W2�h���_ʏ�R��]1��J�*�W�����e���肉���P/�"R5oS��ި�Y�D&�,����rV�G9Cʋ	�к�8GZ��n�2��lb�P䣊լj���3���W ��=x��X�|����G�[s{ҋlv�ؗ���:�V�b�}�Ζ��U�w�O~�b
C�a��Y��f'�=��o��!�8��{����Z��\���aU����ʎ��	�+C����h�E�r$.�{G���ނW`�4 Iཨ[�Ci�P�H����oZ:�8�^)��=Pl�/���c��"�4��l|�ؑ��8R�^YW8����~��.'��;��0�S՞:
��jz�`�Dg~�˳V�{J��	�[2��9~GHk�A|`� ��	B�o�4�}L�"�����JP
`8�B�-��ڏ�2�ab�B������v�J@�OcWoJ��
�ӡ,���0�ɭm��*wzjq����6�\O�0孧�ϔ�i��Cg��ǂd����:���B��[	r�~f;��3��f���``�ҢmT�C�HT1�����	�c �@)q�l�%�(�F��˽N�[z�������7�3��B�r3�k��1/CQ�l}�� ��j��ɲSw�4sܴF�m�C��v��{� w{��1�����2mQ�ve8�
Ȝ1��N:D��K��7���'؛ ��.5�W��*�m�ᵠCᱰ��&�b�k�~�����Ҥ��Ω��<��pD��R��m�F1u����J=���1�pF�O�� |w�m�r<�`���q�)f�i�Ȯ�:�Y@�qD������G�?�SS����J&��(��� 3�K�L�{5�#U���һ
�����L�l��1��� >���'փ�W�t��)9��pj�BX�����%��Vk��y*}���ZKp}��ᖷ�M��5ģ�O�b~���i7�������WuAZ_u9-�����S�����W�&U��O�#���*��U�k�[���cYi�P�Q�7'2�ͧ�e�_�Ī%�F�Cf7��N����ִ2����I>�YK��T����b�.pc�Ax�ڧ�q-����[�ˮ%�E�t�6���� ��C���/1NȈ�(ܽ�;^��Vdh�
 �)�x�8raݦH�`��k��������N_!�!�׺��1U�0WoF;���;5Kv>�%4�?��a���ewa�:�=M�����|{���1?�D�ޒ���T���3�)���&hN!���XtY��3$5��%��)��l�62n��b���swl�V�U` ���'Q5�*��#|F��#��L��i;�d����n�y���쨠���w�R޼�$�����b���W�-*��s2�4�� a�)�k�=�U�+�~�u��JIaK���*������lT���$W)�|&G5�R��m%@�r�^��2,&5�ۺ�H	���{�2��;L���6��>����\�[��:���ԑXn��������xɓ�������r�Z&"�L�1�5MK����
.���>�-{�hd��)���=�T���"�\�)(�ɣ�I��$`��܅a����؀mA����|3W��l\�ԏo����]��f3gn`/�J�L�@��	�:���%.�nH��X���Ǆ�켑�[���}������{��4����	v�Jm��]��͈!�F�/��i����k2T�f(b�뚵½�4rA�_��N��^ʰ�[DȢ�S�b���:N�� ��B���U?z�E�=��Sx��f��˾#
j�c*=�2T�ݝ=�1�K�\*aK���-�G��\;��z���&�&{_	�%�.p.]�)��4���2_�t���c׫�����s��RB�����骈�$"b�Q�X�t���Q���cӻ�&�Wl��׽��p�;`˾��X�k,���l�M�`�@/��h��ٛ�gٸ���Z��u�����a��s|��\�j�9���`�a�K�e�@H�l�A�KTݠ���k�̅�'�����(���L �k<A?<(�җxs���o��DGkJi��J�|C��G9:���/7�6}����������cW6����/f�����*����y����?`X�]B5=j���ko�}�?˂���/޳pG���X�[�8i��o�H������@er>
{����E��u������� %��?�o%��3d��;(:E��ߪ\Nv�k$Y1�hẖ�������E.��:{R�������tV�fଢ�^+�o)�ͣ���O�Ղn�IL �^pc��cj�U�ɶŨD�q�b\nU��N�D�m�٠���pʢUF��v`dpk�B=jV^q���y	��U�.2��!��$y�>��@����:%_*��G�X3�d֔���g�u(�U���)���~η�����ᚙ2��Y氬���[�JW��B�U�.X�x��V*Pm��6ō1�fy��q���e��!vTJ�za�d[= ��y��7�5� ��k��O�7�x�F���yގgr���� v)�ܟΖ�B�נ�'w<c�D6	�j�M�p���0}�\�*�dֳ᰹z�_#`�ܮ�vT��20h��b$F�<R��
�����#�%�(��Cm@1RRHUMW�a[����
~�~�SN�~����N�t�`�1���%+!��,J�_�,�@�lHa�mt�Ɯ"���)B��kY���⚐��v��(�o9J��Y��b�t�pe�$o��M�̫�@F�i=��ʒ�!r2ㆣ �I�KH[ct��DI,��ս�g�C��x����a��Ǯj��3WQ�IcK��1Yܿ���<�6�����"dG���_�q٭��akHm:0��g3���>1���4-��%��]S��HRo%X�En�_ba	m�*ׯ��jR�s��ڧ���W4�N�U��$7�q�R+P����>S�5�z&h�Y��B��<qvS��L�v�B}>����a��rW&)�w�&��e���:���&�K�/FF�6�z����O�c]�׌Ćg�T6��㘔|"v�p�M�h�TysR*�hg�6ͽ݉�?/�M��1�#d�ˁ&���>'JNZ؃�����3����Wˏ��Q{�b�MΧ�,5�P��!��Vs�j��ڳ*�l�����5�5-�x�2���0�I�+њt6ί�C�����r�ͷ=zZy$�������V#?n�ĉ��o��")��jB�]�O#�G똌�}F��_�y��yr��g9s�;�U(�N'N��򼥿`�&�R>$*EQ4_6.H1��ġ3����1_7�%�>0�� �+z$���`���b7)Q�1ұ0Q�kP��)�T���+?��� O�Iք�V����^��wK'�e>PH����q�S��x��f-�h����O�sٸ�R�eL%r܌Z�
[d�|�B�e�׷΂t�3�rvsXg��ӈoO�x�uq!�����M���1��y��H�F�c��������ՔT�oBA�AZa{Sa/�T)�J�l[�j�&�0g�7��!Ϻ`��T���� ��cY)<�_�&vȵf�qD�naH�g�K�|�$NP>Q�)�5�g��Rt�%�|�5*_�x����wD!��h��T~I$�Ή�d�#�٦����?�Ӆ�s�c�,k�����ɳ�0q�\���
n 6�-4=G��O�t8���.'��-��$Ǔ�FG��:߃�$:`��y�|��@��<�jR��?Q��Η�ѻM�VlW�>�?͡q��Պ��t6v?��<�{lcf$;�M��?�9x��o{�R=>q[~Ѭ.���Helj�?�O8�$��)�/�Z�Σ��s�8��M�:�?� c��b"<��2/9�l `7�(� 9�����B�@h����V�{j�$�i�Xf�X�Ρ9�N 4�9=��p���	��D�S����BlQ#��������ײ���~o�!TݲF|T��{�`�PT���B1S����ښEt9~�����8b&y�^(T��ɺXv+�N�)�v��Dp"�sp2 &ި�f(����싪�V�E�'(ƿT
�C��v�\ф1ℜ��44KFnQY^X���f'`����ٝ�+�xG�Q`�Ѵ�vUC8ǲ��F�m����D;v����ȑ=ot]mw`�4�Q{^S)�u����7Tr�ΰT�����M5�c-�xc]O��{���c�Dbd�"���\S^��A�gR����B�)9si�b�{�ZZ�1lFyj��1L�KIB�q)U��Q=�{AY���&�W���ow��j�2(���Q�V��E�XӾ1�u�Bk�z�мp<RYx�h�pHMEDM���D�.G� �j���:��D���_�;��=�/�1��=��f��L-�&��#��a�_�ok	��OV;��U��4A!W��^g�'?i�.A�OD�A&=��+c�.:ҳk�צ5q2^eC)�RD>͋�NHx��h�6��j�JG��,�&��6�dٷ��"�R!�FB[~ى�J+L;z,iq7��i+�\f��Fe%���%���Eب,�jO,$`M����'}}��oGw���2�Cͨ}���w����6�א�����b�y�y��K�j<�)�>�U�*vS km���z�����O��y��&�<����R(�PF�8�R��R�$��u�s�C��/�Q'�%v|��`�| �����L�������Hh����:��|�[�_�z~�����9���O�:�j"BqK�z=�ͿO���h$%8E���j�Y�z�__��J�bIƷ3�m�"إ-���ݖb��sZS/y/_�L�.`�]�ᝀ�c�چ�t�J��Q�\���:�W7:m��*=��e��BN���3G�nSD(���?�"�8q��=��&�qJ�tk�Hx[�>��a����DG�d�-I��z͏5�+/xw&��ᙖ/���|�Q^�4�|9����'/�譱OHP�KK�Db!X�XF�!&~v��Q�M�99�{l�68C����rC&�8&��3���g�pB����)Uv�l��B�O���u�-�ո��)����[�Ǹ�:����悪��B<<崪�ь�N�Lㄚ�H�>Ж���y��Ѕ�J/B�(����g��D�Vd#�����=��N��� t+�4�[� \�2��(�7�&E��|5�N����vF�?YD�|�9U��@%��ڐ�Mp��ň��\�� �$���W���d���5G=c����T:.��즴���6��+h~L��hw�5�+���aV�iό�m�=n�H�~w���ߘB���?x?�U���d]b@�����:��\I�<�����.>H޷��)�aP��Lm��*�u(�y�4f����(���lx�z��_�$�	�"�CY���p2�]d�+	\�_n��$'�H�#�������}��q]��"��o�#��V	��v���!8:\.O/��]cdzM�����{?��W�L}����v� �f��1�~�����������-PO�^����l̻Nz�k/Nw��h�V�rq������`s�Z&e�µK:�F����$���:z��~���C��i����O%V�hR��/K�K,�U�=��%��U�*8� ���0
��@��+�^�B�!z^���q�x�hP90��M|<j�����KR�Q9Cf݆ڙ\�k��w�(!�U4;`��%���L�˺QGC�����0ew�$��>��lO���e[Ez��J�y�`>[9)c(�H!��h�<\J��C(�t�����M��טQ��#Gc��T(n�����)GlQ�J��x�����*�jR�E�0�؀,·�_)!kx�7UN��)Ɏ������u,�/���@�A�9��'��|"�0s��q%�X��7�75�����N |y�;�x��6���h��[�w�m���D�RH��נR;� �)��O�t�����������_?G�a��O���-"��
ב"u�C�_��)F5̵y?+Wv��Te�d̓���,��$��:�%�|��b'�69���́�V������X!|~�D�"Jv˧q��΍|�Y�0ВB;kU��n��{��xHY��)@��v��S1�H��F�b�����J���%0�y�u�pU��I	�{��rU��
x��p�[~�H�jrb��}ʹ���'.g��/0��7q���d�g�4h�! T��0vj@9�h�g�y3��:bȨ�83��@x.���:k�gi�M�� ��I���`��+��ֳ�Z��TAm�7�9e:�WM=U�?=��HM�1v$�-P�br`�/�_�'��滸��֗Ϥ��4LI|�x|p�8D�����N֡��,��X�!%� W|��p��4
e4��Ԇ��s7�!{4Jﺌ�t�i� ���h7u�[�y��j����Pq(:Q�A�mN5��5���1�d?�1���5���-^���/���%;�0;Q�[:�e�Q��/y�O.ȒF�N\���'J#_S�Cz�`�Κ�V�Y.~-�m�*Aw�w}<U^)��9|*(�
j+��2
wܤ�|����I%qt����R�ç�H�˛ l|V�Y�.oW��ѳA}�7
����< ,��V]��j�B��|�
L\Z�%�(��l9���V���ǠvJ�<E�ߋ[�s�����6R�V�r��1;i^2����_�\�4����U>mSB��,��ق�gl�t"��f�yr�?�uʍ�6$60�����k#hW"s���X?]�f�X<r��Rb#�R���^�:i	&^�P���?4��`��!��h��Y�ʾ����������>´�2p z��_-ij%@:������yC�:,@ ��_�%rS%I}r��ފ�=��f�?Y�|�Hy7fL�-4�f"sv�%�[P	���}h�Î����!"�FJ����DV�E�*�-{_㖄�7�Z�8r����u�������7�?~)A0wM/mk��輅�8W�1�j��9"l32s�C�n���
:���+��4��,�#� ���'z��۔�fö����������{�& +y�	ۂ�]>��nEѻ�ќ���EF��	��v�N� �G�]{+Y�z��Y�!����kSt
�i�����7�#�@}�LE�g�IxB�������rpb�p�#��#,����5�[~z��̭CrR�k��i�.i�9u�t���e�x�98a3� �E�.���`�=���-L���p#ʺ�A�A��Q��Ԫ���ҏG_}��W���fN�,D!uniM$)?ؚ���Eԫ��i���}��X�W��3�v��n��dC���򃢓3�e�{>J�R`o�lsT�'��~�.�?���8�p��68�3�,��~���q�%�����.�3�<� ��h�����2-�8"%�EF��Њ��L�Z���u��J�cse��f�u���/q*�2�cS}��F�.#ѹ��Kƞ�9搚Ж@HZZN�]xrau�7�9J1�뿰�����f��߀�X��ϖwIi!5�Mb���կE;������?��6<&�