��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��1^+�{K�Pӏjx��eRn�����Q��#j0�2�"B�(�lt�3�����	�z
^aű��hᣜ��	ӈ�\i��9w�IU�h��V�0zV���@"߬�TF�a2����_␸�1r�p��վ�|+u�5��	����|�=C��t�G{tծ%�uT�J�8��z�>���vJ�c��}4|������G���٘����iz����h�܆x*�QߙG����V�S�'�)B�e�]=ϰZ?�wi��S�ㆿ-�RP��/��i��Zr��x?��i�`D�z�%�~ؑ�L/g�s�\>�os{hٗ&��5L��VSk�}�#'`�k`,�G�iy�..�VV;7�0�󨝊�\_ �"]x��%�-�CL?�k/�~	R�R��K.�f�A�tB]��6Sݣ��]��G5�'��,��ƼFeg�>j'�4�k�Y��?��g��O7Y+
"�?��8b�C���B�A�><mf~�t B+�.�8��N�i�S�'� ���[����*����0y�d\�;10��F��ח�22o�����Z�,^	�eh����i���_��!B	���]��7e�2Ƌ�z&П�b���$��0ot���q6wEW��[�@me�&0�Wi�<�� �WV�jW�Z���e��w:�)4EjNpd�f���u:��A�f�72:�}�ރsJ>hKmOK�RK�1� f�c,���LO��'H��>��S����L��]�8N}
kYZ��]�ۦ�`�n5v��\�<��m��(W�v�A6=8N+z�A�25��c:l��f�͸��{����\R:#(����I�kcV��3gf�����-=L���o�'�`���v٢���7��4<�|�E-�^�/��|Ԣo�KB�f��;�.	_k�p֓�6u[�ڢ�3�U**�-� )� J��!,�U����q�n�ϙ4/�O=}�L_6 � ���Y�e��?�o����@�N��#f��n�� ��'8�_�3��cU���Ч)�fdIP�f(�9�i�gĠlAh��ypk����g��8�l$��ו��4y2�	�k���*E4K���%�IB�Cr�
x�K�3���(���5�+�^;5Ji�2̹B���.n���|Jo�IS����D�C	A��OT&!k[��s��0�=]�Saa�:-]�,��~�F!���f@J�3�Y�#u��+F&.b�ڲ�}��>kŲX��
E�$��@���$~�[q���1��tAMW��L��7����_�;z0�ϳ!Ч���i2<��J�{�9��nWy�:(j?�+�)�re����u2j �u�z��9L��F��~i�zQ}!!�P�ė��|S�B�MZ�_�l b�~��Hn/� �G���� �O �o��|�&��c��<	'��OKs�c(�ڐ��y,��s�hPCF�Ղ���z�{��dt��� 5�ƢX��<�^�yV�U�vn�w_j/�,d��B����ܙ]<�WD�^�kOJ��^�C�g�:TH��������B��^����\��V�ROf�7{�0�A��$���vl|'Aű��̞�"����8++��#_Ӷ�T|
'[>��1�z�k����D�"kR��X8_I�K���WvTB��ա�1q��>�,,_l��k
��C��c����;ζ#���,�fs��\�/�Y���WIK��C�
nn�Q���Y�GZ����� Q2��q�^}�`�;Q/��"���7���[X8Iqk�٣���{�	@���RՏj�Iy ��D�)�s2�0Y����'ꯦ�A1��_s��k��b�x��%�4����g�o��#�1 �y8.��>��b�S��Z~��|W�+�}��=$���XIaȼtgs����8�R�{}�� ����k܂o��Ԍ��ݽ���q�c�T��AQ��϶�� ,��>�\Y�;����!�yml���Vc9"�Vu�����x���Ǌ�8q���8UV�|��m
Ix�4�0/� ��a0yK���_ب;:��f�ax$?�ʓS��n৭kpL茢��6�_$�)����)P/d��vo���a���L ��۰�N�4�N�ikȥ]��(�}֓���Z�0&�i�Q/?�5�J�<Wn�ZէP麼C~&��gI�ʴ���>ߏfr��%�$³��0ѽۑZ��O���t^���F���T��-�,�	�L���$�L|�ҹ�����([����@��U�$����B@ߩ��@�`��JvE5;[8��6X�[t�Kg�赥��>m��B2�]V�[��9��%*�B8eEe?��ë�U�6�#���MAQhL���.��\w�j6<7��X���z�H�Qv.��xyM����Vi������W͸qL�$�4b�����Ԡǘ�m ,�wR�%���6�	�mظ)\�y�Oi�\�+V�Z�p[ӿ���>M/R�q����l��Wu���;5ˉ9�h�����_���*�V�
� �O\ƾ��΋6���6�}���ƹ�"��6m!fx�h��j��!+8�e��XV�Jد�~�$�]�FܓKW�~N�V����c��z����3���"�H�K��@�`
�p!�tfN��.wo;J��N�h^M ��U�E!��]GM����H�m�6�Ҭ�|�\�P=ڥ��ϯ$�>Ŋ�)�7\eŋ8m<B��QI��W�=o������]4e�t=��������'�7��C�$�r�|�4�o�J�Pw�5t��8��(�_#�r`�Wq��%�@R@�Lt��v��@>��.n�	x?�����e�1��9�pN�N����*��5MׅӶ�ֆr��:VZ�_ͧ|�F��Kr:u0��]`vr�S��tt��<0����,{v��H~��]��K�<;U���c�{kx�]�z���q�q�aP��G� ntz�(�7Q��9V��a�1{}���tqN���D
/���o���ܹ�9*�>䡌W]��t�e�}=2oD�pL��[�@2�N�j��2мp�m���gCZ������I�eR�Q�M� �����m��CV"U��a=�h��Ϩ�|�W��F2��m+������