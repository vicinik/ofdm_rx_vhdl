library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tbCoarseAlignment is


end tbCoarseAlignment;


architecture Bhv of tbCoarseAlignment is

begin

	TestSequencer: process is
	
	begin
	
		wait;
	end process;

end architecture;