-- FftWrapper-a.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
library work;
library fft_ii_0;

use work.LogDualisPack.all; 
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.LogDualisPack.all;

architecture rtl of FftWrapper is
	
		constant cBufferLength : natural := raw_symbol_length_g*3;
		constant FFTLength : natural := raw_symbol_length_g*2;
		constant cNumberSymbols : natural := LogDualis(raw_symbol_length_g*2);

		-- Components FFT
		component fft_fft_ii_0 is
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			reset_n      : in  std_logic                     := 'X';             -- reset_n
			sink_valid   : in  std_logic                     := 'X';             -- valid
			sink_ready   : out std_logic;                                        -- ready
			sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			sink_sop     : in  std_logic                     := 'X';             -- startofpacket
			sink_eop     : in  std_logic                     := 'X';             -- endofpacket
			inverse      : in  std_logic :=  'X'; --       .inverse
			sink_imag    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			sink_real    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			source_valid : out std_logic;                                        -- valid
			source_ready : in  std_logic                     := 'X';             -- ready
			source_error : out std_logic_vector(1 downto 0);                     -- error
			source_sop   : out std_logic;                                        -- startofpacket
			source_eop   : out std_logic;                                        -- endofpacket
			source_exp   : out std_logic_vector(5 downto 0);                     -- data
			source_imag  : out std_logic_vector(11 downto 0);                    -- data
			source_real  : out std_logic_vector(11 downto 0)                     -- data
		);
		end component fft_fft_ii_0;

		
		-- type definitions	
		type aState is (WaitOnFFTReady, LastValid, Transfer);
	
		type aComplexSample is record
		I : signed(sample_bit_width_g - 1 downto 0);
		Q : signed(sample_bit_width_g - 1 downto 0);
		end record;

		type aSampleMemory is array (0 to cBufferLength - 1) of aComplexSample;



		type aRegister is record
			State : aState;
			SampleCounter : unsigned(LogDualis(raw_symbol_length_g*2) - 1 downto 0);
			TransferCounter : unsigned(LogDualis(raw_symbol_length_g*2) - 1 downto 0);
			ResultCounter : unsigned(LogDualis(raw_symbol_length_g*2) - 1 downto 0);
			Result : aComplexSample;
			WriteIdx : unsigned(LogDualis(cBufferLength) - 1 downto 0);
			ReadIdx : unsigned(LogDualis(cBufferLength) - 1 downto 0);
			Start : std_ulogic; 
			resultValid : std_ulogic;
			resultStart : std_ulogic;
			eop : std_ulogic; 
			valid : std_ulogic; 
			buff : aSampleMemory;
		end record;

		-- constants
		
		
		constant cInitReg : aRegister := (
			State => WaitOnFFTReady,
			SampleCounter => (others => '0'),
			ResultCounter => (others => '0'),
			Result => (others => (others => '0')),
			resultValid => '0',
			resultStart => '0',
			TransferCounter => (others => '0'),
			WriteIdx => (others => '0'),
			ReadIdx => (others => '0'),
			Start => '0',
			eop => '0',
			valid => '0',
			buff => (others => (others => (others =>'0')))
		);	



		
		--SIGNALS
		signal sink_ready : std_logic;
		signal sink_valid : std_logic;
		signal sink_error : std_logic_vector(1 downto 0);
		signal sink_sop : std_logic;
		signal sink_eop  : std_logic;                          -- endofpacket
		
		signal inverse      : std_logic ; --       .inverse                         -- data
		signal sink_imag   :  std_logic_vector(11 downto 0);  -- data
		signal sink_real    : std_logic_vector(11 downto 0);  -- data
		signal source_valid : std_logic;                                        -- valid
		signal source_ready : std_logic;                     -- ready
		signal source_error : std_logic_vector(1 downto 0);                     -- error
		signal source_sop   : std_logic;                                        -- startofpacket
		signal source_eop   : std_logic;                                        -- endofpacket
		signal source_exp   : std_logic_vector(5 downto 0);                     -- data
		signal source_imag  : std_logic_vector(11 downto 0);                    -- data
		signal source_real  : std_logic_vector(11 downto 0);                     -- data

		signal Reg, NxrReg : aRegister;


begin


		FFTInstance : component fft_fft_ii_0
		port map (
			clk          => sys_clk_i,
			reset_n      => sys_rstn_i,
			sink_valid   => sink_valid,
			sink_ready   => sink_ready,
			sink_error   => sink_error,
			sink_sop     => sink_sop,
			sink_eop     =>sink_eop,
			inverse      => inverse,
			sink_imag    =>sink_imag,
			sink_real    =>sink_real,
			source_valid =>source_valid,
			source_ready => source_ready,
			source_error =>source_error,
			source_sop   =>source_sop,
			source_eop   =>source_eop,
			source_exp   =>source_exp,
			source_imag  =>source_imag,
			source_real  =>source_real
		);


	--bufferProcess: process(Reg.ReadIdx, Reg.WriteIdx) is
	--begin
		--if (Reg.WriteIdx = (cBufferLength - 1)) then
			--NxrReg.WriteIdx <= (others => '0');
		--end if;
				
		--if (Reg.ReadIdx = (cBufferLength - 1)) then
			--NxrReg.ReadIdx <= (others => '0');
		--end if;
	--end process;

	

		--rx_symbols_i_lengtho         : out signed((sample_bit_width_g - 1) downto 0);
       -- rx_symbols_q_fft_o         : out signed((sample_bit_width_g - 1) downto 0);
		


		--todo subcarrier entfernen

	


		-- register process to store all needed states and values
	RegisterProcess: process (sys_clk_i, sys_rstn_i) is
	begin
		if (sys_rstn_i = '0') then
			Reg <= cInitReg;
		elsif (rising_edge(sys_clk_i)) then
			if (sys_init_i = '1') then
				Reg <= CInitReg;
			else
				Reg <= NxrReg;
			end if;
		end if;	
	end process;
	

	FSM: process(Reg,rx_data_fft_valid_i, rx_data_i_fft_i,rx_data_q_fft_i,sink_ready, source_imag, source_real,source_valid,source_sop, source_exp) is
		variable exp : natural := 0;
	begin

		NxrReg <= Reg;
		NxrReg.Start <= '0';
		NxrReg.Valid <= '0';
		NxrReg.EOP <= '0';

		NxrReg.Result.I <= (others => '0');
		NXrReg.Result.Q <= (others => '0');
		NxrReg.resultvalid     <= '0';
		NxrReg.resultstart    <= '0';

		if rx_data_fft_valid_i = '1' then
			NxrReg.buff(to_integer(Reg.WriteIdx)).I <= rx_data_i_fft_i;
			NxrReg.buff(to_integer(Reg.WriteIdx)).Q <= rx_data_q_fft_i;
			NxrReg.WriteIdx <= Reg.WriteIdx + 1;
			NxrReg.SampleCounter <= Reg.SampleCounter + 1;
		end if;

	
		case Reg.State is

			when WaitOnFFTReady => --Fill Buffer

				--if ((Reg.SampleCounter = FFTLength-1) or (sink_ready = '1')) then
				if (Reg.ReadIdx /= Reg.WriteIdx) and (sink_ready = '1') then
						NxrReg.SampleCounter <= (others => '0');
						NxrReg.State <= Transfer;
						NxrReg.Start <= '1';
						NxrReg.Valid <= '1';
				end if;

			when Transfer => --no buffering necessary

				if (sink_ready = '1') and (Reg.ReadIdx /= Reg.WriteIdx) then
					NxrReg.TransferCounter <= Reg.TransferCounter + 1;

					NxrReg.Valid <= '1';
					NxrReg.ReadIdx <= Reg.ReadIdx + 1;


						
					if Reg.TransferCounter = (FFTLength - 2) then
						NxrReg.eop <= '1';
						NxrReg.State <= WaitOnFFTReady;
						NXrReg.TransferCounter <= (others => '0');
					end if;
					
					--if Reg.TransferCounter = FFTLength then
					--end if;

				end if;


			when others => NULL;

		end case;

		if (Reg.WriteIdx = (cBufferLength - 1)) then
			NxrReg.WriteIdx <= (others => '0');
		end if;
				
		if (Reg.ReadIdx = (cBufferLength - 1)) then
			NxrReg.ReadIdx <= (others => '0');
		end if;


		if source_valid = '1' then
			NxrReg.REsultCounter <= Reg.ResultCounter + 1;

			if Reg.ResultCounter < 64 or Reg.ResultCounter >= 192 then

				exp := fft_exp_g - to_integer(signed(source_exp)) - cNumberSymbols ;
				NXrReg.Result.Q <= shift_left(signed(source_imag),exp);
				NXrReg.Result.I <= shift_left(signed(source_real),exp);
				NxrReg.resultvalid     <= source_valid;
				NxrReg.resultstart     <= source_sop;
			end if;

			if Reg.ResultCounter = 0 then
				NxrReg.resultstart     <= '1';
			end if;

			if Reg.ResultCounter = 255 then
				NxrReg.ResultCounter <= (others => '0');
			end if;

		end if;


		end process;



sink_imag   <= std_logic_vector(Reg.buff(to_integer(Reg.Readidx)).Q) when REg.State = Transfer else (others => '0');
sink_real   <= std_logic_vector(Reg.buff(to_integer(Reg.Readidx)).I) when REg.State = Transfer else (others => '0');

rx_symbols_i_fft_o  <= Reg.Result.I;
rx_symbols_q_fft_o  <= Reg.Result.Q;
rx_symbols_fft_valid_o     <= Reg.resultValid;
rx_symbols_fft_start_o     <= Reg.Resultstart;

sink_valid <= Reg.Valid;
sink_sop <= Reg.start;
sink_eop <= Reg.eop;
source_ready <= '1';

sink_error <= (others => '0');
inverse <= '0';


end architecture rtl; -- of FftWrapper
