-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
n52xnOzJ9PN2JU3+mLv3ZTl/vmhoqahcNVn88Ethz3iyubiLCq72tC8kl0EaJp/glhX1ih16BtDL
XEx3hbB3z+WeV/LtLpGo0y9j+nYerxlKzlvnWfAAoa5dfLzNSV0y6LI5cfhjv6JrDUp+zhKPAc30
tHo+MpLbJAsU4j5xowxIKsVpKzpIiSEkQYycQk1H7LBenhwyGgeyIHdT3/fBibmcetOaFvYvQhQv
dNHQ8KDGEa9Rnnca+hie33BL4FpEOzCljwQGEBSvGFE5koks8Ns/CEfyZgtdUd+4ccDAOzOcDgAd
WFq1bGwDvoZVo2T+eJlnFpb6VnSo1rTMZQG4Gg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
TtY6KPazvQdw6IHyrhzRfG+tY6K7VuVoChY+OfuFLVvrKbw3/Dq59GIuZ7o05TutBFkpwK68hWjB
UhJszLLAbWiyipu6stLB7eD6Q0XJy714zbr9lqdQNk7voGA3IBUDeivuE2eAXqvu5rUWFmTIaaew
xXXnRvr9CcH/gYINPGnmf2yAfUOLralLIo0YNtUVgK2fSGBcofRZhY89DiTR/GbZgilAGzNXoacw
7J0eM5DnoTwHNsH5uWyAfHOHWR1NcMrX/BvmBnVR/RfWusLjPlKp0Q2kpslOmH3uzgFy1ic55Vp9
65Gg+BKDIYsSH1oSMPu5lE+CYYx61K7jRmV378y/NogORp2P0rm5ftvBAA9SMmWA1quYHTouUSnn
1/k2sStky2UjVaHmc10J8mQmMKN5gU/Do0AGxZyw7A1MzOCu/y86cfmAEf6+CtFVCREI3lSPw8+v
wEjLpjQtpeZ0V5R9rACp4loEPGQ9Rh7VZ28mTfAK8wfti6qgSR1PVZqOapKGLYQQpdZOgBPh4P+m
hWZ5y+29YJLlEgsjoX/vBuCsTFpnEfEXw5syRdnsBIOATmNLfVPsdNOMJ1Dqae7LW1hWkE+kldpm
cxSeyAAFimG7Y6KAFbjRWVON1Lv35Tdkku/128CzCvo0AjwXg+lsjaWRwEjlmXSGzQZ8pBfpgHSb
ABUqR+38rLz32tyejbfM5hJOYVkDG52CyUgYxzbXsx1qsrR5YgWbRaITt0dNVegWWI0shSukp1Qb
DBhZZJupptmPhRmcKA0KfWPvAdtc/juDQqh2xjpqcvYTv+WEvBOZu42FQLqbbSaVs3foykvphVjk
13YmHYo5zwo53/qRKkax+ksTPmaJR6inuFoGeSofv/ZSwmOzTJcokx7DG17T3A5+EDS1omr7UUDa
xLKI57jjFmOWsxTTnneIma2sWnhjbnBZKVgzzX4MCUPAP2zUpYFLgG+G4PaC02rn5sUiH2+SDVa+
K/ocPayWeOfbTvcGTQCrAGCkb4PTAq8MY1rvnF9XNIyzT5j7SIyABpv682ceMUtr+VRVbblMY10X
EnmkWWQCYubWP6ul53KxuyOw7tGmLaMHWeL6Hz/Xbvn7iOz/t3gQ4tOv1M1QKiWdH1gjMzd02PhK
pHbAdCoH9wOPLdUlfdyxLWYf9Ptlz8qwdurUz/qWVh9ClrtVsCIomRISOM6BU04d/c7XMgJ0TCHG
hBS70J9G3LVmV+0PR1WgPD7nRrrIgS/p/c8QSplIWf0/cthXj6RsEkH/ZgKOO/a4Il7aSYAWISgL
2WRJdS8iJ0x/isxvB8WXSz7VkHgpOMsOm4YJQh4lU9xPEuybUhCxOEcqaa9MIH5QVpVwa9dcTqZo
ZMTn+fFJpYOf6XsuBZQlTHiXUFML/lEIZRaf4I6hAoxvToQjTEKHesPcR7q8wkB/h97fpTWRPXLk
aWCaMXZypIXyNidXFXE7izWIU4Dm6q/1S7ixhqvBsBu63UWlZVpxxChDHlf6lWZj9A2vLlbZiN3Q
aaK3d3p/qSVpwATMToFsl1GfFI86TJSmjRFMvFxLHucuSDgT3vn1P/IaYs3q07bK2tvPUnfFYVFU
mESdEAvcgMVFfsOup92Pl90091kbDG4u8nbcik5fPrfdPvrob24RrfuqHOpZ1avoVX+QHbywrHbd
aqS0hn4tQP12huX+E/kHgAdYlDRC1XVnHicQEm41oV6WRhPajlTxApiEFv790Fc8B3QGSeFwD0Xq
eTmi/IkcZGJpjyYSmJ5bLAoHlhWlHgJI2Zgp/cPZE37NOfWnp0Jmk4LoBGhYAZayh57Ea0+136Mt
O0xKX0dlK5jPFBAxbvaOauW2SKtX7OfiW0SBjCbIILAwboIZYhADtao7naeNw5dyTlX7WA/BnZOf
1BGKLTqaY78rvQ5mkTJTZb7rXCl9B8OLw42A3V2qP4S54lhTreJ09pdXnTe6ShR9JelX6V3ZpOYp
niZQt1IJQVf5Cp2WH/ivS96FXhMrNWqaVUjJS9ClMRJT8Iwi4BmR4d0slLJX8Ne97qXm+zF3DSI/
NwkLGgh2yMntvNpjT08iqel4D4qYtD/lvOJRh2+H/CN1vWoPIDIONXTaNI1rgHuLQ1sQquJo+4Z1
Wk+8Zy3xF/LwyU0lk5EvuS8igoHoFFZglrciXBKybQmFArNkK1ZmwL3jehuL63pa20554JKEPq/y
vpDV84R+ndSCdlUtDp7cimyGy/cXOEqW3e6Cg5MqfdxqVo3AeDbPmuH/gQ8UoCyQ2Jp26QHVj3kj
puXOmr9Qm2kZa67/AZQvfLWVj/nmIMWx44GEQ4nkC61wPIEVQtEUtGk/ecBMJOxUQ2DSZKCSnjrP
GPefWSDWsobHZKkTbthXPlLDk2C1L9Lh4cmyfIdDS6oTV/HhKru/Z7yeUS9TXYSE+QqmuiAr++Pf
XLyD1kVquHYzyAT2hiFzeV/ws5Q+2/U9LlAatqafH4CRN/EZrNbj4B1lAI0nZe6B/tCRmjZsS0VI
5cTidL6LsW/ph0oiQanCxm8e7vXBNYRcr/LFVyybe4XfY+sWBRF56BjONzpoZ1stppAc+N42jlwI
bZXCdeJfgOKkmQXRABiymMk7LuZee0l7aQQj6KzdydCeRQL0qLDPm22w2zkS7xtM2fWtCbN4VSzk
N4xHtCnZEyQpqmMpbjRIbAAD5e7Hx9SG1FIDHMa4T0mYC37ldLeImab5e7fjtUO6+i0XwcGaKYHM
O46FXYIpBj9Zv+xvvcrO8uw4bH6o+4+Eruhurf1iFhObPl9So4u3FrBftr0inwSNKvNhWNHdYdfG
5MXL3kqM3mJjbuobLEP8rLtAzhgfrlqj1xa3W9WHM3sUV1bDTNJf0hXQ61mPIbD3ln+VyKU2pBXO
py3NYyZEX5PTaXRiP+YEXKfLPY3YS7TxK29MfqtTxQjawpy3iQexIABjUFWFAMF5krFOomTz/ZKL
z0zONzA/iePb+pQkNnol0BuGO4P7RqJ+Z/FnTF/0JuouC1J3QavCmWfz9nZqsRd+QCTUqI1tQ7AS
x2xBtINpaPlacZXgvgnV0p91VdgKUJGw/P8GCgmgclH5Tr9Vb0HLCHTe65I1DQOQa8nzcbg276kA
28VjnT3I4cq2oJB8HLDKg1H/V2s8gGEsaNwXWIgUgIJg3pp2WhKJp38FmFrofE9J2dMnxS7mmVuE
99n14ITjdM8E3HcLNLeTq1yX7Z2SkQMkwdLAxffVblUjp5ec0fDNBtBCrCWpCI63ReUBkq7ftF2d
o5lTFZO5YuAz+Q2f7dWfCMOHiFALA4B+A5sX8Ty/h5B18g+D9KZfkSTKKEQR9Q4aeXZfqYBeXQLH
EddjoXAk2HiEgo2M8AxmR/ATzbCuPdR8IjPNwJODweb9C1aX0obk583uxotwUOG/g+rLJ+7owuuk
edD9y0rxrxXTixjv5/4Seyhv4/mUI1DN6fYPCAr9SS+W2AeLw2SnfCGSYHdnWCN471D2DesNXfZ9
i7RyoTmMDf142AzCAVceKBGwR5PjJVI8BhrMcrDz1xdWp3j5K+hHwlgLUPWEkOba4a/HD7lMlKjm
lxYiqaIyjXMSH+7v+JUBXPRYQqBAWGtR01hx3g7pIBbneF7Bp9QtqZV4skLNhxznQbefbzwW7c9w
HZ4Z41QVjPc1lxRqp0Pt5G92A3LjYL2CFnajwX9dLWct0EVsBB1SC//ZvkopzoL+NXuEstkEaRQ+
/yMI+Nwt/WoGDM1B9OqhikePH5qAiGFrf8coizQmBNOX9zHSJ872rPji9SMorYXGp/ei7/wDTTGy
uGM+y78RuzYrLYpxVRPR7N6SiXQzCQky8RRzKLONteC9JvJTcJa3w/hdQ+3RMyOyXFwhj6LcXEGl
vNu+iTDCKuNsDnnPHU8IIblUrY3zx4Fb/EeWpSWQvppz7pOI0oAR+56G6+x9oHZ4FdslCAzJ9B/c
BeUlyEWDz2PD/478DKNicwlHbMIHSG231cYL/WMwxZx6hPY5Muej+TIsGnVBrD5rrfU+19NaTLTJ
xTm248mbTnFe9MUjbznV/5NMGeVqoqjp4tkwtjgwglNeAKD7C0T1qMuliNMMI0AenG/QVZOoIx5t
kONYsLvE7vDbvdahgroOlMzobYlKiuWdi/vVw97yGL440nAtldzn2AV5Qt4dbuLjsyF3XhWMSafz
QeRxn4IsBI3MIq/oic4rXTOO+lUtregkYbj4X4LX64MJ4fN6xkZMlxXZjT8ILP3JwdZb3DuIQhhG
Dxk8pbh84FN+eb527PZpMvuGd4o0I/znG5ctlG3BwrIOo6KZGTrvaxHOWE5I0uiSFR26yPLdsOiz
iHsLXJPZcR5XeEOODuZEmK1TKRxlrC9XvleTehL+8SkuPnErmQ1CkcArjXu/GEqnywJVra4S/nOt
ohlv9xsPiWP00xeUMcKH51ohx8u7NHL8b/TBWo5Z21MHKVrnWj7deSiLlDB93a0pPGvUar5yTbHU
dgDHHtg37tWu7Z91ml6O6fDWx8x4H6uOWK/ItB5y2/UxyU5TYZGEHZghh2IACNvTSXcLtfHMXIGX
CxtuuZV4/01qVnS+yDnLAabzNg8G3WvXBkRBkcKgPboGQD7tQHx4KHEtGCDPtsR2FGww4YtT1eFg
vqveIQx8TgGifP+IGWEkjb5qrpGedmKNMTIy/1GjBOwoVLvPJnhy4KAmDw2wg/avxsTe8BsLlRab
Fxo4rnOWWbPNVebzPkBTON8PaAgitPv6dhxcCl883Hg1dubuPMNhYexkXbhadava+RFGEMBd6vmz
HInmXVcfA991w6K/LYrC5ycX3aTRULEjqs025VpvmPuUn3YLYUgFteR0MScaaqitzl5KxI9rOtBJ
Tx8qzWRIn9T06dCuh0XVxUmSJkqLiiQMMOrZFKHaUVj3qyjkq1N7c5Zi1q5IKMC6KJ9xfdTsaU+k
VW6YIgEx4mKhdrL8DK5SnctX6xANnnBNeqq7XVnkkc/3cPOEjPjel8BxHk6CeLSGuSXCaiETEffs
qLAk0iGf9xyj3pdIOYBOCAnYhBQutXPFShuXuBOa5EMjnYFVd/MZI7c6Pi9bedEx1uhexzml5Zb8
zpZjOwkoXKbBMYsW7B+gMRQ6KJzYmppP6gf/Z1dVzTGbjVY4IsiGYDwLgs+CykJfxnklQlnOasVo
+wDAK1tU0dJkMTPLbFnBxcE9PM1ZtqqlXFVzrwPszdNGK8UIcHb7t1FCL06IK70Esbryy4FjccIK
dstiN+JE/PFnkDUA5MS1ozvK3YYVyNg1Jjsk5NG/DdnwIjwyeIQhDlZtfQcW7tp7RDJZf4o7AI8b
sz573tkhWXkrDWxtg7oK1nPXOD0ZoFCMEe2KYmT3nKOFeVomGJDoHnexIFCZ1LEeqsQh/3pNQkPM
nlkPYoj0YYyWGQezvK2yg2xrKb68Bo9yD48J6g7kMO5ASo7QoENZbhkPb+6pwQtLinCoDBv5/VgW
SJsNMUvEGLcY/8p1SFShQ4Z3rpHISpUsUfXewpNr2yPiqdJtr4US5H6LnS6BUzW5GGR+bltcr8Ld
KL+YT8KtO8EwJT+WWYXI3+tEdT3faTvUxQcOdtSEhfk8OIl6CIb9Zq/wNm/k+HZT3oapE/Fo0/5U
GqoNgSTaYQYHNt2nEUniYzub7V0lNC9CSV13ugb0+P0n/Pa166JujVWJVmkqimzDSDL2YCe2Rnx8
U23wlPxZPo3ESSBsPFC4rok8dj8tmqBDAbH/5w2VkVTjp6Qu25GDzNetde04skQttBnnkkIbjrZa
2KHJd/eL76OQrT97XX3wDh60CFAXCA92KueAOMgxaMXcxbAoUHT2N3BvhRN5z1TEtLkG9Ek4BcHr
hx+xOKmDdLlSJkLo+5E9zX1/SQyr2mqgIoDIo/g1f42P+zwkFyXScB+rcbO5kUAG6+7bIds89ZDH
M1NssuauPkb4qkPS3YCG89Icy2x8QW9xD+3ZSiQG+PUsC2ZE0/tlrV98gsCfo6f0FMTIhZR7w5yG
hIUQLfk5Wqt/xg8O3ahob8pUT4x8UBgdEt4fFxjP8NJnEWsnY2WgF6fAG9oLQatUFDiHo/6/Bh8r
9QcN6/b98NSqaPpkDvViamy5/U0Q/847oinoY4RqiEf29UwcVnC4SbCvfcSBabGfbZcb/XA5r0u5
SSS/i8KHOGffzjVzftGoza177B/WEJ8LAzLkLdMlMoxbNMzek/4tK8ef0/WoV6kQa+wEpOr7nYbq
Zw4R7YneQD57LSMfyJ3DpFFDubfiKhMgB3PrtQpB8HtnvVf34Oqx44N7lw4+BBr5eLF1Pkn4cG2i
Y75NDZmqiP+eVFp4xouB9wMNMChcpVlvgSHfdbr0bc0aBu5LY+IvqmIdYDfb28FtFmqbEDsuggoZ
ohqmZD37co5l9KBiLNHoNHezsRvE5TPKmlI+ckiZ7mPmuZ7yJd3bKdwR4iJFwPYGUjsGma9fmhDF
DlLBEYPSIlzqAKw9JbVjvi4ctAgn+2Px08zs5VjT4YGzcdoPmiHYO+XJyCiQk+w/9CBahRxZtKtj
cUGxwbHtHvFVwlBhdUW2lsc40V6ay2k0/I+nCsVr2Vfe3e7SogGVh5gJVXogPZ7tJCG3t3P52kIG
10iVIaRRmEv1LnAeqCf7Qdq/2sBboxbRL3aDKfcI2fYWlP/ZipFxT8Si+QboE8QgzmXW5kwatnZr
bobQ+tOY1XZgHzAmJ/xavD88odUnPenTf8WUP+MnaQioYv4ZZrB3N6zNi+k8OG/3zDg/3xLenzbY
6sox8/pXu96vN8LYVW3+LcPkaJNu2qENa7fH5sArgX6nOj0kuXb1U2gg9iuM1W+cGJEcNJfnFoCM
oobzGjidLrn864vrr0qN0vq1+fxB/daEJY4Ap5WMVQljydRz47ukCgSlbskanwOuF4/4hrVBBEAo
8eYrTS8L1M5fr7bm/1Z50Kba0lROslqowAys5T9TpwW1wL+youWh7Bu1HuYdv3R/WCQplyv2qgYx
NXqTJjUqrqSC9wPKznzgNZkZ05HglRJ55T619fjPzLlb4h9tX4kwY5RUA1kVuGxKavlD2UTxfRhv
XD+g7DQNWlNbWQXrf4blV8AcVOsQb2bao42ib9A6Dd9smpWteD1wKzBHnjchLMPCuH3l/wDBoQL0
A0tej/vpLBAA4wa8bnpMWZEEp+d8QzYsdvgt84zXK2QktkkspYxpY4w6+Qr7OEJSncG5BoJRbqFi
L2wJurJMNgbHBCBzx3nbXYX/EUYqteJhwVi4tYubq6a83Vc53+YnUT5LXqdxSl75zTo6kjY3o7ql
llzP8B3HQAZzI24u0pn9CrX1gpNAwd37HkJRhUaucJuQ2E4fBCij0q9+v2vKqQC2Uu+8bsFy+06g
i+KksrIEQNNViAEhwg8FB5mMMVeyy6rIEKbRkb4SYXATefxzZJnh3UGLcu+h7ZBNxRnD2wmI2UCQ
Ngq5okI4MzbOLb5D+SVwlFsNU9hZOT8eRmD+CKRPBd8fkYcg4f2hQuJC5oA0S/Mx42ghTJistlGj
hH/g72X8BBV5jFt9QScIjWVJw6FvxGTTJ+I/yY6REKlu36Bf0nBYK+T1CzxIh/aZQ7eej9Eiz7jY
M6EI4hBe6kENkOYvsUlz3jYbDcBtOhgeuLFKoQ3CW6N09qB2K3P6FxD2R+rmVURzvZhgwanC4xH7
pmxWrNuCeydaRui4EZGHAynw+6qGcucFz75UyTdnIS+/UnR4MugWF6ZnqsdBU8w68zkvPU6EON0w
E9RJcsZg56vLSvrr4UarAyVRBhxocn7taD5xCG9cLk7wnZassgMuMU9BxIIg3OCF0mOAROPcOYdm
0Bt83TNTXBPJmThKi+g5uo4bwpz8XgrjIxKxPDm+37XxYfLB56/7zjgWAfC7F3l7QilTMlkEnTEY
XvSYP2yoJ2sG95miXdmR31QR0b65geEtC7Hg/QF1wfidTFSPOrlnJZPqjI63hZ3kYEq7HlnFu671
QysCeJEIefGr7IbpeRRWbYTHKZYehvHzZ9D4uzJyCQEBmbxQZWuF88OzgGnLXY9VpoYGKYV9yqc+
ZAvByxjfbDjolaOtVUghW1eF7IiTl3aGL9cmuZ5TLSxVuYzw4B1L38SeiBehuGTum1JwJi6cf3c5
ig3Ia3JCeVU3RPs1Aqm0NSnDqHUjD4VM24SuLI+MSvzrwHphORo915JH0bLkqOVv6M4YartEuY2E
1EWcNVM9MNR5XL1tGpeB0k2igsnk5FDqI9gpocRqcDjGHsLXlj/wLD0rptBFZa8VXyzE6/KNBY0+
nvTj/pJ4hJj4LWpqK29OlZwxiHuo57DAoI0y7912vs2N/A0x+tGwH5u/P+Wl+ljrcNFAPGe8R6rq
EyKB2SiB4f2M+O8kenAMlny9iyuTW8CdqxWtLIEQQMINc90O8nS1SVXCVMlM+cyIv6973B3zlA5I
8tf6qnvLYF6yJeDVd0ZC8f7/Pb4MHVV1sxwpohi8cFXBDMcODMHeRiUH3CJZjnD81dF/SduqchpW
uyiQsM+7ZViKFkKHZLDeM6FKZvgPD4r0XVY2krWW1uMJkb3sG33a8EGLq+K15FjguLuNE3PHSbUc
vIQ5leED/YxDh3Vu+ISemO8gzf9B3Fl8Fme4Qw/R6Y3MIm6L4iQldfzkb6EXrrNpYQOC7MXRgTef
Oh7h4l45uN0lSONVaPvcyqtJuh9q615Co0STdch/2/RXx+VYDWAzEOeROUtqZr5VBlljma9APtJr
udU0yYlFo/oRRXdCuDMk2fjCPWRuquy/lN+yj3ObYRolPN2H9y10eBm093CKtgHOIDDN2k0viOSC
2a7U5Z+BZBeKUtrJ7AfFMc5zakmxGs+YVkfffCixZdynWnynIucsYpEKrpf77HG7qZSo8yjB2viH
BxOg6/GSyYCQE3UYmN/vGzgaksaKrnkNYs+6R5PDYCNA1RXxx7n3F/yu/XT4V3Qa1GQmzE3dB4tv
d93M3I+owkqt2d7ux4KEjqh4Hu66+JvVixYBzyz6da8KiY6qqkPitL4NcpnJG2yJD/PHPrvtLDZ2
Btj2EUi2bBWateUcNl6MmoMLosM/klE/85JOF5sdiWzhudSZzjCYZKjCdits9033FgBfXzVe1v2G
vlU/VPtjv49PP4idBxt2VCIUngbXICRLk0mXHIflGrE5iU1jd6YbbdElfXqxs6zUV59xJ0/alhMY
EnwU0li8pyYOtG5TYZL1bt/LwB2gODU2k4ARaFL/xsZMT8gGFcOKSs5KQNJQO28W4HHLUlrBh+hS
9pnOPr/dZWlqFLECwydfe+uxacstNqtbECeBovDBl8IuINGbAyQWWSPNbRCx/Ksfusc7pyxSW5yZ
8aI2WxVUp1MOZ9Hx720J8SfOPit3hPkRnnDNUHNRO0AZvVRwe45YEQevaNKmWNPgDd7rzL/V98Lq
5izB/lK+gOQvinRrpABD/qVLpAzcsSJgplNJbmLNiXaZgXjkLQ6kLzsH9WC9qEtkwYhwMlo6rbBv
fzqFRr1CGnUB/rgW6Xj5Fw81/REXRjh90+3/x4mjc4gR2nbkGOhFfPH28OvJF2pmEHGnU+QkILDY
MrKGUGaGjaP5dxWJF2nkwhGJznpEOI4ZDCX7i9IXNI1AoXOC0saCovyulRN3/bkHtK+Nmet7kVWl
aUsPQJpftKkI9WA+uSOqhNIIXZJp3DMFqCTJNLmq03dooGckJ8b6ngo0ePo6MSJALikmtEq+zXuz
+8YtU88i6HFdZ6Rus99bqApvnBSMRwJIw38Vq1d/Ho//Af/YdJVMQNRGSJwkOtyAHyHR2r1RJHTH
RFjcZfZevvvhNqg2/noWksvwxOutQe3eQq4w0xIwnyFN3CSDT2XVWPOfCbeZ4Z0KB+1aIOajUApV
+cz2tU89EGDX6UQlIo39r9G26kNaxiadIcJwXtBdWdjryOAEU4sB8N9CyF62sLfhGkGAQx6HXp7O
HpoOGpGMEmik9vyicOEwHoDUhHuT4ec5DBIoEDDAx6sZlGaepbln3Q9oxXF4QRFxS58Fs1Jv7DyY
x3UUqop1RVmnSlOXWNixWXoHEg0Yfs/fTmNQuIWjfeAwsUR50cUNBUtLOYWG6OLkzyGi+UIl1eWC
xQycS9ZqxiD9KgRtlNI/sYQEojNRvU0se5RvufZGkxPT+8Bf5y103xMVBYu/fCn+ShdIs4+03P5Q
bHzctwboGslc25RORgrFm1Kg7Ruo7bNkZjNDY6y/f16qR3fR93Knd96P513WcJXGVvCJLT9DOjIB
YhhhlRMJpJzHTKe8DsFBTU0=
`protect end_protected
