-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
d1E7t9zP2UUaVsHMTBsjzuyIjuahwv+8mcLvxMOGUtK+zriBhElTWLyqfyPkdmeDjhDV9hTU6ODP
VNun7WWBmw0sDmywPC6cR3oz8/QGAGWDfJy8/4Ho9BreBJ53aIld/h2ylo43ppJdTmFjPxWNu/8j
FjUWmPWjZZlELPyBTv8sZer3ou0zwF5JMmXWOiwE2dLSZKuCvaeLruVXaE2WvSUeRYUl/05FAjOz
Dd0yD7WrmznyQxk9GpqnWRt72p3QlOFoCIz+k/HKIUD+1Lhu7sD7z/g0HhJnDOjW2wN9KNfry2Y9
/6dP3gRx9XtHT8m1iYMn2WRFXh/KJX8T8Dowig==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11952)
`protect data_block
XevYTulHqz6s9rLIGgXRuj/vxvUjCzC0noU6eC3SHbeYuOp2H+D3Bn6w7XgPSQwEcTq/YzkcY/HM
yIgUc/2aobIgtN9cWp3F3I2MBBBbSAeDsATIrbpQC1K4Wp7vL7FQgXKo4Ty37hM7kFqrO3orqQhB
KNFT14mMmhM5fhzHOW4Dmn3qy0lxNZCgCflpZciES+PZdgqEL3Odhdo2sPVbH5iKCj9JFyOKf63s
ajF4kNB/Wybwk+ssKaNrIvVGo9oBE185CtMC62TDuSi0fP5zYQHKQ+cdWoaLzVAWHO7gpOQ3TJz0
yK3czmNbOLYCo183Xsj4TI54JVqVS6o7wObWppg2XSKQSji+re7gaFIBtWtaO3BQr2qpm93c13PW
vNyRzzBqfIiMrje7I8VIv2DqBc4yx/LXhN76ykB4NKmqiQMKkk5iazSwt8rsKAbw1d5QfF5lJQXY
cq9glA0LvYa972J7ozeKe2R7r/K3fvQ8PKW8oTb+rPHc0oncYJUqvAOXc9nyl2GGJKZ9imwchUOH
ZBjHKZ3dgO89JY/XI4+wxOxKKUgqd4gCqzdOkt1o+RLP2nF47o8xvdAlt4dERk1qDmyqyVaKW6go
6sNaCx0K/chadvaZyeRs0EYZZHCxz2SJlz0u4/JQ99lpxjPVc9nrzAZ88wFykoIKC1Z7V/vkB6bc
MsNQGUQJ4oKof7Fva30fMkPHkIOptJv9uvEanB+I1trsP3OIC1GIzZdTYyT4w1fav9fnDSeqcE9t
LhPv2eLTq0FgepSW1hmy+FVMuPK79jRKZNLo2iaFuqLWBESRaOsA4mQtOejFL7mUmf8kzugC0X+j
fFo3R+xDyW3JKAluLn4GqcyzKhDHifR+8Fy3XETUA7Vo9dN/xGi+70yBAKAm5InI/zBfqcuA5vmT
STr+rOXMTH1AcummUziQBOcT6FTCUdYluQle9yf7d36sWcsyIM1DxPQt92OWNM0Xiig//bDGH3jB
I+F2XApmlchB5TYI9q0utEdGEOlkbo4EpdVSi8b4caLRIJni0uje30eYjSFhyQFoHe0XjsRgj3ka
bdXpJBGwQpkPaCYLlziPX7C2LXSAMUNROnnt1Hk24Gqza/vDb6V46bDY9bOYiQpI4SmazlFD7HQ0
rjLCn032c2RfakDA+ZrZniPkOg/JTIStKwMdZr41wZvS75NGiGyIagpxn5cBg70OI36bcJ+UMojf
8AJtzFGIo8M9ehWTsAM5Jdd0JEcO43TEjRSJ/2wwS/80DUdZafGrCzYl+oP7NRh7R1673i8xSrsv
X8T+giC/dSG9OpGdfgn2pMa1SPwKPT+mZgFAZNA36kR9N8ZgJBjo2qJdThVtPlAB+hANMhin2IZD
u8eGeUvs8mlG68ls/G3r8/CEBjBYvkVsbebGPKp48QW8mAfWywcb7zplZEf4l30vx2mlxGNVKnLm
mFc0gOoEJ8+ZbunuJg/mfPgJuBjSPigJD8p1L6oNIvwDBWF0ef6rMYOYBE+d3GkPVpsfknws1gau
JDMHtOZGr83sVK4ucDQhQPDIz2zmjqXeV9BmInkvMivftLISQUa/mIu7asihhdAHHptDDKKfbBt7
LTGPQJpWiMO5CO0a59emDdYCg7L+7l666bGlod3oqJOGhKLdUwsi5jocWkxlPaNO/DrKYEke5zgY
ei5OJ6Hy2+3HKquUgQkhBGRnD1sIdZtA7LhZgqMBtCumJADrKkXYkxi4UZD6fS5YtCk14Kh7RO8e
CEU8hnj40V9mZ0xyZ7q2MNTKLve29Npf3PjHyu6oVnuU3rPdvkqZTt1Hr7RW3nrcNnC4joWzkjIP
8JUwfOdg9sZLthFn+hHy84IvRcj9Y9b/ap6otWCkLlmT8XRuWjrIx6yWJrliFEaM4uGvnUGbHlHa
RTu75CmYiH20JA8Dhz5Fmd7GseBscpfWxiyTXiBioVFPhmCjXtoHuu1ThXShf2c0X5znONfLvNqE
UPgyitaAAlzk+ms+zOEG4k6kwWWYvRATW7247bI3cuPT7WGL1YpkkL/LPfMKQOyl69kBHM/91Xkm
dvglk4zOVibfd4jKdAr4NeDx8CP4UFHLm+6XGoiZqBWtEhcLNiz3nAaAP4XsMxTMXl5VGbVylSgG
vmyPy2hmb0CQTC/7NU+5YaCjXzCsi5XYo8EhCXJRzoVQka4DuaVg1jGOBRQ9+BA1Xw1egNyrnEc9
bswbTjkt7It2ZWBtihebRKWL5RN7IpouZtjpBKvXnBtm0Mga787MUZOxCPz7BJrqdojt63nsfwmL
VmOGAAtQv2QUaDl8bX+1fd/1P7rpGAh68Z81eoL0GzE/lfJcDGrtuzBiI5BA4KspqsKexLbUL9fv
GvxpdnEhc+mqcC4HEBXnQvU9xJBgLoLA/Noml3bLkVoFiGvFtkV0e0+ZuqlvV1XGp8wnCqaRAAT+
jCkAaW6ujLBr5Jb06mVDuOMm9FtoevqHLLFwnHFHIGx+cL2l+stPYQLAPnPMZSNf5suU42/B+s1N
xNRxKHkTb/7w7kHR2f09wSh1SefUUDdP/kB8/uixA0QksxiH4WTKIsK/AgFZOvRMDxfBl14o8IUw
I4cBIm/OUkOWWakk0iztQsMnPaQ4dAYRW6zNVoqxV1AAvgntL15GqZFt2PyCa5ivqDeuGgIH5Us/
tP5nzlqe6g0YPJToIb3TAHCrTwWLHPom8r44AA2AzKMY1/GkI2b/gmYOsEJ0pWavI8SmE5S72h80
m+PW4Wv6jwNQUqaOfIIlObb7ODzfiYt46jqlmLHUdqrYU+RqaFuzVrkyM2qdBwspvbC+VhaIH18s
jUlxmOU80+l+/Eb3O918/oJsvH0pZHm6hex78eak7vty3WWb8UM7nRx3TyvGrFrMVIshWx9/okp2
H4VtA5Xr+/IeDVX+gjWvnWXSX+chivJt3hYFyyujYo38IlBEo9WsCm1p4/NfoKaZzDCpy3CvMrVb
LXHguf5a7c6F8pr9SaJ/e+jxjU6mjYGimMwqZl+bbyG+DG7hPGViPSnZTjO8tgkPztalT70QchKd
p07NEcGlHTTpDvX90COIUAubbEao8qC8Jd/EEBarqatgjA7V4QGmDCuHVahlRgXqMFqpZOCxBuhQ
LuN2hdQBmb9dzlNStR3Q7JeVldXafVEiy5BN4cxA7rZqoKdUQuq+tfJ4OQ69ysOV0oUNR3f4Vqpn
Xi5hLEtIcQWkzm80NDdmw/BeDCOQuKabOTy8HGIEb+EYzsS1glX+w4EMT0NZzao+FhTqEpUhFcap
dUjv/nPBp5+m1d7FFAkqtGAjuHFzQadDmRrzADHIvD+t9WpRUvTKEpq7ycWKYwkx3AXSYB34/yvN
K3O5kTrRNbS+yF3XPv5Dqr3H/5/1toahcecIJR5J+QXwNG2YT0eCB37rdAojnxtGh/qSeeI2NGyx
H+5ONIOOFr3WJPcf835PUspZYo/hFmNrVwIPb+pGlYEtOaaKONDP1gRQ2J5D42EVjQPUq3Xq8xwc
1qwQubNDi3ml7WGSFXyBkoiiX35fMfhtp6qU24LKLavu/sqi6OwMaXL9mfh3jqqK5x0WwZMxifDJ
hskp7/fwIX2PrbkjbteJPHHJo7UgpkmiZODMRtxdSrQhKE8R6itDCV0dmW37zXzK4brTrbGxTZIm
bqggXpwtAEfdllYfv3nhYRHvjssoYK8P2xf4OSimYCoZ1jjpy2dW7XOAkWivzzmLIHqwpI75Rxy3
yuTC5XOVEb0o0+/aq9s+6QaRcUZkjDHy/3MFtSVvwkzIPUzqhaRp9CHT8DJv7THG0mkMnzVMqQbn
BnL6rsurNffuv1r/pPR8eTmmoHswnzD/LxQ15E6xWE7PbV+IO7nO8X93Abw/ASpG1CP2Uv0SoU5A
/th+Chl4lG+w/EelUjuIXt0lnSLPp/rwJL2gVUCAmgPALAd7w0pkHLidDyKERBNyZCoKcTfTablq
vcLqCflG8S0d5P1j0gLW72BcEZnsqYquYMMMvnwRfYhQxMd+Vu4OndYUyUlLiM/J7k2WSfJXhyCz
JhOttAGVwOvuchNIxOV8YTfKbf0NRxMkHeiS9UF8o/g1BlcudehT3FMCcWjIVU4+CJkmP7AwgiZL
Mu+el6InqaM3Y1JTTXq4N8A4j+m+SA/Unp0iraIreGNMz5qgyrQQzlkAVWEzwsGmOCNYGyHFHEBO
VQi/B3HuM++nXIpD9RFyaHS7Wznr0GJbcOkFYoOqTZAFpt++VGRcjC/HUZq4Ua+zto4kNKIQHVSk
/h0xM+QLcqMfvp1YRJzhVyZfKGAwdcDr5NI/tzsITYR6vurD98kX/iUDlTJtqQPYMpId1r5Cadmt
JRGG0u4RT7qTVSfcwxQOy+wcoCnLWFYr0ZLTv+JNbkba0ntgDc3AeRJ2WUFA19UeeqV9QW0CFWWl
FVdLf9Dpr3A4E0M2k9crkGSyHl06+vwXXw5HCdB9OHfEyRT1rzQTFdzCh3XBBCZ+W2TfAqEb8aRb
kUB7hUTHiaI2zDEcCdRIycN6Qu3RYPeDEKluvT2pnwRNjfc1hRUjDrj4UuFmPynCzsTA8zISFuWX
GZ0dDZw2U+4BfXpTF0ebjiqhagE9xag0pZKyYvD112f9xyVd8A6UnnySo8ENfN/z3Fg+dfdBgLtY
oBCKh4xbncnwzMqgxEAajXVGakF8R5e/eEJ010ULfjLoQLR2TQfhfYNkDSpc55q+ircoEG675OO/
z+t/s+v7OKVyd4TIWGDpUMfGKXcVPmnGQW21UDNZPBTsS8VBc7te+0ATOc0uK8aR0IkW3RI9q1fV
5l3mPZ982StGDd3+CPnLXopKmTvZE0fRP0fZSyaswsGVvKp2NH3WYeUZH1MzyrWYzFqEcxvzsnmJ
ZB3Q4sPkLZEat2W2RUECuLSSFdJr106UcBP72h+vwDqRujcbF8rtDJOmbQ3TU5MN2dfJZQVddzbh
Rd3jkP7pJ/1KMv09wuofaZ5etZHGeIRB8XWN1018+qwnrgdRObQD+dl0qU/f0S9lFO+LxsZ2YN9z
fyn79eTNgBywOd7vB8v7bZJGjO1otBECVbEWS6RG6dpscODBe0SF4l8kyLCvOrHYsld1bwpckW8+
YJEFdBSbRUxJYZ3GgFmxbeVGQZ/aEYvkaw3pycZKgQIRNKqHm7Yk4nIMNWe11vXnckjMxnrUWyO5
g7up2VU+QhsDJIoIWnm2PSZS8FLGu63ugg3m3/2LTzBCUwq85CVFJhlaKjBlEylLUMl0Y0ngG/Hn
bJXg76cDkUMIXX9u63O1Qy1/EgWbZ3Cqdd/x/DPFh1xudwiFmNkAetLf1dzc7Htnsc7vJuDvqcaJ
KMvcFbvOUwVvBlxKyEci/czjzVF/8pTnuR5GL6TYBvNWSLS3fOPCpgXxjzbijysw5qjmyxLasYPX
7by8y/i5+kqr6quT1fqZJhKfKRuJxvhbZ8pRHhEDDHVxHDB+rxGYJcpQfQWwHBLgsxk+23f2472f
KVO5XexIO29t0PBwqVlGlaFz7eVdYGDO7OMQ7YCzRJHsqhbdolep/sHhCGGSr/C8P55qbW2AK9D3
ZWdnCsFoxUtYdJE3iyV1HhemoTLlBj/Z9bvHixvi9YlDJ/P9IUkqxChI8E+3rHnD8npBPhvGk2Lb
CJ2RQ2ba+fR8GZF7XDXukOFudP7YghjlF80wG0h2W86jeMq/haTHyoeYzilyiWAKkGoMObjwho74
DXme05NG5mtcX0U7Ig5wL+4abuCoSr+vJtnaepNoUHfW6jfYr7zXBjp3jCgeKsR7r7uoTVbCWwPE
o7C78wgTo0f5wKvgniLp3svMcDtJtM/EZ35RMQRot36JapYuRtWLPHEy5gggp4ZYzjrEisIMZzf2
4J54nt9So9PryrLDPsaL3jGktMT3pn4BXXiBCe9ly//EG/Li85z/5X2XBg48K3xYjC3RGDuLxBEU
xkKJjEsx2mlR5JhM3pai0KA2XS4iRMC25UbRWisx1Rd/hHGIdwAtuKlWmKgtPoZAAhJd96cAvqHV
0q7UwAgUnW5a7Q/1Si+z49woJyyA6/UpV1XqvmPy36g7TYLm6jJoZk+gi+v/vgt7aOxvaZD+Fdky
ZwP5obxJRJrc4AmbsibXoUkPTn8j3igC5NVCFjvBpCKxdsExsbg4FqRRBPt4bSqW9JJGUWNeJXwU
/kgyw9MBLbYX8uVPsFnxsZ98YygXA2nHqyC+4ts4G4lg3x6+nF8/IkK9X02EkRm4Kqjw1biX/CDt
sXDYRvZCOsLUWFacplZsvIOw5UanDLSyo1S3eNufVhFcVlQiTjTVEo58297Ho7jDWrVLwXNQtc0m
kq+pVaVGY5DP+JTxVHI7BDLVen/hUkKyYDeSTXzzuCi1T+0XW0Gzyj3wdHWiwJMfUSByiI1ALixA
1uI561GvjqsetECm6QAGZfkPswf8WhzgAT6oFWz+OVr677ogAaWY9qTQhT1Ki5690fc5eiGjrlj6
9j0cjaWf/obayKisia5/1KvPkHrqV/P9hBM9FzXkfSd3qHdtthDFx51IhsJuzvVdhlTNBXwrR9Zz
crZIgkfVJIc3sx8oQKBxLtu2B3XzMB47YMjS5LjVJy24foRNYi6deVtav/4xoNEE5XNJBfyEjEo9
JNaFTNM9DwTy9iqWtrhosnBe19y23lnDmNiMqWFm5OMiH+VuFJ98VJE6zwT9ySNdWYXYJJRTwBBu
kfs6qaGJ/MZHZoalOormUPSFZLkG9mIzdB9UDag74JFoTtOALeCQM71O3/ja9+xlStACYJBxxxwt
FOomrIzFEhuacXi+sjf5JEZIeG2J8rPJM7sGhgpiITALHqfZMVroIjQ9bnzdEllZgUski6h/R/qf
v++achsf45CCdcyzVQvweoJEek7mKE4L1tTiCzJchSa/hiNDRrn7KW1JfX5NFSC4whXWa3wx0zJh
cSszpzOPvxB1zVqO6xlyxJc4H/wEVoHmgV7DCQfuZ2v0dT+cWFktga+w9ugOOUEElL5aJsA8HAkW
qTjotR+Z4Qv7Z1uFXn9NMLpKn6soWPUb2gQFC4rFreRknWzM4XA05eMocbIpHpdNpSCuz53hxRzq
SpsrcL8Cz4Ui1neI8oksvLGB4IYQ5dLPzcbPNsFKCQiJDbqU8CYJNAJf5xqS7+uSTTq9CsCdcOBr
DPC5pdQe4KV74iNqzFJqgrTtQHvAqMt8ElggzlP8M2xdMBsl0CgEbOxfZKoMZYe0aUNhDR0uMSdF
jFOxMcsfIwPryhKz2TikvyonfVOJgD3keAtvhS0BRcU5Efc8t4MSYhpgAaVxJmp/ZQKJ/siEH8Is
9j+Nf3H7DOAxNtdpjIX8QPxLzMPI3bu58MUJCpX6mptbNZ2rpDHeLEy77bHn0jLzAUDFSelVe5Nh
P8ZRocT/LNR+NcYNfdVcbwXExuWsMpbCa2aHurmR2MBi7+zqyukvi7vLzXVekfO+qYk4pkqAbWAw
6WIUZ31dhdOt4eE91o5NLosuini3vr/2N9gzT7KOpuKXMTgxGC7DVviInDMTHiEqx5e9IbEAvbsd
faY4s2Bj0bbUWEVOs8+lDsVm/LMOGXdFQncIvTM8wtcbwlwZlnrXpczk/LxsMZ57JZPOKNjS81yb
wcxn2QWmHA+6X7Chs8V9MAvTL2h6Uol7eh3Gmho4UgU+cn6d9xIq4neDdftwn/7Hz4DhTE5DThc5
HGepQL+OhU4BFrTnZdlD6ZDuRFsiHkXUtAy/FkPfSSUW4x1e9j/z/Uegppu/NrgR3tAFOXxAAn0q
AfWSNB7ZI0CoMdRz0szA62A9qZB7wPOXWotiIAx1JEFuSqZm0Vl+dVhQ887qXO9YqK5bsU3ZzEls
anW0wr2+81D7MfjJk93Gi41du8u+iEOe/Ss+ZoMcT5XMJoj3N9KcQWk4jgRTgW59zVXcV1uLnQ2L
mEeUOWsmQe1X+XPKCbFW0O76BMEnII5Lqn/WUrY1mTJMVgrrj5V6cJeLYG1Ttv7Hjrs9oRDbR8fv
H7r/1Mlm0OzhOcKdhLKssbQAgYF3Gsg3ui9dcP7Ujcn2tzhPGtBsQj+EXmZAGJlJXa8GAdgW7/Oc
q/6XDVnLpiCAt9LBM/HsBfY+BNWm1Iow7KCrdacC3GvoU4FcT5oncAuWM7K92rUALLU1gqPEpUuO
pYmutKxLsUJJ4YHjSfeCXAeg/tJf71i6wHCWk8Ldp7+Vl1TKgChEjx2U+7GLjRBHR/bW3lQwM41A
YummAVsQgng0r0suScF0g1kXXFviHmZh7UPWDkya/B0lppZJy/4JX1MUjAtmRLow9o5HkB8A0z9A
VFAAZKkPHgzFSmYeb55MWfpuqUEODq6UgVvCdUvzfxr+sz/Xc2h40GqBYwOuzwD5MhDAh+6uZPE2
EW4/10nw8rABNm8A2iY+t1cUVZXVKzCNjEPNYrqTewaUf8sPMwoqteJ/iUNmay8Fij4BYkR94aDk
2dW5yodnE4qul48vXkrGTEcGccCzzMa8Jm7mKIOMt9NO/V2Q5a8TZZzHAkQIMDdI6tR4tX9Mic8M
JB4xI3s/zy3uFYK6LxSEpS+NEuOHtF6fTDqDSPRsDazm4Zl3x4IUoMOb1em+qnMB/hIXT8weEd5X
LuFZLNNPQjxr7CyHfjV2WxUn1MpFPBS8/WV5WJ8yQ39iEM8NMfx7qS2G2zlQ7yyGEGXgQInHKfF4
1tPV9BixYwyRw1ga+3g2FI/7lccTxVtxUP78eMma9o1P3FuFOYB0DFRXRtR5I6r+hKWxxu1FYhVn
l5uolYu5kputjGDmbZzIFNuh5YEA9TmSFiC8WewWbPIsI9dccXIHUH4NRE/1oLqJdccoBDh7v4F8
sdSUpHld2X+85u8hStBp+X1SMFLv0GGptW88zeCZvp6GMRrgzURH2spRh+8tUXOmVOXaxi3AIqWl
3VsvdFIh3cW6uWg790SNiqtIwaoKPmQ2YA6jkiS9UbDrRjrmV6JZe9k/uIbO69fzi2iAS25ryZZ/
iSCg8SKyByg85ySS+lOlsc3C282iqjW4RfI2Fk4zWEBgzIVBYLAVFOXHPl8V7nK0pGXbIs+n3qcy
H9XGbQiVqtUplDVLkWg1umZod96+iMZm6GOsYjXJD0tUZtq2gbJ+sfbaqnV+Qqv9UUCMwWnHpFug
9R/yoNaQBhbBP7XC3htUQmDCQXfRTLMX3X9m9nCKhfKC/vk6CJaM2pI4VjevAttUp49lHe7B81vB
GUaF3gVFvWF/Y+dIkaTFyCaHprG92Vs/NWk0ia7tLRNd+0M04TwFUuSJ6TgVyAMitbM3fNI++wwG
snBAU4j6TWHdugfLlDix3mJhCt89ohQqca7S4g8U35vqxEXwV5aa/xtFMV4BsJnol7M5E0fivgne
mjVNnvBo8DLXShG+afL65A5RoYfH8BJjI51xOxvrLIsTsu+rl3txqXMpQD17lxRTcCpe5UVeaJv7
NoAd4fZIFqIfDOA3SQb24J3jJqf4OzX7+2KdeJ/Dx9Mb5PSzUc4/0Hytojr3G2IS6NpA1Ig71k4X
JfjERKEPsKuy51adCblyXl8k72HWBc0VDlbiB2TcCQR51xQR8XRppHs/3mQX382/3m3F1N/KrNo/
Zi86OGOETaXbP0kPhMxp6qfa9NWVPiEjRRbAbKvuSaAX8y1ye7TDkp6RqZUo27BO4QFVvxwuEKLs
U6DwzLVg0OrE/mcZV757W0oz4lz3kuUTsyVZhtuIUh7fa5VWZSXtqpEUH03eCWJzv3eM4t4L2dTV
Cu4WDZU3yNYzZJShh9G+t6ClNy6wZwjHhXfNMvoY0FMjbU6IRWL3laGpltkm2ew1TjN9zhNedAXM
g2ohMfN4oDgJDmDEUvt6A3gqxzm923JirvOsmtUJIbBH+wuiXZ+VQ9UX2P9F5daE6x1EY5TjlUB9
O5oxetk3m+1ruDC1kFO4sqL9Wk5TnwYY5oVartlyLOOPEgJgjRnVyrjxfF3abrFEDnvTzzDivj1f
qSlT61qM2CpzWYkyTiW11mJDKYxI6KV8HkYXOjyLwpi4AAKHpxj6s5MRMlXKpMmbxLdTjooe4rYN
9Ebd9b63ttnX28npuHX1OVJS+RK25g1xB3rNHw69MnS16Qk0KQcD0xTp7ttOx2P+lQQlEg3RFuii
KmBmmWd3DgwksI5Pewl4RxABQD/ERnOuEenA1fPUuS0jJclQ2/HxQaEDDsgGBnOg22xJg4rSkSQ8
3Wf63QPqccy6w/Z93FQfb03GmolCNqKLgDRfgzaYbij+8OZsvp14vgX1BxezbtX1HcH/l0SG/hYd
1mBPkQGBU3cdonii/YJxBMxhKfpOAYdBDtHx9m3y+7topQYbWolIjFa7bGapyScntw2MDmOtYCaW
scXTAwrilJ4cG69USnmOiS2bnbXSXVHCKoeRTlwz7ynFZFm9DRyYuG8+hNhL/ow9wLwpigIm8llY
KyJOi6iOfId2wcmEes/Yex3ageyYUfUPB5qjfSTn3RCvRXlGZWv9AU1Zw3vMKi0wNGSZLHSYMavI
724/IElWyfIfDtfHVF2/cU8fx6LJxxDhA07nOPnNfHCtpcEVftLANuHRVEqRDMPWv8HYELdIhkRS
J/b43pGO0fdDgTtnX1BeyNUrs7rsy+0Ra5vhyxzSAVap+8TQ2hIxiyBJwzjfGQD/N0PjMQQsKI74
NlHQeO+GNzNK+54aI/TylTJRGVxS8SMo8Jo/B+1pNV7WfnDBOrfmYGwZKbHKr81kHFwFUmcRsklQ
ejjvUqUvSk4SIKw9+BHBDg9PEpsSdEOBbGWShHLiV3UEpicr46crEQEbx0WBJmDvK6BwvGSMvHmm
qlG+oEVWgOQXH0gJuKby9hGJ3UpKK8xCcx9waFoMr9znNa53hXLxtxZc4cPic0UTlBLXeOk4T5fb
6DyysSjYXImjiEdr1HYIXQRTP2wMTjveK3YgC3acg5+M6GUSEA2ptL09P0FbVKxGthFRul1zdY4h
Kg63MbjVc4wEAp1Ip8UUYyiPEPv7+xK/Lk1S9bo6vriG8onLlKYa8WXCn19gctj+U2S+tiNassik
w7O1j2J7tUalY4Ak1NdsFChvIKzBbIqNLm8/+BJmsLovAVGgipBehyPaGijPsKPv7UX9zi1v1coV
b1PBVMQ+ydhvnX4tcC0kx6sjLlm4ccbPyu394WvThwcx/74pNMDZ/Y0h/3s2xLm7oNKb6ma3YcFa
tCuHhfZSQiaD229OweYYiikRHo3AYYposxupYv7Jd8uianqUl8Z0QqwBdvNUy+luFlPqnyBrtRGE
Cf32J0/YtJNOMJkIrCL+Y15umletZYuOdJyMVGtWjXw+1TtiP04yAC4qTRgE3lb4ekSOWdnsbhDk
2Ue9IHqbVyadt1SZkDnPuFnVRrCmjj/zNtTney75+fDVAbVPyQb9xh0BT71zgUaB977+3CH8xuGo
d2CuocWTndzfjJQV4fwa4dZIOmxEtUCdrfuvYT32i96IXCu0G9ikmqUkeNUd9sQ737c3DsB/mBEp
8gFmZidUt6TnH/KZUn54W6d7HbU13ay5NsCuKeZXdohLnEeQ0C3E9L34MjI9V2+Zr24HWpdNGJr/
OxvLIjN34SOKB3V7Y8PM8IJJw3/keanDIZpHqqabv73184af9Ku6zIT+dtwV5VwPQ3BsSBZwJo6q
k/CcqRbHpMNIA6O7twGMzsCWer3gg6Q2ggPUMwB03SD+TI3vniNlCTsRm7+03yCxvETNG7eH5Ogc
JP2jF+IRdygxrPkJWjKL7YvbECbd8pYbA3bjv2A4zcBsKtMq9TIWR4PZmZgOJBxss6FJ6HBZlZFk
1iK7HYIcgzLcaFMAq/2cWFASy4EUqrXDma4uP1dUMGjm+o4CnU8lyUlcNv4/PHJ/wFCEgkMreIpV
IJSwYcsC+IiLo95QV6c++yFHH1WnEMahLD9kSlZ59VbDpopS8Lr92wewE35usX0gdoqMcu5jPI5P
1vB73lG8wF+VGce9Fme36WSIiCCzi63vA5wwZy3KH3VHHRDSOcG0K31PqkjtTal/x0Opgu/DrNw7
HuhiRmT/JtRjb5P+bxuJ84hSC9uMs+29ZJ8vHGAN6OnUYaQSiT6TUHBZMi8GIpMBbIhkKoSiGlf6
5Zap7ZgR7bmWbZZBhJRuuDPD1wxGjGXCohOMAa+xbfMH8JbgyxxAWx7qyqeYOJRPEyczZ4RtU0LD
mi71OTXfgCjgmtrlG/sqzwlfZIN7jGNWlwlMCIh4urCJvILPAeh1aB3ZdHCFE4SCPah4KbmWYXRQ
FdHB1FtC8V+naGIbQmCflPwpaE3idVzP4PGmRBnFD69O8HwdFI6sayAcHQiwcXimcy+nRvAbPt2o
BAshCsbcrjyM0veKFMpI+5HsBka83xvg8l9LG6kk0lznK0j6/gQ3HdPlQRp315ck9Ab13u/kd8sR
5GoWQUycKoYp2/YDzohSL87Aj1qLyqKzdxHBPCiJYbX5k/S6VJcnARV36QeFfbwujxFzrmLkpP8L
fbGPzeN+CCYgQwLIm/IuFRleJbwciFL7F7l4h9hU/ERv7eDAFYRxY6dfLfGLviifQA6wiZrADK2g
OtAXaESwXrkuZHtK2PfwAjgrGNdfqNVb8LwoPV4vS4yv3LXJDNK993dJjmt1vDh4W+59/6gJoVpL
60WGa4K/L3xxvFbkfDXQJjYvdS5NZOeXUpSoIAez3URMHEYjIzLCNAvI0Zr9MUqvBoO+VZ9z+RQh
W5ggK4DVK0+GFOY6+0w8UY9sjeJc7gpZXJEieYkqCV3a5zVXQnej6Ft3WDgzX6TCqATn9D9H5z7n
jSW/+fXWwX6DeXZCik4dGIR5Nzwl4eRtQRJdHV4z1iDSul0WZ9tnOgrmpeWjFYL2iNBzpeK17Pbw
XOfACnP/2Q++KfpHorAxtKJqW52hXvrf60zyIqSH4sMcvH+lUr1oyIaC1YoMUOuhRSnr53ebF3au
KAapOIACiLTsFV0cd2V/SiX14i9pJetAEX+GdtD6ulM5xcW/rfvjZbs0vuBS3Gb38pvLticpJKBz
j0Ss+j+3KIkybkx43BsROsdQR0TeiCd5o6SQhLpf9o/2Fq3uVfy8bnOMcSKh3Aq8HfbnbpwFW4lp
vGDenZVt5dL0AZcN+nf0ea6Z8u4rkGPpL5iTRIzZyxzhPBlq+AZ0jrZsM5wZJ8rz2f0sWo4PzggH
ZJkfy9AwfuY3SvOe+i7Xi+pRivZhV2Ak+ZazqeHm19r2vaiD/fw1P65RaiLHRRq8bKZcKKADYnWN
+aY7JsVppRwZDoOJrVA5QchtZvPsIbx3noWVHtuw0aQoLXO4wyxywD1SanhdqD4bbRDRmifo0EeW
4fXErgW3EawfA/b93KEVUJOz2uenDJP6yLopyAeorK2GAK5HPM5CEoklc2k2i8V+5kIHbZL+yZQ/
MdOituZqY6RV0/rT/0l+tIWkNqX/BB5vmog94l8WP2UScUQyrMZ0wMjAL984hs9hUdr+RwNqqTIs
KkXrbKjyHV4lLnb66RgweUYvgfPZlSTuI1Z0w1e8v29DxRJHkXHMZZCI3DUCn85PkR45UDDyyhe6
Yu2dy5JNU3wibNHECqkVnaDRGW7n9V61afWQyxL6naQFOxsAv/u37VfSdAsdhBaCqZvDzWAuSXN8
jbUKQdM8wYa8QWRyNqrDRb2zb2M91DTNrVqMRUAgfYY8mQggZFjU380YH1TWqVPMGKRuazV4zP+B
12vnV4rCsde9XuSqKt+Ok1kh/0VaV1aAxslOxaSpCaRb9Ip7l0/T602OEgeGeQnGyzhB6ydytwoy
scIRKlvTwAV54kfXyainIopHpTbJj0DBTItjWkWiPondW9bM/AaBdMkU0sPOfwMTEtdgLPzAhpvA
cCt6mFeIo2E8TmRRMLSY4DQ8lN1vp53JVgRNTqEmfbylTQiUipyfWRHs0w1oQz5c6VaorGAAaC8d
MlIdrrCcAhkuY/o2TAhkNh2KxpEhdNPbSl3CDXET/DHwoLWEjatuckgVJDByR8NKJlhMeUewsHx+
+sxTXzeUZbeLtbmdGYRu9nHhw7nzCqIOmyek2ccYJJJckdFyaM0wT2BuwQStTxFUUNo6haiwp1hG
KV75ROdPfrhSDiJ4tn6pETV22EtewGWYaooHWKBSC0ysl5sNygi0bjHt49W+j6UuNc0GRjRnPGsc
u6UbsKhSNtzzhtabBvZHJz/3Nlg34/CjaywyqEEi8B+xKLYHoERBy0FZ6IYPnp4pUWEFUZQGSVba
N+XWbfl15k6IgZj5EKdqGlLMc+KOJw4rZBaj0y0x35D48CMT/Y+e8clyuE0xNjHACcV14fMq/Qyy
TaNbUFtyilzlA01KO1kZfYcnuAXfzLdMV1teNqJqDQ1722l6EMsntxnopSd7wOum9ULQNnfe7BIr
Ox9IVRgDq2bQ1ds2U+Y0puYrVFhE6TCUfa/vtO3VArlzH58Ge4Bu3K7xKzFoGnJShmStuIqvoBmI
+u0N34jixg3UTEQlLt0oEg26cJmYYnD/hD2KZUdpBvtLZtH4EJkf37LpxVuv8EBEFM/jLNbnIbmC
aS8qZz9meE2Qz9iE750+WQ/fxrUY5yhwLhVTOZIhK/pCC/nRK/hunx8lAb2+F6XvEyRUTEkpxRsa
8gpSYF2NvPMuaBpvJGuGVhZtXKyWki6pVbXGchJolLXaXXpWzJyC6LISwt12tuxQaV1X4EnZKLPq
zYs/eXusAywCU4Li4dsb/hanycxweBHPwHbcJzIuz+dkXRKDIivXbYMNAlV7AItht/T+Y1/5ccZf
3/5nTAJOND5196s12FQG8ulKOx7cJnTElQovayFUuHh0hoxYpyclkqf/JUFIRz3Zs4PXnppM8nfm
rwNgAWpOz3Fnf4fZy1PugwEjsrV+gsNb/yTBAx6uOpAKc5a67Sv+WF4WQWYc5wGSj9PbAlLmVCBz
kzhYVtH4YTE0lqxHYrRMW50NKo/xD45i9nVUxExTv7jG2ezwOadm6BKIj6UtIbkVUcS92YPE4QOq
npMZ2C5co6mJ2QA5Jhp/kSqp1RTokC0ugxCPGfR7qP6/p5ID8dm+TFL13kSEkVI7ZYZNKfoKeNLS
iQXxGnr3E0jTPzRN3W3eBv1uz9fmAJzEyDtgWNQJ6iN253v90r3S0/qdCUptuWJuf4ROE8RbkJeX
JhnNsCxR7uRnKj8iwRSeRghPXlprApAzsOM/9xIZVm84YJes4f2FJQRtO91Ns8x8hs4cRUWUaIg3
7W+h2CaEDFL5YWTvPQEJq3jVJiBX1xDv73jw9iVSb/SbTsWQ3pwO/OBkshhkGcechNq88SU3+cx+
B1AlaUY0FiA/fgKl7Ae2bZRr6RFhsWlTX42XnIsFTsq637U6jECNaIqr+t4LeL0ojAw+3+wb7gFi
ivGGRET4EK48Fp5SUgy6NmJQJ8eO2KoFDzx+RpHxtKOwWelqRxgRymYL/LEwtUvC2E62oJhcNpUz
30xXhXmTtEFjpXyNjltQrweZalYkT+Ir2wC9M/gNeSuWXm/eLp81HPfMqeYFPrpsjCXWdbMU9U2A
s6mIZZFpChyXrtSR7f8gYJrTx4gg0vDYoHDUBNctaekT62pjd/BzHGHmdKMF2ihj/Z75IMKCelrQ
+SEChrh8BVH0gQtHAwBLAB8siODob8ukPMxkYbax5JZ7Yn1fReTi+UCa30j79nbtAE1YVcGPWh3P
VRJ01E9uy8JTfwVg6DUFDitMqh8x8+dGx6XV+iwkbumPo70T6826gRjQ/pPKj/6OLnUYgdzQ2amo
X6wSg99S2CYthUop6CBdAvzsKJVkkkza3CMdsMnnam6r5urFixyxbY25xQPbRi5Y56fy8VnUUoot
gBirkIY8lr7XErYn46ufNC40hvVGFAI0Qg2ZxayXl8qMeksH0aT9TpuLOHQyJedaWtu8ukPB/Yzn
DSoWZTnyvCg1awso8j+EkuSoYuBoCUUVU5oRhNCtiCrul6opzhwd
`protect end_protected
