-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CJ17PV+jJK/Lu+DuF5fCHmMhbSPZmhw/t+RA90rz3VirFCnb3l+c/clzl8DnWl6ua6pRH7dYC79m
m6nXkWtbe9/ph6ljEt2doWF86hKEQfbtHwSg+pwSxkt8lVVaP49Ps4HgGYk9cg86dREONV3ZWfCG
wAY+0IFZql8xmk24sR0leosRQbimrxJGgvwnLDUO2TRUmAs+PqMgcWfenBK+/2RRcp7qCDwtumpZ
5+02XjBBc6DdSQLlgvnJqi5i8GovkAlUUxS+WLiz/jz4tUqhz9deZ8RmKuX9dB3XfM/kLRiJsy9v
o9KwgtPS0uk0NNEYhWGqERiruKeiYUKFpmQt7Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
Byh/WFfABgUqb0XoHQ/YsT3zxpbcQbhWASxm73TYK3tYwIelR+PU+gxZEwMHHULxYXW+STid70oj
9zjHCYYtJp2uePe+7f6Brs0uPchSf7WFbhzHgPqphcHAFQiq1pd9rle64BeE2gCUJbtrcduIletY
vp3Fc4bcSUqMe06Ci0noPyLPaqiftirFTYoOvEvoLf+Ymc28ohFfhU6NyvzFm2cqDFZLDKGvA5S2
tBhYlMHKBpkmt0T/onpDnXHeJAm+JnX2fl0M5/alBJGOGPGQ88Zp3usKYzJxczCJZKPopejDjmrP
I1wmkai0CjqkL+SD8kd9tZocp/yNf44lRHVdv4rjoEe9PDY6/PbB5jS57EesjZsKEqxRETkLLCYY
SRBt5JhTMz9frbMyh+GAMEi5NKIW96ERjYZWYAIQUPe7PMD+Mxa0PNYIdCe8C6Ix5H1PXT1BF8Yz
egf7Yq0dp5yOFq47ryyGRxS9nIScbZl0vdIFHgHjsRmvjL3B7SR5NFhOG0Du0MAHHnK0h9s7bmY3
2a1u/0LL67ArqkYf5J1/EnS43q7l0t2to1T66RY04ZBV4u0LCjvY6VT+WrLFYFgxb39AKbY213bx
r0kgGzz3aII/idU2Mz9T4HZiZgw4kL7ZbQafOkpNqTTFfF6CfwhZSTfp3npw0A2OMYXruF00TCEu
gCgRhvfXgdOSrs51dczG1DwxWCc+wtDeJnLxFkgGJpDEeH34FJE1FY69SOlccOoEC5Mg/oFvZnky
BcYEr/+NBCMpnHCBTvOU5FloSPuvJ+je+SKVvPn1Sq51g3S7yI18CPG/rejeqzroOoGPns5r8O+/
D+lLJB8obUhp5Mlr9eIL0k+JHLaFxjVok/qkzsfSQhZIkUo2kTBIzYkytypk7poNxdg/hCXEOfx6
irV4oqZ7wXJszb4kx+r5YpsjHHsbf/BNANmDLv41UsZwTXLkcb1WF98oaxizJX32hJC1TkZ9rbHF
QiKczU2Ibw4X/X+uFQi8q59MvHI9Ya/iRlbDIcnY3aZ3lopz/6E/Nbtt/lWd4RqH74st9xtyP8hp
LLrF1AnaFCbzWWImt+wTxOboQiRn5NMGDebkWjSgcHw+qbWnF1b51IIbvpWVBiywqX35qszwbrfa
ahNF3SfRHVFS6oFvYDUCYrPklOseiI2F8zT1CeHGXTIIIi8NqoDTm31Q0b5Lv814H8MTPHy17y1A
wFBddEi3FSL9Y37ZWi0RGQoVcV3wvT3Dv06ZQ/0zprwLQ35UwJREk99j52RZMLkZDirTNtRjqswW
ufOtL4ICGOW9+aTlLuZhXanYxhF7LQZNQyNfjhaCcQO3xD79/2PzaDxWTTqhwVfIL237UgT3oacp
zYIao8XFZqHMw3KmfQ/MM5EesTm2sfkP0VJ2dls6R8f1/Yqv23qitERoPTSRudTBJoYbZaGK/VKa
X0ZkSSXr8FEGzzURhkVGOn2pOII2DMSIDhrNS3cO6OT7I9t71gjsoVlZ4EFX7eWEqrscSGt3aliB
igWF21ZNFE03BrD8xt5tdqp2PrQvUOf1m14k3C2DKFel02MzUAYNgp+8OZrmr8jXs4xuCyPmjOfd
cNF0V7NY+Bz3+lOLh5OVlLKTi2VfpCGFrGpD1qWMCmc/6iZTM+E5MjoPfUvpX+pj55YdgfROKHD6
mkFWeybj0Mn0B2CN44FY0ARB1TihqAWPrXuu4uvmFFDe9n2AZZHwdqbrFBhIYWxQbcK+1ZR3lgU2
94akXmTj9PYnixMTW2BLOTs2F565wBo0BNaPA3hUMGHeh8utz/LF2gxQa2VIkoHX7cocUpwldOcj
dTpnX7N47QPbXQwMKX1gM0aU4khzoO+Tie3unw18pfTcaj+gpVDldDUFnuJq6OUNmJJVNNWwiHSR
XN+yGNtQWXqs1NrUB27WM4uKTNFzXq7QI46WHnvcowu06mi74l765urHD8x0sFw2skyoSoinfBdM
qawKaTS3IQXrFjaIlD4GuAQhRgngndRsGGXe1Tf7mE75LHT6mgovjBbB31SYLWEAV31DEFulEwiE
2xvzqr/F6q0bOaim7v306tS6F95dMJ1F/a07IgdPvIQTrJl3iHuP3Eo7brsNvYlzNnrdrZtC+BCs
QoejkmuQ75VlpeHe7XfRf210+hfRJs3tQVrhl0jgIN3Pso4TdRIUlNLQvIPxzlqZbGE+XDzCYt2X
a6tqqMtjU0bJfq+TTC1EQgOdbE8CnIK57txeXVSPHZ/deak9Gnjiy26ge2kLaklKORcGTy3zO3ub
EQ5fa3kJ53pDZhRBpRvknh7En4O+6BMd9Zbw9q+WaVEcYc/iptI7LOLs3EoFEK7vR6S2BhAOl8AT
clHQgsIQy98k+yuIPzTwQUOy5CiXU1I3sp7VqSmQ2FrG4JwzaMwhjzCv6gmfYeIgwM+s/RpIzYgK
mz1187Boydn3/mpiatD4CIxQoH9tHoA7b2q1vGmIujyfFO2XROp4chLj7VFthROPSpU00oQajG2Y
tP/gOpXXdJajFdtATp9OhQzOLsk40hPSB2+BsM6Z0caS2KvbX1I2tgO3cuFvvhPQ/rTDOyJk0RgU
bcmCMzNJhKQi/g4NhEfY7hb+unRRT3th/v169mZ7F7I7stT32WOYQlgjz4eyYa4nIXe9zQjBA68U
8JyExTOiAffVQTC7O+JIjR+Qj7bL2xTGXpoICi0TpOugq0Fp1SYv8bm0kDZJLFrtIlCXABh/p7QE
xAoOhkipB+DOoFSYfG/3KNXvW8h7+bEpLqgOYQqqcOjuOcayDVcR3DjZoqm7gksJYBXlC6uXqsmn
LQpTqnSn/0GCdFQ+j+DvRkTcCQdQevQETNojUyVMptu/7Es0hqGdlZEOnSHd8z/a339biphDEoTe
2q/ymvJLpFAd8LLSUDMEox+HQ6pouiDg7VxOflo4ea0taWoU9nLv2XoM7f2idFdDn3SsQtUSNyGH
uOZkUTwVAEu/VNos5qpS3w4GeWNxT+1LZ3XG8w33sLjhk5pytuHytHLarlfPfTn1QyHHPh5SFle9
yGdx0RjK2gANGMActTDet845aqb1zcEEbjCFLqxPfyRI6HTtQzC+dpHjB7jCGJFEne7inl0cQak4
f7VGY9k4mhX9a0mLG0VN5Yg3Ph0YLe3eFT82OsAWOs379d/n+YARD0LipMc0847g3zeSCDu0jQjw
gFN6zJTGbN5gsooQdouaFKhuedBPujTJartgT+sMhg+K6YcDdXHcC2QQdoo1XLtFv9Q7Gi+woexZ
nSwcD43wb5Q40rXUICUV8wgjhQ5RlrIjtURh1q0V1y7vUeuEOrqgYXrcICC3ZyCn0EQC9ybf4aRX
+tDZMW7pmpDbLadlyBejZzntA9ZWc3WDLelmtCdYcA69Wn9vUaXhVfm6gNk4PRVYh5Dh6jvpDLWD
G9ytVR+q6R8Bw/l65GsHjGC/5Zn9qA4x4VHVLfv+C7cCf/XbNTUr9U2hZCPAM5t25dvOIeJ/+zfi
EHtp5no5OC79HYhPRqx4ie0Q6Z8z9CMePyfq0oeL7IfxMnRAfDko8gv5qtdjjLtLblqX4E/KyJAJ
f5n+EBupALn50rBsmV9qCNesEN53A//5Q9ib/2M6oESG5pbeJu76sYxSTzxfhLkZFFT3myJ52tZy
+Bo+/I4G42N2T8Us/s/JAn9TW+VRGnFm6UCiXaJOdznhsTOhpbYYsNjnbBvQPQPAeGcT2rs5pbK7
aSUNTpEORMft03zlwxLMy4V5+LkjgPTZHypN+BO8h2m6K6sROcd897qK9Cecnbnb68AAqa4DBaO6
VHPdHRBhaUvXOAk2r+6GZmk2Jz//3UWC5QcBOWhULQ+UMbBAsQ06t1grm+t1mw9t57zqGNTayvVj
lny5qXhY5HzbURPu473H9uDdXE+0T9FkOw5m4DJV9Aa+bevhbKk9lAgk4zM528z5Sy+FZkZJ21jm
8BGvUZg99pmu1nL9ykWjcvfcl9R9TbJSYD3P7sJq+VENyQe1SoAc4etSM3TDn8smdVwuTgN8sS2r
2xF6mePbRCPH68FSZv//TtPLl3V9X8FIOSfj7Fu9In08TxKQ40fTHOhms9e2grr5B3E/rdi8BVff
NRwvkLDrFtPGWTf+AeoeyxCOPkqv5Ii5A2Bytx3PF8hTxZiyRgAd8EMI95AQ1XrLcaBlCN0Bl+11
eE9GTgiJ6vFOaTTlDeT8GDApPSrPyZUdtAoBxxxjbRaNUCfgxrirTg2VszZAeF/ooUsxjLCCCb1f
t3X4ekxhIM+ihRYJ4xE/VpIdWET66elqW9hHYZrdXtI+uSu5WjZOKu1nHL4dIvk0J/B+gk5jGccn
CV5OMujOnKpYBCcBo9xwt0AI8tcgi1zToSDrKSn+w10pe/H7l9GdPDxEdTw5YgBIVLu1/xwqm3Qb
sWLJufCvL4xtzPqWbGcdS6COP6W8VsBIpJ3LPNR5iXh1yDSIunb2xKuQoK2K4cqs6Hs8Yomcooyv
Zrea1GrWcn1CVGtUJaGr4c91XRs8qg/nYaLvWFQFCmw0A/wreBjokCUwUcSiHDo2ZDjW2el09Pbq
feKAtemF5RUlOt1wo3dV4DTAmIlYEPD13UfJ3Iz/z0fRlFSCPlWwCIztrNhWixKkHkjUPx+q6K9S
L9ZPQgBrTRINQ6WIPfXW8cvgYtNvSPfzwzxi6t82qbFalRSqjAFcWD8uuaglf4JjfCUEg+JuWvba
GN9jRaq3xKVbB9c+FyDYjT3L92E0xzCR/WnvN5huPgYv1/c0f+qiK+Cizf0y01mFSWwKWUSlqfHk
84EkNUF/UQOMRRJ7KczEB1kVhlKqs6sfzRs+4b+gq1kMxEx22kv3DkghNodqh2uZt+JDjEBJuEPP
yRJ7xP2dFe5QyXuIxTNK9UpvnQ5om2KujjGDyTnIy1cV17chP+5nn2m88nFeAWkT53tyxUGZo8Am
iS/KSBJJ5ixRYl1aHM3YO4LraJhj5i/VvzgsBp5GnaH65yLOicuqJRoGyKxjkNZ+AM/HfQefobk5
/Mar6GiGJrcTDw2nUl6vpVz3vTRw0KIWGhMhHaPeI/a9KIBxWygyxD/+l3jtYEb7MvsJ2spqgwdQ
AiN5iOBOLRNt4zPXACunBiRR/7zTayFfNMKKvNOId/UR0U0GMSzN7AEtg11wv/rZoZk2TmbtMUMD
XbPrq9bndL9prXTCcgiFgUOhW25weDYMO8lD3xaRijAtuFId10nOpqZp1SyPJt82Izwzpgi9Oy0x
K/TMEIHNL+tsIMt8RMCQXF71QcRCro/658SQu4EPWJgV19/LOxEet/99hw9d1F3g4l+X/YBcJPLS
UeysuXbRwmnYzmLdgWUzHE8CiTkssrXNY/ZJG84vKBUx4Uu7vKI76g8+ahTt0USUD+e2+wg7URd4
EnZ6Z648R3BBioA9T3GfhtdwOCD25miCiFQAK9p2t1EzcBFuFj3o0VhIhJdwSY/OtTgxCK+RqLmh
Si/SipwXdZEN3O6NoWxgURFRuuVo+MMKZW5GCsRcJr4Swj2kSEs5Om8G4OzbSi64cCsanQBjfX2U
DDO3HYgPXaeU1NaZP9lzWBlgSWDxbOE+fVpb/0aEYVtpdFN5tK39Rvdx3w2Hx2lWT+impHxIjWKI
JD65p3NPKgV976JmYmsIZA5FOzqEJiIrJXQwObiyj9D00gv5vovntRxsE3j2t/WuwXzIbU2ue2eD
Hn1Np/+kse8+3fGLPM8VY/Csmaq3Y7bMLvAVH3/Uxiofm+l0V9RGXOdaYxlxLIlSAJL/jRsk/u6h
qurRojJ3znICKA7oVu9JmGCjKShEQtTXy6OLCsDON1L3+QAE3vrUqoqiUZ3RjF3YZ4cXAGy2dxN9
zssuYDvoH60Fg/T0QghkAn28OZg1sC4SYp9m3/YIRgtxXeCOZXHjcNzyz9lh0FE4kg7K/lB9NAUD
0vSinq6e9Pbau7Z3KFEN7mgMFOP3P1eLBqPl2f5daPOwEzW7q6psi5IpKtlIr/ySZ7iGEox6OI+S
2I3D3kcGLIIrPylgWaYtsDpjKFmJaEagxOjP02dxN3D4KFxAPOHBZDZH8pKH1Uj2p7zytBLlNRnq
UTKT0UCeToGeL9kj0mHo8z3KOJvediCsnA2fDHMLIQlR+INlcIkqGDuqXospRpR31EQ4gSnYj1zD
9J0R1TT27TXokh9o6ZYPpXdQHanA+XglAICRkiIV8FZbT83Q8cBx1mkDex/hRdeoQuZPXWpjsQ==
`protect end_protected
