��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i@�n��#h��p,ƮJ�b������8���e��ʼ�6cy M�gP��g�,��4�p��䑐ISw�cLE��k�se6lĈT|�,�[c,,�e���s�M��B1���.&�U��>�k4ϩ��*o4�+�ѤG�3@��;�����6���|��G3"M5`C(�N��o��>�s�.�7�3p�D5Jy��5�
��%~e	���Z`��U���Eѿ�Ι
FQR�ix�8�s��z��Ѐǆkb����I��W�3�������u:�|����F���_�Et��A_(f�h��(8�R�V+Lʤ@O��T'�`�-04FU3�a���y����Mx/>�ߗ�pD eN��1t�$?�r��n����En6�������z�G�n�юd�����6f�h�Zk��Lާ�r:����J�.��܈���F�r�,*H.�R;ݱ�A��I3��5����F���<f��s�>"ϑ�_ĭ_�����r=I$8�E88�=Sl��D	�^�\����u�7��j4(2TΠ�2#d�l�?�M�=�.Uރ8�ӊ�/1���i����������i�R]���u_��L2�i�~����#	���ϳL�N��6ZP��`�U��&ڣңL�x�	$�zE&�����e�M��A��G`��4�,�g�v��s[g�[.p���@��6��f5~9,	t�9�ż��&Չ_{�&p���b��I����Jy��zݫ����-�S�5�as� ��J� |����G������w�el�y�m��G̈}t�o��I�×fg=��}�?���@���d{Ez9�/��v�h1�)�"�Ϩ�HWb�[���ӗ��h�Ξ�AP�-�]j��k?�