-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vVZFfzBFrvclt7TfhnwW4WcDQrpZXD1i7hLGmlPt5vYyYkeXAzZFV57WrUhyS3KmJMfTnXigJEP1
BvTYaRBqF6a0yX1+KBAxoB0dVbOO1bf2yigIADMnJhyf3ZhooR2tAvuPnVExk3p70AqGwgSpd8Sz
qYjlJ+rOCkvupkL0jejEPCVmtjcJI58lI4eOljWP3Lt0lo+Hh1wYIOm9tzcoQevC20IEClNHqjKi
PvR3cKzXxwz3wJiyvgMR0Vlroxv4Grg+/AViVhqVMMedBqs2pvu82iJZSgjNZpw0Zzo8MmJ2JI+E
qqkkM97/SzNAevw16csPTBf226rVvstBLRB5ZA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8352)
`protect data_block
6O3UTpZYx8dhndU+XzSakDIfTYgzHHl0/Q2zLFqMXxfDXqY8cpW5rbPIQWQ2V9UWKj5+pC0/NQ5/
GD+9AzMOmU2O3NGl5XHrdKZPwoWWp8wqvT8ZSpU+w3LCF8GsIdxmFXVh+3ADqg/a883OV69Bigem
Ko8xIOi9ZBYAQJFL82zY+8B2u6N4MPGnO1KO3w6yWJAFWbxgKz3PAnLwc6XFISMX7FAaLnbve0b2
lZBAqQ7cY3rwyZpi3/3DthFlVHFksdeHJN0WHRkxr/XlewQmiJFxQST4SlWCCbBtnQrFJdQQVmFU
YnimapPgB83geva3/jWhFjdzCWB6kxpIRjRk3cwE001IHK1mXR8kWzK6HMPj/JiV8R5cZ+IHKGe/
/KiaOGUow8Ebaonrk4mxHLCrvAgZllWmsaW1WIIItZuFFxRUJVp41a8fZsajuwInKfjr0Dy7RKlA
ts5fAR0NECiM/1z4+cwXj/3RWBwQuQmcfBBKYGleEdd2ukgI+BD7uqcB3YJC+xpb3S5Uf22PIvxk
iilp+25EB5H7DVNSCX3WsZucyYWfVbV0ana/2SuhZvgOnuoOAaWXy5XeHkANk+0w+42hmtElFRNI
iQSZNNTrhYD7LsCpdalzwkjCTw3vZIBlxTQNX81YI9fV73IXj0Nsl1mmwkYGZJGNfaGct0DdbDkJ
zT2ebpVgHmCS1UWeaEI9ybbI3KL/BJD9HpCS+hu+MwKPYvFVSgHpRiK3Q+KuwZrxJnggFjOqSstD
AstQJGh80FEbkSxp170VniU50vBRlynm2GaBctrOfGjX7Tt3sb4vFa6l43wddWpETPq+QfPoYaoH
W1zmfeq5ehXD818qIjZSjheEK91tALsnmFmc3fZo5YL3/tWlDSm8Dz8tqJP7JI8N8jemkAT2g8K5
MSad8KWmU5Mof/sKM5NG15npPr3NnIIxRb8ZsSw+cPh4Tic2oNgsp4wHb7USCV+EVTszvmLcdv4I
w70m173FMmFDjlG6ZFWC79d98/9nlh8dG9ynmz3qeXYVwVQzS4WyzX3gYmEUz5WldvMAJwo92Xxp
C6JJsmnZRZkwADIui6G5hLVCI66odq4X3RcM+dCCtNCW+hBbJfi3pwdbAGi6ggg/VQswWGdPVx12
brU0SatGdmWM3kolwMvEKUBvfwYrOF5W16OsB0pKy0qxucnWEoK4FSzUQhCD/LKVFKEhalyu/vMn
CZCaqZ8vIvwAAviPuo7PnToZwXHsusqwRrR3fBTNQAt8/qM8asr1jrre3m5iFH2AZZtJTHJOEc3Y
ulE+P8yJhjOVS22jPZeTREx/zMrF8T66E+9Sm1ije0EdPWOCzF99UkZqXROZs4VeJwuFYDCghBep
J+WRVN24+KN4vpw+/xwyKA/cl78UHaKZHSEgMjpDeLBXJhXt18/uhPSiU0bG4Ysmcb7bwfl3tyEh
1cci1jqcmr4uzhiCV1TmrVuXAMVFCAr5E9KeMQ8ixwgPcKhjxS0VzjXPttuDx0eaZRml2/eTGB8i
8LGkKzuPCO3Iwvh2BApZvw2fLU1H9NYl16KfaOfUpRhjB3mwiCJEgPBragQ400i1HJW9VF8JetWX
FxRLZixWNrEmaG+sixoRe0loy+FXjm71Z5H08wtotpflC57q/KXxoT8c16YJAtih8FLFMYb343D2
opmHdGxShp2o6Ef2cicFNwBVsXfbkbrChWljOCqPSibG0xr7bNKHMr+9PbWnPiimjy4Hr3WWBXlx
BVHcgbuMIy72Cj5FtI6aFiU0istEf5iAbP3BHR+zfP3w3ILCe0115xSYeZZy8tsdUzctXJUZK6xz
fki+w6YJpdfPpVdIlxCpOn319lw4MMeFAibC78nOzVRYAVoVCLV+8Nc74iHspNk9+ktAB7WPJJ9D
0k8DHliRO8yk8dhiGkGq2tGM9UOVwuJBkXXydDEKsn74Av9KTrpF8RwLr2QP66rUl8YGe6qEr04M
NPWbLrM/nv1rw+CjnDdxiZ1/myudfN+0n1WoaNLOQGjbHQds/MOQlosMMAy436ZXy2Y7XIYY1IF0
K93MZdZJC0CpSyIxE7TnNPJO/TS3mYLH70Jtg4WhgICA8iSaMSgHks3kaSedMuJC20UtUiFdagLG
yjDkjSDaeNbBMFMfxavT96ERYMYxt8qIkASqQBZgNYOya107jToiEZ56VQTWtN/QviBSGEiySVut
854bdHmsCEboFad6hfbILkvHR2okcE0fATwjOySsb2JRBdvg5+6umxOghzPVtl1hXmUf+OcsiU12
0SHQPMMH3hhfVO0aaGritE3Ry8ynX0XZ3cUpqIZfEKsfxBoOtkgqrObEEwDKS/wpCGyG6nRgfVVd
rWN9R5N9Z3earjvZIjUmCCzXkV/xEJO5EjEIAgWnGYrVx1YxpUK9xS1hRN5IlEp8NJSt/JiUSx9t
ixLHrmFIT4blaouZESURHKdiGbvwO0EKG8ceeDs8c35MapsiIAT68Zp9Z2QEwJg9lW5QOExh///X
MAFvMaS6ZE9VVv4pY0xHQMwEpaZ0e3EKZN80AnOL4dGUtIljqo2rpcahCLOgOzVO6KjGWFkYigER
itYZNcrH1fNHCWGYocqP2e7RYef0MDIIoewAgQkk5M4nRoeq0dXVt06S2I/S99zrMzZ0BQCH1NtF
3JomWLNdYqRdNbQRWpJltEBLM+Ke5msYIKLYN+pLOD9l9277aQVU+49rJ1tYtbO/4vbUP2hhiufM
ZQEQ+xss47vsQl3MT97d0VziVzOI5vo1petR2ZbqDfKF33QLNMFx7oCrV7aj9A6NDPpirAiaAv19
aLTt/xTh9ToHrGAkzOgZpbQdFcCwGClK2WvEdas+DPoJZZ7ZF8dqJ70DQyQZyqLGut5lmBK+/bUc
GXmS7n8f9beYVlriirjGX1NclPONkKpbOc/Y8TMA6lUYT7L+Zc4OrZdVMOttwbOxqcvt9QlmXTla
I6KCjRUjsJaKkBBr74UsdoXCaDAtK6kOQbJa5tkqmb+A7AdzoEaU8ZncBB6yjBZ16blmlLCOFyDb
3XkyxGEtmKjTGHyp8ga2MpWIk4JEkD5m3mA7jlirrukTPC6vJaZ8T0QfVDrPv6g6mRQt68RSgwHM
733kn2g4TLuTJ8YruB6oJrR69ppivZfqWdvBm7Gzj2BX0vsBDXNEMnG5TdA3rSlHZrNqbk2Fq3+c
EKsm6juJqQ/8kWCLifQ5ep7PBRXpE52fhiC7Eev2qCBmb6IFbvALNf8Bmpxd/x3NEMPwaxWbgDoY
pK9jNsFnMvmmh75qGNel3WKLlLQvSEflGMpVOiPBDv2MaREjB5sk08dytarl/91lds7CGACyMkG+
hNyNgnKHYrQeF2RCEnneTiuIvNimN7KJqcBReeIX/1jT0EYp5DWlYpNVPZBHN2rl7dxt80cVKfCF
Jq52hwk6GNBvg2jy4JAULm2yjxDKQxQCdzxfYX73FOZq+aVtNjN5Uqn2uQVk9ELI97CHrcnJVE/N
5jCFUOaS1PGOGxs0YZKogFhazKOQ46CXQqQ9Zawm9G4kDUNLAO0glD+soIPXte3AySksAb1Kf63G
Dh/4V3bKtmxyQJu5oFBdUUVh7DS9wmYMoktZjLCDxNf+/RXOgARq2IzXpL/K/ppFnngSEAg6lbYh
BTSY7XjGyBAxllrBUVV0RkX1DXgStNYP+OvkPwGNI9sn4yLuEGpeEgBADyyhlOIbYrAJM4zmjuXL
hfr7oKphZ8maBpf1UeIyTnFfSswMmTVLbGUVATNAK5EcHb5B0cR4+NkP56K55X4IZSmmOTvqWcC/
qvsC0mZsrBG0KCG8+iUNxXjTTaN4jAsmswVaVVLZsRLpJbcqpoKC33A7Fy32pOFNSertjTweSG3s
ebfMnm0hBhc8ZFMWCShpb7sEXSj5OZ4BF84mK8RLg45iyq7aLzv9lNZ5JZXG/5QfsxP9WGX2VlWV
UqGo8582plojzjcEx4hyxygPgIaEeHO14+dlM6KLkDfRiGTcNCP1p9EL3VELZgur1W/bFulWuSqQ
cLLaRNIspDEtkcKHns/X8c1WXYh+Ofl97yq7xAIVyxWdrGt+wffvEFqbaxbAYYpQaBOsGlto9eRc
gSyfzh3iaNjFf3EGDfdoF1YMAMYG5dA1ct6XH92fgDgyNwZY2kajODsooZikAuvrPPD6H6LYPkUD
zC3vRQfkMpJ4EdzugI6V8gDp8fIW0ZWMoIZ2giv7mMzFCXKtcM+Y5PrG284iynYe/2zPs4Fhz+s2
t5dk3gr6P+p/FP58m/132lNQYK8cMcNl/fgUl2243tJxWblMQW9k19tln91GoWBMhokq55bWq14s
IXg+3Ym1/qgVAjdedBGOQMtS6HFp0UlV4oJJSQz61ljjDJIPWMFY4iGShaHL3k3zq2HfurEG0F9q
0YGqaDbPApKaOnP702vnGA7QtHiPUiKUVYgDFPmVq8wXV/tj9exevSU4n4/d6DJnUkKe9mTSCrxE
14cdcnFdtM/vw1O7y99Kk+l7yPvsKyYr5Cms5zpUkcEAQDG2PmRRwDEdDhNtcyBGMlQThV+NSSDw
vB1u24oden2yx31QRFQq2bYxktX/Atv1RgMXQ36SPY4Bp0JO+IY4n9d0VP0pkZYdoFe7E78mFKVV
YyceRaImm5ie6Y7gunfAx3KA8v+xBauX9LtmLNvGi8FQ5SqjnbsGwp3OX5hlc6wssi+WNmpfYMqU
NKpSYgEIoq5rmTLGqG5vr1emHhe0PrnQRq94LDdwTDc1kny695/gjiUwl70aXrjWfG2p2g/LQVOc
eK5JB4bbQIj56rQcKzngv6V786bSVINha9vKttFfn/9qoKRYSfRfe1zzz/SdoQctIR4lRWL9eBfC
dGuer5BzgmwJdYMXZ3VFHtR0/qWN9bZ3Lj4u7bZjCYT2ZXlvFTQehXL4wy3cug3yhBYq+9JVLLZs
yrM3pQ69bEjGU6VAaDOXTU6/5zEMVFBfNpZcHp5v2YExQH2e8oCW2jd4AnNi6D4uD+mimZBsxqaM
zTHtKm5kDn6LRxwm9qjHJ/P5jlevD/K0DdrehgJuS9tR/g/mCou3+P52Lds+lfArJkH6YzKQCT2r
LSaodvPJAC2f+gEnbuMMz7RLFCnNRmkcQudnqDA7fBRXBFwj1ww+JQK1FtXltYX3icE/UDRIwRXs
+NKJYxLmHouYm0kahz6kZYgbR14ec/6+acFD4FYFSpFpKfXklkLMzjzFA+D1T7UNNTKzO2sBD4vD
6aM7A+SLzqzPbF05BJq8g7Kjj+bYIKqrJgdwxaXIMQqFgzOThWQ1NzVzUTpQNXIJoIZdgE+jBfrT
t9gtcEJYwaysfJxHr1ad9/O1D6zZZWiELpiRAzKNqKVPi44APCR/p1mO5xhNUa+Kv8KnRto7zLv5
L3KsmHhD8SMyE/X/GLhw6WEg+a07AGBITjXcNK3dcAnYyMKSB106DiKMwLBBbgn6jKWFsudEZb3M
5KTY4LjoF8rjudHs49YHL7r4BYOJMck/CH+cznsDmvWTGYbDRP05frV8HgwfQPKHtMNynfpj8SZM
kWRFBr2ii3cjebC3MLoCgFI6DQQ0OIri8meeluF6wDNkTK3YhdK+ucwYzc22sMwVXkUQlzl2Lrv4
CSfJilyi8H4ENn5v9WYGDBPFTfGtzvhp8hRASOncXdQxNTDcWpXEgKeMSlPEbAALIK36tZmP2mmz
v03f3VL0+ZUCwzWRMQveExTYgOmRLdZsOwvekQfMEgWS36pEeE5hnmd01MBfxAViMvIkXJdoPP+u
Ovs0+kTPF8t/STQ0bfgPvYJMS++QCwlMHGcZPZPDHjI7dUcwTrsw4Q62JYbFzT6R6zsRmnLnmRhk
wTz/6r370k077B3M2k4PWNPvBKRuxMgiT9y45RJovi1oRAfa0XgTf+JdjtcMWRjyq4tVRy4h4Yie
jeblpumpIV8evnR6Gwd4JNwzjmpO66TyfOIjt5sw2cQzfYs6iGGdjSXxfwt4cY+m3xSyHPJZ9nHK
IMcP9blBLHNpccAV2W1ufJB9g5WlDoTg1QTGa9JWdGgzUG1tqmqiI94qVbjHv13CjIFdbMsVEPKn
FZyK0e+YnxWVd0s+5Z6gnuNC1KnctJ4ppKVl+HRxaDBG3Q0b9pnwe89RBs7/UH3or/vWBpoJ+Xzs
CShEfcZkmIl6y5PhJc9HLt7waH3jCLors42Fc1mGwMB6W+E0WFCBLqUCviSXkMwqXYZiskgNnpFK
PWxbXfaAtThKNIBSaf+oihJf1FC7lJpLzuqSNHiAxjFsBuYe9rDo1vjSm9JCPkKLiByvDEj1EHUd
FAlCQ7Y2dENvHZBhffmmgfkodM/Q5d5kp4b8jAc4vAikEkuwoxJ87DrJ8/ZMiQrsoi36nGqZ4h6n
IKoCRB0KnAZZZ5kMW+sdxEbG4asBkaxRsLAlxtr5UeSZRbardax3vsZNvbTLGb2Hqw9Cgo798Re8
30ORu5Yn/7TWpy9Vv8/j5SBsDOPO/MTW4JkxylYS3dT/rw2LB9GSqSLVyHjsK1knfw+i0UB61ZSB
zwkloRRQ6jeTJ7rTu8O7aK2X3FPZU343qCd+x8i0gyotA4fZG315MiebilNBO+iLrAWV3NQ0KLCs
ZUstcN1KerecG4qPo3aeFjvVF+8dVaxus3rIAempf5mkv8jhr7rF3A9j9BNuuQgky9Atrgrx5QJQ
8DvEXBb3bEE3GDucydyLHBZ96h0fR8S4z3ML1i5QQk3oBBw9ISziQKyk3jPvpMSTg0UtxvNhfHtc
i0PGPvmord1rQKYQBfWxtODyUrXiX/BkANsuVJRavS2a1rkKrU++NVv1RgCUNDK0OqUce784PVym
1omwNPyNjK2QQwmCx/nbj/O4xcDl0Kgq+4ybDar6Z66PbWd3lfCKkvmpKDpSVEwD9C97gz4fWlhO
Xh82i6wkUfftn4jpPhWWPg3L03oONU6cSS13HjxtU6bUnw44OQHFjSl4am8f3Qb28YQKmNrFB0Cj
AJJeQEB0qUFV7qVFXJnW1KcQvZVObSycCxMwyAXDiJiVXWdxaFmPFp8Hw5qZ8TCyeKaORw0Fe1lJ
FS8AwIOER5TlPC7jjoTPIZaIh7KCUOoerjIZ3rxj28DoJ9pnwQ3cdrUcSgVeX9LFKPvwJu9mKn3d
V0QTiZc20CFtHbyO5vT+W/fLc/ac5X6zI3wgKpv/zgBHPPdvmB+apHZ3jYFB8naHBFSmFjWA71zN
LstlaeeyXBgW7LJHHdY/31QhVo5udiSzUPKJ0oKi1pdTPwWYrblud5ENCqdl2lfcrZtbTgzyiVFp
iWJWYQVvUbc0HixG2QdkluL5YB5MZ6UT8o2oy0j4FclQsQ+JnP7cNP0zR3ffb4v02b1agiEyREZM
XFxr1aUKdnFVwXnnVbwXJOm9B+5BGD5tEgTkjIuH6xj516tmSpQfkwac1AitlQJ5zQ5NjUmL3t2S
yuBHmg3tJfMmZd2jWqxXlZtwEYTRu5QbZpnsIzYy98BKT05SgbLDu7BeDHUKV+5CJOl79a8iYzVL
ejA4g9xOZhROwBmIhwLw9VSiyE8q92lX8NX3ASXnNAvZfBAJcp2jfV8RTM66KFBG433qb31kl1bP
SZcN9dNrG1aPOsKCD/ciVocnfCuz623Gbgqs9tqYjFEnRs18CFZ/tCEcPSOVuTwR+KEkRHrMbuh4
Qz0HgM946GxZcpdz3YWSCUpCC4V6PAIllRe8ByDY13H74vFc5u6lD7pVwLVW+8PTVpIZTwK+4LWh
Hkb4qc4DEXaoecIndA5HwckJzyoy6JW+Cn1nVRXcy6aWaJWfRdCSgrDOBvJlEZCvgcO89eElVjD3
k6BVPBuaPizBKCIcJe8frESQdk/e9+AVWQDxDo+9ilViYhfWg7D+UeKZNYClZc0/30YnW0KIGxKI
zU9cMQlJHz1JOqMTnN/5CxXl2NRgBNtuNlpsex44V+k4Ho2VP/Nk1ohQj7z1JAlJN3v2h6aBCDi3
aF6AUAWXvgI+Z1HFJ9mn5c99ENBJIdZEivqVmojSHyZzkkRpOe0P7g60kcXUXCbxnJePGEG+OzMp
GaCgtg+k5SiwAPL4Dz10qAJl02/w3YiXP0Kc4LBzUgVRKcwGvOuHvAlo3zjUjfeXmHH2SRxuN5fq
mEU8Z3edVzdpM1YxveUmIOCyuhd2owwImU+hhKIYylPG3QHD3uEQaHLPoUyF0nbrgjGoK7RkFgPp
zgvpZTNqiDu/VvQEwOSjiheXygDuVHW4FleNJxyY/DdRhrHb9w79netZZXrUhRDCxkNjJXgjIhI3
d8GoWlYRQP8bYfqCbOQjgR8WdhRov5JE8gC2PwOKY2W42jEbhOYwWmL/osk17JawEIvzKpv+SuMr
Rtq29JtNjWWtO9txpA6/igg7I7w251Zp6gClIoHgp+gka/7wUV8shdEl9OoXV8hs4XLxLo2Uczph
6VPG+oi+O3Qgw2fgckNUan9+wwTYBZ8ejPM1CpkMUaJcv9YvUkchZiSG1PoqpvaYEQOFifdM4S12
rKJyCRoJW+aFJTgknYOX+FKrata15tlTZT5goAY+J4rGJuIYU4DIKC9T66V+SXD2kuzi1TQQOdIg
4TVRFNzwNY7wxrxpLoT6p9nqWdZu1PVkG6gCtm+cqYbnX98FtAspBmhFYi/mdSYzY7bI250ihJGU
517ewl9oYHbZElAAg+sQpTcdVUUQ7FPPHPzFE64tRnNHdMDpZ0gMPn0CSyKTu8rgRfm6wbbTG8Cm
3sWUbk12odvg3n3+qM+msCcCXPe6vBPVnRl4TADeZ88qRN14r00Lht6i4CipXMSqEMODcvQ9jmU6
kMFbeHO2b8c5gITiGkhX9tTPuarFZouahPZiuDuzYFLK7HaORjzKkHa8UtfXZszVIAHQ//m6lbMQ
Gz7tXnzZd/KTbeRNJFm/tB395dEb2pkFPFjSg8/rceEyVHtuyNqF6j7E2SiWlKeoB8+Mk1ODiZAo
J2XgrK41MlWxj5RmafSLkpufcUwjBPxbjfQyRpoq2QAg1l+QEsBK6ezZp1slKFA6+Zyr0eiM6CPA
JRHOoQwEQ4hjP5D+mrG1oyiIK/kZB64pdUvlrdVj0Ok8KqSdnfRc5Fx+hXNKRLJvX5gKFA5oSwOQ
aPmPO6czkd/c7FWvHRemHCWE37qfu1ZDcS9td5kunduJjvkSdvL87ZUtRsDDPh8RkLUKsKA2KOpn
NeJfDPw4DLbBQzeR1ZgMyc91MzfRBo7oR2oQoxdFQi7Wx3x8apkQ43QQq3Nrbxm9LjSedts3tKNe
9pOmDbhtdiYWPswG6PlUDjmUKv9CNtv0vYq5F3QISuhw+A90cUem409zN4hUzyxdNuJdCBZgPMMc
21xY80TaxJlO0HBUA1+GEy7DH3N9HfSjELLTfyi4O0tp1kSW1zIS0usdIB/F6RApDxgclWCME+/y
c90Qj+V85zVT4Tt0uTJuX+MEQSbyQLBsHbZAvVT5Xx3O2pfHfT8oF/tURgH5rVnQCiogivWuwiNv
F/QpIEZCldjDfcf/m4Tc+GmUlRYjDi+4TvXgYBYWwbKrcB7V0DzPNCqgwtLOqUiPMqg/+gJKyfOX
GbKLDHZBACwviOopJdwUG+A2pjeFD9AFHoVoS9CrVRf5hnr6H78gxEvTX0eDK6aLMKwlj+VJ/Rnm
G7pAAxEqvAge/jUx9cw/KziWFrIIDObwgxFB/14yrEIe8KUY8d4KmE0k8ORVME1K4RNzyGf9hS6g
iJLFf0v9MkC+xw4NuxXDApkMruBnY5aTw5IUgPgY+pThBAQjaYS7LLtTMIcDY1hHH+l+z6ys3I30
/D3FR50KgZoOlGlFzqNS+Cw9Z66/8XZxDyt6Qu1Yz4fD22oQEFCEWnlLRV9EqW0GEwITlwo63j/+
Kn8D8XtI1nXic58tBGfPZAwxEh5T2UmgrhG4udm9Ar212xmP/id4W5LbGzHBAW+a9NTOcW/GSTon
2jZv+CJmjQRFXW8SjKStVHxLkCb8vkvQuIJjtUsYYOB50c9EB2bQg3ehX62EjtRfPrW4k/11k9LM
vgXGEKQI3lHSQcFZH03TzgWtN9xWdG9nvJ+bcSgkwe9TK8X/jIlD7gmKW9hZQYdKk/gKKqn2estF
vm7h1b/3HKIGqpbxw5Upqx7G2AMSCZTjoZXQlRBBzK6VawN5Me4Ku2U8SNsrTIcV1sWvScqLsZFP
tbABZwjpb8dhjGBR8EANbH95H+C8M2j14FlYX0PGvWMvmNlAIGYxSqr+yxdRdrrPsgcuXAkFxy3j
N8/Pr98O4XZwvmh19IQs1ctEcZ5cRu8v3zhuBlnyzzuycRvDY8MKY1neGUxAulI4Be9eCuZDFk3m
o1w+FMS7fSpLWxLqvaYvbqtTKQjlp7oDyqJnmwayqr9lw9KzlLLxtcVvhsBpTo5WzlRIaljrVlAg
BBmTxWPuyS6XT3m6FYR7dx9wWU5hOSTWO+WNps8yO/RbkJ/4v7s2xgKBa5f1FMKQ3e9/vWvysiWj
678QFnii6ba+BdRJ7TnAvwpiWoO/hwwLl6V0KbT99KKjupVSnWBT4KKPSeRuUMrwBd/WIFxZe5OY
/h2zEUNmlezfx/cI9tbPgiJ25/v8v0e//ZW4MBXIy+aqSAJh4vuwt08h9hzlOHBUous6v360hpVJ
x0NN21AQ+1ebhlDh1tSW5W5d/mrSctMxy0vrIX2pYHvmhoQ/oDTPbWIWylpQCTpY1mk74AX6zZgp
06RIfNYl2mhZbOWa4SMBMtpKFoqV69oYQWeLQiSgYOayZj1MSFA6SbRMm9RGhZyBFRnP1QGoF9c8
ONlHX2dlkBxpL2+/gdkP6z1AnFDZ9HqQUKzS9UBQbUgXUi+n3C1H4NKCE0zHGpYojc8TvMWhT6Lc
lCgMmDgzTfHAIKJjuotPlKy4rgIlsbe9lAR0VrM6JLqtrtR+D+0B0Ks86jIQTBAbk+EnLfnTNiZT
D9soh0EbJ2jw7FS4NHBVh014AoUaLP9vumvu1Klm+I6sfo+Mr8bV416HwkWUC2DwRrpOAsE44ZG4
CC1ondG16iABTBXBBfZfimd0G6P+k+EP3ImwLYWkY5TmuyXnixEs+hisHtvNhkpNY7DLLQQJ+irO
V5YCqqlWXZR82gOaTeAIQ/BL/SnRacQsI3zVOrq5
`protect end_protected
