��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�#���[(P+s�G+w6m;N����:�)�ސ4=�]�SG�|$�#s��Aa��Jh���2�ꦏ��,NS�`r6Ng�<̰�#����1f��|���Ô6?��&��{Ǽb���J`��h-����R�`j��?�R��bsI�	�M�zy�`����"X=;�d$LD��t `G�ĭ1:���Z>V��#*�oA>>	��$��6Kk쓡(���<	��Y �ӏ�h�4D�C*M�k,�T��	p9�����
�:��G:�;����n�*�o�Z]T��,m���r��P.�E� 㨗<�
������N���!��׼����1��/;�iڰ唭ɚ�˳�Ɋs���v0i�%7�7(����5u�)�����u��82�e���^��8�f�_��P�{U�3���⯞�>֭� �?�F����O�Wv6x�e�(��g�F2(�^�{q�z=<F6���t�x%��y�6
Ub�D��!�;��� �Lt
$Q�AG��$�+�,P��k=�� �0���ۉ���J3�$��0P�qc�p ��nB	��Y7�CH���xG�o�*S�*XI��� ~лUe��a�~�Ć��u�3g�~�0EEa�@��z�dH#~�ʀ'}y���ښ����I	��5���wI�sX��M�b���&�Sy^�I+�L{�h�53�)@���
�`�\�FĴZ�d�=��)�9I2�~��Q�Z(�Z�l>����B��Bz-�JU��s/׺�0�zȋ�8�`�H�G�gU�x��~e�Mx��#x�AyPb�f����#�%c��ݐ��p�Gp��c}�Uc�ݵLv3���ɹ�n���݂_�%%��u�#;��`"��ſ%���Ⱦ�YV+�s�A^�~�!	d`�� ���d����F�-k
E
��6�b�T�&��	@8@���xg�O�O޾:U�����[�m����]�"ߺls�^ DZO\�b��$�f�����6C�r�O5�N7lC�k��t	�{i���!����^�b��H'�z�>�N��؛W�I�YY�5��õ%��)����Q�Ӝ�\g/O;��/mA��DKf+�z��D��� ݬ`m�o�Ÿi�(h�6�?Y{��P�,�%�+�5�DS[a��������$~\����@��[hYb꟤�EH��+^Z�64�2�F��Oޠ?+���p�3�����&yBY5ev��K�W�]{�D8p4?���&g��c�A�z.y��ȷu��U����(��tS�����!����_,�w�q��C�K	��o���vN_n�	��3,���"k!�M{ZX��n����M��<���BS4q�'@ Tb4W��iI��i��/��p��>G&῏�Y�&}Ɲ׹Od�3x��U�?����窨L�bL=t͚�XwpcXז���P��4�{�['����X[l��D���I��b��؆Vs�����1Q��a2�����l.��F G�L�(�,6q��u_�t ��)%�����F9�d1?�]<:�h
�F��mg��Y;No�������a�=�b�PR�Z���3���T����Ov?��a�f�F�7���AɲKVNz���{�j�qY����r.p�} 聺")�T����L���L�7u�	ojkّ1�%��� �f#��ELT����=8R��Q��yx��0J�'�����r> �_R�/����:]bx�'ڎkL�Fu�Jl�H��f�pG&���刎T�[�d8Ţ����u�Iw�!P�LZ0�T=�X�;�X@������l�6�z|�$����+��~x�ra� �1�������Dl��������+^_y�E�G -��zo��Ob�����oȭa��14>vl�p�c�O��u���I�A�*�X4�4�Z�̩r�m�پ��0k������w�Tew��n�K�fD�[���Tu�� �{�z;���ě�n�����R�U�V�7��h������5�{���w�js������DC��)�s>���b��ಔ�Ƈ�>��]Z��N9��҅tL��hO�}����Rlo�<�)���H2�/;s�,��G��fڵݱ�:7&��F	z��P/J�9"�[�`�7�$��rYʲ���d�9��:����N/��gS�pH�X��Y	iRM
�/�h2d�ZB��Yx��
i�dr�#�^�uءu�Ean`5���Z�	���{ ���	�p���sAn�<�c�O���Ƿ��ಳ�GPu��^D��7v?|�.�/� �Z�9g=�0��\��ph��_���Wj�-'P֑ণ��C=Қ�ҍ��k?%2cb2�2����ay�VU����V�*v7&�M�F��U�b��gt�
-��$T[[��n��_9ιd8E�'���<�T�MU����[����~�v`԰32�7�b��tʓ0�|l�5˦�i�#C�Ȳ�����2��{u�.��FR���Y��^)8�����<����������kqGg�R���~�f��=tyd�U#���D~���0,�;|�*h�T����r(��J
ED/��>�7��B{oĎt3$�K�YK�;�p�����A��ۘ����R��diov�mlGy[ȫW>kx�%^��{F!/^�u��f����^3x����U`D{�*o��2(3��2�)���"&��-�lm��,�ң����� �'�JQg��E�rk���|�,��w��b��D';^������Z,S��~��0�C� J�wH�e��1]�1����mQ����|	s�k�����tc� 5�q�%BӠ.%lD��r��pu�_P��*!<#�<���;�9�[	%~�u{y�L��]�}�K�c-��p ���"3G_�Ѣ�����򅤈�[��zV�7h�Eu�9��U��� ����r�V���m�٭[i�x���H6[�Fm�ڢ��x>u*~��mT ���5_l3��<��~@�u��L����$�2^��2p9�+!.F,#L��"�{���Y�i��)��ߋ�L�8����l�����J���*�x�G�4#:҂ͧ��Tuj��c�N?�K_�Y�O��H�X'��u�H��e��p}���B���%��pd�T��f���/�{�W�Z����.1YT��M���iv�nu�� ʽB4���*Fr��(�xς�{�0�Sim�h r$��0�3�o�J���|���7��YsX�i�+�^Ұ�:��}H�A0����r%j��{g��>���ɻ)w�i��:��`t
+S�;���G�>wح6U)�3��2-Q�я�3 �Գ�Z��!S0�;�����sv#C���OK�rv�⬀nJv���8m��lʅ;��<~�����TNm��٘U~A�߷]�漏�?��q�ʴ�� bD#�d�6P�8��w]��pi������f��E���o��Y�v�ڼ�x�uV��ֲ���Ɣd�b���A
�$�43��	H�i� ���
2>(�+`���ǉH�e:�nU�����ެ�p��y�D� ]&�DG�e��~O!��K���� i��ZY�©�n���3��	t8�N�b�.���<6l;���Ψ����n~��#�v3F�sRh�J��޷�a�,X�X�m#`�}��FZJp��Z�A1A�t���C�Tk���h�O�'=h�[�^��cӢ�?BAn4nDe.�ڼ�+=������� $i�զg����?�`�D=ɚ+Ndm��-�):�{���翙��=�9�~d�!����Y����Y_�ߜ^BKdg5]�S��_P��v�`��J�-l�'�)�i��j�7��#U:�{O�d�$"lG�l aM��N�S��� J�/;�#���9�χt	,��9{ T'�摈3��n���_~��q�?,�!"D����ˋi� ���$3�c^6pX�x(.�8��;	���B�Y%7�󰊑(��=��6��-[�O�ʫ�B���_P_�c4��_�X��-k��M\[��V����;Y��&�����\41�*��7Spt
 ��I�tOeiaԖ�X���t`k�q�z�/�qhcb1�J.�?���~��4`��5������l�KbY|R�Z@h絘	V�5�r�.�zǍT�1q�܁��B0��>U����q���T|��˺x����!2�@����5�_'�j##���j�A�q+�v·�r˴�!��M��}$y�A�,(�i\u[�ɔN���cX:~� z�J�g���ޖ�VP]PK�n�X��p�'�Q	
���-�K ��U����
ا �W�˘��b�]7��5�]�)��Ll���y��W�7�^$p�&�;E��4�]`c�VjebQ	�uy����Czu3���~����D��r/��g
`:��7J�������M����~����ܥp���F�䨹��E^�(��&,��ܙ�t�'<���o}��{�*���o���5�������wQ��M2�#��Uu��!���X44�l>��e���La�zS�ń�bu�Tx�(��d#ʹ�`�0�/D��oꔼ���A�`� ?F	IsN���A�n_�|�ƣ�t�#�C�	ԻCȊ�_4C��]��&m�^VGX�(��XTe)p�G&;��
��h����frڑ3c���S{�=HtJn�mze�r��W
�4-0Q/LFi�Y{��[��i"�Tu��y���*�ө��`��Xr��$է8�׹"k`x�|�ZUE!ˣ%Vh{��z��&p��ͽ���3��F�$̨��Lʙ8�^����8z��Kk_�P
$���@(s��ì���\�}�h�GR�
hǲ=8���AJI��/arj\�����X��??	EBc�
LR��*����w�b��>s�B�3j�?�V��\�/e����	�n ��?��[�/�d�'8�@�b ���T\ h��U��G7}!j9��w��J<o��=F�"j��B��F�};���e�=y������.$io8�|�|��5��:N�@�v��w �pN{��R���Fl'�X�y���w8��0`�B�+uC�[�]*�xU�(��"��pՀ�u�
b�8QO1m�t>�)�{��<�H�ٓ7�k�P�>���K>c���e�#^��"Mqr��_l��[�Mn� D��h@�Sk�JM?��L������4Ƙg���L�P��TQ�i�u��8�p$���N�����6U�&��n֏��W�Ǹ~���=/�*�>l�7mh�aF�:��?��
�WmC��Z�0��8�Br��,��>��f?^ j�ɞ3�
AV�tHB�egM�n���i{�a�¥����֊Z�y�λd]7��2��u����M5�@ͣ���T���)"����b��&Pg3H�/4w�l
ػ�aS_ڹ�1�]֙\K����]�pE��a����d�(C������~�Ϧ�4W�i
�`��a�_�o�2'U���v�(�ib�v)��3�D[p��)��.��׿���� Zk��Փc�ύ{�p�b+T�w���D����wdY���K^�٥��Z��Ӻ+g�6�h�R�y?�߱Fۃ������@%�t�O�v��K׭����\k��i��n�C���*1=,%A�t@�)%Y���z9���gP�$ ����~�&����=כpg���18���a+Z�d��E��S�R�.S3e����St87�����;t�[lq�9&{jͪ��5��}iSY�]�ȸ�`i;�h���J&�����8M.�@{��j��-��_��Xa����f���_� $։�>�U��Z�t�q�!q�M�y�Xc��EF�S�A�����i��9�*;U�c �H��|'M|���<�,����(�x(�=���;��E�l��}[�:��(лRW�����Z��2CF@΢��9}�bZ���G�L�u!oА�����I���+���aT����Z�������/�*�,{"B<���I(�iQ�^�ׁ��n�5��3t����c̑�D�_M�(�;o�d��jZ��צh�Q���۔�}��|)�q ��Dѯ��Ĺ�#;!�P�N���ڊo��|(�qe.g�FA+�+);1�k�r�r��&_��S�ٍLm�e�2%��%-Ad���Bcpr��N���UE���e�>���jv
Àx�61j����b/#i5n$�S�v �Y���8��>��e��YS�`��S��S%c��,�8�^���J��z�y>c�t0��w�X��n�[U$�������uMH:�¬�i\���!��iG[����B��+8�S�ΙO�G¦�ME~7����..H�R��"$�y�u�.��{S����n���e�����h)�9�He)uU���c�uv�+5yH��V(4~ӅL��sX+�l�iKv�<v@��3����4ʿ�Á�$�y���h8�#'r�y2�/�|\Y��W�>�Pƽ��뮽'�4�}�{�Q�T3#VJq�)
��v������4�X��;��L��a�N���@$�4�{I)Hy��b�I�����h�it�ii�#�����+e������p��S: �ǝ��C���q3��bv�6�Iwc�B�B�U#�kn��()���{aY��!fV���{'ʐ%o���0���UsV=_hꥩ��j<y1�׏�39yi�R� �%�Y���&i�����x���?�:�Di�N�3d��=��E�y�����%,scd�ۣ�`Yxm�4��v׻�Kq� �v��js�H=������	�?���H�� LM�u!V�칟�����A@mj����������?B �:�V*��OBzy
i��AFƣM^��I���'���Nlg�/���"��s]~��jB�6�X��K�(�	����#�3�,%n�nSK����Y�U(V]�G�9c�d��bx��w��̷_`h9�y\O� ��O�K���?���֣+:����55Ǖ|z����/`�^��_^C�̓}���V=���,��T�/*%����wP:,ߐ�7����P�f�%��t^��1�ZT�A:r�VڸHk�I��şI�&�"�Ŭ��#���2�4P���v�w��5��8sm�m�-C��:����sE��LǾg6�-;�~��#�n犕Y�ö E����os����S�Չ�
U�����cxb��.����N�tgGֹ� �nj�<�0�5���͘��gq��i�`���r2��e��vl��+�dl����-�8Ba��"�9b�����rM膛D/�2����x�ۦ��3�k�cX>����G|R��˪q�i��4c�M��C��,FE!T�&���젰k��ư����o��)���Pg#,).�xРJF�����_f���o1��S �1^s�u���Q�Aj����*+tR�D�#�0�	,�ό���򗻪sBӳ���KZ#=Ox��'TH��ma�/�J2֝�e��̫��	-�,<��d�V7�ܭ�҈/�6�/n�Y�-�76m��<�NK�1�š~�&�����x��	���!t����W����ee�*��^��=f��4.@8��/(��2����-�h,�<i��[�~&Ox;^�帆� xU��qf�qK�_4��H�P?ou����/�]�"|�R,��cDCK+^�y`�G�
;��z���w�"W����;:�D!��ei��I���Ņ���-5�vq�\ ��w&h�`��GW�ܪ�a�:�:���8���k�T��ጂ�������A��=���t���F�j=�]�R�+Z�� �'���I8Ƙ����P��`0���6���#�aV	&��ZB������T��õ�����脌Q��4����Q���(��h*���C?yS��:Vث�f;j��w-MtT���G�"���bVC}Ͷ�;�	"w�)J��'F��J�D<�$�J��H�_�t�^���Q��T��(��'�E����U�o���؛�24\D��G-GT�С��ަb���
!�M#<��.���w��d��{���K��$�z����R!GR	�.><+6�m���$J��؉�2}.���[�@�U�@ɕW�
�K��W�W[Jv���
yAAb����ټ���Ř٤���8[֟�뺡~$#ϼ���dnD�TCk!����g_�/HH����lⰣ�W�ٌ�+�7#�i�UH����g'�����������;-B����fsUF/c��*���(Bڂ��:ii�Eݯ�%/*��~�tdW�1�f���|��c��>�Y#w���0c�(uah�{i�־�M�%<h��B�a2�&`��I0&�gћ�(����nO��$w��YQJr��H+��m<��+,�>�"Gs���-��܍eŲȩ�Xpg��1���T�L�pZ�w����i�s��q�������B��H𖽖!� V*��ü9_�԰Ϧ맼>n;z�����8G@8����i�nɺ#\>����" � �hj�K��z%�x�x��k�_��qI��k���c �ʟVC��[$��ݴ�]��� &�isD>@K�B]d#VV:�lᕠ���1��Ƒ�G$gqw���k�-�Rk�����F�(\���%��o���$�(/��[78��)�3�JD��,�X����P�&��;�$�N-E�����5@P+-wF���I���~�2�E��p�9����VU��R��+k�JZ���N�>$̈́���|�
��F���W�9��)u�܇=p�v�ϧ���+��u���2 g;����n�M����T��6�E�$�ӆ���'�إҹ���U�{��,��#�6�` �2�EqM���_ˊ9�F:/�I	W��"��Q!��bF��m�N�鉃"+r��?�t���:)���6�fcP�gς{y�F�}�j�>L�x�KQ��5�U�7�l����|���F��.��U
�d׸˼�sa�TX����?�tK�\�"!��q8#I^������Z�^c)�f~��d��p�3]�aoC�ߥ���N���w"�����o��5�Ϟ��]Pj�J��%|'�|Y�+�����ꐟ۹|��jb���tE���#�(_�����J\P�h҇M/����R�8Q������3W]��EZ���������$RX��n5*��K+:ފ����V���-�w;����g�F[^�|��=Ѕ{��@�,����	��ʶ=Tap ^�dK���wGu9�������Fؐ�e��`�ؗr�0��т�T:��I�V��������G3A�_#,-�/��J�*o1dȓ���L�Ac7�C�+
�ܕ�_�1`��TP(����~f]ݗ����*ߧ�চ�g-��.ћP~3��4��� Ks9��w���l@�`"�@��i��b�j� ����S�FP������Q�\ȟ�/��	F�ȃ�s>�r���S"k��k<yzO��k'v�!NKwiu��_�LKX��)Ω5�Ąf��.;�Z^�e�W3^���o&�у#����@��M������F�=��e����Hq���q�*0�VS[[�﹎[}&q�+AU4��d_>�,�؏�%S��D�9@Mɫ�	~o;��skXz)cu�sbqB�CAQ�0N�����I�-3.Z�7A��JJㆳ��7���o��ێ@��!)v��3���mUO�>��+���!.߇}��<�g����jw�"�I_15E��9d�υam��n:��"�
�Ug��G��@��c���ӯ ������ �Sj�b3�:���<�*�Z�v#��~��\F���Pg)�1u�ˑ9՞�<�I/��v�nud����j��!�A"��S� �p�9�9��T�O"x��7�}i�y�,�%�.�o0̆\�p�l�:�._�i�6V�u�}���?�T�Թ�<��c�����S�U����w<X1.-��r{
�TD0T7�O�3�(����v��HY��)#6hW_ܥ}@�KR�����[����D�զ��9[�G�mdL�M�_�S���.v�3�4D���q+�X����/��[��9G���
+ޕb2..ՄA鬜t��Q��J����ԏ�obae�a