��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P���S�25"��<���5��+s�f"Em�=4`x��j���n}y�#��g3t��Cq�O�$y�,��[Ј{k�2�jl\��dO1���-D`��/�*��d��ep��z
(���]	�o�9� �^�&v*yt@��"�@��pR��c�)���Q=[�hN��)�L�?2#	�_s��j��B�iJ)����u���&�D� !��&[Q8��}ek��n]��(B�P^4�~'�tg��_p�����5�)S9���6>P7�	u{��Ŭ�
�A�	�����O���'��3$����Sg�� 5��vt�B&��5e�?��6�v��ko��A�
�C���i��+���ۍ$d9�gzN�"���{�P;����#[ފ�(e�H3г�޿l�pfs��Q6m*|Ҙ��?�4��y������H:2S$�S���S,n�Y���v\��`<2dT�l�-6�<��#����9FD��-����(�e���9ZZ-�v����p��m��浩�(��Z���8�׊���y����ע�έN�9�Q�]�j�=�[����K9Jļ�rѼE]�ן��Ф�J��,.�[��E<V�f��׋#+��'��X��cm�=:{��;X8t�����`�>Yl�y��Q�;s_`��(x�1��e�6���m��ξ2���1��5��ě��.��a_�<[4�m�B䚢�
^x�]k�k���7$��9�c��GM�4: f��1�D�k���
yeJ6z���w9��;�!���,��{��g+��a�p\G�y��{��hL�$�h/�ܫ�2�iX<�[���	c?�F������ !u��S3}�(� ���NNb!��H��-���+P�,	��ڠ��e���Bx��ǖ��:ޖ�U]5v��bU�;����hZ	a������@�e��ks��z=�S��Wㆢd9���SM0���1�d>�<�����B�W�+���u��%��&UaB�fkK�:�%|�dK���JN�0GDg=j��Ħ���� �.��=���<-�"��������/Z�>�Z}N �z/�+_��'k��!����Щ��@�(<%�d0R�+�^9�q�¼��PH����W�����=�,���c{w����~AA��"]6��>d��9�r��� �O)����ysm���7�m��3����G@~^NM�ܘ��/k����W�T�%�m���⵪�ҿ:D3����AE�+�x�Z/I�C=J�nF�.�8�3C�s1>S �ek���|X��:�O�*��ǦkD��7�hk]����r�M�?l��d˳o�
�7��A����g���^�DHӚ��RU�%�4n-|n�A��.U��O�m�n]�:tO�S���c��q�G[P��<�1	%3 �^������a>?H}BOban�\滫� s7���dy���� ��sظ��j;cl�o��*��ӣ~~w����"$��y��Ӝ��!y�n���DB0H�;�ӹ,v�6Wc��]�������:4�Z%����a��!�W���W����u���p�k��L�P�K ���IVoeέI`���5g ��O���<�=�������&�O/HK��E�3%��S����ڦb�o^��^K�j��M޸�#x�`�m�(�5oS��wg��j��t+.	��QVe^V���dNM-9��fBr���J���	�B�C�����ڐ�K*N�ohSJ �v]�Sny�ȪI��r이,Y|��� ���gh����Kp�4p�8�ؚm��> �gT!��)m�	��6V�tkQ�O��7��4�ʑ_�)�@E�8���������9^�מ�������