��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒�� 4�o9'�QZ�����3���m���:�Y�_�H!wI�O�n�̌� ��U�[���礎�U>���`jI7�j�ϟqa]���Gt�b��K�B;����w~s����2
]$>�:�[��
F�@j*%SC*}(�/�:����.z�76q�R�\V��:�?RQ^Do�隣��=i�
>��z�"���׺�qĵ���`g�,��9�G��p.��j��j��,r��[��]fz� ��/������B3�V��G��������9��BJ_ǧ>��Z�r��3����Q�|ۆx����"������U A�T@�c�,�W�@����?'�f��zԳ/��ڎ�����/o}��.��Vȸ0F�a�"��L�e������p�Ű�|\O�a.���0�����h1"�t��PD1��~�#*'��""�{�
Yv10�2��\$w��W]g^Y��i�:,kj1*���<da��ф��|�%�'S������6���Ó�
8^��;��s0��ғi�,S�j��_&_�)�7��r�R�ĝ�W���F��0�7���X�l�0�� #<,5���OZ�PR)L��h4��<L
Hb���l����JX��Ȧ���;	�CSz����`nw�d-�%�����X�S���5铟H�	H�Q99�8���&:V����K��=K8�2����N'������=�S�<BL���p�$��ǟ���`2��J/�O1q�6�j0$�����*���ǽ�~��EB��3�%: ���4;^�o�P7`e�J�&�L9�A���1�&aY�H8u�U_��_�Y6����F�o)2 <}�\��	� t�m�����������G�^y�/|J?_�h**�5gW��1r�u�*��Ċ}3��*����oXj�t�:�IA�PK{F/����<�(����ۀ�o��W�m`M[��a�Bε_��n��b߯`xep{�l+�a��f�Z�J˨�$?Q����_N���vNj���Q?��羜����|s�7���i����p��8�gs�u�vXUom�J�^�8��x�
֌�V�iI�,��+L��I��߶*�9��4k�mw���'�m��O��H�PK�avkTQ1tc�!���%��t*v���pk`6��iΌ1��g����	co\���o����H�Hs����I�3?3�M�W�J�F���� �a�e�F��?��5y����"iBNݲ1���ի��b#���nH`����i�_��[��˿�\Pp����9s_RG�=�@i|��FKiӪ%�?f?~�_�����L���*k������m#"�:ƛ�/W�qQ/�0�����&aA^8�}4|c�%��T�;�Y�?��6�������U$�]I�_vg��	L�H���ۂE4�9�=�,R�m��7a!�n��Ǎ�*�C�d�7�^��!7@���m��È��b��(Ìw�E�7��
Y��<!tj\��Z�jNf�s�ey{��Qv.B�ű2DU<������V<�ˬ)���2�qKX�j����8/Vj����8�x�ܶ�?����|���ĝS1�2٭�H�K-C+w�����X|��2�G�ѹ��:��Ru�!&(�� �F����<�W	$@�fϜ�C��P����>���M��8꠪��i�rS�8�ӏ<GY7ij�.��5��0ƒ�&�Ȕg�8G[$W{�oN���L�[v�MBԷjӹ�Q�N����p�7��@I���S@��q��yP�i���	�!Ø�Թ�{F��)^ohA�-����bu����g�?í�/�3a��M�/��ޟ���$ ��0��o�Il?9��;r/�48+����h勾f�F�a�� ��I$��ʙ��^�#���R�����$TT�3��Uflg�U�I1�!gfdd�S1�e-��yV��!>\O�H��	���e0^�qz������G�����*�)(`�}7�'���n�H�&:��EҒ�?rRX�����r������� }��u~��G�Zt7����|Vgй,`s�h�^���$���j�z�;܁�%���M��!^qd6����:d�$އ� �R��<ږ��7�&���O��6/��Ȟu7$�@�,��$���$Ɂ�����l�e�m�K����m0��-�X��Q=��!ے/�}�,ĨA�3D�o���Y���LJ����[�~�B5���:���Mp�(��;؊�@���[�JA×i�L�ӈ��5)�<ʄ���K6��8�[P�S�N*!�j��� �D ��w��;B��ʕ�� f�h^\dr>H�3|����R���C8���<S	�.�����C$��e��jw� z�l�3�'ZH�a�e�2Qw`}�'�1�e�a��e�w���ڞEX�_rJ*X�pV,�eT�&T��`��7BZL�8 �dW&�q�5��y�q���0Fp�=+	g�8��?}N'�����+�dc��#�7�^�G��5��b\[��y]�6=�v�>:&LY\~T�'2�)�\#���U: �vg�­4�/ ��X���7{�_U��
�����	����5�n�=�����F��b��zԀ�<%)jHj�G�`��F���G�
^`��1{]P���T͠2m���ɔ�t�(�8�i���@�p��˨�t�o�0��cWT)\I�l[ ��6�s�����B	�P����C��&��k����ع���P�왽����E�X����7D�P&��n�������c�Wֶd?���)��U�)���V�L���I3h�V_w��f�Ǧ�(��ޘǒ����y�Q"?k3�8ک!�Y;�L��R��0h���}�\yȻFb��@p�(?
���:�4�������š��S!|
�e��"��
ۅGjŊq� f94;Ul�x�!o��^S�7���Y��Ƿ�,�ْ�r:��s� �.�����"w�\��6O�'0M��3ME��a���J�>��:a���[,�L�LΛ�<Z�wh���[f
�C[�yN{s�=��7�pT�ʃ|�w�b-����\�Ǳ�jq?�1&�",��:�j�p�+*Ő�4��ѩ�h=�f���o��{.������*ά��������I���`J�B���s��2w��ɥ���٠�a�P��n���&1'�]{�������P�w�Ij[���8���DX���3�	j���u�Z��S��+���.����~�ޑ�V��g')xN���x�/��������GW�&�_$a�F���D�hOG�i�s1�����ڿ4�\�::�l�Лێw���I��}����jzbب����r����- �FCT]:W�^XvFT�������VU�M�p�p\gC>ν<렳##|��B���qh�O|B@$����zxOS�͑�^0X��@��W�A��~�y�j��)�kK����Y'����>��a��ʟf83�0�R���D�*�����;�<���E��l��^;ݜ�5��$�B9�fc�)��r���	��)��x�@�9?�f������A��5g�C�ؚൔ��NѻQ��}�L�W��v��7�^��e�к�<��/N��z>h~���+%+��Լ�!(�*�P��7	��ͩ��2bR�P�v��ĕ��Q��&�^�s�'���Q�k�o�?�G]��e��G{΀�8��ہLD�k�ʸk���] �������az�³5D�)�8`hPu���xM�&�ᦪ6en�ɝ�篈 ��I��e��t�8�p����*� �S{�%0�-��>���G b�pyڐ�K�>��)��L��?��yw��sџ	�ɐ{=~(!Td�Q�����V�
o��9�|'7�K:`h*m���=�0:�H��(O8��z�@k]r��Ψ�x'��h� �u����<�<!w�� ��J0��\�"iA(�~���h�����b��U(R��HU���*��ʥ�6�q��b��OW�dދ�r�"Wq�7Z���|�����2m��r=1�T�Qd����6B���k��Lq�|�CQ	��Fr��|�b�,:� �+.�_u�%��hd¸�=�m �b�1�8����y����45W�<@Jߪl��<��
����������������'��ޭ�E�}��""����m�>�$G�|��P�{ePM�O:Iڕ��0��|�{h��*l�(ƹ��� �C&G��oZ�*?��F�DR�U��(�eB9PN�~\bW?'��U-��[ea:49��h�ւ`v.��?,52'h2s�±V�o���L"I+�u�?!Ən�ϪCMR�_�NǱ�)9R�b�Y�􊪣$Մ2Ǘ���r����$܇�JM� �������Y��τ8�kb�h��W9Z,ߪ�=�d3��y�"���)V[�r�|����+�ޞE���\�
���`��/�FM�>�Ե��3>���� ��0�2�(:E�)
��H�%��ٙ
��j┫�X�Ϣ����n^,N�R	���L6��� $Ӳ:vUc�<;��+��*�ξ��J��L�"w��򐟎~��+&v��h:'kP�K�۠�<��������NR�^����r�p}C��5��bp�70���l��1>�F�vE�ȝ?��P��<���^үzSK���{I��u��N�)����<���Q�W��˲߷;%��ۖ�?��;|�fp��?��@�����h�O;�}�i�<U�D��vP�I���n�b�Tp�p��/)D�U�S֣���䅇u;�)C�/��4�<D��sY���+4�$;�<4\��+�BZ�i���S�A� L�У����T��c�>�1�v��u��b B� ���-�{�ռ�;��X��5&q���%?��s�� u`_�8��Yȵ%���2Ն�l�Rd�9%3�ӓY͍;�")���u�����&�zWy&���4��!F��ҋ�:&?<�2AE���+d1�������h���ފ��q6�S?M8.��'�}��`-uX��r�q_
l1���'��oj#/�IYi�� �?�X��F��n'���=�x��m�i3�����oo�P�)����6�P�@�<��r��k�b��ppOj�G&��T���k 4�R�&%6.��4Y��^���fe)��ޜ�oʀ�ʛ����i�F�A����V��e��BG� �(��F|�A��a������DN?8��1HO�G�ו:�����(o�5p�����-�tRw����i�G"��{�2�:풾��G�~�2{�o�'YS����[}&uj����b�(�ى�X)M���^jQ���ܝ�=CS�~�PN��0��.�R�z3�����70�C1E��6� .VL��j�9�˵&'���2��x^z�Gg��aۧ���'�Q�U'�@Um�|���$�^�^���'d�F�@s�� ���ѓ2�gCL)�
�pd���ޤt�%�PS����P�τ���"�Z��v"�6DB�M`{���_a)��'l���U�yH�y�/�=X�ҳ��kY�����^(���8����:�����6��V���H~@O`����+B!�XF�r{�֓m��)�F�:��X��� wHp���,@P�K�����o�1}�P{�����Sy����/�]���T��O���x�0c]�T��t��wy؝
�Q挦n�YolS�o��=�R4]����q��8��x ޭI���[�౧E��]��R��[���w�O��D�{�)%ֈi������cB�����N�o���������Ȍ�5��!�=�mo��,�Y��p�}��K2���^�Eل����*ȁ�9�uW'Ǹ����QLK��m��?��(S+y������M_����6ܓ�B��x�C�XfzB�)�Xk���3�a�&uJ������a�Nϵ�5��ݵ$��!�9�D�gՑ��?޵H��^���G�l?a{񗸐;cܐo&�%���k�^+,�O���#��ͣER�~�U7h�c��շ��P�1�KHn�Ļ�g���b�v�