-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bAoX11+eSCnRCkXrjpahGp6+WJq+sEvdTWgFBzoVhe8SjmLr243fmy01Ky93nnwOrfK7x7ObUQFS
+hmk9/gIZnBXVrNlu4WMvJEKB2hrb0fpcSJrx+0Oi1ToMr0inDIHCqY/bi03LzGpnxLkWRynZp2g
7c6JjiaD1+uDK4RbMBflRvzAqv/kOgpa3GPZWdoTAqq3/vLmuY6Lg3y29xqbheKbPm0/ugV/qRWT
b/Wwlk5t/zt+rzOx5PYpQrUjywrfishO3qlIcSuUKXNr+0ony8kIgIpPMSWdPNX5ktg+pWsfaP3X
jg7DLyyXKU7R72jY4/dp6tT3eXkNfNCrLaviDg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
HmCggEMmIIZI2dmISuB0gzT+trH5A2wNWOSQKAVHwSHd9Rt4QckARrz8mprapV0oG3lKUDWH029A
bVHjhBEpXKpxrdPxfNZ/5pLwBiFTsPZxUKBd6wa+qBJTi8T00mc856POrHweSNucWB9tG6I7wkpN
ZQQ4mMGMBZsMikuwqVfIjfNfYietsX3MIZ5N8t8ARmfJuJY1bmlCc9nFMJA6sdUigU/y0SRxCqlO
8/gQac+VwJvy8+sx4vxA265WtnA9iqUgKTHiFjcRPJhqP2wssG34gj/oT7apNaAdJ8FCPH7nxDN5
fpNzVO9e1ty2xlD14tMNacj6W5KSykWqDmem0VEnU2x9KNgyQCrpplGgAe4FZjvijTpQMkYnwkWC
M9XacpoILAOFM6WL91RDmv6iRhcOw61ygCD3bMlxlM3CNE6ZdUvbC3zVHSIE32ZLrMYp8uSnm1sj
kuchpOkYUnRgPWs0UY0wD+O/Q7XkR+42Zl0e1/BmuOvI8hh6yJNyy4iyAQWynUL26CM90jkB4mAx
QiRf9Q4KIa9BJ4MmjChE+GVkd3cIg1qCNOeUblgD7aYAZdtVEm72Z20nl+DFXSAlEdRHf2J1VZeC
athcAUy84UZ7B6XFKqhBjQXa3d4wPhVjbfTuas/TBEeAQwsC/JrA68F7EdbE7HcFmRxuk3FxHeLs
zNwkqkn0HpHUJjn4LPkaFCjcvrGoAcN5sjoVkRd2dPWepO+jivFPPR9G5f6vhzY64AyOxJr2G62V
8OlpliwLgqNx5W2NhtySNMEGtOQs4MPYv4hrYDRTL2Yr46V4Y172bpjYXE14tv2F1alI1fVZloPZ
KJvuDsIcJ57DYO83S9Bot9lVx01nD+8eX5GnQmUz4clGLweJCQ5Cu8Fynkry1m2UB7X7WVqMi7L7
aTVdeN+lKuHSldJvHNNgxqDcPPgnsK3pGygB6bYuBS73yFWlSza4n8J4bglGedNBH1a7yMlDGo/O
8y2/LFWAeF5ik9MunFnA3FbrbB6sI7VtztdAcl9sHpx0U5ACGEVvY2HZtdCF3TrNwV8P2mc+NH4L
zbClY1vG0NAkhjOF585aflw5MBd5z4DBODurotZJDEWIqmQyyJmBi3WVUD8ZctWV1MnffyGvXCsD
TjSCN9QcRrC7gU7faHEQOsjx6mKA4gdzLE9Vd9iDdpPWTFXwu81QSqQeCQ21cXZEVjO7l9yomwmB
az8kbrGqxv68IrG63Yp44ns2gXqMOuIqTEnhQxjNBJHDPIm8sbVbeTTwi5Qg2UhG+7/oKJzUc2YP
TLltJoO5DbVhoIZ9p1WQIwICFV8x/9U1wQ324BfO4nr7ypz69b6EA2JZ60twR/0ZLkFcrM1LaDNs
FsgslW+pej3NtodXo5Js2wNAyDKL112BZ19Ayo1Ess3ZPQFgjvhq1oWhBsC0T32nrbVjPxwMpq3m
siWZeJu1cec/lhC2OeFOBr8hIl/os9wWp0CyUH5yhx6FjLvk356s0+smyQTJuAoD8vEn8pHjyVqU
KI4onbOI9Zs5nWyLqaQjORjR7BanVOOSVnmzn+Mz/pE/k3H8OUiqUNw4rA+TmwGaxDKe4Zlu8Mq8
O+H94TuAlAsHhh9RND0f27rjOD/1pFZvsoy7T/+vJi2wtKdo/1QUl4ajlp++DZIpOuhoD3DWwFdG
FcM64DS5JE5a5gjRMiccLrOJKnMHXzJNpjlANwFZqePUzkt6xC9z+jH+MdK2phThNOsCV/GUEW2m
wui8109KTA3J5c0XX/RryKxioH4qdeAJGH4lzIjaKLkzanITpe1wLjsQCT1eEWjyj+G8TxAeY4m8
MgeEjsBG7xK49sjkr4DWQ6zn1Yx3BcamPdJrVnbGVzv9Soztnspb93DhVDRAy+V3Tkpu70E3as7w
dZB3s1GAHy+vDnqFbS5yLzM/9MlDI5raJLkoJ8iGzpmZDUGW++imwR7hKF7+dWpNWcoqtgOwZXDY
EVfA3780WyMFmAO8letafiNmWO+s42kcilAO+ddRaZeXc9Nf4SYHDgsBaKs7WWE3jcAYWrReKRRt
khgQHa5J4TVPLSx34lDGPrya5fq6T0rEnfyjFgO59PSv45RsZ8G1e55GqT974Bkznh2i841vtJrc
7hB2A7agDLaT4EhtI2ECgQAQQ1ksEZgvXSZ4CdE0t/3ctoHLrBVUN4BSvUBJYLG4YUvcuS5TE63p
TOU/xTvZcx8V4I7jxxVgteScZQUUq5Opp+yQMoWnVkBeEfuzy47GAMDzc2E3ptDZVLGSCnzNohr4
YN2a6JB/GJvH93pyT442+tbxhUpdsVYtf47uO1RoteJHLSSFC0Mj5UXLtUDFoDgKSJiEf9y+4ouM
673YPkI0QwFaqTIfa5RQ7GBp3bfaKNvKLnTnjUqMjqbxomYAEz1aziymEGWTGfu+1/pM+LyYoLfK
2WgvIHiswob6+6U2cw6XqCFWdV11kRhyOeB/LRy4NqcHfBphF7GoWQbn/vJbIirfAa74+WRZmex5
NuTAN/51ldjy3oQ3E7F8WiSDYp7DMq9DlT7fPxpknZTBSpZKWo3xYKW75hC5gVHpWc4M92GudWll
jYMcHVEUCGb1it8XcNwlkHAL3PBBHOKXcm0NbVq2ndSZ7piE1mb11cRk6LkOZkT1mN56pavmfNpw
O2tAsp48H+6DTnu/okQx/3WLAALH/0Bd2mm3nYg5zSJcWdgnXC9o+/rq3smKQa16duKDlT9kHPYi
qk7abmk/22cgxRqitc+28PFvLNlwstpLTAEHM5ym9A8xjvogkPLC4bYXY83wZOUtOegwGXjPmKJN
f2y2tj+TKGB4Sq2SZbtXt6UYw8cp77/JokbJzg4I7no+A46rbjiuXGoBGFRVs9VAox26kEObAqSl
A8v1ZC2WJv8hVrubQHrB0PmX/6RINrDYpcYKzKXRMwza7/7sasWTEwzJjkDrmjuqC9PpBI+lpsSg
42KngBas+hsGin/kOx9+BSPKftKsriVJkuZOOvEpX497zygydmp4n11KeiDpE+/JCfEAR8PueuFA
as6zEllEqiM0/tHjVGXGLoV+qlHBIcoX0akezrTmb9lX1D6mObi9+xFp/g++UVuAGK3GuAZ//Pgx
Rn8S+FwxgYUow9jtbJe2quflp/oKbbZlqnVW4SdnC+4wtqNDdxqwETMDsICEI6n5qbYGDR/SIIm4
nQJzVRuTyaKPRP1AvrB8LEY7wqKzRnUSz7Fe1WdjSMasqrLXmagcp9OTaNSl/cxhdi5ezmhb2foT
7zK2b0rTvhMXQPtE3fuWAgl7K5iand2620d0nq20U8qKxLQAJPV50jjXjhkGZYUSr1VgXoLy8J32
qph7F8HTeFmn1p5HrqbXS9oA1PcFmYQ7ByzBb+lDTWlZ7ndyeALL+7+FXb8v0RRHW24AW2NXPmHA
dV8bQmlxDSd4PWZZYOONt+ZTUL1EBjDQivy7P5P9VsN2DJv7zRHw7LPP86EuOyQYhPChxc3Blawp
EdfH55lo/dG8kMMi0qhjNocCfpty+kwI81y7WTnh1so9nGxtFakvmA14jlMlxLBUM8/I0zYYh7vr
zpZIX0STF+KLsnUgW2GmBqQumYP9yyi3OYypTGLtmzqpC1TP83YPXMXkeJRLPwhM17YlVTWd29Hz
Fd6JwQP/699916VJWZtukE6HS9pZsIAcIw4abFz7hBtKBhHt3nFLgB4EGtHCO99SWpovwwVvgUbF
CvsqJYDKGs/SrGnDSWVgRu0eWeT4GUXJym3muGS9w2gVF3g/l3tWLqOI//rJZU/tNA9dzAP7wb81
2CB7jkfddnMU0+TI3nvsLeRRSMdfeCQl67tnYXUvyTrwPSvnzFJBhn+prmYyfS8HTK95Ey4o0pve
7SmzuyLK2wFC1539lt5vSCUDir/lyjqPucJ1R1HxgV6UHWHl+VB2BeazLz2nKXaOOfp4MkRXQrzI
ZnC+GeBZ45uSSr+9paxlc2zvS910m9ypJmSY3bYoheBLu2bdYn4LwfaWZY2Kiu2+ehiBUIBU6xOd
LhVN/Mg71ftQZjRwersgtbKXh4MZx1TTQ+WT+Wtl/DklzyqSKGaLtwV66nsdBxTCZnaKLuuFt26Z
42LTZAYV7c7yEEPOBcsdzrC5+tjIBPM1daOmS7Y9wrfD9yH2jv+IQe159qAqUl8MuGZuSD01+Kmo
LEJgVxlcHjPWXggXY6XrNb3HLfNWOhfuVckcVeDyOXRt6YeJsDb5E7Y5n1SSMp1I1Enkh98/njPt
QUC6ukylzaslqYldRJFPRy5sIqC8hxR+Nfo1Sid9lm+tbJOok+s8dMdOUVxuD/EbjTOO4ReyerAh
snadIMsH6RM80JGaCy5TJfINUB+kGEJylVw2Ui9VzOwOAnwVXyRpj91Yzc05r9lPn1Rj2mRoaLjc
KujZxfgnJSL/fGHRBZf7iTG0SkzxnZ4+08PWjDxAMUA0/PmqIkaJms9gYWzb62rU8B69X/h2J1J1
6a1hGJ96MwknImIUb90umQxGE28CWMqstNlXot5m+V03MyuqLgX7uxntO3qpNzpp1ZU5VpqNpe6z
PPNbaDvwYdWrHb2tviI3/G3mHqQzn9XhLN80aKJSVCYocn+4KRtSi7SVgW0VSzufu0WTw3FehpDF
SxffzM01+jZnjJFS5tGivB9RY/GgeFQZa5AvEfoDUNSW1DxxA8HWa/IJ2em2p8AQwUqobRUwWYgl
/lV3XysoEYE9Yf6Bc6K0vJG9j933tdv/vqGteyGUxbVFa9x9OADbuEZNKwxpmjRrQQU/s4SuDtbZ
9Yb6KGiFNWGiN5t5MpAFPUiSMH2CC8Yf78i3e/xyk+C5hAKYHX9XOoSJR8Dt2INaYLJ6OWt2niEH
tm3eKTCdCJaWun6w9Z+loM3fmriNKOkA7YgeehFp7uKtv35qYhn5bm1tlVYqZcrBTIAIa66NXAw9
2+mwWxRAcfuxAXtQuPt3mO2KbU+XPPjgDM87VPiXyf2QuCs91Y3VbueIpj5c4i0unSSzjvSHVrdJ
AeBNYMrz+SCUnY3WpTitB2pdKWnGrFOo2W+W6JSDyDw39P1AerBtix/g+qewZqc7hTyeUbAUr1W1
IaWucWcC08K8Xc9j9D5H8sODqJLAsEY9X8Ve1guDSL401yUlcLvYyTqv7Q/6AsGYNEB7HyHuiqj7
Q8BXh0SZFXfVdA7CZxU4dP0WGGJzOVo3qqI6hQ9Y6GwDYmaYGVFgqa8IxO34cHNcZqZLGqM3MxKd
MOP0JEFqfBjEeNBiC1w5o7skIOVU4mAhGjXIgAWSrOTZA1jYPUQqssEDbb8bAMlkWLumgyGCMx2L
N4/Y52w4lUHJxplNG4U5UN229WQyLP3wuekGzL7buwUwq4WTfYXrlE6xGlXYi8PYnn4Bt34gQ2x0
vxpoBI0vZvHaVkmZEbtYb6AjDQFlckQiYE0tvpzUkFSf9bbycnRU4rLoGtPzxDRjJGT05GSIRNHs
xnx6SvCpJGM2dX8zQN2uLl3JWbujPUeKHOqd6jRHNfeg1uhCaPjaXZkduN/TuSQ4KVyGNxY518VJ
aTeABbKe+hrSRAcFL/UtpJbWxhdmMGlaOsUgnYvRFIqrZr4ov0NiIVnMm+EnVHFjfqNYKswSypIq
Ajs+ZKxj1J8nF9M2foLQHLzPwp8hD4s69eFbyfXI+93BJzJ+f1jQWrM2gWkzVJwHCRO4eSs/eJ1o
oTNera0sajFoyMKfT24GsKW4NK9f0Q1bK7jxC6kS/ZxBqiC5wVYvHHTliTO6OpToBJ5LZ7bySxCu
Ca7clwEbFe+u5flzcdKir/ARD+eSafHm2vsHmEqDbSJNtDvVTs9gouwTa3GpGCmGmogVgXPcj/be
QhxKb3CLnwCETqksk6LQwKnsOSfkIQKm1Wxay5pulDSCr1rVgSyE4AzEZKtDEn9ja6Zx+6wJOa43
eLwRhP01kYRgJgyZMQNQEwnNECqGYlir7scYopmCHflYu0CRvIbJPJvczFhwenyExbOkjRaRQs/L
Njkt3TPee2yNhWUYamrWlsOb+3qtBXUH+z4F3QhHl+cstV8xwUD4kXNahhPKV78J7zpY/TKQ0OAJ
AmLvrCaUW26YnNR641ZeUrAXVQ88ne0NKmMVdcJ9gvnJ3xtag5IL0lqcbnmm2IYzdYpCC6AN6pvg
cLwAexKLQlvK4BQ513GIC95hbhv90IHrbU3anJI0bt1vgBGPXh+S9wbtFq5TMS0eyP+YSVcQ+YcM
35Dtd5VWFuQ5ZjjZQRhxB1jOORMsw2euBOd58oXVhtds6piY9TE6R3aPXo+h0/otkpWThpDNwR5A
eAvaferNPYgjiMKLMciGrrJKXqReTzT93B4adVu+6RO9qMncJV7QsISlWbKUfW02QByMlwS1QlTx
kr1YqSB/NcohvonOOClmIrqe5N5Rd1hEcvn+jWPZ2BZymuUUxbqbP3YwUqtRJ0ibJ4p9uGWQEZdd
aYAIqaSR0nNK7ha66AKsIw14mr2yIeeI9DuwLfQkLn7GlbrMHznyaSKEafTzcMxQL1tFnNT/edhp
kBTbj618hjAHJPDeGLVdSObT3WKVAVvt9QiXZkTRpQVOn9RIRP80vcTSDMx3yF6SlCc7gv+Ay/xp
YC1+U1wh8cCgvODm5kD5hyN22ghGjYFkHrB8J0J1q65WTWWIKBInAIWUYpXMC5102i5nKkXv3F8b
lfTgiBcmp8uFWL8dGm4YfZ0QNM7/Ww7Rgmkec1MQueyuIkXfb/ddjd+0FNCEOjIHBCBe3DGQjcF7
PUCeJHCQePtZwW6iUZ9ib4ywlZcjB73hSJ6KtHu+bzFYAyMaLgMYKYFKxjXGr0lf7TfLj+fxH+D8
v/HhX4bJxlFzjLUSLTWj7smnKv2ChZ/LZbYY7kchU5jdf1y9pmsHluszY6mNIoECNKnrd3Q6H/eA
Wr8hG66WBeua7NfhxATK07i9JQ2dYRCsafHJw1jLZ5LxeS6OdHTW0zCfzA1Lm3AQ3GKeJBOMzV3s
9mNo8NHJHHG7TNQCwGWpMXeVdVNHTtrV/VeL/nz2jJUblABh9nQtjPbUBZ7JNnft3P4AiOCKJ9e0
MRLHIHj3r/0NiS9H/jUbCC1uGrVWkEIjxh7ntOz8NYTx/VE67ylBM99lRUYljlj0QRF0o0CEwbs/
2huufO25OU7wOzoJYEKpYJLXuDkTxM7pkGqtodmKv+qfOcbWtvEKIg8H1EX26Gc7nDCwR8MpA8ok
bn3cyjql55cr/pCQ1FbUFKh+5tfCUB68LvV+YSQ3mToXlnHgtiJ7woibq91sYWCar3l/V3pnKS0J
KotmMIkTafWFXL2AbfO9IZEhYQ/kHMEkw+DNPhiThdWljdxvjq+kiM7mA1waFa1wF9uILHSeBBZR
GfbmplazwOmmvvl4msPynzm25GV3iB7QxVSzo0NVpJaH7ZtxQQOpWJwdAhY98vSXGJidjayMPmB4
GZ+ilu85RAMezad9ZCAmKmIvkoTx2FrMib8/+5Pw4CXA/FOPKqRuxfp7C6rhPnX2rdfZW7YwOMYz
UJP9BNT80w/ab2x3Wwpit0kku0dIOSF6bl6vz/KzBpsKJI5QKedTkkuzsCsc+VdEUptdeU+/MUoD
/1Xtg6JNW2gfh7XC/+aSBbea5RiMlq7FePZvSlNJxCbrcDXxT6eWbaQ24aYvXAKqRpzOUG+RPaRu
QRS3hU8NUNJd5NWGTkBcag+ZPo96VoFSSQwmkkoWh7FDSFbKnR2n6fb9flKflMi63LF2FhTLgQ4e
qRNjAfdgDLYHMQlmTN6Lu/kkFahKpVjtNqxb5XSQ4vKoD2yjG3TheNnVytNldRBTToBcK1wPzQ53
/RLsMlwYgcDDWBlfhOpSlBMg7fpip4UghZOmdOIBvnh7baaK3oVX/RwhXNUbkQc24AI95boD7EYW
4AjPz6VtN2zRHtwQ3ZfDpzUzWD9v3a5wfoL+rdE2ezGtEVhOyirwb8/VHXeQqrqsoXyyrT6r27Tl
bAn+4GVAf3S1+Hwm5cDd7miYSJc+vs6PPlNj7+ESNcHVXEXSMCNOyRW1m+f6TZVwBUdqjYR3oYWa
GsgzROwiifSGTqKUO5FCpXklMyp2u5Lj8qKA6uK4xJdROyztih/H4caRGnrHqonoYCSgAygB19oS
Sxu8EJrRvOqCcUVyCjLbGZuhnLvAdV0u3WaNLxwDmK1RpJ1Imd1w6UmL0TI3V/D0Wdj31fdyuaa6
KNRIMQ2Mfjl0rRFMvBP83fXeFJw+5SdWEm4DyrEq8xCZ9KBegiyMK1Ysg2tfaQN4x+43Msl2xmaH
tJ77VFndbg9oIHcImKWfISrPyF6RPjcbEc6EbO/TBPn9xAQgCs+RPHwBmsgo7BvJdbNKVEVtsfeE
5KcmhEKIxNH6aHSig8wTyDvUQTAx/rU7UvraWY9rsaAO9AYm4Jfi7bp/DqpYowH/2SfFYXJ4hgqV
BJVIhxj5KmcslH+YgPg7UMpIDIv2dhiSfJnsRSiKl1RfvIDITZxGS3lhK/PhV6teBboqhyQC1pj/
OqdnQjZ3VT1vOEmGhj1V96bpIstEKE2L9P/aoLFBa5QEOPpmvXwgDfm13EOkLySx6M7WKDmj6/pU
D8/880iJ3JLyOpmcw8c+loxsJ7DW7g7WH4i6HUwhuyJPqPdAQOeCUkELzBXW5ESO7m9wEhoQKwHr
LldxAHW/qxRIMe+wz2ERLCGak9aqoSiWuVnl3lnoN2KOO2kkexDkKi3oR9h3qcoxoiyHT/D0kIDd
1p8K4OmxnTDkGSqDUpYUTbArc+jG+8xqjnnHkAn1QibVrVzZdVj/A1M79hbpK4nIFiQILJ4zaXhS
PhxM8Fl21sTOOgmCIMfWyqtSfLJod3N/lGHuvkOiRxBUW3k4vw2KgjxclQKhiL+Z429+oUmBcshl
xnaRjjFe1C2E1KaGaai8eD7xA98uA3qR0uG/7N51bZarZJjLXbBvsdeCYXLijMGPomAmeLT9BtqM
fg2su/vm9my1Q+SpdB4bocQvmCEcIiamGlLwQoNan8CQsQA4T7vOX6qu8YYG0t1bpMrplYmBu4fi
fUHtCQg/y0uBh51TTrFbjpLWgB+LqxLN21FCur5b/YMCvzwLwmXbvWTgAp/qmagzcJbG63ew7YyV
bRGgtFuCs/EXhbBD/9Sddts6IwNcNCqdDMGyh26jhZ9rnoQH0UYAcQIlFLZjTGNp+8TupyHEnWOE
5wwD12fUWVtHnnJb5Gxq+qypz1RxiF2CBbpjQ6dkOqcfHgyMYov5kMq+b7rkRrL/10qNDIGHZUlK
c+pP/ciwTok0uY6bVaYNWjUjCZwqn5PccuYz5EXxA0uq0x2VcvK6ASmtl7lBCFYLBjokvNdpQI79
IYBybqMqrhkmVtmxf9tn43AH2e6hvyTfrc2clWJwSl45NTXUZFbRT1Z0jp4MsrqZ2dX14nWQTKpy
XR6lH8N8VaVj76QiPPXBPcfdazREE/Kpq4j5bnarkjkldcjXnEVGUhegGldXob9UZ8b/HY8IVFGJ
TYqI79YyUqv0mcLNYdmI0jJ3hf5/KKE7kqOhZlFJfyR+3W34JWmgtBy/TzcL9/MAT6Lwxrjf6LEf
i2Q8p7AZ7AlAn5hKS76PvcezXHraUdPx9fAacORK7V0MBuzxwj8CbYutp300bJOeSQ6ebthkuRdj
hhkz4TIV+6F9vACqJsBFmUM2elY/gnZO8rFbkN7IGQtwzp+AtBoVMK2tzd6aY6ya4XnVknJ97WSN
LRXeE+3SwYC2e+rCF426UGjr5t6lI5dh3Rjzn09jiBL8qzwXvjtME62Y+pO+4emoHXAqpFDYYNex
Z4xhY2XzGipo701c2OJsBQ55dRQ0x4RAQkAmkdzLUsj81kEP06YNrliqB3bpSLhNc2QXT/3SO44H
ekTDQlagcaPOHCwekqhB0sJif6oAQy9H9Lh1wSgeM8DssgZ7aUa7vNKqAPYZEmAzqT9DITHeRqIh
v2cApoTv+n3DMhLpe1rt1AHlxQZ+SZHorEryt8LNvJmwwZggfPe520szlo40qZvtJH40APYYPXKn
KlEXrA10rdH/vMiCbXBzAardK9/bazbJYXaMV21jqKYm0bLZtmO7o3DeR2gqL2TXUujgEEQiKKhP
0hLqhXmFGarz9IG6WfyhfFnLXvYkdMx8crXfrQVU9lXsHrKbLHXjra6ouvzMik/hIe6xeP2JlnJc
LPqy0CM9+it7WDSbNKtWSADbx1UXQSEZ5cNf7/f2bT33vSLktKAtX4xvvqsbV8ZGlfGiYbiC4Kac
1PWCtIUB+C+FS4zh6DiZWR3VIpRPhtiV+HuIaXngMV8FPF+3hWD/mxNxWJg9FNHsyXAvU5SrmkHA
CLizZyoOtIXhhXlXMHtjrUlqsGT8vQ0wG9Li0O8fZz2UNfqn6Rt8wR+WEpxH0A/BhWLgP6FrP4uU
JWse46s5WUGnkcrTFgfyPgI7O8VlquvIMcV+AVDVFfgTwPC2Vtar4T8rvxi8hqMh4zNvA3FktxM2
S7Z+bKjofZqyAEMLuvmtZBCDJKX/LncHg6NTR+8BBRKgWie8LtHyid3stqj5Pv3U7U9YLX+jFQq7
lOZYybEUK6G1y/ELHw8ih74hXdFlsd4O/cNGQ2bxJJGmS6/MfotmyxKF92Z24qk7Un0Zv5lYQTjw
flJy8KbgWQ/EwvYa0J592Au3RMbBDeRG7T8ZuqC5MF3rlxzOKvsh2amuwrtwdZjTqAZ2MoQmINF7
kkMGlHyem34JvJJJBAJ4eL/wITq3U9urySGaRA0tH4IKLLrioN32Afa2cw7G5j1KAx0bpXCwHHgL
jVbVLPPJ0rywGgwco36nYjChiK5C+J0rfI94xcfy5NiPU70OykMJcRxVusbRMrUCCh5IAgquhhiD
Swj//oODaE4BlEjWYrVRFkqhc2OOosG1McnJUMDdjbdZFrmWsBQ0psJzVunXUCcAYvwYd0I9wr1D
gk3PglOGD53qI9yZb2RnD6j8xN0auBxfpZvMJrpOoIybiKodL1KFYBxZJONSwGb5FJA8I5MS95c8
TaZqsvLjcf/ox/QnCBAjYqbDnYkjkt6/D7f8lRtc2LguSkRarBCBc5o31rJTV/EUQLvVEc48ZUJ9
ENIJ+rTnqj2V5FpuO8o7uFJAZTY10gHKZKNkaHafDM+LiwtjCoYN5MygxvbBTfXqeSN11qpRRXLl
0lcTW153s1FguKhoqQN/e3fQwf+5fLd8kheXYd0eFnljI94g6DD5EEW+O9/BsHC2bDrjGyx+q+Eo
hpLo4xDW4q3pQBrumyGEzwb/usUJmCagYKk3JGiIfkP2wtZwEWFRaMErv55yEU5mH7yNh1Ce/TFG
6gRwikIlMa3O4eG7ZYGDk3SbDKRdZqKpcM+jcPHopTTzLDf6yusq7Qy9Fiv0mW+7GeDwX0FF3p9t
XtU4VNj9l4nU9RiRpYu42cWK66z84pwtFcAW5g/k7/OJ4mrFo/W4e1p+4csgaesMt9TM4rVhshIo
ALGA3y682ybLsmIkVxOT86gMrdHT/SNmaCJt2q+0vQxNscb5u35KAnsjoPSrZUzJnFp3Hq6xV44E
5h1lR91ZsGk9s5asX5h4c42hAc2z0hqn50yQ3BoMdOrslLOiY3FvaZ0nfxg1dErU+FMCWBon3g1J
VQ5H9yHU/tNyE0+UFcZutyDO0bdrBWTqry+wkIeFJkAVNh/NpuS1XOs7CQTUfNrM9ieSHUK6LOPl
TaBvgDdKP4ehMNLjf3k20GKg+lcSRzxU53VqFJDmJoYtqn/2PRUek4H+kbbYKHQU/AzF2W81lR3D
29DfYPczc+UD8JPWf6G/1H+6b8zr4/abha3Envku4nCuVx9jD0egKfY5K+7W4Sd9Qo/Oq8hqNz7g
4QPvEzwHcO4wt+FYwSOanBaQhdpucAj5aI2PfShEqFnBvXZ+c3V4QTogEJIiGETb+VU232JjjpTf
eNAvLzFPMNY1akACEm/HbeZLZk1pxjSeRaASEyWPZeGfXeTwStt3AvMqBkseo5UVc3Y12+jnpoWc
wvvrQ8R5dOB1URUDovdNnf+CZp5MDeE+fSqocj3t0g1kX+/r28Lny2hOcnN6dH/Adkj9pb9GIvv5
fNhvkHdQqXn3d8PHCKZej+rI0oav7Nfom/F0tPJtDFG3/0+i0dS62XlwlXfpXcZCPFMaYnIkcTIx
BWEt4JCfob3kgvIgp2EEm59mx5a6Huy1z3lPtfsAsihRru7vKl9tDM2XBZQRh5h6xfxQgw3vaE4R
6XqUv2RqAQefXInF4cMInMFZ520f2jVhsnT5wOSUmNSZtGedxJXMTIqFyZhenB0BZf3dDi8ooOZ1
ckhnW+/lS5eymGZRIHoZiTWa/1P1QhfsZb1xnRZmhCjFMdOsUGBu5jBfINBsKcXIvgUIwtpDidj1
5hUnyE8EY0FKP9e1dZmCRLTJE2AHVvelBPKwErVvV3YrNAXUWOg2VUC8rj+WpkKm073BuNnjZiLL
LK/bdhyf1R94TIcdeYdN/IWHURjuarqqf+CS9CQkfHK0z8iCy3UpUAL3uomnej+5PfRm89OtqJ7o
U43n6oKBmey6qFviLDcDHvvfBmjwXHIQu03UUs8c8YmqfnZmo8+j5T1pB4qE/1GfkL28YSy1LiIm
ZVGehTi6MVVahgFvZmsm0eE21GP5ZJA8COVtF8f/wPMUZEjL5Vd19rUYdix4YBqDW5gZjRadguTG
Z9jVRucfOPXENOx/my4WHu9g2k037rMplToLa2jNbiJ9OQvmwYkRWh/qfLaoqVyMPPHBtpWDgYew
MfC4sspneL9q3ntome3ta/BZ8EiAkru9TnE0WtwOciX0YMxNIPkHFS7L837czFRBLj1qXQqNuXoI
qkT5KByXa21ld5jYDntfAMe6ZmTNZCpo9kbc5M+U6CbiFLyxKBGd6obEKe4SXBHSt+Yp6acWGzbb
/FjULVFP1pNcRlhTSh4//8LzPrtjk17IJ4J3ajKppb2btsr6GLb6Zwcd6J/HAZP3immSixjR45SA
UEElJE4csmgLOpud0JLWBl+45ckWKunQnQmZSEi5HNigxhAVZDVeR6FnPRVNk6nR34W/8T5q+81V
a0ziNfGUU+K5TceWfJLE6myXg2vrWEnvVEDa43DDbR6VMziBPbfXsyLcLuzgbRl8EGH/lHIuMXTB
Vcm4ozUpyjxS1/cel3osHU2YWWL092RvAiB4NfTa7BjC2aHcAY2R1+HvTRAXZsi+cfZpcwKpzjET
4oP9OoezLZTxfgXn25CgTXPlpafTt+n4SCYKNUSGbBr5AQBPen/BIjJBkcrjgN86FdiZ8+0NeWyX
YbrghsCkBJ/jN1txXgRK5qVrYqumHQFkzXWKEaTG6UFBHwrOPDixsuaOiIfy86Pr3LojCNhwwkt9
fOsnXQec58sKAmBf2P/K9m5jtkAviOPBhmaUN+Yk97/OdmSAIjtUgam41Rl8Ettbq9R8jtGqrMq7
GAKSP9MTjfv/KYem0EuVD/zDNOMlUtl/rLCtsxD0WELF/TF2nCT50IN4YA3VXqIlux2rLfDY3zVM
AA+JSLPQlMZLI+sZmC6zVbAM/lM7au76XrQG8WZk/808+ZhI2NdOn9+6Qk9ETliGfpNOdghDdapt
yoxjNgDjcqMyG9e09BZNvayu7TaQ2I5njWD1qnzL4E925gXRbxlFJiBaCZmPbfHYigLX5osZpXW1
qooxh0/xi+Lggfj9fc09GAg+eqM/Pw9WMcWgJzPa401LUt2zVK7a/oq9Cm527xNTINs/SOKzW0wy
/0qsa6QVdL73vm5vKy8qM5i4Tz3ZLFDFNZEocTb+elIhYu+6SozAHeaBo37l9LNtB+nd1Gg0SAmM
pPHz1D+Iqnc75hvof7gG/BZVbTpRi6n84lKY387gbfPI4N+wJnSkkRhWUtW4kwBVLLWXuniRsYM4
g///SC8cs6bREcPWOr4xtm2EKhOReAJyVXNAl5vBUPvaAutGDymGf0IncXYn6TqoqUtc2r+aRe+l
gRZ/vKStrXRrh67tBvw4uPR/TcEMKZIbySRs9kHtLAiHq6A09CJYMFiLXpIDUNhwIp2rVyPArGBq
ft46dqtkn950zriL+NHrpK3/v6rJnYdl3ch0KjY5vr54pVecrLn6PV49Sah+qtqB8p1K7dECzjIm
/QguNK1vpeosuro3/zOwJSUX26iyqatJVycGBSrCjDEcANAzS5beUsCwpewI+cLKsd97DbJcoYf8
RbrodKu5r15CTSh3ZvU794tvJr7+uP1qU+v0vhS4rzBL3NXRhpOcZgrDTa0M/Kk/OHMAVLeb+sxU
Oj6vWqt7p3IW7Z3HUH9rng7/tPTUP6ZDp4HAn/XhrfOSt1EYF4fHbzs5AzAi5lGHLIakB+mUH62E
DSqsYIKAYlIBXRjElu3bXVc7dWzzuJaeE+V5FtnttoCRSojUbSd+bTINjrWyJaS4mNLOLQHjAm9v
feHwcFLbte9lJfN3CXjmSGgg2FieLmGlns1fSSg1i1ps7+1dh/aX8tVIltpgl98DBSt3OLbCQ02B
gcubBKBQ/XqpcLpMUW53wFSYbYcpqZodJTMxQyMpZwBcdgUnbG5lBTBsIWt7g00lK61G9A1BtnR8
l8CVZ0igM4nUhDuSfNQQQbJ3F/K6UCH7ITFVyaC/HFEtDLA75REVj4FpGU3gDFnRQOMkRDO4wE3c
J9Xtpxx0781+e57Hk9yiTLguA+qvXChpEQzxAYv1048oktx5uZF1iTx5D4ItvSlUcT/rF6sAiDdv
h6Wul2yj3vKsiUMnHR47R6RRfChbCLhIQ/5/fhkegtFTjwMAR5ZvxU5NM2GdXBBDP5DFXy/Se81N
4zq4Ws6zHhFKtelwcisPhNLfM06BQpK8c0pV6ND0sd0fPSFTevON4gpKMT4dRw7z/1mM7IeAS8Sz
mePpi4XG9OjU0J+sFwQp5UUtjYQzBXo6W5OHPxD67uETUZFPQMEUkfTSEVHEadTkZwtNCDxIIqXA
IS/BltQoieCx3dwxcmVygjmdFYWilYBhkMlVv7lGCA4xbgNAptVADWJB76WcoQ5WiYRL8tpUQlbt
3p4u5hAUqKrFl+k91+ZfdduLa+foa7BmEGMimSAn2FouPBPmVvWPZNWCnDuXMF3m2PyBpBQzVCK/
8NsrhkDKD+k+i8NwQGr9pxo7L5b9tc/8znNOygop8iVvyqW6PzWR507SzstlvIAqIErKYTaMkoG7
jmPQfLd+kUcGI5spzsn2UzgpEXvg2zjahnf8vwrdTiYEKqOoNYkAw12BGGj3QrxOqQGAcBJkriCk
wqG4BbrMeeibidHW3+mIcCb3OWgpamt0YNQr3UsiYVrVAuydN0U8ZYLVGCb7XuKV1tJLaXrC8l3U
WPcLc1C1oApk92T2TocFp05wj4IWZdymTUbunjbtVz7dg4vYLnKVLdO/+0E5LWZjLGt3VOZ40h+z
h4/4S3cQ1BqNfK1a26mvgRhiacPgOwCQFBFaXod2TfvAk60Ten0Q2OxU0e4RPJZtJecFZefnJ8It
RyVXeqkLnEvfPq4AAlIe5DLaUk1Bv7nHfrZ244M5yFhCg2d335RHmdY9IT3lzCCzTgxVWQXV87QX
HMH4aVtYLOL239dkdaSLkAVOPdXXPKfOT7DJDIu1OzV/Mq28IfScmPZVotsNMaTR99Sy5OdyALUm
lM+9ackyOR20LPzCN8sU9EeS+apRnFBzOh0guMsPat7yrVomgRUZFBNE6qes8V9zfMgAtmVx3wBw
HI/5pz6gxWWIW2kFF333e26iM+6jM5ukH7nzDt47nJIFFjaeZ/YsmomgkVnaaFzgROO8xflL3JnU
QH8uE/Wa1EqqLjrmJjhoPyZHvw+d1gWwa57SV73r8sckxEQ2Dc6nBj/aPsBWEBRv3aj9tKTOmzeK
T5KXd3mCcZYuT4FTujV5Mbdl9/WKQwFUXfhUf5toOhb4AxTTJXf+wOPeDUWEfhUyRJCTQevTHcEs
6CooEvjTXXNykEw4fk8hChVtzE74AyMkLTPsD10RVoeUIy2JPR0IM8Xgmcv+cs9BMGKkKPtoV2PM
qAMOX0v1/fOHU4VrVFtVisjFXpt22iiq03h8BqtwhyTme8Gin8anjrJmh18lJfTIX+wMsFxbg6Fh
kDiI2TNMOyrCkEUHQd45FEyzWvX4Q77BqeOY7GM2bUe7t5JOeVTbHj2cLpISm0jPXhFMgshHDCiU
8o/DOQbyH8rP+e/ub/7hWyYqaqJ3IpoTRh4cFF6udRPJ2AaP8w2gFQRWecSb+MqKScQii9ouJEIc
Q7eckdEzsKhTdCqYR9ktEev4p6eRB5j5U/EVVc7L0jclFtSzLddXuF0WWlnUcsnhPUvAf+Y9ZdeD
jdiNMwZqMEBc/h8tcfsETE3ycIHEtWRv95hDY34CLQIlz+n/0N1XD5W1lbbd8MhJOtQ5Y9rXPKBh
pbdmlTtTy2xQHN2YTgY36LfqN6wvzbjxhLUmpsKoqIGndI/l1L9VzVsXbmFP1ZjHH0P0mcVcTnXO
ugglH/s19uJApPjkmoz2CC6Cy0oQAiHk0e2hO2zVGqMnF0XizsOChjGQupaaEcOkZVCqLOH4DeSt
puCs44ZMqA1t+OOKxsfCFznqzTrWNOhN7AQKsU06YReH62MIDE2RvjpSlFSA+Qj1DI9rPrpEhiIq
B7Mo3muluasc15kCFiSYYbrOOe9667ApuwGDx6KDJ6Hgvd4gUlLkMFMIK4PFrcb8QXyBqwAp+LaC
dMLLoU2lp/xcN/cVTMlP7Zon6D9QMfB5WqGei6K5I1WFgAHBUd7DRnnktKynJsO2Qpod/+TeRgp5
m2506QigFYqdl/99UegBRTTAXmeNJO1O4RaFjweTXkG3KWGZxLzjWOPwZpqHN8hacopM/Gha16We
/XhXUbB3D+iZIk9sb4uIryVFdAVeUjU1uifVKwAx36+uxB0owBoriAPRn51oe4WiRVhDDKcxOPH6
mWKb+tr8Rc9bqMTNnLv8lKrWAmagnt58PP9Jj2iY4cpECFXanWYAvwtAE5Wuj5tM1gBy8Lurx4H9
/RGyz72/NiPlY7lO5ktRN+Wk3XvDqzImvCLJnKDZRHgS4ZiBetc1CjdoMTf0jJEZDizNueVGo7PG
hYrBdpauO4EwYdD27o36n5+NjYXyD2lpq29EX9fV0b8FBN3KPcEg6VlDedhSrN2vCcsb5tZd47jK
sgzrCgekDPVBMPtCcG/3PZ0hHtv7l34AsD7sEaQb1qvJnKREYswjmMvQxCYz0WFRMv3qeeVGaQfj
alNbf5RXxonj3nbIPQc3/MFZGoiMrSCQnP+6JOvs26MdRVQPERdt41W9rfS8gIwGHqVNkPmGbDFp
KUwNPBPYn2LacKwdMLjtuWTMmh6RRiiyo7z3rmqcg6iKWEWJ1l5zsYot/sWFCyeQT87POvOrKi9q
prtF1F0HTqITgXn6FvIh8yPdxry8xIWQzos7r5jzfyDXY35kO9EQwIOhuxo4sDw5ZPhBzScyVQ/K
yP7pV1k+78mpt4Va1DMm7eY5pKmm+Qt7fU/TI/y74d5Ju5+k218fpl90ylJhPW1/H5SA6wVfFIKj
mTczagDpCgRQaww7Q2cMo0D4jpxTkCvDBRaGNM0hRVy5NQid6WecS9JtC6ejM5mTanSo2dl9WHuY
GoeLUewEBO9Z4UHAXH/h6XT8CcHmXXrZq7fjXC+KditovDASyMbH3cFYiBEhPiR9Fa6QQL6YRFgt
MDdatUOAfjGSdl4EXyQ1n1KVH4Pkz2cT1nZAEOvWRIN9keZVCBLsHDbe1Lnu0ZK3D0vIavTpms/+
tWDGKYhowmy1ITwOY2xPWofDN9V+7B5GgMaAZsIS48f41QwHwHobVclLs+StQCiGHw3AJ68rD32k
+1N34ReJaoUnBp7Eoc1RLae8RPApI/Cf7erhA8N6Mk6E6ujlMQaGxZMSNVgEsyHxQH45Xhngu5qZ
W8/eow==
`protect end_protected
