-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UE9OOjsCLB/vbP8qPODacUcwEziqVfPYqbj0HluOg353isxtOheZ0GGvmvahVdxH6uFHUh1gqFTl
F6aRIJx+LFvhqCMlIynW3hiXlL965n5X7HJDskNxK9OsRryhrKK4pAsMCNRHm63tkI71KQpQyO6k
y+rKAmCj0pmwjqTX+e+y+kPaBZfc69f2mtIFwjpOOh+uVpoJrDN21lJd4DaRMD/iakTTu/VNPWs7
xuPoAnNmCqIjSGMFAbajowcRhPj+89GtpaY0rXLIfuwWwu+2vIloOhfOWlGoYqmjpGP1qfEwNpti
RbVh+CU0SlQkahv3B9TXRDDkTP8k/qSZCFm4Mg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12400)
`protect data_block
FAdP7qY6hR+bNtYd/FbSzgNkLg266mR4B1s/21pBMOcSC6DQiV55mgzVDKUcFqaLr7LpjY0sz0Gw
C0vLcRJmZsd9rsyVf08IQJUh1SPVIr6LP5eA6ae3U8tH/FG5wsi29o9Mytu/ur1P+bbt2MI4GVUR
lyI12MkkZZ7nFhSv/umegEtn/KGsRXRmDtFHGkWN9yAHl9ky2/MGBOHYiQJwDdsiInUgjHh7hBZX
F1LARbOrPtI2ERj4/aHzhugiNuPF/62s/u41nJjNI2uEUEtzoQFOaXN6GRfrah2bo4WhV1VjAxnl
rYJkE1TatF05PSI80M/37Xbh5f3VcYCYX+ttOqwO9SnOBZbx4aC+zhHvoxGPnwqSgdZDSZ1Vai1O
A2WrExQ42CZG+nGRYJKNS403u38asKAgNu8ucJRSD/Wva9aOLyxBWAmHXDGU5bc2fKVrw1E9eBr+
yjxVIHowZhlrvt0qjOchwxQAnvkkGpZdRF0S1nXUNnSPs1b93U0nYQnd/EFescuhLnlWTET4lR09
/EEC0zbeqbETGCVhRs8oKosozp9M5f6niD+GZeWbwK+I1l/z23mwMd32ibveiRUSA77uQxXa+0J8
1vT2EeDUfccdsHbiG2qD09py7DIlpPLJPDKI47gApue31UxLc/gDDizfPJ4e9twc0pG3aG5EfHI0
dhmGcxGK2EgIefvPaTcJcV3etCiMM7aj/HJlBV7QRtPulh64xr4gVsvga8DEaNSSvXL8EnU4gXKH
g7RXA8ygUoXxRvrnSlwihRFziHbQq7S4kznbZ2fnekv/xxKmU5hTlIAJlbXIstZkmQkNYWuVncnc
fOHpMRXzVNj6LNyWcsosyFE+NaKY/nk/pjhbupttJI12XQV0GraxZ7q0Bm4RpaQX2UYYhnQV696V
Nv8gR7Z7Mor1V0xuGrOC4Zs79M6ASw/tWYaKefJo4ltFEVEmDrGNrwnv8+q4iL/eUuPu7clNqNAv
zAouabqDjmTChurBKE2EdNH4EQzwYzLH+oWSalR9EWu4O6dIb3xBRr6Fg60+mL11FhJZngjKcw/4
pzcFR2Dcrd6IozNlEM8OjXDjyfyXSCArvJZLcUTj5G9TUxi/rTosw6AeR8T4X3AUjUI1OX3VWcMQ
flqMJxf8J0K9gze/O8aX07ApoFFSObnG9allvWFd1ynPl0ZE7eFqfgbGrAVp5SR9A1n0X7+ajGAa
Ewr7ZVqoTzBt4NiyUyQa6gQVbFIT9wyBjHiPK0160wrpHi6D8atUG7ZhnflNCOUId699bdDEFVh5
SblikOV9F3vhGlc7UX/4lukVJlYRTXnoY2uxOFn4Qhe2SETIo1MeCqckddGq6Ek6eODLPey5bLWF
vmPUWmkDDwtgvv8AuczL3eSL8uJkx6VFBZy+JY5DRwM8St6nYPL/l2QdddF/FejKMHA3TDshzhS6
vIK5ccy6XZnnYsl8HJe9FLbMzczXUfv96TuO75n3/v6t8iMly3YXBt+2Z3mE+Vm2OZNYEbJaK1rw
Qe5XdiyXPa6wbpN/mZrVMqKuqGQl2FQJGgHOPepJQOWoNjvKnaEJr0fGb7EX9IROEwizgc07k48T
cwCgBfDF+S4eXqu1fW2KHIJz8uBXcURn7YG6UXwGTxyIFsdqqeATyjZqmRSUv+bL/fPo96AMAKLu
ziosJwcZZV/652tEKhiv+chf+GwqjAYyDjKg81iLLYaU4nUxda9QKVdEAZ9xKyXFplS3ivOvlQz7
rwJVBMpxXgj7gGy/sY5KnFWGPdPbYXxSdSePVToGqPe0BLljlkZ+mVgyVnsOvIUnFJkwxXx2jZub
eLts5n3/vLApJJx4nqFwFm23yhuRzeTvF3gWlCttcFRDIpoYSahMZ8+/zpY6+ew5zJ0JeckRFEY/
Esp2BS+2InO2pESVEL+pzbKJC0XLqZv31s2aGJaX+y+tCJ4JhdeulI3Xy5smYC2ug1YD54V+5wPl
cil61nQGBm4MSZxz17YKEIHlRAL4WjmQ50B5ze2mj3QtBRc5/WWmswgqxm49P9y/4iHmpK2baNyB
2FzJ0o7824fIXwj7ZNSVV57uuAapMy7GPNXEYS5RvlaCApnvzNCMNhExea5PwxMstRhbq1BSmlR4
EQ15oTAy7ot16pOiraGa702N7gIXn0q/HRoyGXoGj33lnwx110qPgajsZ0nLmuxMIPmFHHT4RJm7
4GZBegA3BRGD86xT0VvZ2FU0R2D5gTLF2oL4zksEKClABth+yePS36T0KhUr1s0ZPhmRP9o5yB5C
IqlqsQB3D/Y0fPBHEBnoniIwCi6mdxdM9LzYsSWUhtxBxfJlwDiiVgyRZBYzFx25hle0DLyJOchZ
3R6bv3vdImOJ42fga+hqg2tVOnaR4AJzAbGfymX1YbVh1e6kJ4ubNRgITLbajRjwdVE2E51IkCIS
WagaTnuNX8riZEpqmYxVInCEJu+iOHOEEe9AtW7O8P6e93reNdA5TE/zgdibVj9i+Uj/qeTMv2y7
0NW64b00COjhPQhVYq5s69dGyqIOK6wEo3pNsnZSo1dCH6diU+HVHO+AZn9t5+6VhsOOUSR7RYmP
rChWhmQsy0E2jztQd8IEVmdxfN6Oms3NCaIpv3iOMbXPuqjumai1H4neRP3g6XeUCYeClc9U1dS2
/kmPWGxFgOrTMcvStliMZNCFbU9zvD23BDiIm30oR00Km7gOhiy5Q6vNnQleQk1qmsjJrBNI7xBl
wcxXTx0c1U0b8dRlraXay9kzIx1dRaFN2lR9DFMYKIQuE87fEMbwir7Hl7uABMhHxKM4mDf8hb6K
ow+VjKiSbqdlUwYgHesqnWOsTIfDN/RxJzSaoursJGNvrAwM1IXTlKMFdAi+a9Piz7Ark0pGy4zv
qp9Eu8pxbiZytGANdAR0NHTVeIH2R63Q7yqnKWBFhGBiIuL85uB3XcfmLOOt2XAWmSU+IoneYIOl
XFzYML6aEhBYgQUHhgTvzhLLfbBDQdZXwo0+CW6O5TziUaR+zUlMQShigswHZ5DYqf/DqM7nZSnM
T8UPTSJyennV8C6wsnVoDrLLueE4cDk1jYw+bucDvu4NhnhpWSK4sidJ3qws9Dtzf1ac+DzEAnK3
EnG/pDMV3b6NKF+Jlj9uT8UCOEnpQWpDm+a+CDwJB3e0Spn1uUSvZIh676/dFd0QZpcKjl6KSsqh
ftQ2mmDEtLIcpBqkQqz1UY69bNOt1P+xfjKIVV7aA9eqL0+CINdwudNrWcWp+HrqtjdbPLeGutMW
Ym8kjkE4QWzW84XhzQOli7QGBaDPHbnSCaYa9V4kddGACGdnPmuF2GhA2Mk/oTcZmJde0r7mj+BE
qNzuL1t+JgoisNrcgeUw6sglNdMnKW8D2tPZ1adCjzgP3D0jlOaeRl5Sdp4eF/28zuvV2PrswStS
HqCjDaWoNBcHXFWXn1BsRdBsuVWdh6n5q0HYeAeWCXh+wrFq2pV1cfOPIgElygYV3t53X8p84eYD
lgZPLTijVLe9OvzVjGsNMA5Gq74Qf140L5banfkI8OPQD5IStiCCSpxemEaEYff0osmJ3+l4fWee
6VpHPz3jrZPZnG8dMU3m4fhcdh036a3OunAavEGnp+CFjNfim8sY7KbnLth2iiRg7AV8Mkq7qEEG
NEGK+QNzEiwa5PpKDSTfVoUXERMoPRwsgWv5LZMzTDBxJmm0cUtuKSPUdFJMkimdnhGw4mMV3j96
oiq5mOoWJ7uv4RcqiXcZoQC7EH3bOAyh4Fhs9X1VXSmD0NdSO0KWpISAzdfRFmwqofyFfg4oAvig
QbC+eJTA5Uul3E5lWtKGANvXMU+1n3DIQDuT1Tm7iBlcsgLQ5gkh/yNicjZBK06wZ2RNpI7bNOgT
AVuIcSRO9lEJKL3mqQj2A9bn3IpLhUTq0LphWolNj3UTMtNf3avelMLH5golMTGMOMWDePWaUAno
2S/AtvQ7OvZRDWwaHV4yAYMa1YbSndy4oFMyU79aAwPgOGod2wzy+IJrYqyjOp9iXW9V09HynyXm
n5NFc5EsXxKfeLM/bzVZ7CL4VCzh7TEEVlNSlmfQv0v+V9/PGpDUU3HQz0QAul1R2d+55seGgIIk
Wg/7GA6nOGF3CeJU7Oh1mc4nkhMbWbZcGeDuVJBQdwK+4KBwn/347298fhVerIPTx412RuhrGHTi
Bi+851/TkuY+0KInxZVJ/EKIrDx4nGQOaDJTT6HA/Mrep+XS37wMAKT2p7AngsvKPInGYxPlKLEh
zC6sgVr3XebtnlUNBFM/fziTCHkpXE6o8/llybFX7PTfeIDM+oaNJh+Ho+eY5fNCQA71FDxOk3/W
jDXpbWJIi6GEqUZqahfu+f5SkdK6+UVXCwRyjd0RWo7LRbS8LsI5frsda2tcNVJE+lH92G87GWln
xEm/D5qzYywsU+SOaFWYR7b6sJXMjzeFOzH1hTA60cfhjoiry8JztHiCGm1m1ZjdLfA3dsu3z0W7
jHyV+94BNJQJQy44IyOQAVzcz73i8ImoCynyP9Ftk04nW0xR5LYBIS3PVV75rFUr/JW5pyQf2I0T
j/0/LyeLeg1ZzmnckPPn5bl6pyFQbVWX0f0Cjt8ptSufsg9sME7vXqxPB14Ep1zOKNQSjo1Wxx6P
kBhgUaNwV3+wZD5uGO2+mqCZfMbJQt+LMn0ypjaj8Uh8p1cjGrrgxJF9iYTuFYUbH3WTiFlgE0p7
Msl8xb8kxlhFxxVJNrM0Z0sQdX1CwTKCgX5kodWnzp1i9y9w22bsTF9Pevjj9Nrgz6/zqi5XiOOj
YMfG/fXm0Y/Fz2KGIGli1i3V7JzZIJz4b3CirPB+IezIfuu/b2CNZ3qdeAHf70tlRW/imVeEmNkP
h4kH2HvXZvSshnUrHRwVnPvwbxfWnPPWjpOR0ACn0oSYg2kmSIoH1maZAEtF3NNlL6W93d7p5EnW
W7CeB2c7s5DdBu6XHSEwOwGhSmAAoUDAaQoLKq3sd1lT6+1M+mm4antebs8d8QXeoIN/sI4IThtS
LZiO1qPrvLHteFk970plOkTom4DmK842Vb3Dx7ci4SzpGCbvsyCnHrsbvj+Q5gt3Y5IeoB2ER3Zq
TjNMaEZcwS40/o1BpeT5JYZtTX9T3mkAhnfU689v+UzzpjOVAmE1oiUiMMOfwC+BrUQSu6ut/qgv
hUvYrPp0xcIuUr4AOI2O73SGPEdYL5e7i8A6oKaGVps7Dx3Ex8xyH+5WBU0KsLsvjoyHslRJsdHK
hYjWQ3HVKjoaEoTHxiN01ENfw46YYkhFcf/pZfBLGT8Us7byEpyE6/sUs+52cFmGVrmSasKAgzYr
EbcsohBjxy3BUogv2Z9w6Fmlf5p3dgR9lhs0inCk2D2NGRO7w3myCbIX/j1soXFs15Zgmw1fxulu
k1Zxgsul8wImGjJGPsNPCSNtREdp3qap5xg8OH/Fs+l03KoWXDZs3t4dcZ47vhmjwloGp2gcWtHN
rphyNA0IA2qTMtyutSgV2jdrK1jJewhUURMDVL4ZtjpPXv63rWjqrRzdvuKw/1jRVfx2v/RUQUlx
V766YOTbn5qm3YzxRzdP9AohUkq35rxDDdpW0qdDJCQz5RJaOPeFweS7f0y7ZAXa6wdcCfrgKNcg
/t2978vmO8+bRcN9xRStWTQMS6JqbfDx8Ch59BGIZH0CHOnEJ0RGlwdmHNprCj7IriGiWhaRM+je
suPF99U9r335X3hUVxku8EV3anpt1MTIEEPlfdiDtiUeYunte56+HqSBLlC4pspyZYbog79nl/0M
GklVot/Nb81slB4PwL1SqWOkqLDUjwE4Fw75x3JWxSNVFofaiXC8gdDjsucrEuDyJ8NN44WRrBWM
BP+cYal+32+/mHCJ5ZK7IKQlYnqXB/x5HjimfqpEbt0DUTUOP41OJGOJmoNMFNuV6qYiG/QCeUnj
rzPFuczX1PeOeRZcCPxgEeoomg4Pq98Sh0nWOcL5BNpp1C/cGgnbJGP2mP5U6koqN9H83iHkZvh6
8guXFKyVToeuq5ODxQFtnoWpleRlM12ZmERPPAz5ZHq0C1vf0Xad1R/IyizniWIrK/0AC/owzRa8
g+zjkolJmsJsqu80tKWAr0X01U0TozK3aN9f9JtHn+jAGq/s8xjL5kpRjBwizmt6a+juqSkZ4fNn
ITYEqp4gVK6JlW9aWVC6274b3paYFTePl5quPkeME1JVdjG3lekTMZjWFzg3yjtc5p3jr6Zj0k2Q
nZ3WstyjzqSu82Yql2zK5eo3DO+okyEH73kVmiW+bfx9wpZpDJNxl6DmlxWeHGMd6swoP3oum54D
HJfTmjrnyiSdDM95vEftYhbjjPIB9fJfmFrDxt5jfYo2NXJ1y1ju6Qft3Bpe5SVuvFy/3W39wOom
mF0uvj7TBlBAondRhYRclG4HrTzriiDhPEHMMn9lg3x5oEYAiJMwB6qn/C+aLzEBAixVpB3dK3Sp
5TacCPGV7zxlRZhyZMgZKy3d9FfrUBpZKEfdpLDRs5M1olVOIOWe7O6XUsfM/W4iIjeoV9/V7S4w
WPUPjVK6Xq+Wa+RWybrjFlbUme5H/s4mCwCuVnzsnkqnDgMkCtHMbyFOym4Epn3uPlWIMqKbnjuR
PvTZRaiCMPaaZsQyxxvsXQFnIPwBUQ3WtpD5qolwoaaWPq4TaloANyk1FrRjYd7tcy98W6Vq33pz
OtxUYAG3oy80+2OuEJxZnvxE9put9zdSZTbstJg8w2O7Qe0P+RUwV2zSSJeLFN1Zzmfhf8oJJxXg
wPyRD8Ku6j2mApRyauJTSO70/Mfc+6/N0idCJ35Q9slyCyU7VU6/o77+zsnofDu1iF/WOHdXQxpt
Bk8LvpPUno0SvWRcqe0QdM1xgIFx8TniGvWsNkKKhQElQmXM2jz0NwVCrlwnhhs15SPPVJpPCq6L
r4SLA35HwbA/7wKNgXa3HT/jtQmyXBSD7VbIwjby3JB4s+jdtQ76D0ERhH5cf0o7js290ZYJ6Uaf
pKTvTgjux3XjwLByLMzLkFSetkcBw8MVf73sh/6TaIrUvniC3Z5nXEVU6V1Jm1aZZwqYwcecvcQU
2VZgDw1W1OXEPaRTXOJvDi4gbhBNWQyOYq+ZoHtDtAjSJAApdNfqwTcjJiFybWvl35de+Lajav4S
WMUGI6iTVe+m+VocRr/S5IDgy5wV/cPgLl7ieaYTGLYyESVKgrcJ/uQ0VbH76V+nzqtb0Z3N14Vb
amQrCaHM9nPcCYoN3OwrMx2sjapv78vhSnqQeNCZvFMPfj0a6VoaqddIPCp0VNpj8mBY/N/vkgMm
JnwIEyVurzOXYRtdsarb5BlfEDyElIDRfuKj6IzAYZz3AbTArN0jHQEra8Choz8JlD0ztGOsj9Eg
nOI/dXDe0PMm0wrDfprnuZj9BJ2v0dM7+mf0Uaw2phkKuNan37QDW64fY+0gKWDYIy3wztkFOPc6
LX5Z3SpWOkxYD+An6KC6qiS+zQJtxa7QFbpay/Wf8jCS1QGDfYwiMtM15oZF+N3FNim3EsZUs7Su
EoE+eSh+xxRV532PifTzhAfyE85JrD6M/j8ii54YUfvuxM6arrSMwOc7YhLBTF/u2GCzrf6YWdA+
OgxPGiT3gQ9Y7Ucg+Rx8fBOAYAC+7C/t9LqsjbDJKSMGW1ZRajOeIN4++eLig0GmuRAsoXNF2dRX
JZLWjaNto++1+1FLiM9aU4C8ZmEsXGth6IisTe0+56LE/pz0vdFSfgXHDQfwDCDnIqxhOLA7BMYV
OScZcJ7CQDXlnMDGf77aZ0ner7URfpTy4WZupCY4aKApDnpd/EAd/nO1MWsDDnPqnxBwuqXUnaD8
S+hljLsCZZqOkbr30uLmMtdh/9lX33bGtI71/U+8GCTbIRzspYAw7oCCScJvEr2T4q19bIAeeErE
4sDZ39YdLr0v1BFx4gag0nSjZLWrRQLIJIcgl8WMUxwB28JHJUT+L591sV53+EKxWkh/2D4zmAD5
XSOkOgBrFwP17l9uP2q0/TvHcb62nGeTmr0/m8oxTVxnodntLkW8agOme7VQVZCV/ov3s93Sdf6w
Od/F9GRvrivzLXBJpYxXdva0ZcKDSJisF2lZuc7KOU+DR+LlLvutlALeZWdGPtfgv9Vq3NCRCLmI
Um4I5b443XYZNHYW29pn5xGzIcGlXWbsC4sgeaNhC440wwlsr5xbSy5yeVQpSjovADGVw1CwHHBj
CTNSB1/jg7yBqWn7/CrTvqgPOPu3ohtpc5mXogkfsQZp3/c6hykjZfym5F3EvODhuty59huipLGI
SiwsCZoXtrPoN56D9pb9frn8S1rggBePdLwCDy56RJMt3IabO1mUvmNS7TWeZybfSSVeGm/S+vTV
Hb+RM0iYPWnQQun7pBmeDrU6mEi/bIhmDn32BamVxll9/MEz6nic5X0AKGphQsRQeoU4YMEMBbmt
bqXeBXw8L4GFyiG0IHzs4ShtoNsMeW/XL4tgdEP2+LOLC89x0zG/hfihZr3aixaXFPZs5bzUwcn1
eUMJ5bKdhOg5DRdExP/nKGjsJaWPFKQ4/0IJfVhcLUqmJpimu9AbkaF2B9yFsCgDa1zI0xxKcXgM
xa4KeP3TnAjlMjYvoIQ2db9RU/HCkOdA+YFxtO+5D1vPi4eOvwi18M+xMKzRFUJD45xiQ92EjqlC
lhKfDYaDfWs0IkdBD3D7Qa5BdiHbxrV0GUTnpu6ZPBQLX5W5r83X5srRLYLfTxwyJfIGsQelNX1U
a1i4EkEZubanP0pfGC9UY8UJhNTxeih9jFqxr6BmRT/QQBc+gcZ9y9a2mB5HEx/+hwYUOj7fZhyY
0Q4mnuP/gm744THKyXn+a3GlYzGUDQbRrn88URQAoUXo9wYXBZ4xoL/fjHB54CBXDSUjQhZoM4c7
FEXNZxjjaE5nEi6yTOdxCuEkGDe+FzG9FJCP2fJIJTQWNtbuBrIo73NU5hXN5am/3GUFAPqWn1hn
IOSzcFdWhouhbBX5woUvWnUdyvEIhgH1ocQG2Oz/fC8J00wTgxsnphW8UdR1sv44CvQP3+xIsr3C
YSkcBylgTYJhpGdDwLuKoavqK7G8acYZlKx5gPw+pM9tTpahItLeji3YBiwA4brSmuUol/pS21yz
xjpUnmwzk/m8MchdPuxUDCiM0p0glLUPc7LO5L1kVKsHc8kTVT9VsYtf/sHPFb3o//0S7ERmkbFE
c2Ql/45K+6WkooiQ+/63nXS+1gLu+nVJO5EScTRg5sxOq4DDW0PaOyHujGfE2wSc7JQJ36vhkjDR
+KDr9abA+SCUWX3O4h6ovjtySs+X6VFmb3UFjPcyBRWUbte2fXVROnW5wBp0n4wQGrZfi3OzLCYE
tBZL/WAE3Q/hcP00I4qlrp/XnUDrrxg0tJhUQ2QddPDP8n1wExeEt9DJtUdhdawUVM8O4rUHFzHk
/xrT6Xi0uVEXMbMg+BB9mvXQjrI5dzdUoBzLzYGyN5rOXCaYnirLhFJB+xroeoa9FimN6LgwAhBR
TV9HlZnZh9Fm1dvR7CVV0k6a02OPL+bCQlQvNp45BxwEUfWYme/9zmodZYfD14H1J4XLzZ0an4M/
Yh2Lp+vrmC3SLdsiPaOK2SuFeZCs4PcFrPXLFLitVQCVLtqk9czQk7smBf5y6oSLpGYnS3Q/K1G8
VsqlBq2JWaUPLivUImzIMvGbtDdWxbbzNVCkS64FjmAMGFcx8vslfj4hvS8574K1WcY+rMTqP6ZW
4HP2rOrAXIKZWF9344muj3lN4H0ssx6TD211eDwTzr6gF1ibc2of7BYW9QQgKpPIhLejAxLxWBVP
sTadKWNTWo4lQ9fCz5v7wGhnmNoNoM86xRWh38/Lbm5mCLW1/ZXfs1Jcagsl/bsxo3SrGJ+fuu7i
CWu9EOv+jfIy2Ne7ufYDiFrOrD5un01c73gRV+pmzSZF5Cs3zy39ezeQgp2+MaWjE2MbzSB6dcsu
ZArSvNpw9qFIXoa9AaUewHx17qVQUy5fO4iJ1NMw6aAZsZxYogkVLEpZIKifGuJbBzSWbAc2Zl5A
ECCCn1AT2/d9ZvuOPhTY4kodaNB++qN1ZZOiQSGXmtlphmVK8g7Tx3OULi6TKSi8krjOf7QWB310
qbijQf6is+UPPfsVL1nKhItv3zUY8ezrniGboPFSEYklUuYPG7jvm0qK5qzEHPxUEvV4Te5MZVDR
Ww3CU4Hf1pbrbwT9PR4J9qi8tejfGHAPBAT3vIHf9a3HnFAaFYQOet/PLcpyMtoFt0OgEgfkCZDl
55mmpY0Xf5ACEtYGOn4q7+rAymMsSz7iQ7FRFsZtkibGjyO+beXjISMV8Z+f8zGMAbSVLw7rkIIV
b7Ge6X16CrkpEft/QmyqXZg6It+BHtzuFHqVXMHu5Ii6mlAAdwEtsC5xL4zmgNGUbqopVU2lsjBf
XJ6vSdqoac0Z7sqrSLhgEOFxzBu6o6I2TFjTCxJRYKHdYIibNVPxw3QeIGD42/VkQfO8Kv+SzMkb
GltW3EiEkLKs8v0aHil2Yrvx6xYZKb9srWx3nzyqS0sI0FJ3qQ5Tw2IAQ/uqRRjJLTOd3a4fK9FU
E9lbjBda8X4fa4zPDbyQLCFqRwolPEH4Z31pe5oTF1Ro60XMxUcMYxtx/QeOrWw84fTcFMeADq0M
AtmLF7ftFTwky1HbxFwUwpAtaeTxL4pnNVqMOLfRnBR4FQ5TZPsor6vUMHARJ95pG2wed++WrAQd
18dF39kOR4z29mXS5WHPNf8CK2iQ/X3x1padpwD7H0sdhjxhWbB0nS99kYcldZoed+m4xnC6oJfl
LhYot4pI1P3fDPquTB+OIHIljbnoFkugr8jmczMCQ5EeLUaxdd69bUllUTmBQJsLPJJbRUSRGr5J
Gmo8la37TcxdcLUdA0XIkugsVVv5JdKsrZwN99VxU0bdV65y5cOO41h7fltD2uppz1Ja+GbgQrdI
5dDUR8fSufWNFdBfRs95vnmAWeds6QmZSYuix7dsXC20pF0iAJQRRCvk4+NtrB/tp3cxxpc/Aqqb
AjEuZzJJwY4PA2P9xaToC/Scqd5rY/BsEiT2++9Nghzu+KwW7/TZf8WFhFCoWlXs4jHDw5Cf5bap
Hwc4FcD2Wc0fVS3o2TWn5Hs9pV6jdBgONxLM6Ou6pfCwTNKatFn0dCCwTsMg7SrzRA6RCoyScW0R
Tt31Gh2Om1YY6C780/Xf7cFUqbpGp4g7s9aGWhUXc8xinvINeCte6gcc3745r1gR6D3CYsdAkgqr
AT6iULasS8qi7enkZ/3VybUGDUwAjlJ9bLH6D3y2jJc1OdehpUvUdYbrz2Fg6AiHGmlF/6ZHsOp6
a4OjQVeAZrZpgk++3dk/zC7H42DQ7OoUjSqKT4vWUqx5RKfS1iVz3I2WHVSKziWpPdM2vOTeRkpE
XLjoMGLjNYAMRd/qvrmmehEer0s3tOL+ndwU/iBFCNmyQOv9JhtzMcvCr6HagIz0dh/ftIhL/2Zw
fAc/lCC3I3epV6UT/jqfkzMO24HX/ROL2pQECuZvaS6U23kaOvKPgEjzca5vxyn8iOfO9KfZuGmP
R7DXgE5JdEkwVI64YGu6Jpcv51Pm1P6dHC/Ji9sy0smEENjV26D/zXn2HT8wUxLNYb+TYcFsJZcy
g6NwX4ChraslsogaSrhbIKG1/HwzMCKmy2D5CM/Mv0arY9Xf+WrhIjh1kGV4idlnEJBD//cCCjq6
jVC2bWMkAtr8i0+SFPPmn7PuBBFoFSut11lsZYNGJQzWWRMJnCFVI2qLMMpH4IufgAH1X9/3Tflg
/ljwR8W35NaWmEo2nDwMt3LpashQPqGCXEsl3sZUAGHNsY6XiJL1zT021KKpv9hw/iNhKDNV8OEh
ypyb9EQJW/AxS1CflM9O7ANijcCTDM+uyOewBK8EYRuMxL5F6GCqwiSfvvrfiDp/MeK6x/BKJOhH
VWn3hlqAVDHIjKclltvK96suygsHhf3HphWw1eYukfTFPpYGSSD/x69qd6T4TeD9GVQPNZJyla3s
gNhwRUOyQ6ROhrgtFJtFw74y5JucKW3J8mXr6r1p62evJB2yAidXwS3sOHmx8d/+OzKHmixK/E9s
rCFeSss+ak2oMetkOAE95ve5QW5zOrBiM2+yQN7rWWs/mbf1KFNp8GItuQNwcaqNudTw2X9kvqpC
LQefz/S79//h3eLPRrSht4s7tXSAqqCNk4EsHyDQ0dDTvcIVm0jgkgKZdXHiio6+oGvhhCU9fDno
Cdayjkz1AUKbhHfWPbBVOgq6jGlzv6hPGVRnG6UZ7oYmN2ZyCjGTxYEsiLh3LAyger+kkeBYL+qV
JlkZ2ZfmWmfP5/OY6Z8WElLtPYYcbclVwUkXD1nTgMUj1cdGNVWyVFReKhzRENBkv03uCVVfMY19
mxMtM5VhZ/CJn5MJX2MT4hh41A9v4V6V7mA0ezhof7bSqHsGxRaOBxw0U5uaSrBae46avJvJyIIP
0nVgXdAxMYczMYd7pFAf8ksPyL2O1TelaYlRfTQllLFzCquYPpDU9HMpmqCfeOFLgTlSfYUwu451
TwmPQ02Lw1iMrnbZVdCBHMtu59PnBbgDag4HLBhiNizUt0z4i7KLQF7v54qV7uYqQ474iI5zwPb6
artDOLLM8b2Ao7eBNPCpo8jkS8MEcoCjr4if0te4z/wAvKTn2ZYlAVSAXJb4rJs/KLnENJrMaivR
oeDCjdcAsF0sASFLv2Moliohg1YbhUTTfvKWeeMhVsF2siYyl4dPIeelAbKPsh1w7vl1OcCJLgOl
IlMe0Zo7fX1aeLCRCUBx15W0UFoAkgYuDS1ddqGge0bVYWm9KEv73olIIdSkeghRgV2K9M1A/yBQ
V88628FpH92rz2dYCztBi1RuVTSyNNC5IN364sGsxG6k+YDz5WBcrR2F4Q6DyxsZAtoqQXcTN1cZ
Zm1MZl69k5hbc3cta6TPMtfdE3acJagq3Lvbpa869Hihi5dP2Lf2UGBo91frjIYRbsz0WaevncD6
X4fIAGJy4i/dTW8k8A/nk4VWVlGjb/xMbe+5HiC7FM8EdPKpAKc/bS5pvRxom/0wxgAHMdYdo7IB
TvZ49bFyZxeft9PhsEqCN1+22pv0GhHG5isonlvWEzt+sfLbfMCC/8UZHFuCdPOPI49BYIOBBlWk
0wL1+eLEkWfv0RZQy9S285aSmyElymO/OOeBHTsRZKWmSB05+RegHNxBaAbBWeqTumDj5zoW5rK7
lRmvWVtDnyxDIM3thWEAcfm3Xk/WV/Ql61Kk8G2e2mG+KvQ3bz5ugammr7uL8wfpisOwkxRzEW2f
3vPR9uZIzQ38dbOCjiNYt1aKEZ9V2M0q8HxsS6zMytoPzQcTSc0GoTIM/otyGaosDHpGbMHgLr/I
x94eeO7svdWlQHmpcbsr5yF/uDzbDPg2YjinP2h/8RaCgF/pe+4J/2PWoXZj1TtvTmhcm+zbkNNx
D43sej44WcOYB1sFGiatKQ5hzS2lR8x0AAHoOg8fDvyZ85DfaNF+y7WV01kCcHoFSLkaZ3Z/JSGU
dSm/aXrbFhRwAkhgoEFSOFcAPCSj4kn+JWU4tQtR0MArhUcdN8ZuqOvOxLjdYb/87s2aLuobf8gz
AHSU0dQ/XBRaYDI6mg2KJOmYZ5gpS5htFeSgWt9nCIDQu8pCS81D9kNovJKGNT6H782ZIV1OGV7o
DJkqRkdJWcCPmCRAnKHZq8PJBXwD9PnckuhIozC/H7jJ+Gr0TH5B4HcN273Gf3Lxsue/aSdgazJH
BwLkyEachNGECQV3uFTEko4huuXQis4hFaGCJjmT6Xyam+BKDQulTQmx0mNL+TFgVR/PHo8Q9fla
zDrZGaPXmlaik1nghs4wwuJYr4qqnTpkI8hzqGA0zVHfskGhO3FWE7q6eTTzXtDaQjZ99lHh8ol0
7X4dzUNZGGZWO734nkKtRHHvXyJYLdi64qnco8XxLmbjiFSg8Gx7TdFXzLM9gmTfgz7P1qkstqdy
mo33iqgDom2eQOkxUV46Rh9zh+DXHZusDoLfQfe/mpZlPxNS1HAwUm+gq2jcwVl5i4rZ8vI6fOQW
55DRVYaSZQP8N6FivMPm57KSKpzR4zqeXPfzHmsrrSFt+t2XbeMrLsS3NusoO0Ol8nXlXxGDHpLL
ZhPj5goU1v+vhKPpQClG6H1/2bOiNFKkZ3OBK1HwyDKM9ySWNOkfDLEMalpJZiAOYFiBs1Hzatmi
HOshO49pnAXGdLwVGJtpdgAFCrN3lllx4yyLpnr796i4qERs0f+SbWW2eSlHFny55f5FafrYk9Rb
MEtL4f9pD7qqiQAOIvLjBN7bOqEG5YF90uq8s6trE6MKKGNapAKLADr5QSO1+vcsuErLkXS0h1Pd
GXsDvuGWmZ3cA92TePclG+AWwQ6lXj8CKes2koatYbKr4oRCOPGm2S3uUpQZXO1qjGWlXuzO22O/
HDtE9C3gUs2qKUaXaMCOt73/seC6x9mgNAZP9ytlqC2PSRrONYqm8fu3Ulo4g/mpWaU9JMr0rHNX
M43d+YhMTcuQ1wpTfo0oHKheH2Ur50+MWigP7Mu3JFrcOrOWJrCbNeclNe77mPcr2751eWrwGQgo
rq7kvlkB3KjS6saaf2ZFXcCRk6U8bHouzkMZbeYNn0o5QoBtwhHp1q508BWbUeK9dAKYjMZon5+P
WLDcJ6DorCYTdQEHxE+lkjtsEYnxrKJKPlnyENYz1kd7FkPzYjgliOAdCnkI8HF9cDRJ/5mzvdp4
TLf4CA4DI6Q2hGqvnTvknGwPRRHXNd2GEBK+LK0dOzjqW85iG06ixvl/FdZaPrBsf3qDLbQvcg/0
OocYv1H9okUABCSVr2ol+/XHfK9yUuqqWt7Wv3IThtzL6xxvspY2E/3R5UkEN3G9rn4hRDzAGEKW
nGWZSIUg4c+4OC9z7B/1CtUGUM78IJ8A5N+Hv40UNLsfXeHmYD0+fYm4gVL777Lb4+bL9QjlomRj
QIm9wSeN7PZwfWth/fIzcFR63NaMAGbxb18BJ3a4Lsaij30NX1a8YopX22zimvKeue3oQbeDHG20
aWn+5DYdBnJSPynPa3XrsCz+HDZbJBhM5wbQ3oyugGt8aCw46GkQ7KNoI0DXLvSX4FXMxZ+FJHet
wWl+f1l0X1iQi4u9aU73cAePhdvq2cgqXdbumZf/pjO7BWOOkKyjM7o5wz58723kZGgV5gyEq9Ew
0oPdCUgQZeR2WqJzP8DeaRJi3U6l43B/gIhBzVl2sU+1thJXCOZKSQ9JiuZVcr44ET1WsZk370fG
ulquqv4nur4mJt5YPraB32i7hAGrMWIvpw2HraEJ6IVqNO9bCqjakFGxFBkfA+ckBnfDFGTPW2r/
twFbv5K6yywXa2GAryQUa/ueAYufBxUtJobL6YBIsEBzZr0Ydb8s8sQZXGWBcRJGj66ddG1aQ2lP
zs+9jT6z/AviOuV/TZCneKO8QOtKGiKh+x6lqGgVNWWAGIYnWbq4/Rp80K0gf/09W/HCyqETiE0M
98xAR6VObGbuyqXCuyBp7onbzGqYt+xZY0vvzl6JZkxcF6jt4+HFj/P+9c7G5VU740jjQv/sM1dL
t7S6iKWdYIXkydWwCRfLF+s2x1UbyFehEiDU3DOcfTx/QvKM0R3ZUCwaMMGHjNA/XAeiXJma4wnZ
YR/Vu24HQOt1ejowxRzYhgGg7U8u4mSZrIL3vFjY3JS6KhiEIVpPd1ptH+Hu81ndZQrPbtQsOMyx
zne/kl218i3FeYCKIYbnkhQMq3T9WvVxVVJZbO7TMgdjXUzSSabiK78zJQmY1AulGUb5AhXdPgxN
r2e9cj4lc06gzrEEqkDPQILGIjg5r1e8eaZvJTPhfjSdOdMxp2H0pJgAuT1++XrMcbWL+aLYkWpL
8ZWTIhuQ6bo1shPxO0dW+c+UNXppPpP3/gNIf/KbJ2NrKsmrBjJZPab9Qs6RbWyFeoTRWH/0jUa9
HusoN8aWZUYmQyN55Zdf3o00ilIbrtONdQ/EfPc9fu76YXh/hhk6q9onYSTOzRh9TWzVp1z/C8/8
NPL4vCaceaevgupEzwbz9da6C0BssEgw30wmyLSP47VJuKo5XEgGR1P44zYSkktTVpesi2TW0Sjs
7HKWMWL5iietOHnlSJSGDxn17zi0GdeMq5wqKJW91Byevzz/6yPifWohdKIxqogUT8BBdIGFHLb/
4LNWQmx8FLp7xzncFmyyYd7XAvcJis6X+hVb3DZ5onSNstN2uNwC7d4UpxVBdRf//uRJ1xYS40Ld
Hghsyvvvyut5fRllgZZY2ET502DvG99QOFK16GJXA6+LvQfHP9Fd9kd3bI8PDjIRH3arSzoLDXka
DF2gsKmuZK44OqmpUXz2HaWhbh1FEIzgGA0u1+14gJJzzOCN/Ozs7bNhd2ft0P/+F+bRylaYUAGD
ieyoHoH96r6Fo51CYNz23N2lA5dcGx1GX9DT+JSfuZsNBRDE7uk+lRkodOTk6N76+klZYF2/sp+n
VVG57rZEsTxUU+8/tUp27hDTjK7FOSPmxBdmDhYFsA==
`protect end_protected
