-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kktzou9BEDcc9Ii39hqc9c7OaGj7MQr++PS34usPcIP5ramY9dl61XTjo2nYAMorhCru/nRVabnl
CP9YHWF5LNOWrcTxgEGzODYNzIPLdWff65cVpP9Gl1d6s7Q07lNPaXDH078uKIELiJksPA9FdTC3
b/HSbRLwZNvdTmNe1vz3vLfuRjy9fO+GqJXuDz1R2c8OCuaFuwq2g9OZMktyw3NYIAPhRTaG3trz
+2z9rzLc6tXQSxB3y2A2nIIBKWwvhPkKfpjNwZ40KnnKVfVQ8mnvtAYA3/nT7Ut+lDsJx6IxkLju
ymY4YH0Qu5THKqi76PamAsQ90mwdtjoIOqSVEA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 119056)
`protect data_block
/0Nqjgpfh+lGsn8NLchlmHL6Pr36/WjqLKbDnyVmtcRq87aORIUDMDEJOnHyNodxSXth/zucAb0L
OL7hDGatzPkOH+TqDIoxIdGOPwFkdbxUGmCcH3p83x1ECLfqBiyNsOTPuf/v+wzQA900lhZ1/Ro4
QsGnBkVjBhfHMJHURuW/Q6VPmk9kOY4Mq0xFjk9q5FAi6aNQtnj46M2fle2HH/Y8PIn07LHkflN4
1JSzgT5olVEXB43vyXk23mPeAFYolg++8DbAiNJMcEfsoaQAPCbtiyG+hjkhQN7o88OppyBVpc8S
AHD7+fCxReUqu5f5t+LCQ+EBN3L8RUphEhEWyMOj8QUo9sxOAHUEJxIf+XyQv5njWlOpxhwMzGb8
gnrcB46pb3NB6HeOIdM0XhT4jRpTggl9JIkcduu6hSiq3yLeiaFR5VmxEnCDZdl+u3P06pSgAfDi
KTQpUxTXzakAFz5p2LSJVZQC4NHwcNkDquLajVyoeZdtx3NHmdw/ug3LqvSX93f48CQvx4Cypg5i
9Z04GI0XuOq5E3vVkjEotGBl6v87LHpNiiDd3Gw3PfneG9iOP1CXlt/9LfRqefCgZRoQ3ktfDyKR
6PyPBK5vkBpUL8AtJ3LHx6KVCtUYNytsadkSF4SxFjBrguU29e2JH/TlfTWr91bOYpbERR+7Di8s
14YIQZbeB7018LirRaU67KgksSfIaaQBl1fUL+Mjuat+zHcMAz59nGSQFatN5MYNBWiunUAJNFOo
OE8RuRRPS+0u5R5Q+F56X7O6EnpmeY9Nyk6sJN1OWzgCNqfkR4fMvrX+JLkPzzIiuip2HxAXFwsE
/pgUxSOaAFDe6RFUiPyqUdq5741dHthtAaggz+QGje8wkEdRqywNsi3+i0qSGeL50UWHMp6hUUrD
X9X+ox53LCe9nKIMOuWt+Y1T9BRoZ3y0OapcqoxrmowtFHVEi4L3qTaUe/0ynI1AiffWPPUVsWEe
Yff9kchmP58HAInTTZWnvva60ddHjt1NagK81sJUYOvo2Ftzm3IMyCk6Ew+JKrfZRo/eYtzEWpit
ihKx7sOOklDs3QIwbSrJk2cFvuLKLyS3PEVZfG3Dy+haQh2VpzTvHC7edldoxADrkqWiRWBXMZOx
rnn+Yd4bkbNncSm2s6Q+Ecq1rfF+UuIv7IEsVyEN5p/PTtgzpJSdo/q1jQ3KgFsIJ/pMmMmK/rWV
4WlRPN6ga8+3D2yWEOHp4MctjFrEOOpmVi0XgHcxb0eK30KPk65pa6aoH22u52X16SHJA+23SONh
iuyfjJCaELRDtYRdTtDG0bO/dZuJKGqf5PqCndG65cpO4484X4xHQkgghBLOoGjIfEF4lwPi0V3D
O3Uz604MlbdzwPHgYrrB4GKZTUTMYp+ADcqQUm0o5FzMtGAsCnCnDuFmSYwFymdBaEs1hLubpYg/
RuuqaDAAV8kTu8ZhWYNQqWIz2zNXy7+p4N/FpcqxdNWLBEPEOBNpaA+qfxteTbuS+wxo3DHQfVTG
wB4dkX0BD7Jl2dnN4zn9EYdlYN8NpAAeCbqRVhl/ZPjmblm71RFF/L8paqtjJTIsthAjrLh+d+Y9
hhIhBgUhlJOkZBSdfS0iu74KB1WYJ9n3LLEINYYQWyulLBgrs8x7S3XSAZMiR70f6LsBoVE2ZNBz
Q9U3IInv8j3EZVaR6KWql4A9WiA3O5dMMpLbmGyTb2jV8CyRg4QZpOLsDvgsyAyPmtg2+b2WY6PJ
uLf53YiVaUz3zxlPS3M5sLveoqlihG2zH78KqnX+QHpMtqgX3ewyM+4ezxZaM09dognK67DMwRey
qwhesfxHy4xDujdnc9ZygmZGCIwTVceQUwGpyEMdvpfoyF23hlfO178CF9qc6v7YiVA9dhcEG1yP
g9Pq4nEkENwZTU3DOHaPIjbeJem/EoIEhigz3NervUZkE4dPNGbkRbNLNKrHL8aZ2M5yyDIIK8Vx
TD260x/aoNe7QTLHzDXV8dxzFKwp2ELLKNRx2ieTyhCGDGNjdroM6HDxiw7nOvRyWlpypg2V3MEf
wpH64kIwko3YptJxiz4lQf0rSEQvXoyW0ZL74hfcAcTrwFW/8ZYcN8HSXjYGkEPyQ/fT0v9itw1p
cClWRRirkk9dYES0dbW5rQCjsVtVW3fOE+/qGGa0untEAhcyife3L04KJ1iFmQdHByNN8FEkvE51
lsfKV7jusjCMkCJd2DDYia2hR7kY36VacWKYqs2YjVDEKekTmmmnkKhrHgxYPDZzvPB+qGpLzLnE
ifsIMs9yMFs1fKauesvu/a2ui00U44Ubro8xmcREHb0LcwUhRm0+LZVdzkZfBkNX/lDWun/97Y1H
BafotX44HHNfOhScUjFJ9TgEAr7bX8S+iAyVxRtuLqh67LQxWCTJLeaPzAK12b2m+CEsfMPQa2qP
Fq06MewWVZrmJ4aoCbsvYKDtUI3Vry4PcQOKybbFXQ/AQv6uKSXtTPNUi8J1K1NQ4XjNk4UruTk1
N4sEpNL7tr9bg7CjjyxfKTs3zqRAtkDEJTxeSQnffF/Hc5HAVLptpwApRsG9m7DlzzxcXD3EChnM
wdORAmnnQyVTNZI0Eypys3lGIPp/gnz6o1uevgphmhP94E66bNg5BhWxFjF4HuCqMmosOCjI22oh
mUt8MqgyQUEEVbkS7LwEJB/fVlg9KJQPFfxe2Q/OG+JRlSJT1N8GrUz/I78aR6cRaA5gq79ZQfxC
3xAh4aC7iM+RTLDqyyh+5QLveOfQOdUdi3MRVWAIUo035lZJ4MqGPRgX1J5gt1++aCisp4vyzL/5
zVZ3s/jriPIUk6BxaqzqDwVw8b9ewfYmMfJefVFSqfZlOKU0badUKbTUOGEXRPh8LeRh/ocZllmU
OmWEJBuUUVWNtGrSvbdMe7T8r3OM4NfB0fL2HPMUbrnKukAC4zKdMMqYBoO9bBpKklZinu8iTRts
70+UfwGxe28eJqKFgKx8BjG46AX7i2aatlhN3OXBAOk5mW0qVK0X5ZkP63X74PMcKQhEjQlOUbIw
H9EF5LQEYIZ0clDYnI//Tx9drDgkin0Hp2uEHW5oBSY/4vEQ4L8L3SmijBVrDTulNl09S5u4nNJe
lN4MVhZIQHASSjIDxwv6vYE46m4b0Ur4UPCcOjc4J7FsdRG7WqXcnREJHLRD6kZwE8YVMrq0yV9a
3v+lG4KQJTs0OFkcewZRewqBf5xKgCV1B61SXSrisO5QudWGnF7DzNdpQRaqmZEimAwavKGllGoD
oVba4UOIOX47WZSjOcEKzboU/hMdn3YF16lfxzaIYw0+pV8/dHBeasex29eJoYN7+J9Dfqq2Zn99
5muAKwrl7N8lFoiZjN+2k7PSK4Qx3LrjG36/5NseCaTFkUf3VwMgr9h1rPnjSPQuCBmQyxxhzX8P
XPbLOH1NYH35mN2eRthenpwSh8uSlbSlTtxl3OiB5kdkJkXZJDHeHY6n1dbxxVOD+OX7qRF96HGF
vTL/7/oqrKqPjnxqHK3U+u/y9gLJ/iUn4VnQkEe7hK6le0oYLIEb+8Zc+IDPB6ca9TbrERvB0Ubt
AjWuNY4Y5wakpEGud+JLGP1H0Mp26Lg9jOiQksaGt9SEtv+VdQ99ahGn5qA8EorXdEDzd7iwF1oA
FFhTgbS9mnEGX4997vUkXZh5zmLzXVz6jYBlmViuAzoilK4HaeIpGrXLPTVvq9RL+2wDeOTt53nM
DFWPP52DSmcqyD9MbEAzJRbDqxK+sPAWNpapvifSrOop81cT9BntnrJ3mv0NK86MsiAp/K0shZQ2
5CEQhFtB4qc3PiPCgEcXn0BQy2Vv7oB8DwA4J4l6ThhlEtt8WFwniDGJsjYY59J9mDVtAN416WWH
wWXegxNVQl6LEkbkWJ8FUS+8PQHXRqbv3xDKGPG1VBGLFUllyHeRo0cGPYa6P7Fsw7PBKSUxbigg
Q/0KySicy3BAGXeUjPrMyaJ8b0j6w9swQVQ2lHn+BhPxH57VEZu/aBQUITSMtOvTViN6iLPEz80k
rJNy7xkQVM5PJck1Glco+CrT71w1yllR59IxshMj+bV/Zz1Y7m+oJxa4JGV4jj5YvfNb0X00oHYD
rJsIGRU+mOz/1d9g1lFW/0Uw4tZKzLJydFzaQQq6pmluIUaQsJUZ9J5zlOIAXGYZHTqkd9nCbznr
QonNdkhFcSEA1o2RQxJJ3k6XrmmsAph/at/gErO7ivh2Q7Hz3vL+KQf82sw/7NfwfNvY7Uz8OHVp
9PelrKvmvnuJqu69Zpuwq5mvmvvoxjPIynwt4BvkDWbeGHMfeo+F6ULH379XE29cxB1uBtAGm9b5
DH+8y7eY4WIZpcyX+Z3brxmPEBJ93XQRK40GRQy4RXZKSw56GUpfYGIgNbyR33IzCrxhdZzaud9X
DZ25WCjI0JipyTBzV8xyJziLI0MvejNs5DgUycq5tT0nSuY5sf7rfzFPnBbVz2EL5ZFTMkii8U0T
EZPUwCfbUmxmaJeU7aap370I6v0wXnvqpanG3HWVmn3KsWGwjNbZF/vhIfFaViRe4GKHyzVWbN4N
KiZTIBRBma1s9ivqxkByVKDwgbLNp+4kUxGljbdFJu/NPGOXDPPJwlgHHIvobU6tPDLwCjym9bsX
2L9kk/Hmwavjxr/RRjZGXnnC5gK7FHPDXUuNbxyUVqNuVq8TMFnEC1UsaL4va7L/zPfJ8BBoqHsP
BpEcvSQUtrMANxaC7wLx1vVp5vvYfDQ00TH+QC2qpEkuXYeTOpceQzGY7z9DxI/i/wcLpWSnQVFt
rKKKUYoYEUsu0xGvCN/nEp25FU1+Z9AmaUZnnKPdqMest9Dzc/+jhn7ku9CWB/ZsJntPhVY+Q4C/
mTAhAns/hIVG2jvk51WvWizLhbN1vt3WO78QMJRP3M4S3lESGapsR2YnixtcAa7WK5iu7ZdJrDlc
rLl1t4FcGnFovY+kr0eI3a75FGrA6mTZxAd4AwTyLK29gC+oIou/QLMHad7AjY4vyS44CGh4t7V4
dZkU7dtfvPeGq0rEXTOBEh7DI3TObOGdzxK3Xj8JJbIyIJoxnBAQrVvi9A8B5uKUIa3HftL9VNuX
hZvFnOQIHKjZS6o2/5omVfRBSHVKb8ajw4Q6XXUPE5fW7/eafJmzb7aU/TJVwPfqKtkp4dLBMGwp
t7Z4QGGYWuennn3LcAqCF2bKMM03s7ZykWyS5ehRJspgyKk+6RxjuEXLfR1cWLRtHAEFWOjq3olF
3hfz8gO5mckqo0oCv2pe4cEPuSUTGh20wWTHiNdW3yPtkyUceIfxe0p8lSnL6She/w7DsTrQooMc
o+3Ub/qNt9SAfpCqo7WYOmTwtaq8Z/ic/taLXwDJagknNPrqcMtWKHbNL0YuI0aUQBdmlFlqeX0r
dvGSHs9AbbnLM460+amPgN7G+zFhK83yptJ6JS8M/5U9T3L7HtaYCmmud5P6LTHeD7Ve4eNo6q0G
sMB+pcBcrnmHJbErNC4aYfEuT6eaBcZEXcoZE90QbNJwQKSz3caqNhxizF/LpBO4wMuvG1DVLB6o
BtGE/ubpBhFBygBkfTmyyHPDBDGiSu0wAbdzdIB1hUTkOZe1ic6OpH5a4segJX+av9hU27zkjA1z
pXLvn1QsQtY+aIRPi+XmSPLkprueuyHYL7ly8nUwmc3iwbTbtPXNdoFytQ9J7p9XS1ns3RtXPzu+
6S0DnFtSxQpSlT66Y02KrH1COhV5qCeFjBl1rKsqsGD98OAdyAcsLpNDhmLqAdXED4DIjI+99pjP
LjSm6lslIDkye+hLrQPxq/m6qg2FobCvB6xlp9ivQO1sr8J0XrK8ZVH5gtqwV+k+b31XiQREX+m6
RZeH+iJvR7FSmQ+dUkrre1Apf4+ODcpD4eqbHcihBi0ZYBPvQ9vcvTcsKCT865p6kHHc4ZEcVXkr
V+ZUOFV+TQLJ/NZalDIRVyRyusDKu9NhGqle1/qKRy2wsGiqZMIw9dpRnqLA2VXvjokR4akFnsph
ObjZryAQw5tTDy+I4iedWJEqV9I3RRPvJA6kHVN0Ufrog1l/izFpS0WCvu9oZFKgdbq8xGUeTRC1
NNGmoQVZtKBQL6kdN5CIQFACSVxnYF7mBrJ7Q8xsLxiaEXSyzRKZbSeM3a9AngmTsGugoaYUId4x
yEAvjgsyv1QRyaFJXNiUzvVauR42GzHuYnTHU5hPvJzgyjFZvlKHEWw0jKuca/zH+glA6oFqvQBw
sUa0egT5cy5KVKgM81QzAGA36ci9p9q56KEGF0THQxlEAvSVfIxcHty4roi/8TLHT/uzWIH7UFvy
Wn9dP1jjHYhs8MqiQaV+/koHGgek9npvH9so41xQsVA7fc/ZGTq5J8ggqsKhvD35k3avBW9yIWdp
TQ6k7XwoMM/3jlJpKKvrp4VgUowzrjstll2ttIhmRraY5TbXMaItPIN2uvTrkCPlkjfyodGGCH7s
ATsqLfdtZUsYUvawkQOTSOEqu3YWL3fiLQ9M2h5SGITL6PS3UPTfq6aESKrL1J6xP9u2xcuS+nZw
teTJYCSeK60j+ViwX5scW5PA73qbn34yfJNymJ3zsxSQugAfIcn5Glhz2H35L6mY94DY5Qv/v6LW
pxtdwdszynyFaapkDNQPx9gCuxaOC9/2e5TdH5nWx7fzPCc1QUM9KpEwhLtCo73bCSKE3Ey28bPr
efqKXnSA3ap6Ww75MhIiSQY4L2DYh992gklMKzM7yQPndFVlNt7OauRpUgjO+kGK0pWRjyDO9WDT
7j3Eri3kRTlJFmB+3q6XOe2DYgfSRhbOvkDiMpHI9ynf2aCxRfm5XESngdLA3+EwKepJO/zlxbLK
JaT9jaBvDOoQWXEhmriJU7skU8ewdEwPI368ipzb9NtIw0yPfmAlCW1jeYzpQe9d0iRlcOE+eSdD
HIgIl9tQ4L+CBeoJXrw2r7n1Rlo/mq6QEpm5VTWUUEDawhDR2j1NG43CGEDIe9uRd14GxLjZS8WG
XUbUhsZRw9aD8JGQahMVHYhpDy/tLctMcOhC0H+TKtJNzm2FmKFPQZqv1hcAtRHkaeafmLfZAOLX
mVl6Wv9udCc/PukY4riJF/ETT/BMDk0yPmNaqazXW4Jg2tdMpfjdqDVw65+GSfHhESPOkUjcZxOu
76pMgd2cswVXLYHGyx/JEvKz4pQQ6oY5r1fXipcQiClLz+wJa/UuU2JLS/pvrx+AnnMx6hcKsUbI
3+BN/lix05f5HMON7wpbEc3QxK1KWOidTlexa+bLoNpAAp7Qh1Bez8sdrcHHDvhDmmZvnnzrnaRE
xoYCAy2eDzbSLiNHEtMsHobs2JkvbRTPLbkT+dERzAtbZa/mCmD1IzadFCohV05lM/8oP5gCXfu+
HUfaSmWlAYQLz5hnN6ty2dnE6/r7dGkQk9OYhTgCKHZj5uT05/vK9ApGD6x21OlfQg/VmzWVI+xb
qZHUzs5i5Kxt2Rsvvea1AqMtdSvq/GZzXNyoYmVe0FfENO304JfhzuExYFhQFRbGFttLdeJskn+k
G4rcOnme8O3XdYYieIHPtPmI/hj3KwAD1oBVqsEofLQFt83vi/5v345H8LgqsuXgHGK847qNY2ju
rrlAXV47Huj8TE/AceMhlRGmnkU1u0A09/3ALEsoaCBmZs2gULQ/xHcwB2EwcCcbgb9llVI2pOy4
Wbc2YfBuCrHu8t+d0F3sBbeurEmoB7nDdn7RIzDQCbQxwVE45P2E18RGxcNOpk5rqQ6SLiiI1TQy
x5gkLvaQB3V6qp9WdAbInnAJw1UBzCEvk7fvgJEp7PuIkzY4scFa9CH0t6Q3Fl0tnN1ZwXgYcdPl
6AZYRfSzNtEyti0yp2NkFTtY/3jMqoHSUgL6c3TMpye0G8tV9eiQG+BQMHuGrC8sePRg9UQwXSvS
httDjSeJz5sSB4Io9khmV+zA3Gr6mobb/bjmpnpMBsjehypDoMH056rLLZSIIMP3CrXiSIuKN0UH
gaEhjap6r+twjkv1GZYbg0d9cDJdzqCOwgNojBdDpsx50NaQedSEduIDY8S9RMLR+4EFOXTWz8Mi
jQWhRC0ZViOaqhc1pNEx70YQADEgtKrG6617FwyiaiMKuHs4oScaFNxm5UpNJxS+gvoRrWSwjzzK
tbqLtLoLsUJhh+qVvx8wBK56ev6iuMRdilTKfH2Me5gHtNdxR9VMU9uBqOjqwFkQDxjfk+MgBoTl
6mJdbNrp00gaMjmxcvHSb7LKAclyajQ2tzznplGJrJRSN7mU5KUQo1ty8E7FITFy5s0sWryTln2l
Gls6+Y5Mskc8aOGEgzchF6e9cMOTLzM+qUz2kyb8kUgsW/R1RfuBMupx9z4oD+uuhYpDuqociQSR
DdN3KyCT6DoJmdoh/nz+ztSRpwQcICF3WjOlbazVV5AR+pKiYYdYWjTNI432J8/66RzOFIRgFzx6
x3pLNI5Fr6IMsDinAU6bU9YHK+dYdw6riiYmi1Vvi+MdLiIeRmwKywqs/CpecSHIlhSybCm3pu7i
OWhfao3dVSPpYAw+H23AjaHar/fDorXYFBA4IQT5JMn/kh1hBln0w4CJdmcgkhKDwgzkZ00zA/XS
VzQI/tVnkjLjfmmQVIwQXP54RvndFdGbyB6g2REcefyIqKFp5qTx/qwc7IXQyxUOOpA+QadrCqkh
QSu6ivPO2TjVTb5p56UEJE9pKn577mCJDq+Mbc084IzFTqcma1JcXT9O4IL54bbhAndx7yd2ygbk
6jK9pu7abpKIKi9k3MblH4douXqrmyxl2WWgPREYdTKoUoRXOf46myHjR7UWLHE/92oZdHc4E91L
zjqnYal+TGpIjRmn7Li0rgheDgj2SJFHoWCsahN3Hhaila/7iAl0y8jM4TA8qCqnGGBYwxqnDvOv
SReuHwj9YTXv8JmY4SWmAC5B4gwEY+1z9riSiFtBBnNUoTrIGWlS4wfriAHUQmhO/wNUVxECdqnO
JxnFoMFF6sqmTfveaAo7OF7l2CH4XrPWriu9qxygHAZBeNMuMqyruod8UONEoqwqmQstTHErXEH4
z8VJFdlj6mtN/IgMdcBtwhrMIkbMIxZuHbnAF//KGxBitYpYH2fgehxQq0BgoTvaryhYGokxvrTO
B7D9DPKIOO4wCCrAeBE8zjZ907fx8lq9c02bEhWxPirZx/8zG3b8Bto9y4o179LAeTJ12bNwD2/j
MfD8th2oCWPeEg2zYbY7+pxFPTF2hq6SI1DyRe2lXZRhPnDsTRYrhukGQi4oj00gvtDLHKK91lr1
t9swJlJfTknWbLshuFEFh58+7zILU2leZ5yKeEWbCVUD4POeSFc4qJLVmqnVlushlraGDcbvVhBz
/yyxsIo/0dvzJcehu31ZUSUYYz/uYn/RToAgyg1WxScWXwXniOX8CTzcjrvGuAe/5+N0GHwBgENU
y75ziVypYOT5xFOndeHDWh1aCcrx2+7MsquXkzd3Yl4TO/G9WBLd7/aC6eyZlcMP1YCSvIEsDl14
iGjsLetmdjAOoRTd5OF0JsGltSd+1C9n/xsVRYZqbQCNLRu99474s2CoJoddIH1qEySse2n4eKV6
3FN6hM59z3tItCvMBNNXgwBF5catO7EIhVeov3ioNFFCa2Jo2GHzxc6yUweo2vPHiw8Kb4Wa6+cJ
qRfQkdmHPV1UXbLAV8RZx12GAJRaeMUxp8s+faAtQxoqOCAMv95pK5hRiKmgoOn6fcck/ChYNI5W
izT0+kQ6g39xMuGeBJ39iKv4LUlo6OCi8Adzy68tvEHQ+wH1RVroCp3/0pIyApi610QUTbJRIn81
kPqXmasWtXkWfvCYyqObzZIF1ggyPIlVwzGNjueaN4Yn5LwVn6o+qhjf1IzOkpANm6oDBJ9/rTp5
zPFmPjRdX1GhWd0g09wm9AWjclTP/t54gekTEksD6mXPpW7GokRIDr2epDHPBI/VY39EH6Hd3rfP
RBRn6ciuXMTlmh+1XT+fBE2t6yjw7y14QW2pl1rt1RWZ72JOul1rlQFGcbnp3wUaXH8pfpqpSXRr
2Z0KOtIe5dLmEkmRw3Y6XGtW5yR2k8BAkgIQRYG+h+ZzPVf4wI3fg6QB2bpW+BPgM83oZsEwcSa0
aBK4sawME4maTkAES9sSC1RsvwZBWVnvKPdpoy9H+kSed0WeMd4sSeNpCB6sUHW1WauGfSpNmwHJ
fp2jvVe98k4DgE1BzVDeotuc8jwtavl6722dGby2ojo+75ApiyNx/MQX6tTBYdti4dI820IXzp6G
gn/eD6hXuQRJvI/KxFjTPf6S5WHuiMtDxTIQqi1xVEa3u1KxMN3sncH/fdnPU5pIxxaAqIr2OwE/
hM3A8dE3sROQuz1Pz0pcGIEo+MsRygj0rjDfzoTmMYIn6oaI4tpOPf9cHZxkt64xXWu6a4sLqeiw
lDxrXBXsAMihN+1fVPZUIWhS85Nkb/hyCUvnpCOJR5deYpmAQAjYW2Ec2NYIVGZnALXh09WPpT8h
Q7EJbxWNOcFfAw0KKmBUFDJRa+QUj1QGthpGx9GZD3PspSKSNu3QSzTk9CFuErhB5pzgzIEpuwPP
mIJRJj7o8ihnH8HpBMW1TkqZL1yxgn9U40NuCTwvSoDJj8kc4wmH5H8HNdQ6cGOLk1eohCgsaMsb
p38eUbW3L1rEHelGrnz805y4d7L7rbF2SfgwBsy9T9R9xnmGqPLItWED23qdA+yPsnfPfMxSYLP7
vr1Z6AypB6sUKTfYkayoJrA+y3sPip2X7SrAymFIG1NLcin364MxgXSsoBsL7pg912TRRe7/mcA0
aQXOsidmpjT83xhZcel525/qPEeeGI/AoPMEgA1k3VJaJQc+0kE0+OR7KzdK/1/4d4oEANNjFOKD
cjovSGFfvHyA6Z5mUFO4qKddt23I0z8zX5zRYej/g8lknPU/oNutCnfmoGTzHAdiYa/AT0SJemAq
CrgiJzSIaxFdNHwPnqFeL4PesTKuyJG/6Q0djm1k7HD/6xYYZP/wIewC30how7TX3plH3E3K2Aqr
fNxIJy0tTuuaxSFMLXXi2UetFeVnjiDaxuAtq4lGBMU5+1odGk3v8/ZvrjjmmLGOQ3PgMB0YB7KZ
wATplb7tbRy70zOcNiLQxs20eFkBmO+N43D6eA3OXofvmH2EXoyg1X9cktdI1yGjXQ+TGJVcHjyp
KrpFrXZMPxDyl9LnQVJF1sNpNHdHviSQ+D62Gxn2xm7izjYW3tp/JyqJE1kkhcrGtU+DsunJovHs
quj+sN3QMKtaqQZV+JpqVk2LecAUMkxy11gHfO4HwL4LVXqq+M0rRBUfr6Zh8DzJhZgsCbHJyKWS
iGwKNImqIFZV7TSInCCHUfuRTlxltZprcTL8GmI8yHRp5jT0vmTk8Nh1Fp+yXyWp8bSLim4roZ8S
LL6DWesAg4SxH3dmbgZS50ujQDtd9lpgJQjp8eEGUkZlZ01VtCZ4my0dk1jpKnYolXD2P9EzFJaO
FWY6eiKW9aud+NzSqX7t6xuSFJi2UsQ4p81pFi6s26dxNJRj5CanL1nNgLU2bxQew5wvCroK38ON
t3KUgtU3KUpc5/4KG3bx49hbCW2F+NsBZgP+L/4zLyljGEwbYEwdymuqOXBRofOM2J049MdRAWWc
Em1WTUHJmEtZAGZUowHdHZQtrV14vVqI0j7TYiRR6SoZlpRVOWHuiATObWLfx8A/0FPoFecjkXXW
92wW8QZMLdtl/l4rsSSfhPRzEmE6JjfpB3waLhNAs1w1YmI64cimyUt5Z9kgVM4TKdiroPcf3l5E
zWdBV3BHFHoQKsRkUZViHpnwxiaOLR1XgtjX/DhcJnK6C/Cor6Dtp2mtpLcdp6MCmMJTsHsbLmcz
v7gQTWolvpiumZoiSaPzcyNtrhZIPFBI/bSG4WDXzZbAhRYRGdfvFwSt4qnHAhTUUW8J2oMcZf6U
OfIvMvLHXfc4Ml1zUCEd6j4JnmiO4xKFnxvNB9Q3tuEFfCcKx+79SGYscRDMuRoOGJc7bBNPX+SM
m/LcaHhOwO7MUvhStujvD6ZvSrCkL99MOhF8YYY5Lc6spSY3RGYm/8uYymmk2rwYiiKJNHUBcDoC
ZE3rQpWvdMEwC6v3SPtW4Y4SQwkUa2V1dij5/t3kamkV46qOx2XdExTs5hl2RC+ILRKKH9ggMKAV
KHn+2GbsinjKKJDJj5mWPnf4eiPbJSTQm45P8F0xoLsbPIT4gfBgMWgsoEKuQmHTSCfK517vQz2V
3qo7HF8mRo8tLqvMCToq7kV7QK3EJzjUewGnPp5Owq6FEejL1tS+Za6mqC0DRPftF7IvJ6MtaOr3
u0e2/cKhg/0Z/6ModnUhmPMNCCsOSpRWn9VImGyA8zSCS7w3x+3VZC/hhVvnlQ9tvSjkYKn93bsW
xnK7Bem3c1fbFaENksc99gZTke4IX7xjk4nrw/y3w+ByJFoNCrg2fxlS3LdfEONJEt+l/k+M30L/
1BUZrtE5Dyt6+t7ESBPZ8brivxCWpOTKhFvFpLIgUUtsFthbCDrvJzSuOq6yxJvOmfFT0WqhZp16
j3VSoYW3whZVwYKtTs/5FWb3IRCnonw9JJYskiGIPDPrSgBrJyiP0pkcBwp7d/jRMTvLxPgTmPTf
MWK3PgIugQEW7VsL2uO287jnpxj4luzNjDDaStptSZYts6bjy07C5r49+Waqt3Oh1MKoYr4FM0pc
bPIoVYuJZ/kLP9kf/ZeQcvKF/L1Sq8dIOvx4u6Ps1CXkJINyxo8c9C2eO5z+bvWfR1gIYjgncazq
cNQh7KkQfkF9TOOmfMciQuwUgifEEg6bfs93sp0PPWAEMjwORC0cvPbcflf5ERz40OyUQlICNxTR
PciCjpcx6cJlXbaxc9+RDCY37Ppaz1mhMdZAacUmMnTrhXiCTOMEsYVjEf4G9Z25qiV6skFtI3sA
9K3WGpV6LVAWDRtgemCKsThDTrmJ8pFHCkCX/zuoqNFNCUJ/qrj6YvDwDb3nY3vGt3n/oxc23dHW
i/rkgLg+w8aqmtZO1Da+6C/F2dhvkQr5TyuA4jRSdf4FgAhD+RZmiS7DADfG9gQ9Gv3kCgHpTpSZ
DAvMaiaWypVLXBmxW1au5Cu3h4eQ/iWzZUeNh2mO2JCmftgoZW444CsjWFWH2T916avrgUWJD9Y9
EOoApvC2NVw5jmCrZsKp3BgUmzmRQ3B6vsD8ojBavJe77HMKOiwpT02VOV+Lva6sFMbFjLBSSVBA
zudUY2t4UTmyqFd77PJ/U65iZ8irrw1xifOvN4QFhQvclX4kcOrSvmVnFm5afUkEsuG6/mQF7D5W
VyTvRx4XRNp2rsFtHNmHN4m2n3wCYF5jmm/SuhUrkdKdD5NQGIq7jIFsKAdj/QqzVh68GiFoS81u
HtuSGxjwDKnu51h1Ntd8Zv8DNJ+9jM1zJ2CBzRre3FArFXA1tHbF8WYX/q2oFSp3iQHOXui0XkoB
E4YDOzaG1k2HZklwnR9i+JL5KZwqFe746EEhBtlLC8hg1WWOLY2E6INhLyC8FGymq0bqMUrSXFYc
QRobAj6BRmuh3n7XvZudA3LbIEN+ZTyYVzWuAcp2sf/OE6QmQfJzI1HSOyxgkT5WMZOfJFcgmDxy
pj6GdxZlShHoAlZ5Wfe/fq9ZzFEW7br6iuXyyvloqcb8sJNG6Q0/9oGCMz/++LczTyh8nG758a3d
EQ3o4MbR9Tho3Xa9aHuZ/gVmKBCaNX6rxR6LVIJE05+pCB7k4+6IgzYRY/JDNI0HOV2cz9ppNzf/
sFLpHu35VHrsChcAWgmY9/pcHzxInK5A9RFP9hvDyOWzPTT+24fhQ3n5hO5eDPMAyI4Rss9mqvYL
hxWmQmzAX40cm0YPe05/XXvDCunnEaXAoySpbQvgbKmw+lrnszwYjwWEVbyJJ5vxrIN/GCEqKB1O
9rQoxFb3kiRbLwaJgaA/MSfMX1V3A4M8lkqWEmy5HMWgKikOQ0YDyfA1gGuH6s3OW6mUfiYpJzdf
DU7bou9g86+fwGgUwSxSBvX/DnShfM3cTFBdmcXSLJCsnfy0x/UuHh7NO0sgARn1/R8kk6bkvSlW
keHZX7HWB8YU2xckfstF1b3P8/K4zHtwL/K8efK4c/61aBMRzNnraAPDXBPsErGSA4yWGvFnaODG
BF2N06CEc4Kx9iToIwuwhncg30D4T5ytaN9CtWZi33f3RK9mg1klTsBTk5FgGUoG5zPcZTmOxcad
OTj226WOomQGj+v4T6Zn0g+L0sbvrl0vYlYAXG9jpOGNc7Pis0PzS+LU6wFeNofAuqjlM4exJ/dj
PBxpqrA/foyxkwjn4LFXgcUF2j5eRnnlIBje4KBkrlQFL0Yl0jLAxHUED6B16Nt+mbA6xoWpG9Al
Q1RLVbTsBapGDqF8QmMy029iNjBWYuGZRg8zFQknO25S8iVb5V3PaX7uGK3Ta2JuFyGvNFcdRzMK
1WexdV2Ngo05S+h2yWiHYr0j9lmob63ftMZbHAl4Q8TqBiJCSARxGJH5aua1W9/CcjIOop2rj+ic
sUaPqYmSwMY6fLD1r0Ihj5+OJQ9bkJf4Sv53PMWRriLuIJT70kNqE0TN/KBceLtdTnmXlIohTLlQ
incNgXPPl1CSS2bZ7OD0ubGWxv20OgBJadgQ8P8UOgJ4ayslaFoOR/EVqUaPl1z3ymeCvRrIGrUG
ftByPylfnO9bUg4I2h8spqucO/rm2m3OIBHkSQOkjVjCCbiNxOgzEkbdshUPoIe13EiHbrGfDWkd
yhISv1iYOQ2MH05tMSPpov9O97MlACkiAdUKgWko2llNpgxXe9j9sMjwsUfaGGZNNgL9Jb2aeYKP
LlnRdZUA3ZB2gX4mB89htvvKLqyKtjiPZmC48TuYpmtKyXJ6wX7eioX7XMiSEVu+y1B2MkwLiKIK
y58CgoxaTUh/COt4phN2rj0ZBlbJZCASH9+Fi+Lgz7hPhlsnmY6hsftiFaz0mbymUu9dpjs/10UW
DU1JaIGH92UpARksOVNGvA/krMoCc+yfudb0bNRgY6R4QVrxpDe5DBKwLvgbvMCmd/ry81l9VuVJ
1pGmvJ93z1TW5jLvhPyDupaWgKY3wkru7XLyM4eUekJFxPIa+hNyoz8ckv9tRaZljcCZrDzU3JUq
npchUsgqHtBPB39rG9uIKxEFPi81j3i9k0PwsoG84HkCILuwq2JMENYK8zkdPHSNmOfXQSaW2BDD
pcWlSDtiH96/WHeLLpFOS6XH7DabLsvTy9fsQaPKOsC34rG5fpp/LYnUvhVTVFpqhJawNlP/DmlT
EaHzOH6dpSvG1eQ+B2fH23ti6YyyPogeSmYA9oJ+dMUY9Yj7Pri7R50574DIPaGlbpLJFSzk9120
qreAuflCWMUM+AuwipXij9u611py/Hzl8dCWPhPpT+Lj1X962CohLXtGpD20uaoIMRPB+2RJICvs
lMeNLAqnZRhVPIcVflRywhx4b3kIvb0OA9XvxZ1x1jYGHdzPD7nFleFW7P9O1+jI46CcWqGDkXKW
BJVNwCgpxJKs1IF3pTluxhPFsVw0+0DYq3YAXrS7A93wD8kEJx4nR6qHr8Pqri2GM+KK8rv4ytFs
Kw505RMDfQjGc3MPbg1Yio65Odf5qr6qT/yZ0eUW8PIMg+p0i1dqYeZJWah4YGdZcvnHsneRcFvn
IyF7ojXmumb3KknDrlND4XaMjhvgFUl2fra4trU/dKlAMqKkZNh+iqZxLIaruRVBe4n1kYO5trIw
zyp6Iq6e+ZVS9RgTS7KjLNwC82zGAWCR+Zksr3VOxGAYwnFIWqbB21rUlNIiNZp6jFYSXfC90RHP
KevQ9gHw4iMpWl3/ELrR1NzANXoKqIeZ8reZSYWkFd/xuqGG1+THd5mh6xa27ucQNADWFgxgsMYj
LeciCcvAy6BEbW7Yzccek4RJ2P1yjFnIzpJqOhTr3NVHRJMisVhT86FWZO02UscbRwxkGFPMXaYJ
xSc55i3G16QMIq+dZU6vF3gNQE4dEBlE5WlsNPIIgFup291DzdViKjQsz6Pu5WwslL/x+RkNOM47
HgwC8ARAzLdrwQXxqIvyUy/Tm7NDT79cGHcVpne4Nx5NSA4tsNczFJpsew3JTk9OygPJS5pX0SBV
ZW98G0Ka8o2GZGTHLr2cSUWsaUbb1ILK9J28K892LaVgwFj1eY285shEkA7ogfEGWoQq7ksOi81d
p4yMfSkKEYJuSKEk9oZp8PK0984kZHuRIfNFH6tX4lNYnpPKtzqGHCzO7KR41p1Jg5RRS8ZO3Q7z
s4MSeIdgjSmFwk+41DfgBwG9kDqRtkZ0rwttIE+e3O0vKEE/JEb6owXvbvyafxzTJE4EG9UuW2t3
sw3KFh6TsuH0tNZmWbVC/S8EHxhcFJKAJa3ly0IjEYjhp9wFfCK6qQuY2oT9wiUxgoEZNTXkLCvR
ST/urdH6yt7lvmTBBYTzxqGU7N9gElw9j+ZPjHAmael3uu6tokAK5OxYILYJRoJ7QjHlGPYc5EuH
75r9oJhlyOL5vsyV28aFzmAk+bvg+r/AJEVcGJHF2Ln0X0G4M8TTayKksy9V9brjD1mzmFCMiIdB
ggP5Ihh3O30L/X6ybXShFdda5tCRN1TNduqM3LqOZ9WU7a8edvNwj3VAwY8jeV1wF+r4nrHWxC/x
aeHmsWEkN7SCn5gWh4/lbpxAgyagqZPdH8TE30KjRDhyalrfMsaBqATT05xOfsiqiqhBvgy9x9rp
S1mp2AGi11l3K1v5WW1e1j7Bf9gI7Xiwy0tDKqCgG62y5376dzy9O7IkFbi0xO4zfjqjR//Ve//K
4Sk7lRjy2iRzggXYffUwjAQKu+Ckpf+YiyrOcy/11l/7rz9BKsshvMZty9U4GxUErRhWHk8leqzN
WfA+BX5ypVXnv6pJ9sf/2gBQdBkPc55IZ+YD11veBJ3oLF7/P2Y3oNNdybn4+1MNZvibzAUa8vz3
px4xT9D75kxNLs9ejWnjhfZwVIshLEn6MMfnZFM52RKxcQDnjJYZ6pGBeqv8o2mDm57rdMRaVU/0
mcRu9d6BgU/hIbUu9Yg8Z9x744jl61EG5ntIcffVNyLIMTV1QEJQUewZ0mwFebMHWhm6IQDyRDJG
Skb3Y3dPQXVQlBTdtiWcHPnpo4Yg9Fmp1IQbdH48x2G0TnGkcpG79HrE7yzs02YffYOnUgqu/zLB
z2q3ZVI/0xOTDqUJFGLgDrOg7nZ7DbAXTji/1C6UO1lg+6kSziJrKHzfkxiWxNqbmcZMC4YdstNl
KLbYwIlqK1nqFFMnFbN2rMINoiYiN39HX4ovaOTK5aeT+2dTx3I4WVq4WXO6TNbTRzqx1PPfzgRZ
49arUrURxNe3z2N//2rO0YOUurefLlYc0WgpYaaBwa9w9XWdzjjm67m/l7s32DlNQWhTTAA+ZUG0
kPimD5wmmqlh4+xcperr6n22YijFhhUKiq7Cvwu9pA2JvFQt57Ahjn5kgFGbowgatdM3+xn//bn1
KnjMNukP5Q+ZDgZS5bfsCUQtZOkWzzFvhSAGQ/ELUr/eYvUoG9g49lsZCNlW4HEfFvH/AqQZbmYk
sdtT5R1p9UPB7EiLLaBl8h4ZpzeQ9DKWxXrDuwaCpc1c5JHys1CRVlMLSEczwdbTYbsKGP3Wpp2L
6XBwYDg5Jn787jWM1dDhpv+XazbKYTQNzumk4wzMybh6rxfLkgKAns+WmXALPgSvCNJ5ada6ksKw
jX4CyHhJ4kig3wRx0kPkabrTps9tIkoRsSrCr16N3poz7FxuIgAfq7M8psb+evccHDSbeQqYBaB/
zurSm7M1wQ1g8cOmBLM2i9fma2psTdPiEfHwXwjOMy4k9nOz5qjYexpm/JbxwvmmzbfTHEfzx9jY
8LWuNHuUbfQnIDSJ/VUiFZkDk7VDJjyZt7KzLi1yHmcGIHs/xpfnEeO0RYctVgee8t5019xK6OnZ
fKCqUPZeFjFSliRcKSgavF3w6DddnY/BhFMVRdTecskbpVAZGGmO9zAFxYTHzOSQyb3/REaRQ1Tp
7u9GlobEWbXgJXtSdiBMRAQIzwgg9bgCkSNTHDTZdtHfacWY767xYbiTu625c9Y+RLE034s9eAMi
u273Q2ue8MjwpyeOCVQ7V7hXFe9NkpJMMSPsXfsyiVwWoL9PNR/Nom6UtEk+6tyhwL6vsnCDiXFM
GAV5sJuhSjxN/8o1GS3ef5KIQvr10nDud6cthrr8J3EL/5/eyE7oFFAoxwOlgYQJ/9EifyS4aVkW
enHJHU4Bmk2M5OFudzrJPaTEFvFo2mdMfuFScjjc6cvs9UNM+RyOWmUL6xr0QzNfulnI1tU6sBN1
CcPeW8CRMN2J19e9+jeNKJOGukgLCnox/TaoyxGGjKygThYWNcCbAyFMSD0SC26jxTFcenR+BInM
IT+11IH2oGrDNicr+0F1wc5Gezg1t4jSdLrQOxb3UWCprIVgrpZxeRDInG/b/8irdGlVaDkwQCt4
+GIbiyQzuMpzl1ZGgk4WI7ZNnyH1EDSPtJyigh+EadlRMHYK0ikwxzTdSu+YB03zDlTkDZzcfbOt
xnALk+JU2d6pxJSrBpGZZvVCp7HbNW3JC+kP0d6FaiboJ0/20Yxh+ep5rfwHyQXzrgv3mx8HS6T6
PHid+EIEd2U8rpHF9yRqunm9QM1nV3/oOSzaU3OvBLAgO0v5AksxslZNCjyFnhrr6yRIpHHoQ5ob
6li/ln7S3nNnvx2Ti+sm22qrVeVnQTX+QjsMIP8iZs10b/WyIFxF3I0FQ4mEtGGu84aOdIuRv7km
a6k2XvR9aKLM2JlCw+bPZqYe0E8awceHpXHmVraPrPAeT8oAsPxJcNiYEzEzyVKvrTFbsIOmvABp
2TyjhY51ocpe+puyi0RDe7Z+haOMWGiOO/KIN+LjEHSu1TAtE8egC1mLh+Iv1JocnikBbtt2dl1i
uS5CyxxM64yUdTZDczPb/wPqZt3jmFy6dTEwwr/3zkY/+U93mDZgpqKkXMdaM3T/DCMtW2IbMzUB
eszWdM73A/u6q57pqMNHfAetDXQeJKMrCEYsoPCvY0qiur6x4TPGJKG88W5b2drbRZ1LeOqgo8LX
zuQA9l8XWFZsBsDCb/x6BtDBlG6U7Q1SkVkYhCXdiZ/Ftn4U8PJTb8Vs2LZstt0Jl0UfQTiKn75r
yG0Bi4E6OIQWSyC8ejNRvMZAbfgVauCFBhxi8bU5Ewt8lLoL+gwlPgY4HwbWxVsjpakPSiRMk+Cn
u+Y+/xeSbYr1yIzGx2XRfyXm+emtc7ZDSMnHdVZmcmTkiU1x1l65zSJgvxu+5vB7gfCsMy/q9WGw
WQGfNm1JU101t0A3vHYlZ8FJMtPgGLGap9yT5teyzr/IuXBUuzehweX334sncu2V/LVpc/L48tnj
lcn/EtBf+w6/wOt6iacNSr/Exj5cKkSaNXGH1W69tEyQ9HFLz68YEIBqJRpqvVFhA7IujHT8I8Qk
WEgSPKCliPmZ/UtKuidsPiLm7PxjiLDW0Z9TaHBpu5kWm0eBfqHH7JFNWs0b80PSpIjHCLE+T1t8
1CRRfcDf4X0A6/e5FFEkaIovwt/veYfrI5d1oaMzG7vVVKWqRPzyOC1XU7StgoW/vVh8O/esBlgp
eznr+bqBlnZp1yj4JbHodEeB936+HeINwrMyJVs1bgLWXxEDtv0yZXFDA8je9Rr6/jzjHbFgqnce
UZZS9QBtIMFb2LX/piMqZbrSKu/aB8ujKDHsSqXnQGxM5BcF+0QLiQMLntr5p9BQ4BcyfTtFqLsL
e1AwiuVMOer6aE8n6wwn3UBC+jiOL+HA/+2aw9clKDtrFeWpjzk2WHl7ch62SYUmnOZX2YruSPih
O0SOOXnPmugqDpJ3UQfJUL8soU3AbqIpXwrYmDc6M2N+fWBli2Hyntr/O0OgZZVnX9Z9QjTtRU8B
G2aQr5ib8DQ4RnEJKCa7A5EkDJNDJPkUs2vPiRaPRqRQGVjRv3C7fPgMXVj0aSU4hdTdWWqLY9Mk
hoVPpvz4yf8P9RUDxaesGGckqW1e+l1sR0m430XftyY5oByQQZVWs7kh8RRBdSmH+ibVBGF+Bqpi
ykTvFfK8UJhkHdqQZDjEvlf/tr0FfvACGLZmEROlo1WcrkURengLoM1N99b4RcqITqGQJcRyttaJ
XxQ6c1YYLy+0/uEP/UjRhk6Zi/mAm3dgAEdiZPCdQU5/XpIYs9j4KEk/ie1XKGfF9CWp9IrayzgV
TrCSieFRG3v5nOB8OXgR80ZD0118yYT87OcdgIFhVcd8FY2VP+JN5FGk4fddb/Cj3/JNQRXzRM/3
OsD59ftFUQyblIr3clxX9mUOHnZHpbyHTIVwJxQ2Ch0eHcUZfxviKJKF3f4PvzXWiUw+xOrGOe1w
cP2yTahqW0VHFATyOs1pim3ZGr8ew8AzmKJ939ERDgNY3l3kyqSErNG9QacX4tK6DRjKSr8T8n0a
sVPVoImLLcLMYZ3GKscqcJ82U1jpPvrlelY+0rn54VrJ6lYhqSYXnJE8l28dJcyJRMPxkei8jVUw
GuOkzB4EyXe4pv7D6MOVpFXNyvzUqhn6c6m4aoTQMWp8i1/RezMBCL4XiMwnsg0ePphhZc0W8NuH
POF8X9OCyAx5//zz+thVkvZbuTRe+yYhSwFrQPrfLPet1IuHfMYKIj+2HW2KzlsfkeWZiVqH6WkO
b8mZOdl6VWlQ4DS8pytpliOO5FcfQeoOEmFODTAB3tpGPClrhbR6upVBtjhEbE12+Wd9Suc8ZeQ9
yhBiC8BSEOazjinIPNho4/eSZCF1UUvqUxKpx1pklObj2etxBAwYNXqtm0705pEYPmCw8Q8VDGAI
nllpTUdQFCbZP4MocvLxDLR2PIG7qh/6evhYMsh+v5sMxdk6INQq/53L2T4HbrD7NY0wuMig0hiG
wz75I3YyZggTkVfxHby+JhHdiN8pZysraZVsvjjIlE7kganx5qoXrN/pNW20rS56lB2hzjuz8qpp
4aHBUlIdDLxxi58BoM7nOhfDjYIE1EhegAe/kVEBGI8jBeds6aZbEAj8CejbsDB1UsJifbjWzUfe
OGLJNGqTHWcCXhKk8PEgPpFiWOAgMe4D+jyX7OXPnAlURcsYbPZEaIqDkQ9ubQKCxZxLL8OHGEVL
Y0DjfgvjX3XWs1SVHpfQQiq/OURyYe4WtJ7nl6wF99uKcXwSd7UjU02bRF3eG9TCvceE3a33+wnS
oDbiWo6UZo3wS3LrEh/NSQz2YJ6e7af5MVdejPXkO6l6HDEOdiEsoegUVTJLXMWTv6VMPmgGv6GY
d3fbQHJrGREM6xoUw1x3fNoaKf7bj4AfMW2AzX1BRBJ87lXPb45ZAN+SwXdWMdaSlv7pFYAESS0O
gp38NzuJZeZK5Z8JyMGDikP+zuOBRftp3GRU5EkL77OQEp+vmwHCtHbIumNci172xBeAphiOLXjc
RPuH0CtCFFtv/lVoLaN51xIRO/k5WAXi8e9vKC+LObopOOddzeFqRRdiRup4NU2PHfMIJHmypdBt
Aw/5X8Ypq9dAH/yDACQ6NENc06YAOVlwgPz7qhhZ+BeeyXkSWhL4M1M8JR88j3Uk/FwFnkwMcHFS
IJwpsLo/Y/H9IxX6BACancC15zE9zjmR3K8wKtGYYTg7MgpwPrXfx09/ZUT7M5z91vx1sgqaAbfI
rMVXnDbXMM0M+Rj5P6PZFOIHGpckyq8ki1RSiw8SSX8dVwkTd+Hmt/ASumBXoqvPb1AtlHnEfwhv
pPovl9QaNdXJLKQ/iDrTg+16/TrUb4FkxVzN2b8MBYArVjVQKK05yLEPqfDxq8hMm0hOtEU59kaQ
kpHzH3bYVB749W9161r4S2wfIOxqimlmQZdLIXr8tnGLfdi+KPG8QY+2TIW/eob1WVZCGthmp+Gr
xT3HVKk4pSRes6yrN6EBYNXF++48LhxZEkn+GLWsojLvw8QTNr7Y1Ub3SNDqIXdL2dgaoM/oZWpw
MDvANh9/hI6A9OxGdEbeX4hGs2p/iLRL6PoZt9pMROKX8t+AhehQGoejo1T6xt2W2UJquGl3hXB7
NMer5mXq2FqERbYlozutLtenqcJzRazkFGkx851VSAjEuJPU5s263iDJ51sTa4WyqCDIr6CNL5Fb
XYvIGEqLsiTZElWAmy4LfM5lwCs8DQ155UI2WdopO0IDV/CYPpos45f5KdiEX+IBtXxvCNw5ZMif
uuOlpetTpbkEiaaDXdmPl6mO3d3O1rZK6EJQpA8N76lb0wiMkSVnkkfoQ7rxryMsVPqxw6AqFIrV
HxiXpxK+vIxMd7qFrQ6SE1poG0kZVALBHmFTsOzVqZrg7Ikid2VinXUbRw6YvOZh5llpePiChiqZ
iMSiFfUwDP+UQzVdtBQ8XVz7BFQSNwSegxERohXw25Nzt2bI+GQRMXRWFUqiJHIIW7yB8HWwP5NK
RO7QPokBfKodsCvKOqnLNFoDDPOOj8K1LLXpQ2I7iQ2b0M4rNN0k7lbPCMJIed0JzWYsq2VmWoyN
8eBfE77rXlySjUtMnZ83GAOaXuDStNiTUTdyIM+DRAfE7NZ7crJDsNep7kvzMOY6BXwf73mP3ALz
AvBJJjCduMlipHsgcERh6TFu//3MFbT3ycDMI4FS5Kp0GeAf9G32SuPE/VrWQKXNKlL6BZhhpnEI
VtUv0nNZlsC/iHlUGKe9qCYvt2p9J9V9z98DORNrL+BclZeGl0ItSkm1o0JyKkaB9F9+1S7o/rCH
4TRZ7gjdDg1xinu63/tcNn53LzOjNJse7VsKxOlF67uVnVsvpuQ3CrqO3yub7m9feuCkSEZ6FOfJ
CGwXV0E8XaftZNxan87hKBmj78ZaeZijoZL09v4pYH+Yargk7LRxxSa24N9R2nWpMJ0Gaj/9h3Rn
T41lC+KAAczlOG9VGxAH6nuB0tWWZmDpTlibOXwqwNIswuv7nTOOf9sej+LqNBTi1YHFbSEGywQ0
aKlUozVz1ld3bcH4jl49NpgQNHipz90LcmVxMeb5wvXbNBm4zwtTkS32Q+dMeOEAyxH5UyqHw2Zs
4UI6CWO72VLi6uxWE3tCFFre8p+LEBdxUJwSepNFlvzvnpjovzPR0F5eWjc+iHwGC6LZa5wDtlfA
oiymTTGsF36ge2bK+gj87GB6t4pUH9sC3saP3YFB3NHVKeZhdMh4Ge2bzn/ImuckXANpMoY7aThH
otk8WyXZmdfoKXNsfRm0y8f6u+WXwcHRToB7eekDKQFZp0rzlA32u9AuRz9Q9U3rCMrsGTjt6lUH
+lhuBCPVD1pYUD1fMRo7sCNS39I2nv78MQrJnw6ZfgltOTYVDSdL41bLujkaSF4i9fFlQLAJI77/
BVu7vkMRNCiTfRNm94LnRnnA1RJpH2OKQNjA1sJypDEvyDyIg4jvCGGLefwtYfE4hpWSRwQWCXK+
6/Zew3BSHCTDYy6U3t73rmSP3GzOsCrXzRrlaMVyLXEr9lFSsfcc3E+uv9UWQ7v38h88+Cuj7GFH
iaKmjLn0Vsj6m3kNKmQ3vAikmOCVIX3mBZkY/7SyxV9JZZhXDgA3NeFBqKbv+rupiWG738y21Yas
SckDfj2kyC0t3stQYwzf84Oaf3WxQXjrBTpFsngBlKeowW0mbb8n1CGlxNiqAYX/EcWZ438xl/of
CEhXdqcq5AxbR8m61ebr8VH30AVzOHCOD/cVxgd8zIuiSPLQA5rLiBjFqsnNTobf7CWVwkhrQECe
fCCfuHYXcH0thmhcWbiZo2i5dPRoHtT1/L+J1sMReJbh5AkKRpQcj6lHEvUtkAunnd9B0jpEYzJ2
n0XylyT+jDEs39OPvPlTfQXM7gwYY5McNLfJ0Kzcso1d5IM7LD5X2fyvz2gUGz2VRiBcSRkeVaf8
XweB5P9rsxY8TeMlr2DmgjbsctyqmIoNaJtJSHAdSoSHbYuHaopTJyvCnPOGnKAXfGaaH407JlEV
Ue85//yxU+0XbAFxZmnUDMyBCxfuskAuemAq62Cdq20GROPPIuChKPsja0Ly14ZjJ2/49BIYyBNY
lagwvz6CRtIB7LroXJnnj0pDmo/h37dkOK/63gtpah+7x0KUK/uAuzCbWW0bzZWjFwvcZYUC477v
QC1qLYNRDzmsSSri495Ri4U5sr0wLAyjShR4velA/M/6Irjqplo3ZZYyi2teOQX3cIH9HCMoEdUy
2dRFU3iiC6OV77J2HSDeahc19xY86mWsZxqhjVQYpJ7ydoqfG3MYoaC8UKOFg7Up243e6gGItCuZ
/wmeyHlS9MbyeN4+YgnNcS+k7JU17ZdFCT2a1Rx/ShYzgHhmmVMUsHRWMVpdxwtVV810P+H8RTX/
d9jQ609891C8PhjCG931oQKAbD6dUuPGbHtfbpscw1aJKYYYyq4YMdOn2OsUVf5jbtdAd83Ax60p
wagutzhLt57/vDiiXV8Ycx+eMuzyXE7QTzIjZiMW5E5jxGAgJYXl5ng/kU+J6INfwabPxeeVmeyY
3n18SJiZ24Kip/m9w0+hiM2f8x/Ewyc9PeGt9UU8FQEFyrYF1QHejMdnripRarPwahEg0tl5Hmfh
ze69xDnyGGRLSzxU3b6+T7ASvSXhOQPOHO56BBa1fHtB28fOd6HNoJgU1rxHL1ewjRaVx9BnodEF
U5Ay3BAUzn5aKwHfis2+rr7FcMf/IuARYc3JvtuZNmQb7hSvDQN4L8ND3WP/W8lxWv+L8SdUPO/i
d14fN3gsrTXQ+bz0e7PEkPB9MlLau8noeS1spG4UBkqH6EWqkN50Gt9LFtIMpSOrm4BA1Gr1kgac
EQdEUUDsVcTslknm0WMGFhLNPvw0YNgJxlqlGxZ4JoHf9mSc23dU3kc6jA0kDbWNx7bBlhU93CgE
vHMmCxnGz8c2KO7EZ5yAAna7H6EfV6uSrJ3ZcqayF10sOTKe0r02Pe2sb3gx/KOHC3wMX2I/j6nj
xQP1T9WBISjM5p2ORxMcCa67S73ShsLO+z/Na4/A19nkURypfnxAbPwdfbxrw5D7B74LP0RjgQ0j
EeSmqQdkv81Rr7OLpaLbewCYuEZOAdGahpEm4nrNskD9dfZOSFq5/YLqYjFYO6bwjqvpEhwX4TNz
FAWbRIyFzj2RbGXOivaMDVRSjdmRaDYPBQ/oqJaOLwq2xTqCPOBz4NtZeCPTKsoSwIRJipXctj45
Ix9nwrDPIarAHXiGJt2hlTJxPKv66wQD50aJT0CAU0n/AD7P6EbD39zCYvRa2wO3snwbJQlLIHhv
Op3Mm649Zu9HChfCHdtT+tP7JnwixwcUSpd7R1xAzmbGvqX138JNBGIZyA2qmc3NP4VH45OMT8QW
e4CD9AvEIS1c1twWfKkL50U4BF9QbgyrqLykx9Q08MPHXWuln1dOkIykRyYcapL8Vg0nvWD3DRdf
YgTmY14qFpVxciXmunr0EjnkBaEZ4GtusbJBYvrbT7qaD67B16E4uXzMAsd//8e7QjJvf1Pifz8Q
uo6CP+nHNA+5sB8um+tKB18JFgBjm9C7bTSuxJXEVpR2uHJI/1fJrB+K8Csf+1SWb0Pb+vz5EQqL
kKtszNX8llJgktPDlOtNHSQYgjXzyQCukl7BMe4JCJirSPy+Oi78AwDfTsFDzx7VJplnUcAdyc2L
l4MqdCtFP68nwN9q1Giw9xybt6XwNoSHBZ1XEHNlsWyH+LnBHcG+n9cbxNrSAfmFWnZU4WIh/JNF
VZhX4RE7cS0xxxLnWDqFicuJ6vwjbBX5mm/RwbJVJrHpcCozBxTZlIrETTZuYkUAiKiTxEvfkEFl
pSaohptfCwDHgW49Z9W8dgGTdi7P8x3f/vz38rfji6rML7UFVB2XbiKEBFFgFcNY7XIFeVUwWCfu
RFVmujuKB+6TfxLPLjTkY/oe1H1VsSr6TBr4mBHzTFh4cpqo3+WO1oMdbCx3ky2BjEoJ0EoyQVS7
VNqPy1CKDqdvhtF1Zvo/wrNbTifpHNuV+j9RAPaWSUUeuemn8qk89rhIgwQ5Lf6WzGIa9JOeMxFz
miYJ6w/024jlf5Hu6F+OMSCrFVqhW7jLybYhFyCgihMjnTWvV/czwbls4N3n1h947G0zcK8qtFni
G6MAPvfyGfs2V5joQNrBZSQdxm2bFRaaEazNRqcxLyDJYOdsytWht42VBXyhaUBsXncc8R0B3RSi
dmy/JKgXmC/6PAGNS1JmegXvA7SeJR3KCVK25d1NOLg/XyeJIK5DI3Ax1WvEkulNxA6M/jsNKDZT
c+fxHIXzlBGOeyRMTFauA3oSP6c7crqmtUZvVl/agNPJFZvACU8ReJszuyRrpPzSKOJuZcSie6Rc
VEpPXguGEE9pWvxHIEpcT8k8VE2dEXeGTssfJ2v/nrx5S2OqFeV/nJUfc/+HMmTDulxYN9+V3xzY
Jk3quGDnV5I36LJ9k0mtxRuUZfxMpN5olibwsRImrWQ9zIqeS+UU/LcLdU8K8Dx3jyAnfrjYUmE1
uOaji7VHDkD748T6Vj3/KTXmfQNl73MzsQj7P1T/2EGBqXZAKB9x/H16NH45H9VgiYS2/ltPfbYx
roWDFUxsmXckk+UhVcI4QLZ+vvCcwT5sFFhgQ/d5B4S3rKsdgkKN9xOHJqI3lNT3PT2LV3j/SIqg
GNWuA795wb5NEUfsqMAZU2eDvFu5C1ZZIiEMI+Y8uN9+LbULkIPSeVqW+AlOo3favpLqN5/IhCJh
CxXU/ZMF3iZUmCY2aupsZkeb7cLFOkKekg620JZQ50NgjDRzhznJqgafMhrDmhaJSNCD39PdQgSx
mdtZYnMEEkEpKVGduBi/EWZhTAZozChQAhhxQ7ROd+6DmvPbeYmH+pq5KR/2ZkbPrA0IQ70M5eoy
96SXVdXJHklP8ViPQ4IQwJfDLm1T7+ZITlBdZgtNyWzvjPA5ELsOLDPVcgUif2INIOWpVqgrmsM4
U25SsEnO656x6BwxMPT2YA8e7CjKHIuVlwQ09/1W/73XR1y9vhE9qHKPU5iwP862z0nwymUNk+1J
LCIlD5TahvxW+oNZ9SYY9yRDAVJ82kbJGVW8AINTyeYU4bg+/FzfVEdtC+yFFyHwaqkpTTaLLBCG
8Q2T5CxVLotS8HcQvboANQJ2iwcyvmyigOkTTuREgqAci+G2VGN3oQL0vrJRFgd4o4f4wJG884c4
JrEebb+AhQmiwNbyi4zKGq9IVNJIIqOx2IKuaIKrGTFtMKw4ufFdiA8P/f7BJm31OU8AojwGPUqC
xglc91TlixYD7U+sBDTVS6Xyq3ptWp52jO9sj/tRhIigGA70CJebF3bAij1OuQwhb4HOMXrmjees
Df5qROgoPWYlIRn6knGLS/Zp4b6mTpSKBHoAufGLNusx9Ww/gsgYwA/ky7CQk6LjcbU2Q0WZ/FNw
k5xiZIlmt1qSQkhwEXqmbKmPzEN5oGjvsVrgZSV8rlb6CAhH+oOgCXtZ2+UhJFH59BGKanYxId/o
ffr/CUPLzhMuEnFGRPEW4yu1SN7rZ4eQNr8A3tTEdzObFkk7qu+IE4bNO7Fcl2QofgevzWPnxgXw
CGp/RUoc4a77bBj1PbSWGzaU4/kKFtmVWPoKY9HD4uzg73AQxXpJpJisj4Y3Wj5vGjgdFPZD9gSd
N0NpU4LDN9dhUEUmOsSwEEWxzktQ3nOc3I8lUkVUefQVfNj1WtZaJK1qCdvC9gtGiOQyPJsVq10h
H+lU/IfdCR0LnadOxi2nlJasSI6pl56Xqx657KcDYgTyRm+6E9bbErtmu+DgVZKu+7SyXvyPu3pF
oU4hq8QY5aact5Z2FhLU/p9dj8099atPXXfssJJ3kmHOAXeriN4u1wdupQP9WNoKHvDgmvyiMoBC
BBdrxZNwU2gaQXER2pfO9xuvlxa6R0ZPrYPA+I/4Tpd7OKoStYA3DNFx8xSYRlw/wTsmAyujJ0K+
qO/pI2i/WQNsh99JQ8Bw4HNO+m+pRJ1auSyky/ubyAdrNGrqL/wirWoRd1si+I5zzejDBUm8WjvC
OOmHeNp/OIxV8V9nZWBFdpt+pP8JlfJU9hgx8cs3I9BxWxcVsiVcCYW9tQkUX1O7p/Td4QedBKwW
egtrwHISyK3fAM6v9QlYANZXF7XnWW7L4LrnmEBAK1CxEjplQW4EQgZgPLlGYspmLpqEYpTPpYuJ
3tLKuIhrzc1/z2kq5pcNG5INLFRO2yCMh0ZsGRmXxxet2O8zQ8lCGFMO2VUAKsXdUo7qKgBCqHeG
4R0p5iHnozP8Hbubx8cgpvW5CdYjIwcSKYDVYngZ7M1qc0dx35fjoXkN8CLgB+9MhY9DsFMkdpE2
fT0GsL7rFiEoaB5Zi3crrAiRtlFXY6AenD2/7SSYF3pQwhhV3NCPtBKqv4y7tnSuJrZ1aIpk9rsQ
VdA9gmAQqI2MFmi2GAdMpOnk69sefupn+IGZ4bTd4Cj40eC17YnuK4SpQcH6TVnWqxPqWCJpoyP5
HjEVTsups3UNeFgQd0dmJyqS8lQy8967tJEkNu75k9g2Jr6KFQQ69GVhL7jkNOVBCvTmo8TNToii
EbJsATyr/C9hC7Sh1tGdSuE7Q3+MPnFHDD4Xfaet+1tXiHAgMAYkIcXQZe+anuOc6SHl/Fm3yYU1
d3kvHb+N1w08uZsUun2HSggGAkkEoFiCzStTALCj81ZUTYwqHKkxFcB1wdQkBgtwU1NTs/+vF3gC
8I4HFcLfdPv0kNpj6GFwQYVx0wsPJ4L1d83l5z2lPGCAkTWSxqR6qMVs8XeqY4n0nNRvj7xdOPX5
SHD5SnKBZVUsWteviOfyA+wocPKmWzu9dsDD3tT6fI03He7/KpcK1X6dNNdTLXFQAhNejU5LRrh6
L14f8B4SfUSEqgH1S0SDZJbboV4O/NB+bpu+wG8EGn1FwEqWEU6vK19HiC8PAdOVS1CvDTG6ZBPw
h9bG0jiMKYsd0G/eko+Ial8qUO+8QUMW+njvQSzS/NQw4BdIeeZJa1pwE4GF1XNmA5V6c586OV5v
NUlsBp8rrItu/xynH/Isk8SYS6zxHlnQ0h+mdZyJejLTMh2QeizqqLWGf3xii4yS/F2MW9in+XFR
Za1guz813YLhKus5g4s+bkhv7eHCl8mHVivqtN0UCUhP9nXCeCQVPpsC1FSje0BdZzNeg8AaKqrw
os7vT7dGiQwuKNhLlVID6OHSY2W+Ar4HcmM5LkIRYZCtUwuWhgniTyPbgyxoTFMNv5BByuUdO/AN
4tuzVodgJHPejYpxS5Imh3oRdFRll/sBpa3GLZYy5SYILFfsHJ+7fC3iRTvAuZfNqMZgu8vQ0NLX
PJNvOC31enA+RpL0z425PJV8hyzCSEB/qwI5z62YhTZ2ZiO1EEZ9Y6t6Ev7AMLJhtIJ6klHX7AN9
uX1UQhKqQD1FIghYhxqSoeIyL9+6ypb5xQLmhkIBagORWEFHK7+sxUXnwBOTXerzaqPWdYZs8jEQ
0IML+aMa+0LQnYfpx4li534heeMuCBlZ/8cE85vAo29TLr9Z3mDjOCk/ADx4qM01NL5vr5XJJlg8
9mgAljFh/GX0kqniiaBJu/zxjeB3F2eSbOV1WBfC0eYZKbHf+rqWSel1ol5nqiMkfueEl04W6x89
MAYQoc50Rb90WEpQWJGMz/zGnXMQZMOW8mnRcueBlexiQzy0Au5P1719CYoYMb6m45x69LDpZXWF
Is1tfcl26CYYLcPakCaxBueOGq3qTe4rfYQ7iBfZgtJd6XNGAw6sefJgzBgRAbZeY0DfzIInlApx
eYka1hlUFdqbrLrMlvPH09ey1G5ZGaepJ/SF/kOeP75kSioo8V1hLSFiDlbC7lJ5gI8aw/9bFwgn
Ky5zTCqfel8p7iis7gNuVQV/pxmAtNtPj1/kNdsacxf84gYJCuHlS+UvTBzblBL2teSwM80x2Uv0
7OEbuvOqkeeBlhY01l9S6EWv5a5kOv8YRJhS4tti4+kG1cyRB17Vionaz9Lq0zsaGo+jlfkLuUUT
HhrTtApOic42c9AmGMf5z7EyH2IshnSjrsciKngGX7wS0m1A+SdG3v++SJdZT2yJggEISyq8M9xH
auHjgfw892SbUlxrbSut1dwba6JDepuXIZxbrhcgeTKYMMp9QSoBKVvrujhdBSEr02R3AdRwTo9s
2Ku/bHzUVxkm5urMc2m8RA7SLX1XHzE4PuEnTrmUb+0ebJdjOgrJqoAmifiGRiBqzUq+jIu2veAk
bjSPPQVXFZY/ZuwL0TlIfvPfuuBWpk8hI11wQvPzbtIvveRfu9BNdVP8uNmLTBXtrp2oh/G5FxLj
7LqkS0ydn5gXnSzVR+/tIRko9zDEBLu57OehyVKPPYDTDZy9W+npWJJfrUy3jqooHZXExu14cHrs
zh5K+7guxNiykGxChUw+0tkkBC63ApWW5/s24QR7Y/PBW5pPUFdR5oUDWUgQETIb2OnC7PSS7zb6
q2aCYE53f76uQv5Rlas32LwUbkjM42/QS9tTIhhTa9pTQOxhEwWuS45eTiLtibVrTDy+qoy4kfWs
H12xDcBthHWOsLKYw9eIdvThIugurao6L4d6z4vWzQGMV4xThCw+ckNzfpbAyylVltLSzRO11A2T
syXT9Uh7hMsDebnOKCLfVonx47jERAWHxpONEuwWDLrt0WMwGtQaosEgiZkGWF8izfoItdv0K+9t
chHGtk5KZOVWuPrURWWsHtlZ057Jhmk3lot0o3XTSg0sdny+dJGbO1Y0xfTElOGXj2ZX6XZzda8F
Rle4KhZMk7ggK7muytPQiiigNWqBz6eS5U4+VNfKR1dwbZJ/UbMfvvYUKLr9EIA9+qzYja5xU698
kP3ZVy7P8ruDuDG/qOpW6L90I5ibIP/GImAYRDUlpN4VlAHS2eCQx3wrMFrRv/rsi6buBVVyqkJy
6UthBkWAhuzvWhVulTjOSqD9NMaBk75doHGSbA9ZfXP4dxMhkNEsoSAi6HfUw9ETZ4kS3cMAAz1G
vF57My4uzYCIU575unpzyYMQ63NNZ3ZnLvp7zsARmconZPRoHIAXYbrbSX2MVxKsDSTsAwn+Tm2+
PzImyGP1IVoxXCt9SEJkND7nhTXIrw0Tf73BRqZxUj6poidc/vb4BEcKpBZtVZEAxVsYMCFksFaL
VGGKP2NNCQ1FfCrvd6MRLhQEtkXUhGA9HJsXN8NwJgOViTHmAS4IYpJjRJbHa7mIFY9CuwcROMWg
0b3h9dkGOUx4jVVxgPmddHJdBsHSZeefbNbNFrInW9QQIvJ309L6u5CbmdChNnry2zCCvWVurluF
hy/qCvcT/pB4eOypyU244QE9IsL+ZxakCt+Ds1n2vrwsO2YPh6uy8VhoHQXQUaqz9SdzhvQjv3Ic
aDlBN3j/yiP9XOwY5s4e+/1srutpAT+6KVKLrdex2YawubP1y8jGM3f/UsqmpZZMyv+pcR2hNOn9
BmrERNqMBhH3Za5CIoRr+PpAPtl38x1QbPXaGeq3vqHqT/WEKcEdEeHdPFpULPPxcTM2slmlfNrb
aRq7CBY8HA0EafM0p9vRn+YiXMfKFUUJ9DUr5idTxMiwvqUg4TEi6yJOmDXllyS8/SN4B656Kpv8
tP/eOP4+iO3a4Rg0zuCfYMGjcthSEmkmTw9wRRUqByaKH4dr4fDxhTts/6Bi444ChC6KbbN4a729
j4goOkhSUU6eiti1JbGX+wfuj54FnjjBWNWnT8EkW/IhnOAbJA6j+ZfR1Ywj0rNlGhhgjs8hMFyA
I71y1lQUL81f/jYHxFvABxWRsj+g2HDv/t6b+SJUOPRZDCSlal0NoRnq8q6nPkgGRAkq4cSg+/E4
eib7gYEMgvzLDYQ/kNrkliUK5bbFEMC/iJjwU69uWIGLG6ytcQ4Tklzzh+n/h+sq3bPaO+xhmWKF
y7MBnUaINZqfapcpaLtAhDRbSuSsX20/PVvdobyvAx6hJ2THESgN+kUmINoDLjiiZpvlHAYIUcoT
omJ+VmflopXProfvsNrmOt099uBwibOXOt6YymjP7p14kJKPSGiiwVF5rMx+XSiacaIvu1X487Sm
7vtWoYpx1svgt8Dnb+GgIEOpbt8Cm/LGuMfVNSaQBq0igQEswBrrWoPlhWGUo1jb52FkIBcaoQbV
6XMjhHCOjSrpCMCKSAfaCmiP75z2jRKUnEXVvQR61SzmdnXVik9hq4iN6QPDEaq/VzvmAO4YECbP
HkSMPwMzBsuRq6hUaC0hh63vmTOCF7NZO+r1F/iL+hm+8jKHwQL39fWJbLuTSESjM1V7L6xlah5a
TKp2SLUR8vnclx/5OansdAZAxDf9UG6l75uSq9urxgcZ3tInAfg9faMxoEejG463kwWRwoUfgc42
zeDTa0miWtK3nKCV9Tb5KIPpIGF2cSiGwvvyn3FW+SbPI27iAJDtXfm/kxoA8oMmIh8eNMV33ULq
eTP6skl1xPIrMsUbu0LSw8ipZtxjEG7Rn4SoHfEDLJLjtAGtg6f9U85niWSb9296LAiM0sGbmVXh
7WkWDLpt2HoXkIThZIGtvAoTQKWydjHjKESJLmfO6YEUBMf1zkWAA9mamh/xTjlDAKrIi2Dw3OKR
8sWhx8WagsFATTkli4F0RuH/GjGMI5iH6a1d35VFjE2BK1eOYdpy5GvT3XlvdwEwsct1q4LAFpbL
J86ZjOh/tUMuXAtxC4hDrKrR3RQnJ//yJt74vCeKeFaFiRz9Z3ia/SXs2WdBGJG2AZKM1xgqLq6D
GchgwZLjeXa7hFL0oBAC5bgmztZ1KlFR0FWYKCDouOjLl+K84tEK2WnBTQ1raJMjgm52pEznnbLt
BKDobFTp7UbGGYB+xsJRpEnqSw9yI29RzaqIUuMV2N728DhTuPKsDlXymGfMW2XqNSa4Kl3BmhW6
s2CMUMJ8OAXfNntAzXFy4ssnHTIwl5LHsoDdFbAaJkGrvvabsoldHX8ARiMwdF9nALqZknfiWK3x
Ax4eH/gxLN7rvZNFumnZv3Fa8p2VQnjkLQoim3M2CoVBRGoxgi9kG8x6y7R5YCPBBahbeP4XDCTN
N5M6OXn5gpyx7uANiLrSOqs/cSDViH1Tl5lFL0rTss2mAVY52DgCwNt2cO605JqPcjSi15Zj+UpR
G8ZNvQlG0P6zDuOzxwc+gs09KSbDvMuu7acDzHxnWK3KE/nd0hGmzxEZLtDgneNj5WR/Vl4KOsxk
idsVlfkvJgGqLUcRM+kaSm2zzLc0GQcU0Oles+ZHK3J3iKGU6IUWHau2FwrBC7N5z84a1jjKsUMm
bOVUNz8SHawkDNw2/0FZrw5xLdj9UbEsn77wMbnKd57rXiaHQ9R0hkWYEhU0oWqeiYYkbgNj3M7g
TGLeMkADU2+okiZk3ZnKNsVaq8+6z3MAJ0RU8Hf2/PBUJzsDOlr/20oMOHZxK47r70UnXiOxK6Dd
gQ9afSfd67T85BSQARMGtZe6hnXrK1/qSaB3/eUm5Nrxbz0b0+xis9fjt38YZXc8dazDFt1OJJ/3
vf2oaq+yHQl5fL7+TYJ9Pye5aGt7hcDvwNMj9txLIvpdRkaSAZUbI3Tbep8F/HUfdUx9zBssJj/p
b88k/tSIJ4tY7BMMkH42IEdKt/TtYpsPbqnUNSjXVE1Ywn6T4EKBn49+/dOgy2WlF5VI+D5wOznh
nbOqOEwzVYmTdW9+s7Ryb3SeLOGWZFSylyDjeKfayDz7tx49uhQRF/fhK9aoZVDEbdJIi2KmP4Ef
hvrgyBLLfotilbqoXuHZLNllSQKBPbFGs1jTv367IU90Azy/jAaOWBkn7AYKQhoFEPPCcZUTWj3h
x0opMelvYDVU2YmM3Ge4kSjlIJn9hXhgedIhPs87vWw1fdCEXwnbLzBvIpJkvJvgu2/R3RMIwViv
W/haKOMW1CRAa+XyXskQ5n2/alxFcGe3B4IM7SleRGnfiC16WX1C5GZN98VpGHtAmjcQxcz3FNQS
cQ7FdYvNhn11dsbJb5AQOlpscloCfiQS0pRi7+8tbpg8UiWmMAx7/R6yKV+Kc0DDeoCY0O2dRVYK
mC6+DaLN6ewe/LW+yHvNtJlExjw4XnWcFJ1cH8GMPKOYiSCzjPq0djI22SfXka59Dr4aGcKCbfoQ
wScEgd4BgRKO87J3vx6sEQMjkZq0Jb6Cjt1kspEYKljah99YTVAyKcRayhLbjslMhq6Z5oUCBGJR
/6ooq/nbuZ/UHguLRZCGl9s2iHQVlURb/Z1OtuZNNvym4v3A2fwyjiyB9HD/2Dz/TlrfdcsgVgQG
d22QAxKoSYuKCE/C5TWYDHrmLHjyRWEiybNMILzVVmzWKysKBwjxH8U7rUXMCm0NFzKvLBdS037A
Qpl5xHn22RHXwF8Hz4gvy1GHBl4ty6nlsYFvqQq6sJA+vNOYSyWH0vYDdy+rAf4hjWdc2WjqcxuK
Fi4G9DCdFicOPoUAMjxSJw37XOIbuf+mIpl9rITuryXPV3cIsm3owTX3GTU5kVWLp1SVZSqlgx9Z
rM85mb8b6iON1ogzqeXed6AMEd4U/FRun5h98D7EHfMq5IlZXTl2TyacInRm4oM113wIpFlezYuI
xn0tmg1gAL+3h7r4bvJd6AAZsQhJs7FKbwQK+H9T4JDmnwWjpZ0aOb4DiHlDjqm15r0JX8/4h518
L43yTWHQEPiu5TaAug6RVe1AYalyKvwQLlGiOnwqFK85h2IOnuS+VrXjLjzq/Oy9NF4cX3BvpVhx
88z3fxLLqaqSOY0odK+bPod0pzZtW6MK7CYmKz8tQn3GPDLDn9ZldQSbZsxRGM0Yp3juMyoNK42f
t4Mf/MoTln8G87o9qK8PO7CZvN7qQCbz+YtSTYn5TW0SRtve3ySEl3WHs7raO26C8qp/+/2bGHTp
7axNQ5GQOGPN9XmZNMIK4PG3UQsQ4sZGqGPyeZfr4x9hTLiTSj4dS00l45BKjgKCmXi6Pg9J9A8k
P50g98Q1a9cns9Tl0xxuGrKzWEZRzBt6kzgDGeZKtuGLr31T7CCd9zUMg6TRHdBYgDKmVQvkWUr9
7YZMiTby3FVCSk7mF+/d1Ri3RhVUSUY2aPeZanPeyYjHO0Yl2p7wj82xstQWIcTjI4yehUauG2gF
dwLm22CNZAO3zVE9hG2a4ipvlFqb7XcAbSCLq3HwcE+agISJ5L4jSMIA9c2udp86KdeHJ/z09QBC
y794rkDqqd5bjVoN2v3o/jWvRtQvsSFWQ9bfy2NLAg4p/4bB9vQN7CV8o3HwEtfjY1JBOfsZMPJf
S+gp2e2xU1lc4Ct7lD1ZiAioEjLGZATdAYqK3TQzcV8GSYO39mtirvQMGqFEtABJauuVqyKX2/5i
tusfuTWFR8u66pEefNdhxe/3gM0gCmxsIsredubKDGR/YY9isb/XA3xEuwHSuCNaoKi+c/0ntqBm
1bLkZw9J4k5y2eZXGM7gsO1DhKKcZzYQQ8cPUfsE50J94EN8me6IQQJHg3jYBEghmbVQDnZ6kK9B
dm9OZ+wNhkXEs06jfXJsspf/kTdVH5Pk65mbWSbfqcF2wUB2RXEfzC3ScFo0Mp4fpZDJXxOIqwDZ
ypzC80t+9mltaEsWqRO4JVgLGV1r/vBofSH3Ca4Hft0I5lCi1DtsV5OKWUVC/ECbXNAmprO8HnXo
gfC8yHqX8do8IruMfZmUrPnUAzOQ7WKBY2QdAkGwNSa6MAEXT86wSbsSov/wYAG4ZLhDKPxWuGhk
MrSgbUysA7bBRAm9eQZhQgNw2S/iwe0gpkQ3Ho5Gcas6PUZm3bx7yiZpxz62y9mzvXnU8wnJAOKw
MavTLidwkJXVgpTXaM4ZC3QF6g6/Cg5au32udpfShlnkvRaTaECkqM51FO8WfVN3BnwuZ/WQ4XjY
kxJITtuckCRsK+F82RCeVePqTu0iouuxMqEnIl/VE8vD6//qGQVRpppaphBsml10R5ETJJ/PayAu
1PX6y1LjAOLIqiCjncut+XfnpDLfb9n4TLK7UvWeZLxEJ6IJRTV49RyIdfxEE1h5qOZWcgJgkCb8
czpG0tgzRFdX0578iCqQT3xsJjMnG6ytTwqYLJcHrnGMvR55GEOBvwZ61Gfgm5pRDDj35MoAiAJ1
q91KBQyJbuFQxkSeMJPkyWwnBK9/OXS7ulPLPEtjHA5p9sylTHeapvO86hE7BppeWyRohrjyMGvO
S6tmEZN+ITIvt1+j3QnAr51aG9goP60qUDc3VyCF6C8g6TS3c86s5VKFKfgAoilDIxyV71YXqEE+
m9n98NbjCu6HvhCIccdjaZ5dok7rHZxrjiP16FWq/Fi+yUKpJ92y0dJRfDwp+6jQBoO/djdifFfc
LmnxP8Nhyp2OkLsZVNONlx+8cdComdOwUwZQ3sKjFOFLb9pPwK+lRk6HmYTHez+ujtmXUWZxkTWX
333MHD5D/iKw9AKZm9PprtBlD/Y04m4/Ym0oiHL9shDVZrxkyFjrEr85TMMB7QF6UFBGYj9qp+bY
c3fdIHpqVzl2xaZeA9tX7rYYBU6dzYKlzxw8SrV+ZVtvAPLe9IsCbHr9tng30QfSUc3NTbsgZm+y
Kn/yyHi08aFqBp5mOQctVrKF78MHXMcCh+AggPCdM70uTp2IEy23YnvSx8l+etDLzHroWW1OaJon
RiBAvuniREy4YuFNGK9qRnlgqAfHBeY0USk6fIImOVEEtMBABcPCE7BXrRYrvxNU7h//8JgtbQHk
UsZIR/ardrSKy94W06Vt5K5xk1SxyDJgzV/mXlqWnPNQ7UDbMXN6QZrD/NlyFzuZn0WdMi9i58N4
LVnbgEdxP869WMpob5uIx81Mf+0N2SKkSe9NgywaCL0NCiOPhSV7Td6igyNWAXP1dDVqNeVUUgd+
F5YBgwQ7tT6BSuJ3dmY/SFyMEOL/o5k/CluiQBxwusIVv0yDh4jrZaHZyh95g6ph1zecsjCyXqsH
qMPRH3DQ0MucIGLENC5X7GmDMV/RrHabQTiy+hRbSuWkUkpDLOMb/HaET7IwzLpCADkGBvDpnjmJ
N6SlbZGQB/HpUY8Ywg063vYwSfzahUIhDhqtctxoVjbs6fpb/KoT+8o6VkmfrhYgwm+PSdiwC7zL
2+aV74ScH+NIsMWJzLb89ZoD9E9LXAOSBCZ/0d0a5h4YIDe5fMDW3/kfLApo+CRrSfHxal7c2I70
6WDz1Lvodxyvo6zS8tO468kFABxY/vGfEQDcvHxj6LaxBrV0/wjqsLv4mCfRPs0i0BehDlVXJNCw
NfS2wJnCymod9UhxMAIjCiYdt8w6lXzwPrsNYApjGq63+zj61b7R2T6J2hb8Uvt91NTxkGKDzSpW
4LFMU39fFxAKPAQiM6TQ5LogUJW3cddqXyfkZtZcoivhLvhL2DrDW6W5RZnxIPd1SYLR4hNXTSAg
NGN4mErDcPxNTbWEeQCgiSw2G+bp+YjTtvaPfXfTT6X4h9fKLAYQrR3SDdU2sAGeIGfjt65QlMsw
A7/ZdftpV7O4D1h3mJr2WD69rTAmNscg29iVwiqG5w+74wZwnV/1CCNbK7L/mbJpznZDpNMNac1h
kpVvbd1lUrQo4XdmDUnaqdmbG2J7S/3ZvIzozOymfFYDu1jzfNe+CjGQRI7+aWII7vxqNbR/gU4k
BRRFWRZ90nSls1iH03UV5q1Shba9gVa0CgbnLq08G5qOzZRN6w+RKHGkVHbJ25WZF+0xiji5X/bV
0I4f2g+90wkMHSqHR4paWDH1UOdmfl0UWTLzDQVO/Mtb8RXMIhC6P2IOD7SdVeZZi9TNpMjDMpI/
nojAeulqQu0TSR0cnpi9Wf5haRQvHR1Lx6psXE7gu426Z6OIEp4qhkJ8/4e4EQMdHDYZK6rTLuMF
XBNgISn2RqKkPmoUBCqPApP51/wIXtml0fO21WOmS2rWs7YFBzuYC/RDmCJ1tlA8KMdxmNa6+U5i
01ltLvMIONT9nzQJS2rINrwgcPopIPY4IEuWE2Shw3YKWVgTDi/Q8512BecXqP3Kucedb+dvc7Zr
rnFynfBuk6XiBSa4EJ3AsOU8J08AkArmzrsBNXEQP5h742tDSQLCLoLOJBu4mDO3F52gDGR6qKZL
B06qpcG4ETFcg8gaEq2zK/MpjQh4oxKMtgosfK/UrzaY2GtN44SJJzOHIRirCiKWhYbUlNoljqHt
sJ+2xtIibkkafdYSAmvgJi85dWzR9W+lpG3sddx2E6yw8J9YX4+BvMrCeuBsCjoDpBX9bCnvVRr6
HaDPyhbbzU+udMdR3P6ZNGfw/tvSSa5nPnm3ZKRaYWL0qn/EjnlGwJhff/Vb3wJb4ERfD3OHh1SA
JzweND77zn1umOP3gTsRyGUIcgp8fLEi96n61TEyBk/hO7QdYWixXkLShjYAK/QSDSVwoM2SZjl3
HxmRJViclnNy2x70AN3VgqaXG3Blq5rlgzuYM9mIddO401RoXM5o/7SrZnsg1V7ZRAjeLUT7zq+e
IEGPAFcb3AC6DvteuSi4OXrTIG5pf0YMtmPt3uvQkLwCUmuf4tNwyG/S25UStJAbJVrbN2qZmRBO
vjWFh+69cgKunbJa8qLJLueeGFo6FiLyzUP+Pic9L0jpevWsdZb+zFscxQgzaAc93vHjMDiQjhfi
ec4PMIT32Iq4GRPUBw+OW5cqS6wxpMyanhVLzCVyOSsxWTzynKWEE1JGp0JuA4TohxlkMDnz0gQJ
wnWDdRd2YihohERmy7Hprk4GnlV5PWvjyIytq13aBAPZdqd23aKE63ga3Q9UBVLiAU6SQMYH5hf9
Yy0dB8K6dOss9d8/BlFS6JXFOIF+cpIaOvoq/Fb0eXhCGdCN2fe2p86iw/KIhYgx4TnWNnznL5zJ
egmG6cT2iVTmqG3atL9JwBfEGnJX3QOLdR3FcTlJsgqHXzf/WHWHHny55qP+ikxHfgyzbqDiyPMb
QltCLT8rN4ergJBCoDGazamDPWjBCvKZ2zA7TmtuZaUQFH3885eFRLPDallrmxhY8YRVdYTqAuRw
07KKTASWbqZy2bjA7PZ2cVSAa5DAgbBdSKL9xebZDjdWQ3L2GGcsndqXWq8wmBEKd0WdArD6mxvT
1loH0vMjbRMAMCUW2hidyE1RMHm/BisdaDtLWam8U9RYDY59X4zrs7MlIvRrCgCAITHQDsexFSrD
9IlSWH/j9oGrWcW9ESZ+SX3Q5IVZSllS+Hk4L4DbvacZdb9/zgC8/H77tQetgS9HXj4xdalKxwtb
4mJ8D4UHyEoCrEfj56P+ISs37jrAWHAhsda7xqrdjU9aCGHzUP7NfZyRajn7uN0T7l7/hflaW61J
Fx6P5pKPWkQA++o+z24GClvIcqBOpx6PobElbcLH6PYn0jXgsX5Emj9ZkhRK4FOpDijDV/JDOYlH
Ix22cpavFVzdhMP7PFis/p8Lh9WNr5QhjB7KMcWWLq2GBUBC7WrZpmq/eXYjBpEdejfdeNL4pzcB
uHK6xMRNzw8wBZOX9nACGiFxu6LspqdWlhYcmP8iGTVPgkUwC0kuXjjvBCoD5WOb0Dy/zTfsUCuk
fKTVjPKGplFNlagLZDQMMV1Bt4nnfEel8fyECgllA+/gOdqq5HpGIFvJMQPFHHLphpgoHj+KUB5j
ZZTSBu9Au4jzIlKU3Q2tLq5siJAFZ1gbemyoMJKAIdn7j0vrUkB9Way2hgzcAJa8KH/mKizUfrDn
rszQ5X9QCwZWsMa522RMMNTafBLE+iDivgkqMPJnxcpWRmkMk//IlvSKuKHXumGTOxRNan0gkHke
xlR7UuTQDp+07L5v1zi9rhMsaO8/X1q33WNXO7NQYlhbngjy1ePnOcp8DP7jClihB+K3ShQ4OEAA
ZZo4Cv71iFikFRfI7+x+CjK3YBeg1tsNPVfcfpepsD23kNnC9ePGbswGHjxICON16rxUpHNtTrsA
TDbXzBeYAiOobF787GZ1LYrLJk1DT0EKUcWw6djrkJkiL2fEUudSwjd6RUkemly5hwVNKuOrIxip
43kO/lY0NTettIC32oFRe3yEK5W/4xUJWelgyJFXE/sBKUIPsB3Y77WqGpIi+eZt8miEiebuwrWE
+luseS/UqZ9OF2CCNIHfIkvNmVVzGo9EQGKfuZF4yCLIgiNtalZEq9xzlfBUhKOozDqZnXkQdW5O
wq3J34mbw/RT21Na7PDOn+cgsBabOBfs28HkAgZD0ioKlWOZC4E2ARcJmnV3qsR4gQuM3Y2XfttZ
gIPW3KlgdGxw4veV5307kifmf4B27yz3xeY71RixRAT2MEMGAPmrh3OmEU3qrMKRXho1M/ED+D86
ouhuTfk76+JXdM89dfOJ2Uadi5iPrNioSrhcLARYvg9IK2qlNtWRpRmRgA2J4iyPXhM1qt+5ZEkP
EFZew31gtKKhzl214j9GK5g35g2ZfBigmvjgUtrEQPygXr0QjrThhGWlLk3iC5v+fdyJ41KCGypw
AsQVbEaTKZlrNPRsXC1Q2sShaIidl36L6UM6+dBrSRA/vhTohMDTGpLSR+xKtOe9zJc9n7Mslbin
glPmxfIS7jxmYtoykLX5mJYdi/d3LiZUZWE/biYTmooM7OKpk/7tYpXXuQBqNP6mopipzXHAObX4
eFlAdg0XPoEcb7eCRLeZa3TBiDLqIm90VsHPW5VPgnFAK29JrCH+W6Zr2CBRWKmNGRp4FLfgan8w
R9soYkA6re36E4VthmEQCNQ2QyucKWNTWvU1pkPac7ihy/NiFajgbCZ8PkeGbYSLDxDDyybMMqg0
CtpQKcdvTcu61nCVK6Zf84fgOF3LsVxjVG3UYbVSZ5jxMSugFrFKegIBDIXKuGBcM7J0FGta2RQg
t4kCUkS+rQI4VzgwuxPdSNVwCFts8+qyxj+KLfEAxGuAT0Ojptwin8uGMa1tavHm421OmvrnQPHb
FRFlOYtQybfxDth0u9PgH848SAhCm0ZlH75IKcjI/MP6GR9BsEbNEY5Z1c0jQBr2EbqarqRu0EIx
jY6PNzfW5GEg9TjP+WQ3AUNe/KdS5aMz5D1z0bnFGNspn8UyARotE33kMhyss35fuzFUz0ea6Dp0
dp/0+5972Dzlcmbj5WgJmPC0NYscwoyHHh/Ar6PDIeGLvsf37aNa05rHXFOjztJO125tEl2TitXa
NOTu+AfLo6JKoHHW8cOqFt+/6DAEKFMJHDmHiBDQxfpFgDWjXPMyhM3MLPzrhzvQ11y3EpkBPf/x
6ZSHDYtCWlURUIafFINfST+JEid2Gu/Y+TuGpIY+8en5Xd9Wkp79aZxM1HOp/MQVeve8r8mcyY8J
4aeIwqSrptSfTUYtuVTLbNfOUGTw6E9yApx1afs6PkHVbXOTRUFqY1OF094/zOHLqFmkpR/eyMMp
PjutTrqeXbx1CnD0j26ZrCiixxoSqnHKx2mZFIuZqyBSIoW06GvwKmAcacKqkqvxTwh+XjVaz2E3
kWojBIwuFkC2Koc0rnbS9/LPrNtFz73VWoBZtFEK3HR9TfKJxcOtWezPw4z+9Ps4jhEXKHfZPAkc
xjUKd/88PXDQvbk6bqfmTsmgE3YHBnfOHrvFGAAckrIOnYB5MHuy/vp4gU9S7lpi/8SEy27CPsj0
g8AJcVEq5MrKyFT3GP6PAlSuRVkTSwkvhX7aXYs6F16lN0Q5+2bj7rBWVmIa9h2btzPjSJpvKMPK
viAnFMWhCfung7bOi46tXhOVW4OGXyV3oQNHtWmFvBF6HWQamyDRhnWMrE9xpE2FZyrxq3VoE41J
yGBskvjR0qdrEm5TvX6euXiMFp1Ej2dKgDCYWGIwSHo3BVXzoC3sniLkE9BVfkfaCe30cFdIlZVQ
4TaYCHqSp6/H/pn2XjybUTILkZarJi7lf7iZ1lT6gOpzjz0dV3HS2v1F3rd0ofpUdBaLZK+BmSlk
Qp2kwJjzXYrUTRe9yFH16r4FibHCigtI1k7g4y7o3ZrQkjfS0QRDUBa5yF57rQ6owsmzHOkf1vNA
HqopUDUkXmM8HPOOXv4KmtXF9JAiXYWSws1M5vyw/j5lbc/afgD5InVsjUAkGGmpRBPtOHAnzzlx
RU2MCsY7lNHaXMgHUulQw9FF9HX51MuEHBr7Nw6W7epAjOb3IfcrmfsU6X+itVCkKJ0IiHNJc5IW
ornkTkPUmrFOWQ7vB3UlriMBZyGRTvOBBDefR06PucVXaHDSkghlDEAs4VZJKpHH7d3Vl38b/BeE
qZZs8mbrm4v8c5ann9d00JVyQVG80fjzagkxI7fhjv/TiTdoN4373oDbqpgnEN+WPiWAxgs2c3I7
sjVpPJ+MueoSdWHYd5lXmk9NODmVqL7JDZ+RwLkk72O7Drqna3lsen1+J7Td8pX1dcxUDGAJAGRr
tyv+Clb8zm6Vu1tQejWlT139MMRRAkmGT4U+XvtzNMrNizSIZrMcxKr7O65CfuApMm8cuj2b0RCU
BSC4Ms8kipnrvgKEUZtHIyHvpJmr+6dgVMCZ3YqLmTPxUM+D/p0x46gH4EZNKFO6NF2ITvyFtJGd
hORnaa7rSXDbf+yjze+N1SGRD1zB+xJZE4eIWLc7rZy0pVhPOGx2EAP/oMvZQTbDQSAHnpGemSyK
K1m8t7depAvfrHInAViEA6wQcKvYpYgOByzY2gwvLrFTcQuAV2/Uh4mM/c+jspwu6TilBCW2h5y5
DvQu+Bu34FGyQlrClEVMDb3UTwIG1gF7FShQd/pCksbCNnuoLLOXbGZsn9w3S3uvD45NBKxPi6gk
GK/RTW+CYCGVUCnTXD/1IEPv1QvifF1YU4Mfimys+SWnryM2ciUlhodRJy6xgfS9zVloz3hn4b3n
LaNzULBXhY6Wvm95PEt31Vk/Wo/P+3NEYCdoxYNTSNMgMy+luoh3CydfOrRDu5g1al4b5/9HceTN
YRFBDnjafhAugMSmB2eD3jkqqDFaggJWrHZI0Aseq9akUBCRaoQTdx0YjZQrkP8LsolPaL1ywpQf
MtVXLo88GM4vACFTWae2hxCyuQKmZDdSQVbbpMWl9bW0i2xFDLqLi3iv8KUBjpNxYCZYqolmQ9LS
JD8MTBtLMEzx7vCALlqCicECeJ2N/dFgcPN0eiCABFcrahFaoAlXBQkiMEh8fS5TNJ62OkhWQ6Eu
8DCW79pOZtUqfJEVCdeYBZ/XBgSVOYlqXq8OjB5uE0ZJH1Zq1h65A4vAtVPos+6SgMTjIdtegPPp
m/clGaXws9qv3wCtxy8gYRFxYBk2eWEIz2WfkotRL0XFKNVpYgn8Ix00pUAHnvmQA+GUkt02Gm5T
ENcYz1kJo58Jo15CVwhmjwOeD7+s6P6BS7uh2iqGAaolbvf5vdU0/aw7CGKTaPHIPirOBtay2KZF
yF4Lob926zlmTVWb35d7d8pK5/Dc5l9nYwtkrBXPJvpqL+3kS01bw3oY/niKVeFDlynRyWLbpX29
evGY22MawswQtXz4+CmwKW3dcHu0m6/Ss45BrXuK5PjxC9W3cuvEehSp/3MQPv5+kt9ePiMzJ3Gi
eAj48hDfLUnnvwv74gAAKJiJDvE9y2YqtwDTahrEgl/bTTt+RKEAbgJ8mz7eZJTQUXtHb6UXOHL1
66YSlpoG1n/VHR5BfgxPBlwbS1nFDMwyiyZRCKI8Pk0fW5YTRYXS/5SToLXtxq90M5PtHCQfYny2
jR3PVyw+LdZ47S2ueKDKt+D/My63NYG+noC0xREhqOZw3zJZl9eBwdGu70YgZ1DHUJkdowJPJG8G
jFPW4Mx3sttg9gE2EzPEMKv6y1FMzqFIQ88XulV5Meg/FcqIuCU8dDmCuW00TC/UZK6QWuLgq3w2
saH8BvMclQQvt885H/8/kUgF3Ovu5sJSlw2372WGEt2vBwEXzStD4miRCScJrxNWBnGy1uWg561j
tAZEpx9yBqz3oE5CYkmEsu6Km60Zj1FjxshZsgmzXbNQ6sej4NpVdjWtHh5eFxyB2uMtbiGWIp//
A38mylff1msri6VxkVCmigYQkuwhVxuKmv8E1jyHM7mkgWC7lteGmGa4z1IlfKFG3dk0bOqyiESY
Jc+0aWuL/rKFn2Oe3U43mKYwYnnMEFE03mRc6fuAocaABjklnanAzupw00w5PTZhbHy1Z2h6PSsJ
dRFEzPpNP46jX6+bujgp2fC6Y6M90TvP7NSfr+fetHpKPWIfPoIEeESQ997mJtJM7haVrrHKsJUh
YwDW0FqyA2ZIQ5zjWvd/u4TMlk6z+/+oGV/SlgNWycFyqKFmhaV0HjbvEuZEcFGiHFsAv9VYhHvU
cwF/XLZJ9JctFJ/J0ERioQhhLmif/SYdAew8/5JrH4/HrTHujUSHH3x3pcnvUOAWVShYSGxbbmg9
wzljEMDJQBmvPJ8JQUmRA089sJmBw/l4pGopKOAfZG0JxQMF1ekXnxuVPqe9ORluGwNmcZJkZo4V
jMCzXLHjzgSXKBuiYuAVLukd1L/ow7n6mC8kV+NHPbJuHKhsiV1hP8atMw0wJRDL6GgSi9wHgENr
chbyYF5PBeaHPxkK+zXbRhzle41o7W6uWQ8Ea5iQ+XWlngpZYPQ13PIGMUN5ezeduRazqe9GS0SU
M4g69OZeES1kpvqaYWxxp/uPinB7J05QDzWD70BIwtkh4vnPDLhLdb8zpdqd1dqlfbQ6kRsEXb2X
JrmAxxHT/+tUmsBzvlhMTS9U/tkWVmRWqEgHbcY7FSTouUUiCstayqbgifqzrgqCHNJLMgwR3Uoe
NacOsIr0b06NuIItpLUMdEmilU0+CTBvol7l/K4UPSpO5/eUtU/jrUQHod4NZDmDWh2KtT8iqiu0
D6NmRKvATx1A+kPMg33/yq6eHOoyCC+6G/jKPCUKVWAIo0okh1/KZN+3kFdvvnsD23b49A5h5gwn
noKrmwRHO8DAANbhjWBA2qIvqo4gwdK4N+377zI+Qbwkw2mKXpjTRODR9XPqR/YjduVQXLAnx8Wu
njfGTLwMPmMonPknpIAVOgqBFQ2tEFomyYvM4Y4rv0Fp3M98TRL6ZxpzJ6cFcMzTcbTkfAzIINBW
crItT2PnWvD/QRVlvnbc5wZnxvKlpnhDGuMefT9j7fJsXFu9eIr8KCh+24VqncCvqxzEUqnX8XC0
DdWEujUhuNdlRVAWoVd8IXaBIFOA8JyLNUPkFrN3WiLCmNtPuhQRy6a9PH8W3WdAAKtbYs6+Ki8t
nnJdpsz+FTWJSbWdgoWfhe3RWw0PrbaOH3EwdzXYz5Kk955WPNK1HwXFVMlWUIKpek9PfGYBENWk
6Tb1bPfV15GT0/5gvlcym/TKdt3h7WZpKLxsQhd+9J5KlqA0ENGVUCFwvcML8KeVio204f4nQP2H
6m8VjFITypQMVpAgsSuixiX3WwgZVJlSlWMzCF4pHltgcJkdaNh2E/rUpDpQmE+/kThvXk1HiCJ5
+gWlGjteM9LZhpX8qY0PuliCCWQsdSVUc8O6CwZ1tPrSuyS5YCzbO2gPLTrBERHHmu4UbeiAwmM1
7l6cJ6n2UzAVu/cFCG/iUv30Oh1iK5DAE4idQWsMGMhJKfXiYBWa7VT6JSzs5Lc6Z/0CiFqdFkq1
uYI3xv7tGH7ogSAQObKTb/GlQgvusbh01aU+K3PGJf7swR6Z1qoUb3YTwGzHd6m8m0dRzXJnLfvj
9tpUQ8CVbcGA2HihqtmRqtuP6UeIped24iUVD0wy36auOmDXzk30m++rz/guH8STsrQGhjNcAHm0
Txt8R3/ZEHEsICWF3JenlOWduHr4w4FqEcjd7GzfVChW/UY2K8aFsC/J9I/AyPV5OAnKc5oImEh3
3FkpAKtyUdKfydevbUO/Sd96m9kuvfZgoVRGu85QVCwQDIA35MBcDixePZT4cD4eQkOmOVciZbiR
jfKqFUOPg6Kc/HJtfJKPICGY4TVWizUWmop73DxVETWTaQCTbbgc8TIftt/iCQJjudptf45zKoK7
Q6bnZs1ftEvEVqc9K/hZVY2DHk3977j1vQSVPrgTpNCuh1cpQc51zfYMGp6Ses7RFi0fhAm/BXRx
a7tsXny9INjP+Wq5drFgN5O3ZKh3OFG2X+MMlMSPuA7DLMPzBDmogbbvx7g972pScgVECx9kml+0
Cb/IOh55Nq3q4vOy7AoGZaaSC+Tv6mvEsHV6DI+Rw+szsG6N6RAah8oDuLkrdRJbJ5+awiR4zwG8
RBCKfi79KqbU+HUVhJHABy7jyhNpRDJTzwWKltQauZ+ml+7BrZdLFaq0bcMJ8fkFXdcoDIGzJ+oc
+qPe7RCehl1Pi3E/AQow2Ea9AXk4x3XYgGZdaU0CFAClo07sBZx0FZJbPlmsZxSn37K31+qViqiJ
Vho1qFawx0Yu6Ov3LDAfRlPPjLjRNfJp4LDZut0U1d/OQUkH8FtvB+CUuRKJ4j/whSeADa58TMko
ItXa2iP7FsjUqlWPfUSmQx54dyAKD4T5W/+1sGn4XI0t7gHQpsEwwvpsxktaFcpVosyGopDMTFoB
RKqYjylArHiJmsLNHchYOoSctZew68FOzeHXDx3Tn4NyFZYiWugF6dUjw6U4ttaMZPHag9BWRNoU
SOHJzwIzsVuoVXH0Ebs4bnK1OS847wPR/nTbKHSkzM2Zqhb4+93JgxhynOLzV7K0ut0XQ/3eSqHf
vHp+PxLxgtKprMu3zlETquMEx1tQ/kaGD/WvpwpdU+MzaoNtIZctHXWwQR7Djcab8h/b0xa8OVF6
qc/r4dv7oeZPWAmG+IF3gpYxLQ1mwUIg2FT0kTFusUzjBRapqSOKc0z1KYS3DanX33TdCtGi1JWz
r6W5gKDMxb5S5E3XXWX8BIDCGLrfIcF/m5a3VWQ+jXVeP2SOwf3hEGm3IgOue/RtgZa4UHfycFek
rBVImWgnaE95D+/1xpFR5gNM2goMYvuHvnK2pDqfyeR7J+xl0t9+j//RaJDpjiDOUeZbQHbTfKI4
N8K3VeyV6qALVMnAzgS+DbfJHcipipqVZTaDwq69uKRedLlVdhnHWodajfjiWdF90FZ5diYvJUqa
ddaCcBJvVvcww94idbSDu+kucLjhiJidxV9QvFchBzprgV+8His9vMPSdXkOeOglE+eMu00e8qfT
l7jV2GkUNqPKaKDeORcapUKsjnlmY9ogSA2NvZLEDwRnxAQgo59MZx1dm2q+9Euu9WKU0SwCpgU+
+73tKwbEPLxk45a9Ct1PeWQrplhNNi2DNTUfLgsgylME2CNnDgPaAZP27rlzb3AdKHT2hK8d49nH
ZnvEm8vC35tDcQ+TWHoUb2CP4qIKvuDFpYnIIXVGf0jWiixZki3FArh/MvJ9PLQB54gAHEj5YnTj
+8XKqtDPY+boG/NOeXh7fhAbhRvMPxtzYwdTPZsh89TzBwpXkfrxcaC+YZz5sGuxO8ERVoLEEsQl
ZtQ4jc+wQOTYKAiNai48C+Nv/zxnP5Z1IOPYJnCSB+/S1K4wyq2tKmF6KOfj3APEWybETTCU11OV
n8eWflKGFCZjakOoC3gXKiZ70k9Lox77C0D9hlddL2abqGB5h60eIhaZWmJ7ZPsdHrF5deUJfCLk
+/F/NM5vR8KtUxf2t1CSgYb3lLruC2jsX795DmgPbDjEhtkWDfTPEQ+OtCBorHqG6Ia4WVM3wkbf
fXI1lrFyMlNlgC7qT6xmDcjqRi71aG88JkNQituJu4aLrTwtOvoSxLahOLfOvvnQQr39b6Ie5PoK
Tm3A91jH0hHoPJS0uyM2hXVwFDJVvTB48YUyfxX/iHqmYVKw51EEKiHKFETlXyzyzYI9CfHGaLG9
qbcpgZ4nvUxHRykvdwU/C5goEftNBOmLSB2umN1t9Qrpv4eYtYbXMVRFajMqcgkHoTu4zj4G/aFO
9nbq2XVsMv1n/pTmg1q254HeYcbJI0hbsbzLaMG5OvCuJ2hBDOs8LYhRsfl2QVZyv+XraK9iIpyg
XNtxPWOOh7m/OnYEQReZ0PVg0mOdNGm0ud9SS9AQwa8J0XAJBQ0a+SAG36r3JOL9+clIxfbsHV2a
vk1jO5mPx5uOM9Tf9iSmrbShWzkyCrMifdk3+413bCjJZM3LS33ebedFEvklxe4ksFuy5JOA2C0t
obAk9t8XHx7miP2qcISDezlfXfsPgKEOovk9VP5gE2TDL/XDa70dIoeE3TR+i8Jb8v69vrz1yIxv
4Lzirui9lMoCG6FV26i+rgGIx7k+s3ac5/jBXyJWcYB/kcFerpWh5lLkPtlhgKE8jo9qw2k43anG
W57rEfbbOr3FTaQcl/SfHy9bgQ+O9GxtmxQlT8xaBlKUE2ZnxaxybWp8g/R8Cbj2i5GuGBrmpQVj
jXF+8q2axpV4CuIwYm8y1QxBqzXE4DJSXC7D5dJfRXiDx4btl7PlJkUDRAGcXJYDZ4SuDVFbU4yL
KKxe6AWS8GnsBcd+ZJESPg/7ODpvHqrJSqnlHIqVaHT1am5DpHWz4+yakxhbzvaKYkBQ9H3/u68O
p/P+RI36eEMd8FG3/CnDVhDDsvfsuXY567fQeDVKgwyP3xyXe6wYR36kD40TcEN76OONRXbCSmtI
APaDlQgG+q4J0z5ENMgYJ/GQk3VmSHDycT3kSwz3bB6w0PWHFjGTifg4U61SIFlhdUl+/uBOiduR
l1CpYEaFz84GvVHrAl6PZjwbV5DHLjSVl8qf82d70nyBm3sGBuBxh+VitvltWaqYfwjpejOmdYOr
UtETDQGaiQTXyUDa/I5Wd0vT/wkmE57ghZ5VY68PmxXJxRrKQRX9GbTfhnyM9bobAeeg3dFuYw0k
zvTsblJPMV8B07v4HhsjMWo3gpEAsJKreD661XXWvM9Em3uc7j9nTQDURIlrXQXoxiMZUbu9Cfky
zC+AqAmJqcFA7+rbGLkVcNK+0o0/CF6vUTp8YZ6tQRzrCnTwIY9Q9FOZ03Y2HxU1E/hNLfYE7E9U
t2V40mapDuHoggjP09m6qmKginOUGl4QPfEz53WNn5NVuMSPO0y5D6kBobQxxjGt8rWyMi+2dYDD
OUHxljzIEQ0ht3Cp/l+aATO4q+HUhmdpchJwZAvmkqRU/Rbj1EgBrdE5fZIkfRyS2RoA3NowAFdF
9MtMYFVXwdiTmY0QByKP8EfTfI3SDrqOK+CvIPDXBhKW6VQeqBah8l6lA2NEFJfBsq63NJccBrrs
4xXSDiwil2KozvYcsotc/2aw+9z13uvgmBn7yl05GjeuGiXmbHeaX8rD+1S/4MhUAL+RN8+GLLuX
sx9e5rLbjGhxviAxSWMVLOLm/eTpO3M4UMIg6AVrQHfRfyRHciHmawFpELCLSyCEr4cNK2tG8KvX
IMIC/tMBYb7HZP8kaQfpVj6hVCnDc5HrQX3eFcRzBr/oahwnLRyv0hmUZICaVzbNJAeoTN2Z/msH
wShtCMZxZof30zlHeTmbgx1ry29ZlGLVWXAD4ijWT1sq1q20ocSwtieN0d8P4CA/GGwZfbXE3C2J
WQ4Wcw7/Kem3DtERFtyhwg2YjsNjMlyvwf7AjF1qyESqBpaeRdx07wbt8s91fmAmDxiZzdCUAlML
++0OXubyEq55qA7JfAz1AvtvkKxH5j41h2PVxb2MBkFRO6N/AkKrlqJLtWglx+IJUWaeuayZochh
fOl3TzRXeAQUvhj/ipWT5nVW2bheDFlc9A39vVI6WKDPUVo1uVOb5N8mSxNwHfjpUEMLjnwlhbOq
oeJsvN5Gfq8kXt+/h5uApain+nvXMzsXLExnt2Q7sdhTVeTB4QPlgRk7nbXNDyp1upvr/5xFTH6R
BYlGLSkWxw8TbXfHOUJO9M1kcZvWVuQ8sw8LMm8X+12UxhIylNA5zpNeAzDJM+8RNsRpTKrDJeyD
Ty2QY76hH0XoRNuui0VLRAWfl/jK7H00n7LjLfgTPqKY1xcQ9z2ytixrQdY7UQbF7+RetXLVm195
RoFclIWjJC0e7QxNBoPDSZjvohqtIeh5FbU7vF+0uM2TKa+hnnqf7gicbf6vO32yE5h7/M77plcG
vEGF/AkHyv+I3vnZgIt7qkDTPhYuKsGtCT+HjsjimNfOAhVMX6u31LEVoGAbNiItMkBm6z+cN4iO
b8gnsH2Qb7MFwgjYopWBIKGEvFTJmy0S2aZzecg9pg9/n83kzM3ZQr24X/R85l66t4cREtlsjaCj
Bzk+t3kz1NDtXIX8Ry9T9L5+Nl9PIBUh8ZqwgBs/FDlSQxmRExE3UG+ZPCemlmfrbgPr32vhjK9H
3c5kieHsbOYlCQS+qlCcFthP3WC1PL+TOInF0Qn2iOI2RxDiydp/jMVYojk+vWszv4UrkhXrftdv
OFXRc72TXdtMvlnodDMIx6T7KpxBP8cU+3aCtgsw0FgL3RqiAh0ntVDfz7OexjZVBMrVQkAyc2/n
JQhfUo9WxtSnVrrPlQI1hS9WeCckc0OeIl1qVKQPbZa9xYtvC9LD3QadbPAeHgjCEPmioWUfwF8q
Ufl54c2axnd+Pkb/rc0tGq5c1F8R07N8TiE0ZE0fYw68eFNb1YgTTRKTu5rlnFdHU+3Q/8q8/iCx
0n8Wp3di1z/6T6kBZsOO92SdmbJieZk/k0/sFUEgZd89d/h8zKsQ/geCjRr/AaOKhnXAWO3oXxO7
n0rbVBWPLZp5Qzc5ayojAtYvpSacWnNRlRcWCKNeZmBwilrZoKSj2CLgX8qLAT1kVmfk0GWAVOe4
AJyVGWfKXZnifBtfbq6miUZ8Qo0sQDT3EpmN46RHmaSju4YuAAGAJyYGDwwIMnxmj4nr7LKhmAjM
WIHyf/gD6TfR6SKRnybCNfHKKRsFJym/nz1/+mpVsnxS7oN6fWEGZxFJ//GPPvihjfIff2DALTC0
jnIsD4SaAXZCZKGdZIb277+/EdDL0LCvuG8nzKg3ctSSpJRZR1c6JXOvWUPDXMJsp2S/T/oY/7sD
o0GufQsdDT9xz3W9dAkGacld70+ksbMmBx70Azqs/tS2mm3au2dZSJ740NpvQjABQGp292mU2iZB
v+Qynagr05Ia9JPqXJWjc3EAKIKlSd+8XBrQVRRWb40AVXsUK7I2vMbpp5ir8wgeUx02eb1E1UHh
iOAQPlUD8gKXBKJYtzZ8tWxM535ftbb8JqaGlmkfOGldYfuF6/wwCp16LnPs7uilrKw3kDf6MVue
YAgP4kE6/RYm7pJIJv8xqcY4stjPdtz95MYvjdX29KFABzcxPLx6YCK/zHM3HR4K2a/URYFYG7nQ
149fldGZkU3343omMJ0D5l8eekC66hlBsQTkk1r1dKc16cOlOD4EV8TnK50oBx7hFM1pNOnHiY7S
lQXeH2Lf8ffbahyTzxxXRLtY+fnWo6Y5QkmM/LklXj+nKFmG7gqnyByWXVFuuIjsyBRt8QDEILvY
ch74er8NSwDAXIhDHCOj4558RdRItwL6DZkAEyksfS5EgVrqRpQuUlB+KMLdAxmnj6CoC7Vwx6fe
BUdW9NAG3WquQLONlRVt4GGf5L6caokh8+DQIdnncFuh3f3otpZsKApubeP91H7CYm+0FGxZYpGg
WnutIZDwXFR64ICoSZeoH2q9A3xXxaBP6vi7zFdoFCQjSHIc+qY/GKM9U+IbsGgvR4bk0XTBnta+
so7sVNqUZppB/9w/LOzU3gddWQjmq+dgCWf5NiIDt+olSWpDfGop+6EHbeZnxeiywrp+Kj21UmJk
oeEpvUrHJLGDkJEJEhdo0c+tfn6YbJeKa4brhK5zJ+XtpultyDMIRDeI38GV1kg3IikRhmi+bmXO
Jg3FbjsOy7ZS33MhiQX032QR2ZdiACCiTsH+Z679byL7h47NBUBemhpdZIlEfK0ZQwlfvFUKhewu
C6zo40PPQqtengLJNbkQcDacLl0VIYg89JH0W2I7a/BOMyswUCemu3vLZ+YeNbHWsFKrZ33HnrN6
fDj35Rzf3HYiaSRFWstV718ivSJPe4a8I3XeG4CETkCjNBuKuaL6VSdS0CHLeHFFsSFDB40YbSNP
r28OX4MLJSGHdQhXbe/1As1kCR7VaqwCciA3gS0+tNoSNtMHToQP3F3c+IrMJs+KdKtg1I3G/JeN
o9EvlVuS6NFpLkiFQ7KOwTCjl9vdvkj1caMdwrTFVaPSs+QMRnoK94SdWqeUxGRvSm9Lf+ktGrbY
dydl6Lr2sUxx5KKDDPYJF3zVCtTpSS1d+kHWcjsMtRn3CthbfNl0NDyUFM6YFqUKLU5WrYGBk5Hj
XUY6KE2BAUfwGbjeShU76heEef3yAj6pa0bNGp01WI7imvgjgwcuocYmpA7qdBfWnG//eoZhQhUz
Tl3HlO6mKZvWXjNaFz/KPCkilim+A2hEIBPzmShDP3dipz1G5PWJe+Ej1/gJq2OgvluLxNAUJYxv
+6purh18gy0M3JEtNpS3RF5oGQFWvIbnxbvSfbw69Ba+4goHQmNia8gVdZO9GsMZXa02cbib2Mhu
qdYJ0UQWJ+VA7Fgp8Yinkn/yTJCwZqwxzlACMF01odp2+FlOyuVhLg7Ft3sMuPcyW9YBiY5/V6mX
3EcdGDy3YWbP5tWGnNrxMGpnJ1zcr6h0CWx5egF2T8BMrXnPgietabAsEHXDfp32EpJ677nmJxKQ
/9v+F8kU1PEsEANSCzVLv3Ggg+JkCZhuRXAyG/vKTn/NK0/TrasHjIZ2ZjMqm3Ckeg7XOaOXSqeB
/bMnCoZxaU4r9La3Fdw+5mTJs1XKi/rzqPME/1BD5l2KdZitAWDt20puRDea4VtynCyJOixfK6Jd
kbsJs1ASxirXpE3PeH8GYjZXAGrzBNKbq4TwMzrY7V7/1WnIy/O75ie829H5tjthW5mHG5kktqnU
7s2ZN9wkXOX82+eESdo/h8OSsuyy+ghHrOAty8OVLQ/cBaGFy0wY5RCszz5wAYEhBwdMRxNS6iTw
xpQyFCndJKRDmSyCeHzIGAPHaccMX2ev8nTRJA6GzHSsdgS4cEt/jbTGtjriZ4wsO8U+L22hHya4
oy82VFkSftLwHnRp/zHdDMJCFc+BcsAnB1+VWQCLb9eZ7BPcyGTwkZ3OAB6Tb7+DuQLhphRudAij
x9xe249TU6EWcIKqeh9rNXC+1PPEa5iFBFrVH4vn+/+iJMLjJFFxljSOeUMrpkixqqCol68urLVA
4o3da0/vki1ZYaDLQ4Bw/2DRWGI5pgEojKiKwqcvSWL+z6sfp+hGnRPFoiOlfLFUuD+BGRYXg5Jn
oz16lhRvzXeA3IeOfYR2hPJMTH7aKkg6J51NtqscMlveqp/mEvY4Lfn6O85ivXzAl4NM0cMK3BkW
4u5eJRVp/2JhwS4BIENZh9HkY9g6vFqXnJoFwYryN5mHEDkKh9fNt+K+nUbOhRHYkUTtxIWo73lc
DT7wfvjriiKSclhilary9IW/V/wJppXR1rgdtiVPJeIWZ+6eDvqIBLtsMVkWxf3zDUzb28kF5/Db
rM5wrv9YSE6ce/zHGgyaAhTiZJMNVPX8wyTipy4hhF4ZN6Vcr9BzUxeo8hPnq2S9O6ufanytaNXU
3R1Uo7Ucbw6vXo/CkYi3Pdk8h1wWHa6ABour0X78weK822AfqFddIS9Y9TdWC/MVnO6GpVR0Q2Xx
iTITStynjUxkT5bqN99MNL+LoXjDBGTNVvxYRJR9FbGDyMH/NN6RddiOTfxAVl0i2Z4xOtWGxxHu
p2Y313hWmTj64YZcF+MhR5i6aX9slUiPMBhyjXLuCx5pBtrOjsFm2on1Wit5bBia3zwZl9PIV0xG
sD/ZQd5h3MkWefbzYz8d039Ljw/Ac9VvV/uksFCz4o4/FaN1nQcBuEzkbTCCKVErOt8cWcNePTS5
RYM/+Cz3WBenhz+a/MJzDumIwntMkGYY0tCdnitBRXl7YATPqmv36r2ExXoFREKqMVJFfVPyox02
cdk5wuIH2CBjqcU+VmvPfHi60rGNuAkUAHZHxTr1xZp9my7dAeh9CRvl+48zY/SVN6B8mzyRAj2Z
W3fzEDmFZ2PqUZjkRE9DKlkzMvJI0qqpCMoUKoamNeqvA757CL4clVcc57Jsit2xIdywwPUcQN1M
qmmPHama/Van8rvnThv7t0al+BvR3a6vUfvZzk+HZLV3tr1lqJBxdSLit2NwrdiiaJ/6sfBWMRhz
zWuIv5o55YHgGDMyNWwKDm7HSrU/hblzeXhQ7cA4KA/awz0aqlJ3VGFFWdKi/CxbYiZLj+9K4aVc
4YDvqlSxndEYP+IJGcSr1UyM/PV50CYoj0tp2/l5/nNWrH9L19LBOOeT9D7QN5T1aBYGN3vtg5Fa
CSmwzOfuDPhkmFCEeS/Ax2xDjQt/zeV0AW5JanYAKwL17CRY+JziYjOFN3ra/+oa9PzR0w+SPasF
mk8Br8MP8t5taIeBkwXht+rR0O8fRDSn3SibNfyo7Yw0tF0QzmGboVgEodLcn5EPI801D1kFygVE
fX+EaDzmgEKq3OxnM3c++6X3tyQoEiSsbg4u6bZkceloXsF5GD+DtDlL3xszxJj29dRAN3LgBjIR
w5tDCX19cZiVUbfFSBo5x30gjB5Z/qgOrc1SCcSZg0eiAbXB0LHpKCxmqeQmJNOae9WrgVVhwKqH
t3hJviTTOtdqmgkcxpRSt38EhDiUmMajF5Jrt+qc/fVG3XnxrmvaCSItwrqdmXi5PaIqRdb+jl1l
SbImJqQw3cVsNNt0mmFlCjVK4t6jkZEu07NotIRES3MYaHbWzduKeKabcr5uGF/BF0GMCub5T9vu
YX3uQR1wNRWYMRrLlZcwL0qyNcLsxpuu7VvT/obstUGEzKY675gYFvlZImTNRsQABie4uBjHzhWI
hrWlzcJelXpLOkNYScDhDzAg4sSpXjDSLE5Zw6wxEkVhV60knaJh8LymCGrkGLB+jeFh/3RFKSRr
iPJx0iswt4zkQNUgFz+rHcsW5VHVv1irOMwgn6S40Xlk3gJVtpGKOia6NWycrvWabtc6BcSwqj65
2SB45Wtw/Okxjvwnlr4b9BsEesDtQRFzV4dK+EPATX7huY13R2WTd4caPFJ0V1aQ1CymtEtyyXL8
nU2gRE2DR39mEJ+hNuI2XLD1JlvBGbTkERddLp0sFJLhp7bvuZyI7g1ZnsgcZ5lBjBAFCUOtAdwn
AG4r3l0Kb5Bz7LqE6+vyNQPwTZ6mQuN8bZBPNZQncDz/T2ORc6BRkoFIcTyiPIbgmY5FMAmPHuRb
bvwjFd2I6AOvF/Ei6CwLj1gI6hEfyesICbgTOsoHY6iexbqFhyqxZi+7VfHbD5kjAXNxsAa8jpMR
xyALwxVNirkXbiX6Skl2W5MQtN45SLC30Rb5g15OJ3ijtH1OWMpbQ7/IlOE/YK48SpX7zjP1bFgE
yIBiDsFN6iJNzlcf/JpVJugW/0diXIxPGYgU7hsCKNSsL/9HzXGGePK/Jz2qlqI9hje/+e3OEnMV
14om+CfcGU34OL0wYqFA8N5bBOwZYHymV1w1hBsjpKbtyod+bD9SD5xYQ2TFwYjmltaoxmJDrfs2
n/Mptj8CDnWrONvM8Sn3RBm3Lwo1LR+SFysmkMn8xqpc5+bUHiZFcAehzEv1uhapWrITlCmEdSYd
mvHpxOqcx1J59+9vrveDQ/qgwBvwxclw1wrP4R5bFntNnENpHdAxaSY5zNTsdkmkBSTir901r0V4
efn6Zc94Wpgb68/e5So+NY9IheybeG+MdoV1KUjMW306ymGeEcMjG1SVivEnOWikiRexxXBYixFh
mF6lpGpbj4nCRlCcjFQj2xQuFJFKudVSKfFt3PIQbBrNc94JPLhXQbvuc6wkvKiasPXOp4xB1BbL
mV8wxAxO0SP4LNZtIxNom7b6VMBAzrmGU9nhh/EaUEvoO8eoOscb63qVJ6fXzUVf8U+9tXx0ztto
tjGMdUQy4jfNw8DR4pC0qb76SJnlYRS3VX4NtuYaFwZPlcEl9to+DhABf/jDjnNYILb4pZc4y9s6
CgNU99UpYzp5jW5IPWBXIIfancXFyTnqGno0FmoHvpQHDVFwhhfxpa7juqY+cPupRKeaVMxVAkjp
+qVo4AA+uN6in1JjvytMb+x+p3juANWSUWUtxSY7YcTuEVHzsK3mzYLHGmlAi5jWhuFfMq9nxglr
D0j3QzjMadzYigNqxRh/0CyZsXs3T6Fsey7KBzdabnyXI9KtfUeYGnZL/Ci8ABi7dsAC8gbB0uyy
EexpfnoSpDy86TLfMvj1qqvT4srAhtsZHMPAoZgUwz5AuMA5MZ7vhp88sukXzgdwKsVX5VRPyGn5
oR8UDLf8a+J5V5AOIGZl/gtTlO1tn04qx4pQeF31U4ZL8Og36xm5KxkLwSeR+fWxQ/GhDnc1DDPl
/pCP5OJMmKg5DUtxH7zNk4M1BBVXSf6WXwFibfT8rUYrBl0X0j2KFbeF3d+0l1fTw44E3eTnYsS2
3xJ3eJlulIYg9kV/3u9nlwgOMq1aZTmMm1HDMJfceppaEraG3LZLz5pwEhYWiWDLfy4lKC79tsBI
AV7CQ/5XregBdEmk1S7E6wngVv54AUUwpe8mmF6SIMLevRPMzaabtkTKTYI/VqM9UlgDbUlhaypq
JT7+cKEp3JNAtFvr5p+XFMZCVmIBLTKHFNQ8ZTfD/sm+sZxewxGQx59wbbRW3fFDkUvjXKiiAHFf
82+rZZlMePNBbJAW7lbKv5O8Bk0TiIQvrsEVeP2VdWRMx1CsPDHTTEUDcZ3Y3+BNEg5J5hT/KbQT
hS47AR3CDNNqSnr4Avb6eag59Rz10uhsRyAd82i3coqMHG+XFJhdQUb6Pnn2XYjgj2I4YJCF0Vhb
F6nZC2Glp8utZGvz9jE+4sIj7izBCmCm8c1xAmmvEB9uwtASCtzrTRTtykymt/Sr3QlbWrT0kkbr
ycL5cM37GuSCNZZtFBB2lfQYjjXtI4xc5t+HTtAhKVJMQwAgNEdNNlMFjODCxxyZYW0tW6UbTH/q
I/l9Z3hBmqWqbojmhb+FxHCs1+Q2rb9laY7c2urjadF+yw0gx001JwAVm6fBerjk6ZnsWlgLEE0R
VgCUjt51qLwFtrTJjJpLQQj0/ZP6yBFq945eEoVLQpbqftSUbk696/6nOJK3OKj7kZ/7ie3BIFsa
gqaNIjVKcujEzG5S0O1UGmFwlJ9+XzirAPs2SAHQRJ0lOM3xTK1FPuEnbap4Elv+aFdIFQa9KL0q
ITZrY1a10me0CAJZdXZ9NRRpz7fnEOHdL0x+8SgrK1j1dPxvHpxu03EjsQQMogPo77HhP0VF+gyj
jk7wzHPRshCFFJn8DQFW+/k4Gx3U7tsohpEHErqYdanMbwrEXguEHq+1kJvftHImzd/GWttm0MML
jEgqu0oSBwMcjBP7BFPyDMFNdr4pHGVrWEngnF8k4SkNdkECeJLnnPLHtBFCz45SYjuQ/gxTY7hF
0GZWzrgYBI3DsHSpINHQrc2jE5CSz4xJaIvajtoeWGcZheYe0xpz1hF59WpEIPe09haZYSsLV4N9
c8qZ/r1UodBGKvDLLAPMl50kxQcWJvd4raBnDt2+i1uLOmRQcPSo4Sd2LKXCDgseyBEuIWnmgpKq
nU3cmPQGc/Oq4Fc599BsVXkjQtnz5Y0EBvn4T0PX5qiiDtMAprg2AGo+AEuTV0YPw5l/hUAivDB6
GpToO+ICiF2S9ncqMVX4gs0vmeIYpYD6Ed1RUgwA3JBF8xclAq/HCMt4ptU6stT1Hwa7+thBMO3W
P/g87neWzWwz5KikCBBY8HJOqpZhzhXNDL+N9AybOMpkOYf+qHFPjIpzAbRi85YKKhG3l4v0GqNa
+rJLMafPwwnbCrsNKAje1MHRJ9+NI9HyqY0jzuZYs3UBaVZYhIkAnz8L+rWAae+SlTAshD2C1T7S
PifzBdrUwucy/IaEXyC9DLlAXlLcLLFjtX2W/Q4tYC4fbDelxaJEGvxHWZS1u8NIosev0SzWniYo
+FXtblWa7RsGKz2pjjkLUmLCacZHggBMdLneWcsWqb5skyDqIBqKar56R55r/saEcZdtzhF5nopM
sRQvSKDDpUePZthjNh1pypx8s2TCLLeY9mHtqiPqyNJFJKuCwNkUM4gi13baaGGkyC1rcCJjsu1h
JP3BXTATLd37fb+Rb5ETaLNKHiiTG2PfHiohkX6zGdmlPZnM0nlZEKUpoiuC+Sj6LLfaO+KHLuk1
fkFoAKw3BKKU3GOpQptYT91YjMGU1WmAp7BsElV+d83AY1Lwnvbgp/W2j+OS11h7sXqFSmocRZJN
VuLAwXCnL51fddF0rNLabF5V5x2QtSSojjBhg/eFkE+bOuz2Ado185J8DYhTIeGrRZo+ysR8lGqs
W2xL/E2wN+Jv3dow2WfrHrJSEmvuzH3lXCUHv4X54e5eOFsd6mcj5rKp6H1oBbLs5J5JNXyiyClu
2B2dU9eOdFJeASk4U2nuux+VjSiD39x/qEBaoSw83Ng0JcapH5x5P0iugcsgxo4lfivuX+Rz34yh
krA524O+fiR3qcIBIKBCHAVsBElEEUxwUGwELs/PQo28orjUJq1vjId4bwJmXDn6TS6e8oaiCIQ5
UdWX7y73dSg4BpkRHkGez2et1PlNYG10kQr9dlNUpQOonxlMs0dgHo62HkZzjLmXHebyQdwPByei
u5VKT2VF9C7cDbpCvyxGjxtbqLrLoPmfCV13blqlCR4K23JKsUHfAKtY7gsID8PjyjaRVCLOXEoF
mNB+f/UNACLCZz5B4epj+csRFeE9dN+rzq7XIWpxT5dYsGX26teo5GpZCgmDUErJMqlvOT9wSIR4
Af7dL9PaVwCNAm22VuzTC4Cx0sE72CYE9LZc7XYMVUzDJQRO0rxiY+XFTA/hUcqeBEkEB4cy/bZ6
+DVfJDbjKhwG9UGaQeW4K5MQryEMCFneDEc/LX8YkSCvTrI4Iqdw8gLVCO/DtVEQlrSNif+f8vGE
lZkz0bhMJjf94uTMPDxOJortaTADQ2Z0xbOjLhq82Q2Rc9pT4sWwG3xKbhepX1/FVWnYUUMluvI8
Ya89N0OEPVEAiOuJJNHR2LHfZSOQupc+DsA9FojRZfus3cZ/4yWRsiUkfc5EthM74H3bpPpImo7E
aDQCeYUXtou+dWNduDEji1OKntv+mHxe2yu27hFyPa2Rth291YmkF9Y22/h4egq4gipX4iVPTiEA
rpdyUdGs7A4J5qjWo9r4NSvdxrUVLKjCRF7Z4793glceImmOnUhYDhWXjhwP5YTJVjq2FKtQ3iSA
TL746yf9a6k8T8B6q9RFP+uH6CnJ/0QREbnkd7/mv9Y5XwQehkqPMdQ3nOSMcDXBzc06wgAO5P1X
h9/eBqSMg+rO0lLwCwCArVmt7bEEUJLzMrnY/E4tHa/6ex43bceUYmM83ew8KcfAdj71G7P7mFFI
B1H6NsphmaRMf0PUuKd/bnRxXpeU4wBVTXnZagvBOhiOPFswcxQvOhzPZvA3WXyOTcYB+rAW72Zk
wicySKQi/1fl5ou/Ijp8AQaBeslZ6yVVvlTFhkcwoBxuyWmo+BFcD+GX2OeMxhhdS4hJNMINSBeV
KwCm07Rq0LuVovRm2HKyGh1G5yr3oegi8OV4NBZdY71TgDcbneUbdiNiiNhGB+vv3stUL6kZKLAy
7elzTKL5M7+CTco8Dwq7lRgIrOv6tj2j93u6YsZd77tRqQWmSBcVrr2ElalhIiN53FT1IP/7y5FA
nZ+Yme99wj6MG073CzMUrM2tKlJapOXBQtor4V//jIV2E/e8Ta6Vp2FfC7Zl7brOo4+cfOhg343F
c8AeIPjwqRDKD/VxYPWBLxww3MxP4UEESLC7KjsUu+6Y7a6nTqcHqHY/MJqRemwAP20kvKKZ+CFR
Jh/YKEp2u948dYzCbLa1/Acb1SW8dmlcDRUk3Cy1X6dCYrZc0y+m6dLkkgpywUxJrAhisRPp1002
wOTFvMvlW5+7fwCF9KV2Hh4JsPuvahE/WAK2xMkqZ6a55gY/1A9qtOgBpIwilXStBUgOZNXE2Hm+
GJw+oMFTxI2ygMwlJ5S0QRdGBECEYTa0AQRFflCbQnbdsf7bMHEcZI1dZ3GksGpKvSBo1KCresin
XMDYHIRwEFNjABNZ3adJScu2PO6S2gNu+DaWHs/+fpMmo5HHgeRRrMFIWg8RxJLTZmMG2qT3sJTq
/2PacyOrWZrVye686/rj/R4WXYkxXd7S4mKbHjahFjHNGnQVEiFIXl7FTZsJSnuTwkWuqgyFB0lp
m6ttvv25m+xBQCwXkob7ibMkiFexp/kNI+mhQMa8ag4x+bhSLkyf3OJDOujc1kbQBfSwOz6aCXFg
BmBe2q4uJfUgiAyB1PeLYBaJoJ4OpQt+1zmNHsOcHLds1hBNU5Ib3Mbk9VKfTDNY5OeK6PxNO+pw
DX2j0OaHnf/PU6HT42SURHakMfIa7ABQ3ykEY5JJC3kdZeJL63m92YT4GrdazbbNpUJYiFZOUKsw
ZNmUrknKpTFMDkAQkKCvt0WblIJd2FLVCZU8Nz6XmUkPcifXy6dFzihDMkhoziyXvPgsyy8a14Ee
DGIdmO3/Gy/gacU3eVTyBqRhEx4xcygzAnqPpRdNLqJMKzWXT5fIR1bi9wY415YUTg0dqXwUxpkZ
7/QCJ9UOM5Ybtak41vj+9pYLYa42rI6sfPTD4EdX3PsKfcanndTANvEa21OU9evGsmQKn53ixgTL
8ZNCLdju7U5Tad400xun7ZhBc0LyZJvebfBQC6U61bHKSQfrUydBc1R5uvWBhmJLsNKp0fx6mWW0
D6pzr48ug1mgEqEkifzQ+CZIdl6E3IB+Ab9vrK76iOROFdjOVCw0nI/30DEqcocvpYvnemwkxn3/
uaksokqim+aHxfv114G57n3eFiNaVE8K4RBVjUPEvpaKYnWSL8ens1nV1kl2Ilvs+hznV+w3OK+K
7J+sog3hb3mh7vdtxSZiNYc/giBzf5QfW9yYq0zsWMwz1k1T2/PP0xl0HOBUu5XGfD78nDMhqbeu
Kz8eKYsB9UY7ZFCRVe5xC0vU6jw1CEBJn8ylKDT1imKxMjcXrxtrDLLX77+QQqp0Qw0Uh09m7igE
ZmNFQHzXXH7s/oqg3EsSpAX2wVO4FMV7V+F/IAHW0AIinoFpE3OYIYPj5iDsJqqrb2BEJsmnGWj6
0r5b5RUgfyjVapLdPtoMVCJkUjDY9gR8/UAUi0H4BYSKozNwYqvc8GnKtrZJolun+Ux7ZOEFw7tN
X5pNT/V7EIavh/8jfbasNMHOOpXLzNpBI4ioBYyg+CE/SM0a6OUori6PIa5wHk6UnCQX6Gxf9jPB
zRAD9uo6xyqaUiijkzE6QfAIhdaTPPBFB/1XdDDVdHC+Y9LuQT0fu4pbRXrg7xG1RWe/M5fC5poZ
dL9ljIRgtd9nW/1Zsd/dnnayO/6HfFXnAbN98iX2DdE0azfq0BvUb07B2fjMgV++reyAvRGd2NLz
Cqcyf36zEVKcLKJ9uo/E4ucyWlVfmWm+lD5Z+GO5E2pXnw4T63j0DdhkC23Q/rkM9D2Hhxp5sN8s
NEcUUllmPo42YX5wD0IxCvD/hnnbxWX2hZovppH+hhHTRadbsnqoqaXmumCBKgw86e+4G4WwnT0e
wGnVPvxtsDJ3LC+ChDjBegmbfzI5Q1Vz2Hdn4nD1Thc2M/6UeXqdp1p2DYTivmcTw20kJMWZMHum
v/6KhuWPatfSwz6IJ0qjtGM/dzHcJUNtHnbbCJixd0Pp+iVyHNsr5C5PE3R4FxPAXQpFzI91u87S
uQz7asNsL868mq8zv8JVWpet2M9V+NaLGcjoXqGWdrHJ0684R0YY4KudXNJoFPieTYTPfXEnEV2g
QcVAI8nG9dnVd1qsgqRlwHNP44TNjxSE0duXoIrPY1XVuC0swWJbsG2w1QWxJit2NmLFN9zF8iQG
Woit10RmEmUCc+c3pEe34S2mbeiqSp4WlplvHuVjebWT2SDO8UR+ytDHfhGQV7kFkhwGIymGbUMu
gLuos16/kjnalnkWtIRYDe6AUBV/JSnaFxjo/44lynwwvOP0GCPnrMz/cFztuRb6zHN6h6PgdBqM
I24Kr/vGzXD1pMUX0J8QuVRwrnMAdS9m3QyPyIi7kZRpczM4+p87Y2T0I6saznKjS/1N8kzi8h7r
kdWqpRXawnqat59htmZ9TUc1NOTyVdzwp+o6wUfYOtcTA0/kWgKpcXgkdbK0f5y8rDA5PXTcwDJW
UxWcf4+I/cJhuz7DmxC8D/zjiXlJGgekX39WMpqJ7nNivlBQVgCGdi0EXgqsqio8+Q2jhkJiswob
9SZjPG8/o2f+I1nbyKeye8eDb+aOeVN0u46fRcg/eZ9dB855eaXPRmQadNLG4sFB8Z5zx+Pw9EJ8
jMy0BhIb5VbDJ680IT4P5ayBGP3HdFikyYB5ttQxCo+QsCcTI+zduELxJQ8H5+SrC+hVXqqD1S5Z
BPBrH8BZTHxKV7R56LdmdPoYkY/PLkZBs1O3IvRXlj/DI6LNVwa97MT5oa1k+oE9jHOE1z3Q7p9e
unbaSmoQfMbnOGUu7ogGXU3eoLd0pthQKDFW7KnIMoVHFBX5lW0AT6tYHt4DfMJM+iEY0D1Mxvmd
WM3UfD/6g+w9Xn1b01YXYRlQN9F75nCLhqgTPKVCSR0MOYsNBu3MegYN5G1VbqSjNSzzD3RC5lNe
nlIUVw2qclCFxFgNqiLew2iUsbEYaXXvsXClr3y7v+DyapfNcqwu9mLwiCf+x4JemQ+QnUz51i/v
yx7AIJalYqXMkyFHeDxF1Lh1L4oyHZG8pxv+STwXLbu1SMKZAXxPaxWp9f7XknIOcYKgm8Jfc/kz
g715qOele1k4Dh7aF6gxVmO8WZXMlitVZZQqdtrK28MPqaVGGfNspT2Kpg97eF8q6XrO1O/yD7Fy
PtFRxrZILXp3hjY+3bUlY5SkdQ6RgkD4mwaD4UZFIHsQYOAnpLa1Uf0qcFSu/EgGqKIW4Ey1uvAq
iJy6/IhBgjY7Zn0ZAMr9YKA5TyeGZ2vI1R+hldCDFuGfrOj+2a2MeegZWT4YmR2gciFKrKqIJEo1
TnYiNe1kqk0zOC4R7KWKnRvHkbgVeQJyf8h9UeiHQ5OVbR6TJeN1OKv2OK2KdiCtfQWYH8GnMra5
id4loTPqS7gG6JrxdXdl6+inX5PENEM/s/ZI1zKZ8kg4ByOTmFmY+UOeFnl8uyY3bexO6j6qdITG
EtkcSTybBgPlIoHjLH84YxX8d4Z9QGIvKqlCknIi7whXBKKqbzRr7h+DyrxPqaTrrRjjiggmahDx
nhCJhv/qGYC//8FbgV+spnmFBhMcmDz3FZC5f3Udu8zI7/UbWdckkMwgKmumNauK9jLEwchKoTsB
yQbJ8+ykbU30yc6GnbJOeABPrLzyt7rqo/MO49iET07bEhS4mPUIOQRGpJnMCNQAUyhUlACfNNi5
TWoveN5Jj68N3ZftPzXYKIUEZ2tAd8pRUrDay5P+e13Y3dIT08RJ79gDcQdExGFgpKy38CiiQdc3
YtBrE5kjgJo8h2ZbG+Z0nPXXoXBXloNaJtQSKpCr2SDGkJiN5dpHM04oyOMgnsmc0ZI53Jn1e4I5
jh8SPtmQJbG7e1zabTNg9XFveoYUK5os/yHK1JiEF2iMq4JpdN05u5NkX3Byc5wB7sZzD7X/c5QO
sJDgAgQD/G48ngyVwxl3eMYlGt+QdcknYXHAtjr7iOBzdOFfKz/qdK+QN+xloHIQ7Isiu1OYoNjt
VxoOQ8BMyM2aL0ajY1fA5cgwlX70Y+9ZzGYliA+XfyuODFnh2nEG1XTEpqZQ3F2x547ZoGkzjD9H
75qomZcLdWaIRN1vSegURYAzHEluaGkopU0ORGNkbOarJo6JIKbuNc8FzNEivax7b8i+kDzWnFih
0Db4vNIKmkQRPqcEVw213S3ea3rD/jaa1IoJ8Lueveq9ktZZ3HuevFe1LYHj8zAZm5REwGr2AMlB
Y9ojsIsGHfTgeD67L6HTyomlpy3LZ56bJnqDyhy6KIAFrkj5VttxPqOiGFadcJxskU07a3n3q8NC
7d3pZvafhSGGcvG5mpgREsmQKquvI5DZsjXGkUQzDoE2YX6I3r72P5GNTn3vxw+bdy3p8aPiSEZw
bHlyt++cJkl00H+YgLbzFHExeKuLSg9rvJ7dvDxMEiKHYknIy72EPl7Uwb2zEw9vgKKzF8Ua2/MT
Cv3rMPu1V+c2Rl5P0cf8skYeeQHiAKGMdrYa1XzrB0l1yZz5V5mOqFmwQFVtjgQE5f8R4bLkSHqh
YtsKNFkyqa4AnSi8LqUbQfC3eBfCXBa0ZpI+2jLvH81mFhVvbSFtYjGEPrmAXdgmM7PGqFd8l3x8
ChNQ8RCiILNIi+YWA4WvwvjKi6tYrkbtALFJMiYEGjaQhEKLOn2kkUNhGfgfcZ9dv1EaPTHDVqDj
rOs4zDcDsWzKkdtyQSNRSCwyFSIlyP9e/UJoPcBoHxCbEu45+quf7c1MngNfkk3NRfzTo1cmCb2K
XjEfZrd2xpbD/gPSr5IINdBV3iFrBG43/oRR9oabShQ38jxKYxiAWnkIs2gl5ur3k+gGdP2hSJfH
nBCuWjkx719x40pIbt5vFdB/Qr9DPdbkN90VjIfULRMwCSj5HQsSXZ6w4kqszPrBqaqzMcAFSgoH
Kb3KkXpoLZPxhTOgte2eOiR+tLzpPp6xRy0LqPvEG7LFry+6h02MsP44WJWSY9Dn+CutbDUt75DW
YUh0pIrwNhJdW8fUnpdqqtzdPmJG8CYAkwbZgk9L5lLb39ybkLS5AhxPndfaawS+PGqSkNk/oE3y
ZLMxBjnAzS1hD4ppgge1QO0SpIh0ULxyEvuW3tuMwms7MdpEgkeH1K4PddrHS25FsW81nBJkrqgP
lkHwqXFG0ijJ6idLwu1tIahCVhAPOygO2s+kAo/Erqq+GWPWSpJAg+6a8Achim6LsmpmCvrdEYmf
miA2txd5TgN3rn870Q0MMV55Je50KFvJI/egfQcce/2Mzn32jculQRNvPXkxOPvgVU0cUau6vh0E
199bK2GwIcznPyElgZIJ4vpuzhfNMEXNZjxw9sy/fri1tdMCjFRg8xRB1xItSU9njLyO05b6ClBI
J0jZ4QKLzd5jI78exgJmH42DN2hLKeMkDozxYrWLu9Sp8ifMlquZ5tXs0/FZS3xLxKZuISm+smaA
+++BArP2UHN8NpPD6Ov5LyJ9QaL2MqNd4TQzdFU9vviymi2SKpKMMForchd0Kme9TmE2DvTQA1YX
9Rv1HJLW/2OpZAxk/4gl7hIgaDzdIIEqeLCbooBSV0HrkUf1C4r0p1BOHyNlshftbhKBLDn4TFVN
vUjQ0jcI4rWlVVMW8X/U8sJaV5Jf10DBJzZDpavP8vUJlmurxyMR6zE8dU/u71fAXMQAgvnQlRH7
U66uwY3/YOLeZNLYc8cyEz8fGXrrTgbOBJbbTfnDLru4wcId+vOrt0tMO8KgoWr73icxFpO6BtP2
in+2YGmhuETGDcPqgyM8AdDNozpC724VZVa1M3A1K0uqCIpnk3XKQnU8Gk7ZWwtxZ0hj9kDa29Tv
N3W/EBThLsrw0pTq/zLJ1KkzUNy6qYlaTtCmXgdd+Iy2k1ks0vuDxrhXYxvawpMvmcM+IQ5/3hAO
2d/BgDzAiW0fjtyyN6xa8xLZqj1gCnl1dKOCNgpwbyf3TCvz2uAjJ8d0/HO7Qg9uluB3Aosj7Bsg
6QjXWRjl6SGUDRo4ghli4Hr66N8djib9e7X7Aguh0skARtDMeVrKWd43/MH8GsgEdZFTYowXZVdq
XbPOszl5wQKskTjuqz50ME2wjOFdH+/s8fOjtLNJWqupi4kUVw/lGnJK5odJhi2cvySHWFjKAE12
heQcuzvxGniatIHPQAZ0EG1urDwXv3JspzCGw7W+v2P4QQQTlcpObBSURDEjMoVQqdq86bze5CJz
U1mbaz88QYn769JW/9QD9GusYQr2M2K9EijPLpH56JRUEfJZRf5zsZWtnypnSlLLP7syA5oRj+wp
LcFq1YiwOP10TwuFwsuwsLrm0H8mjuGWH2h6qNNoo1/esbUAo2yU0rn5txbQzvVu0rw5BokpCeoS
W4x7Gy7Nf7L3DTLTNScGIhuVDjw0pwcSYf7uw4+EFZLDIYkwDOaJe48sXC0Xh7EEnPfrHe7iN1Ce
j3fUD6jHIRNimUwLY3MB7HIZHvVjhyBBvS8799A6Xesw5GiGHUuUVl5k6c3B9ia0h1GMCXHzFft4
afahCCyRzsIT1KGbtp92W2Vs8cM/DYCps1cnBv5kE5g1qDsUMydwNqtUEa3hG7DMrZasi1ZLkIw3
3EpEZz8jkrrAHIUWVv9PIZNf8izgn8epGWYuXGUHrUWwLEK2J1VDmpmEeu+mO0Clr4D1BxxCx/fI
sLiTXucQGLd6/lMWoR3jSVnawAuN6wZxBYzRqTOobNdoK+TodXsN8aTylrBSxhvFYO17HdfC86fN
toN2U8Oxafp59JKZJVJDH4+RVZSRplHFYBaFV9AEXIuKPZadvWX1YhMqGZwiIAoiCrgGM97JOKLy
Mi9+L6SkI5p8D8lnBNdRaDU7y9IkOppbg5G6ZVF1q79wWLugZPbsnYUeqwNsIgY/WMA1sm1MUW57
0okM6orkc7ga1ONHjR4RB7ieDQFatkEKChX6ObtCuLjOgb/3p7Y/kx56PbdZ+6px7ekc78vlIp6V
vRvkxT3wAlE0AwKEH06X/giAMfGNGMlmOOjPILGA2vFcld1HeUtcr1VGt1G4Xij5Z13KePzrESPk
FopFztnLDJs6E5u5WgSYObRm+H6rLGqZqTpd4MY7xGGW/fRRV8cOjdPY1Yrq9NpwfrX5sau/rD1X
q+F0Lw3nU64QJD0x5VOvlUzRcmWrh/6ZGo++BZisTEWyqZcD60AR2yeb4wvXataUIkLPJGmNuzTj
NdXOL47POvKSso/lu0fmmAX5CEHoayh7T65/dxc8Ac406ZGbb1v7egtv7rOyHyUT0V3UGaHr7RYd
qNipOMNH+DDp0lNUCZAjn2OgfI4nCvkly6+xWEOAAKfTwTNGiv1SgswSH1dxCg5psq+MREckpYNi
sN7boV5tbfwSB1P1nYk5NumI32C57RWIekjdVIWK1EEXvxjY8Qe2IPfTuzy+Uj9QmSe7pGx4aOmB
C587RsiGH9mBhKsXdc2oZT7jZEk+4XCj8l38ON3SCJNDQPpiVfsay6bT3H/XnwtuVegSoSi6RG4B
XHk7UkrcVv5AJC9kiamX95YSuDmj4qEAVPGmFFKVhwjQE8SrIIxirxKsM74IcTRlDiboPF8OfU86
Ut66Qh+NxdgqtBa8zuYIH2rcOxACZyheAAvxXMDeTLHKlHwSj4EYHsDfUi1VjajMhERfFg1aFrBG
ydDYwY/X8tx8jF4L0QyG0JuleoVAqQpOlryX+NuWas4kCNmSjUMzFfX9wUjkwS9lBuUmlLpIXtf2
xtOuDBy9pi2cXP2Nd8JF04s5g7887j1dZJY9IBgNelJVnN6x1gl8HIHUBwhgNM5aSmVpSH7TzYT/
oWsPr4rdTILNFJ38hV9ggUFSztAdXiNuYnuoDpUjMdCm2blpq7q3l4royCMDe1jcoZtznbN3kEVN
9eQ7nzfPrZ8y7EyYKDxk0x4mfVQl4+YZ3AmFUhIgTBdvsvG78DaLM1f1iozatRIMFrBeS6N1Q/bn
q+PBQQEP4oN9V1RouMSWU1d6uvl1S2NDs3YkpkNKBxqdYJTRV6ZVqDotoDWyDBZ3lIJlJegCOEwk
cUVZpbdfEew2NiQrg4X74b+jTgqw7Y62dOhwez/PeAqnBUl6WPSrN+CAKkKYXu1ps8+TJohxssCu
Gr2H9ZQIhPvBci3EqgyuCX4fV/nFXixMblyqcTCG+V6l4T+JBGhwSTAl3tABjwZookQ8v7ruxEIO
dFfxBDlgSRShAFpHQDeXY4kQH8xbO8e6E5bobPOBWR708SJfJppOeM6JOc97oHnwBEP88PdgQPgn
xuVbfrW3Dwl2rHXWH5/9rp2fPg1guTpnkuBYBdgu9AZ2Vey0LWaZ7N2/Haum3b0l6L84ZvIWilRA
a+mlRN/f0RHzLeEBk1D68eTJ2CzddfG1c6h6Dei2RT6SZrftyFZwF1IOPTXnflPDQh8pKs0ANl+6
MCLvsRdurWx34cbpB0IwPUG29XbxaBpEugP15lXo2xFQltgAJmWVOYBhsPfIKCHZn4nP81hQS4nx
ym87kALOtx72102/WhGV6bQ4sZY+fFn0sr723HCxEQZ8gwco/PIlmvb/HjDEMU0CwSBak+HveuCJ
oNagCkt49W/X/q/evGc/142nKAKGshFqK/gsZAUgb/NzoEKzFUW4D51EKHWe9UP1hrEgbAqd4Hty
5/QVkpHMC9ju1TDnNBMLNl4gC/FnpfZeyyCF3ZWlF7sNJ4tTVGWeG/VyexrZgiZf0VGPOgDH6gaV
/CGQPJ8t0ilJBcjrXS41lnLDBkEaF2jUVloOn5ULCzeMqSEuskNi6FII8PF7W9CKLML4/r8yZ/ym
vjqt3oO67BBVg36pR2xwMk0hRh0sEt9E+Pbqu/EPlU7KKynmVvEDc2U6B1WVtfxnjZOIYj7HbNJ9
LX5OspHNfnTeniQhqyepgUmfLXPZPBWE0rtuP/5rsjozZO4zv5k+GKOaP3wv9ggfSD8c+xShzCoc
IugW6LOFpcdrccimz6GLajcQopLn83q5UwGTDxtQhY0owEaVq/z1rofmPJEWtQnOxnhzEn4ARZQ4
1oXitFlFY0Xw1qDGWE3JTXUa34vUiJVdC228zs4P5CWs3OYfM/RDZ9m0JjCiOBW0fC+16K8ASuMr
KvGWL6Kgq4NopuKRaAsaVp9KQRYM84wPe8Dk5/XRKc7v31P3V5U8JYzCKHocmpk2XTJ625wkMuaU
wMna4x4N/H1SBkMnGYHxc24915rixn7vMueTfoAI/arifLst0gdzbNFGWc3zotND5YSf8iL9W0Y0
JrrqJs0rSqIcJikJ1ETaIkG4PdLR4+j++RhSZnh585EHASJBMUaqM24TvJMf3+UGPgO+l1mkM4ZZ
7QBx6donJImx+zqeSmifYgAfkuq89aSqekTAo+pJ2LtZO284mU/rv5uKbLput9h+Tfj9jQOHcqoF
IR2OTHT/zJ/zASZ4rh30yzQD7M0/j502e7uVKVggjDOo0Agz+PSMhIJGjb4mTxc8IO9U0fjgkIqB
HRGE0jgXKD2cKOaGoeJVLfEGXKqmzj2yDeCZNeA0UnQCjOEg5QBYst00/blovLvuiGsP9dcdJ2OF
Po6zqYLCmQfFXBqr7G5/TbfnVCMeOXYBHANVhR6Gw5WkGBukELe6Q4DGe7/K1EZygGXDHOkImHP0
D+Ezc60xpXBROJgBwzWi7L5bSNzNJRL9TQN9KgQeJPUNojTD2vGr3T4btvbxrX2x0eeO/HQmA6uF
H/6MRBGnAIaoRiKo7F3sGLDD7+l29dTmmxhFjBmU7KuqJirCFJPAbvWc1MoL7oazq+nEIQmr6AV/
bqLBA3DyxNXH9Y3+TN/hCaOiQaM4+Ryl/c/k/0IpBJ7Ya479u0mz4eNojp+Szc3Wg2jcPuPReOy9
Gf3uWg1Ipu6rXbtVGlXek9QyWQ7D9DWxl989ATb5CMlGDcBdwprbBy8aBHM7RncMXsSx3/jbWvyk
nni0r5jbuXWjy4pw7sU6rXtv9xM18lr8XYco2G5V5ie7S6eBjmWzKrzOcsGaeCUQ4LKGnR0Z4IVY
ugFoqDVSjOB3/wrII2XSpShIJaJmBpmEHoZkYC+Iw9ABAcCJBsFfzLHEc3YrJk/1o25ptFBWt0LN
WLEiFMQ2XQZCbW0j1LG3mplbhDHVFZm/TTk+JZa39GeYCXBn55h4j7zSHif+GQ1ETI6uDmVP3MPn
8A+W8mEEAV4Igc1DoT3AHtIW/a81djg9m5urONbiS2dq/S9kM2xEn4QB1QPmelgieVWfwjp1a6ON
4ErgCseIthKOYhsRgx234YhThzqMXG6PUaMNJC1H3+jHB9cb4NP+E2PUH3R7QSNNEeT96zuSTAJl
1rZnbrGgQQTW29lhclUuNv8JIBrCkiluZTIm2QVq7ew6JHzxkfgn36GmP8/cD3QZQ9ouSQlU/sMy
oY242VyDrOtEZNgjkcPDFkgeR1ND0rtRD/FCxI2dSF9z06fkgcHvUN20IYZeljTTxJesU48bH1gG
1sVtS9oWcxZN8mPFIDWaP8CXHxJECQO8RYDndX3wUaQaO8a8EHSs2TBpuWVv+ARUPHDM18h+wu3x
4uYpn9jILrb1+xR465teMxy3zZc+K92YoSxxpeKdQyCC1SfPRIlX6fjq0IA/RMu4e/z3Q4vy67mZ
uEPNSyKsPDxlI2oPTGRTEG7HUSRpX3dEEZTzv7psUscGiUhC7Wl6yjbfB4ZvD9YIernsN3gb1EwW
g5GPqSopY8ILnxNYWHwKr33Rr4Q1agUB2G636GJ5gP/FP3sJX1O0vyLHfIDY+Uwths6G4fgYNPT1
+8r3E4qJgD27Q0RO75SY7GCWXeQoR3qIjBQgRPxE4OKNf+XyYXmQJlHCa5jGzrCGWrCg0BIhQSEG
/Xggy6pU3GTkYYr3SQWz9qlQ5ueIoBASSl2DAh02DfoUShPFI0MEGZnxOXatk80IJyk+ldiuIymu
De4Aovmdw8fxTM7XTTGDLOov83TupAF1B3QYBCCz/rQswRCnZhwY96k8osClRRVyj49avS20FOoU
ideohikTnOzQFPxH1PTH6Ct8JSoZCKtGzWzJ+e7zdU7KvSKWsOh9wUbXuBGLIEftGUAnEqPsl7Ux
t1ayCZGquWPOII21jzObs8uLvF29SLBGMO5+yf6WVQX3aWE6cEuMv9o+XxbhksjFEYvKlUNNL4+C
0oaJnJ69mA2L1c/YjrpNo4BHn5L04dpUvzqHp7U7RPcGpRlnvFs6KKsbK+GauFkgRAjS/xXRzC7G
oHXWhISIkGeLXHMcET1BCDwDKIVXfroeDVQH4RH8PUgTsBm22WPmCSoz4pbOlgxsN/opn20PjT43
YOly2/442F3hSqwAyiipEKUJiS8x/O0EgiCrVMgmoVtKLQ8pxIlMXrJ5evCTKg5u0q0fYliaTcgo
NmUEjqki5kztqmpDwVqSu6i5G21yzslB5crJ51IELczgMv0rWvAdBJcw5rBouWVRN2J2eJb14svL
AGwcWBgO4t44ibNKhfFF2rzLtWtuIYo0HqpzOeJEn1ONxhtshdrOfD0sw6QTPEYIgVyt1HejziC5
BGKts73LRLtU3Vtgi5oUZ9AZQFGwnxtCLRbUkUCMFEdM4Lw6fds9PNsm1TzHfvM/zTWEGpSrMhe2
DolOCcd5OOTnwPAAXQUdGDMnpbkwfwbF7lvDo1xiChJpA9n6dfxfgdhdD3rHYmB8a+9pHq4E9D/A
8/wRzitqqyhgXKgwtgvXn7jQjixWj52LNDZm27SLc8QkJtUQAElIiMnDrW1egzhB7mqOJE8Ka++V
x59pC38GnwnoBpySBt5BsuNSl6loHB0cIK1REiC0ETcsBIErJBYiHECOSWZ7K02GGihOh7AdOWaC
qyDq8zuo4inaYXyQEmUdJoADwvjb35M9J1Rvtux6O9FUNA/s9xT+lIIMu8fBSqW9yXBdWJnX87Yj
nkvL729LeKhDSZO8I2r+YeLpJU8hN0kUFFz+v/HDVFzJu2YUQBUnzktjdm53In0apXWUaxP1U5oy
dLQ9yoOjL5eroO63ALO0OQV2lBvCREaty8J9rOKoWjvJaHHKGm5ZRXl6d9gKcC7NNBH76PBGOfFi
VkFeUWJ+roMUQVrFnvb3jT83Y9uOsv1lextFTLBfDGYAt3jXemZUX2FcGk63UdjW2UXvP6jZ4/Zw
PJ6toc12BynMlp8ilB2ZPWDRlV5hPuDIvCFfLa4oOQof3ZJ3mW/qlsu8IXl7I0QTtRkZcC631nJA
Mtf21IfLGYdKL9pQ3rUocZj9uRoeHvfHhQQAw40dM/ALgjmMPTcS14ieKkZRwEZZxOuxrkcyJ7qq
W/SlEEFcfXZQU6bO9RgqhVuVjBHi/lDC6N2dyCZ4bPIgHeW0o0eJyWeA8R8g8uo9uxrveNAChEdU
pGKbGnyUpKXd0WWkZSC4/NvOTnVp/GftLqoTL6WJH+MrYsEFHP5DkA/ZvIyq9BUD2GH7kswcSp3B
5GjZP5/A5Qz61XTvxUkq9waBR+450QIBRtf0oPvf2r/niuRWBRyLaZSrqb+VYH19Y6q1fbQeNB9S
BZdEpblgWH6ZWKmbPKnRpMJ4/yq3zJwJyFJTpHpxqsh81kUhizlTGE7hHWNGL17k6NjL9RpoNw0R
gmbsB4Wh4WmkJvhvTzj+hMLxIfvGXYol9Ma720R/witPIz03nM61ppFxsO0kWyuiuzTFyF2CkyHw
OndN6q2BmykoqHKqhFyXXkS/C2fmFxAc2e5DnpaSIGemoXBALUHswVrcW932ofL2IDlqo0Nl5WPD
7IS93MYUsnQosqBuDqYZ7C3BrIifzBGoe3mUASYoYgZ8CGX5mDGVgKM+2tHEbsu6CAXHNDQfh++3
NgKpZbOp43mqMJcZGAEKVSD2ehxBMX876Ui3fq9HcXFFu/2/d3DRKMqZ37oHWZbShzRrQME8rk9q
WsttzQoOm+ME40C6gHJWdZ53VVO/8k95nN9/NR3ecYUOhJ1NzQV2Z/NJCugBrPpOeDvLqe36O5vv
Og04pEpVVzRVALGwq+EySMuECEutPiADVbjenKjHC27HCNrwcdRCkMEc5Uf3tye0Pdl1/h1uQiyn
Uz6GPBduGzJfnm96PcNJQoRPZzcgrv4ATNLFZuh1dM1C13HUQF+ok4ZjSCiJudsIvYohUhrIfK86
PO4gTx+a0vpvimw0fIlC2Za4Mbni0WTDMZKf3TKzBdBHK+uolUdnI77kQkm3PRZ+WQ+vl21cJLyy
ilhc76YgFH8ffWBj3aKwsAd/4jGFaLTnjh+LHzrDGOimOxlX6akKYp98uGZ6hayUhwt95N87TEiP
lS5j3oK/sRtz+VrZyEh5UuUMQUXP7XjQlBsy3BCsJL10HiOEUXWEV8qpwcY9YxWU9Ox0YUyRZADH
H588+RUr/Gag84mhNlcwVLkja7GOtA6dJWTJ+7KjHewqV+P88xhzseksWe9YHxkL6jAFcVVonhBI
0ZAjCGCc/mjgjviAwgovV2CH/kXWveunsc87K2yLPHJzse7YuMYqEpp9ngXfuaHAmSJXnd0FKztg
JAO1uz3x/Gm6p8JZKMT/NTyeDeW5U6DqswsaD6t4yAx+hDLvCk506sLY+Ojf4mj8ccIjEL13OgcT
8b9JviOcBkvfgmro+ecoZTuNawfbrBrKqzAY50r+FTwf6HVRweFA4miji+Oz27p1WR2TnsgV0IZq
zPLjXTZm4yp6vJRUg/YmFlOHwufy0cV9J6zRvjoJqxR/naFFLxPxkVOo8LnJXQev+XxnapzejZAQ
3ru0Mj/414raIzs+xN2P7IQLTX0YTxIUiqarXDqc9s/e3FigEfZ9WDBXBAJWX5CyC7qfvclDfVC6
YTPJzs5lWEwpu3iEmNtTjsv9Hb8Lh5RYR4HGo8RZsF46fMS2ajmIlkKw090/5uJzo6jBv01y1fpS
I/oh/Tzm3x5UjDKCRaHKkcSp5l2W1YwZ+N8E3R5dsTQasUsEUWUjUev3SwTNPkiBoR9Ag7k4cQ+r
oMITgCQt+c3QzgE5E2egdthheRTbUwC/ss5M6OAhIyOn3vcv6KMI91vzg0okSu875EL8Rv4oiX5R
d4ManvgzMRaFlDN9L3lyqamZMoEfoH8OMJXvbiHX9/z9gJNwgACMyZ7q5T1bqugyHlKEaDpoFQDO
eEVrDaM8clw1U5Rv+FVH6hGblU/Ymw+nVAXdkD/yjjoeJT4DWFS3X/6rGfaLdol0YK0Z46u52B4e
O61vn8rQJkFZXrzEjCchPsJ55Eon6u20s4evfL8Z3Z1aYMT9iSW7cn9DcngUCkDTJi+L5O7i5jM7
uiAVgE5x/s1Opj13sbQo0Gcr1H/OwCAtNxdxSBSuOiCTLrmR+7WMwpJ47pHtZyD9t+16HcHUFmBW
U+fCx14VTduK278pRJWkIIot9wWDkO5iWRHjpvj3B3Lvu3nCR4PSbIMKLTYGLPzMuLYQGWjxwQPE
S/sZP3Kh/uRNQDIQz2LUtkOrNlj4KM/SzOtT10YF+NZn4b9jmPXwYFkBV67nL1Wr01Gb0bDPYoYx
tX15QaMOqetNVmQeV64/QOWAk7Veq8SJqQMau5GnWv7FJ1D+G2ZLW9OiOdTvraR1olm64y3i+2+R
DHq44FxVmXxq6g7Xqae9LcSK59LWrV4/H4hGR4ZzdtEgcbDsmC/O+EmhUaYUk7cPVd6oKuB1pGgq
e4moXHA03A8FhfrVm9pVExfr0kPul5tos3ep6A4AWEefJrZoVgPVKYiooIhL+FNxyeStnEpasvjH
aC/j5TEPaK0jTZSkBJK/Cbn5PI0p5PoXeehrFIcb1UCnGcY+MiDL+CmIcMipgKk7Nv0QsSu5k2yE
7k6CRKuPiuo8MGQTkg+Urq8tdQBhrtrxo+YdgHliLRiIpUBeH2gIIBL69SHex8LXMu+DbPfqcREg
zzGGL9scAceNddfBFQel8Xt6SRkkmkyeuAghsoe7FSf6zSIueCyKZdQlSWccqlHzQ0/bRHQRxXQU
nDDzVfGmPZpn5HWV1sn6W3BBZJhnK9HtX/4y5XpvaHb6izCYek03NnUO6IXi8dbS+OAsmWgGr9Uy
jFCCy1iBb7AUgY6/AxS70YaQA76gcqZKx3LejCIysdoKavMo7wW1/0OYXItalVpSDZFPQwpID07b
9fYYgHwVZ03NJRwYFr2Lhiob2FwUTntBi3V8A0kLpjTe9GRsRtHHWMdjjLQFNmK1ZvmXU3DHNnKH
/d7FyvKp72CGD7qkAJ8eDC6YqwgNQkhrSbrf0nmi7jCJKdgIO60kV3fAxmlk7r9TmBjPLGVwnopi
zt23mWX13y47ycD0OKc2/OHqkkWn/s8nExkdFnMFOXLcEYy0NC1/95c99LMNrV507OXmhcs94dn7
WGaOHT3Jgx/IrjEzuNSt0d0N4E+sAEYAaAUPGyTTH57i3wJUegIvmQJnCETIn57FjGKs4RmCdJmC
eAP3XIp1XxWjBNNn28mktWKgy8K3ByAl4wHOrq2I4N8FwdI92qHP93lwrFrUY65xzDgVaGijgiou
1yfzTV6uOXj9tB2szDxR9B/MCjGhAa4URvv1iid6vpCxVPs4T0rZ8WmiSLBNPKQLUOW9/jPzyY8D
kBFh/lumpkKfWTu8Sfs2Z9VOrYpIcF8X23JHCCGLRCmr3K2bOzjS/A8UUS3ruK/isyWA/75x4rq7
avABeCEgLg8+3XgQBxFhSZ7wUlnWRIqX1skS1gDvmL5Cs/BnAWjwxiDa2sDjRAEGILDyyu8d6Fwy
zjidyuiCpqKcINQ2pwvusGq/p/a9fwznrkpFNXyT/BmYN9AriWdTzO8oJMmrF/5YGwemQqQvac6G
UV/YvjQu7vp3g2YQisJZLGglYA6tt0MIIeoFDvJrE5e3YwsTv/e4KCyb5GbAaRkIlMeeaAb60/Zq
qEKy5q4G69phT2O7HS/Ekx20sD54myGtiLtQleQp26DSz/diyqpSd6zAUn1EGu4CMEMBHpIvDSpx
e3uaLDrEmuhonLY1moydn2h7YnPFoZSTEqWHLWEoVBfvE11kQ+Wmphjgyl6RZDi6Bua8cHyYZ/3/
5X9Q3gGIG8kRGddDgYitEk7OW1Xj1YyTZRM48GOfn1vEVna9kuErNFJpdX7Oa94MnThrRF65bYps
MrPIqimP33fbCv4hJkCgbWf5edZGU5naFpG1gQdebmKv90ybmh/j6IX7tNHjElIRW46+3F1B2iJ3
39ebo8jmA6OHABcdFWHcQnv/WzuzejyqTy95VGzpZqXSTEnngyWvjn3SRSiMrw/UOMgfpwpF1eQW
sbWx8GWtJJqWKEFv9Kb2RtZ7hOP6/Y24RR4XOlwfWNimGprXhNYP4sKThfi4CaVb1w6OCdLROXyi
g/vKmjlsepDKr+bKBS2u0S/Oeq4ekh/gN5+kqglj9UuvSz4ioK6RYGrt6/0zudCbKH6nGBnZ/vbn
fojPkJLRYCw1FpHgn/LcwGrZSnvfkCVsWsrHQsCXjgTrnU91WrTWxyMxiPWekKVWnND21DrQIM2S
9mZLwDMTBI/rapwZdMFks1xXdk8vpPc75nXikcVhy/I1Q8mYvYkPYtf8BtO5wKdFX09VILFkHoph
Hxv8wQfyCTANIEpFaFVeOJ6zp81I7yq1pNm3jpPSL10tiIugNoQ9UdiyDXFmoHn06n6wrVIjm8gJ
bMRzTuTxTUchKSwUBGWs6KNqVkuxDex4USbDMFSVJiEtCCKNbJlVm56hZAU3pTr2QeQj3PRAx7/s
8xK+PQHs0TXB1enkkkRTHWSpiqGnDzIks20O5KGwwl0OTYRfW84W/QOeLWTn2+rkNMpR5/F2fALY
fWE8JLiuwHUMAPOcCrsSky41MCxRV7TU/T6TdtJ6gwXTdhEepe4BL3pRK7GX/+wpZwkVUMHX6eBp
H4M205tKwjM2d+OlRVkvAokjHoY9HmDlsYnR1uKhK0fpwdbe+QqND8aeCAa5W/99omdSNmi+JqIf
ya4+D6Rw+yA34HcJSpOkYz/sAlt5uZ+B9ptE9fwL51zH+510VahXOttYSbs0nz0lFY2Ao4uz9POy
eyqSO6qkyHbwvIES7Ki76nt3I2OfksZH8uI22EODaB0MDhPpTyX2OHQFMog1YdIuTDpE9JXRJlBm
9F2K6hrZabbvHp5tLWCxog/MPKq1nK1TlX1OovZaYZsWuHsRi4qOQkcVVyiWB3hbpctL+aTVVsS/
Qs8hYgV59FB3ILjscFcE2gR6x+jZRMk5LweJYbYg7yIjrc/GYBwccKv/OfwMx5LwpRjNUNEkQi4y
OgYOgxgU5yUTdjt6QqA/2fjMC397KSzDAJel92sUV8tSRoQX+wQ5JmBP3Dx4got6znMlXu3iNRXq
ayAF5f4e7BOGTNEsc9OcS2xtjRlyQgTfl2MMrnUz510rITvEAfyN+Z79o8uyYopYRzO06nGX/5Ql
3MIAFQHVWJUMd3nZORS/uzSM2Ura/UZEj3R/OCjC1bQi0v+ZiGB41g2NEdZsB7rI5A2zWhMQdQ7d
4IFh/qVEN1i6h3tyPr/sObb5J/IbKBZM8iA47JNtp2sN1t5Zv5E90jYMQqXXAyHNv75rp5AnnmA7
91RkZny1TQyhdK76OMomrcazHlOab+tNAxnG5EhTetuwo91QNOdxcpL3FVy/1piGAhrDtisPu9BX
dQT5eLwFh0BHMdaevFos2U6Ar8RMJFXvChDcDcu2ZhG1+crA8vZKIF9YGL9H2KX4oB2eunv2iy1n
ZO/GqzWBgvyxqjgRXJeyBjGmrPjGgPP2hciC8XKky+dNtxkh/s3OyuDX774w30V4NmHO3GAkJRyM
/R2F3hsQYOEgXMyTob/Ji/Ans3HEMHX4DjKD7cgUdES6Xn9OQn0qJdY15JWfNr1fOtz7Txq4pOgu
OttWnyHNYHV7z5wqtFbAUcL1hMrqJKUwYWntzr1RZdXapnXJ0cW4gbdobkN4U64/aST2woNQqYlj
F/hpP/32giLGs9rly2gDyqmxpz0aedLZ+ElOFAg7WW4Rm9XA6EiqDZw+yxc/XsiDJl3QAeRbXRcL
K5AXLd6PAqHbSDV9yJfrZN9Vmwx95CzfOb/mmIOVb37HW+elPhyCXN/vyExvvbISSbtmQRVAXzaG
r2nCCS0e3QYPjlJQcvwVn5h1g/dISYMJ52tYZKoojMVJ5SEvINwngXqjhGK1bhdjK8J2lyhzLOrX
rPl7owc/WUnjd6b6xRovbXZw5qeS6QtbOma615hkbCoeCuTEhXS1Yf0t6xk6UjUC/AmpdvGecnc9
mA1CpUjN/LZZgxnLbZf0brXY3EPdPXysPHzLMQ2F+Zz/uOPlStL3esoXN8B8OnwMnPOGCKXk5YOH
Jp8eUDRon6Sqs3GMrMuHF7uJt4cspe6NTN0gqJvCuI12GZsFJbRAYcE9nRIExxrjl3d+XG4IZnXr
P16IgMYsnLr10sOKS0o7UpUtl6q/xIcE99SyGwKYtjfp4A8ILiNuF9eQ3qnQumiT7cTGZ70fIMyn
I39UzX5N0ErLUF+XwXlB203M7AqTBdQKHrDDvZFsh9b6leM5gTonEeEl7/KIkDiriOIOeuXxzai3
5gIEnMCK73ZoSYU0Xh2Q2omRU+ZckI3bg6p6cNpwD3cYGQtYg2MR2V5X3gW/UXbyD+l8sN8Y/P1N
CtUbi1EVzjELlvEXavJn3NbMnKaFg9sHtyebhwBoutAFsGUS2l6qiQzuES6zp1ZtqnoXSNwDpFTh
5RYu3turbV9D4GMMup/KZfSx3uuDGhw/358IWBRpetFmqXgiGkCMZj9yxnlbMOGv4wX+X/6FDOLF
BxiCM5uUWxdD5LpOiB4CJ2x/gINPxBwh+TQy05d9TPpoqZBFzmDYs9uO4hZj1A3i25aMzL4fnkel
n/j/WaAiKsJSjkflmrsVxdTiujn1ojpjBejwPxzBz2lf0WRyNrHT3GnjDIl87BkGi1SNtzJKG8k4
PgqiQusnizHzZ6HOg2ZcNAEMyd8K2y12mY1750dptH373cWGIln8zJKu6gvn6dfPbbL0KunzjfSP
5Y90zQREtMvhEQsNmLFN/6ArcvUV2wavbhHNF1ujy21uL3SObOgEN39wvb17sLizMT/40Z9xBVlz
nCz/C01DlJKQseUbSwId3TbrDkxWB3Q3Vy1/nEVzPUTeE1RB8qS9yO12y+uRuxJsAFqzkHcSEB/C
nuxT8+VkPvm3ACSevkrGJ4UFIh5HK4zR5a7HZhO5KQEw/GWYzNHJKQdnFzKz3AiKoT8nRnbtiCxS
XWFMBm8N8SipcfED48D3fKZ3x+ENuF5eGnbry9QM0AXldVha9kZvvFCsi62Z8xg2A7POVMNU1imU
qSBC9HALY02sK1jA5g7zOtss6uRgDwxI6VTNJAR3P6Dbg6dYOg/hFCBU//ZYwIA5mDIpxZwfu1qo
zuQTWrOsKu+Ba8eNYFeRB2hkib0XFc7OUDpuVqQ8i07w9w8Wn3omlX6uW4Hi3FTlxMPUPPFuPSTp
FCGmJ5yAUiaBmyI/+BG26i50weKci7Nssg90C5X+VoUoAisdJHs7zAez+1FfjgIgnT9Q11oqKE6G
t9K8VUTw0b2Grula0jnZegP3hCb9SNil9yNpTRzbugikW3hzashGE1BhOa9hMPAnZFR4OTA02U4B
X2YhlajxpCkdXMIaeR7P6neCcjPEkr97wJ+Q9R6tYu0cATg35orrTrriRHd5ON9QEu9Tpijhv2iJ
Dl2nf4uB79ivoe8j12QtUUbA/F9PlYofw23qwzyiE4mfL+5LtWGzGkoyscs+TD7soEY1JdCN8EoG
Gw0FnpAO3cNBV5sqWnPWq4/KZeMS/P+sgIiSU3wuokaAqUjDiBHzuL9iluq9BPpce1zNsO/OyN/u
EuN8ujd4HmueL5cZVXKGlLvC7JHM8n37jR4n90iB9kpCnIdQ+k+s0Db2bXV4rWvgKtUWWG7pfSJp
1u7rwRHy5BsA2BG0/Bt98bqU2HTrH0jMv+S8LSCwXBfsRXc+ThNQWORIBprvw+bY4zi1dZ+bz8Lk
vf2Uz1/f9WfJuy09U8FpU2KMIneHXNlQaZDnv4pMXyPDKFU9WnFeFx+YMi95JR+TJR46CJ5xu1rh
55tjjVY/5nZzGmZUiCMOtP51siXV34Tcbfp1qg0yILa5PXDXMjtWRJOj3gYiFO4/WT0IocU+kLQa
NzuqrYG+3B2V41dW/FUVVY1kG5lnbYgI3ud/kP5mfoNi96oWcdGjY3ZhauIqCQi3p5MYu4lPNb6N
jsiaUC7D0S+13lSt261B55jGxVNmKW7KD8Gz6hencPBZIWOUQzxP4JwK505qLHoXWV3wdEzQQscm
QN87n1ZE3c87H11+eFsnBCMoZcPm5+9r6MJnJNwNsxenkVCaN1AhkPA4oR5UWQTYuXv/e3x65Duv
LWVz0FIiUKJdtDJ8jBb97kMCNYbwlqr4zVXkK25P+h3ko7/hN0riYJD/mPEU1wc6vezPmNp/glP9
xnp7LiIODC2qxGnfdU3RmKzmIOgcRfNWjbBR9KqhqdUrgn2Uo9IMpTpwmxU4DeZdLyLoyToCdGOo
uVb+oWI1XJnhmmj7G7s3lW4QaJG4yBM42aK1TCCKlbeWBwVIJuq6Z/s/q7lmo2v36L1gZcRWzha+
JeIngMJy8S0uYx92ASKydxWtLFfEnSbzBH2ZEsnFIM38UGovfOBhSiMjZcbvAtSngfxnhAoEJyGo
15jbNI3czQaOBHxVC9Rqa8Yq3qh8YQRZlYn72R4sfCROTNLiLCWVYSbrK6n9eBh6XS8DrOaAk9KH
JTDke0f7zTrnhs4Uhu5L+GhJZxioJ54oW6Nyc6Pl308iwzjWtNrFrzlk6GzlVfuovIx1iYdTG1Pf
r54FYTg4K6ldUiQrrgacikA9Tpp+FKHRCl2sKpdM8ZgVluuEjaQ6COnfZQg+1WWT79IQP5QFW+jS
oLa/8gDVgP/tSYQNsgpub3oyjdze5TFXxaiBVmph5AIT5Ohd/qp2A02yu9v9AgBi2M84xPTYyL5Q
L7IDVcct19hamw7uH86vUII8IcgNHd4UJNgpK5DiR66QIYfhgrRgsIr9juWCbspK0E+0IaZz/5YB
IUhBo1ND0BeLUGRHuzvJ/EC1+sINUVuqK/2AvixgBDDiLrLzkTMNQMSkpMDqnwyAbRrztUlTPPuQ
T4cLiaHddy1V9Wca/GkulThuGzAsgNMgoNIJf4ck/wHj1+Rz6LsYww1oa1oRm0kft1XAh5YF806J
ThHwqngHDdAZAjHt/kPVx4M13HgIQTXbtN1urGfsJ6fTJw6r9CCSLu1uYGR/hCSYy8WOyh1frGfI
F3SgqKnRjtJv0MjxWlqdLKIQD/p0dnImJ9QaPDDML0LExcN0x+kpXMvsBkWuHECbfgYOpUztGxuX
YMoxPYv8OP5vDTJY+q2II1mcPVXmw1+TesjfHYP60kyfZ4QoWjQUZLndvpYuFBcfV++bf/MP0M0K
Ziur2oyjtrOKILiX8jyYWw+GZp7Vve5bQF0PL7o8XZ8aXUv2WXx1/mvz4vXvtQqqr3b0VjWs+QGI
oBmLswUyzill2F2TkxFDC2GNt7OHiTQjbvpguuMHaFnPUzLwykvMuIVc/QZTi/JzP4y/8XjKp3Rp
WS8LcyoIwaZU2lFbv/3KKO6YdL6XxxdKjEjbZ6PulxLxQB3jNREBdgA3NRTcbFaAMzDycf5f1ryz
qXHtOG8sMFPogcnI+s/+nCbnWJmoUdaK5WVzw5vDop+nhWN9uvALYCP5g48/4teGyT0wvJZE+Xbx
PVrvWMKrln6vWwOlRMgGWfCYZnsqr8ClyC5WASQhKSBr3Y2hSsK15K99hCmX6IOWhFriK418YyiG
VbAvw6oGhyLb3DTtHLkiBCjTX5G+sob/2Rno1vojx5/WMaYxijEqxAh9lYtmN8RtHbOxViPvrK6a
eJFkyGFUO7lWhUdCPdduNQyrA54b9XEAfIIulnwVTZaNJtRxiTe8ZMWucaaqtMDRE6Qgt2vp52U1
hR+a8sRfekNXHtQiGKfmPgz5eUcwfnuDyDpC5MOf+nO/iXn0Nk+a+KpyozgpMUt42u2dgHhrnUgb
ERW7ewFUSWCC0aLEpMQVN0zxN/KqmKUPf2cRaAqxj8kRvh/aO585u1Y0ljrB7q01T4u2H30WUTI8
li5hFSCLARY0B+O069MmE9iM30HiedJJn/xYriURNUSuRajy8amY7u6CukXoPCeGcSH2SJB47LZL
NJhAAdCRZ1PDCMFDsQc8BGkbe7VFJLpgmBnbHFDlO8jUr30PRc3RGH20QLs0GXyJXqNzHRkUINLA
8PiVY5+lKQO4gBqC054xRum2DFZe1NvZGwG66TDInA2ADLsXpq7b4IZIVppEopyuxLNneRQeDjxS
0QiCBNsj/Fc/iiNz5EV28bMOOWyyv96j9hgZUEE7/FFCNOflZUopg4bnCCwnKqhe7X9wOSt/jIfi
lEVjlpN2cbnX7zAgzht17WdvcurwSWcOR1UIOKAuu+olByCGSLoS9w2FnGNAKgAnVeFDdTCH2Sdw
HrA/bAO9DRqecpuFM2gzH+Mx6ZZG2KqRMAOubgoYl2W69Oy/F9GNvwymSzyKPsmyfOECngf+8ax9
JN2iaXPOeQf8MGIjnBuey0e5Z9izM7KIogKVbL0ncUTwqLOmpMH+wnZ8mQZsXvBSue8MgZwiWVYA
FwBvY17KmbsGyiDzju5YtqJFqHUxN1NaGaMJPMMyrjCuTiHw/1+icdIHErvWAcJhbTPlx+pWDegd
6VygW+j5aHZODN+OzgwoCUtE/H8a2A11Y/DiHYbLxkI5wV4aueKY9Ktpdb2zgOwAvBaXp1pm+36G
asGbB6dOvDwsByrdD1EGp/IkhYjFuyCfFGQDiYYFE65jEkZiHDcvgq4+xt2xKZhgC+AP2plos60Y
y9y/MkfkQwjhYMODWUi2ec+HwpU5k7O8h52oWoJSE0PWdWNe4CAoAxC/7N+hCVgtFLmWdvwd7SKG
DY4z7kB7hQwQ98IDbaaiX8PNyQGbXtgwy0vK1bx7gTRE/xaHDh2o8RAxbgc+OkycUAiV1MAmXXFq
tC/jgnSafLqqH8ZZszTEgtieMIVo9ePwQW11M+0LdR5Vo1qRojGGdJlL7UmHXh4hJzITuRKLMFyr
6f18zBvAvIEbFf5fADK6YdJl0UchL9E3rchYlAGh94pDJDwwVMMFoS6kfCRYrRpa/alFa9mEpJOy
BOmjVqaQq5Si+DcdAMan8GIacU4sPPahtDw+/97VUB8Ga6cu+nv7NGWFhHzVAvHUw9kAG2bl0sUL
5c6joIhDcyEJe1EIJtg5xXPVbEOVRNXDMbOwv2ACmTt/6GsNuA0msMN/BNy/fwFjCp9HqpxRRrBC
4QmLSBE7UpjQygRKLYFZRkK0eO0OUBkSvTld0unWwTmBtWrAlrHhOHDOHNblo3zzaOWi9pKMnJ6/
uHCjpWiUc0cwivnJtQI6QHhhmaiRKOUkW8Mb3l7+Qt02zgH7Cqi7FSaYDR5BoAsTEH0du/gzXiKp
Pq5L8hNUUdREv69YbPJzgHzW/Aw2Z8xND6QVNiFQzn0Uo4pYwJZMAA9We2aD1WPlZjwy7TcmHEd7
AyH68kG2ouKx4ajwfqT71hBav/RTvl0bCvwizVx88IUVqUDWeyMjuUlQCboIboWSWKYR58OS8Y4U
PD5RRQiLg5IW1yDDhojvJfu5OtFNe23EKzAZihtPDlZgnRdJ5IlDqIvXoa8fSe1TQ76s27tK7ZQ+
5sCk4pGqUxkhJHSpEdel2Px4wVHU/RCLd/bTU2S5seOuptiFqKH8ShdsYct86X3cg0JHkAE8zj0I
7VwKFjIog4lI+AsVU1mWZDE9CniC12QP2K757IBZDk0OXT+Zq1QZKaJIPlv4bAXhgLPlQdlqBGmd
+NgRYyULXv5SY7QuarsM63NG+q+NA7cSEG7Q1hRHLs0aoFN76lto8sk65epKjClggRiWU6gKjo8C
KpumklztAIJqnJgxmcYcCqPdWVsN/Dt7sE/aLlp0LHlvaZUx7XVSjKxX7zHGxlXGrZyrH+RscNPV
l51UeqpEKJ2ChVqOQANtiSuA/nyTf4F824xz8TTsyv1J6jTYTasH9/mc8GWCQoEUjekzJCD3cFD1
FTFphVqDiFaVQiV5UdDexQ0kCdVMlxTPBwgIsuzXFAWP/l56onkCJH30YSu4WblmsqFhSXujDZkQ
Q1cAJnYHRP0P047z3RMCnzitMQ77/Aj+ZGePTwl59RDQ0/kWuRZ0mnaiPfxWti8XEjZ5lle4Eu+9
BaywU4ghLsjKInSCZayDGRYjqqhhFacxDTwgdqXY4AKD3vxHTWv5hmlvhsxEFl2KYP3i26Rglskv
2JBRl7AIsq/LAy+LCBbXT+fXYfi+EXigJXpPsIFRD6zzXyr6dbDdhacBB7bKJj1Zmmc5ZAeOo3Em
VWzujhoBtdWH26swJQRXeADOdVV8/lU0oW2VxTn4YHGNOWIpoTwxEe914G1nZx2+ZwCVEGqBt53z
UqSlo/dzyQhobgrSHpAg6QXj/ODVa1fpq9j0q12r39AVP/L0798szdZRYzs0YpYOuP481jog5m0u
zpj1pBJUHffbtZwuDKyh5qK/+zUg8eIo+AE+B4OF88vJFJuTVG3OIW4LEICBDk15qPiw5+gB2yAm
iV9i0OlF/PanwOpmGidA3RMfKb2Z1b4Yd0gciL+orlSvmlF4DeUOZpngA+Mhowy5uMutbFw25iwM
nXiWjECrt6nrZ6LesTqcZGVA3I/0G+ZFsXNJjMGK7gcvq0n6rj5i/1f3yJo5htS9IwtjlYdqaqkk
fPuNZxtqT7BcyFNIRZgNZTPxuEN0jCaeniNtPTHOQaf7m+8ktLsl2FO4VQLfA73jSFlO7QFdtnZ9
ffA5F8SAI8HNyyFGT8dps0pgIefiG97HP/kLWEGkuLwssAWQcA/BD99JJEN0fQ+qsPOTaap9PwPc
6V/La2uMTPCrj1YrPSWVhIWwbm9gPK+Sp1E+4/L/ZPecZuOZWnUO3xyz48fmTgHCIXTCURJtMh/f
lDs9kr8mP0oL/1YHk0Z616GG/nOiASrnLJuRZM91l/mmTU+aZZYHr/rbcCRiGlRk7+Dxd9OL8pF2
V0m5P20BSSm0iwP6my7ucDF0+BgEdxCaKR2nlLSGkb8tdM/r/yFNT4b7vFnF9tfS+YdxFQghthq/
Jsf2Eld2nEDVnSAWIMoVFQ3ul3ttFlzKZPRmLyfhRBmlEuimhBIIIl1XoJyHGreuPP2Js5GvdBaA
Pw1FxBzOfooncZie9PERZmttPE5DCLtdo/wfgdj9ZJEa/3z79gXO+v+aUDp4g4n4alRHctar4x3A
f8DNOM9D1oDjYfDZQMJ66axJCQsrkXkmwIsgvth8ZwsiuWhPfM23XEQL6d2cAztLkFJ31E48kfk+
PY4GfD7zjJOBrDu2IiXN4pdHs7afWkkH7oaP8FKpgzjePi1TbPpE8gz9Gzysw0qAy18DyHVzIfwL
Z2EHE1luvxb4SO6MtRXFC6bLExFzVFc+t4anxecm9LxGmvO+09U2bbInbOtKwRA8dEM+eZTIX9xI
Bo4sprWYeT5puhLIFW0VQNlNThTIBDRxyTforrwSrCHYaYGNjcpAptEmsGkwxqcLd05t0vfjHdNg
hklZ9asQQIgrzlrf72bgPS0CpY/kyzL4DMCcmqdBzM/7pKcgzavAXhGzrQeiY3iUHF6Xx4/VarlD
Ps0p1KFdeg/crExUx0Ck6KV3KKhgdrefT+vzafAB24D5oGbzuwWAavetpl6cNvJm/ODvZKkfgPdt
H2hMJ8n6je5yUzwouqLilWZusrJ7e6DNaQ6Krn6X1VQIeV9lEx7340TyJrpO2m7EWaVhW/zuzT+D
WUv5nzG631NpdWlAf5ROUVFiHFl1MMndryodOWnOgt/T9K9pxJ5TYHr/bQ275Fh9P8PWCw+JaKtH
Xlh8Z3to2BMaOX89sclonF740urnJVsTOZPjlz9t/pgzDEqw2+f8u6moQP9ffDc6LSQL3x0okrJB
CLTOsN/ZVUAJRANEBojPf8k2iTAr8oeewGt5g81tZOp1peSuDqKq/2lE4xuErpt3uQux+7pj3LZR
dPviiTkPIOsjVST5ZASjm6O/ATuR2/8GhFPK2MF5YoBhMIPywfVJ0h0UiALPEOcw5OXiMbpuKcwO
YLQtze0lq35ikdgkd/65Wxt4NuUXz6zw2od3q2QIx+7A2Pf1O7KRg9zUpAV4YKTFfyWHIj+73TEu
YHK2tMzGTnY4bINu8YgE1ij7vE7UHiXfNzmizeSgspiqXkC8cppR0Vnq5mE1PrQq/Ey1F8WcY943
Z1Kv7FeQTaBvoEIFC721vytxGlzw+zty0plkEuECW4uDhgPFzKdKOzAgJ6uiNI1hZ/OSfrCvKfdr
xMB6Gurl+zmZFWqjkKTd98UCF0RHjgzFeVQvaZhe03B83dxryep/Q60ZTlv1neHZzG5H/COllD61
Vka8wMBwhRD9SpqwYt9G0uHcSVS/ZUO+0CzdceqzNBc6Nn0Xa8sT9PDjN4O5azKlivjJMIoWy6TJ
pgEe38kZHWN4kD+gPhHf/NBI6dOj5qQ/jsyZPG66+wNqmeM8HTlBWMRVl/ID50bDKF6oS0+KGi59
ur40BGC5OcJNhbAPKACgXhrFVqMcxGzV6Zgg6ZMjEyz+UfF1Z5XWqddM2/u+m9S+OfxM/RXGlgS0
gQFTmLtjQ/Da0yf0tg18p6EhEFiH/4rUKx8jl84xjsOvK/W8hHnW4hUZTtLbKdcugV/3GqaCOf2s
RzCSymJwuqxHdpGH5J6NgPxIczJIKdVd3fi5kA/O+BELkapwVBx/oMgqXy9GvDXqeekQ9SQClHWq
sCjLsL2Hgqsi6RsZZjGT01vYtoZ0sDyOsfV6r7r8RWYTcgg13+JndBn18hQiMx4J+qHzIWTVTErO
2w3KBsCyunhGmOBmoGhkT04VimXyOcpg3qnwrmxw6hERxGM79UBw7b7WPGsSrJfxXN+P/XJsWrgA
0jfxTU4/MFYl9a9FyUXmg4+zhdKpzKrHhKD7JIJqU2HzD0htVKCiHL7obRA+Gn0rxMDRJAsTsuAz
ypvQcX8hSIvt2z61Pcgqaug5lBHG1X8GgUks9cqblNdUf9NkFY42bNxbdZjdSnUcwwFYGMCI1r6e
N5WBmyXoYOL12NPjpm9qtKy8sPBrtLO9gEpmfrJS7EsKssK0Tb2b/Jo0qf+G+SX22blZR/3QyLmd
9ueoDUAMpa4qoxujBYliasX+ExgKR6Xc1hLY/AGXbFC9VqMTgUOpHy0KpHqowUns+6c4r1Oqr9Cd
LOO/b+bf9baa7ysccjGzjc+HDJ/gSrXdbfQa4SLlAXPV3uF3y+J4NIoJdRbBX0G82AuEcnCqE0Fp
KEf9uiajmT2i6iv2vd4gnf7w6RXlxKdBl/9YldTkGhr3IcfvrtZmt1orBfwL81zV+sWp+xCFlxni
FyFni3d1L0ixmjfY1zkD8NnkISo8RpFEmEOtR56RvZiW3aUiGJSlFTgaL4msjvEUfL+b3+/FWNAZ
jOs67zOkE3N4EFH+rJPJvZe3eKeLhmSMBD1gODhyX46iOUNoN2GUjcuGsnp+IOZ7tYiMMSpbbgRd
VJXbbhuL0MVRfLI279YEI1iEJmHYx6Dp1TMYelKn3zBdRplvpLGQnc5/z1tFkOUnUn/RspSkjUxf
I2vnzIwP8v7wTt4OoGn5HTBG9jQyRiPmy4sOn+zvKoJpxNblvoWA+mmwKamtXNtkD0ZtxPgZnXaV
gifZ9B+7p0H6mniCYRZGKQn/h3mVwln7MGMMv6A+yjGBt+ZhNKAC8mLc+AqTLdxBbjlafqT0/Njd
ijWlOFABnGTxMG5oizrDVt9AhEMrU5Fy/SgR5VNwan1L7Xyyk7uuich1lBPtKojwdyhkQFIfP3f8
SFsV8PJ7Z7iohfUbMoyp0cwkZpcZw1BXmC4JGpbxwQxAGGZOwrimBLMkybVQ5a7ppS8gO0DJAYWm
RLkiHs0v4MlIad1w4LUTsbR1X9dRCBnHBnGpu1ungDuVKK101y0UzEYPspUIR4o+kS3hpWQLP8LX
qvTIsEZlNolpN4tF11f6Ynv6E/YfBiiUuxacLH/neoXlU16R61NIqNPRIUsxZGWheX9YsN0Mrhi1
+tFIuN/t+NPUWN3dra+JaJVXainez8FlpbQv8tkAPwRf1JVsp1xmjw7oUa1CJomv1xAltmPGdu9Z
EvsJK8y3cOd22LwF7LoxhbVzXgDoSloj2nEwlo+q5pUQTnO7Sep7bLfFCOo7RVpfOqt3LoW9HUsP
Qs7+9dkwNfWnxb7k54ubZSBgNM6Q+2KNPzFT6iTo8Iwcjzkl/sbM63Q6XKW5zNITlpidDdhKivfL
yPxDqXZZnHuS+QtHfcu0PRREW0qNqoT2j/fyzuXQPH1JvPo+ThpHZHXj9z+6QV338pBYCP2GAQDZ
rgnadbhuohHW+sDAwJpaU2wDDGqb4iZLVkkYwlrbS/foXyhveV06jmLUHpzPvY210x8ku2+L2jy1
i1lxUD6rD4RAi/vX7C8ovUX9GOKpVDCFBxktsfLqhWvoWwlWQMXMO09wqq+KO3XvuaJ9CWw9r0iy
jvwrGYqcJOE7gmnG6HcOkBg4TDzSpHb8vSLJ2+reuTtJx1fOIer8sIcztLNOs13ljinbq2L5fSI6
Zewc2v5vhHwQCWDjZiL393dni+QH8eY2DkKog0keJ2f8azhltRTePUDM/E9rrOb8NcWLSslH0tNG
KkZa7V57NCGvO5uneb63DXafySXLQkVHDn7H29T9uOJYQ0k7x4nP6swVv+FlicZAFB+HDAYHLX2Q
uMKuUSKFWIvZbbG+Q+bFDNw7Zl7el+DI77lx406zToSFCLePv63XvLEC1f5ZkNEVhHd2ClajhWIE
4oy+6CxOoTeh88iY1wbiaJ4Tw5iNmbh69wWIF9d+SxEgB+7i3N69gyWFuSmXviy0GeZ711ZtmhKs
TiD/0GuzOtvDaCAMjlOTkYR0W7zVXQJzwK0wovuf6+MPVV6NCWFRx0cxmJtfhDMmes2hTylIeTl0
OkldcjAYBvI0KNNQSLA81HiTKk8Kb43eoL4n/MZy0C8sO9xBmP6ckiqUUVftPqrwfRSuyqfQSnX2
nLxGMAqBg+xFmnu4B5Bhu485z34ReBq7vSVAnquqD/eMRNkvPt8hNd8zP8/8tp0qqahEQC6u0cRk
wPKrHiurvGJ1yhnRCZfNdZUYECN9V25xYiOIaN7HGfA1j0PRRa9F80ddBSKUKGoBQA+anJz2Nrfo
hmeaLKw4i22VKSaLtRGHc+FHt0hySaqPQiNdahLt3aQTzB4UG3TQxxc87+CfqHfbU/LF1EPl66vW
6YZWVW8cvsvIgqPQ6Vi09B7Dz3VKo6QTY3cc1v9gU6qTHB7Ivzdj9M7rZ9jeF6r9xuukVc5qLhqf
vbFzjfoDImbhbzd+1zIIEWxSsDRp6MTw9mLWIrvFPUX9q+12uNZP8jhkM4Ca5dao0vq8SqSfGi7m
SuJon5VEI3u4d9iSR/73Z4o91M2oZWwwrdx3UEGv/IxHDIB8uisflEWLkjmNzeWJ/VapTcJQmFe/
hGkDVDQOCIPofDSWCm/+4zF15HMG4gdSUyrpK6mCoi2fwudfUha8vmLbzIe8kUEdi/rwcPeR5Ydg
fIHIXK4SzA20ZFpYtBcBaHF2xnvTBGJJXWaZtxKdLc9hfl1RXKo42orWGr7Ad5XrOrlRNHQ8dhJQ
KZta/Vj+oTd8p6MmFlc3IosvHf4nms5MqyVGzh8/3Xp1u7Nh5BgcrSxSrHamqU2T1ERg2vVap1rN
Ym1G8QnAoyOr7D4R53DmOIKRdNdbx69t8up5AVP+a7RANY5MLHsIIrN8ZTua+63CVjZkwWXaVDu2
vbb2OGR5yicALe8k2hhoGL5Yl8l31O3InChjOzSr/dBsseiPwvG0WdAkuAj4uZDWa/1ICluwi7s0
e2ihCpp/ya6B2tCWA1pqH+gXyeMBzXaiarChtm2b0ilJ8QjeI13cfkPGsjYre8QGOP+SqSyJ0Bmg
S1JRvxtPKcKad17OUlsMz+iG5oXrH/Zm6iz8yxj9uBJd7W7s+C82ODyzYiuL9O2UJP8hwe/TAbUL
kYmkVhkoifb7PSYD8wLsjbqR5jdnd6O6xYwCfu5qhyoX1MAOPkqKehl+oJE2KYfTxEn8vICBrIpw
r5HbpbpInarO2DJUV30aLIwDcWTAiXktAVAFkVbtfBLKFHcBpQkmmIakGot3IyELWZLWLQevQQVD
z6F73OKQeMmtg/tts1orWirPnSSq4GwP8XtJXKQnP7C6+j0qIg8bgleX/QnXqRNUWzmvfu5JVxye
zAZgeXNJhSnjvn8veB0iV9MReXdBryQgE3MHaP8r/6T9qS7bGwxFm5RYq8M/9pcYuDxXbMxgoyY5
zQa20bHTnk6MdTQKiifeZc7eBJWu9Z69hqa7jgH0pZ0d1lNnQfWk0HI0BLzyaEq6F2k665nunayI
ZOV4pM1RLEHPs7r/9f1onGkNqACrlsC2yZYib2ZBfunzw8dqqluuxWP7iqLLgFTRMYRmK+FM64Fs
J3xGWSFq7sMKcp4AFIXDozq3z7uooEHbBGxmmOeIYNnWF9a9wIEtXI1CX0H0QnqBoQN00g3chtwI
qsNe72vHPF8mlwmxjIZACQa5HZqyrVjG0KGQWYW5UYyOmC8OSp60GqRwdB9eK34KB77HEqg9O4/t
Z+5XwSIFQmAxHvj2gNXINhH/W2KN67pBIZKzf6HX42jl799n+NLT/lUtHpVaRKttqaWFTDApV++F
rkgDvCUnvoLf0NZqPuBNzGSVowV9NDHaaIYqskjTaIZ4gzxAF+Qy39JPLGgts5yxMrTl1+7QlhsY
U+jQHnBA3qxKcafamlvpRMlbqhM3vj8wwM9xfrZ896pOsoJNBZ8brbxsOootsV2WGhVJf3gXF1rP
p8HTSCvNETI/w5vLhl3vEJx5I0KJQwDIrMPrnF5BKNSZAK8U3rBsv7BiOEJJFaVkM/50KVlwkWhy
Q+ATnihRdenxF84d7e2Az5P0QDgFpXJyttNVfpsNImLU04YxoJF0Iw2Mo/T6jaV4ICQAsJ653ftA
BX1XKuJE8h4puZ27vhlg5dNtxX9eLXWlxT5+/B4bS3h5Z592kF7HJff/saTnHS9pNj7ZWc1nSMzM
KwHZ2hntqS0cN+eBxlJYbaU6fOC59dDeflwfi4deQTc5DBLyzl/ofK07pRbD43p8Vwm5R0KTDK2V
aVn9cFHY5Mwdk1zEBPVOmjcWjYO8//LM1oe5vAWY6TBEZVyQgeeT7T0w93Cz6gHFc27JonHErej/
v149AGQbJZHBn+loXnIWqY3pjU8OXDUM47hEvBHjgllxPiy2Uai60eZ5IP4kw12Ji76UdWh+llar
qi3F06jW0MPIl9FU9pco4Obz+3SviDUpBih66cbEUpcPlWjDQ0rSaFEDhk+8Ri8FnMNHUNPrp9Ez
uvp1zBqDb/Hf6/IEQVSA5/A2Lvnfa1tAv0gtJVLydA8u3KhOQkyU4DMBg5WlDIjCre3+g/KYY1hS
gsHfzdPuz5ZTCN52CV1K6g4sBVF9NHQyiDpd+0OvHIoPDgPX/G49HfUCFcae23syvBuzfu2Uzi1z
9zgtIDmmv56nmgw4xOzmnMbe4tWg2aLsuGHIuGZGoOTKGDd/UuY+BtTW1Um8F+UgSwDVn/HBYwfr
KhQ9M8OuRqQYoJQR1X6rILXzMJ8X+6DoC9Y/GrrizKyCn52Tj/dBMuXCgv7sTwihUOEkEutcjJkg
gMaxkXK1IArPBpFqm3q/l6+vGvF/9dmovgvrbbEVNB4pIaI7s767Wce9uaiiuWp5+iOOT4kIMOqw
ITZkGssuznDstG2yf46yRUe8YjeYCY/uux2t2m0BDkbCCEMukOUzT7uyxQloQoP2040DPDVAtBnb
CdqKtHC8Oyl/yu09HqY4sZgCSgY92ztqBIFDDdd7KHNnqK+yPZmydQvpEzatkQdDHMH0hZXI/AlD
eZBQWuVjV5aaXrzS1Y8lgDyWzMwWits3DNra1gyeO4wse3pP6LVUErbHMQuwql68EuiZq5vB3MtX
FPtwEOChHZk0jE4u4Cs8LsgxGbB22k+OhaiL2ffDw41rTZedneqk2EhDVgvsqwwKP12OKZD3n8C5
45XezmswxhNNODHSqHfsMbqDb/5fBXk1zbMCoT6TyAauBApb/jg3f1NjnVSnwNCro9VTdL8g0Ytt
xuohr/lEgfk+spBUMKc9N1hzcotMio03GpK6tzHJN7QFB7xRsV+bcxVYpvoPVlv6ts5tSlfnoMDy
SjjG158a4zBK0YBfTB362IBVeAQyKNhhwXEfEVNh8FYGgJSp4HVa7nuu42+bUaSofjWVuxQoS6nl
riJTHK476cKWXAB6B48Di38NXCKXjdtDXHkn1TZXn9ABj+hFJDzWvnQAZ9ueUgHQXc+VIAoFdNSv
7WiLAYIYWQdMI7S0birvMAMqxJOCFp1iqOYAaYppGb4ZODsc1wB3vPvElEGCX3ux4c4RFvqLnckX
fxVHRBmB3P7AIs7DZYQq9KGR/Es/+pdB/8/nl65NBwmBwVs0QLP6zWJJYK5khqRVFxQfnaqo3xvF
j3zhEjcitdZSuZMuYh+jbKWJSEmUxCve6CT2UqYG8Ln8PWxot/zP/T4cPIDDbncKjUkEPWVbmqRx
5iqM2iZNS2JcAzTIDr3dkUTagWYO7R2fl+vO0QgyX3IvnFZsFwiaB8V6u33I/+OUO+s5R84bMWl4
CWvaaVYAEugq9HpST2BupSKqwcG+frbBL4H3RXcNgpAoHrLiI4PSZSVuQhnOnBMjgZxZE7o0YhEu
qK7AcDFXMe99GtuF/ZoQ8ZndFq4d/B/yyXethKX8tiJUCYW5KzyFXDBulc21gNYfinfFpMWs3k3J
PonbWbz0H/6iRccetYQdiNXFytyB5ygMHSSceP6yv9Dq/lF2/lT6sSdDkjn2H5x9zjWwe6wIfUpp
7/AcD5o/4N0PL7E5AgAfqt0RmfgirKILq0w64Xxf+AoZoLrM/kGd8OH1pce+EPp0te49EywsLwff
7C2Fr/EjKEiGmBJmEstqBxMz4LgUDMMGIBUEWrpEB3HGqS+tpzuxIuJeEpQIMqoCEgO37NGxHKgs
0B6GZOQrWbvLpMWBRH1is2ULUOAUrjU2TUqF3i/FRLi/iDVpB2g3XoffVKEGMJh1RB6v7064PZJO
pa4WlB0S/IUkNz3RvPTb69SfVdMlmBfQSbz7yECDjmuj0St22c4XAc0xlpLdgbRGoOZbjhWS/Cn/
NyWxyCo4UsTZJwkFSY8z4fYp44bhvhsD8jkvNJ2xl4Uw2pTQpjrijriQ8dPZrkz3WUk4sfS5+Q6J
csXoNYaNf7uLlNOjtuDdziokcOSjzzWkEtHgMw06RNsZBc5VtNcjG45rpwtCqYrFAjekRMxP1Jgq
iuGEyGH7IKtFmo0S3szUv4JIW9OyhDnoYlpBk83ihWGwb9nDYG7EpIIgTcvpYy0Xebw6bXrE7sMV
o23RmziMgg9MGM7wCYxULy9hj/Oa2vFBURc24C6BUUiESqSC5OhDb3J4BadOwDtHm111ZChHaofq
XE4qv8G1bdiY/FWQSV2AxIunfbZhHlvEEodUBKudN/uujBiEfSzwHq+BuV+7MkoA3RjLD4jPIbqv
umL78U7oPk5aOA4HE3Hgk4hvW5P/n4qFCnwyA7pl1MT2E5o5AaraipetEYKz12gFSTYlSWEKGu8v
qyrGXL2jCp/PEIKw4QaN4oC17VCI1xgvSxXlHHiBRNRtmJPwNe4GY57tEQgsreyMuoFnFLiQYnI5
SgParc/zI7oaAs0VNQeBXQd+KSiAw42c5OlB3HwMsYpqQXPUOYxMrQn9jUufFd6+wclrvgweQjDZ
sd9Y1xKM+LzqakJqAZH3+bpFbWqPSql6Z8oqrVKBN5dSByOQSMhctoMw4cc1600cyURBkeSybsV1
Omq14CE5zBP6eCF12WCThSqd7sf9xCk8SfaEehIAShtGYvYloOa89TSb4LULmPsv2pYbYxtlH+nw
awsIagWi7Hf1q7JaRRRFjTN0QuKJUKLErPLz43HOFVyj+JFN/H4HzHDUBLOMB8Su4bvMyl91DC5e
uw4ZlB9PUhUCnLQvLHgCOEq06ljvcRCMCvLmFazQBa8rjmrqDli8hREk8TE54MlX5y+8uW23ZqMY
yFFPTQ5+8JaNNsMFY7AXFQzzHv8LvKJUDYPsgudiBQIpEKWhNJuFUVPUoKW09mNTs2b3hhCSLDVi
bg+YquRugoRjiOZ3dTIM3hVC+w9oPLBgCiZAfpXzHi4jQKw9q4NSL/rD0nfHEzUgu+G8JAlzYMwE
1UUeh2NDXKKwZ5TTcFRG9sVUWCb0llEW4ua0/UTCBhDEHry1t9Y0NZZdin5/o2x4WV2Sj5dXyQ6r
p+Xd7uX5FggSehn/995tE/VUVN8Bc50BX+kmupYw6TUS7Waf0iUA7uPRubo54FvCgbU/rmTszrYl
B1Ywv1Rt4AeVau0waHAbPtyMiG2vS/4Fu+o3G9LeMTxGsgNvHvFMEMRWchNbLxU5ZtU1Qa3o8WUL
VH9JtbCBEEQpw2Uj+53DvY7sxDPXZVuqJfgfcv1wtxjPAXI1WnazXrzy30B+9QInvlUGE7ykbAwN
SHW/koVIEaxAyJk7w5w2vRQ0ovGwjVUV+ZJ89GlW9jeeaRWfzQjMCWkCCbENMjT2dGtBNpzG47zj
wgzC65nFauQJ8iBdVt8WEvXpZokkhf9FWBWMCQsjO/GTv+CuuEu8x1XJphY9bBGzSbVo240zQbrR
w/F61lwRfOcPej3MW6Rl4fenbkfggxCu2hA7bpmBoZUheBukslIv37AjTjbcmyDmkLdB13Gnuopo
tlJY4Nl2ciQAqWNRnOzFF977djz20BUi72MaJnRkh65Nusa7QvLlqhFBVTUqroVnI0GbSR+L7bPU
Jmt3TFw8O+/6XEMT8Y7E9+uw0CCkkQQG9g7yLR9Hf3Nvt+HQ5tWNVsLSErrdISEHR6JpPK13+tNz
pzAggH/1kkD17cKWY42kyGM6NLTbq3Pex+1WCaVL5f+W9XNc/MOcNTLLDG0yPNdw0aS79LFSbzjx
KPxQKUmnugdOz8gkA1Cgee5+fmBNTQBq02p043D/A7FyWF2y91qa5fRZMSq+Tx7qHkntOP5hIc7z
jdysxngJ3zvAP5rmD1COMKN54tO7ue76q54qdfzSoNqSqRTMVADlrg9taZ2eepisU0yijLbH9XuX
UDSCMrtdvkvRcl41GroS9Q/J+R24jZoEuriZkgaZtUVVdYUmo1yCcqWS4f0k3Kkw8MqmVuYGgoJf
f5fLQlp6dnFoGTKH7Z84Ht6aw+OlkMDPsGeZ9Q7NC8mUTlKK0+5H99KzCp3R3uM0oLUIlz6wF1/f
YsHa/DPZ5xQRnY/3KxBzWZW1ddEiLjHB5NRZLxH2LWPFy7R7bMLICoQfSXa0ahxvESLyttEa1hY7
x0Np+HQUDFwsOxSPm44LY1SjciI97Zur/zQosPaaqVmwNiWJputVQJIRD8SGOml+zWrTfvcKw8+j
KzTsmx/Xt0U2mwemqM+zheanDmmO+lBbRdewXRss2FHdq/BE+7a9J/bmq9M9GF6oLBILNLY9pi1P
+mxDERamRHcWG2XnecYD/piT1hkHtFXPqVeE4X/ZMkjUlsJbHt6M4lX3xWBOIkKvy6UCq5oKyhzm
GCfcgw75l82sJg3QJHoSBRFeKeFX7GXD2ExvXONTDdBGGlq9gZk/+xqrgObXirv0nvoYiR5JdZwA
bXC3KnHcJhscWE/p4Zbok6bD4on+10Z8WuhgWKGqR+KLX6JVpIgLvLPQFAWQxWe3wsv6NprLAA3i
2HRSeKurJmc54eEiPX26+XWIIPgnw82lvNGJA8zcETAnAT+ZWeu9Hj+N67DIIQkJeJO655ygTfJt
b0iHFc8Yr2Eqt5VKQKNiwZK7/DL6C5d6fMKKTriTORLbo5SBKqbq9YuX5Ei5TpBrQOrunHo91J3Z
3lcPuafdYz3NVuUdyh9S+tvy8QX2Z+dOKdA42eTWOGc+xzHhK4cKjgHmfagxj4ZdXyoyp6FvKNkc
g6v4NOAingAtEmw04Hq+JDHq5QFbY093NTOkyW2j/vxBKvoXrpi3FW4vPX/h5XUIyQ/ITs43a6a4
OpVeR8zLQGlVA4eFwtKXpANWKUVVT40oltXUmwl1kvA7iKq6lOoj2RFWQ1w146pg4DxXCtUYYiMm
nCH9KiS2wlGUI57wp8tXuB8/s9BYcABTDPEdjBXLaNwdDaDs1iadZ3Qa0GutDxfXCkiede3MZNcc
XV24F6uaJ/oOMBH8P1eVUtGlMOWarv67nTRi6bDydbAmnUiEurSQ2GdBpZxArZu6jhdcK0oEl94g
ufVwIJyoT5U/mX5lyALnzhuM3FdKBEKQgnT9BWQpZrdOXSrh51yJsq22XN3y/xtJZvh5SrPLNPoj
TXwvZcEWeNV1stMJs/uYv0uQampt5jlvgMAUthYw8+XC6vojyd57BXj99L7bbNg1op25gxOqFRp6
wsLpPQJ6MLOfz9ngVOAjHiGTsXa7UDQQ5WJl0x22dy/JOLQ0ir8gqonNzcqw3fzcwh9+cVRQZbxE
YtWg65eg6gajKbhu6JY94HBD3W2I7dBeDCa/b8BM8zRLCeGq26b83VfqGhnk7cei10b0juic/+HY
zVQ8DlEzXiqWDHz6Zp6dH/1MPRkF3En0B3YQx1HP3IP/W3cjHBGVqL6gJnerTlCZUOo/BpHD8J81
nvOcEtglX31fk91AUozg77Rv6zRObtOCAVwkaOXjolsvK7qm8fAk2pZ8XLQerNDHE6oUAeLIMgxW
0r9PdV5CS+OpVQcPhQZFgwdmldfQTGy4b8YZra3ELq4Grhlgy1fp5r8T6WZm2Up6abQXsyV4aCei
OgLIa0PNA9B/Gtd3u6swymOMQp2Nwkt6j8qimeNdRQDN8oRV/wkYEsx6rmi5kwJrlkCTYFOSPdZB
0p1AbeRCH/j/M0IFs7jfj5We5CstHC3H3SFmRQcpPeZeW8Dw96Upma1+TZ4UeMu43zsJ811h6LsJ
H1Z9xCvf5N4X7X8BSH8YOj/SJlqeXHIvCUls3cY+dPtWBTkMXgZ/fBraHfkhp4brmQEL7bLaNIZu
9KurcOB6hbeT+1c91nzjwIT7IV7L+VFkeuUj1X0wlrekoPUliTU8okRU3JH2KbSTGzUpaQ7QGpS2
PhPu2RVer8pvg8l40fX3PO1INprfxcMXmGGTRw9Sjruzbshj94+MW3rO5pl2nC6LC1pcIbUKeNn6
mPQdzPvYqw2WcvERLGZHKOszCILWeyFbjU8Fzh7ior0VqOdGha2x/T6JH9MGbL8NXd4sCq04m72l
LAvyensn8hT04IAcDOSq22GZlenRwZHPT5k/IJCOSR2ixw4DaB+e4QN61fqjeMVZ4BukOeSLvN1i
g6HNHB4ns+DTBFEwQ1ydZrOWdl+JRDst6lkeZoyUQRztf9zJ42T9SRepSSoLJ/seQfPf3h1HyOTM
CJYCQDn9YSIOZSVP/wo5pL3FaeVm0/uRD0Q38hoytIfFdceuxrZC+ma7peucfcblDh+Ds/2IuLvt
GWf6R+o7amkifEhorGmQtNLis0DxqfTyAGWhCap3yNdTospdot9k/qp/ERdlriD0i/nW8UaE3HzB
5EroicPIH9sSGtEZV1fP17i17l28UjGh3sENKAEG+WryRo2EDTG7pEEAUmg2Jsj16R3NBywNe3dr
jmL423wko6E3i7tMgEoN9vGQFQSKKAMCNsU/0kkGBeeBPYvA2QYf/DDjOsT9ClCBaXOvXqAcTH02
GeyVpXFEr89O0H1DpbQWuTLja1BqmaExOD90yE7WDskivAvl7kN0kAub8rCthurbiI9ECwOUTQ+X
HKtetj9NGRrnGokpG+hu9sZRFc2kLrxtVgQSq3sTsi7jtSP86CCOOR3hGjJLZY1ByFs2/d626hAP
Cd+C24T1DfjPpf3DI7PukfvgNi6FbsQeL5ziMEnQgdeiT/NUCt1vyr5zkk55+3ViZkOU4ZsUsVWQ
jHNX70nr56XhKVx+RpXjEeL7fA3D9Qzgngol0QJy4B/z3J2LmDhNpF3mNXNWJp4pe98+rwhPzwYz
u9rZjpeNkc1LzmDVTgU9UtXyB3PUTrgjoTFCvhLNb7kIXsAoNpz3Q0rG0BvESu0HNTpp6cFvQk+K
8678RPNnHFg7Hh8UuVuu+/kEpx+auqlSJKWMoc3+ALOsc2Kbr7HZqFqPp9aEFsoxrv9Htm+pU+Up
nsmK0bQXn7lWtgvWMgtsdNyyqupKaPIHyJYe4WNEnrz5QPYShTJjwuSgaBXsU5peIsLBNch8yRYP
XgQOwZjZef9Eg2b+po76xJZU7mp0teVIjc4v3oJuXwj0bu5MccrE0S0QXk67SxSihR+65S1KwI+g
RT2KVdD8cI8m86cLelfYQUu3QYRtw6zAp13UyQnaIKJrkYOqtfqPBmSgCrF4J9FKILKiex2oRNYJ
FdeXHfPobs+EotMmeVfl5ka3Gyim71Dhj+3wIJ7emSJCqu0Xjw5c0UhbrBk+estTPTtWwckJ/4t5
CQ/GO9EwH3TmczTZxTkcxWcz84hPYbD6mPCtUaPUkec5tOZD5Q+WCakTRUYjJtdOaxXEml5oKJm0
syP5OdF3NTvjknT8qjrx907kMi/dEgXT1/as11iL6lWcKn+1TaemPjvdiBpgdRI0t7BFOZ03rGqU
x6KZ4xqRnUkntul3EbaSII+x+0nRkCjo0Wi2PCDd1v9oJIQHNdOGw/SQKUpF+VlXj/q38UWKI+4D
7V9KEd9RTqJuk8170uNTW49c/gscY+5RRmE1blGrZgrjwpsFcCK7gNWGIwgg9TG2uTiwJhZr+/09
PI0a00OAM0hX7ZUL6gGgbpIRxII3Rc6TyDeyEXEee1+kxSuFn9Oi5BTQwb5vShM50zgFzAaGtzBE
aTPejaHT1G+moegam20zm5pD4J9YxB7hkP6g3lUht2c+7xkoDLqQnoxyIx0vmc3Qg50HcE1RNsXn
HGquQU5Vztyh7+LH0b8Zry9lVpebjmSpJP6/9Y6cycMKOOc4Nswi6AD11RReNJc75qMkeXFf4B0K
fkWACx6vLiFbHxtYAMqWBwzI4OWtKgEwJYeZZKLYQKDeT+ztt+79bhqejfJ3sm1VoGpsjb41QD/5
CBV2TXikKGGpYkZYmnwW29CRwzQq++NDg13FEiEqNEOyAiRHJq3pC1zLOUcxZkn0FRBOEG9EgswF
SlqyuAKJaD2W+mbz+0QR7Kx3hLjss0L9ht0bi0SJlXmNDgy6D2oiDlkniemkkBAKxuffF+cBAAuI
qLMZM63/P916L7IA/8EkK9wKSPKxFR32cayQbUEShNKZjLlNOBRCEkkST9+4vvtRwnd89ilbt7RS
RmudZHJvSa12D0Hai6ZiZwDXYYX8Bd5aenWbB4d457HSefYVFrO/y7nKGKnPKntSdGYXSoLWSYsM
xS9OBLFxwK34WSFPhc3j8PJ/X9UzwZ9KzAo4HQNCHqRE+onfbQnSJRhnH3Zfl/F0Tv0/1/ANuyRT
j4OjdLXpwJE46B+SQ4wc8vvnE9YYp7mz+sDq9r0gt4/BxdrwTlwo39VzfEIPG3AHQ34MM22Jt8KD
U+hSMjLIZHZ03sTy2jLtR7mIZ/DS09l4FC0EcBqMTC+3pB6pMgqnNo7QRsNs9CZ5U6aHN7QB7Wjh
27J1HW0IlIj3XCyZJCYUlu+X/5SQ4epMts9oyDminqV9itMc9nrZ/sSG9cMtPOaHTz4Mx6aNqK4N
zqHvAygL/9ZhDUKjdNx20yEDI+jdDMP9CkQ4noZkpN8GEUsl7uiWs4A7kTBAjsfCkCHhUJ76cnFH
4ASltKnxxQVKgicYNs9fNfrPO2Fl3BNgsb8c49jMd8GVMP58RRWCdkZfahwgiPuXCroltVj/x6JJ
uBtnJw3qWIAE8iDRVO09WVjn2kR5jc1en5aXXUZH7irKJN/kzu1eUWFwzcZLiB2jdNAiIbfCHDLU
bubpLgOmVzh1FT7thD89nt5zJaUd6qSObSoQtciaxiYhDogVjjaB4nwhLmYgWH0QYFfHjytfwu6Y
bpLqTpWyHyaycljHs31E7za8WtpRz104n7k5/chXBiTmK+s65Fk0e6HT9Ee3X6ojo5uFbTN+EamA
dPruwyyX5hdhmqY4x3CqnDga0s5G20YzLYNxKotT1e4jfpKjdoT/6cOUiHc7b6Y53DrqsbURRRVA
LQmFPUhis/+JBQv5R5++LY549ilS9zDbn9Q9fp66QxXWV7ah7PFg/UK82VXJm/evkOc513/z9OO3
o40pMPv8SP4tQKCOwZwTR8Ekb5wk5h+rh9HR9Rp5/QqwTrUd+AuyWSNTjlvnuJIrsPR9jl+Ai+h2
i92dMMTOIJKALQLnLQqoIpoHXvcoV2UoI/LBNvZ2u9a0mDhuXAeUhqltaGf/fbPpFAoRiUQoFNsq
yQhH7FXeMNowhyTSaS2Fyx6bKyXJPdbeiO+NiDBXEQF5/5dKj0uFksM9aC+1+xua54vD2EvLmb/8
jvJpVzSSTDewcMG30d7baQ+1tDX++hx8JQfLeJ79EAdeep/3KUPOJCmLDZrwfHczk/06WrY2sSk/
06TuCn1+m18sdq1XPxNeEE+PsRlqwRKScNcOw9YOnEB4GZR+DeZ5pp+GDlP3VOqgZo8Xt/el0vOf
0/g0OQMd6OUIykT3ErGUqTJ9zqivNQnb38nBVBJRXVqLYxXGFBo5CFY5UiodDAsTSIGFb94YyOWL
PI81r0YB8044oI9vmd3Vx5r+gznlYhGgGhQQz6NThowJVxgffYpOG4SCAVE1A1Eh2TBVjQaYUEJB
+D6GF66jsjkBJMOPf38e7ZDJSbf+CvbF3szxPE+rPo1gJ48qxRRnSLg99D2ssfcf/g4EIAkxknEI
P3u9i5defX67G4SggJAbYGPbi6d+I8yYDC3arClkGiB2xJ8dPKOo8DTta+MBzBKj96Gz5E29yjBs
xR/se0yLXExGHrdOUvRt1oI+xb56lkrF9IPfyC79XApo4pamxKLy7bPAkN45AqD8/otWcP/L64Su
JPv8GUsZ8MwQ8iAdOyCKnms7cd6mgeBFLMjVHu5ZvbyMGqrMO0Qrwt1ZqGGyK5shbQOyHDVa59Ek
20VK+m3mXSD5Rm9hDeQoJKaV5M3a2WzrbH2mHWWcojh9CzSEU7Z24J9u1SAo7PSaT0lZE+l5lVx0
h8io+pdwXd5mZkHcma+keh5nCzWFHyyD/421JoWtjucbU43fGLtMcj/snGLQoaVRaDLXwzpnLqHw
rYba+3ScZXLG2oe/lhmvY5/JtLLYCZBp50dFokZ09e+0vAqNDNAVNIyqjXJPJRrRrqKbJh2MKmYv
wtWdA2pxLZNgHuI0wDxogIZyK3omypFFEKp99Pxcc1NfKpKFOHd8DzrEc0U2/7XsPQllu5NpDKEb
v7i1pBDQ6yNRUqjmowKPOFrwr2S+c8LngvrXYwQzmToEEMNFDlCiF8s628mlWRjTcJK68XL9YoOa
Q0IXY6hqglRcO6xG7eFFDwJID0RKGSAydCR9rSjuNQ/u+a9difvoC4rgD8Cs9euev+mgESarAhlR
l+lFb39B8QEVBbjubynWqvbmN5zkshMg0FdHWKi0SlJ9aL1+Vy1i9e35GvU8rNdBUp8dCx+a6elN
GafDR+mQjlJ+EHx2e2lLWF3V6LTPCmKCQ28AonrUzI8l04fEoesjM9qLOXekTaNUUrATqph7R27b
5wqJalHJPwcJR3zMIuB9ldEPuLQhU/PwoExkhnyKhp9WA+bRCY9fsnT71rMJFCN5XWlCSkVVJJin
NVPQV+0bkyDufQ+bxheV65pnUlrXyTnZk9n1Zi+VqY3IBP+A3jkGhMGs1D4IUEVoakokIrYkt1Og
5JN/7+U9AWZTVeL+9kSqTh9kfKShRPdYRpRasixUs/77gZOI7uZNcVBus1k1nJ2iVM/WL14bznST
dB84dll0Rma7IO0q+vErISXNt4HnPoyc0jz3FJ+oIz42X52p9bnz+jYxtl/ZTxPxN0NuykwsvoMw
0Np4GFE9XmHH8dS6W7YfyA5rhxmHyF58wnmXRwbYZIsUZb5GKVabBrvRarhBMyR/J5nGjnI9Gs9j
hPPTrB9QkJymtIctwsBc+cAqwS6iP2bhOu5cse7Hn2eOnH8UV7CKaksKNXiOnclWgRdVTqomjSfD
Yf/F79Dj1G5U6ya8gtWJh55PGFiTui+GgiApsJ8pF7RO6gpRUWUlkRBdotNdQnwrg0wyzgQeYvFo
0g5UspYnx5ioOPMgcVZsgXXrTRS++oc1dc9ryIphCqkQ3cWEqshKn3A8/mT7Z5hneI7V48I/pNLv
ODfNFr7/d7b4i6ej1dYYIgH8BQu0ceUZBRHC4Q5ZlMqY7dfeI7JIGhIih/aYiq3MtusWtCRc3MXi
IPokjIHN/goN+fbPbqCTcWG1j8ttdp2rZsg4gpoTexIdVGcF4aefRVf0Hj0FSKX9ybCvb6fT+MdU
be1jh9xAtwhZ9m72XiBjiwyitr5CZPdP1AOps0uu4khB4/RfS7QDQfvMZ6lwQN+bmr6AEQ74a4oP
agY0nOUirMCPJUK+OgxxFtNzs+U2lvYBpEl2gI2ZHc0RvBcaj+TUgYbKkJTZnwApf+bsawTgoQx5
oMvg8LWsDGLCv/XTn3N1KgEaZNsZPzl2tlzghZfETEeKCrP5OyQQvVQWa/w+Ee1iIDk72+F/JU6h
fWgAQTPEMqDYZOKwC6rRitydjMUYKcEfqudbA7khqgdKhgh7Cf7GQdeeJyAfHmzXpD9q4zHyas26
B5xrWrS1lRP3SA1x0hKG1gN/VriG1Fsm9a8y56VoHQzLRi83z/tcD6kJTU3vQnfwjBhGvjY6FENE
UY6A1cF3CpKEoqS/DaI2271s5bDwXYoxGjPKnhYFvLx0zJVZ7xrgecd29hjR4Mr3MqT0TzzDJk3V
5Mpwl9Vmkcg7rbxLm4bc+UmTK8WdOJe4d1wiRW+ThUz5d+LsZtonD1/OC2q4HHbXTfB/doh5TEYh
T4OQD2IrMdjc/Ny0DlB2vhLjnRkbC8iQaG9PWfS5MYOLU+ByQzox5pSaLTgj0oYUku443bt9GCtq
Q6MUBdy1YiJnESK/aTGhgbtUq75+QaPGSniWHFAvsL+DwfN4A79aFMurXKjT5f1pO9qrVV/mk0+0
l7WdASf5o2AiQV8zkuGfgvarwiVTetILrU+c+dgyA3RE7k0iFQL6cSUNyqDaaJUpBCyGucqAYS/w
SfTZlfSKf78cx8Wc2bv/mOzPBq0G41Rtnvypd0czTX6HbFU9v0FzNEQB3b5Lm6JzWGK+E9WLzowj
n61CmbaceKeO/Ern1CFNoovL5JAKaICqgC3BPEIRo326DDlxVnE5iW3irZBCl6EQO1fB/vsaIl/l
YxavKu9J1lAWPZZoO99XoOxigKFX0qT/3efP0PKkdNaw4Gnmeib108T6pVQrcP6/oMuKGflvbVHl
GpVLKIsGIKr//bi05K4uP4JqToiYky3ziBWEkBfalGSrAqgWykYnWAl0nAF+FJ8l1w/KULmld7BK
Y1P56vLe7Y13s4jZk+gDvT+8//YKtTafYChg2Ta8EEzvmpanjSowPiGXDbkdPEddPg1OEsHz8IFm
7+GuTUW5LCF7ScGCig1hmC+ecBWq008XKshxVLJYYsRSF5CT+18HdlhszzMl9vdl3wXiNYm1pOpJ
Ka/3CEIyqtPAI7nWzUyR3joOEsjituXjJsWQX4QUtMriVj2ZJ6vIc07R4FBhTiTwLC2Hqh7/6zwu
O/595y7GV1tL7tZ+1HjLD3OkLLm7onGHA+7ghjMseBLt1ar/1riMTlWhyGrG2Ww5QzZsIfi3X0I+
V6gmOAtOmEEkPpFmlCLq+r2ySZXEdLoyiuPA0ar2rzyhIExroVCzwL6nRNdPnCFha8W8qDhWLptF
vK514Ita1XHPDd9sAaJMgSVvWQO4+VZuJXIMTiVEyQ1JckVjyO5Bci2ioonq3LMxqnCbVAygQ1yc
B2LU8XFxsI8sylnOGPRMetUg77KQPZJtw85tvonsipwDffvYjiOiNkhhjoTDtuNOAUERU5zdmKCi
R5QY0BVrXyigbe2JR86AmByM4c7Fa1CSSCcvjcbfXNduiYqBuImxeBVETNdR/LTDxbX+m5+CM7U6
uPVn29YyiKwzlg3ixlSUIvmUxXTC2CcE1qq2zcxczOmDnzN0UAwj0BU17ORLtiQz+go7GtW5Hamo
RZubg7i1vgu9qLqsMsY6Sn3Sy1mLQea2hWcUxb3L6reEYbwur1kgbvbhDiJT/vAe8moE1ryXYt2g
Mb7qSWnwSlDbaYyPsiSLPjA0p2E/YiCyUK07VwfaPU/ZTuX/GH0GlMwZ8EI9VugliIC4N/pSxGj1
M0oeCbc2j0PhFr+sieATW18ubz0TTbpMtb5kFU06YGx/fKglcUbOW6H5NkBZuFuXhRAYq6YwcwpF
F9xZr93pikJTbqrpN33ji4aYPEJ8us0cQDXuNVLK21x1afid4hBRLi8/uU3PeRyK9rFaLgO0htRp
UK1Z6nsxuCnL4zKaomm4U15HUlsHaVvIunovzRxtkgZHDFTB+CQeDN02ey8qKcGsa3DfUMxeXhy4
Fzm/Nrul15GL96lYUakm+cbD8G6vSO205+ogVryxRsNc1VcwWxeq8U8lu25oz7PcmBa094vkwHDY
hzAI9TVzk3iM7/yjXn9zGK37wV+ow261v2xO5t/FH9qp916Spoev3t6FsBHlEO3fTyWCUm8lpW/G
fHbgA3vQJvpHYqcKiB2y0onw937di3/grmjIIefyoh/R3Jmwnmn/sYbtXXWwUlumUOYJ1WwoEaBk
5UOi/TvgzLiLvOZtuMY31dmrJbfmszfZlA1sW3f9d+zZQp7EIC8StHkiNPr6YYjeHjujyvEGpT8c
Nd3hwprOawucfaNcgH7sswGPs4yGakgz8W1mFDL0rUfq3l839j5dtv/cXMxuQKG0hUFPFF8F6Dpv
JAI/JD25mGN5Heww19sLsnk1aDsYKJHMcE6JAgCoua/wBoHKmnRxRgT/ciAEdihRF5M9fYfHsZB2
JuZnLa55NVF59lJzBWkzcimYiD/Rj6TvcRXmSqMMyzNLNUoA5gg1eT8Z+4MSM+eUt9M76kyUM1ZG
l11ZuptE/VB8aJ7vwa1m3D9UlXnvO5jNbEqhgZldMMWamKOOY7Z13TPkNS97TtCC2zykHyCeIEK+
ngyOLqrbgbCXvrRQ2+oTQT3apCOgTqb6vBtAD3T5u72+FKFSXd0g2qhFdI6vLMaCFq/2qBED6Fpt
ok4c8xjvD/nKmeBPlk5NMtWFtY/e2AHwGzFh05oB85XTwZQOSfJz8umi+wAGb4QIJORrrra1Ebvc
l/4KwrxM+FdGq2vnot7f/qCmF2/yKxXy3XsoXsIii8poVRwSp3o/WtgH6+mAvgrxq8d6LF7Mkk/N
uU97eGo08MtW62Z5yCtBUjGvGwseFYzpvvqeyTEu6CmNn3cmEluWkokSiqnNU/f4ArQDYMvv0kow
H4zn5SfBeu0urytz7C8F2jpS2IY83kj8rOQ2GRULpWlZHcZi9tp3JBkAhTVr3vxFcaWeBvsCt/2o
ZOQE9SPN3IHrRvsbV2mm+synKtvWGKYvjS7DNuEqrj84H/KX8mE+Ja6nI8J0eBCSMBPCf/I9vXbH
pRn0SilDdugCqEzC2+JKZElfaEScejrgrz+OskEIJeyg+0eiKftS4qYl6Jw8Oneg/11ztruBaexw
VfKaEtA1SvDkjUsi3CgA5qY+hvI7p8RmUVCSfj+CsoL56gs6sAglKwVFBFO3ohMcUoK49XW+0/r1
lmn6X7oG9kuh1MO0NaAptowvHm/xH42tR+Opobi/hU0myV86XELoGrV86gk1nOXxZhMmOFkEi/xo
BOkfcVyMUd4fA6ihNhD+i6ZUiYOF3nEbNBz2GBy7ORDBDueQObA2Ks4yiWMBh1M2UhgxDlQwzT5V
VSZTcUMMRGQ7DcMyqFlQDawDAm4lsfTVlFQvlt6Hfs9cmEhvrBvu9Qzo8Jyff3HfiD660oWMthup
74BoyA6ouIq0rEnU9N3g9QQnU+76Maej1SvAhNOph9jYlLhR+Xq9H+QHnGu6a3thsK5GI65Hg2Qs
0ZBNy+AoixpSPjBwtJUkuUdEJkVLtS81BA8T6CrGMojYi3/UWQ57wKS8gtpx/cVvJ0usYC/9UMkH
GRjZ4wCdxG4x/tvGyWNsFuXST8GRfyfMsPaM6CY4gGPNEeI5iHkxbesddw1dRr7yp686KFIEjbhh
VoB2sQFtW3owkc+pp6/6pg9TZvWsYXfZNgEyJPpwlXm/sIvZ8mIabQ4XoDBgbBOXsyvgjeFPwgpF
q94tDO7LOUZtDRQPxEzzOis7AdVC5o/1r4dulVP2pHOvn7UdYTmyRan63dG8Ya6LWj4xaa3YpGFo
w4a2NcmnDz49IOlGSrxRY1Ml15kTudwQaVdwkNho62Mj87dDzguhn9YqKO9xUI6qsl68t1hEfHbb
+WQYq58DbWtcT3Vtxd13R6cNrAmEPcbZtuA+vxa+4KVTovLJw76LNgq30zvLZFxyUz0iNgu0RNRo
T3acLgFQ0oyAm8xKGzd4Qhq8ftP+SPFQljNc0RmZ50vI7Ygz0FF1d3TRCX7XvBmSIiedI5PIquri
EdItyX5RKYRQwa3StbY23WvItH7SOv6BkmVTrnfsVP1tqG+uv8BxYDVO2e2kUEEavYxRxmDcLS9F
aVlg9i5wey68uiuTX6RQvbUNM2TYYMR31SzeEEBwcPdmq6+juLHLyJZ4UwOL5Ul4xt9DJqr4bhhC
aG/n3mOoo+26/8em+5XkPr1iqiCDB0X8i6gcv4GV3NJTdYTYIGEzVdTkfQfaDBjNrmWKarzaSr3I
ZoZpnzmUAp1wCaxkSuFM+AC55Y0SyEAU25xsb1NWSqE3LF6aiN/5AQtfhDp+vtOMurNMwmQgh1ht
sJXzktrd1nMhMFclGdCn9smkzCqEw+BOa0osFc3N5UFFaUbzbvp2/9DrEFl/AFaW6Cv+vAvhIpjO
vtDEsIRoGLTExGugGkRQHHqqh+Fbco/O10wpdqDQLByY5RcDWt336YYigdGhoLScbGtfpFdiu3V8
7K1xbXnqdgP3lhb0SziGvK+fCdRzem7Qzq7/CV+Uvu9DWasTYgKsawEBf2siNpEZKFY8i9oLkfIg
MoxWSzV4v8NL4HRur+2cswLFrfMPXdFsXCnDHNNKfwGeOz36fM73b/2CsVNZf+M4ORWvHzStCMqH
o9STEhWznHMpeK5vMP5kz+g2pGGAB0f/ajyRxcQbqBLJaBhNiVEehKGGPtdP9iI0LSywufFgQ4Fi
sIg+B9gRA5XYy1lyWnFObWH6105z2JnYviOrmVUihiJkLhEcr5MgimcbtM7mucaifOEgvcpSoZii
i4Ztyi3+x4KmFiMje6QoAWvz+w0zO0xdbeTNYLa43x0/7jClNpdv1tacitK7INLnz1/xVVF5sTVt
YhOHOcWYZWfoujXPpbgjAENmQZs7ZfnYX7RkAZj+xAji7MkbkncZSyzpeU0eXmgU7wQnmxjfn2/N
WolBWvA6iexqWGRnE7Cn9K66LbsZw/vMEZiOVwFVBcopX0N3Bw6taEXNetyL8wWrZBv6oNzmL7Bz
1qf6Rz8vgogh/Hk676mVVKtPSQBUL9ea24G/EaUn4q6aiN4h8CD+wzsxPidji51u0JHSu2lf8k1g
gV+LLFHCxYMxrMH+L7ZzRxwUztnvmh6VpVNqHKDdHj4wZNqi0iYLAHiX4639ChTSodY5A93kgPEb
FWdjP6F6P12NYYbuOCHPyTq6VvBInnE/d/1MeSwy1V6b7QJ9UmAg9v2YOHLifCVJ2r9IELfoFpy2
y+Dh3tI0OaUUFr3pthTOHDU1uoy6ooGHYs2zRVJrU8Y4mqAY3VhoQSIXQNC09iO9Vu2SDoWGVc9U
1CN48z6DOHqcPNXanX1yiXUW/IVIWCoP2uiq3OzL79yBjQZhT74zkGa9dV5OPSsmr5kyc4qVJGAi
3y8gwDCy9HxIqjbIlN3RjVBRtNN2sJx3uDT9K34cE14Eqr0NBUUdBnQRbYi1ZtmnXCSAy9zFxnkI
e/pZAYSlkgH3GH1Ty+zPp/5ILBMTislAIVHFX/OJ4K42J42hn8wQJ/BsJs58rdTqW3F+xk4K5pAn
3LCXe7QT7MECwUapMQKkqyqipfTN0e8DCpLxfUmonbasll5+Snew/aTN32f674Xtmmq66w/+Kq9W
zka5UiuXlZNU6UXC8msvuSBj+ih9Of0/EjXsJu+mPDOzDWq9ZNdzgXfQswUrQyMFhw/H6+mskm/s
Wnvo0rwDkicUkEJy8dRzIvhbo17r7VTAcdvO6EP8MMajgKHo4r4LUx9UpqzlUhMem0DRWLDaTl00
foeKcHnkCQe2QP9NKwYSrG9wBGqytAwZUHrGOaRVCe7mweeYNlXZYe378fcKRcin3jNUMIbrJKbQ
2Z9mcYrva8vdnIUWN3rHHYqXN4Y5wbpFs0RrzdRjijhyNUB2ppG0iOeDQvDZJL7e6dhnHr8G/pMh
iwo7JKIoGRwg1GWQBHdmf9VazZnhH9/ZlWq5u8OTH7CIqulyuD/TLAoKcDbp9AWTv8pF74Zdu1ej
evvgYloUEP1Ah63nVTR88p1Mammv83Npx3GbhLRTAeK9z/+nHRHiTPs7umr0mNRommdzoN6QWLLf
E6rlHiO4ZFUcCyp3kw94e0mswnQ4VgVs2LUE6lxCBfArxCW6w8AG84aHH9tFxK15TONgH7wm/FZl
NXVKFuvr9bARSbGR+o/evJR6XMzBr9CNbUepkl5NGlADcAC5x7vD7eaN2HMWDm2Sp1yeJpYtgjUc
HVWglf0ZNAbDeV2kI/W5Al/sjh7rmYVxSIuR8gjeuL25FGVHMRi3PMsSTAbFU5egRj/NN+O7PlHw
NIiIv40HB41UWt7fMYGaLyPuEsH2k7pV6vC/ZOefp6yBfZQq3+ry4/60Inr/jxe309eR9r1U7Y8N
/HJ2mJjU2un4fDOSjMogJHjkq8cmKY16aOgOCvMKXq48GuoxGQEfX6Ku74siDuuc+iEt+TSQbh9a
e+LUEu+OxtySfp24MqDgYCCF+GjtTeYFLhYd2asx/toYXffRZgjmilbxPabiK2g7dWtlumz62giu
aDj30j7LLPVPBgfMtekTqV5E3vyfRKlZdq7q/HYVkrS9oaBS1rXk2Pd8omEUqc032Tm/g2W3m8ji
iw2FzDLVuA9HeUPkgGkzx2hYHTHQ3Eckg2+ShFLDmVIwymn9Jz+Sd5z+cP227xQhj6Tb0mEhw3nT
b9HVgPo/rxkPgThyxXJn5Vzxl8g4E5xop9K5ZrjhCkLJUKu/6bGZgFaxYFg5bcMQkUfBsx/zdzy/
G4PI4X/qX8rPsCm1ECvM7ASaMPA1ky/R1oKNOtH0SH6biiYlxSkHFFmvnJXv0ynSkClf2nM7ItyL
nvq35GgZzMSB6GFiMtBeLp9JfkFjrZkUIVpHWyQ22nrsKXq/EQf1HgeQ0PwoklueXvNrZby8vNXu
SfTty6WkwTf6fGnu9/iCkksQW55jS5DB6zCwE+W02FA/Lqufr9IeXM6QaZ+hoiKIVm3iTCjGsuxE
E0stRj6pZD13z7vDu9EvI++oLv9klqX3R1lH3ZxRnr7TxlEequ6YNKYBKc8EtjyjfQnriidONjY8
Em3Xf1TGq0djLkM+aImK/PE7u3Mz9iAwgHhzhH2HhVe23h17OSX9JIXKGBpDe3RxwNR4L+iPf8xi
E5mOh06NQcsiVOu/0UDZX6PLbEfH7SjspyKLzaeETTjm6p9QWE/ZY7/dWBABBNEznb06igMSTVPV
fNYNx3VPTRIFhHcsccsEyox0sweNvAwfMzq6kOOiDv3t64XARbUZLh3c8uVC7Z6nikGeYYGt4Ic+
TdiEL1khf1eVfu42f9LW3D1LXtYbU+VjhH27rWkWAI1XOgdzLwFVvdP7tqxr7tHYIbWbkNaB/n1p
VTVs+RG46kDr6O0dYXXcQMJtIvjkdaqCOO0+xhT3mnvbn4Zo7yjThjsiR0NZx83QncPZDhaXHg02
PFfHJA21CxNGoJj5PfDuiNXZ5XWQqVmgr9fGJQ87mzxqgopa6Jq/UFpQ3mfHaTaV/I3IHprii5kX
Z9fD7lUyGDVOVjo7Giht1igFjXI9SJ0zM7jL8qakV+95olXtsaAfC+fFGiVhUySLfA8CQb7P7k4R
8HOtyx3HI758b5uSzM0zGeNKIJg+Onhc5edIPZaW52z1pRCAtESNonhUWyqOhzUm2IaDjxkR81Us
XuEmibk6844hYkGEVQxiY2tgf1AehBCfplhpRfE8+44ssfWw9E6dsOuQGx45FtS4uVipWSTI7glL
f6egL7P8jL00o6osDU67jma46u/9R9GXfCcVywZlvunLm0Rg50OpqtuTNy+3XYUk4tS84A22LW4f
a1h3zFV7Ppc+Dp486FFg1fmJjz0Ka8dwvTcC8g6IKAs0Tak3Nh5Oc4uhI+1z9a/WLSzceQODuFt4
90fcEW9vVnb6QuY5uOiyD1X+yKnyGgAD31iMkDv79bCjUl9QjqEWQc0kj0oHEnwTSKK6DXfC70di
A7iYhZ1t8Vyh/mx4U7J1SZ01AaZzBnXMe9E7TFtrFapehbqypd7rzyJQrEIF2rEGj+AoHDr7XQtF
78OJr+n046B5jhdz0H+tKKKmezb+U7IHMm7cZJPwRX4iyhsb1eEmCvOKm6yDGN2ECbIV7ALJqN1O
yWCcwc4t7+7zBfaQXF87SwC0IherMlpaSfozjdL1cNIhh+rnmR+PkBG/K9951H1ihW8l2B9xo1QN
dODBmw1lS0RjteGCcLzuis2wx78xVHOEj9QUL6XDRaKFzDLXeLCjBOcUTR514haGR43iCvL2/pjU
qioH9+q5sOdqFvpkFhH2t/jtenh2vXPeFw9W78C8twRHIA8O5Gte2S3Z85KjzJGq8rS8A/vQv18n
/09ED932cV/kpBLZFIrjnG+0mhOeD0DDkZqR5+uJw7596coSt4y8EIhUPafAzMEj2VFE0V3WUnH0
iugXfEuebEqgCjoTVKRBjubCdXojVCh4SHjAT48k6HoK2JsN0DpPQ2MQt8f8LHfVtEGvFQ8X1PXG
MESl0TgbRYOnO17M/k/J2DjhicugYS8CKcpMfjZSMJT3TJ8VAXpVqDHgOVZouq3VwwrUvJkDLkfh
hiqYMLgpTFVwyBo7Jn8yP637Qe+7o9h9N3T9AEbVg6GtCarKjd4G8bK+nFEhG43YoYshYFCEstHj
aXEIIVFV9+Ni6zXLAPR3M+AroG/nU4t+i7CSz29YDnbbn1+Z7/U1a7/4IqW7bqIDdPyf/eueem1k
vdP0WiNi4t53B+nvYaQASzIUpBxfCtw5QYVwxpieBNbmQuXm6PxJPpDm5nngHp/UDMwsP4iqal/Y
9L1kAiaO7UIKwQmUOWd7e9QV3sN2C+aKo9SV5yUjBTFuKhIGDhV+i8FsNJYON3rhreAuTxc9fpFP
8bV6RItiADe6qT6cmxR5b1oTCIB819BgaavSxFEG8ni3cuFrDoAj0IVreqW/amYcyx3tgcBnvzKZ
9ppGCgazCWHjtnsMbfyCCh0TZpzVZoOtx2s0XWuxJrPewG+p0b2GkhuVYW9vrVIFvhnjiyT8O+Aa
84Z52Sf0JfUE/yE2TyAQVykxwcCZ8Rwd+XwRa2Cr0JYE2S60r/cOHKClVWgQ4bAWfCzwuJnWySWz
5cTFcz7GCqSbTuW2cnHosnBozpK2ak3HD28dNkpBPwzrn7meL01rmirEncYr7Qv45GtHDf7jw2wB
G0BvCBBzZ9A7Mo0seT9SnEgW+FdD10Tp0psBnbRbKranEQ5cASAP2DuMntE8h8d4OyFEjR7V5c3s
UpYgzoMxyv9TKS66N9H5OQPkOYF+8FKqLq+qRo/Oqfea37NvxKN1Ed3sYAbRjkRh1TFzC7zOayiM
KBKBcx6WVgURFRpzEd+DehLYGp7UhJ5e9dzfIasacTQlSNo8UxVO7yJsCB4K1wZRk/0DHvQozrul
q0JXVUdCv/JSSWgPKMwgsqWvkeEYvLqdCjvwkalAHCo6ZEA0rIDvrCGnjn6FDPhJ/+j3iFqgH3WI
TqhpKAANhO80uTerCPG11zzqpC1/qqj2ZZI9IQ2YDeV6iKH18w4QC5F0TPdhH4eGYTrMqh+UDaB3
Na8DNLI/yA2NXKHbeCUFsLxL7gXRRMYN2dNi8NdwnHFAn4AiAvdalptFnwABxVponODU5bfnUBOI
DKbFk7QajfNg5qyxQruqz28NKTONyZL1AN2UY/Ww/z2ZCFtMYdBKBCHzIBdnpukgeWgNYYxRCXAC
DaM1vGJ0eImIEXMYDBwf79/f7lWTdTQjVxfcBtQUA1tpmubZi376mataSnVf0hYJ0Xxbb9PgMRbp
RiFYSSyeAOXa6osfm6rtSW/Zq1MV3yrAq3drWYH3rYRzZwH0XQS8AliuhXyyOpne8PlcOLZDvkzD
CYzGEmwjYbSQaVs3xZy5sges+olbcP916fxR6T0YBUL4O102GOMWBPsjPI0f5l15QGqQ15FNj/Yy
P/PRW/RXN6kbvIxQ6Bmh0u4wNjOSqA3i+Fflhq/RoBNUXSiKQ2mZKkeVe+ZAyCEmMGpVo1YFS2oa
dhFwtTlRAnBUV5nIiu+/ZJTi1dbYokgLbtqSw2/l2G68hfIwYrELaCG9k8UZu4fCFLFv2CWA0vRI
yLird/zXmiYNpJDwuoDFBQesNVUqOPto7X3IraTCZMaYQm9bmSI0ysDE2lSchW+w4ACdbT/ZxDCO
x3Zzn70git5/0ACpEDdzs7/wyB0QwJO5HaHxlT4rljc0bnTtaRbeh1iJ8SCOmiwg2NyXqH6Eguw3
agWU4x0fkBKQVeg5fOO2XsYtL4CrXl2vPH67SpPAodbVrXQIoz8F36pwkxL3JfXEO59IvArockl1
x1CZQHGXhx5i+tPVsXneVfgOpmmdw8/aBhIOI+hKVkNyZ+db8hlgLRKR1TzTpsp2wdTC9655wd9/
H6QErSbrZ2vYVtJ/7V2olZx02xyzYYZDVPGygozxSEasjS0N/a+AyAQ5FcAzb/qh9OdQi1gM1R2K
VJDpuSfe298k0XZ+yRLHH4+N0Hif0b4Y+PchsyteNlmD9otlQdoGiNbnV7CrPRDfgNqZdbObkPSD
7U+of/e2r5Pq8tJD236EJbR7IxG9kn6i2NBKHNV2fWsowXci2AoWUPQhT7GoI1yTQ56XqWfCfFbs
mLLdAbMmjGB24jrWyc5e6ebmPxGwxmQ4zAmEg6ytH/u6UwRbcDJ82OXdFDqO6UDpxI/WZkUFAaTv
ln9LtuaoAB/gUPNPjL9drkjYHfeKZu61zQ7WvO+O48tZGq5kYZ60Ouu+BXKASW0ErN2opnWQ34aR
/TTMZHqSy58UoKyjjP0kfDA5QG1J5fYyNctVWyzfZoXIlsb5pvp47dvx1gZFShg7zpl38Ag02aex
r0nQYdwW12oW+zfpAGA6M2+i0Se+a7gW7QALQUrMxU+VvY7S/4yqh8RotGFezLjyZMMbPqdqw9OL
0SIoJyzC9V65PSrNGaXUK52W4MMbJlwf+gcDyHGuF78e1PuLt0Wf+FT6oKRFeuuu9XBeF4kVaQ2w
624qvKVVe7ccZRl53n4phgqiUXiJf4tODRb8g2zZ1FWoOruF7VYonQfAC1lYqJFwTAbttfyGBBlw
tjoZqOAL1iCVM7fY9aiQ4EuCFhc8XptNHk+T0LGFtHPv0LmPCC6AosaKjivs/rJaktsrrAN7YLid
Vde6Ab5Ua5ealUOVs//lvEMbZ8eVejf5MTGyVls1Kyopo9LYMcisj3U1vUQv0AufKYsWtBN5IHvT
CAgoxZGRcF0R+orAoIvGKRdSUjBp9euV+72uvYp6fTjBIPHSu2SHMRk28ft8LQp+M06mx/9HyMUo
L3YByNZph/cm/BBsz5KOMZ1FLgLwMEFgH8WPyt0f41GcLEkUhFjLjUAQRHfuUc0hoWD9EuxD5hAw
s6utMv5nkHkbbPXvQ/Cigy4bg4lh7hl2Wp29JpoTHbOTays4XraySF1rLwAn4p2Ix0kxRAUjf/Ua
fF9SnoK6cZ2X2725CU3kFGAlnYAlgPaTOpcq2ijILiRZdmMHyyKTfkgI54oXGMH1F1r5NyENYO4q
y7eLpykswNeLnr27Ic0LN+gWVCwaHBzVF2pvoemadzay+QRwRDVo6PdJEilr8qbloA/UEW5KeBbn
Rc9F+NUtRFidx8ytnIAqWcZxxQK7Qw4MZGMz2H2alw514dY0P7N7VUlD5EjAYRMZtWIMMWB55VWN
t+8MN9O0/FxFIayiKsQnf2ST7XPelYg9B17vY4JxpEGbjMzZFxdxiJARoUg8z2QPs2RZxNYU7/HV
s1g/+o/b0IhGIXpEkcTgLPYjJ9xlpusI4Zz13t5ony9f8JINbLKR5khOd866VVce5YRxVsjvkOfe
60RQAM5FgWyLa2YBvvfyvs1n/YCe2VSRdWKnZ1EvMM7ct9pIim8K0+7v9hxx+j6DZGQD+UTXRVKX
Ad14pr9VPxCWspYXEnSZky5PQiLReUYUrg6FZ36oXCTlw/v8ht2Fy3uG+44nrrAoIFtszNFPS+/k
TTI+iIDhy4x8wH40hQDMr6GgzZkFZ1AX2Ak7PK5nYmtrXINQJBGDejEipT5NmpqERLCZfdghz5eT
ZZ8yoyPP1/b7+yP/vuDCDSMfetEes6R5zcxDhsiqpU2jaI+WDKI5zntdntnhKDicDSUg9ng7p4DF
HCM8Wxml9Y7qATImyk8I5Dt8r3Lesp2njnr7HTXcrotWNZWOvpLYjluJxZ2oQRqDJYgCGprfkMXM
c0wTDb5qKL3TxnCydGu4aRHlhAfssY5iG+Vo/CwmT1hvS8K8ule7GeHhTWTexTF1XPdXoH31hoW9
MsXrL/K7QGWc4p9lLFFhcxppGl8S94YV/9Zb4GwIQTsSO3zS+86X4sUg12g8sNVO8wZSkPqa0Hrp
XH5Ff9fq9ukCnS8BPdF7YSYQ60EHCf1k4HcX2bHBMdg83pzeydIewMMVr0ENRN4tbzivl5hMusfA
mlVm51U6pE9IRJQcpkwYRuTe/feea3ZS8W92vNXLZfHK1M+UwQbOVkJ/+QHHpzNfmhKp9WgewjuA
W5JD3UVCEGdU9L+KmifbMcwdwk3hTnnvW+aXUOGVF4fTWFRQtWndviZptOcFDsC55RT+KJNHxzWu
dcFdOJxWzH8El5eeq4+wYCDbQ78YJCR2mfPaq8K6YP8vs6euQ9O5V+kCoTkofBm/SJTNZDcMRlXt
2DHGSv1SHupNuAU1C1qx0KNX/mlfJ9HyewUkKqT4UjGJgVhMb8uEecQnvmot0781Ppvd9b9h0ciM
t3A/xKHAJMfB5ZiIuA4SLfGuxUs23EtNFvMLhuFP9Kmap0rczk86hQ+DJbLXUzRWYMQ01cCzFWnN
Fc6TdHXzepjMeULz5/J0Pktxphn1AoFS1pHmfMfRnj+Q4bmxmN0/6ZMIpGx3yxc11ij634wBv5rt
AtOKDwJM+fkzGYQhTve6eDhsQmPae3McPuvkWW4q3BrJrSUz/NcBykhMzZZx9dS/XL6Fe6cCPA7R
g/hOnfc0sbplGRmLiIvFBSb+Ym/Exa+nIVODqzWPZlYOYmK9+Cxn7VPe0z7NK9eWH8vUjdYO+gXb
v+fK0+Sy+VoHIQkeIx/GJELO92vCWkyn6nyPKNcVYYHqxZdZWDlJRRrp1Wolf1I0zidykSWh6QSR
TTyYjjZ+t57PLc58WfXkj2oDB/HogyO7lHfSvUOQFQLhwRT6LIrWmxNzEBneRGR4bVjyWRbOTwoK
PmbAWdVQ267AlI6hwNrOc4Sd3fUuZGaKyzsRzk1GFTvO3WfXU7nO3OgS7dwB847SYyvA7ZbldSE3
0OAV4Fugn7tUCe7B2dTs3NpE5VE3jWOwGzKmAnH8i+2HRRxEWUY4m+r0S8iNHoU54ayTfWCcwxRL
HNQKbE/WuGn5z0JgAdvuMU3RoGm82IRhqZI+kFulycUZnDsBH6xWzjdhH5U8TGo0+jiaedHdEECZ
CyrgRASJDGKkPKL6UKtUtW83fYSIFOhBfaNLA7qp8DqVUSETbWUZ0uwuIW/vnJSZDVw6pAAU04Ey
6SwfVoQEtJq+r6lDmHZDC9rb2/3O4nkkgnI6Q9A9R/O/NwXenKTRAfNuGTxvn2M+x6vsKgXvj8/0
Ufs4OfvZEbP+hSqOmTLblm4k8UY1+nrh3lB/GfI4DREZBh5VnmybwNMFDkjb6YBtwgtDuaZHx6m7
1bPmXEB0G7LqPEsYqEF4Jmb/w/l60ccqfLfIbiZ1aqVAk38t5mUTavfXcztcwQODPYRLKjN5TYQ5
5s/1bzhTIsnEP7JynUgMQR7bl2Iydw1weAJvKm2oyT+Ap+LXeLr60/KKqDevmbtpcX2Tj7ACTXgw
mQpnWzN+nOjrrLl5ILZ3OzCymWiwbC+JRXfBslYl9R3qvx2zhAUOI3AAgpvlEIWjO4Zk4hSbCYK4
G1obHk84v97dZGcEHBC7ueq4rgR45N7rzvcNUDusEFeaOni/RGtqbv+9iTtvYFj9NcPKG9mcwV96
Erp8ULwOilUzM6aY/YiqKebQbRJaFdJ2WSWRHR36bEfplxmkQhYK/0xwHbenGSRVriMMJ9UNGlqZ
xczNT7I+LqOjBvHjZ8fkgF3AMr82BAzgm8QPismtCun6Vjc0X3wDi7l4bkol7UHo22lQgsfkEmqk
mIDDKDCLb86IylGGr5/E432WdEaBw3+Yks5cAVKx1VCJbJxZFsbArFnsifukPEnnYYsU40yPt9yd
aFN2e8pm4ruKGZHOdUX+IvP4W3cItr+giIhgYuSR/sRFVqzOQPte/XTBuPYPSDopQAC1Bm+PWnCL
VDxwMlnBL1zZKhavO4cMrbGMWn2LGLkx7rtAqjPiNRzkMYX7alP+Yzt19CdphZMQ/h8yVHWBr0yY
9PxHpKGG9jNGai0NTp9sN/USZhDrQ6V53jYlSPCgMEUMYAh6mhVjyR9ZReowAp0wLj2ethV6D5H/
o+aS74rO7go1D28dkfUeEOGmu57AQjsENMRDegi7VVnQZ8dxDZDhGVxFLB5rRcL6NaZiCjwI0sB+
dV3iBFwxkcqjXL4RbRWMCEh4jJ1IsBMS5QOsPaw+lVJiNC0feBRlyE2UiEhMeMYAGkom6vTVeQdC
GuMi/pUi2bIwOcQjRSJ2+QJj4PHz8aEEER5pqtP2yUCH9+n84nTLqnvKMONNR9W42vchVF/wQaaE
jRAk74NrkQH0xcP/Wy6Cr2p0TchjVdpTbz9zObXywtQkzcx5rm8sDIiZbGodbheDYDPGkIxaGdV0
hWsDg2bLJc9pLv5eeitAZeAUcysWGrOoXw2NnWVUbkI9+yGn7uuslXhH+KnOPCXwqySzTVPXzhiR
IAC4eFij/169S4pytZnF0wdrGcszcpBhfuILvsNPriP309man1Jp+6JIrTepWKicTg8sZqM/0fhO
jnv+mWzn9MRtWndMv664X3qPsFdC9vT49zkVudRbrHdDHmBP3mmu+YTuCL3Yndie1o6Uhll//j/e
SXSofRaIbbrwHWhfowVmnnB1y534rHVRy6R1EoAiOT8ofHg0YqcZnwPPfNsBjkdnIN341M3h4GCf
z6xd8RS4MHVEa0P830+ko3JL7oZOtZqpYMCbI/uoaK0tJ1tzURvBCjTN3WxeYTCpGHM0+eRt7ltG
nLGctYI6UqdWmwVRgxIoppOd2SrN5Pbega1n92QQ1SEDtVTCx32iaDXtZN/sKn31bEQIS3Q+dOQu
Ilfi6Xav5UTBP2+nLevRHmcIyGLTFW+dfKZp5T6VpIQG/nrvT5PqzNbXD5eaC+ehgxddkaIPUDfV
WQUlkd+ZFPIN3e7hLA6je4eMQTtA1Q900odtNJN0anUUAxE8O83bYlwXR5kEL5AAE1/d7oCso3m7
dShBUC1d7b9CQfPWMJwj2g0vTe4y0k1h+li175sxF6qUP/m/tN438Up4H8u+JFntPPYseeuT+H2N
Qs8lGCBsYRHL4n/oVikUuEmbf/x8VlSBAhFCbW3LuGNAb8FOG5icCiHeGMynLlRHMGr93iya046h
l1yGLPVmLy2l3HcjQteYS3almvPxUco7OBsFen6QWUPTkOGhDvP7L3gWgqDxOn72QbuuD8DJ4MaS
lEqx8MSTwFSxvQGQpnG9WguePMKRxpUD14k8v0XoNYm2r7yV1cJimo8JGSGQJ9uXjxUA49jl5FHQ
gr8vH5qrZHXoNY6Sx9W7c0uAB1PNDyR6H8Qg8OsWR0KTipain5JgXiHNIG6fSJNFiLwnPbwckq5j
1IHxUBJXXn6LRgX9uHMfQLLDh2SDudcOi6ajJE7ExUihgBLA6p6M36W+I8jTPefNGcyOv/GG14xt
CH4EfF7Xs+wuh/XAE2QjpXrvDCrS+eumf2ITfP6n3zsbbbIgtk15HbotRGOUYc0nsc8V9EhEbg6m
Xw8I0fPZziI1jZwfY06PqlWgHdYow8Z0sBxSV/BOz+Be1aXbYcMBI6NCaK+d4CG7eXklMXoR6OmS
RiAu2o7+kVVDs0M2BorGq0okDgWLouY7ytkm951pYyvhTORxIBEEAM63MLZUU+eV5bmouqEtx6On
vOnruNk+2TBQHM7IoGR5omXDOwQ1kdwtzv7/CddZsXhpwgYpLefdT/cuGaEGK14o0uH4o9751FFe
R+pB1SJH2osoH95qJBA16rE7wv3X+a1pn42CA9KqiZFD3U9GMoEBNyCtxy44nANZvQTJo5daNj4t
EwIGtprxp16CmL5sTtYxrhrgqYghxjds6yp9lYdTCaTsw/4JhAg1Sq4Qp+m3HaMT8HzKGzUPkrRW
mAiqYeyt1cqyyfjVtOA0AA5+6nS9E93tzLYtsqtqvEi55LXCkOgOg3HqBz6ovBgynFtkJnAB7Q/m
Cdv2NHBVhcc3HP0TF4aynhpVxwLOywq7CrE2sAo/fgGwRG/u0Y9qzCqOawBLSzkvhy8dfh83MuKD
8CpdQKcSLfOIJxF06tStvGYTt7y79zabo2Mq4xOOoUXa3oMHnkTXlxGlRe5Q77+WZktWB6ICOACx
E1ABYOdXbNydFzwl9fZBdijr9bnQhOFhnj49cel4SqpNWSSdtN9d7lFG6QUvimPVTXSfdoFAmLX+
zsTTWE57kh/g6FG7TzmLGTWwt1flIgOV4bq0xaJJQ2A2w+051beDZyVQTf06bRKzfjSQW0ouVMz5
4Hu2NlGircl0kTn0UTXej9qBQ5WdDpkkGmX1oQwPYMBmc8TSJ8iRHOYEmmayAXfJTqLeGD1ss51V
1QIhPuxtDxeqB/I66hPbXdTd/0U7JRlSGjeeUM81yHfGTYG6t3lSMtJmI9QLqNRHYUbqnNgLgZAw
GGw9P5KLuulK61ea1MmtST4r5bnouH7OKizgJ0EXUWQirCiD7aWbcjBknk7YJXSSSf94bHHSJ5Gb
iSU2VwAB0GMdOR6u1df0x8/7YPHhy8X7gmAyghGYkc1yNzv7hNFtqYd20vG8/4D4OeXO9hl4yQQL
syHxv5x7UnD+cDxA1OZvAO67PlfqF2h/CicdsEGkjcVhDlFj1PAcMqCgj+LS7etfYBGIdOQqRHdH
mCVZemISDUn38A4Y7ug8Cbh4vxYEg4Pk31qRroFtRtsIiuWDp5h/vw5O3ttE0ZiRqzuloeH9w8D2
BVmBEM1VW3HpYyrraGb0Ht+AOi7AykCBC73B9/+0uSQzNLQnXsI4MgzVKJaOCeOBIkMY0/CLtxuT
vpVkxd4cIeo+McLjOFFB/+FqyYr2hqZUpHE/BF/6B2KMLAt8SUNqQErYouX4rjh3FavqvY2BbfLF
5cpI/6hIqQrmRoNhHTb0PF/0gAvdN60SRUf5ycAJbHncU34rMxnCgPGk2yms/tujC8G58/+7AGWl
iA0UGFxlEaIrEqpa8CXl8hOnSf9eIt4EuJrXv0HT9FDH7yi8sEZOO9EtwMWwdIRW3ExMSikAFYS6
0zqk8o8FtXbuc8DGgGOMD0VkcZS4ldAgL3Ozu8ajQ8HlSX9wAo2P2beuZEG1XckUDPttynhsTI/c
5vnuZdtxYBKaMVccoTrEUMj3imNdZwLYq0xgeXj7Hpuxqvy7hvtu3oUi7XYCq4dJJEtzXxsoixwA
KXlRYjW/PZRXYpwUSaGdsCNTzKBdMIL8XfYdAc7FVEW/CIt9H2GYZXXx4tVCt6hq1Rd716K+TJKP
x1yvRdUwQBVVlTdWuF9L6o6l1/Nj270uKCc+8hmERdIY47kEd/EgSggB6tZn5UHTVZbtcIzH9V/Z
vr3PGKeVPtArMRY+k7sA3BOmCyhed6zLV0BhnBiUi9qrf9mrMzA8s7dTNEl3Sirq6z8I2DOaxH6A
jffOfZ/9aHyJwphEEx7KqyKhUbIw6shT4cD45ae/d8yKZQ0gInppVlUKRhG6wVtUxb8wmrbhvgAV
R7MsyCiLknf1Ymzjxo3ARNycGe3F/64COeJayYOgVOxEogvo7KjEwDBqycHf2JXQPLHqB/imiccA
UcgebjzXL8DK9jPwU8DJHX71ejHw6lxw8/R7F8mfA+Xp+GRE+if1GjPOye4Bo5/vk0ICyjst6A8Q
wGVSkOONT9w4HM1dvCOzZ+LYqZhRK7W78AjoohOK3cC4rQihyiuKxDWJP5UEx8faRaEu3fCMN/XV
yrDd46dBzIKONvbRhZ94PbfY7WvGD3HS/sAKGDbzOBBVx4THNZfHPH41ZpYJm9uikja4rOgi7KoG
smQ+pnMB9qNjJ33OvYKXMAXApawkUGiup6mkzjqfBqgXE/nmK0lPreM3fePXJ1x57w2lhgCNwjIo
XamsQBVfMJg5qwj83R3oh0t4lUO2DAuhYc1fNz5DVZyJh7pjYkHyqmQSR7s7a/yTic9uCCs5iBMG
HKXkaYHrVEzU4FGlyG+/nhLH4ajnUWOSz48X2dLdUFAp/iyq7hsU+S/8APwIIxizhp+cF9bQI3yj
NpvF8nVKNbQ1JOIQEpIjXPJFVkTSaDQmr3T5lcrOwnIWHBPvwn49rxrViK9MB329FNaZB929UuXv
36XULhxQVNEnqN3fbHJD2OSzvA1wbAbL7FzabiCfUj6aMT8Mei/ZsQp1VADC0QIM3TNl/f3C0Jbw
+CosqssDq3RxSidiu/a4bCAZNsXO63iU0JagQNqDmHg70UVvdWFfMnfmNURchJVss8rBtKqSd6Ce
ulEzVDIfqqJveLJzW/MvHpXM98b+UEVSLdPmeAHQKRT9rpntJAityEuIT2+KmbuvqBa5dPncPEzj
H/LldX1ll5yuEaA3BvoEw7TS2xTVRbLLO2cLQiKDrcRUITUuPLukJ44RtX2XNvoBwj+6XyrDCrho
WE6wZszlDXF8z1rK0Mp7ugDovDGhk1IsRrjlZCj8AU0i5ZQXoxqKC4jmElKEFNdGhIwgfeuvCPes
TRiz2cFM6rRrIFURUpOdeIp97RbsHacxfo3LKD4pYxWMMuzTbI1Thm6mU+KjwjfQwIiSQOcxYc9I
Y2t1vFjeQJqrEAQrVRhg+rkrmzjIZMy+E3aT75KpQQM3qlNiQLBJPzS0yz+hc75oWBBQ1BBE9QeG
SYFdJQcJHQKsj8zXX3DjJb4Pupc9gOSwEJCe/oTv/MNRiImm3zIAykHBUp0WTCQ9mr2Lo6tQTFgE
HrWvMXWHgDXdw/oNMPmIO6TaJ0MZ7qNk3K3gsiNX+uouPwKIQitUXBlL+DG/sCYcpQdHV3gYgQRt
z3p2FMhxog+T/9EUEQhWet+atRXrCQHrRSzEHkSFAHpgw9+T3NIscAw6ioWj0exQxz4QPjWhMtot
JXEqC8hpc+JhGGFgmp2Bm+XwdA3hEtyrc3OzkiZvKyNBB17FtdJbzzKoncFxTxjVGE5oGCH8VNjg
J4vs/dSScZVa5r+GKbkNBmdoF/dSrA4fMPSf3jj1Xl2ZUjQVbFSeG2qva5erPjfnU4T7WZeB49lg
0LqpZlxTZAmHFGD0DhFwYUKW9tf19NvpvrKofqms2wLpYe5Q+lnfo0PhyVnbEeq++zBCHW5gu6ko
J0XfCTYha0jWI3RacLVLkaskWbvU5Fd6ATgIqd7uY8gkqMQfsqwpzpgZvYyp0tyJlPGUHCu/qERk
JD84Fulut7tVvar5DCHsuyZPz0xuLrcf9BA9fCMZi/LdAvoUe/JVwDBVBkQJ9DR1itV5K2NhKDAG
hGpshoycMdMu45rp5d81tQt8uevy6RNTFVXJqQMX3U8Vhuay9+KoM/W9NHRfTUcKmrUiEi5ceRci
noqHX4oPWbJgZ97juthbrA9be+W4BuxzYDbCN+YL6Wc2weVOrI6HRj996BeIqtqHkonspX8VxQWm
X/vlSm1qY1hDsqM+L9Rz5FSirpGGLBe/RXHKAFz1sn1ApUGWdGTrDHFJi1y2Ed2D7rXXWehDCGcM
WOYB9sgvkLjpb9f86WVtiNPU3jQ5ZOukNTzfKqFMlxsy+yobCpJc1v381rnGCEUC3AokvTvD+NVw
RoneG15oRL94Q2YVC9FsWpFBw/q0jpsQ4RtZpw8a2jRAeB0V4sqEBkkxoXmlxnvDWpcfH0d2gcFw
8SihvHSenjbyEEQMt0Gg7RtBpb9hgMa6uOeOKE7Ww9EqIbYztrQxxTxxzMboCV53xKRztzDVfT4N
4ysxnNzTrclRj4GKy7HZKoYLv9Umd7sUD7XpekcvGmVUmURzJAowzG7PJwvsYxzHuMG3VeUgQtNt
NK8Pxp5DZpWn7vSnExBpE6H0GnJfPE8aLRKIS4ChXqXRFIDgQo3baBi7vh50QRpn17VoT3Fu3gV0
fhfw1VUuk3g7lds4E1FdsgLY//DbGV5smXk+EX0Bg58xLycCNqGcPiRaqGJPMLW5guAkrKnb+o0v
HYl/QjltHwgzrsBG/uj7MV7tsPJgO/LamJPA1LVeQmh4sy/5PifPY6laYGNBUUnyIvOBGh5TyAdO
nlAuoS5Ph6IMXEx9fzTx7z+O88S6a4fV8pIoqYT0Wr1JiEDg/hqGm6xpDO7SYbrAaUvifrK98LdK
i6qltfD1o5/SAOMozJucrlBtGJSyA/VuzCcbR7OwNZ1+8lyo41n1GSCgp4M5r48gF0u/eb9cm2nu
4fFf7zKWpPyUWuOKrIJD5fwrM4SXzGMOlCAZuBhLx/j6tsR81gymQw4wm26W59UjY0rHIReqqAUW
SZ8A++FLcp1539dYwqqQcwxW6uzJ2z4rgC7NYSZRrlubKB+gnvkA3C9T93spJi+8mv3olAJe1m88
bAyMc1PGLpop9Vupypi7QJQdKt3lJ6z2NkR9ih0sjKwvBywra1YqrMRY1oON6FpxcknOOM2RVNs3
4/11+Co9lH22+0DiPS/PFgCMf8yeBp19rxB9QgthL6UZzYbz/WIEPWR5+0okOZzLh8jSyiT5VfES
OodMRzV2A95UJRcRPWAeLnhzAdOAs5bwj+cMm0VGp/Kde7pITtvCtKNM1uoT8VL6582EfLm41DJE
+mxLfgLDrGhoXnpbiz2G3iH5pVXX69sMi8H9gny0IiCCedxyTFm33kHpOxMVbsGEFbeZaUCBaQfj
JkMR5cxZJbq4SVXZeiQPx6Aj9jg7cvzg2PMsXOx3W/u1aUYtsw9AXQVGbVVZCoN/I12pVSBMVo1E
JAOl2LsBzHPd7wC9jO+nfr/OGg+Eiy/94/s2mVjCLvQr5SRoQsrBgT12ZF52IgXEuieBcW5Yxazm
enq7Q7elfXDuyTj2VHGvURKsOUifxQkaTEND/icoAIBIh6E5I+0PDGCObtNb0GCoQlbk5N8EuMNA
q8KEnt4i6BOyNTk4ZKKyvvpaTlxo/o8TuaSDC1NcUB4T78m4anU+VV/4WeteLzUVWqpWFJzUGjMD
lpwXd0MRntPbFsszTwap/+VfN8RaOIJwQCvu0PErYq88itMqTWc8+/G0sRIMUx6Yd9FwrHQN3393
trXW3jhkUilf3TQHKO27Q4r1LctDJjAm8LUDZf2NBka5wzm0rUe/zxSlLNXkMaiEtjMc4BrTEjjA
ugiuCH3wIwP9TNbo9TLChvqfI0IDwRN1mONeC1gwoe4CAwjnRihpx4wmcORuUg6+SfMbD5U8qvrT
qCCbgsUx9XfTKhA9oYUTA6SiN+GLJgRx4ycfx9weOwiqohZNxDhssj11ExCxHtLY8e58UN9BT6Ji
O8QQK+5lozyDGNVUaYYHRjPvcYvmaILIfYP0OHrlsyJE33ZdX7+6/OxA3fTlbeIE3BJMubjZ94MA
2AmVelMOP5iGKeGE/0lpN7A3lFJ7xJymxXj7wCoUo9b2qa79F9dN+wd5WLETCwUmZpRsDD3agor5
bgJkBxAEuN96kT+saG+DNbAS1+wTgHXfWhYhQf/bzZWzltog1YvS2lK7IRu1Ik4WC0jmO7vNeR6N
IXvjsOycbj1ecGs52Lbz0ucBQ2NR2tczdfO+jBURcI2VPNa+OtJucZzE51kl/VDd08FdhD5Baqbh
E5KyvUlpP3Zxc2TQEqK/4c/ThU6+DCPFZsxspm+nU5XsNAsquJMGUga1Q9l3DuG8peTBC35QznxD
UT3TL9qmKoglokr/qr38aWWRfJOzs2UzASE+Xzc1blrg5gt1ZkFEcTTVxGjzYUv9lCjb+HJQYs8x
X3eioKHmtF/vMfWApgPDQ0HMtTGcdJtcoJaRpqrWKXQS2HoBsqyfQWKtZvA4nNLXmW1jxdlQ6l/b
uRwUi6XvHkz1qn6jY8shgMD8GJ/UEzqH6M6HyvjN8S3+9CwVQuIfn4Mt39qd/Ge8iROUDTT0bG50
vXN/IW99AyaYjRdXbrxC939CfZR2YO1xBTW2XSvvXvUnUMofaPK8U+sGM7lPa2xIiG0Ot23ovXbQ
nq/PraygOoCDkOiWdxtniXvd9LsivfX6NRFz40c4TA0Mobd7RXJOxn23ebS8505vl2yNZkiIl8k6
55RsxAYUu0lH3MFz/iR5ej4/PwNpc+McM5eyFwEn3HI7zjkUJZwod0lEWmJ2EsO5/pMt3zUamVmk
T9chmXa3yWUsPlvyNd60670+Eyvzinz6C7Wrgq42e8wV90VtBjiDFLphNSwznJVKHiyPp2YZ9wBK
z9jYrxVTxPdG8n6eWqSxP8ilY00tEp05Wan/sP+IWY6Ji2UtrSjnl/4p+TT2a3jgYxLc7cA+kTo+
UrZLLmpjOGmM2jBmeKNi116xrVaynQdDdGYJInICNK/w+UT10TDTZM4X/whdwI6x4J+6C0j0T0C4
344YTJL2mTM1WfPNrkgErrFBoAMfzCYdmvAuwZ7VLDxaTG0fbbjwGQE2c6aV/b610DZ4KhjBssnN
GSXF3jgRv73C1/kA3vlFKTsBz7ZpR6FgbzS/9nT3oGd9foJll0G7tr162bzIjzH73uSFlBEohZN7
KY+bGYCFiZC2AvETip9VTfsldcLcfK7Pwaif0m5AkgPi3pPocsd9xgwTZDsJ2TBfUTQMOVOFX1Jk
RZQsSh5jmDtdum4j+So1pk5XR6iymkyaWW3G7i4FhGb/oXqikcSFwvIemu2vXGpXBsKxDwzOwaHP
lsCfxkjDd+uwRVsmzJSHZOLR2blDmtUee1Vj+eV4abnyTu4LBkJFrqdmRNP8nffcvPdBKXDoKLIq
2NMIW3G3ixbCEL2x4ZBni5t9EwS7C8MtW97LqoHF7wuQjb56YBrj9a+OkCTrWXJaAany0ilNxJb8
v5BrR5LjCVi5+y3po4yb4HoPxzzF1Eqm+qEeFoc7UTpxHNMh5YHxoOueXYfnu+QpDU40iweul8Uk
asbwibU3O59BKgz7P70/cAEpbs6ABZ3G7qBggXLcVsiPKkjPrxoXBmi1ITDJThrdvGdF6pZpg4Ww
xPBlj/knOrORG11EJam/muojBsDzvYOES2oXgvo4r8M8oZ3B6rwqSxyJzStlzoQGgROuZKGR+zeI
GQKtqc0RtlsJJeazudKWWWLm90mj5cb/H+fC927RYz14jreDwztr1P6+Nv9AuqjITm0crjiVOH0e
bGFXE/DSi3KPZiQ1oQTl+mwrRQD+7LwS4H3KtTwIZpgn59zX+el4sX4ikXtKmMfiSCl0sC53AdYD
aFwTp2W/qBV12EgbZLVSXYVDW9qZ28ES+XwOEjNMl7obFd7AzfvylWVbd9rRoDHLdr4oDj1IH1nE
HFHW+A6ZtobthWEG2Pxp5XOlUCdumvN7rxjBrZ02tx/oSih5YQpJ0zdzAv8MCAw/fj4dLhEpK5jw
7xe4fe84pg8KywfHpJwStNhVvNbTqjt5LO5g44IdqvTzrz+j/oYg/us7L9QOOIgOVu2p98qDDCAt
9jt9gD0nXdDFljoYVjYpp8cuNmMPAi4DMNoumV5tNE7qmL6PpCwrI6JHWWfCjxl2S20NV3Y891i3
013MJg3HEXrl63c8a/jWZwsWi+dbnokCwyETHO8m6BhyoeNdrkfR+O4tnW7OAP1FZnTrDpCYhmjf
v8grsN5H0L5K04T4t7d8y3hO/HMxLFjba0t5tXCzROMXmXTFNosbQutXH85Z5Q9obiMHrD2OQPvZ
XIr7tgJmuxzPHLkswArzITROChWJWMciyirbhYRb9TleqJJK1T72eYz1ibpaX4BtZXYWoiZ/aXXX
fH2E67zmYzmtTANrTCuTeT+Thx6sFmyNOJyvNdq6j17iCHNCdITH6eRsnhSJNuRQ6t86igG+K0ZG
FLvBu8phqTUPeYAyRDgTKYmfZ5CfK0KkNJ1/Ne6Wm7d0UgsI6RV8sptyZRPDmPbhJhdrSexS1iWw
4oajz5plrVtaCjgGxN3V0ATfW3+BrcGRt1z72BloaxswOkHSnqQ4ZrReMtre1saEDaVc55ls/1Vq
TmGFeqmnzNdQzf+RbayOljC/RrYTfl/Xfh5bq99hagZaEN3enqIUAYOwePu2ID72vlg7C7sx6CUn
fjtWzPID6Q/Smn9dqkLmNGbSXrX2bmhCz8FtO9z9uz3c8GiXdNeyeGqvMoyhIjTR6561Lun4PGoi
Ee0vhGjZRU7LOJwTGgqcvjvWUBneK+nXtPT1og0sZ4xdYdCtIjK9XnVL16hMe7IkOiuR4l3I6Zir
w847ApXfiPvDmrrmdD9RzIbt2Lqwy1XI/AOpMM3TPcFRVOlD6wQj2XafkWRYYC0LW/xfOLKWnZHy
2+IlG1z9CJZtmLonH7hNaNHIgsQU8+G9RYTER2VDL4y/zBIyJLdMcZpk9E8nLtbHE03zX6D3FkNS
cU1OQgw4hhOBXxuZOoS+EOg4x0wghFxCxHFUfgWme3DgoXQmxsMrunOZuL1n99PdfEwXis1z8dZ/
ATRve4eBUEwDpXo48cLjWdIN8Cm9e3B70gTsAmb3JeDI37xtEtql7p6LF+QUShPfXVph/uKSWKHD
6YV7WwM8WHXS/Ng6hzllizG3TcZyzgPWie6oJrVleDSV6iV6GSlQAs2mJyk9rwXpDgBpC7Z2KTkk
uvA3IVk40Yhyx/PR9d1bodkyfrrtbt5xF0lxUDMaC16fFeKmm4jYif1faNN3EtJmUQBLQkR+9Yom
cXKGpCwsswVuKX/TxyY6GPjHtH8UXj50uEEFRzWu6ce3q8eWe52YbqS1Nog+xpXmw0qo+XP1G8nT
AoQ1yvCjCbgeb+ST7lWeePo6Gf2uqkl/m1b2q1TLAal+5SKEBluw9srzXwDAyCqurDqUAB7Vq+Z+
5e7BK3b4RXMVu4fpADc2Wqdi5SpKw2PKsWSjGGN1Krfc0sqpdeczPs7vhBjhgVEZerdQcs39i+fQ
pVHqBaCOwdyiT0k6b77yLMmQ1Jz1ywlzjSKAhi9u+MeHuR21C49fEO0fIioLfWFFePLAQTLqIcz4
86CLV2ODfIOHEg1bk4L35bbRnO9izP3aFi/Xxy3EMV2BV9NS0gTloxWtsg0pN578vHkwiJBYXK3g
ZuYORdEdi363gpCzNp0aOsK0HX3jOMm6vv+Is2BZyTieDQIwiNZidbyTYvc9Mt6TQpsz5J6HHgLz
kRGX/C9VEmnCVKmolv8ZTSmZsOMdv+jt35SLwja2YshdfTyc0kFgBs+w9xlhPMB52WEyB/JYErTL
Fkb/gWybGq0Gq7WP5/syejCnWpWC3uqbS3z7UPc+Vc5h7ubZU8RSMKzcWiIMLjRHls8XXTX9gyDw
2jbWTqkEq9mDyBs3qiUhq9jwLZQ9iuf718K3yRKTuTgMvZX0nq9U3Uubm18AAcZqpirBI1AXfmPb
tTORPRrioPK3FV2RuM+tHsZpuu7m4WYv5ai1VrQfSRABOrEIxhVgnAst+2bIRBdZdidHU4fWvnWG
yA4IcA7uDcry1l+6TVx6R+eahpfZq8bDDWDOiKac8Romcx8/TLJQ136v7ggs7mPh4fe7x1mo3qoy
VmDq7BauWSz/jL+1uxlM2RVL49FkGVXAkIDNvQmIccu/iCfzXbU4URqnkc1HZ49NlMMsAUjfowgQ
V58NETTnKIKAnHkvYVxMPhYNqmf1YgRo9tSv7jAU/4MSoFdDS2RYUxq0U9+y0PTV7dBfgHC+byi1
mpFADFhxmJsTCb6BXPbNJGgYYyRikeF2vWPq1AKWNOwJ+fPpwZlgeUQaERtsfkwUpVfb3ZDUkl7h
vH3SqOIoNqUF63g543XDQeVX4NcnDmhgn63PKntFinFqYiXach/pUfLRE3dJGWIMuD57aqJ/bEud
oVhQVNuhlKCo1K+30s2cwtsaUZkTcXt7H6pj23Z52uPr26+BoFDJlfotSU/QvQuYhZ3tByv/2ZxL
WC1jbSb2/TVHeWX5Vv3tv7DsvxkoKM7boj+dnNrknJDu6CdAUPrVM9d9i6Z4Y7MZLZQNyFQQCvn7
PmfYVxRCzp+zDtRZmDahXeOyhBoQ8nfKc0MdpeufqPuLxRe+JzNimlPrp9/J2TP4/t/o79EGkCJK
c8QV8O6fwMSDBHAoIZWUIduAG4KHC4CA+m5vPe7x3Hc0ynQ5Il7ZSIDpGwkhEwTsg1PDXCCIr+Ik
pBbV0l2eUlSU1UAtdsAQvwMivxIZqmmgs/qkWghivjaSdkm8uLZpKsmEfGu8v+13BtYaFmTURa91
4wQZyrWkCW+o1AdxdnnwRZORf/PFMp/B9ZmfpN4IpbZZtbWz+9JJwQ4iYXEBz3szC7Z8VkaS+fEy
mzi7jOXbMpAD3KPs2wUMxMT8brn6EmEE1uWrXerfgb1ZeoinVGUBqumrBt8QDncU+zKHIiDMDuth
K++b56nc+bQ3LoA7+3dPL4J6OLAJB9Sxxdqnn6I5VdHQ0EOihLx4dVq6/bVnekxUUdjzb111vmV9
SpSJTHnWFfT3Gqul80fHn0nRXUcMTaS10ciQrYHW/5Wwo292X49fIjKCyH8n8Ybc/EN60SB8K2jQ
eY4HpX492TsvVJXGXORexJ0bL/1EGMM3ZdWgISWaUflMwZpjpyEUh6s6sjnX2eN1oHf69Yw2bvKT
JU+OKqSwmXVR2xOuBKiIioXs3AfOqnmSYlhTWun8DYJWBt4tClC1SzwWozErgTdzmo0KQy1+xmCS
9HOeNNKFa2+BXwMivt5cfOc9W1XoEnnPyjyotX7Y+Q/WtWklJ6lmmGSWR+wHWyXgklbi8Y4S0pAp
8dsWnXH1b0xfQCSl/HNPidz4pkzv4aQgO8Gir+KFPJRYAUvqpBs2xcnPq/gMZWIpwuf3Kjx3yxp7
SFpDR5V6HcGrHf+CmAcTcB7kIVkDXLglHkO5Tzs7eFd+cqzQPD2P9HtpeSWYcVIr1kjorYKorHct
+yve1+DGDPddFNhsuzhQsoOXie3aOpJtjeGU7jFD2RhX8oBD9yWhsn2MqxK0faVtbYrxv5Iccd4j
kUxl/j/5mfW496/jkiNkjeUMe+0UoU75XOC0QHJHbCcTjnZzZuBz/5zcSvZ36CfcOL3SI3eITg1M
SwufG8e4e0+7L70ZSKvjs8TvfuoMlUIEEiaisK5D1M0SeMhfbgVfd+7C145SG/N47WUfQkZutDL6
zfSxdI6jyqanq2eNE813jPLTBZUdwKzrW21K5OckJNSC73RCVP78zhedGqjh8O3ZYjBIs8Xg3KMw
A5B6UJV1anoFob87zteX1qUUWyeQ/S1KL6AkjQroncug/i/v0OeYaF0zK/FZaKc5EEaN2UJEPqMF
YjUIgMHl4P+xidl2wOhmnn11TWXuotYJ+TCx9/3HqdDClRAeVMnLjLcjESYKKQhIrNbuZIpsFtq8
vRMnQkFY3Pzu63fj99Y7I2QHESJsehbANyd1X/IoweJFIS+k7FcuhcBe0yTHH/51QIPYrTmcVtPe
Kj9iF35MwQcpvmqd/T9MKSogXGhXvekLXd/EgkUINThJRumZaXXaq/CFEVwXpJcFLdxWBeCwQryF
Wt/y7equrshECiYyjXxK3X/ELplNNt8KTpzZ7csTn/uZWcbGLegAjXu/G6GCxvYb4qRosInISpPq
u1S6hSOc1DqjXhUrfIAbjWDHnedrVH7YtZCqUmk9uttvJVB+uuLjqvn39rSp8lTw72vcuLX+rBEa
PbYGETkUFc9tFR6zIaAYDqWfcaNW+sEDH4gFfsnY9Wh9kXLTukIkjbjCwCFzVINdRkZTm0f/pDAv
mkv2ICWATg+FNci2ulp7RASha6pz+bY3ZrwsuKu5R9Rt0TJR1Jv5G+0/j7Y83eEI0mfBQ63JiRFQ
3EqtVVLrezc027bv+LPgvt2UTw6c7rdbtIRL8Nnmb1V6V3JVm48hVJo4KlWj5xxucYhjnPPyJW7y
xZm6Y7XyDO+F8N4vasFfPn70kU4M9wdBYfOGzyDrIDESAIR2Rzvu3rCFxJDx9tj5JPzUOB4fPMOT
qvlRYc6BkymLma1dzm6egETD1nXZ93dKTmr5OJuVcqtEp/X9y0DCC92qrB2eXqFmxiL85vQ1r/N2
z45MCd2qezuZ+eUUdzq0jczPp1uMrr+OYqYW5e8EisLPyFl0fI7sEqMAczRpifTZZH8DLF2ewtqc
NyIBtrb51+jz7x7H8wS9vxrGMGiP1AfVpGBQ8U5Zj+O7GTPer3EcK15Yy9Gs2Jz/yt0a+r3K3+J4
QzI1gr18d9jWl56zyHEpt3fTW1krnxIOdlkMtPOPSmYJjxpt11xEJCbtgU+a3/diFLooo9/KAupY
fhEVwtbQ+ZEfWAec+2Kx/NnRDK4xIw4FhkNA1xbH1uFanZHLv6Pj/WgICDZUYbN4DpkstoECMysL
vhhV6BF+1wctq7IN31of2oEQQV1qOWoZUO0JWt1oNrcuTUSsCHDkedOenkJUjzf/FoCqO7HrjcaH
GGpKcVkVx/64g+2Qp2esfkK3V5sUwaUsETcm+6Rb4g6ZK1kTIsvGKsLejH/Q1gA1p+hbORAS/ETF
W3gLpeWoS7gMhJL50g/GhIUcgmzTEhAJgVw0GXFfMLxS9l1PBtd3H9bPZgYI+LQmhGPpWzbr31az
j3ppD7DGsIxw/XmpTEc2Nnh+NxJ7ln6XgshfpF94uypYPaUUFjKjEWVN4aWQQAO8gvJ4t2sK8xId
qdyAOZtvj/MQgz6z+Wb8jFz79Sarpdd4NImUVDhfLUgwKuWHx/Ryy31YfUC8u15G9XAJmGtBsm1L
KXAh3IkfkIxWU1caMk4vwSEZseDtKLD4OWXl+3jAhzB/qJu3kgO3tfeOuwiIH+OXIK5y8y7yl4/l
ZvVDDjLdvycXAbMq2EGO5zkyVBCI2jEoQ9s1c/hWGFuZ/a24RiellvJnEwo0QY2y7v+GpqJ3TIdq
2gSWnu5lWRblBosPZKJmMwiisCisJ7SiYE884TyHjrtzQjz82hE09hw4IeAC7J51heIsI0rMf0XI
yauVosKtBgHPDVmlHoofRwtcw6/qbZIW4BfcNkX1cpVirKNiRHy6NKVL48Kl7Uo/z6FhzyIPg6Wg
IflsjBDP0pGc/jSiL8qsYjDuUgvtXBQ8KnhuMCNDxurJhGUXTVky4Xd4tGmfyGGjE/ix0gC/kTiY
+vXGJ2FIFD/REHmJkmBqCCMIyQLKfJ0tq/IvJTEwBgaxd7ETmQ2MSGxw3R7PwTSKjpLl/eQhkR5K
coqSj9ESnu8DTQ34Jqe+g8HnzX5iAQeuJGcIi2LeD42LQ2ljavrIkqczNzIUteK0F82t3ZnZ32k1
VuTPjhTQ+UnIORj73sOr9YOpZ8tVqtWKh4PFbbztf4PJkk6AxE+NCpw8uWenfDSOgWgNczC4fsZ+
TpCkpR085/CKLUh/BkaotpYpu89LfbYbNDKvmFR8hnjrQu5wPjmaP2sCV1tSeS1j3rMMfHeM026A
av68dDla7bNe6NHOokunRKKNyb2mUg4xhaB8v8wf/+s0hCVE5euu9zLR6CL4Q0zpfPflwdAjvpl8
Bx5Q+UZrEjd3Lyh2mb6cC+yp0TBO8gYV4la1dPFMxYdqREODsnIAnbTJruaitq2S7YkqINaWpPKm
XZM8DzzqXOSn+JuzQdlsWgHFJoMpI45/tDkU5B5n2NhIWx6rY4xKzOLBenAxK/o5Ng6boj5lM+nt
gV+L+4xqi2KYhp3f9W2ohtyliPDIkE9UteOiXOig91mtzFOPQQ6/vntaxf+5410uCwbQIVO+lkHI
KUW7NYGZ7B2/LBBtax2aJs3ROLPh8Gg+s1I7FenBq6g/lexzOHQSdJOgcYlyBUuJhT3+ppc8Gaa5
Yy1xvEaO+RVvNo5JCfIkrSFlyFMeg9z6Lc974RCa1xETCbWglZU9F3k2km0v19NPDfxyfp53maQ1
ZaZJ2GFKruZcKRbmsF7F25osx6rYy/cPa4/CByBRSft+Pi1PATrzrgzqBHZHfBNdtb9T1FuVuCUG
UB36cAh77/Sfyxk4PeeLhPySS9k0L168/gnzbOcnXDyCC97XfUIRBQa1zII9z2UL0a4OGZpF4LPi
m3AIT+RKzqmcipdqlPbdgadkbnptCAZKW9CI85USFXtskcd5hsoiVo/vPBROqEutzWNmbOXH1To8
jpkzRFOybVIWE5iybQsbINrCWAe0T1pwZhmUH687AbCGgtXhWRS3+rMimvXQNiNAyd22n1bycY/+
7uFDN2QcyE7A+YJoP5AiIWqCGhdPxsrmXiBPDNboPu44SuKVBazsDS95wiW1eGHSGEdK8FGr2L+J
YnICqArerG5M/wW1sfA5zu7QyfFT0jEllrn85d+OqPbSaXcJ9htAo6UMiVdP6ySeKKgEEDc5umOM
eDF1OiFmuqjxpit4sGOaR5NTS5RrCS+D0RNI+1JMgxJJ7C0jCg4jt0B24+xmfJzeSpPnWc2u3/YY
VDrcsNYX9Lkc/RJBE/rj8sezZhcSlVM1euBfdFcldaAgZajiN8IdVquoLGngyLh+xb8mByPefOil
3CZBzRTBjXjIqCldpQDHtlLw9i6+o6zOATHnJFTVZxpDgbGtOzi01M9BFIgHicVBmFqQVeSqma+c
3XphEa9cYYIEGvXp/vRjztCYweYCGFZ9j8rcULMGrWA28lrAhe15FGCtxgHg+hbZx71Tlzl/8YVQ
4y+UO7O6r+Vjj61GECgf2bY6xkEE0mDFphjGHZVjUdS3s6opFydWCMRUVA9VjIjaFJEf/XLTprLC
dhOc9TS40tJcCX/Ap9ykSgbLj+8Y/4VQLu91O4XtO79Ed/oLACVSUd3DI0jLhdoLs/oiXchQWhsT
ExYmLblK093QEgH7JoNg197f6tlOVYvqBL4ECbU87z6DdJeRT1LDxeZXgGOdEtTgvV21iDyA9ddv
U6g+Q0TYOUo6+fNEVZr++VwwhkOwV83yKZ6XT7n+NjMhOJMSiM91rUtd7aafMHZWmMrsInccqUGs
OZwoAsu7swI9WMw2vQNptCrzh9Zxku76UaJN3EPU8MLmNCWaJEj22pf42SZWnpqgSWVbD3MxZNJt
QvvTAs3AzLGe2GckNitIkec2Ffg8VmThq+ZTCUQ/M1muyWX+9URDON/GkDWskSBgfkbKlcYThMba
GEGt9QRZC7V/A00Rppl9vfMxv/ATPESKkjzJJ7w6BsuNr7RKVtsj+2CHTXlEfePJk7H1UfFmN8Ct
G8aDEj9m2LlMJ9UsRnSQSi1NRXKbk3BeQ56OxlEpsd074RPpBSElIRMaSYWf265mfn5H+TnGVaAJ
55gseUb1DLAWSl7zGRWASEfKz6/vpY5X5tVQKpiBfNWJIOmzoIGihvCBx5h9LcEJHr+vjbCbrAdU
+Z3UcMjB1t0brRKq8gemrvGTXHUqkNvwOWGE2Q66H5hbBmnVifRQ7yLRtCx86oqU688kB5DmyagL
o/ynSDhfFuiuA3YJ0C/rE+2s8B+arkzumyiMpw4/5OsZ9aOvB6VUlVrEJTEgqpi0eNstMAilwwp6
EDKAcs8tD9iYI79ibHauFZ+ScDdRWaF06cqJYox4pYzW8MTT44A0ZkMFCBSxmUUS7Pf0Yq69qlq4
9fW3xmPmSBLfoPcRkouViVPoKUnlO1iPbGebMPXj4m36X4YFicvwg+Jt2FYMQhO52X5G5FfqnoC6
1pf/tsgyP9w5P2WdVWfR3ssmA5TNunHBNrTJJuOBygenPtW78NUCOfuP4DlMU6jSfYvuGel0XjUk
kMs+6mtk7ifN2v37NdnL/fkmVW9o2elop3TOyPBovHkniWHdjznfuoAlKdrKxM41asr4AMY+xnMT
Xzzq4WIO8nB8lkwb03PxCrqbk5pWNcNB9e87x+JKL0lL8/lZWW3yX1PdEbtJeRFQL8AjGX9A60Mm
ffqtX1OzGCPvfC3t1hJuwMutxinPGARWWcJMu66a7zg9kQFhBa5PJ9LYtoiHAbYVdWLe06qKEVtC
5fvcS1amP7qp7iXhhqJ63yjIcnN4qwjD3zhskUE1l+1XkL0VFZuUVBP0VljLQMAB1mxAf1t7rNme
KJqqLQqPLCMwNbzWXT2CttYH4K91eC60SrXZWnF3nofb1rJcRj9F32bi3v8Ln0mEmMBq80G67qP9
Hpgine7dXUtd7TbabH/QF5XuzjtDpS5curJ+RamO4SVNA6FOEaJwvVR6mOWu/VOa3sVelLFcshtX
w7chYwu4o041Xefr+AVBdPlIOayIvkPPSIQyukTLSctpCIENVJtS2n6w6SXVownM90VBolNXRDuq
muzWn53rnwC8MBiUU4NyB5IEsSZDXo7LiUkA5WiJQS+PturUdWPytrRG7DyqxXCRsVNFtU9lBRLc
IGeWXDLScJkejwAPOcz0gn3hlxPVy+PvwZ0Ofdsxq9uzy2XM4FaykD+OvedaYF95ushR9w2MUnbN
lkX2VzRv1Q6y/QQG8bdHRWGviPMDJmDIcFl9kJN14x/hzmt2M6xDkr9jTjbQrIJYzLn9nfzxtM4d
+xDMPV+WfJted45WStgpyH/a97JPy2ArsIYjS9frXljFfDQn4WQpLJjmvKD8gJjb07eJqYxb2FSA
/y3unyr0V4hby2ZX9GDEZrYOb26OcZW78EyhgkLUcn2HN8AvIFs+yDJiuF/T3VB2hG+WQVGqLHfS
gc32J439Bj4dViyIhFy2cTCe/CgT8DKotk2haixfsDvv6nZYYO7ssrg39LcWeDzPnQM/dEpaVtrD
XJfsNNRaL2DTZRVOtx3LIo82qTtHfGoW0tDBpQPDmYIrWCB2N5/6BPWFpYbEVnuZX2CQgpu9FI05
EKFoOehagSq8zBNsNvBsb1hmVsG+lGzTnY2UH95tCvyRIIIrA3BQXTqpPgkJnWkw7dQAQlIfdycf
UxsFc0JD4FWkbFxIOExJs1Xz7+158EMmNFl3sBKKnTdtQdlVwO/7EZOroD2g0e3DAzcc76+lBD1/
ProoKWurwuhxnxs7F8n4oVy/RlNtxRKmcsvsUuCwK0ishwmtWVqsmuSJAGi06l2f1wkgYxAy4i2e
2+CqrJumEb5Dgse12pKd7fgl39XxF7xuNuiORylT8zRBKUkg/jO9VjN8xIPfTFHJGBssJxqO3JYJ
Ddcn4wUGWWU4+zTXPw4NnB2V0JhWfhSxeWGs4Gc8WUUdU9XCGBzGT4lWEwEPcxCZeD2p/rpLTK8F
AnqVpD7EcUTagRFZ+nyb+aMsELyyBUPs+T854G3OCH2PvGpfLiAGfpJjdgDPevG9JUBkM21+rKrv
1r5NWYar9C43nH0NXu/MD37GZNyy5CZcj2YjpXmxXZHPt9tcXyif1e6bBlSW6wvE7ZJ/95HPXP1i
qLKPGbacID1zjAspU3iaYi7i+EMtHU0u9R+aEXCDY1tv6KA6sgAGmoLRuGYcepWuQ/Q8soE7lR2G
NeLqLRC62QGs62AP8MfXyJwkmR8i07B7tjXmQY2BpB5p5aQ/vEXaLmy+s53KC7cw//COZr8gZfk0
7Ahv6bBuYWwbvRppS340SyMrzYvevtq+aNGi7+pC/1yewbGN65kkVDvVk7HfwzyZ67wXg8q7T19f
77HvUeAx6azWN9i72zKpnI2VeVz6OEaBlJ/76GrNvE4ljFDu+u+DjDEHN77tqm90ll/DDXLCdBgV
vC1ZDtjp0vCaHUrRj7S8GyjkjfSDZOJHEZFQAjdUTvKYNiWMlaEh4L7SJEoVLOrKLfTOrpdk4yTX
sT18BQNJX2MPk8TgJ1jJ09TQZP46HBOE225ME9blf4WFxB2gQl7aBaffnBmusCEo6xReVhoujDkw
FmoCAUIglbLeRLMaVp0ETGzVYLAqqyEAxsi68G5ZiQK04v8vA5GigrufOJMBCIfLSoATipWAGr+I
zg4a6SfMKrpn1rZQje1HANG/wrmpp5HRZVWurq6XqgmZL0FS8mqt7F2TS3z/x5U0tU7s047yWAEN
7cubcSc5/mdArFClnBxexe0JJkM6FAdQNH5GWt7OzgIy/xjl33pFpo1XL08QDGOVjFfXH+3eze6x
b4RMg60exOhqRP7IqnwqAJYDOwISkGWqKgJvErHwzteutsz+gUe3mM9pUHbHjGvEEbSjQfiOUwHH
UPPUu+dWTjBZvjoCjnqk2Q9/awziVCyJcsrYCOl2N8RT4APh4H7FWZH22SWJUxgjq6g3gCdwDKxR
THA2dCd1FY8nqqU/90p2/vFwgLK7Ghv5CqQpfrWZ31sRW+oQ/HQwlibe38AJ6w5FyorYvvZ+XGeW
wwvTFE4dvd/cpa7V8BALgeu87eezfN0Z+DNXtniKOIZ59Lea6cd1fepOhC4sArXFU6Qdyh+JP9wR
CxYcFYhuh2pdB7XdhzjmbYT4UfQmdD1R28zQaRy+dsoY59qwEUfuFLGoVjah/50vUnfxHeLb0i7Y
X1L4waun6SPRphy9M+aTy7cPZZ/AFpATCmOPOsC3rVGILAJfbCNCv0b3EnPvQlV5wvGXXQk3vhG5
dDORXd1EcAAvnQGuGPf6YO/W8B9/qvJwzK/6NiSl5UJf95kdHx1IdF0dGew0mloZfyOVdpxWpcZ+
qxX3M9OF/r0zgV9XCMQ6/zZghkmksX+S7zDbI5q1T/UTOgD4jj/4h45ApylRLwlsg73U6vLpq0hG
G9cwt1Mje2oRknEix0Yh+k1iJN+rNZ3bxg0kwC3ADYg24PrIlfyI+iINN7/XEK9y8azNK4YkVIbN
KahUU9gNxoyjMwveAqJorZfLyTYIcTY54Q5ga4f1ybZXqtvJ/1IEJKUxES2VTq2BGAis9I8quabD
KPkBL8izTFwKPbCqT4/4PoQ9pC9rRe97iCDY9/7aXE3ykJ2RXVVQaEKeR0bJzmgl7v7kNtoy4p8v
69FTYz2pr5JnKsJptYiGj5guBu3yllrcr71Vy66rq0Z88Q7Xj4OH1L70lzjo3XEPOEZ/6p9gWyDB
JeDV7aKKsynmkkHxrkstzD/m13u+ljP4cvkb0Faa7rpZa9EXdikj6YgJg2DIXAiHyD6Tr8QT4mHi
SPxayPum2/eCb+X7wXmvdMHHhy5Qv6x0W+iaGaoksmkjuz0EQNtvyIYg2ZQEEBeJcHdIlnK6g5/d
Yyt5+5t+mgu39xTZWN0tiq3ZUFTlYNu1DZp1DdZ7puU3Oqhj0cNAzPpQ2EJEZW+nNv/5B0ew7j99
u+/gII0hIv48YgO/eiJr/hhqhVFWFTrhtRtwYSZMJyYpeKl321mVhLVXyDWOZjFEIE7D4ijLIkvK
y+rOLPZ/vj31hohOfLJxwEgiYnCygO34KuihXaz/zYF4gDdPMwB6P22tia9S0IoihpeZv160i7KE
cVpvE3/JkIe1mBHbPOtdx49/iDHtFnTf/YEGYAoictG3+VIQSLrRKrdjBZ3OaH5G6XtQZuXAkHur
E+cU+24tk+8MmEneAExizUaNUVjTMd7Fsl7IBk1nEk2WRp9h16+GPGl7/l2W6MYwCYwrG7C0JIRx
SO9BUJ79Sl7vP9+a4jtmmjzmYDll7UB3wJxRnQkUcDWctr0mbDqarcIjhhXAYqh6fA4kg0NvNJg3
olqpageg9ctZBSISHOhkX5l+ful0MCr2YTzbWJeBeBdVOIlEvRW3Na9vwdlTvyZTbCHw0/yMOSAu
lc4SZtLaC+d+D1hWC8m6vaOSdyrwqNyQokJg6IvPcjZSJ/PhRmEqZRH5WJkXA9MCMR+u3zMPQbYW
IPM/ti25bMx73Giwt6nsBlppytrT31N5cIqJGGNVler3C0ahBi94PGhB1HBAmuEfUoltjZa/a+2o
Fz7121l0DQclK4zyJ9RxY4b/tnw4tbD7BC9GkR5q+7ciPOFOfFMQ1DaigvYVMxM2znD7XVxQ3Yfr
LdkC3aR3safNqIJTeOVvoyyQSagrCCn6NmZi79MDKd2L8PJGby4gqiimmuiRfs55+Q+VeQGdAXBj
IhbuprgaWQ12Z4FihpVJ1H1wI6bl0x6UZ+B0BlIgBOw3k0JG+MkaA9yzRurZJBsY4OuiN12doYBv
4KmJ4N/j48bOmfgJJzJZ1UbrcqtMNt0Jz6QT9nb28zcPLhIbmquOi+m0GvPDkp4NE3WYrazO8hhf
13N2pAipOQvv9E9BysdTA3mTofBi5ky5WTUigTkdjddt15P4D15XAAHjBrm0ZO45YzhEWObQ1mRa
nac1Z++z29D6Ovk5o1JXmshXxwyHJNR9T6kMeReb3UPBRx+4eFHCKIuAQtb3ovwnf3HL3IXl6WgG
HzSv2e7LPvsdbNw5g/FMYPV3etsEK1mYsi1Xte0zK5XV9iXJddN+9yklItPBdP+IWkrsa8TwmQVc
IZSQMvduuuVYCh+8MYi2NdnsByy0gWyWYXMwgSlNO66enmiiqbd8tc20DbVt7cfh0gX3RxBEDSTl
x7shCSA8cE/obgGq5VgXjVB2IFBF/mWjJcuaP29p3fG/R1Fq/0Szayc7SdbsRqwDqFkivzxdfCuI
0Q4kfvtQRC0UE9ZZQhdhyhT20V7y1FLWB9v7fy10LBbpCEXShsPEBU6S0fhZvawXf3y3d597zQZD
nKKm+usLOCUZYDWKdDnYSE7d6w/MeDPsjnOsPGsueJNg/uBJWOGiw68ZOm8unfE7BEYbKCFwoftS
PHqkZzA0470JFxuuAvsUuTRRhRnG+K6MsEmAWoppaTmhKO8QsbKQlsAIs3OzwMLDNBu22oIvm6MI
BI/4FwZVE1ESM5I2arERdo+amICtV5fTBnu5wb53pBhVxE9kQ75UYqyn6d54KbEaW5YDdhsZZ0Jw
VTDYMXx/5xLkB96V8Iknle6J+zB93pBTmR+ohXC2vkdpvUo+9GG7+1JlCG8RvFxtpvLnbxQn4R7U
5DtJU5svonIJLA+d840cWcqTd7Ui4fgvqLeelQ8CjpVsXErqsl7SIoGPG4pfmhuLe5Xe+5OsljGO
n104a8IaKd89fY01xfMVvGOBM6/juHXYx39bYgbq8Gm/ZOR+XwLs9tdcZO9R5V3rcbJBFSbsnSFh
Wod7/8K7AyFvdiL/+UxqPn4+LKpW1BMyv+kY0EA7aGb+i4YI1l5JgsF60mKd6l6yV70NhoEwd9gY
WAEsi0eHF6+zFCy5yklFgAL0xxhhIUUKSTVERQQhLT18zBT8apDnadhs4IgMTPuTyTPJGm26Rv1/
4vkyadYYoJqs6jMNEJIOyRg2f3iqDNmY6YNRAfEB2c6oReD/Ni+pq9NSsXMotRa6lePnGhIU+iBH
RJXL5GP4gYzba15mwZz6kHaGYp8ja2tXrrnTFfPFKRhAjPudje1knn2Tjttiofa2+lgKunAU1EM/
TYALkrDX2WhuhzeH5wFaL+YaWkPMxoYlc6IVRoHu3qAJY8eq/5VRg4ZUQJMxtp5XQt447he4LCKL
T7posIx/BU/eWrsCxx3jF5BcLQ1mpm7XzEzfyMPJzrdoUnbv/6n61r8UBP5pVR5dO1U4tpT0umQT
x8KIgR22nio+C8nThRpsQT6IvD6AMWFuqkEgnzCHDl1QVhU9nWd/M4zCPaEFwOvd4HK9D7hkgfej
FQoMByYdwzV+EhvpIIptFmWroDmu+BbfszwN1jlqxVOGR6UDpw3MqrAsnzmsGF9yaWgG+Kg0PuZc
6Z5AX07Nr8J8VvM8ltmgpFCK2mB7U9skgFpNZNitKuh7hYK8kfMdq9OkVBgdhRas53SH63GswJD+
nibU5ZTtgpvM/oB8tbQYx/059o5va7SaO95xqBHdawiuoyMP12JVq2og5aTQlbHI5/HIQK8g6VIV
aelcY0p62NPoihNFS+VFrq6QZSE+ilZVL0Eo9m/6L8/aQcypXBC1YvMT2hLfExFXrJY+RCbQjL6c
EF1w1wOx4meiLdHSGG2WonaMdghj5RCDJbOBDUmGsjevsEg4W3AbLwKY5r1pAgj2lCjKKMTOvNZV
FRZlQwIvdujZIQgqYa5mmXeXRyEaWApLfLw5OmuD0UaPyA12unfnw3sLHRpxNlApBTqoXO672j+o
r68L8AAogr5Mvwdm/7W5xXf7l/+UAdAClTF+QJdHC2fDg0ygGg7O1KTLx9Km8Tuq0bMRSK09ba4X
DB0DB2Q1VNndqXdpuR/IX/W91ny5vxhffmS5mCpEvsY1bnEhP9DobFgVIv77vPpxZicn0BIcDDPf
wjy38e3Y7wgfEcy1GOUpdzaulaKr+fy+U3/YOlWNVsGFTx+NqcJ/EyQduG/Po4VRmHyXyxj4FemZ
8BV2K1kLZxCMU4IJtDNKu6A69QQp7nYHfFa+8PW2AFqVD/vca5R+goHpVmrJthIg4+0O5j4hPCFK
vvT0xqwR3RoU7i2Ugs5QOMMgOeGcfAYyZJw3paREl4RG2WEbURWVntuOM3ol9RjFB6L0Z+h+w/5i
Wc+0XwwIuNfz+9499xGKA8ZBOhWMiof+5UMqKP0FDS3QlcLGHoeaswLO53HGkg3bPJpsrexFC+J1
wE2BOCH7lDDJVxRLwIfRZ0ZrA9AaiIAnz8iWDVDmGyBWboYKtioOJQQCI8DWlsebK2X3ESoAH/+J
yudAosYVvEfRqs0WfLqh96KytTJ+piFHPXUgN/YCb0JsNWhWO3UEowg/ir1NDCnErEybozOS8diF
gM6nk/TOLKfSU9VmJC3podkFXXRxTyS5KEYBR/m9qxvx2yxAuT14NFSmb9oPedRafbrnZ6Wif9Al
NUboLMNy9HMROx1foF0/5RLRtIAEfbChS/po9u6ndpcoHdDDphyHWk2LpBgk9w/qa7F1GqP6Dd3N
eBjPeguPlXnfoNHM7Xdt6DQOvCqpFi02cJ4tsEqam1YbjC9mqMF1roZQyEYw7EiMSn+3SjD47JAa
Xp7AnR7rclHedxB057Tt9Cz/+Z3N9rG6rA+qMgEW+plM9sQyHwHWMYcpdjeiH83qQ37xD/8UfCQI
HSfBWRMJmb03Qig3wNHX7QS2NaluTkzfG7VMb6JgA3n3stQUYQT0RgarO3lBMV4Cp8ObEgHd7PU1
ehjzdhgnu+VGpcVY0hy+DLPMY1Q+iDdw4+ZlytfMI5x2Khyvxlu1zsn4jNosWB4uStO00WhOj3p9
MT9w6wfN3otHIQfXpDjUr2hKnrXUHKAREbkLnnpy6D5hBokTz40nW8eP/wUV12RPKHsdpChZKQ8P
48ykQuwfMguqV4leRhZHGL8dw/iCQYYuXUxQRqbUjZCre/oz282PEt942tGnEEduvqsh8I/pquPD
hgfzPjS1VRjz0yoUEN6N5B2E5rCHaINGcYs1gOcCODTcBkXArgmsloC/24mtJ7xiC1+5SjhOEmTM
J7YyJKJfX+J90bwjP36ybZHcueFN4ZPsv9/bWcc92RChwAvP4uMP+kUvDxMaNCnNB9UHqITcSX25
csvEXTboXtCQWGNWbe1wW9rOtjQ9sZWfc1M4dGOnsD6Fp2TdQ92kFeBUblMTcE3kPIUdLBIguJvn
TQos1sHJHhrk1y1SxYG/KwOCiNKQbddTzwNNSGvGmJvpWk9A5mfDjrovzVCP8LQ8pSxVfT0nwUYp
BAhFp8uBabq2WoAnWTuYvO4xD5C3CAWpWyywHL20cGvAMIQenAezfj2KAX+E35uNJ9NicBpbl4M7
6no7DrvvI02UzJFdLy9A1HI2zKZr8Ouy9q+gDe5ZhrnGgWmfQhJ+xngmDbIqXu6q1/Q6Hmh8Z3Mp
flma2ioyYn15iQMRMDWvlYMObukwtBu2/jDt6j4P2B1qrWn6mAjJUVjsu2FWgeBw2Wz8asmfJjB+
fzk5+gskJYb6ut4IGTMv61767j8uQ9VP9dvCwYrhG+frz0TtnD4ncPE6kbQ5pNZPcVHOdkx8GFFs
JOG/75P5q5DkzmiJHYdv+ULgkalLhiMv8KpqVdoi0B/n7jp4aTkt2BZGIAGdVKnN352+o4TPAyvn
05aMsbgRIH6+xtIhb7WLFOmDBe7xAbvz+otLNxV0KzWlCVO/6c3GTwvh90zsrj9oWwgVtp6rNWQv
huNrX0BAteAEYkmTHV542iiVa8ns1x0K78HY9mq2FoAgrNQSs9iKPqp/3vf3yAeOzOYB4zA95KoX
YWHDKofvfMZFf/WhrpwfkQVVpZ8ycVbmbHY2pDb9HrE8VVgYcGYV9R24TaUohUSpRyYhHq2dLrm3
SObEIqBwNezjunm3zFvtur450YjdXATI9ysK6kXNiDjK3FZJ06EQYHxMNVcvC+M9Xgz6yt05Osam
rh+7XLadn0idQtLLUCOla1LodYfuUfQBYsQsBjkiV/srDDD1TClsuCzMdc02uR5I12VZgOHQ49AG
fW8afwNCeiLf/Cc79q+KMOttG3BB4MmJFlDzzCthbSBAQ+0Gio8BK+WuDB4xTiNs8lQfcMMTX46R
5Cd4EVPZB6a86cGzPfJDAqA+MHVllbYc7wnNt4/hgF+YRtfdzfzjJ5qohpwl/vNjSm6PiLiaetoD
1xe6mN/uy7+mhsnKgKuT6Lj7NaecfAiDAcBDJFUSH1MrdS6AmTPMUngr+Vvsb6YFORqgjUJodKKc
iwZ1t2x1cM+575JqZfTF7MYltv7l5xf8tW610ptNwK6uKod+QGr1lJS/4Ro+MGenpv34vrDVT9DY
gLbWZAM2uIbiwVbaYPgC4xI6ZTyZUu6RrVj7x4tyNX4yPxoUSmOE1AgC+4hUVRQui24QS4MOWiPg
LAZbw0jByUOkAqVn+2+79mgDe+dvQACY2e+sBEJcvcDuh02bTE1u5btdOewbvqT/H22AghL4dLXg
Csyp3SQtXRoyLwcnm8EvpiJtnvOr90acGncpBqCEo2TQnf8b5cK849ZzkgZJhLPmc5MTce5c0NQk
oD2m3YDy+Jisia73pUvBZAYXJ0TjZ14+gYriT43yLwRVvUYbGgpvUxoBZGo1geOFUhCSBDbL1P+V
M2UqjfCSv7hGS48mYTrKZqL8Q3scDHBUiY8erPAbv783SbcvkJbn24dHIB51/dskUFsOm/NBKQnD
1Nz5PH31JrGclCM7y/hLwMF6e5Pn7563ZXQnz0RPUmu2JQhe2yIa9dcuVj2eivnGOsMgruP6IFCL
xiG45xmj4LVxZFJpM4FYpDjbTIESXcWJxplwjAiYdeXFf4Cz8K5kEzSGEHM3RiMrDwjFmHUNqzlm
YSLcwro+fpPH2+ygP0v/VICIh0YLVgexA5hTAQoET9pzN5Eutp0+ytnLZSsftp7xgPzVMrtsK+KD
K2bm01NuFnGbXJAn4gjxwCmurPrm6zUKoMXatjDd/QMGZK21B1j0h0f7scpu084SER1Jp8KYnVx2
QOQL+3+0RmZntD1bfLhMhbjarEFsL00bC/JoPmZxLIszUgk2W78CEybFyY4i4NrS5Cwk+Qp0NtyT
nnQNL2u8QPfyBpLz8htUsz87iaoVLTJW4KuidLjcgeFKvkmFBD0jLy9BwLmuU9m0ltvuQzcumgA1
Tr8tP9xsGt8I+0su+oMVHnWtceyzYuIWLSJXDRtdjrCu250qj0QhY1k+Fubirl2Ql5FNjLKfXoF8
ZsElOQsLmF+7674wMXFzDSdaPyCQBJyaAxlUYYqXS+2yoWahKnY6HGKGQ2C/Sz6kWI0b1sfZOwpY
LDClAswEoLpuPIYfY7H0597sbYx8CbwN7W7Ef06vqbrI2gDZpIIkXpUow4RdEW/kIqcBXjqw83E0
x4XUUeDazCb+GkwvMsGNbP5gUenJg7W5SQAqlyfZ9+2KayDTZdFMJ5QxeY4D9rhoQDGDWiHxaFPT
IjmvGadH8aDljbn6rvGDlTATlZJYc1adKy3j6h3oL1gmiJmvZ6tK1O1cnRn2baFyxjcy0jJIb926
l1Sa2dXw/mEK2vi8JDMJwkmToRabSJA4iK8weY+mXEuAV7EYtI3dUx0YR3/KrgYGQcAtfJn8QS7i
Gm18Q+Sg+NySN0AZcLLxJfQ1FyNMuKmG2Dk6HjY9jGVQzwIPEmprM9jsfMjsm8SVlziV76MIXtZW
d20rmFUrt90QB1qgjlL+G1KKfkvm07kPPEIY3h7Ea2dpde0epnXicGPaXKRrcHyoz/Z4jQQ3Ad1e
2b7dywYKHFFfXMhwJOiM+VVH7BGkVMXGKe72VYPx7ing37z5qChaTHd8//TH4a6lgDOrtDEVLR56
PiHwm8quPiAdgXx/xqTHLF/PEyapPNJj/E0QKrw5/3+MHTl0tTmPoqIIVbj+yElF6Sq/dJISzZY4
hek+5Aa/+emSGeLmHIr0LJhB3weQx2iAQrwHxe3pmkFS78WRWX+9IAEJS7nyA9Q4QEL2ySiTLcyA
/OnEBTdppUeRij45JdsuJQ3gb2i58DmJ3Vj4FkJQP/iHSiQEdXNGDlo0K0kR3pk78/vniFZyvjAY
BKRJvezZTWv9GN+rIfS2SsUB2JsJAAj9eQJyDQVlSOjguz4hCTEqkyzQjuDiT5f1HbGUpzRu2WTq
58NOrGBPWpV6LjuHJKMNGushcPEvA3RxYhfLtvfryVndt2F+D6cHG1tZuLvxvgwbJRbLWN0dCTO+
vcQZ7diep3ZvMUe9E3KDiDq9o0Dv0EysKP4Tw5Jb7udpwPaIORyPRTEJCBq/czxeyGTnwg3L5VPL
qlZV/2WmpUuugO3/U8D5BoTmbk/PJgV+/lSdSerhEfDkLNXlQ+P2yc3+PdGR8cejl0Y1DTYVIK3A
K+fOA3qDZp79Shbh9+jZtcLnxxzH8LOfKHaSjKTZd6M2E+6kbxlYkAFqqHjeiCJ8efETsBTK+0gB
sGCHhfeX/DOBqXwj351bs3eXyGQAd0noSp6pNcUvTt2Ftm7sa4GshI8X0CLdlPJZE6XFINnJGibZ
Oj8Y1z3uGMfV3US0fbYq/oPEwaR2Od7otIbJIbrVdzetrfcI33KezycIMs/sv11IS2c5RSWS8INC
QGjRHD6tvsQX2erdtE0nhmhgAH57p0VY+VR9ZLQnbhDyE0bdIl1yabWn34UCsR5CiB2KQUM4NSoJ
wfKpENmMSOtY9syjdwqQ/xSYx1j7yQPMJ8Nw/QlUdooxhZVygH4Y5mLgUFouZ8UQjHqJ6E17FRiA
Q0HaPkE7PyC810SBetZQtLDwMQ8ZWBKTuVBorjYEF3BiGucPNMACcvnVVwwV+AtbCYI2vCPugZHW
P7eAT7gP+2hR2crfowFgmXrDkBKixDezH6u/vav+mAsfFJGD+V1kx78f4EAkWuXgKybAE2Db7F43
NkAPjjyPkCj/qn8TC79kf3wWrCYeE41PqYY4LMCuUrrfeSYesAN51p/aFqJ3kmMX5aNohYDWhnCB
5+MPP7E4njg93TLLR/8jBuiaEekegDjcx8xH/JM4b8FOXbXt81e8ZAcGrcW//A8yQrHG426bjQiB
1DkEacyD4gzkQ90Y6ikenC0d7rx8eoKw2aVYh906U9UY81+PdPXwPMC41QbSFyNuenH5q33lw/33
tjkRh8lyyXcO2WO4oqis98D7ZA6DwySAao/DLpS2HlKPTJEO4EPbS0OqDl3epoFs9oRt4WilWvXF
Dm4wT6F5VR1zCpMoDLjoeP5d3a2MB174Ov0qYuZiJw8+CLc1h/+OxFlBe/S2BHYLFbnymenu4ct2
gwju8dz5obNRzfBXipzzSOYje3okgCUjhbpR+uYV7GSuiGR1SkJ/2KaaMMcEqnkwT+J7hhuX8EKE
obAoFxfEf5loX+DCxTh6oUW/lL38GlxZ9sHTiCiFGA+ecv6V/wExzcxR5q/suwDh+Asodkks3llk
fcuJmrzKsOCihmlcECYWBqvUT82BE+UXqhguFpph0hne/umJzTzKo4Q3prNTcXyd361B/6L29on/
w/Ez2oEU2XnsKhaaVk2pJGiwdHplweswILKwzO1CZnm1E420srsMjEhnrtCIVWbCJljxJldo4k9R
hBdnauyEt0mN5NrG6uBr7xiSsPu8JXszgSMVs1tt4F13Vss0VqHhIjSIiks1j7XIR44rbQ4Aw5Wc
LG3rX5kI6OZtrtrWTesLIG7BmDyShl8U8p1tPnxsWmtPuoxFtg8soUeM6E1V/H7OsrZ2IMYChNfh
cbZq6k7Bzrk4T3R2p2U7/R7xuRkugxD4CDP26lIy1ejj8pTRBnoCFt5jQypigpnF55v/sKm8/a37
67/fZvn2/RiwzfsbBWGOfVayvZixgX16JwTolA2Xab4aZeXSpqozYAaCKO3SaA/4YjA/ZHhYtXVS
jprUs8/3/9JBOiPxhp6o8211VDQmw7kouw/Q+iTLFwzugCb91JPf4EJUBBfgL73Glpikr9wHE/e7
0wPCTFy8UKKdqeSHlZ2rRxicVKOnQNnsgWjFNchrDZFz0rtxEZZVpmCZAKQG6YFxmbYpEQNQhd0o
8DYp5hG6rE0nDCofS8C0hNAutXcClINF8LSE7yOzreqm7mawFL+RbN6KDM8xaDKkTCL5NAkrfYNp
zolEwGbh8wElWsXI/StLWetnobC1MUQ4PB8auZkoHTvwGcx8L/XqfsV/piVtufTOhQDg/xQkcAuR
p2Aa7v2ROSxnu9tvbvU3LFJWqIYmtRUzs4PZomKLvpZcIFHUkRRKN2ICGcPXaWTCKztTz5ZfPHSZ
/hnWLdtQnhvluPDIJZtBpMhU9y7fe8I2s3j9w/1R3rLzGblUd8/hj0IQuzHMyE3ZtaolD63stB5O
LsTSLXwQMJVWL7QEgf4mD9HG0M4RDtUzG85OD2m9d+tR6fJrp4VCUpdKBQOgSL24hNIk3mWeo/s7
dhZKoJap674Mrsvfr0XIfc2oOLqYxJnRt0h86yM/v+cOBfb9tBnIw3zzORLzo2nAfDMDXdfB2oms
64PYnkbKUNkyfwZVFk0zwS4izK3t7xWp/uIHHepjsKqzRnAFHKbwH2P8eraCZsP5rtRiBaDfhPqE
GFZ0tAStG9MoNFuwtxBtxfjS50pQwHaN/7WBm0g216T8JX+59U8aCUPPEmCMPwKbjPmF/88PM8Bw
JvM1i1JN1RAtNOXKbPdGKLKOPMqTb3m1MRBwl+bt9SbgIx7VKoqkLy4olxtyfitxr+sqU2zrYbtB
I+cU4UJ08WHsAug+gO6L3xCqkYKKEo0AHLmD3EvfAiVJBJX46iSVZWac4VFAQcmWCxtx5pFj178G
nMS4in1Aokvt6z3gu/BQSSCB/Q1FlPL0yopY3Y5nC+FTRLe5LLA+25YfVGExkufxr0kmCA56IglQ
7qfg/El2JvOx/lSYGedf8XFoiSJBVQRgou2iHKZc4dyNs5blpql/dOEjSXUm9eTePsjM9TrIk+pQ
8H3/pTOX8rbPkfVCgQGqQ04hrwWY5SmFIsSiicsigUq39lNVq+65fLYPfthH9iGn1eE+NLifOj1I
qq3Ho+WY+0Cn5DNKDh2TBDa2Xrklfd5S7Rz+LkN5uYxEi0OpuzN6x7JzHXa+4ufQy2VqbFqL6rqJ
/m10TUg3wQcS1ikQ5FEF7VXGtyDcS6jeiL37bZ8j8KmMqLKMy64LnnmhXnQSZZ8/AVySuYFrBSNf
BufZiXXoLHO0xi4kXwZQ7mEAx0/FQesowPVFFtDs2M+hKracOVn/vjMRmu6Ocq8J7SKnbBVH58D/
FmnyhENyygbbbsihq4xABHGqSqgg0+UfMh8cNv9iObx3u2GBKUv+fdRH5A2aRHacCOHjOkBfW2AI
cZvAO1RXIxpbouWYw7f4SZVC3C0YgunAV02iVYwuqbzBMGIxm0JwrgT2p2GUMFegLq0OXjlQqVl+
34K1asKnGyT3SdEahzYx/j5i2P0ShDaObfcD2FH0tpK9rM//UGhgWHjmDdCTheTMQ4JyBysJzoOZ
zY55XOTRQ6WNXWynPhOPjeaNAzdpVBUDASltn6Uv7V5arncHn3lzLqzxMSxPRfwshZfwJA5We2hf
bhs4zAXEVE7IwjrlQk66mBhObWajjEmZUtS9xFolVTHKZNAXDxyJW7z2b3qS4dTooEtfYTW8BLKa
K9H7yXTKQPWyPaFOE4I/dKa88pA0CO4K0UWXCjK2IeuXDNldjzJ2NriCl3dj4/PHDywPCVh3vSaM
d+cK0hzlU1uCGFyDWUzLaGNOYphxjAAcGzZrvbWLWYyBTJgCmcrr/wS/0faR6GgS62OQf6AKoGbQ
C9jBhL4UAd9w+T0p2rzurjEAUveuqKTo+FJf9oabZ/iRgGSuGb9glH2wOXdmjBq+FBUFhH+p8mAR
3K4E4uk1eer3P1tItx1sgHouETiLCdIyI0N9GFQKo9REreYt5tM/zzAbnESsJGqXI4zVDcetRxdS
t3M8iJhKnVb8vNlfqplssXoIT4smcfRK925G4S7ocgR98O38AG20j8Rw1T3dKvrFOQs9pig3AVPP
0mHYR0K5wt6PS1r7cBWtzUwidT3aaKxss71u+2Tpdojy4jn7jVTBmo310xWUdMjSq7X5sEZqhGSv
tzhIrOnMS/aqg9YI6Cw6arDq1JkC9HQDBiK0u0r5UvI9QfXxu90h13c+KrV5BnZcHAqmcn3cCv71
ZwCsTmsPw2ai8bi79bTUotzC8/c73BYr4mSc8QD/VSNaegQNQhqunfALpnY5U5HmoJBr67iNJ/0n
9YLGRt6jkHEVhLsNYjRJeZfNeK8Sn3CbIl54uVLi5G76wGEC1qx2BEb5xZF+xKioX04yxsSgqipw
qi6ORTf6BLQ6vSpX1dsh/7IsG3dgBhEgtDpDrha5W4vuNAcGgqiYhPrmsGBZHZ/ayc4qd6AfxeHd
eK/w7QkxPEs9RUUX7nkoiwW4in2DrO7vUNbqgrGBmmV4mNcDbNzf6J4SNWoyoB7YZrrk/b0SpNCJ
NTIAPMSwjXvM+vKpB3QpcudPb96aJ8VYAOJoU5PqiAIjXPwmIomn6mPZzT/tQPf/Rh3W7MlHgXve
AFgVFl4GpFcM51tHSarWuvVmm5zugX+ZgBnXJZC9Eec0LpgvrJ5/MoSG8DZlRPy8UM5EKup5Q6SD
X9WH7Qjgg7Ua27fn+e7BJd0/HZ4ussyC2BDAOKU2OtaFZx/eiSEYXL2y6okjq7fzIKP2UAQmXDka
0H+uFnD+xricN4rAkRL3rc1YN7D66JaAdGu9DIrbajbzuFo+qpqVV3R5vEEIN6hdfHif2l7PXFrW
TV6J7jX8DhqzEi2WrpJX/wb1D225sCHmV2vzf2jJEIgyaFPxrSUKuRtv4XV6nW3fAvE1BHvISwU6
TW79S+P8ECfVHXKkrwFFMwBKLsbAiB3R+bOlGex/rUmlF4fRhBKYF1jiyMF5a3V+jcUvHeG9kEUL
S3zxIiPb5/wwf1rl/HTfTmK+QCyleavGDYnYuZA+I9Xt0BXlYps3xJ84jjv9LWYeFfV5H9uuTh1E
Jjc8KBvVfOgELB+PHBZ/Q0Q2drJxlaEC7Gd4nq5oeMsnj5AU+KsPEU6hqLHtVrkmn9VBj6/KSoL8
Y8qMb+e2QykhYo+dVapi71EJIMnBlp/MIOQd8jWxydWZ7cMJ5MmzyBHSWZVEe45Gt7i9OI1rSglg
/jSyp3TvvDGAWVdHYhlqs4XrVTnLXhpai9QJqjHn8Lytzds8xB0GEBM9T+ukeyJXiKIwFR+HYbWI
uD8L/oP7C2K8koWPBHWzTKB0536yd+xr+qBGgD5qRPQWXH9UrtDPu7TObTZSFHv4D8mmWqFTCQ/D
cb7Egmg10BTTaOm6Gc9AkbPNnL8LDVEUteTrOn6x/mODDcQGfG5suODNr6UZa3vc6+o3W4Lpej9a
ECYWrNNItYH0Ub97PdhhrpvpePDhVHgMAtyKMjI+DW25zoCiQDEOa0ivk9AvOhoj2Ep4TS+Q4a3V
2EB59oPm3c/E/T4TTPjhcQ+Ut5Kq1FjzRJeQZwIR91MQOWHLcjNBKd5wNElHDetpRghTG/aTmuSD
zMfGfo4tGBjD+R3TAeWcnhE47vilYDrY3FO8aWcx4EvCPbu395i2tW1WzxxwGjwIdhGENGZpk31F
iExI+cBv7UOq/lgePkKyaJtDAtC7PQnpGe/5qppFVaoHG9TTS0L0Hn89xzfJ+7lix0bAAwQ+wCCf
E2hLX4Uv0STjcWU7Od5zLbs8iBHfEhkk0Pt/MjgYfX2KH13zgTYAqMxOPRkjjO5p79fKlDIslDJ2
DFsOinDhgMfqUMDsZc6pEfygAB8oOkLDjKycchhL1bB51TIjrX/dq+97STnimGbaHiZ9QfufEvfW
HNyV6WQt4GnwP5lfBXQqAqbl8gKo1F4mBFjrpLQl9jagfX5BCXDPV5t5PyAbrKf6tKot5rXySnYI
YsPSwMZVRyWiE9orFFLt95519ZzocQAm52PzE5UKlDEOIeStqUgbDsBZVtXhwz23Xx/p5uc89R42
wxvFsp2rHQyhhaJuWaSqrGlxt5KVqAQGmB5bRFxO7aQh8MBtuRxH6WUfnqgC2fpASvTGsV2GztfY
Y6gYdZ5rCKXJPTXJICPWO/3DQZ3xre9Fwr2mITh0Z8B2Rw+Ggy6Ysb6+i+YNBZKx7GQpStzcCE9W
T9PV5tT3ptjFJdfr7j0v8ZRGcdbcAaC56sIsSYBUYXMtNYUN/rOiPmtbfuimcEFOJI/CeGgNOnAy
16WqOuiWS/jyJT1XRfTm6Tit+yAIi+63ybGAyn3xTL/tmChwdTzpqSOwctksgSdi946phUWplpL7
B3dBDKkRhHeNg9tArViy+GWW3y4uUJy8zZ0mVTg8PXmcl9IIAs5nhCWGEKGk+BoKgDf05a4XH2x3
PnEjw3Jd4BWHDhafYb4Y1z1BsUFOZRghnxZo8TOxFT2rBSZl6FdPWVPJ8j7zzOZpR0OSHMKxnBQ/
UW1Mc/baC60VQ1hsae8khsjii03FGq56PvcyAVWXq2hxrCUOyf5CeZjRTdqWoXOdPMitE2/MlzSL
s1/Dw4MpFfpLdmrl3RWLsaPxobZisTm9iDYpCZntS/+VJ5r4/Eoi7Z3NZ6sZhanD0Ww1NhLMSycm
IuhRP8HuQ4caoUDSwDxAXrBlIIk2lgUEobAQE3AYi/zgzkbJrBPo4j4Mobl/ZrGkShWgY1vdu4O8
EPzVtu5Dh0xpmlMHAib4fQN0gr3Ori2mAryIiEAfrYAMtKOE8+lhHl3+wmC9UqC7LhvdIWfknLzN
/zgQ2aIeQxflQgXLQedpcZ/Nhh34yjEwvFN7EjR8/Ki+MNVXp1YhnfHCw73Vodq0areKhQ0p7PAA
99OeQTCHBsWKRfyQRQexi544hIG0PkyvJrsMMxIg3GaUQzbUsETlnoWqAMoQLAX8Xum25PGaY6QP
Io88teEfckIrja37G7eZX0XZMzKXpREoqmiD7ifyNPDW41SGwOPdZXKLlW/nhxQMTvSKGaiTqVht
uiycf/yNDwYRatgw1EFzGFGPYoYkQTJpFuzhWrzuC5b2bOmFdpknCYWFvee1YcAdRHg3KIQxow2f
TOgmEkO8w/4cSiOqcLgD2lE9TEAZ/F7zwd1ErIA3VvGBXLhpAzvJPm6t7DmQSq9KHLenlVXAAu/m
kIYQpZTqKqdI20IEx9I7T3G8xhV9KBoiooMBpDi8VB97TJeX14U0Ae51if9gPnxbGWKjNE9PENtB
tbvAyMttmsu32uj+jYetcK36BYn2TYRs+xMc9CCbUxIw7DNCKeN5wS54UEGRK7k3317jF6qT3sDk
Alfj8q52Ewiw9uLwIBy5b9Y3fidT2xu/Hk+7cJ/ZQoYLUgMBbTRIt/IRe8o6IsakZmjDtOVY2Io0
9k4/LRwopFye3ONB0RkCxLL+m+VxuCqwaPwSy7cBllRCu6tfrZ8uKrmEPh6l8bJPBZNrfKMsy2gL
th+RaIxfbDBPfo2hNuAlucWcTjYMpEAUb1xMa76Fq6mBsiT3l7YSYrp5DitFogOMxJkXMrDOkpH6
XzeGVnPmKsMUraT7Gz76TH2sQ/2XjYSEMSk2oGwAldDdrP2BjuUkZv2wgmpuwya59BCxbKOMzhUU
iAtfixRkxYI0czOlFTvGKIYRcpOZm+5J0h2yvTY0f3u/4DB/PunlH27NDpk2LOGjha9CFTA4Lxsb
PzN3oMajApM9dTwmNTkCjFXTdZ9hQhqe2eC6PArKfOwnsIJ9zqmHHVkm3lkqUVpl5J1CzCoRKiNH
mu7BVpWAJX3dAn4mDEYNkgBUvSZWXtAxJNsW/Qc+3k8GFYz6y/LlhML64pQfLCwrQna5fArgzm3A
FYucw0QWF+vfa/TEgycHadRM7lXbedLYNob4qrPJBTRXM66NtX39ijIfHDDJmLF6HFvUKRwF+EW5
ZW8uGcpw8qkxsS246upQ8S7TM+dp3gxMZ58c7blxUrSPuugaMcHlBAdgichm2mDU7+Z7K+T6os26
CAdS9HE4zGI67RaqbA4OPBYumDj+PAhiM6m9++FYDXkL6p0fe6CF/6+TfLbKeF+i5CHAgzSF8J/s
i71IUyoiYUGPUDOFjICGhbge/VmS4kveqIF70wZ9hzQXGo3eaCNjjMPsuoxPyv9bh32F1MwnMnUy
Uvsa1m1zzH/MO1U3SyMxLvAU7hIS4gWi82aSLtQ/FY+jbg6+EpUwm1DBiVxg+ZwMKVW+qTEbZM6s
2AKbwo55u2fDBuI5wIuveCZKqlVZ+Ld47uHLHdf+lpRyXHC9uM1ZI3/h8yoKsBLXOO0SArjD60iq
hzyXiqGVNgUsktaszjyvIauw+ftJWTjpHvvd33fnPil+xQhs1A6FUBjsvPB/ZHSeAUEy+EOrD9as
U9SHqo5ake2OjfJzNMjeaeR+kGe3yTtJ0yBt8LLNNyhVQELQAFzOwn0au6V58jhfKwTn5qHcMHyA
NlGgoewbBorI0+eBLXfAWaC85T5bBxS8Co+o+ztN3lll95dW7Z+pyxU5EeK3VQYr5HNPFzvNNhDh
05wsCWkCWOHwUrS+1mL+/Zg1J7on7wXTglhA9HWGSNnXEh5hyHOmgLDJ6ng+DvNajrWqkpCycv/3
oghUhF11Vw9CsWFt5JTj6PliOQCFDqhIB5W8PTy9YXIO/aVOtHrQiAlUz4IpG29kR7iyzFzExga1
9wBB/yLIpfQdR+RUQPHbCEuVyQO8B/7eyVkSXjCBvUR5hToa4733tyY4LR13+rSrcL0hp5EGIENN
2rkww5Mw3OpEO9p8j9Mh7JvWvJC2AoJYMopNt9tm8VJQy7MfCx5oWkK6OudNpIspUh1GRa69UmLK
9fvgvay7Co3XBIkDjrg4Dorz/ZTkO5/sSawR4nyb6u0mj1t+7cMjpKW6o5HkOjPh3ZFcJ29ui0I9
3Y4mh4gICqFS3ZNdnjxfSVSNNEMHaNX8DJi7/azI/Sp1fmxX2q9MH6O+jsg9SvB3gEHtjvso1iWy
SjIDOLEBiTn2Tx9eWcPmRcvXPCGjGYK9tHa518aIdFa/hktaYu0zLhIL1rWVQ9zphEpkwmFERKOJ
36ChgbIWcKGWcVV+fi0Nm2YujFNoESXGtugqZbfDxSTbUg70jC3VomhxBBn+PBu3L+8cu3Ubjti0
bi/VNXWPt0ZrjTiy9IRO+61oGQLSbx6LbaJ3zhzfrf0lBTX+0WCFbIFoub3aDwfcC6R5XDgdwljj
PgZj12UO6ddqJdtV/n9s8tooHG/Fz10FH5Jti6kO/bsBNyaHpimVZy+kjDDCFGxRXC7UDconq34t
HMi9iwqAGoqzJaSjLVuv+UeYlluOmsDjZJvq8k0I94JS3F3p96qKpcqFPvNjM3k0UgoQirAW2HSV
wEyJ1+sXKIcdsHEghJ+QQLizy+8pt3Foym92HdYeFEt74ymrU5zYbuQXoHC4QEj75Xj8yp38gHl1
NSDhm3iZRqhR3gdoDwAOodDB+EeQ65J/5myy/mgGl0MR2k6atTMs+q5m6oOQX2vgOCwzv/JKfFC9
q3DQouQMYo/z5ul+3op2z8aNc83X7I71Viy/8OqsuDy2d+rWAc1OTyfYKzH3Bz+7cT+OR2HPZEHx
qK+HC3N/gcXMCvDya2ei+mlhudqdVbjEzSxVj5vxxXyIB+MiBIrghVL5pPWTmjciGDYiegsHzXWg
hUG3T00LxYZ7vhnTGh1l28SZGfpHyeFAQ4FTZskLaV4u9Z5U7DC/6or/JSHIOqotm+s5CmCiyiXQ
gkMHYh6ocItQuCJGEdVrbVtIsRESbrvtsSlFRYmhRHQbtf9G3ENRAHaFCjrUjx5/tsQaEeyMVzH1
DaAbqhjUuiLrfodtX1zN0M91IvPb2Ag6hAkR3elA7aIeTkVqo7EM9cLJQUIGRjS7PyT3eKQ/g8QK
8sHN/e1ANr6fjOVefjaty2a5tCh1HjS1+2da06+3wpMp0WCF5nn8ruyspICiLlRECsR/zaJtgM0r
B2Km3sQfDkTxIGJi8eo1LPtpKr8Iry8dSytKXRalS6h2E439ut3+JeMb+tr4szP2zSrSPDB3TT0n
Q7Ty8/FSD+oxG55VzLppc6iznnuwGViMCGhiUU51P1pWz1RrZ7VNTnPWTsxWqZmBuZeJqOv42wAl
V51a00Hgd0AniA2mZNHjPwqo2KS8VAW5GY8DabThD3eck9fBxniZM9H+mEF4Cr/fbCmg3e86JeNf
NsxPdykdCh//b5vFwqfZXKm9iejXKI9N+HziBC67zh/6mhzBw/zXw+2E4B5MiGO7GEFXL7mge3QZ
tbAoI5c5avPk3S6bbeN8Lm/PlsslP2/ca6EW+VTV4bRLk5Ct96staBXlE0pw2e1r+fxXxj9ZQ9Cf
81i3ni9Q1HincUQvNgsMaG99TwiIZ9XXH0fmcZNIVXEUd+ambX+Gl+ALYZhA6Vu5P72JbKiqgCBg
cs9lDGaAkKL3N3nNysZltIVJXQQ4FDJ/K8dDSFSlOo4oxbCUm7OerW8J+3gmk4AwYo7TFCbLZgeH
a7QFoZ96ptanOECmkHWFvkkJNSlcn5Fs/6BwYQW9T3Fs8kl3wmAyOqL1UFmGIzgikTcXBoIHhEov
teNxpSob013fo5lgnZycn9ca3gZjnFAu13uuGW3HVuUFZLu3cfZGfUIROwrqf8pSXETQ60cuPRGA
Bc21nZm7J4QbjZLlZXxZ5HCiWOw3KvOeOUHsGU9MgiLHd9CRPsVJGE7oMIGE95y8Bc21NSmsPVgF
NteiWH3ots+Ktu1B7ziI7iyTPibrdNTCxnIfTRsjapf+9tQ5xKv43gBU1VH7WGFRWdE2rJZxxN0F
38M8ySOE1v+IrXMvIl8MRRG8QKXV0XE4JYt0y9nRG4CeQwtS5EvJ4w/TtcVH/1raqMO6g8fDAqjY
5ibpBlwL/rWVpB4Twuf3nowgq3thGV/08L2/etb/ZJinsuVDLFEAvBG6XmHk/65TwKIwpEVFzy5Y
zhj0S3SvKsk/nHlGEfZNUOOraUyDbdAHyE1IRqvtAYP5NGBuUl6SmN+6loByfnTPPI/CDnCRF1hU
vClCKftKLGppcE4yySukuXWBN54QgQ5xnUccXKwe8Ji0efDIi1xoLf1wrxzDzlZLEBD4GTdSkLvp
SBFRhn9Tmas/CTZmPmXiuCdvXo1swbH0+WCQhV6OejSbAHPO2yHiC8TGzPDkQRbKq6u5Bj+9SRoT
Q/kHkxpQMxWe0kk9FYoTCi1vbBbgVxArevxZsqQMoyRq7GVG93b8HGtjDBqKrz7uUtzIgTVUwbYt
1eXouPruaw8Kyor6YFuFaRO5GtsBE74wtbpvn5rWLSRyze/33j4a+HazlyxMMaibOP2TujnF9JRH
A3e/WjQLQuoE/MT6jKIzfaqMDXnffB0v4/A4RGyjBA8oblkfGoTRPTFj/Xp95iGQqrTlIZ3sHGt4
81EspG0tP29/QDp/6aC8uAij8c5tyv/KHEYH4PF8d1LAfqyZ/CWWH6prlCpo8VHS5SAHPMTnWPhm
gjptbV5DlGnDb8sGFIsOsnhX5g6dYfZfHoULSmY+wawAxKKAoGG2EIRGAF92Qo7P23X4J8xPLhvd
2hbYGo6ges4rHTVZVD8h4CV6YsL2b+6Y8qCBWWhlGoRE0mMPKhWODlVY9vHlBS0crc643ndr7xhY
wXYRf5cP/H6mLHF8607IjOd/Sa34Fjbh9EBKg5Kb6jhS+QeCK7fKx4Ofv9SqlT3MA1K6feYSJHgW
sXjG3kKbupFBdR+uZcYLUI+7nK0U0wn2+5IE6VpLDngvwIohnUhc4IXFaddAMYeDXWN07d/zG2tW
oMITLy5gnklew3UK4CGMso7Nbz+yGCvsoehd+FAJqyZJaAQ6iQZJFFvB231OQW9NB8UY5Mw+kmxJ
E17nQiOt2SLwQJKLf4I1ryHP930NMFEXMzzRH0IdOTLcnhcLrcG4wLWxsWd+zWfETapwD2S4HrqS
OOv7kZo/EEB+B9n5bX8Z4pZr/dCgatXhE/lv1AouU9wLZ8t89bBk3+VJkPspDPzc6mHdAgbtOKoB
VnIDMYEijR1FsBHHe45q1H5AoQ52DsJEKsKQWXDdFbp4gP1QCeV60euw5HYXZRHtQg0Juamo0/Ji
GNgiDq7eg6bGUe9RWyq67aijxdmZtqwmvOvjLKOyCfHPUeRZHxcAu4P2S0blH/LEgsmbX1iH3+oi
flIrzlOvJOHLAxU2slfMuN1ySJoOKDKfJb5r7uD3/iTWqaTj+PXXskdktO2lc6g20RJn0w5GwwpS
L7MHyMraCGi2nS0jTVXm7ZKrWN+KzduO802kiBBru0uUiApGXeq0l5bhUZMICvgdKubzPI5tbkyw
RkrBodrh52FrjyrU+LzhGZlAW84zY9/OLJ6v/NIaW2EtX95/9tXRGRUwBqLhwIOQHbeI5su9h2R1
0ar2Z3tG4bGMGBjx2jLwEz7lEtzAVmrOKEhns82Vpn37huFyyj5dxsU5lJvm10sz++39T9VIDIey
2ASHychcmKBJq5CgxApJte8IphfcxaHs4im11aUDa8b97iTaxQpxipKBW9urYbOGzPSCPGNJy68h
zVYHgFxY8uxENDxkcnqYgYOwjjZ2+FElxlWfX573OyGzlkRnR4owM5yOWyIjexPQ6tj/rhbj93Do
IBtqCSHLQwaDblwXhTe6pDP0K0A/quT4tNC8sEG0vipR/abAq/AdTh2P5bfN9pzWUi4Qkjr/+tQb
cGRDHPhR+19XMYwhoILPou8zmcgRSE7hN+VURbjQ4Ah7Jh7CNOTQHwlQvyCNqAbjn55qS4PbJ+Fy
xrQDcr47bCf8zhpaQfHxM2GssG8nmQAvONXYp6TNDitcE1QTX6LJs3epwzVs9NLPy5q6rMF3o+T9
BQFyrtOqrTx6ptOtMR9a/i8mXyZwZQ7oJDb1NhvGCJxgv7TZDwVb6ugK+a2jZFbZPV+k1JD654qx
0AZFEkLpqbDnUuyeop70jNlIcGT9xel+oi899/HqAWFkK8Qm26vO8z6VXOxcYsKfEDpSxVn0GS2p
TjGJr8hlir/kiH5u4cNxCsQxwbir9Yu9fZKcBaJpeG/lllj5jhYyhyD//iy8y5/OITFZfswRWBzJ
nOH0d1X4Tpgk0omn4NlSzskQLwB59bpFZp7nF8H6Kz+PidTUmFZBB8HqkMc2eeodKhKtWjdGzQlr
gxydev1Dus2bzmfF27meXDiwV6Rr6mgGAlpqJTuaZPVOZFNc35PLZ2dzaRv3aGI5H46YUFIyJxLY
MwL2CJnx6tX/bDgA55ZqI2z9siifpI2aiijf3GeQo4QYAbLeIjNsd6hOn7QSPPlAramdIDf8s+3l
pSVCTDIagXVvycIjzLQ/Eha/AZuoZGbc9kvKVbyEW39lDa3rsz6bneLxPK4EfwQ6ip9X6xgL37DZ
cxRg9sjb+liM4g9/MJrtQmLFaenaQ2gArj7GT41815IfUDN5rAKtKCJDpGVP2g8ywQxmQuvKmZWB
iYjEZ1KswV4tCCPKYu9CeiZ/FYyC2AZikXCSdziwgEUeY0udRwwIUJvl8VzBkVijiRfEELc7uW5V
2NpvqV5pabR2fGsqs/nH+fAnIb190BB+nCKN7pK+BZHhYE6TQv/FYebtLQ5Af9Rv0fp9aAjOs23R
70EBKv/Dl2xt9V4cT1+qr37hfj4YOIRpxKIbTPmobkOXiXS0OsuzvsWbqeC8sOpsPEdGKTNIx16c
T2Qvtkr/rFf34C68gxQBuLbKvTov3eMjIVlzoI8KxECvp1Vq8WlJqExilAZ59qnQQPynFxdQx3+G
jGYC8u4bQxGp7fDe2v43vNNSp6Q0/gAdVfFuuGJCO5V8GLWw+hq5QXHSeeRcqj+y/MyKlh0sqQoH
6855FXV0kuLcrzjqLVcnz1hhMLDjZp1UaWfI+UIv+Z5OfZS5o7IoNqUAARXQTlU4d19qBpKGSScM
eBnA4neQ7HHOVu0NG7Hi0049Lv9wD20HTuLutZ653xbuBf/NMjcL1ToJdnvOjnWyhfyw/KjrZhEr
0qExYMz1mtlcYwKaulwgosslKtcULu9cfl97XN6voddcNZRzx4odYKvr5hsxZNjXMnJLXeJAXua8
HaQ2d3PXPnCqg44PVWeM8bRwJzy08cOxt39pBQTyrKfkuN02vcbUuQ==
`protect end_protected
