��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�#���[(i���]������ ������!��`���ݧ�X�B
Ь.��-L�
X��p��!i��Kڈ��?8��zA��)Lќ!e\4���$m���������|�Q�a�OA��=*V���6����
O���C����e�y�WD����>��i$O)�{���-�O��G���t���E���&7H��MwH�|cu좌�б�em$`�q	��؁�y��	�!-���^����m�V�����D:}[�P| ?�j^"@b���@���gF���A�e)>h��c��|����*��а�~a���]cOT���C��a���.���ٟq(\�ʾOt&��4�r&��o����͚��_`b�P�&�1^�/q[�AQ��H���:��9̖Pv(Q������a~Kh1T�o�B�O?�	;�v��q�p��fw��aer���m��&z1�tl<7�"z	���躁�i��a��O|�J�����jO�z#ط�P�K����.$��/��רi2���M���Ѳ���?�Z�(C��K}Yjn4��%{b��9D*�_IH�i�U������@u`��mJ\8����ZkcA�v�����ھ4ܷ��x�����Nu���\�g?�Q!�o}�K�<+�H�`��2o4�Pēu�T�U����j��-i�2~�՟-A=i#��-B����l��a��D���2���������߉a�o����?r�
z�h��MJ��K���MnN%=��gh��ZK:�)-�X�9�(^s��FX���}d^�Z^=M ��� !�N�pPΪ�ip�v���5b�
�mƤL�����ok@�������#0��Q���e-�	��F �r� 0=(�ex��)~�^Igx�8/!�%�Hw�TK��	d��G.�M�Qk�����@[oe�Q�L�(�,�*pi�����bO��JH��ڣ8���5*��)�xzzQ��n&��=[tÓN�(�U��{C����G�QZ�8~�i�w����oAZf�6Ӣ�Udg�����L�A?���'C�8�!)k��s��R�4��8��zm���e������VK��@�n��b��\{T���hڷ��08�	Bߵ�X7]i�/@lQ�Tȯ"�es�4
V(����:�8�m@
�K�����&>ϻ�H�7��2�{����k�l���X�j7�yr��p?kC�ex��M�>`}|5��9�v#.Fp;.��;�3"��H ��da�U�ƨ����Z��V�#�mj\d�m+�3gԥ27* [I*s"a������L\+6f�C����L)=�ނm���8j{��:j=�Z6��[$a��8t�pw�	�]i*y�	zŷ���?���'�D��U'E~9Y�Ff�B!��ɿ�/�1C�`IP�����n��ˢ���Z�Ctv��|cum/�;^����Wt�Gi����~f��HP���+ʍ3�zvyl�����:��[6�v�f�ЛJAm1{�x���������JYɒ���7�&�C��B*���f��_u�`�砑>���-�/�y�NU���k�gaєf:�g�����_(l-X�BV�C3m�]����Ww�o:��g��Mփw�/��6v 	5Q�DE�	Nϻ�}u�9A�0��0�X�糗����c��տ�l�Rr/#���n�͎
XX2k=��\�|�*��8^w22�D}5��'��ϙK������B"�3Eb�x5�Xo	g㕆	�&
,�k>뭈����G���w���{�r��<� ԕ@~�d����U����O>V2եr_Y
�{�_�%U�m�:1q���5�c��#-�S,8�Y��\����m�*��3��Y��R��YK�$� �V�#��}Q�w�5���'b�_tw,�~�E�f*Kz��b��s��g/m�u74��qc�OI�v�ܟ,�;XrW�*����4��]�o��}�Q!�#3����sۘ/����g0
yV��E�~���/3?�yF���7�k�L��z�wQK��$�#ث�ӄcyJ�Q��2u�wP�C��e�>�8������X�m����?�c��{��5 ���H�xƃ����#K���p�����CNҕW�(��DS
�f�@���F�g��(�`��O��H��H�>�И���~��o�c,wR����4�.�x�7L��\Ӵj"9V�j2���I�����f��T��7�NBO���1Px�8"�Zb�l*��e�G����FZ�|ەo��O���C���q[�]v��� �̜.&��?�C�9��{" �s���1Ҕ�Gf�Va�3"�?��riʢ:B��d������cg5��o�`��p�A��!ߦ����G�k��b���s����d��N�����̯7`)�'���2�yt#CY��A����:0OF�a�Rp�Y�S8V��m�MFa�n�T?�Li�-�Yk�<F0�w�e!'$����jXzZ��u �)���.c�-[����KY������|th��u�Ԓo��NRDU;�vc\������4��7�]��oa�˚�l��	c���GB�VЂm��h6��r^���͔-����?��cL�R[�Q���p�]�>���jɰb��+`���W��$�$y}��i���/ߪ�i�o�J��e�?��X-�(�̒�:�lwAE���g��>�Â�i�Q��JyX�g��h�̬��#����]�^�(��9� ny1�8%u8� #QW`��9#� 	Z"�Ds����O��Ou�Xǯ[�̹c�k��%��z���تY��*fFW�{̯��\��؏>��L�9w	R6^8���V��e��t���u�O]�B�^��wѻ�?�~����S|wؕ��_�B��8���Ne����U�8u[�]�(-�����&�'���Qycb�vm�{����H���Q�g��ą�o�0�:l>��H��D�[ �\U��/
d椨?���u��6g��<�r;H�	^s��e�k��3J�D���!��0U��V ���	#,��*%����|��V�� Q�p�^u�o�@�b��;�R��mϕ����C����+��G�S�xX��â؊�O��{z'T�:bκ�kp�������(��r�aZ��
]�'�ԕ5ܐ�e�_�T������e����:UG{aCE�a�pI\;�%ĶQ���u�g�V��u7S��a��"���
g�1�/��/S��d�~�;ӹ����20��T��N��vl�R���5#�w�@t�A�35��Ķ��/�+�qY��."d�u,t�Ö�sz�j���"�s�^]��G�9Ď�>��ʑ�e>���b�:W��9��f[��tb�F�v�����}T�tj���=���!�6
���,�rUY�2'���)���s�qkqov��N%�� �hr��ZlH�Q�<
���$a��n���g�8���4���m��L�;R���U�N���a��1�٧ �?��*{�7��i���N��G�wI�6ux/�L�C����N���W��?��yYz#�l{�f.��{u�*�<Q�C������4H:a,=�_�	?h���X��l����	�������WȮ��	G로m�n
/x� >.�ˌ���x}���Cn
x�O��kDZP���
���@rSRr}��.�E摗�i' 
��y��en�����;(�A!���R�C��s�`�o�'���	i�z��9�h�!۬�c ����b\wl<>R��߁�~|u��5"{X"�`�G(��� �]t%j�AM����m%%��<^a��$%���R���*`�U`='@�>���|��b�Uр�M�X�n���e����)E�	𾲔��`��X�I`hD&�^V?Z{X8��A�VY:Qj$��'����-�'� �G´^��aڕEN�Ф߸���n��:�K(u����X(�Þ}j�w$�&���%g%h3�#��$&K��K'o��@��_8�O�Ľ�4�H��HxXb����"��ۺ����t� x�޶	H��H×�$W�Z��'��f^Ɏ�e�)l�<ָd�8-6����>�@ �i����`V7r-*G��ą_�Ǧ˲���kN�
�����4<�@��(Wqk�^�	�x��0�h
W���w�G�
P܏GAM��7�����E%cW$��J��u%����{媡\5�5�{_�yP(6�}ʺ��:Cn��	5q�F~���h��� H2�<��v�����N�ݭ-I�ok��kC���x[B�zү��FIM�W�c�����H䟚ڏnI�*���2R��,5���L�� q����� ��~X��0�">��pψ�ޠ����$�AB���@�]����������b��84_2�v��3��kQu����UNRN0�[Ű�Q���[|Ϗ�~Y�*汤Z�of���Ff}Hp)@�m��4�qvBzj�
���#@HB���@~�~L��NZ�����[�q�Y���bws�����n�7���ÝT����ŗ\_LR�����W�]�����e�O����Q�R�0��Ȅ��=iW X��' ����X��5�H`��n�/�T��i�����q��8U�r�T��9v�����"'�Ġ�:��H��vk�7O�@�����{�TM1��iԩf׫A��1���!i��jR�zS7���Yb��ڬ��X�G�1�̲�bE�t�Q�;���\�~�E.|
����0?�\���O�7���d8V#��xL��Q�,�q3w�ljӂO!I�s	�|_����A��H�p�OÐ��Y��d�G��U4����@M?�#�S�5���tQ�K���p��?�zhKC����h�}���2���pR:�5��˗�N�a{����5�@uP�?�������-�Ƶ#�^� ��y��S�п(�wv���/,-�Z"�'��EP��L����3���^ނ�Ӂ�3y��