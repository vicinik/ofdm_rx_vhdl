-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XsxE4jL1fEeMmSPxmZN9cgIlL/4urjviIclqnSjDvUImegPBxbO58fbquRRoKpyXalbYV8X18oYn
J9kzXTOx7qOOHtFbPlIyxcHZzjggJcB5uZ5nbdenYnYAZM6fagz5mmp0seLCznqM0N3eq3PmsToW
R8Icqpg39GKBsEj83cM+ScCFicw/g7pnHEI1Sj9plrLOcjlYdDY8+F+mDer3ye/A3Ar1HXKZusAX
NTdeTXDZnVgwHnrQ3E99r/h/sMij1DkntHOOcekaBMdXgJP3jorBDYnnUs7/1oQ89G2R5RI6G7U4
Rypvezt2i3G2bRvGSA32cX8EA2w8uNl9E6oFzA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6224)
`protect data_block
ME6KSTxauuCmeAeRPo9iLg9i2qaw28pd4rSXGaZYzQkxyk+adxIivQu7kMhAnRY1R+OgCKVa5aDk
GhWnsuOrQcKTDiT2qqmabpP7+EhSHYdEcMygK/jcwEkf5enNnUIyEZgKk9ILgCGGqqpXW8nJGt7l
4TdLNQnUBEllE6J8RT6PNANH3O3mzQQMbwT5vcRrB1p/wBgj7AQc+wmW/ZkQO17YWf5YBdAZ0KUp
1w2OtFYL6SyrNduvfTgIH7ckWxGT1dL5YkZLO/xII7riFOV7Ng4S4ZUUS9C4K3ovV5ngVm2NzrlB
LyQlr+xxvGnQ6j/K5uCc4+hUXLRZ047hOYOuT27PmuzCMoihLE0dHXeNtzYocGV9QaO9Hmjof7UL
JHU6VYlFU0vHQKeh1rDjDuycqheAH9cMnGnBoQS5pKT58eJImtre3umEaE0Ow2kmq/FsBh1G3gHC
9oh1dYmTzIyJRPdlbwYFtnvixzjcY7B8TL9eo0wFMWADrgTGFSb3ibLIwIrlv6wx8MRuGLyNB66r
HpCslAKs8MX77iWGsRFSqvKOnv9gbzzhwZdbLU8r2ofOdpIyjbTQDY8qCxKgqJxFFqwfP/3y9jjo
4VYl8gX4AQ0gbXpW92IWCivJgWTz8R1lTf+7iXS76iQZTZSQcJaawvqrUBIHMV5r2SPjaTufikIl
/IUEHAbY2czhRKdHqy8eKS5CXkjinZIsZyBS+FEpT44Xw+FSFMVO71CFVbL7mQAShwwAWsq3OxT8
sZleptYjkmgf2R3NJWDXaRTNckgiq0srVqIfu9BjrGo3H5IKsaFoRv2WO/noB9XMefs/leP5Y7Rc
Wrebu0PUskg8t7i6HL1ZkqYBpi2d/zHvJnhYPlzItPGhQ3poplmxZJjMne3o59eKiwK7OdtTioyl
///lHuBvgqrzkNDznqI5WjnkvrVjCbg2Dv0pajW9d3UZ90NcV3ZmUIN/2n2QHSwIJtHGzUCKFqhz
yCjW6oFpnRcjLkQlXtxizD5QljYv/1vDd6H6rXh2DOGlK5SiZa7MmNHTS+Xe8Uy0h6NSTgGqrZoD
TGcwM0Xr4D3tpMTg5jktPWYZcuu/PKGY6MZWJjpTHmKLfXUCjzoJSwYIvytrvMHcyIBd5hcZF6Wm
jNBrVaKzqzk+3jFMbmuuohiQa57yUCITgD0dm4KKBo+Vly8NUP9SA2cB+7GjDU05sb8ruHLmcoEK
qUiCunDHF6tWB0aMLsa/UkStvCJlSeS3lXl6u1AR/Vw0QztsoZr6q90nIhbaxcjIs+iGwetwGJm4
NUZMAuw1L1BM5F206E8oqjTn1NfMeOW8iXaKys0jktlRh0DMP246QiGLbMCgxHxQi9gbSyRep6nq
/b92UioovNTh8R94xv+rUkS/S3PFA1nXIe9NwqqGgMep6tSAMCneZZ+hP50KR0rWPP5sQQZnPZvh
HqsPpEr2c7ptRYuy+cJeLVDPr/h8kiarywqBtlril6Jc1F1anTihMIcv6OF5YQ4Hlds+oUM5N/xn
8a41bS10ODNamWEuvSRIN1KQ/vRqpyzOMWZ9xxJJqO/uopAxNv9ym8MSb+Y9nMESQmmLxMRv7pCY
eWw4JFJ9aqBFMs5fWedK/CncJdrvAKTbpuBDmqXWV1mIEgbhbKTFtE+ha2T8W95MycCtiMTneF0N
u3gPK6r1SLNvrXxOBNFn85VPZJU4FqwQMZjBp/pfTOBorYv5gx03AQ7eNbmENC6N3S62btncB1EG
9IOeP9wUVeRFSXhrjMdFOcYBNjYLzzYEazo+RYZUmabdz3PwWv4K45rCyMv72W9t7QxGSqezk1bx
duSVFRUhnj2U6ktMe0FWbhkQOYdqfGQoxddgrvMymorPriIhiXIFdf9UzAP1UZeVNNmN4FS4rYif
NKxdp85c7V7ptEKGu9N5AX3qBmKocU/nhaxWSn5jiQ0qxoC4lj7nf8a6Ej/uYX4A4Vyz2tR5jMgo
arIJj2t/SEqyjCqy1JH3QFyxNlSCBUo0jJQmhzJ7WmIRSZqo/mZX4sZWYkjjJ2mUsPkmPAKiobmU
rSR9+56Yf4qwv15xTfqChxcG7FqHe0bF/bMHWaAdabCZLY1vIN/0VVoKVYO/9nzm2ZQtJ+2LA6hC
yXLhobOoNFa2YtqbOiV7bJqpec14ZUcop7WSkUaFy62FAMI8g5fhAU0d3tkRIlfcMG6Rvk2mOv8A
3//bXe+piIIjnhuep+WYDsnMskcEo3uR/p/uRoy5F2HjkbxKhGusE6H2kQbR9VDzlOEzm8F6jrpv
guzHP3DYX6wEejwR95gpmug2XE8ps5ICPevdPrwBKhlIelQz6JD1rewIPGWE9l8T9Nz0cHCvwEnR
5+bxYw5SA8Eft33DeeIbtMM9WQS4xdsSIedEBEAFumld/pvfLVsuaLlv1S2FetKd75qyuIIAngFB
Bqz7sg2ebordjuDJPefDLLn0cGsJ4RjTbJN7mWKV44TDqTTVwTjI7bXsrxYk+nhkHOF7aB/uEG/L
PE1xPbYsAiE1fdicT7g530SnrHpZjN9avsAEUmIVPil72ClgVHTwkHkagNl5l+m3jZuRZsrRJRgq
jJHBx+YyGDcLOBybPy3n6yOuwdN0xQp4uaGDMvPYkkASjjhUjk4VfI1Y6xvBL5ylDodwWUez9rwD
02yF0ZwcnFR9YlfZ4OKGTIM3qNM9xaO7c2b2fIJ2cXaiHSRLJ7vFPvV7ka+OUeMnGEMw+3KKNyko
1EBt6smAlK70sKQIC26oYP/6RboN8mvUpFsMzB9GOZX0v62020WXFQPdKaVVEBlaor5okUNtCxbE
7h42TCWwQn8wXUhH4JAKT3rOX15p+kxm7atCT6kdjHa5wOy5ESrE5bdZw/2S8PMEi9ROXJge143B
9v+i182OT7/WKR9CgjulJ6+F/bOYIypMGtgHxcEPW3/7uYhINM2dB2qe+nQBY61BIqheX/+BauZz
crMLW3LZr87NzvV1QSSklKIBwbPjTTqSahxR0xjv8Kn/6J1aVFRt/9bapUpBGzN34f/nm4QYfXB5
ZfESsqDuUgWb7d3IjQBP0q0SLFi+BzxqgJf1XPbY94AWJ7MN23fhZYT7hfPpRc9f1jkJ7pHdvbpi
q7L8gHCdNkaCgPJixf9SKOJnAbYHDKSjneeZFhMFdaBE0Be6dz7//rNMgo9acEcNuaTAt3safv2y
O/xevfWyrrOAsAQIZI39fqS68/f3+Y6lK1I46+ZOldF2JMtUaJM6ifgapB0nqxPuW714pa62aMoM
VkcXPVCWNrmO5fOpv8K8AOE9iQ9yLR2k6K65wWTq11kKo540saqj+S98Z0z6DFFYsM7PD2wMUzRU
PrG4j6RuAtd3PhQv4pGnv5fojnnd6ew59l70jsVaVJpifH4eNNttD/ebPnmzDdckW0W3OPPAs1AU
mxwJpidRDSx70pB4h8CNZf5mBi6mwUjodlqcWcKXRMl6CpKJWIhty6BCUmZzjNO7ZAhYrJONj2H9
GvQSVngCuWPh69KKii3KU7aBLkWZyERhRaUidBIBWp/TuF47qv0gt5t6kpmhLAaGl9lhvQeeSTiN
1pdmLDQA77MZLS628+2H4yKU13/bW6yfs0wanwPM1BdhxhjpYfljZPI8LA/87xuSL3JtS60ReRsW
36mI+4Go1q/khHrB1lnfcTo7Vmth00ao8vrs/6psqyFksuaR1kkJg4LNUclIpj95pRZ8J5Pn8IcI
5bon7/70fy5X8BHVZxEaGV9Q2tUow59A6ZdYhHKiQYWyPmm2w72KhsPWJK0wvTqjU138oMZFhrTr
JdXYVG+zixzUDj5wFORXOPJSA8+wNDhspBBC3wq/AJUijtJl079IatBHhAGHN+MTUE6RFTWUz1jb
7FK2r/2qwOeJurqLfQceAhbJmUPnU8Y7zs6yjtqwtY300tl0b+w3L9NC1mfWorkXmmE+tRxbwgKz
yA68+kJ7JUrAAF5mkRRHwV9ev2SLaj5y2pSLcTMJR1nj+anoln0mVmZpuRefmEu6scBnoIBNEYY2
b5819x3yVC2UJOv2Bvdb4Wzt6gSps52O1ozLqfKEZ+9995YVpE9ZCNHNqsydD/IA7ZG6SEfgDCzs
MTnHHxepUpJ8mZawl7FMyVWpQOD03QNd9RbRqmw+KuQNk+YRPRtvH4/3ITewAYEcEOs2bYCmif4g
DpLu53RkWJsx9i8i6QPnHfZzh5IDYNEGpX7cyoIiTDAYW8Zabo/nRb1xivsKXk+ggA0Gt0bD5mFQ
RoLtUph6j4FVsR2oxN1d3SPV6jvjfriEpi1h0t2O1150cCsRvGOgvnBdzg9h9JIExExRKhcG4Ecr
Zxrbs2rLs2WrT1wFdLrjS/d7dVASWMqmZBzV/9VQJBKcFs6O+Lg4/M8x1LGzAq/BYFWTBcYmcoBE
g6WvFsr8GqsBBs6FenPkbNUlcYVrn59Wu0RxSlUKLxa47/VWxI4llhmiLbrT2B5NO9oBa3UbXiK5
/tfpf9HRj0eyzpNwolO7FCSyOMZi5dUAF5b1sSDEYhxzwh0a6j3gmriVIZx5TLm6T4SDY4mDGcEh
aTDOXiukh8A6MSAazAgxaha630Juy275MRmWNbjN2O4/zaHzJ4NWHh96BbSeKqnWJ3J1SZ8EQ6s1
X2EeZFUJbqCNyY2in1DFvWU6tYUio0QhOa1kMbq1cwmj7Xu+qxyJGB+i+wHWDeZH3iLu338QAEyK
OJcSbYTBlJ63k7770+a2KcVj27O+RdenJhB3pJiKvEKDfYn3P1Ft2LImixrZWRl/5qsQzly23hBV
n5F9IyJQWAkp4CbpwZt8DKI1kZmmvNP6FDfBpiRX85j9UftGMwaPTfVmPF+BoWQVmPt77Vnn7psA
wn4dPRyu09LZHR5DyXCOZUli9RkXf/AJfpRUD3y3JvVaYHZ+gtihS1XpGmQ9YoK5qz6qr2HYUWhS
/Lxojt6PwmFr+d/LHcBjCEvQMq7XUmDb6IRgJ7env5AQn+dAYHoqqq1anruijU6dvC38aKtWw/iQ
f3KRhQ/wTE/fSda9arS3wTCQhPSjgCe6YCKDxBesQx84guKALPowgzeg4cfkaz1MAjPFbkdabt82
jHemn0tAqDYV+TtOrYLSHIL11JtcT1d0isHsFFzi+3PKoZWUlkUKMLODYHg3r3En8LmpgmkwIE7j
7ljjHG9uELNJLfpHCa9w0gvee4w7QZt1WrqQbbgjmDymrfsp4tzbKfBm7HZ+tlercVFU5B5sQnP+
UI5nwGfcpMHu7H/7DxoQZuKseCgaY40YQPB+EcY6v2QmChJDsAkWX1HoYdAwPRo0I63MIOIabNdz
JvJjHoOgOJbeK6weuGh9deeUt04LTYd/IG2+rt11DTnAGC8a/A1oLug3l3uSupyAuO7K/c4D9Ac6
XmdN8eUTmYLMyhjvdsrmdZNwkVRhcNTHSkZzOwX8dWNVlXY6OiG+xzCMY7d74VZwtwt4a6FKKcqW
mWEkQy13fjpgMj4JOxipATTsmBkTcdLI+TtNH/7CmOmDBgm/tF4dMDWFaUdDOWJGkzRfwUL/NxJr
benZAalG/GW71sJEBw5HOSmDW0bFHmPwLR+OSCJ88NVF4bJZBGni003Nqog2UBUyxBJpHwYH8nYP
jW5gItBy8XHLiThYJGqTliAlrGR2mLFdCS/z82AaZwmfEu4MitcN0WPeS7dkTld8MmfyaKQ60KsG
E5gDbCEhRA9v0E6+R7KJrEBBuJUT8SoUuR0ceZnHD8N0q1i8MyVlOE5FSnOscd8RdzTLwMVdg/Y1
rZtWA/EStaFQk3TnFbEJ4tzx2/IMW5GM7X7lcIIx0TQkylZH0hqDTdgQJdkHb+w4RfWsbeJoMhsX
/FEpoZCMVzHh2uNNuasFEkqVXgDYRddnPJ0+bfGhSEUUsUnETE3NG3hs3WHnA9pnbugEcrECb55z
NbbDisw+fWUa27MgKsG4y3bWy4I+y19AlRTbhalYHlxxHJ9r1r1R9MB/BPTirk3hBV0Lq8VIupPT
Mq2Re99Vk1DEfN7bl3w0bQGpnTffb7GKvhuDuwov6c55ZmlhfvMjAp+BC/5Prb/fLG5Rr44E5eMg
3geZJ1UfuXWyVoUuuNPRtjIgSzoLWkTYwhzIg8nu9R5RDOEZc6cOBMtCIx5QVUSRfRUB5G4LO3We
W5bEk1QE7s5H7dm+taqT/iQHDdGzXojFCr9Go1vHYMSIbTuBdw8chuHW8VsqzgkI8yo+f9Rt5gJE
NuLea2l+c8tVLHobpyK9kG09zmPCZw4EpYz854rrZ+nUnHZT30AMB50viO2AKO656HpcnIYSjTca
nM8bpp9wz8JfmzaoEPKI6F/XBpjttNlUT5xq3irVw4iH5QWjIVxoRIYDhYsZeXxWbLUKQLfeqN3H
WZ+DCERWe5hoX7Vwp4vhSexKXWft88/LYyFBiSfiz8D0NCqDvmo0K7Y+sw9kxD3VGHvdKuD9eRwl
rGGyKbpT+igM+4517epYzwgICAJ9XdZBOpW/MUMWXVxWwrRUe3Id6+rQ8msHUMTBscdr8QBRW3qP
KVixeG+MWS2gZu9TM+/mHzBceAcSRjh/cLeb+aiVz4oQlF8JzSu6aPRhBjLjvk6LYn0zoDbM1yN5
NPmk4R3bcAAYuXoVmZIRB99hr0Hpwq3ao9B1RO3mvTTjbWf75fvzffyMcfgpdXFHBqwmzRY2ucIp
mZqhFiGC78OkOF9xtc0OLrC6xzPTG3LPkReNF608sXHoq8A+FMNJKvfYwJ0KZ3xoaZEYyVvH3pIe
nZSh3FOPPoQEyzYeK0RZlKKfTib7WIy55QiChKBTnDuCHd7p9o0WXWqpdO0jMiBy72ic+iVjBnKn
xmkfJBB/yLTigJJ5NJ36RS38ARBl+O3tMABChodbQA6xDdnNxnisa5BgEHGg3j5//XN/lWBjK5cC
ZyxCHk4zcabma/9QlvpOt9Xuyy0ydyg7MueQD9teWCu+nWWk8hEwyEXNA5aRcLtN/kiMS5R47SRd
JXTugsN99TPvdy9dLQIOXKlp7lJv16JdBTnjMFf5EC4ntCBHB9Ew0aism0T9IIogNv3k5KmEszDV
F2pcV/iMeNZ+DCFxrIKCxXV13P7yrwU9sOV2c4IUTyhIOBLaHlW9PrD2RN26iQ1CDbsa5fVDGj9M
QrmqXix0CmvM7UubVb7ceRxadY4g3mGq1uiXFabGmhmcPtP0uSgftFOaXx5CaTdG642AXN4vD0en
3x1bAZR8E0OYaeHDmy5Y0ZPWSDcPkP1APjIHGRZeqxPISiH8xmo4cvTUbXnsWZaPOpEvxQbMwU6E
PpzMio3Gv4ew01SHvl70RnMVRa1nZMSXV181bt0KfK+8cUPdP1geGgw0ZawsSfd8oLGTRwnOEriU
cAwJbN8EZjn+V8mLlRmYbLfFhb2n5BQbcQcxet8EJJUA3V/zao8Hl6qVpXk+XQS0QIziRPcPMG/3
AQDgoRW9SALcfhp0lDJWDHhcraf/IBXE1k5PYc64zR+7tzmDN+YyCa4yFNkal9WkZ7/54o9uwCbM
Ru39UoDl1zoDNBaeN3KlKVkYleX7H9/tO93GJmKejvsOrLhv5vz0B706JD9o9Uz3Ln1Azlw71d9s
QqbgUv9yI7aKqJ+ITPdafp650ITa0nJEvHJkezKbW0BInaU+o1u3FjvUF1+OTJT11Hm5SnTG6ZSx
4OKrz8MwzyN9mp5E+F06yy40mewXpk+q06ZBRNes3BuZ3hhxWWk2z5wwdL56etF9CP9DdtXJtpfm
lvqI2xLY/T62Ulwv0BSPhvYEdD6RanHqcvjB5uO+pk+HrgVgvfHPpqEEPTEDkStwAWcYeMJNVpv8
zgwdB+gb2UnecrAO0DnEoW3Ej07aYOLu+01tZ6NoxUcDtEkReokeuzahTBld0BhbJrFMUMT0ltcF
VjqbYhHrqdQhosxJRSf7FBLLLqixgZGSyjsgzWlGhI4NxXMS0pePX1dnGtWe1GnWyZ1j/12DlV7q
6GfC5hYueA2xbeY7Xhx5H6Be9VVOtxP4+DhZl5WBjZXuaNwKWOFi4ZrpnN8hS8c6pdu26T6BUFRC
Rns9VHd3qd3di21kgs8gE8kl86jI+e86+7vhYY/hydlZemAXROKyOVk2GJeR9l4IXJZb9/VsV4uj
vSe5ptvpaDCxBS8m54QMzlY95Hc603flGS6W/zR3l0QTO6FY6kkW5r26f/mMQL1YBFLHP6ZwO67T
lhDpHMqaAZwRKjjiuhZ42VaX813jlPp+Fh+OW1kyi9TINo+BG9Y/hya8//q13fmfk10sgZixJjWO
xgJPIyhgJMMTq0I=
`protect end_protected
