-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S1YA1oOgKp8vm7+StNKbL03tTbSbYrbNgORAH+iexYUKpCfPKdHpDoW4DW0mbgnroaH8YPMFaz7A
r0PoaZTrP0AtqQ+2MwIHwUZWtEzZZfz8v5+3ucMZCQiwG9O5vuoKGafCXqPWrbtTRfQ17RIOx7vV
2XoChIMQWAJgBVNDZuKMmU+UZ9Lf5pSdTnAXuG6p7CD4wnwdBzelBSWLef8us3Ld6JvQ2Jj/5tlN
Vvk3mXgoXjO5oEbsKdsgvACsFgLwkQXZBGusXORZ6y/y4rcFrVk9wUHBJCuGHNQzP29iHNc/iLT5
UqIcBl+pD0/OFjOAv/htdJWeYE+1LryiAa2hZQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9424)
`protect data_block
dq/K1TQz8VIB4qbOymFvEfRk1zQmmVjyICncFUYLDrze6ERR59UxPbEJFJ2qsMhJWKcf4eUm1oci
mCDNqCXTsxiqm5eGEORCcSyl7t8cN7mdJGe3TEkkSC0Bk3Ltt7/UYV/sFTLwd4Rd/Vy8GVXfT3aB
duLbWJd9cCu/e/g+kdoXO8Uac/AX2yb1kcT6XwwL23WXI3CaZv+8EQoIwinVYiQ+zaGPb8lVzSzC
naJK5eN7eHbidKqyo6w3ZpsAmD8ziBjTj0wfZpQna8+9DQ8aulYYQl6fWX62h5cDymvpBlteRY86
BpeIU1lEpLpq6qln4tMSA0XJrb++qIKg2SQEEca47570xa/mVxUYg57lMMxQ0IuqQAQI6l/8bMMZ
eO8MCs2hrWEU8gdyvQbY+jzqLUQZyOQHxO4v4i1FNpATkxsy7OqZxNqhyp+dMB1yp0vz4Lkggtdn
xndvIAKh0A6l4W7oVHaUFwiWtNRLeqo5KkTgg7wqpRqK1hL2k6R2J1cMuTIbDUBUTJs28D1hFIe1
DgZ3Apq3UokVhvsF2vmaNTWjOEiV15OgObxQ2KEPdsvLA/unvQJnmb/ClZajIq2mr7C8PztthU4d
TEaFGBbWJKwYcRc+jzqk61iuodM2TMWbJltABoe+CWBw7HvnY+v98j7BfKjwn1UuTjxpJqmoI13D
ew1h4YP+fJ2ugV7W5Ccg5AwjdvwIWwpYWGm2WkeDnDKGfnwj55djaUvQfrTPXAh1TlXb9flVevT6
hmSj19lnRme7OZRCJdRZLcDs+iyqJVoFrJzOv4tIkFByYSDunFRuNM4TYqJhdpQBuv5nOlUIlQKS
Ztwc1FP9cr5dXD9CVBoSqS0DtNXh3AJbGobCqRdBTND9oYjbra8RhFU/3Y53zqWQFuv4G5fK9hso
6ZYIK9NIT3XS07SmuHPF5WmXxO50XtVaCev4mOWPatDp/CRcbh5xtiEsI4np62mPW+Toq94mGqcz
6osQNNwc88EBnvamnob57SNeCuOuyPm+H6YPzKX/peJjreUWp317v6A28dzLXuGSV/M3I6PrZTFZ
K/l67lDSSfxbZ6u/ES+a+qCKPASeUhHshtATB/iYeyX3AJkdO4D1lvE9ZHNN/cYe61K3HEBd3W/4
+APzG/npcwHHN8t0qj7RAQpLqEvQr25XmmHMTIjduEAgvHOkB0VxmKopzCxQMP5c+58aHXvGznC3
JY0/8k/271xbwS3nas58bGY4Xd2pBs2uXWl54IQOy4leQE5ueqyYWgzdR5uXSCL7YtoO0Z3ovCz0
Zovk53gqPhHDc+0qDDEK1657H7FMWTr8HWwqPNWlAx2aQ/cTA+CGU1+63CO3Dvwl8SYc7kGH7IaM
xK5RvVrDIqdn8jVn1eM14dxXlgeAUfjj9ACQX5hO3xwyWV93Y3FV2bCkyLKehZmDfAVvQrdwUBkK
jIMxAJTGXO4qs8nuDrRvTt5QOdKQg6kojKJxtI0VusRPalWdoaVXAeaYwixEr1Ol7pr7ZJ75xf0G
C2BLZin5SU8f/MESn/WTCixBTFxTi5c8Nm/FJmJaqTWSlGZEGXpuWrcRjk4KNKTzNPtjlcaWU7HW
OoBXg48zUcZiOFUI8i9+eehxxZni3BZ7vf1yFl2xL7UXQvgrBXF3qL5bY0JK3LWrwRV70bIH6Vz/
Jj5lwkiedrSLFwS5E3Zt8FcfEuWaCHuQ0lpfRdHsll0Q4xymrmWJZhoH1R68rhm+7O2QLTjhFjXz
128XmCviPTMzXtkxl1gyVHu1Cc/X2dnKjM97mslOJAUEoZuw84G5ljlJwZePsTZ29q1CoROJVn/X
dBgx6EKtkoXUGpo+5cM9IZjt/5DWW/GfLQUO1R7OuKCYz84ldZF1BJq+vOyIGBhAyIeMCdOODAD+
RE4i8bMsmLIGkMGU7aObwD6ezEd+bcLnrK3ri51i5ny3GyZROOAhDYrm3rE4x9UdhI97mGWLcbNa
MDsdgclZpd9UgPyCvuI9YXwaZQ3pyqAB29iSn2SGm7uB4TTRWphivFtgWLLWKLcZ853asxpyTvz0
fFnhEFWq5YLgrAYQT7rtDGfppIdpNtq7UFNFmeuYhtcjVZDP0+8PPaKQ3MnAAXcr3Seh7JjiLoQd
pBM8uU7UH+L3mWhAkpAx/1Ty54WlQ4/gMuY0GLqoHJm9tikn5DhwTQAzG+UWBfxXQkCXuFLyqOOx
kfFkO8et792tWqNzb/I8QPCpyc4IQ/MrNg77V8itYF5Dds+Rkug5fckjX+ebQaOg3GLjqATSdvR1
DKuYRyXxniDUPQstpYwaYvvQ/bhQJyiIFWVlGy30IPWL15VdAwd2kzsXYZMvCu891udfCaId6Ugx
6Q8k+qOmx4riM29F+TNy/4MDFBoe/PS2viFKw1lgG48KWrqoVPkis8a9ePVXCAna+kip5jFh1U4M
25iypCTOibIyK8jTOwYWIF15P8+8kSwOoFFTQRIw8VV/3dAPogNIRXYS1lFGGnW0JNSJCvEt5Nb5
JFM9vBcJVOqxrF8/KaoPYrb2Ut/0tO8h8kEx/hCNm/ZwyVSjF11t8ZeG65r8mIfWZ/URfc3eqPEf
eNTg9xzfXnr38y4DFamnMHs2gbzhjnfdkBPCND51/spwzG9OeiXeYSQ+TIWLlHZhIm5IhQMzSAWw
z7ncAp6OfyLL2W39lJ7x6WtESJvqOjzdjtdnMjbtx0fnLhrsBYSuK5Rit4/ym0J+daPUD7m403r7
JUs8yTL7nQuZUn7kp6R75876yjFFTWJ3vcatd1HqYuoss8nzVynzrRi4q5ONXNy6I0nzZ2DljNSo
AkN3O9n9XXIUpeJuGjlnD5qAMQqYn9jtcdOD3MLUVYPvwg6wRKL87gxMD4py3jkbzq/Dv0Daxx6H
pmEeKvinYnaLxEs9k9vvf+HF1iQiw+XyyGrPSME2j1n9UOfW03JFq4s7OdlXtNPaZWh49I48Zyf9
l3ockjpRz9Km8OH9Vwc37JS9/OR+Rt6HEREq+hYfaDypbF7xsh/yjumQA3OgbHx4Oq0y0nrwd0dD
Sba3I/zpROuET6ct+5BaPuwKtv/s3xoOUI85mqYlbWXWdYhLw3LS2NP9KYW7KO7OGTN1Z4ud2Q7b
Zz5xX2A7ThI18IdHr+GzqfUgR4MHEaArwjB4kVF2RQgZxfp75+67oY8zGQhYBjNiqWvlJ022DLpQ
vZ0z8ENL5TfIXqyg361vb+qGthrUG4+x3Uks8NJcTTinHEwrPDweaHGyGnkof98yKdOLRX3XO7WL
YJj1zW0kFtMUjtWSHVACYbGZ9M0IuBM9vaNsN2tcbnam2g1oVewHdQd4ogQgvuSEBqP56Crqxb8D
NZPOXoTlRpCuVf2Zp3GnEncHhs321ZJAOkfZAo6rCpf3Ya8agzDJ488HM/zz95/MNNTCDxmk3mCf
dMxrs56Duqcwpp+ub19+5b9crXCGX0wd/fhTFTzhrHi0FqkTmZnnA5ytcKuD5tHvSvj8s7fUTqJE
fQDrqO1aFIJ+UZlSnnXqw5QtHA0iy5V3oEbte7zf6kdImjRWmTxwvvIbx13MA7nefTi5Cd6qYZ9l
hSU9rmZVhFTIFgMOQPW9Z+qgmhbpFdcwTOdpqLVsHXMA/zNKLOiQN0t03chq6ICMEGCo5WBAkf+7
AT7W/321iVcIvagNDNBDw8TbqJtp7ChsnL6XDOx54z1VS60CGEtZyh96zySNXJ2dnKr2/Ztw8Rqu
ut7KllA5bafkYZIG+cQyVXyJG0WxrOpYV9zo97TAf/vqBnqWmB/djyAp7xPi+coJCs0an/N0kffP
QWqRe+tFwM7IKJEzQgtOGnDETIpJrvUufa4hR/jyCPWvEu5jNqURfGbn91CqgXqzGLwwWYtVVur1
HerhCcTT8VrghWSbnefPOoFTGkTgCQeClflrBlKCjHhaX9d+CTw5NTDMKssEUXpV6q1rhC0V42aN
xtMzVkYI11osPCJf7wR2+G/nvajaIuFRsBJw6hoclgpGclskaOd5AazGRGKyJLhhrPifJ04OzoY4
RSoC3JIQ7XredwQxqDaxWfKaTszp+ylVf7qQNp+SPNw1F0+Ywx07h+E0fulB4S3Md9iUfa/P5A5T
HaT/MoF4hhVvvepE8KvYaZfx3ZHnOHkHxJN0xgLXCGic/6HqDsD3vWA4ah5mrhlnIzfOcwmntcE2
Ok9M3k74OziEH43r1tzl9X0ypFOVmXEED5R0h/PvFbwR2pfZDyDebEyi0ooQh4xNwqwZpON8gHek
pjWLnGgzuJp8+0geO9hrpnS8WZu+xhQAsY5cJ7RQFnTDST6KBRf9C9ShpJqe8NJ/i9kBs8fEG9fq
Co6sg85SDa75u8Khh4qIuEObP/jK4Un5O3v8j2gpC4HLKZj6zSOkPJog+nUYYgEbXV+pF9Xln7iA
HI8EJtHOGuKwfvLPg+pFExe3PPZmT8kHijLrOo5yXOOCxJ/24hDwq4sQpQA6EjbCLrhL/XRsDRgS
Yty0xxQRGn2yMaNyWz/ooy7Zp8WnL34qzNIqQLq0LtG6WPSlWTnsl6+tL6O2SmL27rwYZyfFnEU3
MDcy2hDkJquaWh5if2KWYg4R9TAb6vN3CaAHIv4EhNIV7QDlLlowgA2TCT83Olh8nRAoWVc3wtuB
/UbCrxRscQNHGGkl4uMiDmh9Y+uY3w+99TC5SLxzykIIYeXBs2I94fv+x3rQsKfHAl51V0ADfw93
ltxQx7iQUrsUWnikZNmPHZTGh6Fwl0/+2cJ9QVM+JpyD6Hxhk3FdPfoWDWdD+inmOu8cpNSJVWFR
tPanCc32sG4QLFH5PwZ5lmNzqgWa2kLNkWWEcSN1hp40+za/R1OarZeyDbbPBKkz8DfMHIf7x82K
XCzo1JR1uyWTfkQd8nb+jLlUqQQ499rCr8t0WhYjcAcXux9hOJUJx2v018R27Ibuq6LRU5Sv1QTs
UIOP98WY2IvFgArCoRkNTryym7T0TWeGw8Qf3lTy9eOC2a+x96X1+QoADlIF9SoIuK2ot3CvuHBj
aVHZBgWoL1rzJOetXOQouinHkWtUErEHNenWEg4RlKJTTTjasVvBxb2uKF3ypBDWxvIDXtzxO3jA
C9TgM6qpiz+/kCAEjHw0D7FhjV5waOsiSn/FfSYuGw3XgDAQHt33rdw/gx6DxTt8d/gQjNlvLez7
beP+9s1lXWofRBaeAipp57WppAJz+BUhGgPpu8Ep+vbqMpty83VRtLpe6aoBV7I1afDcO3HH8QLr
yqJKAnAitRcqj6iDehe2jauTTUdZ5mMDSLvNCLnSXj7ySZB5K7uRa8thDhakiX9tHCy2iEt+eOwY
7sde7h3gl3Vxa+NJZTmJHqO0GZMLMCjMa1si+mtz8gFg3f0kC2sEYb/qI2qGVSKLJ/IVpDf5Ubiv
wLE4LwpBpZw0YffKznk49cg8sO8CGSYc8tuTe8HfFhoR1PDYGKvvfXR5Wk2UKHtM4J2r4TeMR/E4
GM4Zzv02QFzqvQmg/HXzErR7cZ8hGRSSPp73mhZvLsmXqT2do6w6TChLidlOcMsrJc/w047Nq1QM
JFi5mIW9jOWxCTYqFRrhpJRuU+rLnsqG/U6WbHiEI+Xc5dbk4Sdg7Jng7seHifphMq20aZ8tB3+T
r9GDaUY6Hg8hrTbU/+WnKw4kgYdK1J0YWf4HZrO9q9m6G4i4QO6T/df6DmoWGLEjjJHGac4QENUv
/TAanbghb0QuoLjBgE0fYRM8shMNbHTzY56ZNlG7tHFRPKNmmZbtyG4TF7Tdnbp85XslwuWz0Cbw
00J5M48rNRgzCeAE6iaAmyUI4ykwu1VOzbc2NcDc8f5QR8zrMNZVfPQlneU6B4ZMS84COdeqXwN/
LgrAjz4wtoR1erfJ7HZb6zDftXJIqfqxyQaxoxzDYHyw0LVYTNruTk7oEI3Ze6KKfConJB46aqsU
DaajH5U9zze9/QFhn3xeZWkygFomTA+SAwzfVs8eQa9cW9GVoOQ308WIUNMLMNi5FYhQuJiPOFIV
H9afNHmOpbtZIdMovylGKbQfsu4jK61WQYIO5c5n5hekOmmTxU/sgcu4OfgTtPPPnFN+b/l8UtIa
xdsuoi0siWTxhWvzu3qW15POcVc3UDn62Mq8jhRtrbpQ/FyFhJVRMxbn1/mKD0JcKwTUicB5U3t9
nbDADD4Pz1Rl/lt8VqHuvyWDo4XHjhQGvGsMbAnbvqZhszGvoDTl8fhbRbkrN+Y1AmGG3UKn0Cs5
zrf6MJ8736PzcHURI98Apf619Se5rBGzAvCzTaQ7xj16n27SE3AOl16/3I2ROlNWPH4904wcxIja
1N4GtW3gtg+JKvIqIwxn1HbAWHomASDxiArPIog+FlbCRGAc8QmzzncTqhsg+1ClVZdyXTgGfPSL
zt7VKXqML12QJcrn1nkZtautVUkvu7R53llblHaKE9k1tqAIyiJSo/mdkhdcg5B0+4z1L9BxipAL
2n26DgUJMZz7fzHGvBxYoQIV9i2tZJCZ3oat44keGG6YusrU5aju1+st0SncE6w3kncngt7CQXHq
TpzFUs/U2+Yo0nDYdQcmsdKZgxTnuCNcSARTZGjR9O+sDWYtigsKlK6hljzxFbE1WQhZsWa6GRW0
OWsw6tnqDLYBz08/+M2llCrPstGWRs9bMF5YjTxx6oHNGIadMNDzWxQyWC2X0HkBspJohKyiWQXP
AUAXrWWg0kzh1EvSbAgzEZ1GUbQ9/tQKbG7MEZK1QvxIPYt5nhiWPMYjhwsYqKnEzt6SWTCaDwE1
VCnqnmbp62jCzeRXK8nVhlN7ouvCyRo2RDx4Zjw+wi37UBg/9p4bQtwDCr10k4NYnbzPKBaBd7nB
ytIYoQqG2/DflMxvF9qXePOBgoeIP3eS+r4uraHOOILBjD6RIZCkI/oOEfG+yxXjDtPbGwtviAXM
Gg3Yex03mJE5xZkaZJ54a/UrRrYHlcN2K0cAKlFco1UUQ2GpgSlSSORB+Vyh6NWwMb34r2ZvK4dr
iU78iBoDPOw5TjUfM7RA4ccjLBy1Qg1n1UOE3wjGHyJ/frg9/S8qCeQL+9buNw7ebT5RHtYD6YUi
78OGCBLM5dY9BpQFe2MsJZqoVR10DF2NBIk4ZXGfDnDjM99U7uD5hL+YnnGWFLwZeAtE3eBkXHeW
aOaa73BZ0LAm4EJt0hjZ6sL119A4/j7wFdL22LSQSoonfJMxK7KCPFR2E5NU8kX0Hx0psg4YRMrI
oYtzDAeYHv/B88mQNwzJRUXiS+Nlp763oiIZAxziwlNKB04t9dsaP+APQu6ZQBMlYKI87h195qdX
jvIzH+Lw7ndCruDKbAapZeGwMTzCqdyy0WLV3P2GqMJy571BIIGEvowNYDFduIiO+2eVHdXXkEUP
hj/cRtBXaJYJZKd2XcPvRdzKaqdDn6LgCKrGeVN1IcYh4L4OyDvkv4v/XIyVjy54YYus5JotRRVU
kE1SksvD074a4WO4u08HEaFWM+PyrVF61PJo5duW+7Emet7E+2JFLlNk/Guzto+8RK5Sdi+doP/d
KkLzgjWUYed+sxyWnUzRmdLaGlWLfk2e0WOi4sebavllKLyaSpWta5obPdzqWUxZMMAQTYsPuU1w
ivGsQh6HempONnViXnNaZqyVuEmOm7eV+VrZiEfCyXQZI4UTRsj5mXOHH665Fbb4YeyF8lhs67OV
ojs/mvIKmgPAyT4v0jvMyQRQU9rN8qciT0al+H0719EwngHSU+cDDPIZ9AG5rgPic2cZuoVz7xGE
/0AhOp1THvnU8m5IJJDmuawKJ0vW1QQJjWhXHtsamQqC0BmcPohjHA9Ec/jcJCzPHSO2XcT4/0mn
IsRnl3ZkwYFhqr5jwji8HddOlvPVA+7JclIcq99YSff2zFv96CafQbkRDfWxD31Xdh4tC0ETk6uN
CZz45OkHw9aGvh0jZO9VryfSjFqf/u9+oXG/YjCaXjOPT9WqswrnqIdxGFEOCAn/W/ARzFTMDbxz
DfHg88ZTaygAo+B14pVgZ9pdFfFWZQX7N4MHpHnAGwHKsKfF5nVYPk7yMQ0KfyUdJ6lbEjrkUlgx
B1NBH/Fp56PtmaFKfU8qnYxX3r8YfjkTX9uadgkokKTTHCRRd3M166gbWNr5k1ZCNI2Te7+Wu7za
aDE2HXiuar+9Tl+rYZmxtFl4c/Xfb0T+HWG4RNY9jnFyyAqfU7ue1t31tr9H+Tg1KsuOG9eDdeC9
4MFfkBuAq/mKpNIixjnCurkw3wSKNHE6pD2Lv9s8RTKoftGKDEcISr4o7MWX/YPJrwvok43dM/UY
g+15YHut3B0USZ0GABuKdI5yMk9u65QWcL5+1MDbmOWvWWC0hd3Yg8GbxbiNLrF9qZKjKDTkT1pR
E5vtNn66UPb3ZOhw2+pfxYVd1Cn1LGe3NMN8mbSRFA4xhGAd+/BMjwXIU4AmO4/7Y0SfnzDCjIxJ
3WAVeDrcgGQf4qz5QE9Zgejr20IU/YR8u50xRN+Fg1MCbLd/wKgKWfIB4eYiKRRZpscjjQv6mMU/
lmhLYEBW3TkBOR8se+ug4iF+JjOyGSmgszDs6fF8cqUpzKRqy0obLY7yhNZcPFbe+mY6B2NHSjcH
NOLw8HJidzB3n2itAaprN3IOpQw5lqfxuMMikC3j2J9FtqKrHFbOuEn738NuauH1mPhmivROeXal
3KiZN6/OXVG3Gcg9ippaXHmKEUab0563pQX4Hdqbu9HWWnLEewAuoDnYsRuhF8My73Eiy/5EakI4
dOleX8pcRPewH4wwB/Ch/P0e3U/rv6HJ0W2o8/JgeebYPGtQfiRGfADAQVHUB0+mk2dkOtTRunk/
dskFrKmULm5KdpRhkkvTJRkNCCj5G6g/NsQxIhNaitOoWOiGAc45oey8bKInLOGVyCA73Cig2CrP
d5xHxs7sO4IAuY78+G72D+UCW7eBIx+hoGrOj3UdrloJ8EKKyh74d8DCpoiVER2pUPSuaXHKBzwH
QYreXkbJKqjQebeWh6WeQavaZAsQdRJ1/OM44gj/IegryMqkTWDu9LgsfKy6FufYStj+uqZb/TE7
FV9LHmjJ+cAwi1Tg0x5r83cRGGGBvNcBZiVhhUt0tvSYN0wrUiBkV3OM3F/Vq2mkITFP3hVQa/Te
hybGU/CB19KC2vdn/BJM1IUbiEeQb3668u6gsPL6rJOaRPLa33J9lPnduWujTlwq10c+kRuyg7nh
LmDj9tHXRyspgeTGDXblgp/bZxb4MF4VCy6wuntoS4/zy4Qbu1o0d4rNmwF4fETwQV0lIKzHfmgr
m7vemDWMvVkYkiqoRMQtkT1VRbuTV9Nl/mqO32W4KY2ha0PVnHyHKsDR1EIMQmxQcbcyyCKRdNMc
fdeAJ/bErBILXecXOpT84bJxJ4XhkY4NJdAVqIeirWbxliBDHZNmWlyvzLZltos+Uh1kYDRL2vM1
an33ZiYiCMtqWVu2qH9nScUSI8uNhNdVKm0uAGfVwAPjUFRfWjftwoKIKLbfwF1zTrHid+3SkIQe
f0ap6vur2HZRKq2979MD9Wzw4IHs1U4s5d31jEQyNyFMK4eIAGiQ20WW2TndrDwWGPwzEpQXaErJ
U9+D0rTJg+FX4rFSrCRoE0x0kAJ1ACL33uSOIlUhAErOz+OH//ZY5RBM7tUUzvyX3OcD3D/v1Fy0
LgGiuhkBU+/nIpJrFaOXPRCDs3HiP4XASKEkFLlNMWlIHj1tKQ8r1ca4E0EGwCIGWylkhM53DFZ6
K3NoHGxE0H8mQd9KXC9A8SoA7GgLOXXfb/bpc9S+ERvoplmAepiHi7pRsLkZt2q/hucaGW2NhwkE
AIPeJ7JpaaGis8h/jCq3YQAt5DX9/87wDsAQ0dgvXOdXlP+2P4RGh5IgexSCkt3tpftOc7v70DZm
aFlKWwQA+rVT0HhYwn40IcXo7rGED/x90bF4efX5l5B9+Pm0mpXVkYFJKPHogKCPHvVBKGnKSuvr
Px225PHDnqJZNOiH9tYJuTWHBvAUEcrRL/I4/qrm/luVCCqiuHI6nPK0CMxSY/PzerDCoRPi6OwE
HHHOmmGG/f2J94VvSbvS3+iiu6jM/uicN8qaG1ApQZtBQ1kBZ3SLXgW2YVNhPz8dIYprOebvNjZD
z5K69hLlyPq22YoqgF4ZS91cwR5QDoVFfj0mrEBS1w4jYap1hVfQQ58BfZRs1rIQix1WDwx2xm7r
6Y59TnaIBNWtrpJqz1fUsRDYzpJqXeCVTfbpJTCY9YX9DgkeXO5zOJAfXg0xPWU93pdHD6Xn7Qlm
QBJoaO1ewJ2+igKBSQN9crtZNDm902y2nB3pAquIQ/Vb4pLw1xhb+OzhlNkPo2XFW4vZKUrsrds4
oxulGlVj+W2/7gWNZQZ4FPsT4XHXPyDpUTgnAm50wTIHnZUTYzeEKlauIBp9rhq8Nee/st8+NLlf
zcPLlOziseAGq0ElWgNQPE11LgEMcaRiN+mfm7JIM/EPIrSY6cN3odvDG8JE38KvSfklzy1nTzur
7IY8CSZW3ZJVJk+dMiFpSTPy/l0GGzPP+GsR6gSjc3tFZfY+l8ApBiKtNCd1RtflLZFJxecQVpr4
KscxqxPO7GuO01IhRiyv65fL9DUwZ22e3HHXQvJmvEHp6FF2b8DJDk0IRPic8FY0fm6xbyIQuAPN
jEilRTZyievlazgcyohcKUU0wBQEJ5SNA96wDKzgrSRezz10UzxjwGfCw4SB6svJEEc/P57vqJa3
g5EPwaNTaMYbOA6YzDiG734aOKUvb4SAqWGCpyDkgnnZpRhI84ij8ziE0tyW6pH/UiiuyJydqXk/
8fhsdO96IDub45a5ggJzKBVpnrU1s42mK14ao8YuuqyHfL9n+tfnfpkvr4iWq1gNXHW4tiLlTZAC
R7Z9RgZTdLP7Adz/EZQs3SZGCnVeEEu0adnAch9S+nZQuTh4b9nAeGV4Ul/6tZHBSCpvUYjmSJTi
i31eWRetXvsG6RjiETlhTgjcnRfpGeQItalaFUiDzuXMcumrThit/TM2tTN23eELqOH0HuNmE6Rf
tQwsq3+TV2Rd6zbxMuVAFUquJtc11QdkZ5WIRP6Qk5TcGhdfU327LRR1IfjTLaiAP3geekXSGEJw
DY3Y8rytw4lu2XzFPqo+YJzXaj5sJpsD54Bh1ew7wfZAP2R/UNreAMj/vIlW594QsriSIInDxk0d
COMMh3mML27KsKP2Q/JIhbwMh85/apmMKduuyBXSZxNDrGtkcJ8xmaG4cCeA2kvNeaOsM22jJrwk
A7zLR1fzJYDbDBtyYQm/8r5M0MMG9+kLbL+m4UFmPtyNhasZ/WvXwzfeMQOdyQ6Lh5SPcjpUx2Fl
PXAZCxe+Rd+YJoAZWHpcGHEMbyopd44vmZt9wsML/CmtfC1RTiOMTMGQ4GtcwpyjQyRjd8YcGBWt
mrMLyRJj4i3g9Aa4Y2Pe/KKUwTy5Y26YdgeQqBdA7DKbCISh/3SCYePYJruX8G+9UlQjyTqVjNPv
Z8b0ye+N+kljBWn3VggP0V8xHCC8cSitlqDlAyukE1NH8vMM3SwiXJi5Zp5OJzV7Q+lqMM0a4tDT
vPEISz6GO/rIg1nf5vW+tsoJDVOHQpbr0YWvW0c5nc6bOzKR03SSoB0S6TdGwhe/vrLzC5DvMk4d
0s2DEOsJ2D0WE/AKL6t99E53l6OQPGXfmYibEcY/BZaD6RZCIYSc6aDoCdu7QR/0g17g+cylv8Jb
uVKH8+5MyViFXBYHxqCRYFjFuiAQD758Fjwaq07OydRebkPvea7u1alPoW4ZT2D/EWiLIxyWmRnn
FqVau4J7Rj/fXsu8aW+ETiRn8fYbUqxYkqUQ0YCa4NDLOkvS4KJhrE+vlBziqZdBMHgx+Mr4F3K7
AOjerio4Gx4MErvzawCjo9Klz47z09T45aRDylEkCOQQwwOSa5+CfYOTAIy55xo21j0BMYomk7wd
cw6LGU8aCO4sIvPJySQgQgOK8Tu1FYgft4U4QIYUx/deZAXC0eOK8RxtXWpiedaKz/lkH5NIvYAh
ihZqwtZiVALBVIIIx+T+dd4lJVrMGcWskCIIzWyJ0U061xjp7W9/aCuJg7OLri0HTV/lI4Ph2SvF
1LQ8fpua/bXVFAweoPofiP4lvH4VxavkjZnzXFLRctyAtIt/acetAW19bAHlBmyunX/AzbBp10m9
y6M0pYJeCQ6jAsNSe8mLf4S2ZT1uu6QZoWfBux1h3L3E1rbsrJv639mljRKpHW4m+RKbTs4RcpZ5
ho+xPHo/inx5kPaQM+4q9yPtFOmw9sP2thCme30IOSEqbHXuHAzwsKEIke4RbJAb6uwdJP9m8BbZ
dH8Rf5NgLsQuTqsylNvTQffzDFQqB7lqc1gUvYPJ6bqt83wl68aYDEd3Wr3kL0Ic2E/NcuGhHJm2
i10ZJ4AWnOOxC6FzFXaBnXKeT6SIE2trouJIOOQ7iX21cDCtQFTqOkBL7pL+qNYmET0G/+IY8U4X
pZypJSl4JIwLvMqKRuJg5uvxbH02b5+OwLOZxDe1G4kHssqdasUFJAkzUTZfHPXpAxn3U4PtHm2P
aGLIWudzCI30OgktARtuDPsEnw==
`protect end_protected
