��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P����6��	���ǔa"XĽ�1�]��3��`�b2*r�z�ſ|�=���ln ����VH���.Z�р-�&(�IyO^�q��#�nv��<�;��r�)������S�kÖ�N������>�0a?Z�+�"�{�����t�0Iu���j,�J�B��d�|��!�j{t-�j�����{Vyÿ�G�W�P��UoG� Qϛ�U�Ұ
hm`���.��iL�a���F��	�^T��A �WGY�*��3���m]�S�D'�>��gil�)#���u���3x��A
t�����wf�^t5��k���;U�!��Rkhrנ �(���U�f�b���Cl6��7m����?S�h�,&@�GW�'���B���F���U��������W-y�N�<��:GW�����wVN��<)�����h��?��y���u�c~pl����zP��}�^��X�l��<2=ˀ��N�C
(S@���.���P���G���txJbo$(�OM�K�#���o�N���Q���p�x�l���ԣ=�������ƌ����\��B&��������P,���z��"el�o�=��-�=���fi� 'W<�RZ�&��͘�'q�@��x���c��W��l]��� !��XCϫ9�e=Z%��P� �S��^��:,�ųJs�煏�MyJ����� �l�ܸ	\�֍7r
�8��PgAz�X�l����r���sS�SS���VX\��6+���f� cN�Dmҧq�G��葕�0kN*����F?3�2�$�ND��X��4k���0�-;���h��a:ߴ2��p���V��7'.�v� ��T�4֣#g��I��ԣ���-4R�4TÜ�w��������Tm}�"I����ς(�:�[33�GdV��� `�^�rN���C�F:^r�nL�����@Ȳ�ma�4��}��gj����u\
�����t�8�'t��:�;������X�rM{�R�C>#<���l���94%��(/��u�WW;'[v�����C�jW�5���Az4Ou��؉��l�d�S^&����S��r���@뿳T�x�t�ZNL��E�����1_<M[̫h!�x�g�#�iz�/z5;���vh�����_n�P9��+����m�;w���A��x$n�Fa#r����:����t����d�
�.c0�eղ`8:�1��O���*�قRW+ǘ�-����,��hG/)�0���DH�������CdSfv��eU�X��{��ii�LA����qa1V�fd{��n���Kqx��H ���~ >j
�:�ҡ�2h$4�G|��wY-Φ{�l�q�0��K�ֿ�M9�c=�Ջ���D0�=Z�a�~�βM��9��Fa%��FH!Y�i6�uY�'eX=�3��r�1~������3�C���QN�@j�<}�9z�I����l���+����%%��Q����)e����|�:���$GO!�7���3Z*7��� �d�:Լ�:˓���s ����tW�<`<<f9�L��ӂ�r�\}R���s�#�NK��V���,���Ip���0����yw ~N�i���8���}كow�����߻��3�&ma��	'�JSJ�Kf����Ea"B�%�U�%m�oi5g�s�)�1�s�r;m
m	r��a�+鵋7�	���h�jM�<��y������ª�Q�$xI�U�c��$>Gi�4˟eʋDO���'��_)�Va�B��=��v,E	�8=y-v?�b��M-F{��a�l�W���h9�Ltpl3�\��:+�M9)���ӗ�<y���+'5 ��~����1*�\����>�70]GІ���i|g�4���>	c��c]��7���zoF�kSM��/�ӝ��
���y�r�A={r�
�D5,=��
�B3�NBZƏ�$!��N����@,ö*L�}X=��H�~��*rw;Bĳ|l��~�(*'�������&a6мj�IS@�p�-����$�kPF�Y�m�s�cq{�~Rz���pf�A�J&�q�P��f/Ȼ�&�Z5X��&2��z�����w�M~���{)3�9���ٕ�5�h<���Y����#ީ�>�x�&�}�����Nl�/�+I��P-�$io@��ӌu黢�������}DNXV��$Wn�j����9*���B�;c��o5{�N�N�����C���Y��
)\��Q�$ʴb/z=�d���$�:Ӂey�zQ,�W��!jj�ah�oC���R�[��яZ�iZG�`����9��<���M��@K7�֛ɠc�^�������B)���d}��,�9K�g�W��LEl~�﫝��\�U��(�x���,t�������uD	�1��9�2��0+$]�H�B%�Y��R�.B�5��;3T{�oX6�g*�n}J���0#��@.�,%�L��E�Qx9r�����`�Zrf%rm
��S|�Ԝ,�����4�p/�K@0�[��^j��z9
�5�l�&,D0=�p��J���jY�0�_�;�@�����B��B*��~Ɂ{��1�p%Տ)�l���$��qY0�R�k',Fi��z���4H�D�' dw���NQ@w��[�'����c=ӠSLY<��{10�,%��/���q2U
)+��Pu�L�l�#�:��@�ؾ^ٛJ}$$V�3���C�p�8F0�����|Pt�����n���nf��G-�f�ᵄ�NτG�����NP�^}�����?ۯ�͊Tmk�Aڮ���C]&j���3���#��Qxc�?��-@CG��*�(C���ҫ7��&L6��y�֧~\�(�a�Vеn[�8�<�@Ep��2�8�@L�.���?XnA)(�pa@'����Hq���gm0������U�$1���N���w=��L��h,S�V��C=�� H;P[�*��p,���B�G��!��A���@�y�ߍ�q�Py���" �n��c����Y��]��D	3\^a��W���Z �Ì�	�\��� ���ۥE��풐v�����Lm޲V�� ��Z0�� 4�e=(ܵ��ڲWy5��Q�2l��F-(]y��xXc�1�7�W����6{6S�]��ʿ����ї-�_���\[��3X��?�"��E��Z$�H!���>�|�fb�!,R���Bݧ6\�ݠ�Z1}�9�6����� f5<�7�VL�=V���>���W�Z����IF�=�Tx������m���Sq`�ސ��`@%b�4:�69�;2�AӜ���'��۷���է'�**[P�3F�7�|-�Fz~`����X�P����g�aP-nBH�������@3vbyDH�8��h޾�~I/��5�\�tn�Tyu8� ��+�hLP��b�6=�a��N�L��N��h^xP�D���&ʖ��2r����(PР�[���؃���4tP߶|z2��(�~$j`pnNA�0{��$٬��ڟ�Jݤ�p�W�`s�6���B��������Q�?�h�a@�İv���������}T>�:�R�+)����ԅ��xq;���Ya���'�}����V�4Q�����՘qo>܍G�&ha�b�6�y��(%���d�F�;J���/@I��	�J%�X��La��頄�b�����MMu,7�~P��8��&p!�뙁��D�\�_&�7��w���נ�A}f5���;�5&j�5 }��_u�
P�:�v�����Uy�o�_U2��\"��*�1���P�ΊpX*���L%|Q�0/C>>�� ����M�q�����8�x"L��y]4
�ҭ�㪝��.f��n�h+�7�U��n>a/`�/:��.�V��uinh���[qsˁ�$j��̯�7-R��O�mk2�~g��L�c�JN�2kf���
7g_y�u�./7��n4�/&�����l�f߰��π/l���2��(���H���3^[��|������-|�-�C8�1�p�`DoE��~�r�0]��N]�L�w��1f���)��*77߯�#�9d�R�c������mB\	�u©M������8�No8��k>���یr���\7�=6|5��i�j�/|�+���������Vh�G���f��@��-d;���������2�S �>7�a�.���=�'�nkM�d"����ķ���v���ewTVJ�������qi�K���BeM�;2�~>��XF �f�ul�>]؝�S�,9�A����Cɬ����3�D^V6�A��� �8�&�JWPH=l�ՠ2�G���`�ke���'�
��P������v˴����R0u�u�(�9�lH'��$"��k��.�]�iT�^���)��"SN�{�(ط-D5e��(���1.�!�{�IŗMBG��&�4Z�fTN�ۯ�L�yRn(�X����wR����C#�u�*n�j��Jw�?�rr:xâ��ˉޯeO���9� ���!�H�j��Byc�SxƉ�|Zi���U���:��E�=�&ќ0�/Y~-���Ym� �k~���^��Ji:�^P�#P�U4���s��N[�I��b2�0y���\`�i�S-6�s"�ϧ��/��t���;L}9zʥĄ���U�&�{�@���c	
��.%�?υ8����>W\��H�풸��|P̞�;X^6�2�C�1�E���S>$	y�{���Y��{��f��vչX�2	D%�%��H�ĺo��<ځ������^���sY#��OS ۼ�#CV�ŧ�X1�`G�� X�u^=�nE���^8��x�z�~�u���ݿ�5������,ԅ~����pL�V�H|/�7��U�g����KZ����PM��p�PE���J{�?�M�s�}) x��8_���V9޹7K�@<�����_rҼs��(�"ĥ��ɧN�"�5 h�]��\�$�7x�±Mj�M���W5R���Zڐ�l�g�g��X�/O��m3����D[�E��mnW�;��o�g|�ݲ<�����U�9��Ň�~���s.�Hţ;O�t|aFpm�H�~+��|�ΨKHb�!,����� iV��~�s�/��L��;Y�����a���oU[Swp;1��g[\���L\`-��aô�:�!�	�[�A��كJ��gNY��L�4|�e��t}[>���4�
������m��3t�t��7���Bb�ľ�%�"w�C���U�GMo���!
QW� �Pr����2S'���g���	���1˅�٘�0�ȟ����g�M�Oz�w���PE.��S�k�3۵/3g+�q��-.�K\���=���/~�R!j��M���J$�ͳ��h�W���_���@�w�����D�g޽�3��]��f��e��Cɞ͊+*���TD��������nnl:�;��z�o �|>e�����J������lxTK�X���"!����_SH�9���܈ժ-%B��YD[ȩ�\v�J�C�	ލ�]@�?[Z���2S4�v�����6Ӌf7)��z��4��qw��g���l�x@W�@j���cg�l$+�Lc�Ƒ�jm��u�7�ܼ��K�N���>mV�b��*����;�̂N���j"t&^��}gϧ��.�4�(�~�@X;�(�?d����D��cJL.��	04n�O�:�V~察�ݬ��Ob*
�<�w����ZW`�1�_'�:�=��C3�.U��4�@�8wH.�^����:�#���J'0$8�z
���h�g��p��g��1�v�\����;���%���&��W�"�q0>�"�����c4��ǂ���{c��2
�Q�x����u��x���.�:J�폗��� �ݿ%
@L�o;������7Z�Y� 1���Fƻ��A_1\�0Q��[n9z�m�TΪ�P�t�hʾ���v������W��Q��b���q}$RO�d�}n"	lX�M�]�K�"����*�hj�Hi��h�on U^��=��KF�#�=v|:��|(%<#��תY*¹��es��!�31��]�@o���[�}��m��*�!�ɱW��lZsޚ7�E��`;|����o˳�Zl5�	4���y���aw_)��{��swc�{D�^v,3��,Oo��9m�����$&�R�K��Ơ�;1�������7X��r���hİ1�U����"���b��y��S���p�睭�.�9�kq�nLA��7��I��K	��,��en}����ox!�U��{N���ް,I�>��,	h�Z,�����Ӳ�b��
��C�7����H��\�f�#��ϡ\�p|;Ҭ[�=M��&{��[8�L]��0���b�����x�7J[���&�y)��8��0g��i
a�>5kK����f�q�L�^�_�n�vk]= 
+���p��T0'Y�뚳OAMl��BQ�ш\`�Fc��I��L�Ӌ6\xǻ�����ة�Oz��OϢ<R�5�B�ýk�\��<���t� G]~p;���L�L��zQ�����{��&$��"�B�*9�v7��h�T�d��x0�����5}�t�m�c��OşEZt�w����L�v^(.��Z��f�OOh�R�%����1~ZU��Bv��o.dxSP.�C���2fW��<�����X��5�/ ��ID�Ln S}��k�
K�:��H��0E�Zw������?h<|+�L
X�����G�}|&�O"��KHF {��f��������K�Qͳ/�|��٨B��p�v��9^��؄k����_�M��7�����Z��w��2�Q%q�\�.�6/�}��t�]G���WUD=��|�(������%ȱ�:u�Ԕ:��u �UfA^�g���Rt"�Z��aޫ2�ABǽ~�M`;�7�N$oX�xp��#ͻo��;��m4�X���y���[��ǩ�@�����\˹�P��g ElI4$���ʺ$�B��O�4��!��!���/lֽ%��$����h�z#RL�U:W�&�WŌ  ��h�XJ��9�C��Df���XK�8���>��p<b��"$�!��+�e���[0���+����cY��Gw�7r�4ԟ�G)���TuC@�sn�r��&��ZM@�̒���v�(퇲��;N�6 ��A�S/x�MH���<! ��K��;"�ذ?��	�{6��l킋���v��6�LC���I0�����XV�BÈ��&1WS�y-�Mb4�|��&s7��;�"�E�� �m�(�we�\A�����-Y��y��,E��6m�զ���-|{�eh"R5�Lqf^�1^�:s�NrU��!*��^�!(�}�=�o��c����a���N�aӎd/D|���r�L��ĸ�c��T�w�C�+X��DLbMyU�Y���`K����+d�Պ��ʅݚi�6�˿\��=@�AaT��m��"��� ��cO)��-Ċ�a��ʻ@F8�ŏ�{�����y�9#�2�2sV���.$���A9�����5��]�>�������=3�%R�L�-������t�g������R�s�I�u��j��V�tQ��M���>��h���*������+X��C@ ����S�@@,�X
��&�Ce5t(�Bȭ�����;�+�*׭lEaˏ������X��s�v��q&���)פ1�����Y�5��_WJ��l4mU��$�M�g|`� Z=�th�!N<)y���V��
k�	U�^���K���9�F*�Y���@Z�3fy9�G�����{�d��a�L dn�2}�6� ��)�«¥?������W�I��wѱAh�>`8��#�膚5zb�M ���E�r��+���f�8����Q�d�1��D�$5ML~�/��6��+���i�G(����Mb:4`A1o#���+��r��Uf+�Re�J̜CĎ����Α�IA���\�nI��v�X? ෦��i��eqX��_j������G�6�;���!<��� `�I��bx������'^
��x�^�m>�#R�t�O�&M�C;����ˌ��Y���xԫ�Ӆ����Mŷ�S_B���yV,p��/"m`u�䯮�HRT�5׷'zZ�Ĵd���K��ܐ�,�grjT�8��NQP���R��Gh_G�֫��Q�ES�C6a��)�����ZD��\�^"�"Bo\�|��G.�7�C�_�q�TC���E=&���]�[]s�Fu�}E�����U?C�J������&���y<O���X�9�|���ևu#[�2�Ef�1�09�6o���:bXS�CY�F�bz#IL��=b��e��&���b~ҿ�L����l��΅Z����逑��Pj�6<�Cvp��Yǎ�Sl�r�KC�J���˦�3ӛ��⚌��Z̙A+�á�ڽX��<��(��I>E��lE�_�
y�����B��]m�B���N��\���_T�e�`9��G@�2���{l6�;��u��g��?�}�q%�fv�P�o�����(Vsw�`����7�O5lS9`���J�8��Rط
�3�}�+��+�sx�F��-.J܉3�C��{jF!����`�ǝ���L����t���E��o$w�}�wd���C�܏�,`����Wq�E�
�����!�n� C�����6z}:ڔ�vU�f�B�?U��v�
B	�3@/ l?킐&\�`��{$�{������P`�����ɋx=��;Z��Y��+9��p/�$N0)�y���d�u���C�=��q <D{�$I�����Y�`�궝S�d��(���n����'�@Q���%Z�k��
�A���V����?�n�D����b\�,�Jl��,5���� ���r
n>��&(��K?1�Lü�1�:-V�Fnd�.�j�b�}ܗK�ذ�<%=�%	��܏	��U�0@�Uj��fÜ/^�?�:|��]�p�`��zv����,��)�C"VpG<1@�6o'�}}��5���tB�
�@(y�
��{b��Xg��,���c��O�s�? ��9�[���38i��+O?�鉢('��n��╎��Q[�gG�_n8Gkq��$X'gU0��ϩ��,o��Ǡ�k�|[�9��h�ݘ?`*�����#DKr	o)�!p=�=��M�W6��W�;�<��HӾZ+)�uo����l#��c14C�.�{��$w�:v��i���q64�:����
�� $�3`AK;	c۩q�wņ����7kѽ��+�Y�>N ыGd��Af5-9c.sO�Я��"��p��s���kL9���=��\:�N�=-5��(���u3��lj����"�	*ox	R�#�˂v]���=o"ٗ|�t�|v�Q�R���e 
��h0�z9<��m���YM�Ǹ�1�g����P��o7���iϭ�_��y����QI/�Td��^`/[ಪO�F��Z9�w�VǛ`���>����̏���HqT.q�����~"uw�·Z�oe{����T܀'~�ɍ�JH��+��q��_Wc\�3O�<����p�x^�o,d�����>��1�t�0��ݛz�/�)-;�ܺ�![g<�Íߛ�����Y�D�ސkc4
m���9�GO�DdnR���'���
�A(VQj�6��&��_H!�4���ٽ�jn�2ؤfŽ6�����,�-�{� �~Y��8��-��54�0��/�yg�5��>���i�'�Κ�,eo5:�u�*Qx��Ͼ�j���=�3/�ϻ@�~�늹~�	`4A�03�P]�]�4	 J�hN�Z�_��C5��-:�l�U^��P"����,�.�@T��K ��!s�m���4���v�=a�WPH����}�iF9>tRL�ܱ�E���RȰ~���:��a�����~�*���#���c�9���%>��e	���ĕ\��������c�q�7��O8`P����5җ��xF�Ѩ�՚��k��E�4]'fՎ�Z5O#a`s�s�<pv����)���xG��� �L��+m���n����[��H�Q����KS�Of'�k}�9� \la����f�1�t�������'
�^��.�i�^	�����]
�d)��b�>�Hg�+�.BpH��lK�>��k4kRJ����rQ�'\���!Y�V(vG��$�5o�A�-03�n!a;�\�}�}�h�k����%7��|�R��:k�c�������'��I��?�BʧR���q�����u�颅2)EU��/�ZC�!��2��=񥛹k/��`p �6|D� }n2�>�����':5�W��[��#J���`�V�A�ѵ��E�Q�7A�/����\2+F��>�c�����rg�Ҹj���y;n�7�#�ӿT�U ������@�B4<o���iҝ3@�.�}.D�l��T�M���ꊕR�m�M�{O+{HOQ�]A<���� ��� ��{p�%Cd�R�@b, Z;����� ��9!���g�aW�S��kTpA��Ӆr��PY�8�j�@;�����h��=���dw˟:�`�²Ywq���OWq���c��x�/d�'"��#\�>yq�Q���Aw��ĥj�Ry��[�8�7k�:]���!�B�z|���h�\���҃�a2���q��R���[-�����S|8�g�e��Cg����f�!]�O=�i�جf���I\�,@�|�7Lϊ;�C�ô��!^Zm���A47'8MI7uT��$ô��F+�񑺱���a�>��##�(�N�0sh:��Ω�r�ޏ�0Ta�:M�
�Zx�Sd������d}���0�P6U�Z̓�lj��׬}�T>^�z�Y�W3H�u��=]V�HmA�*���4u��2�����9
��d�� a~i�(yԤ�h!�F~��t�z?R�yY�9��"�~k�`w�~ VQ�x�рT�������tI�xp��`�����jնYC�������r���
���`E=>x5��L�;} =MC6�D	���}'ݖ-e5�5���z
[hE�W�^0�i�NM��ƃ�]7��a��`76��+5h]�#�SPb��}�K�Y�0�J,0�H�\�8h��Մ�
F�բ{h�(��a���5p�m�<��昗���s�=���)���u
����cF�G6}]R)!p�FǨ����ƣF�̟�"�$U��Sb���H"�����؜��#O���蚑+��Wz��远���Jy��5)5���I�I�G5T��-]��Oa���`	~)��Tؗ�ЇX���N
���*� �چ#�5�񏉆�_`�U��$��r���$'�z�Y��^�,��~�a[i�L~(�jxy�1��5h���pw��δ4�1�������J{�-*ƍ��0B��Z�B��E�9�&�L0�^�=��ܮE�7�����{4c�$�.H��+�Η�^Z�b�ė��{�A-s����ԗ�S�e|g��|�H��Qt��K^;X1�����b56.~3��]�(!�~V�R�?y�}����݈/9��28E��@�]ϕ4�r�cj����+b}����Z�0���W�SR�^Q��T���.(��x��tzm�-۴],�Ďm��N��z�$�o�l{�Y����G==�A|�����/�+�hP;j��2��g)B=A��
#m3�d�<�IU}|<�D���=�oWׇeFb��aj���h)�f�OU�����7�J�\�:��Ad�	�_oc�C�k��g��$B�z���轃��A*¾�Ykfǵ�B	Jĺj�%:��ڥ\����C-۶�R<�6i�]������p>,��}Ǎ��>��Lp}��Ĕ����&�B�w��i�#t���s��5"��s��5i�r{m�0g���;A�wr��"�ۙ��`*c��^z�c$)*z{(&������P��R� `6�=���>�g���%J��qwū)4�ǦM<ɹ�r���d��n1h�C�a~M�����P��ċD�$�Ȍ&"�g�)���"���ܢ�31SP�����,�D�LW11k�C(���������I����(P����Y�ͫ9���b��\t�u���L'1�;�h��S�kj�\O�W�Up�]Vf�8�F|�0/����@�ԛ"@OhRS�q����W0�����F���k�RD�B��9�ITi���@���ˣ�pH� ^�D�7��� E@S�ph
r4C&�k�Lܲ}�o���`8f�ϘK1u,N��蝜ij��:}�h�('���Xt:�-c�%�m4M�6�?��
�;��tg����8lNA�HB��
}x�����Ǝ��!;�@�D���W�$	
��j�8���8�H��VP��o\����/D+���5� .8� �f���	�L�]�{,����>
m�6NǸ�OM4������� �g��ݝ)=b� s�+�	'�A�ⴃ���F�9At�K���q�����5����z�6�읳�Sl	L��
ɳ��=r�ݍƕ�́$��j���>�#܎L�I����j�d�!�?�X	�\�=�I�I�#���Y�KX�E}e��8}^�
�)��s�'�����bE��-�y!�(+jHR�f���V�<)k��`�C��*6z�=r�C�K��k� 4+�AV+���F��g�tE���lh�;�Z����(���V��<:�V�$�o�	`�~TjT��V{�t�kvVX%RR�x�r��V�o5�������6ճB����e��Sy�X8M���Q$����z�͗�An��0���[��q��]��Ay���p����:8�?�b���XO�.u<n��	2���y#f��S#£?��7Q ��1u�^d�����{k����'c�����D�>ɠ�R����'��'m���2�$��� rǺ��^Gѷ0
���!p>d�����q�>�.�~���z��$�mu$�h���b'���e��sӉ̴��uP���yZ���h��Ex�~����7�`�l�-�o��ilg��XǇy W|)��
,ξ[G֍g�q?y@�5��M�w�W�E�ZP�|ռ�C|r��8 r8�QQ~��V���9u(so��kغx�����L�(��7��l�l^�����S9�^E��e�����jc���˥|<�Fxj�Sm�M���ƫ�-[��G�����K��i��J��iӯU�? �"����2�!T\���O$�L��ٵ?�z�%߶^b��0����B�K��� �>R�T�3�������)6��L�j���ψ��W%����	bQ�@�&C�󄤍�f�A��9�@�3�y�����_���[1R��$ ���77�w=xj�¯��H2�uI�4�_x24��pK���e6��n��S��i����V�U�Ӡ�����[2J�vG�gqo�J��.y�[�?�N[]'+됬��s�g��ܴ텺?n�1��n���%m�5Ĕޣˍ'��-d�#H���Ԅ�QOZ�~����N:�*���_3�o[�XQd**������|�/�+�"!���������]G��A���iV����2"�l�t��Cѧ��g�҅ �|S�+�7bMx�W��*���k~��c�>��!6ד��E�\�d���CB�1�x���#�ޭX��E]��q��O�f�.��7\�ubǰ����t���O]/w=���"o ��%�'���+w.�ȝ-�W��L#Ij�8ݛ/�z��ɪK3�d(�( s��j��(@�r3�\$�����NW&zѫ���{sPdLU�c��:��u�`w�e��[:^Gܗ���Ak����}�����Q0v��%~��%�R��+�γ-�.������*;���l[}@��D��ۣ�!n2��"�j�ӭ=~������|�f ��/���S���_2��; l���T���
���8��ĸ���.㺓�Qs�t�DlO��E<�B���P�b�v�6�7`;���+de9�Ui��k���B�ǥ1��j;bS����N���uC������������!RS=�"�ʴ��P"X�j��N���^W�ǁ���-����f�~Z�hB�6$`f`O��[�c��Q�X�	}c���'�<���E����8�|�{!Q���U��Ӄ��|��6�����3���b���7@B��bQg����&4�s^�j�2�^�)?�26k��<3\�@8ͬ�DD�D��P�iI랦6W���&r����#�k]�g:��J4(4R���%p �J��L�n[���(c�-h��H��������E�HC0����[|� �+��m�H��?�����=�o����� �RR�
j9fd�	�1��}1����X���h�za�/�š��q�0[�޺{e�{��<-�TŤF6qA��$�{����<���,�>KF]���/���>�'���`��V���R�]LӺ^�ʝgŮ�BL���{e�g8�O����-8L����]����cE<�t�n��B��be]�W�������&iG���X5{��Js+š?�[���\^4��;�|���Fg=�x~2����������hq|J�Lȏ�:�� ߥ�g�����o�M�L�H��kC�`�o�A����	�P%K1-x�5���5v�0�V;��3|�ʄ��K���
�7CY�z��k�(Y��$�K%aN<��f���I��ϣ�G�����uCw������U(�|ѽ�<�<A��WHog�@Jb�4*Vݾ��ѽ�j+��+�3�hO�h���$�3`�Bާ�Sq�Q9HC��:I�VC�#_}K{�R���sʖ�ޥ�6�d�`b^�;�>�&>K���u��b�M�^C���{���F��>���^~z�x����W_�};�g��R�hB�7(jPUi)(gǮY�63�l��ZYeE�Y�|7�C���2�NsMo�nOu�w	��$=I �����0��w%uݵ�_C��?���Y��b�:�*
-@�w��&5�qX�0ĩ�>�m5��f������M&��#4�žҥ ��| �J���g͝'��v{��n�*6�����ɌO��+�u����/S��x�J�l���nᘴ�48ܖ��u?7Ԭۮḥ�H�~`�"R�!�/��N ��}��̵���z���rқ��i�L��S�?�6�,�J��N�",Y�gӏ`wko�6Ewz�l��{�/c���!��*܈��D�Dy�(�wJ���2� d��>X�l���j;�^mU�� �!&\~_�M��L|���X���$qE�C+�ڟl�x����+B�!y�K�ʰ�k�A͛剫SR�w4X�*`(��D|�m3H�C�I��ώ7]dy����~fQ\���ڬ�֤�\���$Tv��*�|�yuO9"���i�:�؆��{~��s�x����[)n��U�W
�gD�ĕԘ;4� �l��%����dt��Ob���ٯ�3�-��0?/�u�b7���ࠍ�H[�J�>H��p�]I~�į��7�_���+0/?�{Z��2՗F ����RJPAϴ�M�S��%�13�gX3��:����z\��T��ز��B�쇒�MD�P;�O�v�����
��Xģ*�֡ǅ��uc,l�Y���
(������0 <����):o�e����\jѨ<���${�D> 8���\���H/���i,0�����3��]�[�m�~��-,��%=���0�Ը�H㛀x4.z��5Ie_f�X�IM- O|	L$��#�*�Ζ���Ԁ��g4��&�x57�iN��O?ۥ�lX��\�?���7BO�.��̑C�^��3/?�qƠ�x���@h�xKP�r�VP��@�[}xz���A�a������n�d��aN�<���0��u��U/Ft�7���V�����{�hC�i�85��9.��I��nI�+�%�hQ�~b�o6h\Zi������T�,}��u����WB0{Q����K����>���NK�e��d��x[�C�r1�����!I����kr�����\����.:J�Y����Ơ�@c@�
_�cƣ_l���}��-�TbDk�C�]���AɃWfu6��	ǔ��-8�;��]�X��r�ya��8�D�E-�����f�k�/)�؞��6�E���TA*\�בb:�D"w!�\c�RkkO�+�AaqUG��=���S�>�0!"U�N/���1�Kdމ�>b�2��|b1D�"��v��}���V��g��}O{Z���ˇ��전i�����f��]��Y��N���n͑<�ݏ�8�LZv"k�d�R"�.��3�*db��~)��	?��s���u�Tj���9.���b��W�ׇ�������83��
3�g�Wh�[D`���%��nZX�\G�� *�P@�W�I��6�, a_j=�6��I"�C� ��I�1Y����ދ*���?^�oƨ��]��ns��pq*"����������[~�0��;�jmJ�ү=�P�)7j?6�c�T�pÚ�b����2p��T&��1 h�NN���oA�:,��V@��K���a4�����������!�2���oht�-����7�=�)�����1`еI��⊂[47�����F�QQ73���o�6�k��[UAY���1l�C�;΂�����{������<S|�ۏoF��!����OQ���^���@�@?�M�]^���eK��T|N��z��#�d�b�ګ�ib�6"W�?��[��N�ڴ��L�@�c+Y�����\'A/�;�����+�d}���L4�D���6��h#�܄h�
�/v�b�<8<ϫ�ă0�֫Y9�VOWVI�A%���4�/�6�z�Jˠ&-Ra	zyv,��}Tz��h�U<�U�����u��nZ�5��=����9�F��|R|�Ň�xë�U/�h/w�.q&��������p�LF��X�iQ�ǎ�������v0�+>�wl�y����������RS o��	�h\��a�H.L�|)<,��y�l3e�Ax�K"@�X��b%�zc��_ا�����n�p�I^���ď�)�#����
�T�	�m-vD��B$�N^�I���w���b�;��p\��m�r���SB��׽�R��P.N�PB����vV0r���������Br�i�X'�Ǽ����.Dsȱ��q�pR�}�c/�$��k�}�����fI��>lp�Wj�c���m��*(��}�����#�?E�5:�.]!�+jeZ2l	y���٤D�S� �� �St���*M}�N���7��r��?{��bW�r�
�0�$��NS[^��pf�v�>�xH��C�ʪv��;�j6���3�bs��΃�E�cU�@�+�י�E�"�F�-��v�>AA�C���arlIQ7�U�/?�	��i) pʦp��	+7��/�ՉhzKF��8��yU��}��Ĭ�+��y�h�kh�7�<�OO��	�`�.����	ځ;�ו���5��A�$�L�b�kp���L��ǀe.V��1��;U����nʢq"�����ǯ��d��j���3Z��OI❎U��yֶ�F#�y�����I	:�8��N��a띍��(���B�z��D�t�_&���Gb5�݊	q>dmSY��+{��x��� W�rp�^b��[���
KW*̈́�Nfo�����o�r����?2�����`Tgj���-�/r����f:�l��ޖ��3Еĳ����3��stj�S4?�;�>C�@��.�Z�󉷟�?�!�t�-�:����X�4d������������.�����G�Pu<]�kUU>�33S���F;
��v�ܿ�o2j����v%��$o(;�-�Z��j ���u�8�Tj�3�뺘u���q���Ղ�m�eO�KY�&v��N�e9�'B�5b�ǭ�2�+�gc�\��0r��ߋ��/���^y_��FZ���F�����P��Rh.6�+�N�!K����k1�x���o���K� ���C����E���n�|�&�m�Xq/]�'6��eE�&��8>W�S�qVg�ߺ�.���e'	"�i��9��~�Y�v;��rj�tA±��,�E|��F��h�u�E�����(�(��9��5h4�5�E�4U�Qt��ݏ�7��Y�z �t?~������DΧYY�'�o7��rQ�!�a�Nnz(����pXOW�����;f���5�|d|���a�~���{��JOA�Kl�9��_+uk��Z��K������Y�L�-z�m�OX8�dh�/�.��0���ez!]B0��Hq��B��i��P΍�և��B2�Z��OR��]�O���yo:]�R���p,T�P;vˠ�;��h<�5��H�4�l�:�y28��yx+S�@�+���(c�l�CV���:�-��������P)A���G����`IV�()���R�o,�[�/�L���-�d$�_ef��� FF]�+�GԔ�?b����<F����;h�(pvS7������ߞv.�H,� �>I�-��a|��Wj&���rc�yªO{�%��t�^د����OϨ�o���U����D�3�-[�`�f�-����o����ᴛ���]z�U����[�T�k��L��×W��v{'�~eMe)>V�oq�>�X1�^k����`oԦ'�S�+5n���~��`4�Rpg}�`�wI�@ܖ���+,Y�g�╷4�Խ.��]HU¡�8+7DtaԠ)�/BY5!PH�v<$���������Ma��n�s�V�F�x:����G�&�UoT����&.���<��b�c6���ɽ�U��Olw�݊2+��^�S�"A�dH���f(����l(�d9�&Y�Fn	k�i|�6΅v ���0���a��4�\9��H	N��4t��;�5.muYu�_�(K����#U�|2��e�_n�~<t A��6R�m�͉��0��a+f�yP��5CPa�{�����WR~@b����W��'�FJ�B�,�&���$������Baa�N�n�Ck��ʬX�p���\͐�������LQ:���3渍�;����Nʐ��s��� �f�E,���y_J��GO=񐪹@4�ڽ���j�y�}�;�'��7喝B�i����۲��P � �,��i@�a�4�qE�L�|��}�����̝`�m�̐�4�3m��gq�0�6��C4�n�"�*�/�1�2�e�P����A�l�s5K$��˓�")�,��������}��?.C�n2�dQ�������5g<�ajؗ]I�]�Ww(����:1�'�M;g��u��os@����h��78����[�BNaVG'���=h0��B�=~�s� 0�$=|%��y�p/��QF�ڄ����yB�]���83i�|�׉���#�=��1�s�&��y"OmB�^���R+2IA���f�M�$Y�Aޯphm��Y�'�)�Q�v�o��B�l�{�)��p�.3�hb��_|��-�Z�íǾ����$d��C�������6jLD_�8�:�DW�Z���_5��*kR�:��c���na�;st	w��N/��K��Ch<a�n&h=ù�Yu��E����L�h٦��_����1V�g�Pv�-�,W�vx�v{ T��$|�rȁˡ�ߤc.�\g} �u�3+�?+I���b6t�Y����	]1J!K�㚏�TR�><!�5�C_8:� ��v��f����ͼL��~���Ӽ�
��S"U�d�Ww�2=~���Һ��_��vZA�̼� |˽-��Q
 ���¤�g��P,$��
6���T�as랖{<�F�W�'t��;@<�>�7�n)���RjY���5��U�~G�TH`�$�Hi�?�6�Z��gT�f��&k89��jyݒ�7����;�����7���?�o���q��o�4��ty�:���ۊx��M������Kj�5F��%�x�S�S	��Bpfΐ��׮��Tղ�?#�y���h��]���6�i��G���V�U���#�[|�Yﭘ�Q�[�E|�WgU��T{��@�:>K����Q޲��HŊP�����y�3��6����=,���9J�f���Ŋ���aD��lԋ��ﲹ�y�Pm�Κ���a���T9���O�]{q�VleKP��g�Ԗ�33[���pTR*��h��r���*)�@�P�/�;�����=������-cI�W��-w�k�
��z��&�bx�q����or�l=r��T*���o&�N��ڏ�r���a~X׆P��yUxv�T;LP$��8qb^]]��>j�^�G�{Z�a��̄�P�G��|%�ӕu�+���e�2g��UC��rO_N��-�`�K�	]��7!DgU�3���0���]5۠(��C��X<ŚUR�ȵ��~�?<����v,���Q��Q�T�6��]����d<<��H>VS�� d�1�媐r0K9н|�G�}�$�乊��Eο�Z�Y�T����ت ���n���Y�ĺ1#�T�IEB��ٱ��T�tH-?��[���w��l�T�>û��(��o�q#Bx-1Z�Nl�E5?'/G�4Hׇ��
�nќyafs�}��tC[H���	�Ī�����|8ʟ��g����޿��z`�|�N-��3xa��_�S�ˈg��R��l���zET�sxO��G�]�^:�7�h0�.�RK1p�� ͽg�;��6�/J��ukՕ�gW#V�&
�z�q?F��.:#��u�Ж��!+[ؕo���>��C�M���q|���jDs^����6���u�g���֙u�5� �Ht�px�c���k�WH�+�X��.�UV�~lO-�nù��ڿ�[�STکH�e&=�(T3,�iE��Pi�e�z�ԧ��X楿z��:�_��~ N�����������fIK��W_����������A��	;8�P�#�R���&̒����uR{��XX��Z�;o]Sʼ��hgE�I��UܚG9����+�/@�^o��#J��-����1��{�e	��)�G�ɟ����Cg�㈊Q.������	����#=��c��e�+�g�����ޭE$'��b~����ǩ��hB���YGF���)�zY$y�ܰΦ��~bB���Q���a(��I�lo@ی���{��c�Cѕ,�~[X�M�/�B6�/�'(��[,�7����K)�Yi���m%f�3�oQX�8�L��H�0H^T����������`Ds�-f�O~�����vऌ��w�ֺ{Ejx�j;\;�&�P��IN�qH��f�����W�f���q�(7��7sQNR��7ZF-��+o�TM����i1�m
�(�;	�;��x	�Ǌ>�W &����.^	*l�nQ 2#���1�2z��0���5a#�ڷ��e��F�թ1J�������5�G'�V��ַ@�ZT�e��ܴ{�i���Z7�G-��ʲ�"�.]���HWh�
�����dCp͙�:u�zV�1�uZ&������ÿpa�K�
$�X[	�,H����x`��r�d�����l5�F�O�����⎄Zd(9!���83<^�Ǆ��7��b+D"kp��X?=4m�Du!5������9����]����<��mf^d0hM1-No?9�!�^q���P�H��kB
�E{�� ���ar��.Z*q-�_�'*>����"���1j�hj~^O����Ϻ��f5M�C��p����=-�^Е��[♢~v���I�Tz s�M�zM·�@`nےz�����
�`\������~���" 1.jğ�Ҭ��}/"�A�4�ɺ�~w�%	�C�p�u�ӆ�埒�ig��p�F����K}CF��B���~l����y3<�&�k'zj�jA����(]v�X�-�qi:�C�9�u��>Ŗ��q��:5��~0��,T��?�w��w�WfĔB�wD"����������o	BZ#�t}ͽ�`5s�h䍼Y~x�h˟`)J���"1au�#��_J�L"�y�'��<n���4��}��)r�X�D^򰪮ƻ�~$���W�����)0qO�(;:��?Ot��Z�w~ą�wP���m͋pn4�S�ӛ��]��Ʋc���ojJ�55���a�J:'����U��}�eRf{8}`ޥ	��N|�X�)��FW�f��-��PV��{̱��ɍ�ك����C'0l�Hˋ��j:��hj�=K�ݔ�)D'��LM�6��k��� �Ҕ�iS�/3.|�RX�mW�e N�'�~4��u`!��g����J/.����K�Qt^�>�Fm�h�K4�3@�n�2�g.1��ˇ�R���L�����,�z�#�
��v�(�%��U�|"�ڈ\��_��˾�t�AP� �깍��w�L���:�{83\��1�]r�1�=)�R���hw ���B{i�c�l��,���f�g����t�e�:*�b́)�u�ǜ)���2Վ��Q��bBhɓ 0��X Vy6/O���?8f�Y�#�Ւyۻ��!;iҲClF�$�#�q!5��[II�H�.6.��ʆD���F1N[n�2�4�Z�'= 2��j� ����_�ց;�)��{����V7��YlE�Ox�>����a�(��A��4�՟��o�Oq3��s�Z�����b�vP'_8��Pe��A��z��!��bW��UcA�L߬�fJ�%�Ҕ��segg�Auq�U��v�HkT�r�v	�3�B^6�b/
 G=3�۹�T���a�2֚C����2D�ƀ�h,{���l�P�X.�'KCUW;�=����v�����|��X�Ktۜ��Ɵ�#�/Cg8�O�_�u�0��2�P�1e2`���%j�;У��L��_����.�\�& m�g��^���ɍ����/����]/4q{�+$�Մ���]vK;�V�b>��	0���l���fyL��D<U�d��Sf�Z)Ǩ�F�o��P�؆�������������d[��66��(N��Sr�=8����>|�O	���������Mщ3t~��Tf��������E�'V�zr(Lk�]Ŧ��
)K�[��ż��o���7����U4��x��sxO�e�uoVUǝ�F*�a9|�w�,�k���9a�O�oI�ˊ:ms��1�x��}����@@P��!L"��أ���F��E?�+g7VȲ��ƣ�m���#K���S[}R�a����$�2�ت@�?L��v^�%ꖗ��vWZhp�|�%T���o��>Aiő�.��Q��=��!�5���ʠ܊���g��Q̄�o�݀�فr%��(��N�7,#T���+T&A@L�&h)��%��_.��7*^j��d���e҃5�[�/�=-�������������#h*:�3 �:K��.M�C�9ڬN� �Ȯ��أ!@tX�|�>�= ��Pر�S��������_C����bʿ0�ZZUI6zx��Uw��E�d=��I;_���ߜ�.f8񛙚�/�n$��K����?���Mp�"�G�L1L��ޱ+ۤ8���">@刕Kkw�OI �"�y^JX燒�%Gy�:̒?��!�~�x��2�H#!��ƫQ�:g��7�И��s��hs3 �"K��R���d�_�j�+t�fbNț��}z���l
�r�dI����NU�q3�������W�v��ȇ�}tj����El�'X9e���@$m���c��UG<%y���arB�Nɐ#�JMfj7-+�~~��PF�k_��<��<�}:�I�y`~l&DLC��NS���ԥ���f(��Ӌk��Fq �c��X4;���'���)֙d��WR�ӳA�"p�[���R� ܺ^�'N��/�Zص��u��$ۗ���V�Ŗ�7���^�ZQ)n�.A0�勎L�^�͡�"�ǩH�e��KV�EM	��Qn+Ẅ#�1���Zx���$a����o��*��nP�:7kͬ%zF�W�߯�=���j_kq�C�5�f����_.�xc�{+d�H+��j�lĬ��*��U?�V�E�K�4;������M���%��PE=,\�!M$ь�Z%7���fٷ��/!8b>M��(�c���,���8˒�n�����v�L��
���^�ȰG`~���r�2f^�@T� fN�����xw�']p���F\a����]���J�kٖ�俌�\�7���v)b���.D��ϭ��ݚh��qy�t�����6"��*�)���EкFvEUw����a�u����N��x�p�Z�0dHC&��
4LxSw�Iq�'�n�S���
�������ǖ�s�������['@���;o���~19�*`�$���ڏ�S��2hᷘxS
�
H��yx��Ç�2`��-S�͚�r#33��a�S���Ĵ���& �X�V��D�d�F�N#YĐ9���o��X6+=�%�]�!��h�@��^��»)�r�LeT�"<~�Ϝ9G�?'����Kz�:���96�e%����"��g�uB}o�D%D����(ŕF��$�ҙ�R�Ě�CQ4��|��1�[����{��e���x?�lM$�u���T
���Y�Y�BE��=*������1�!"F�w�xO��!��+�q��*��F�;w2:��,^\k���8L�XȀ��^J�c�I��*1qA�6V��Y�2�����ƅ���t����B�͠=�N���[��9�l���(�">e[s�U$VC��-��}HO�:�]��#�U�/:!�оu���y����!���D�	�w�(lM��jS��p��V]|'�Y�K�[���:?�Ŵ�H8�r��b�s�l~Pց����c`�|�'��NFZ*Mt���-Ǒg�+8�$b@:c*Xyj�/��fM������^}%��@�o>^�&d{J�s��]1N'7E�#�5[���gc'\��敕ƴ(�+�������-�:u��9E@ȟ��
�7�i#1������"�����q7T�O�Ů^Wd.c���}kf��!B���/Y`�ȕ��yՅ1Z�`T���l ��ֺwm�Z0Y���j��sA9T�7�es�� ���Љ�X�a�pnrL��t==�P.�,����TØ��*J�J��~���*�CI�V�ۏ���3fy�h�ĬP�R@W�x�	I�t�R�\�T�I0��ɍ�O���<��GP;��z�* �����߯�*A�#<��-��՜��.�tcf���� #&U�*vR��}�#SP!�x��G[!��/�`�8{I��U�Z��An%��ԕ�=h<����N����c!A4>��Z���ɐ��c�m@�N-�T��ǫc���AS �!�4rm�����l��<��T����/8�w����M��q=��9\�+�13}��5^b_]A�VH����A���"��֊�n�*p���[t�:�c$��e+���e�ł����i52^���I��xS��Z���Q�ȉ�qR_ d@͞�g���%�Tغ���k�Ч%��Ә��jy���I��MaX ��;���9Q��m�4�,-o��{�.u�3�Kg��|����{$8[���g�Q��y��Y��P���/]��_�塋�I�F���c���%`��E�	�Om�:���Lv���0*���=�s�?<���h/�� �A��:�3��=�x����nx�U��ܨ��@��F`:�-_�	?L�K��g^rdEY�dvS�.�)��ſ٘����A���G[#p��r��V���g�����mq�Ǘ�.PUˡ\%���bl�^��nXܸ�1!��L$f&:����*�Y�SCkz�9�ӡ�_C`��]M�?��g����b�rr)�a(��;oC8�J�k�jE��+�@����P]Z�[n�&g&<�d���e��y�k��D?�Ҁ>�ann|�T0�@��j�T�ZQ��a�]�ddk���ёTq7\�	�_�KX�s(DK~��mI�pjϰ��O��N�A6��T��~�|{8UV@<���b}^�ߖ��%�pl�ɏ9�ER����'P��ln�t�_��Zy�aԂa[U������om{fQW@����t��`���T<�QRٵ���f��h�H[%?Up�I"� s ;�3B)?��� �)΅p�hͨ���=;DU6y����#������p�ɓ��#��sT�1��b�-��l��R��Q"��t���t���nr:Q�#��_��A���?7~3�iǎA��S�7F�H���P�T�6��p5@0�k8ɖ���m�����>y���f��EYz��їZ��A��(Lqca���O��<2m��h
>H뢦�(7���<�3z�4hL����>���u�Hf�����*L&z��4P�[�}X��^M 4t!�Ց�{>W�؏u߮���]������(����TPH۹+��w�7�yT��l$D 7�^=�D��ky�O�np�E*p���:��=�����v����,�=�p֩�)b|�M8��\#��n�J'�M,�����^ �v��α		��Fܜ$sd/�W��͊/��M������A�[�Txuyew�R�i��9�7��M�����As�|�$lz�vs���E1�ޗFS����~�*20�@�M�J˸�#I��FJU�.X��j!��x5vP{wI�C����<�o��։�U��2�q�Zp}E�T�&��䇺�i�^ZR�;Y�#R"�.cM�	�)l횕{&���J+���e�Ǐf���5�|09 �*�SW��G�(/��b�d�@"�����9����-ݢ�ś"Oh�W�n!�4@'���jzw��7����R�?���Ʃp�����'�|e�)��yP�[ D����Ά��H�ST[W*|���g� yT�il*�n��V^�K?�<d����TD�����4Xu�%�h{ ����Y,�[����&%$�zү��+uy�TI+˴[�e�c���� JS��2�V�(��*@86#�k�dSJ$ n��'���?��0Mh?�I�v9[6薥?�r�5?���/��,�������:�`%%���=4�Yp�Ԁ}e�����(���G_�p�T�\Gz����T#=��W�.*_S�MB�o7}@�6��4(��&�����x��"�;�݂�����ϗ��1�J�(�4V����«n��>��"�L��Jc ��̛s5U ���!�5�ofA�(O�#O?��k��"�w�ٽ��,�
R��ARDgzz���W�s��
"wb���p�<�x�9�������È�`��7���rɟ����LOj����C:T��L-y%�w��O�CKGVĕ8fJ�f��G{D���i�V�����+�W@�{���������Ye������LǍ	��x*A��{4��Wާe�ಈ������`����5d ��1Z�ګ	���[r�".c� �7����OSpNe��* <ű�6A�+�A��6�Զ�z��S4I�R�Z�
����H�iB���r=ᓥ�Y��k*�3s��#R�S���8��� k�r��3�E����奿?^.��,(��b�(�>��`ܾ����#�BMF)�/n+� �����b�9���̈�
q�lm�8��f�YU�V�W�;����԰�-�x^���E#�1t�����E_6@K��V+��ev���X%�F�Xl���.���]�o.��8����$i�eZb��[��}�d,S-�����W�:�d�X"�6sڊ�: ���`�\ގ�W��$�38�����ǅ�O1d�Z���4��PeF��(�+�p}��r"H��+�W����<T�t�_S�i���L�}~��∟%Lu�c�4���nN�zH���ŀ�댛XлC-L�l�V��._/C�XN���u:����}�F�q	�Ԙ���n*�b�.H��]"y�X�v���@�ؙ�6̉񏦭���w��BȚ��	Ӈ�8}f��ߎq�+;~��oD����)����|�MBȠ�3��0c���@,72W(M4�� �ڲ� �!>"՘o���J�6���� &�E��x����-���ϼ s��E3W�����"Ķ�^
�s�j���%�HlO������*���6����<��~pm��&��='~h 4�� sJaQo&�B�!7��(wY�����B-��+��z��f�6OUB�� �KБ./�f�����E�G!�����ހ�`R���'G2ܰ#F���͹��;B\��*]	��b0��葠����}���K=ȳu,D�z�S���l�@B0EO���M��QL�5=D�� �Hc�is�J>���|k��(I��������]�*iV��<���'�h���3���
�Z`�b�f�e"��*�b{q4d_�:�:"��	�q�qT��my�gOj0�.�ۄ��uGA���Ո^($P��a1���[3��#C�\@�`ʋ�B�>uݻ5�22	gM����y=�>4�/3�?p,xY57 ��M-ǫt��� nj��F��cuW�wʹ8��[)��Z�fz{
���(\��_�f8�7e�������Z��̩8S%�J"�PG����p�������F���K�{����R��m���B�{o�/�ۮ���KP�爊�J���?�� .�7�M/�����ک���,�I�yM \�>,��W�g������!��V�
n��-����uYCy?������f�,��0_�g��EJ$e꟨�Ut�D��}"�u���K�zNUF1���2�T���O�����W�8T�jp���a��.�X�N?�S��\ȡ�| UI�񳿓�^-L���a�v�`JS���Fcڟ�gvJx:���Hv_c�B��'�p�񉁡J�1�*���c]��j{m�+7W�&ۮ��yިcXr���+����pˠ�7��F����û�Տ���b�Sm��5��p�WEra��]��0P-q%���HIOq"/M�w�����Z�r\���v��sB��K����F?�e+���,�Hg�Ӧ���/(�l�h�
�CA40'3ŦK�3sp�3���)F�u[R��e�AGgu���7.��^_zkT�5��}6���=�j~*8g�m*s��Ƨ�[S�[\�m�R���̌Vr���ː���/ޓߌ�u��B������?�=�i��~Q���=���Nw��9���K���HP�h���
�)��Z���O��&&��O�q �*�R�ĕ+O`ҹ�N����^��XO�����8���l��^g�]�U5�����3�.;%{��KP�1Í+/UV+�J�8�$��F8�du��>\8v�:o��Lh��-*�t�xrJe�dI�i��!r���I�6\��>��0C�QQO��,�x>m1����2���Fy<��H��y\�l��:���V�:��kB��_&��»�\z�������R�������~4|�"�ܨ��Ne���$B�;|�o��]a/R?��K��x�42𽭥yQ��՚�y��抇�g/��!��q,�ܧ�nN�ΨO-���1Ǎu}�#5N�Rm
�p��@�y�5�s8Z���I�^�0E�z�g#�0�j��L���_(\_ooF�&��BN߅$�I��GH�owN��a�(L;]]���2c��A��"������g|o����8��7;ݵ5�+<t��������p�0gO&�~Lʽ�E�[K\QOz�'��G
���C��I����_v��<�����O��(㽼��@|T]k��樜������*�l`�
��}`	�����z��D��[�����Gg�]���i��� w�(�ΥyU�ttX�[4�*�y�Q�U�j���g�l��*�fjH�Vi���f����ڗ� �5f��� !�Ϭ��z�N_�u���r� E�ɜ����:C��Sa J�D�X�#����j}&��<=��<�d��_;���[ӣAS���g��ڨ�]<�0�I�J�ޔ�f�N#+.�5�s��jD��';���|py�5�>��������J�foo��b�d�@�Ȼ��d`�-�J�s��䳴���e��?\�?��]��Pe|D�(�#�vr����d:�]?Ǳ��yV+M3	
P��K��O�)ͫ�/��<�߈mZ���d��5�����e :ξ���:L
|���6��:�*+K�"�����T�<��ye~�<BE��~^M�vp"|����WO��U8s�ؓ�nѫ7�Z����-����z�K�햑�B3��[�<�3��L7%Q%��M>f)�Rf� [<dZ6� ���h��#�4ضU��F��D�h8����OU�m+�$����?�L���P���_������~l�y�:�n/@����{���<�TV��F)�8Of��˟�
��W���3d�g����(Ja�W|�r��Pdw��\:Y������z%A=ș�ʰ&�w˩�k E�H$t�{��W��0v]�6zԝ�v�\ع*g	Š�<9��	�,=�X�e�Vk��0�\/���	�J�Zʌ$���T��i�S��i�al%-'�o=��}vWq|�#��߅y�d��'/+�y���9���Y�01%K�fϊP�i�5)~9-iWT�!�$���N�]6��>D���F��oF���\w+�`�p�7��_:�x��͎�\��n��&P�'��L6��@��_ި@I"�}֮��
��P�61*�L�1���.|�e���x4 ����q��P�����V
�牴��q���l����oǎ�Q6�x@�����gx���/㼙�>��%��n�m�7�q����I��8z�Hx�`�L{�5U���G,e��?i�9FA��򗒯�i��b#OT��<n������W�Q0���&;������y�c�᠝r3��3�W?K�5��;��vT�Λ��,����)����q�_r��W�X�7K�MDOM�{�3/E��#��� 7��V�]��6=V����eo��k�#��To��X�Z�$�(֟�0�RC{!��G{��d���9
E�>����*��pF�r�.��SX0l�v͂B�/Љ��7���i.����W%����<�73N����gWS'4iCzi�Xi�.�m�玟@��I�Fv�7����m7&R�('�����5�yV��9
=��T�0�@J�U*��s��zU�.&���/�¦�:�d�P��`|������_�m��0E�M�!�q�y�:���,�X9�˩f���U�@H�1���l�:���>3߽bE��;�L/�L�7�R���N9�@M�~2����_���C(�x�����m�jH���擕$<іcn��K!Ց�B n�f=�b|`�f�f��`�VSU�sQ�O��{��b$��Ѓ$Ru�5��!q'j+�o@J��y�H�8�7�A��)����c2�\AS�!��}��������5��������t�P?��1��E�c��u��i����(�X�'���J�ŰvHV#�A� }����yTN��?3��c�R�����G#!�=���CD�f���������mIG�06Y�+T��\�IBU�Ft��t%� ���ç��d�>�4�e�m��09s���Q��ʢ�hѢ�J*S��''Gs/�n4W
�CT�����ݵ�F��BM� Zd��������&öqnVӭ�F���f&�N�l�~:���{�顡4�°�A�W5��Z��1ur��Fݥb�5n�#�4�pt�z�z���t��02��V��t���qb���nl�B�d������6�:fp�p�X�W�=
����>T��{��6�����D��]׬���q}#8��&�>�Ȥ��;Ҍ�vc���z쇫ݜ�,7�Y�u��_�8�Ц��~�x5��\�L墛U��y�� �sj;��ķ��P���}$2��o�{5�ON�򐰚��%w%ۙ��� ��I��oc�<Ȼ�i����#f�y՜��67E��-�dp���WK�{�Ԅ�%����E��%���u��[)�7F� �������+�Uw	��HJ�"�L��"��Ӻ�ܧ��)���v�����j��<=U����>*�|=���xi�"�~��
8�HZй˲��*u���(�(h����gf`D�1.�|
�ҷ�	�^"�>����k���sJu�z����E��U�MT%��0�p%��ι���5�|�LͶ�V�G��pܬ:�أ��`������)R� ��ר|[*�C�γ5[�Qₕ���Г�s���z���ZX��|Av�e��Yb�Y���ԑ{����:-�2������V��sb�,1;.��4y���e���5�3J����{S�*�Nd_oi�� Ҟ�*������"(ڐb�C�fB�,�,��nJ�x-c�jy��pݵ�Wlۯ����Ukw4F��F�j��X��&'���L(�[�Y�\ɓ[���Vf�5��9�����5JϤ|`��ګ��Ϛݶ��Ҩq���!2*
a���ם�LBL\�J�C%��8�΋&���U&�_[' ݄ B��N�j�,��ʲ�e'yb�p��V��yv7����۟3UGx��zY�y�.�m���wε���LTu�����~`b2A�ʀ�9�-c��i�>���wy^��H��/~�d��"J���r;dsa51���vM�]?Ț2B̢���:�oh
�T�4�TE����y�'gLJP�N��.�Ǵ�\Nj�~N�dJ�"��@�Er�5�k�<���֓x�\*om�2N�C�u��Ϟ�KX��$#D����I&l�����3ԁ͚�X*I�^�:v��X�0~���a�p�2���Z7���`�s��']��r��֟UDQ&��r ���e~�)��� U��i_�8d���B��S�]�/a��Uѩ��J��hlR�-�����^+��e@��M�SB!C�<ԭ/t	�{��.�Ŵ�|F�*l�I�f�t��j��e�\�\S����^��7�D��3����	|�1 ˕wTi�*&L���)h���-�U�ܡMIi��P�<T���Ym�aɢ�޽��p2n��R"h~��M�S=�m	���+���ͭ��˫�_T���6E�>:���p�6�|/��BRy��B����L���D�y��hJʘ�Y���)�������*�0��`B��t
�[F#X�EZ���}��Hc
4��0�[ⴳ-��{E�!mz*\ͺV��"�H�a��5�:�� �j2v�������S��uh�7�YV�Bo"��k(B��
X:�"���UJKEP-�g��4f}n�]H�Skj6�S��/V�
��Dr�ަ���ƌmn�*�uJ7�^Ë��ܔ��E]Qhi����;Ip
[�8A�G� s*�Mc���������{��N�6eՔ�J�+�Ćס���]�J�NC8Sk�p>�iv�������P�L�O�F�p`|]d��O�"ԗ��ii�U�z<Å�	Br��z	WK�ܳC�r���R� ���f�@{��dbkb]�!rP �G�|c��36s(� �����4�~n~�x �b�2d_h"<��f�s���[f�u����0�2�9�H��S)%�,t��G=��`��%�#:^��j^:��+�Gq�b2nXK���f_0�s���)�
1�&�+���2Q����E�y7`��P"����>���j$"X�1��﬊�0h&J�t��NG�^o��'q"ߡ���ᐾ�Y�#�%,���LD -��f\O�j��1�i��-d�f�x��Ɗ��qn!�Bs�.��o�$�9��In(Bv$�1݋;�-ik^��Q{��:��"ý�ޑ�� |��Og5F準���+�@�ITY������~�v��%C}{-�	��.a�e�|���Cvo��4!6%6	f��^���󊠸.t��I�8r�k�6+Y�Ԅ��%a�-�j=6�Ef��$��\n�
��N�t.	[��u2�-��M�(" 
���j�X1Ӽk<��w:�����fvq�X�0�����LK��U2.�Ȯ��wa%���w�݌e@D�9�UEL"扪] A?�s���/�"�`<�|�+Σ0	r�-�_rR���Q�R�x�iH�M`hH�Nt�1��P�iwm�+}$j ���a�� �6�Q�ą��E���3	�L���l	�}E�QS����V߀�=0���bV�Ak���[3w�no�&�.; �Z�y�LL��N�7 AB�I��e���Qxn��Cva��"�]����i@��,I�xK#w����U�J��p��4�������@Fyr'����竭�4p�жt%y�!�|ȃR���;w���p�@���$;(�M���@K2�\��Q���؋u�E^6m�v�Ǫ.��p{ږ��ODh��
a��nN�Kn0.�E	ɗ�FN.֖O�n>6�>u}�M��T�t�z����ԛ�d���M�Ȍ?���Qr�g�*�j�+�[�%�����晽������d^�7�l6��.�̘%y���*��~�� DB�'��X������ؙ�+�*x����Yjp1Em摤wKu�Q��x��^1�����(Y%$��msF���wq�o��v��9�U]Ii+�#\m�O�Ѹя��o�R6�<|��%���}#� c�/KHG�V��Z��6��u�NC^6"_�|b��0�y���:��3O�;�{E��]\�կs����A�I�yHg0Q�n���Ԭ0��s�<�"o@���
�L��_�z:8��{�3�8ϑ)�nHR�&��ΝQ�1x�6ۍ��:�����#K����4ge�/�qꋩhU������v�o��J>:8�[����6�;}QS4v��;������YT�P�w�v2o���e�L�2J��0$�uu�q�OF��ن�,
 _�9>��n�8q�,?#Y�u�<�U�j���4����Z$�!�����ds������+0Jot{_]� �F��bo�Z�����2EL�HsF��8(�0� ]
���D���r:�b�mev5�죍�Υ\�)������^!zKP���8K��e��h��J�S�l��/5�p�i9ռµ�u���R�v�i�2�P?�L�e�
~��APwH�����Ƈf�u5�@+�]y�p�?|#����~����"#O����C ��t���^��a�љ7��c=V�T�+7�	��}����dK4q��,�o�|���J.��0�����>ì��38�
X#���^�`L�mm���_A��^X�yzUK���Ǯ9f�/��`��B�&��1����G��a��Rh�H�;�3�c��7N�	>!�g�x竴���ܔE������>�*Ş��ƍQ�K�n�w���U�0$��z��$X,��<�,��ju��(��i�P2�W�����܇~:���v)���G�C�̞
�m\s���"㈨�Ո;c:���iw�������rJj�&'����}v��ځ��"�L⪵O
e�����C�����Zv4^4ԗ�S��yE"�̕u���ǳ���]����V��>7Zqs���ʾ�,�SY8p����s��N��i�z(�,"pX-���H`�h�%�O�Ӻ���֚%�}8�ĳ.ŕȲ˞`���O��9�
�a�ASw_'�GKKW=�M��[�|0R{��6� kg\-���.;xE�i_oY�2j��c��^(q3|��J�;s�8Y���{MJ}.�]��<���ss�q�:;���:�
�M!��n\F!7�J��Q�P@����\QmM�o�1�%[�o9��Up�[�H"�&CQ�;	_���K�e�#��Ikl͹x�^[]�o\G.3b��9<��Hd�t�żNۜ4_tBp�R1������ku>�q͖\3��CN�4��\��VЪ�a`�B9D`���>���&s}׺Z�Jo5}�9�m$��������8F��"u(�@j|+�*]�ͼ�w���� ������{v����0Ĝ�4[���?����&^��"�~
����@I6"������@���&��Kl�:FB��u��=�s܍v�)fTG���қU���y4PV��;�e�Q��i��Ұ{T}O��T#Vh�U/�9[���>��`�ɕ��D_ꦎ������I��I_�2c��Xg����D��pI�<F�S(L8R�q:K <c�E]ܛ�B�w�4~u�	v[�!���b��`Oԅ��MWf��~\P!��/�I�t�k�ܐ�y�Ѳ�����{��Rl>E^�M��Z���9���,���K@����b��B�B�^�#�&yy!,�w`X�p��m*5�t�H�W��D~]�/{�@]���U���tO&`�����M�$�h����/U��e�GSC�z )e��� �)n���U�\�B����(�JKE,4y�a��=�5j���VpC�R����9H{���/p�T!���ڮ�a�2X��$1�(Pv�4�%��u��ح	_����g�iܔy�@�ǜ������/�6X�.�<��)�ǡ��v�?��ȍ�Q��y^����8��鞐�K�=�BI�?��E��z�!�s�}5[`+��|�8 I٧�1����r��B������\�3�g���3�X�b`��u/'ՠ1l�{e�1�u�'v�d�;�^�t�]�ڏ�W�ٲ<���i�l���2�`�݄����G#�x�o��G�uz�w�>�C��Hث�~}��1G,͒����w�	��L���;���H ���W�+Hh7�������gB�����9�{2&ͱAX�Tc3��y Z=#L�S��"kj���/q�A�%dWN*e��|�+���	�f�uiu�������ͣJn�BuGA����ۄ���T[�4���!J1���%EO*L�d(>q�a���t�c~Pޏ(�B�a�o���	�0ᄄ����#�fY��uD�:� ��n9_e`��4�l9-3H$E�J�7��,��� j���6�!e��"U�Sy�9�U��^��n�I��xpR��ې��>�ϩ	��"��R�; ��)3h��çN��oX�X����,6��<LqC�8;�6:�g�N�#	�$�M��/P�T�Z����h�wI�K6��Wh��7�����E(�Y�o�e&��������iR�|<R�,�/�������xS�d�8m�+ؗ�`�m�)M�hsE�չAP�+U�����{�t���$�C����9��>������)�f�Q���'ޭ��r_h��\�����ޡ}�J�VӋ�N,(��<��׏�=y�|'=1�ɒGβ�4k�=�\I�9��n#���b^@\Sp���~VFm#��ޓ���e�MR�*�k��W��廫��	��	bٵ7���Ix����e9���Η�%;쑿Q�ȍ��P�Q+t���^����ʉ��{�p��4h�|�g0g5
X �b;g��&�|���m���{eh*D�ͺK��I��e�PY�j�Leq�((+�/�G=W�$6�4�3���[�;�n�XA�O����?���ִڳ�^��z�؆&��db��^D�p��}�,���2����n(�M���7Gvu���h�>�!��Е��
?���uEqm(�i�T��y�kC^*���.`[���ly%C�:�"Yk�n�p��a$����)�����tӸ����~o���T�?p��Hg�PZ � �am����9�R�U,W%{�u��a�&U��>��O<>2��?�X��'�]�����%�)ª��e���O�� W�x&�!�~1�u���RV��@|l��l���&"�J��ZK]�4�A�	�d��;eX
g3�z��4, ;sޜ��%�#�����J���'kcIH��k�bAP�Uai8B�Y�R�����ǖ���\�şK��	�Q�VI�$!0�� ��dJ�E���u�2�I� �pZ������Im�׸4�m#�H��y�In�i��]�V��
I�J��p��Vބ2;�P�U�?�man�I��H��|�D�#�M����/5*FN�a�}t2�w'O�f��\)w,�_t$!��/�Be���j��ŏ�iDˋ�]m�z�̹�A������kZ�+9̈́����ck^�T�C]����2�3 �%)��~�s�m��S.�����N�i��\t�W�4� H췞����:6��m(�����JkHl��>��L��W�J�e�F��50�_�jǽ�f��t��7��^��33� �a�����ZRf��d�8B�,ˢ�U��CC�&�63����0��ς�G �I�����k��٢����U��@���}�K-9��n��K��@��"���C-̅�$�g�u
"
��/����-ьl�/cˬ/i�Q�u��6%l"v������2"����5s�t7�Z�]9j�9�{}�$�-�J}7aq9���_�C�>�[r��p(%Y"�n�k
���;���S)�qp��b��&Ͽ�u&���m��Z���j$zNp~�����EI��9�h��؛������������pq�.�f��uX���f��}�y�����~9����;���(�c1m/�jōv/\�7��h��b��7}�U��*�0ib��v-l��Q�B��k�n��u&�X>��Q�D1*Z
�*�=Sa�z���]ޅ0�v�	6��L7Gt�f1-�9�W/�>�d.5w�&��?^����w��d/�u�������<��l� ����i�%��d�ܓ[��Z+�'�$���x�!��8�|����>l�n��=to������{=R�"U�s��*
:& 罍���.d�6�.����}��EMZ�uT`�r.'l���a�� �&�֤)]>Wk�F�~��"�#�N�X;���1�0z`=򸔑7�!��4�!c����0�&N6��▘X����s�h�W-on�8���(��=�O���3%�e^�Z��[lc�W��>,V�ާ��W�g����1��x��K@�u�J�LkWܘs_���v��_�����|/1>Cܨp�9�\B�s�hW�-��jd�pԨ�,kj3X�����
��X��?���4��}I�?*�����s#����@���a+m-��W<C8�)p���q��T�o�����
�ofנm���gX�&�Z�8f?�V�y"&��_�K?��a�pi?����im��;�n�FG���NtLua LԵ��lN�qC����4<�yȕyK�=���[gk��L�z@>B�F�ʱ�r���d��r�E0y�옯��������Y:���!���|.t:^�H��je��$�Ǩf�Y`@4�����ݸ.m���%={�(���ԙ�D�cN,�����I�~<Ƨ����s �l�!�J�O<qR��j;��3&˳E҉�l��۬�${.7�lF�[Q��4g`�v)�)	-�,�_�~60����Y �4���Ơ�=2�M>���+-�Ka��Ps���GpXBJx80�)��F��?9��r_ʼ`�W�l�0�jd�n���b�`����'|�s�ؘ��#?�jM�.;�`�^�����1�>%��n U�.��_�YgiN"���"ĵ^��dA�bȫ�e��]�eq�	@��XC���b� ���^	�g��Bya�'���l����6�����p��jzk�IG�"��F�!I��1�|Q���pq�����`CU+`:��惋��*l�M����D����>bSx�j%}ϵ��0
������6��O\���GVf��$v�>Y��Ͻ�B@���L�LnQk�Id9ܑ��X��{G�cq�l�l����bRM�����]���`�1�U�+��"�z����%!Jb��_�0����Ǿ��?��Q���/���������Hz�yQ_�ڧM�i�:�5�*A@�o�	�{�DS����^ˮ�t���"��NR�/YR��[ɉ�II�>A��}/����El�v�4�� }�dnB��|*�%�c����P�r5�ݕ�b@H[>t��������(ԛe4W��ŘgI�:��H�����3�Q�Gk;�WQ��y�C���.�r�h����Am����+6Z�
g���}e�p�r��a2ùg�)۵ \�����YD���O<)��9�0 A�gjs�GB���Mxs���b[,���p��n��ᒎ��ʨg��tg�RJ`3q�;n/+�Ăw�� �M�@���_�op�ǝ'Oh�8�	ۖ���*���#]B<(���B��J����`/"��>[�3\%�E7|�NB0��y�mD��}J�w�k[�k;�aIPW;�G�_GV��쟟�?75%L�G�bQ�q�%+}h.-���$�*?{�㪒&D��Z����*����uY
�:� o�d$�b3`��ݛUx *��`�"��xW7 �]��A�s��|?0���_0��!��\Gv��v�<�=l���+| �ӿ��ۛ�ˎx��������ʫ���V�ф��t�ILե�Ï�:�K�َ��u6S�%_Ѐ���8t_����S&K���E�Ӻ�j4��ɉC����N���u6��IWo=KB�H�J"����z�
U��\x���I2�N� S���L��F���BK��-�+B�F�=���[�9����<�g�b��LPg�vjvcԝC�׾Y�S�j���
��B��.�^��I�ӦL����y�����qE?c��"�*�{NS���4d*7����h�υ�U���
�&������n�M��k����'6�6�U
��~3�ϕ%�Q>��&���EO�<yj�\_;�7>�d+_���{I��"�o�G�
�"+܍W��O}����U�趔urm�a�W5w��5�S����o
�z��E�D;%�j�H,��O��uڬ!
ģ�r������m}�ni��o�@��Js�Q曼ϑƐ�:k:���Pw^���9vJ8����VZ��L��M�@jC���ULyIO��o<�I�
��P���t!�&��������(4�B�w~i����kW��dMC�H�!)?���T1�A"F���-c�zb\�ǫ�Ew%�~�y�ހ�]��	'�_Qt�xc�_d!�>����e�zϞ���J�k"�p�5"��x�&{�d�"Z�}�����!�	w�f���s�Ö���ŗ�Z�Y7L�&_i\VQ�sf�^�9��ԁ���S�6 rhom�c��ޭ�|���M�MV{�l)�"��]�0E���G�ι�O�\=�?a���Rʢ|�)�Џ�"��!ɩ8���͓���?�/�=鷛�/R*~��o�]>�t3#@���,�^Rf[���wr=d� �2G����� �8d#�8���;^�z�3(��,��?�"���T�F��7$j�ymTT5�%����T� �Z{;ˮ��(��?Y6BS	#�}��邎B W�������WB������kT���>����Y�Y�|;�}G��8� [Uyi?ST�_��Gyپ���v��f�!����J�#Rg?o�-9�.ُ�L}��4J����)V���O`���������D�QD�!��n�R��9��2Y�=ܙlDI�gw��l'�d���>�m/:E�!h�N�灻��&���6������ݔ
�/ ]�G�'�d&5��˩�ʺ���8s��ދ8�?��p9\&e$�-�X�O�N<_��Z�s��7?� @�([?T>V�XIS\a��)rr9��g��ܬ3��r��`%@��P�GwV7>����a�^И�Y0�c ��6�����u����#��L�)K2���p��3��7�s8�t�c�7�d�|�}gY��b��{��4�	�|���9Z��&�J�C�o�#��.x���P�dZ� �ܝ���uB/��`/F��܌z?����#J!��`|�AwN$vk��/��J��K<ݰ�w��}�ܜ��!ŊPJDr�Ѝ{�k��-J�F�/�}ur�z�Q?��3�� ��,�NTcIR�U����<5}z_�wY(~������-���=��L!���J���Μ�������B�0�$�\@:���C�7��E�G�Rױ�l�3��c��^���F��!���рD����h�� 	2�PD٣�Na9���7��p�����ҚQ����yū�v�!DU�_X��z�^
f�rq*�7��*���;i=ѦY�o��d�=�8Q�y�g+lv�2��!�Wx���b���4��Ň3�HG��{��R7x��4��]B�����`�m�!W����<74��FO¿�@ʅ<d\ �k�s?�p���d���*���oi�T�)��A��%RspW�8�B����Q�����sG�Nah~@V�m��`��J�5o�jk� �XG.!��i��c�(�m��g�<&l�_��?�'�q6U$��+�؄��qt���`�]�t�U�"t��jv	��]s���f�/~/\�%_����#���w���ZR��)�m�7)�a�H�nC@�i�?H�F����Ӛ�}�g�ھ�o y=� ��C����UV5��0�;"� ��d/�փ��# �lm�b��-�K�(���Ѥ�@$��:|�Î#%�S9T���� ��V˅x)��hȳ>��`�wß�VI���ȵ��P��������k�b]�L�����c��ֻkTx��V�<�-��d�U��>|I�M� S�.�/l�.��:�}w<i�ի�t ��o��Z�b	c=j]]bs��`���X�.��`��-�<!LJ�.����Dp��ǜ�S���Y�M���h�o�[&R�u/7c$v�� �\�S���S��i�h3�� ��d��)l$�h2�f��)��+ZĎ��D�ox�*nk
��^(�ު��Q�}�u��ܘ�z��氤��Z�Kia	�\�{���6�}̷���X�X�L�+�!���B������!��v:�2��Tk_΍��t�GN��4$����%v�VbZ<=�*�J�~S�q�BuJ�e���1��匬��;$>����$A�E�X ���_]�nd��>z8p��i神;�1HN��]O�w�g��z��f��}�ҶZ���[��=d>���X{ɔ���?2z%y�e�A zqǆ��,Hx��,��4�\�$qQJ0��(D@),�`��wwp~R�Ѓ��2�!K�������
�I1�|���{�:�ܻ	��[�+G�wg��� �ȩ<TT�O�n��"�H�ڪ����#�ж�1	�%�?P�T6�	�4������K=0���������$�`��B8/��0dZ��+��	9�ܘ5�%1&�{��k�;��1�/�m�������$F:s��\��y[�dY��ʸN[��(�%r��5��m)n;�k�ܠGy�� 9�T9s�o��,�sR��u����օN�[�r��!-1���WA��������c6��86zL-�*�&:Z<�3E�u�W!�(��I���Q�<�B��wmb��R��o��	Z����l$�A�ё��%��9W ��教Z�d�h�.z3I�8�iK�9I�����
{�\���,��gà�,��p
� N�w�l&�1�#8�C&��k͝�.��QO`hQ��b!ſJfz�d�{b>)��mB�>6��.�Gu�q��-Њ�/[ ב�s��<~���>$\���İ��D`;���?S��-z��!��p�>1�Qz�C��Q�����ͺqn�'�$e��Xi���K��ȟ�Z�K�Dg�
}�r	>�g��q��?�͇o)��ˇ`*'-��a( �X�'1i69��� @Y��%��4 C���˫��7Ċ�tp���)�a�b፻K�S%i�Ԕ✅��(���NB��!o���������шZ������c?n�����)N��g'�ə���=�w�j,^:el}�Gp�1,��BØfZ�)�&�v�����;:B3m�����9�~���z ��:g(`�k�
/jD�I�duf��w3�=�c���)���c�Է�LD�c�yה�#;����p���-�7~�Ԕ:���Y�/S�L&o��SjF;�f�n�뢞��Ue�_oo?�hє�<����^��u���T+޵�Ҏo= �bp�
k��b��eKFh��Z��T��R����$���#�J�gn�������E#�d
8y�Rb�,��u��|��D���dD����]��M[w��j�j�5�cm*�����l6���:���7��H�ێKV��q���M�o�O< < ��to���R���N�)+��֤�P�5i���96��y�[!�OI�y?'ɪVLL�/Q����F��
A�4J�`��Icz�Wv#�đލ���6)29�M�$,b\���c�`	�4���2�E��uZ����x1��;�tX��Wi�0����T��m�/�~&&���f=��P���+�0pAf��'�N�ش����X݂=��9$0/�g˚��B���K���-�i~#u��'|d�vһ��6���|֎
�$@�vkja�N"��[bJ���7�i�>!�o^����@��R�Y)��~��1�ȩڳ�A$2�.�m�9?�5�Ѐp�Y��*d�P���DĮ-'���Υ���Q����{*��	�g��~�x� ��O�H��?�^�$6��S����x�����[f��0k�^B�UL��$N�SP긿 �ڝ��w;��^�~�=���)~F�w�M{/�)
<�o�r%~�u����t>��r��{����b����$A_��nM`b�yEw�� W�E]�W�mK��r��ؿ��DT���7���8g�W.E��� �,�d��!*�H	l �i�6�3���K�~X%�����0�r~ד\�^�ok�˔�����>�RЈ[br9�V����������~����?���G���*�˩왞� �9��T��V�[��� ��y~2A)^�B��j�_g�xVb��c�Yk��@"�+������1g0�{�Y��=T�Z`�;e��u]�;�_���Ѷ��3Qy
F�2�6���W��}�Dn��-����G%�A	~^�5;��w��1W*OzvV>� G��@S��I)����z�0�"���黹aR��Hn�Sj��$1�bI>���dw�ŕ��O�ڀ�"G�{�k)�﷥��Ho��|�"�=kt%���E�*��0��%o]�k#��)�_B`[����!�F?�W;���I�z���B���D��5t#���6 e��?��%J2F�M�Eu�\�BВ�b}�9F5�q�kA�0/����5U*R>�3���(אP���<h$��Y�nyB���S�����D�D2��x�9�����;��0�NZ}Of�N�#�4<W�%��|�x�ɻ�U�c��Џ��1�41u?����Ɇ��{����R�PIoT�3��m<-��0z�4�GkQ�L_��� �������cf8,Z-��"T�f����#� ���ͤ˔C�=�찞�l/��dI�t{���?����r�-�üD<1Z@VI��O}��1�؇�"��o������r>w�9����Fe���%�ήXn�RC��q� ����E��8���^�\1O��8��{1�PܾA��J�� ѩ	�����g��� ~�����*�%��I���7��eg�5�T3�^k�G8���nNq3q����P��8���n����}�`������=*�_qn(�m���u��sG�����С�ۀ�f3?��v>>��f���Q���V��M$K�5���M���-�{�g���p���ڴ�y�ƽ���!�^��Y�}�C�j�.`h�հ��b�-���r�����k��0�R��b0g��_S!�1H�?�%�Q�,�hj6���3�@�!h��]PY��G-�R��k�f耛�r��ҚB��7����zB`�J9©�m��Y�V`�"XpB@��<D��{iN���z7��rX�������6�O�Q�gH=����9�ߖ���c���j�'@�����Po9��ƒ���yqX��.�2[q�:�S��H6GR�����	����m�IH:�yVÃ�;�e1��U8#*��H��oT"�c[4d��"�	���*���ăf3%���&o�Z�I�G�F�������9=�O	TǱ}�^L�L��&@�4����](v�=)����:��_�m��i.9��kH�$�2�r��'��#%���r��Ugꄻ[9��I��30�+Ԟ�ӔB$2 ��z�MSh�y��>������ ]94��M&��79�ASD���.dο��.��4������	����O�D� v��{Q���2�fKJ�r���򭝽E�����
Ec/,>��/n�;��s�&{瓚	o�i�J��w�m�����ys��H'��W-4ڧт���V]6QHmL,�Q��R��&;�M'�q@�D�O�
z:����h����A���i0�d���zU	dStsa����Jڤ��M
+�����e�x�{y��rEE����&�,�+�]r��e�x~\}!-��'�=���E����h}�!����Cv�(JޙN}f��ź;��SM�{�/T�E���+G$����v|��X�/Q��z�CJ�<��'D�x�W��%c ro�����|9B	u �є�.��� �(�S\��LF&�}���b�ӧy�2z@�'6@"�H���眬g�a�����>�X_�)��^=��?M�>`�l�ow�-kD��|����TM�Q�2IHqZ�&y����<�� ��gɚ�E��r��1��n�E�x	��bZ��X�9��u�_���	���6:#	�*�w�2�D����vJ�e�P��Z�g�[/�8E��x�&���a���~_�й��S�M:hn�s	h����hJۅ'���c���_�|x�j��geb���;]���(��ypg����<mV��6�ix�Tͤ�#-�0V]��-%�I�*�@$�#�1�h��G6�F�ox3F�:x1^����t�����GP�\���N>O�`+!8�s\���M��8�uㄔ�Q�����1sp+�P�hX�9��T�v�~H[p�@����H���鬘���
���>hw;A��E�g/��A�g,�;M�́bx�jS�X<NۿJ��Hj�&������]":+�
���_�x�\��]�Px�R	rT��Ws�{[�Ny��Um'����3
V�܍%q��Ʒ���mTމ�" ?�7�n2M�AhJj�9~�jz8c1b"A;)׆n�ly���q�?�� ��%�$�����-h�N�KGбsؕA�DdF;�]Z.d59Έ++]���|?�$����ִ�� ��o�� ��$��8
��R�i͐���W��/���qXߞ0*1#J�\�R���������%��aړ2#��tQ4:�^�ü-F�տ�$nV��9�_:��kֳ`�@{��3�9U��H��$����-���h��?��ɡ>�/0��ւ�s���,��@������b������Л���EL���A�)/Џ�ݖ�Б��JЁ��"#����yM�4���~��8�
,%��/!��v��mpި1���:�Z[p΋u��}�i�P��VT]L����ղz5Ȉ��O#n�a�!��U��o�;v�Q��W�l�M�72�5%G��ZvvM���F�T/u�xG�Lu���z ���u�����h�W��bT�Xr��
�hTK��כ��+9i� ͆����ϑ��#��=ۘ�r�{k�Gc� �y��E�N �Z�YE��20���k^]Y�O�Âc?v�nF|&K�vs�~�2�0ݾ�5�b��	��t�w�*`9��Pp�	�g�S{:��xJ@s\˗�\0ħ�K���P��߉�I�nOL�5�wp<�3kݟ�3>��ӵ6�����,W��[|�6eZ��f�ޤ���b�D������M���b#�\\Fi}��خ<���c�������z����zo��ͭD�J������Y���W�m S%S��Yqo��kmPOnx#����mS|�f��̱Vիh2�C�B�����g�D�Gi��#"KRIsn&�܊�g80�;9��Ă��,�,�?>t}��X�v��g��
��"`q�3���x%�%o�<3�WL�t;�e���ō:�?Ԋ�C6-��v�,
T�f�Y������}�EWH]2��5��q0+J����8�Iy�[K� t�0�4��!�,����J� ;���kmy�w�1����d��KQr���lc��F�G����G�T!�(��A��on�ҹ.F�K�xO>aǠ�}�[���QU���s�Nm��ȾQ�bdv��dڅ	��Bw��4�&��~$h���c�ΗQۯS_�I*�@��_���\C��Q�k��-�zi+QGk�d�p=��)��A�*���<el=��E��
�{�Ԋ�!F��A�H�=�`�#K�6��ܙ��{�)]��Hr���S~�dژ��͗���$�i�@��X��q;�)��M�Zz<�7	�����vY��$�3/���?���Ţ�	�/�U�[ΐ�,\E�RW�}�r��䪧S��.�S�]�`KD(J�E棞�6XqK�p�jHF��%*m�@���� >����	�f�z����,�T>�}�}梗��P?u�1pa�׺?#��D��^���iW�����>����'�Z kMÿ����Qd����g�e��ë��X���-)u�/�z���Uв��ck!��RH{��v��;D�n�V��-�ۜ5�>Isw�t1��n7!��ҵp|N������;�g���N����:�&�-��"��<�
����W$ɛ�;�5ի���҂q�-x�7����v����;��T�28�)x�r�,=�e���g�H�id���� "����u�*��]<@`���]���@b��j�ݏGڌÙ\J�£���߶�\�k�l,<���e:�s�h�tM��_� 8�dx�N#�\��(1mJ
�j
1t�$��P��Vv9h��h���˭�|v�!8��d�E�w�S�;��¬�xO_��!0�#�G���@�e>�_�j��to����7���U;X�(�a��X,�����l{��o']�8p�\"nz��x5(n�0*韍E׈P��M���	����:bЌo&ց3�m�x-�^ �2տ���`ī~���W�z=DC!W�[��'�7��y,��t�)�;ǰ�y���@=��jF��~vɫ6*��>����^���7{ �I$K :��9$�[Ç������C��4(&e&b�J�xG�'7`rM�<$U~*��|�`&~��7
��"rL�݋���枤����1){�7>r�2��!C+.�_�����d�TWi���c6LD se
	�5�wc	d.�%��e�ϸ 233���O-�X��5���7}H!? �91>^����]e=��be��Q)��U��y�ڬ���5r)�p ���Ћ��MNз�[�	/�D�W� �]�:��A%�Jp�BfRC�_!��B..9��aqy=
�g��-����ʦ�gV��7o᳥KNh�����j�{4��o�����[A���
-A�4%��B䊛}�-�������{�϶��.q0��-��r��5Tȸ�4�7��E_y� q�!��l �f`S[����������v�B<
�{6��*bl�;�8~�0;6ٚ5͕��A4u��~���QZ���u�5�iH>���[�� �G �����l�r����k�u��?��ƬY̻�m���	��]ܚכ���t����A�+��w����$��qU4��qC��<�E3:��.��+`�/��</n?j��p`HM��_��=j�k[	P]ŷ��J��G�t��18�-��S/��K��B�F|���в�.��&T���+�1�1����1��W#��æ.m�7T٠�c���"{K#�M$X1�}w�������܄z`Nĺv�2J~�?(�W���?�qY/nL��9(K0�o\����&��d����:�=yB��j�S����N�i��D���z���Tw�B������o[�:ѦeǞ)�����nC�|P#�c�=|e�D��$-ǎ}��/��}�����J@��cldt���FW�_}�(�r$RoXL\��UW���γU~?�l����f�{��`��0G����v�5��\cp� G��&��f$"�����#8}�������I�Z�ě�sS�)��j���A�>
��N�Kv�Y����e�@�hs�x�N��*���6/��M�����:�t�Ւ����b�hM_mч�F�iey�n�Z���b#2��b���e�t'v�]	��U�i5���� �Ah{�^ŒV��s&[�a����n�m����l��9�
~Z4��RF-�/����oOJ��̓w���d����M*�3�R��
^����c���'"h�dT�#���ܟ�Z���N�V���`�v}Zқ=���>�B�#�h��6}���/9b��I]�;�ݺ�]-��Ǯ�fR��N`���oMB�[!
�9��w�h��|r���WO�G2�n,�A��~�6�wm@c�l�[������׌�?�ڱ
�DKB9[M��;Nn�>ޅyk:��(�5�B����[O�֕�sA��l���a`�S*,#T���r�M\��|d<l��w�E�&u5�؋�%�j�{a�0b]#'?±F�J�D�TH��eO-J��E8h�����z�j�|,��WIm��o{5���ُHCDs�X�u���OR��(�N_��|o�A��35�?I+m����Z�'�%��'\� ����U��"~݋{������x�ݫ}}�(���zLi;���Ľ���z.g���?�yjH<�Ց�"ϱ�)6/Qǜ���ؗ?읤>ՙH��:��jz���� iKgq�ƎpK������4$�P��8��5�60#����	�dZ��ɚS]����i�+��n맿�q�Ɋ�8�(5�_���!F�~
��!O[� v[$�®/��/���˓�lu�����aQ��+=��+s7k��yl�B�7Z��>Nx�jg*(NHc��-�zz�YW������4Ў�P1`B��ʕ����>G48��0�)�zC�&�OF7u1\�BHF��y��\�#L�� �(d:�\^Q�xH�e�u5�{�i�<�ؼlh�j����4f#��-,�l�L����������G�\E�[���'�
�+�hd��pg�%���2�˿�yy���� �	[�P9k�}�"���b�J��(�a�R�a�BM�54��`5��x�h���	�N�y���Ƥ�a k���d̀��q��74��
ּ{�����-�{W�8IL�@��br�rp���d��K����4�o.NЭ�zo*�oJ-�	�Z7�.��$�XW����1s�or/c�O|��"���-h��	۰�Y�v�A!��4N�����:�D���o`S}���y��i ���/
[j�Y��/�[�JKO��ם^C�˃�<M�HE��\I��
����+�t�~8�)(�#M��,4�S<��M��';�d7.X����H~w�/j����2t�h�UȒ�(k?�X. "���	�r�Ljj�����T��mV�_�M7���L� c��.�2�5�x7Z�1<�T<�	��qd�f�6d.����W�ii�9������ᥟZMw�	,,o`����d':*�W"I��/7�������s�.i���		U(/1��u�
uIl�_wA�}�X[uU��)Y�7��jgp����Z��  5z"�u�&��mƊ�8Hj�P��{�ﺰ�f�C�l�Z%���'[AzK�&�7Vl*�u]�&��#�r[#l<ԃ�Nꯎ��$��EՌs������"����`�oM����@���XnmH2��rԹ��3����K!�y���
��Vo�<>u��Zݔ[F�{Ѽg��O����|�#f��u�ɆW�5���<��{Y4D�}��Z�چR��-<v�JF���
��`�*�>����r�gJT[8���em�Ǝ���s���c&�(Fsir��E��څY�7>��_��V�Y��Y=�����-��F�*^�k��������-:ri��կ�
�Y�4=ԕ������ &�F|��5	>���!��#��6��+�T��G�K�/?lb���r�]�bR{1D,��?;�ɲ)�#��S��[q�,n\|
^�o�o�O0�b��.��LV!"-�|��"[X�)�C>����e�e/m������{�c���{��s�mɗl|��y�2����`�[R�ǔ�GI?����&�*�==_�w[�.�~rCb������<���䗒�������ɬؕ�\?��a����`Sی>%fޟ(���1H�OH�~i�BZ�[P�:�	AG�Z�����u4	:N�K�F"��d�p��U�Y�C��̺��4��4@-$-�۟X%�Nv��'-���P��׌��h�+����L�z/�w��%��|�H]�F���h��w��nrc����r����S����E�:D|_m���go2�0�nh�C�0&#���tO�;'r>�����fT�ܨ��;�H���
���^�,7�/�O*�<����}k�2��D�۷�U��6�$��s\p�M(n6���J�Dm+w^�*`z�!\��5�U'f�������Ы��@�.'��3�� 4Len�׷���V�O�H�C�o��G�0��S�n��. ܩEaQ<�����/F ��P ���y������RNʝ9�܋�7�hC��9���ɢ���	�b�p�Yև�� ?�Y��d��ޘtqo�-�L;xC��O��D�%��ў����l��n{�3���=?�6j)��y�*F���;�T1��&t�^�f�}��U�pJ��4�e)ȱA��L�ْ�xK��D�Iۣ�9v�H��T!vY�#��IUi��<��L�^XF>�P�cxQ��L=��&���1v�A�8��z� �Fe@�|�u�F1��l�b�&�ʫ�˃W
(��?�W}"�#(��/ c�u՚.�O!�J,�x�ggT���R��$��n�q)�8�B�ӿv�k��1������]��5���I$��D����?���s�ޞ�Td�]{pܥ!��k�\�C�Pe3Z���>��j�<4��7e�/�0� __w���� �7��j�WY����l� }����
���bä�<�7sHi˾9�g�9�{������p�Q�^ɳMf��&8��m�mX�� x��iKn�R�ȡ��޽>��R��9U���W���X�*Y�oҕ��?��!�<�x�f�*(��K���i���>[L��N�FQ5ࠆ���w��n�<j"C��_��6:��D��8�(5�j&K:*p=ޞ3�J���p(�r6hB�uV��(gb_�C���ڎ�\o����$�������(#(�7/45`���B���8`~_[��<Vf��n�{�qg(*J���q��gX�3�Ij_��nVw`]l]�n+�a!D�R)��2M�ezY�y�걭,�����&��]3 ����[������Jݙq��s�&����M�~�S4$�ވ���i�Ƣ��Ohg�%<��5��)E��̠,���K�B%�-���㹤z��[����|-����$~�KzQ0G�-�,�O�%�h���!�������	xh��Q���zN3�t��^ ���O����׏�g|/XA�_b��%���E�!�D`G��l\
�`����?y��0���sE��tbv�(2~s�aTz)��C��!%��x\Х-�e*B|e} l��UQ�����Y��]C�� �l�r�K[��y�1�8Nw�=���	�����l�Q>E�E+�Oq<ڭ�?c�m�f��i��Y:K�s��Τyjv�X����$��p������Bb�w�z������0ݠU�x��/����-rT���+�?h��~���r&��7��rsݍ����>��D�=�����ĵ7��3��}�(���Q���7�\�ѼYPN�&��,�� I���`L�)r0sw�?�Q��g�q��r.'��o��c���k�l>X��M�OBA��;�> �Br��
��!�an�����ܪ8ܽ2.��k�wg��LU�O-�d^Z�f�#ֶ�tڊ�*e��k�M�%�Hh���81�BM�"c����BCIoI��"���4��r����%������y�Hʠ@�:HJ�Fv���T�Ă{?S=�B���I]���g��ek���h75@T�G���N��x��v{F�#�n� �i�H��Gl���hTh��)7#���<Ɩ{���soa��*=�^���.�u������}����ض�&5�X���u����v�w\\�tP 3�\����Da�v��i�+	�-'��������Q�]?\aRۺ=�/ǻ�v銺��?�w�����f�9�)���������v�&b��jY�.�ȝ�����8�"���7�|F>&���)�������1�4��
ٶ��g��tc�����]�V��sT��^�n���N&[�f�Y�o��԰wd�~A��,N+o-1��������~݆�tS?C�p�\�M`�+6�8����Վ/��.�vޱL�?��/��W���sԧs'���:��0��NPa+��|��5c9���Bh��w �H��;y�W^ ��)J�����.<�M����W����=��K�O���*��[̻MB�Db���A,vlНf6R��>����-hމJ$֎����u8��"����]�u|j��R̽鼱ywv"n�s���+�jV��+���������]�4&���q�ic�T�ٲ��X�s����W��R���)�ݕMo���b�N=Dz�a��>G�ZD.�{���]Y��fUv	�#沀58GQ�ʎhj7�֘�sV9�y����,���)Ф[���1��� RKH��!�Ż�z����Xd���f5^�~rm�g�N�� J���B6Iv(h9%������'W3��I�`���Z+�<v!��#A��5����ŕƷe����=-�2�#�g��^g��s�̢��`��&x�7NM���o2J�t+�����J�B����@�rj{�d����1��ɘEYh�C�T�f/����r(��JU�fb��N����Ǐ�g?��;����C5�)n#�(-4#�ޖ,�a_f��i{�����={�.u���1{��2��WI�,����/��X�n�F�:-�(5���
���:o�b1�3�9vE(���G�``���������3�v2�� �ؙ��G��߹�3>LW�7@qo�Enφ��]��v��Q�gY=�=R���+��
*�eΔM���v|�4jC���7��t� ѽ�`{�*�a��1�Z*L%���=\T�ZkH����u�P)�Y�m�����HZ�{����k�� ɊOF�q�EG���م�g-0���x������.ZՀf�ƽ���n�I�)G�a��,�X>��j�6��7���q��Mvwj�uOd�[�l�G�"���V{	7?�h�D��(>䜤�$���W7� b��Z�]��=H��}����w�Td�p&��!�����T]���Kc��݇p��K�p�W��n�����#b�]߿s�a��*��:��@?�
�HJ�!r�����l���(�\ڽ��1l�[<��}t����F^�!I��X��� ט��hJ�3񈱤K2T];��4���}������� �#9B���,T:�lI"�1r�m��"I�Q�p���k4�Z��@�x�N�No'Ƚ�#���J�sf��6L�e�aQ/�\#����G��l˺��K���v�&e�%>V!�@�a J�Өy=�;s��	+ ֟�ޡ�~M
8E�� p1�f�����$���<6�x�AY]��-��:\;z����S��#����o�»�;|�~�wu��=	j$no���#�/r: ș�p�®�zI�"+^����(ݠ��.�*��t�]Rj�I� �;����	�R�mi�N�>���[���ew�3�k���Pp����x�fN\�C+.�v�A1�� �kRz�#ga�}�^��g�ED!��ef9��З�b�p����g`��z�i�7�҉�YF��C�����x�1�,{ld����@�����Rp���=x��M.\W�4T�����pwa����+7:,|����@��E���Z|S��w�<z��C���@;k�{��k��~����"> ���=�����	��j�^�'s\�Ə������E��Nۓ�t(�λl���2>n��ހ�~��9�s��<|B>`�j��ho�#I����^S���^|[�a�Q;����g��T�o{Et���L&";�^�)�i9�wV�����Z?.��/������x�Ye�m�+�)|=̓���'�)����i���G�,#;����w�n�4z7^���t����zt��/5�^N�����vv�:��~�
Qߞ�����^cmg�q����`6!{V.�{'>_y�֭p��Z�g��Ȇ��!�H0�E'��T��v��%��X���wq�g�kt�RM���A�l4�n�K���aHaw��Q���,"��`MLTtJ��f#ٚuNO���J��j��@�©�WvVOzu�����R]���v<�'zY��;�	�_�c3�$"����>�. /��9�~;��)�搂};��ٰ�߃�#���
;�l�E�cR�j����<Rl���9�g������>N�:i�Ი��*�Έ���3�}�,���$n��gz���8�흂fL�o�_w!G�"�k/�؜YՔeꍂ�C��(."*3М���%	�}�8�;�6�k��pu�X=M��d\zJ�r��E#*҇�E;I��[�*��+x��q�y�,��3�RIw��\�����})\�f%�L'�	e�!Y*�a/��RV���4����zb�+^�������y]l�ǿNM9�
�_A���.������� P��&�ڸ���NNR�~�??�=3|���"���B-$vq�{N~P��Ɨ7ؒ@v�Ԧ5�|��X�%�zL�1�����u�ڠ)a���q�%-t�3ri���|I�Eb�ԇ���b���'�<�<�⠁{�4X~t�Yf����(�P����]î�z�LHSB-��z��;��e+�ip�Q���:X������� ���r-����Liڳ |�߰�^&�h�L]�lt�{)Z��1��)u���s.ʐ��.����u�n�vDt�+z̪�+���8
B�͌�c�$	�'ӣZz��G�kB�M3r�vpQ��V����6d.����X}���۳�.I׽DƯ�w\��%~Zb�T���i�����*T�@ˢ�)�y���CFv��ͩ>�J9\�3l��$�h���e9M0yKhbn��i�����ђ�>"?q�Ǯ��2ܔ�?t}�Ԫ.��<\T��seЩ]F.�Z���*'���k ���k�춤��<��Oj@~�q�nY9	̐Z�e���蚐���"0���f��9$CvPĝ�7Q&r�m��efϫ➎h^Ӫ+|=7s4��s~��Ѝ�L�u��/��s��e��WM���>�m��������_�D��xH�SxA���Jt��4��q^��1���S�2AU��?��Z"��q�s�ݮ�� �^��n��/s���߇H�&���h�n�Ƽ�-i�9�Й�D��NZ8�&1)k�
�� [/ڬ�~I
�m�e��.�q�~Ҟ��^�r'l	*�d?YbS�D�%��	��5���0�3z..�P�О(#�A�#h�
AW+P��D��_܋\5+���.�c�YU la����o�Mu��B睩��m	佂�E&���a��IP�-��R��aD�"�R�+ҝf��,ͽ�v��O���~�qp	"�iBX���ǆ���-Hi�~��?�&��:��Y����H�ư-dw����g����7L��{`?Y4=NI�7d�V���?8kg��;��x�k	��wܥ����)}W�P3���^�	k�E �3�q@J@[+���J?G��󳣪�`?�Y�D�����OX�+[\�΁�\�Q�����YH��<�5��8�uH�L�M�F;���������v���jg�,�o[�[]���go�c�C�4?K
�ak��A�n�:��#-$���KePoƂ,���ƒ{�|�����\�$�u�3qt�	�����$��5Hz���懍/B*������q�f��Lyڟ6��_]�HR��w���c6hޑ�r{%��'�ށ�L+v�Y����Π#��ٶ+��� ��\[P-2НM|ok�����!<�Ɗvn��+.FW��1m�)�� `�������b��z��<�Sr�R�v+w`k*�y���,�����H{}��=��1�)��k��t'�QN�+J����3 "��'x��(������H#.H�)��4ou��7�,A�*r��8B!:>+�{YĒݠa�{��m��a}/T�9��F�'=�w�AQSэ�EMmN���c��So�Q0� ��]<ろ����Q���¦�Az;�8�V�����K+�:��R��Y��O8��b�d����a���	�D�Q��rh�%���;mF��p[�3�j���R�4꓏p�ϣ��}h�嵾���6a�ˆ�)��@�@�{8��v�Ity��#�(��AFpj���NM��rP!P�}������{Ӣ˸�N8����Ab�W�Q�0��I8�v! ��r�ɥO�RHz��Gu�N����}�DnyNY�e�*$ύ���@���W	�P<1Pp�п`�h��N�=f1�^���9�D�Z/���n�)�$tKJ���Koz~Q~ѬW�*Y�����w̰�c������2���8Gq�(陜]-���t,gy�*t#���$�ʗ�G����^��Ϊ�:0�LIǊ�K���D09N[]9�����IҐur�	q�9�(��g�Z�����܏c�|���F�)���(?5d�߳�$�\�默tA�>b�'-�9��u僚sY$A�s�L"���{�H/ O#dI{y��k�S��	�K�BN��_ts��hԈ(�V/�"��$�.�Y��h������D��L���]x��f`�Np�����8�ߧd��+|���J]
(����#l�|����r��ԩ˰��裄��I�i�K6-�P���Շ:n'x�{�	@W'0鱑��7Ȭ&�sJ�19�S���l����n�ֈ�)��X�z��9w�9��������/o�Q7��&E����ב��=�  z�D���ü!`��Z����1��Ɓ�Q�yӆ�G�[����N[l( ��ۥ�/���x�-;�e` 2Zj�f��g6�L���*��1X�L�/ю�����J��x��쿂j\�i'd�x��E��㮣kۖ���T�9��p�wOpV�B�l]�g�
9ȴ�%�����-6�7IF�K�aJFs	�"�ҳ"( ��QJ֑�ˁ�����d`à����`���ϴ̛��K��OVs$�+��!����F�: w��{\����?�j� ��� 	i%��u��z���{Z�S�h�ӛ�a��I� ^*���ض�!� N����碠)u&S|��>��9�wt�/IYw�6�_N���YUn�@�h�uN�X�䬊�3��S��`��c�tC-yG7����W�7&������-�q�KO�Ee��'�,'�H)�M0>��BC����I�[7Zki����*7è��Ù ��Y��<b�= ���	J3HF�	�S��	H#��/m�	�~��O-����XF>�FR���rq�����>CQ�iܝ�q&�磆b~���WV���Z�r�V�~t���ˬR���ul�b�z��������	��=|�V�Q�A�(������(�N�o�qz���G�Ǉ3�������g��Ϻ�GҠE���e�*ݲ��mv�x<g��ݳs����c�-��z��W����8���8��C�ՙ0��~�E�O�.K�XYcF�6�`�+����N���`��?l�v��O�oeW��ښ��Kn������Q�4�:7����.�ά*��1�4�ԡ�Z�o>,�ۀD߹#�䛟~��CվV��Y�v��NI��m����d.UZ�Dd!��	��Q��%��P�E���G�{~ɕ'�F$�H�����,�z��?�- *H����S��$x/���)��Hh�F0��bۙg'�WMet��k$�mx�ŵSʘ��ZJ,r�E`����͵k�����Je��|~��~�"<oG�]�g��f軩DDjn��̫s�h��S/>�(�E��6���;������F��THQ�$v�`<�T� [�����bՔ	{�3��GWz�����~J��n'Y,����$4��D��lw��d�Cc�'ď��K��'4'jOA%�&��DX�NT��R)�����E���$HV�pb�rֺP���*G�Г���7J��:�\�Շ�xȆ+���^	d|H	�ۭz����3���i�	��쥩��;rTA��#ןRP�7�xI÷�+J�]�jv%�?�с]|[�7�)����{%�P}�g#�M�"��_~���xY�%�g���7�#���F��#��1�����@�v��F�I�d0�>�^{\�g�1HBOi	%W.�?�{Bx�d����4����3y��^v{1[ ���@D�q�OBhi�r�h@W��A��D�软�LI���O�iB��D��UY�HX0z/�5s�ӹ���Iob* �GY,�,NO)���@I7�&L�yU& ��7��kD$�	��v�S�W��ý��;�6O�5�}�̇�R�*V�������+w��NpR�˪;Q߯ڏ�=2^�r�t��D��6��(��ē���x�̭OCd��{����2)S,@� �}��Fț�\Ya���3xKSq`\&���^c�Tz��Ab�v�_{,���0'��Ͽ<�c"�����D�nU�R|K��0K$�I<�:�##R$�|�{�NK���<�#�/�h��Z;����T"�.xfW�+�����$
3&]�����^o��aR�҇`Џ��'��Q���wL{���u;����@�_�s�$r�Q ���V�z��#����;�6<B0y�ϻ��C��%�?����9�2�9�}޼�,�ԣ��ih��_�|�mx;��'�0��r�a>��y���P�"2�A�$�����:Sx��Y�U���.2����BQU�P�@b��,�t�'��6K\+;m��J��ͣ���8���#�Йc�aT��1^7����%Ȗ�ME�@Ǜu��%J��k��K򳾽�D��g�P�c�ѿ��0ͅǥ� n�E�3��Ri����v�l���&ݺyu@A�V��@?6&�W���m��Y/�K�:��1�#a$�<wnvb��sG� "��j}���F��rvzK&7Lf�����i27Vp�={@�d`���-�x[.yj�ǻt��#�-�7	�%&e�U�#I�D�/ԫSMi�s��N���y�A32I~�A�wu#���l��W��#|�5u�F�KGqk?�M� �}��8����c�o�T���7x��&�������{3��O�+�"8�����d�@�'?G[�6�~B�u�nf���:�,�(D�+@u�$N�z�l�辅 /F�U�]w��\6��z*y*�W7�)�[/�P�-������� �5\�y\|��������?�Yr�$�&�Ȗ!l)�%Y\�,q�0u9d�����f􋼬�_��l�^�C`f�ޟ��;ؓ�c��ZyKK0�9�Gk���\��;n?����'<���ǭ	dX`
\c4��!J�`�u��mw�$���K!�nHDD�z��V���� ��'�"l1�D��h홱�Sר�����/W"�H7Gy�e\������-[ZNR�Z���AY���hh�Y�,:�S��SԻ�ј����l�8��%������2}����X> �0�蹬5���D�e-��_��1.�@�!�FT�R�!iO@ٝ����8��6	�[��y�Eb�b�P��	�l5���
�7���#-1-ً�7�U|}�2fȷ�,.��Es@��o{� ��w� n��52I��t��z����#.1?�m�'��O�$����E��|5^9�i(�9�g+U����-E���+
qD�?.������ �>\����=��@�N��G��iX��W���氛��j�;��qb�pR�#�,@ �9ޑ�6d���t񉭗w��V�6˹�;����8bx&���5�B:�[0^@�}��W��.��d�r&�����0DZ��A��kr�<3�>�@��1�=�"���C�Ư'TVL<C9D]�[���S!��b&�C�S���K��ʊ-Wu�&y����!��t�x��M���F�MW	�v�{Z�z��ܕ�8�0��ö��d){��1�c���kS(0�`f6 %P�8~��Qk���/ƜE����@��幋�1D����<@1��j*LF���~��=���l�w&�q�k��u��`�7d`�.��7����=@ Q��ONL�\"-�L���);-i���������O�"6ؔ�1i��=��엨*rEj4Ic�#���bR�%t��S���G��f���k�l�n6��g����"��E��,ikO�b��@6���(��X_�s�UX��e�1t#:�kʵ�f�N��ڇM�V$�)*���ݎW�ՂGp+��("������)�B-Q�&|���N�[N�P�Z1��`�;5n����%��U/e�F�u�V�Y�R�pmĉ0R��K�#�t�I�{i��7��#�J##����'2\�T}f�m������,y�tx������ʖB�`T�����ڽy��׈���ez�(N�YK��}�Eԛ4A�x	���+U����09 � ���~y��^���L���r����T6{�.��\[B��s�Je:�<��6��Vr|�)1��@�(���5�Uo����05BΤ!�������A'��?����i8�2����%�!+�R�%B.���6dˬ(o���
#?�1C�Q��~Kr<�y�Y��F�i��m�����L�U"���骠��٫����xq��*9[ǔ)���kJ���+��Y6�,nV�f���l��K�)�3w;ubQ5�_�&�JS-�/v�fdM_;ƿ�)�yj�i3j6���.����a:� ������?T�~\ߦ:���c\�eFs宷R�!Dś7I)�v7�2KIRt�����	��RB���|��e�%���ܓ�̻�@YL��i�N��\xPBq�)-�4��r7#��z�W��=~H0���,�[�l�.�jB�W>j�{���ζ���Z�n L�ؗ�*�]�~�ɻ@V�e>�����_Ј�|�4���
P�ϥ����x��޵n'$�T�Y�8�;�]� :\�ͯ� � =�Aʧ�Q��~Y������}�e�9���P�B�
�Io�\��ؒ����h�R��B%)��&� �iu�Y��P����&&���)��CZ���A~�r�����I���Յ�؈�>�UJ��q�8{G��9qn���@�Ł����;nb:����2ݾjٸ1��O�GJ��e���Vc#{e:ЦQX
��hv���)d��ɶ�$`����؋R)�����·��J�{s�T�!��lư���{�(���4k�[jް|�{�Qz��N������X6�& O���O���]�np����ꆺq���$����g*tB�u� �no��soI���Kg'�ъ����`�@<
}z��Tc'��̥NH���W-������VG����GyJ�z����i�%),7��^T���Wd�P�d�[8l@���h1��a�wS�?����*�QB��E��7��9�����gJ�B��$H���F�1]=
���h�,�-�ˣ�#��~V�-[��^z� ����T`N*u]�"&�S�05�\�@�B�논s�/��C[���ߙ(3N�E�q��{(�V�7�����r�x�:B_JX�uO����S�e�㘌8�#�K?7E2;���U��|s�8��{�,85Dm�Q����^;���-��)c�oCC�O�H�*���t�fDUvq�:�Ol�򗰥���f<ė1n��FNO��ɖ�*��7۩$��P�T��z:&�Y�;F�ӌ�Z�o|����+31����9Dt}�ӣ��0v-V�R	v61��j7%�����r�҇��4�E*�Bpl�ė�5t����h� ����D���4dp2�Y� �a���,��_r��f��DP� i���w����]'i6;t�����Ĩ��3�hs�n	%|_�[�f����G��q�]A���h���q7i�p�6<��K�]t���������k_`�;{�$���Y��ܤ�?��Ή�orq�Lgx����%�[�xVQ҃zZǜ �@��Ɏk3{k� �s�H���(�u~�H��Bs,�wBC	!��˭�gA���~�r��Ücl�⤾����h���3<��M�~�P��Տ��'��#��;�;�N�
 ���]7��k�
E��|��~���k;Ti�������zdVUC!�ct�����	��o�[��p�,���ƀ��TjH��1�x��Q����_	_����.�~͂m���sc7~����e�D-C'���%���GyliHO۹Ev��\����W�d���ȝ�K���R���K�\P��-���ݒFJ��T����O�ܱ�;��ʇ��.�'i���]�KY,Ǒ�)����G�r�����yX�ʐK
�u��z��uc_$�6L��2V��l�����-<r�;�4Ӹ�N�M8Kv�ހ(
#M��4n�NT׉ب��Z)���U�tu=���؏K�>�G9}N�{`'���/7A���Mq5lc��N�	|���~�\���'��å�"^!r&(@5Y��0Y�����ep�U@��۲�ߓ�1Q�n������]��Sn�޶�P칇��$�`��@Bo�,`�:��h.^r_�o"N�ipѐ�R���6ͫ�J��G�9��|k[i8�icT�Ɍ��(����D��|>��7��&X��q��<�+ŀ0�A��#�D�7��b��W����1�È�a�k�#��z�Ȓ��ʔ*9 =ʳO8�)O@(o�/�#�$��Tru�!)
�W����k�Jo�'}��x'MH �M��oY�*�FB����܍�k�S`��>��|Ui~0����Y����J�2PeޞQQ���8�=�ӖR����s�t��P�n+$��tR�6��KSb1l�l�o��b�A��Z�]�U��1��I� z�X,4��o�� ��;��S�i�A����vG'��u�4���[������q����ua߷q�~NO�"�\sTb�_�vM�����-��Q���h-�`K��A�G��ٺ+aEngw�J�l�&@D�I�8�ַ/�3�u
'u;�b���I�!�TiS���͚ӗ��.xe�L�/�E�8�7b�zH���G�5�c=&���۝O�$�"�� �ͭs��{(I�v�*��{�ѯ=|� $�q��F�C(;N7�&C�����׷�%�tUDHHg��qU �Ue7�:Gϩ��'���{�1�v��lY�W�p���[�.�X�����H&oZ���^�"�l~{U �?P��7��}a�#�V!�GEm�FD|tU��t[�VE������	�Om48AV� i��է|Ě���k���XR 7���x,��&���`R��/gv�q5P�Uٹo���*}R�����ج|0�4% ,^�`Z��� _�)�|ýR��P��8]++�[=	��ʲ7ŀ���h�)IF��� CEߠY���<OP��;y7����]BU)0Fi{	����@���N�>�i��Ĳ�h��^���d`q�8^�&���A�OmŦ�
�������+c�͊�R��r�X.ץ����qD|�~U�L�}fE����u���`�P(���U6YV�ZQPJ�@��:�j�������bkz.�7&:��#�T�.{8�{�>m��[
9�#F���;�G��"oM._���c0��:���%��Ѻ��O�8�,�57xTp4���O|ˍ���Oe3
�����T�vXK'tzFm�.�[E�jB��,��%���O�"p_���5�ȿQ��8j�s�����07�{HT#��V-f�Є7J�\�Ny����L �u[���5�y�'8��쪞
=&ϫ��]���S��Π�%w
��Ƞ��xQ8Q���Ј_6����J}��c |?����������eoDU���J#�Q&K=F�����cڕ�~5�P]����o�/e�ɹ!4�vw���x�4�c�S��5Z�`� �����.�.D�.&�1��s�(uB�����7�9��n�9`���}�4��N?x��~p�(.�{Y.���|����]X�<������
�ϓ}���G`A>��m�#B$1o;�NV���>m�>�%����	+�����j��c���K���gUz$�Q/<�a6�s��呗r��H �sp�z�6�vch6�<B���<@�i��~ݱ����q���c2QB�^�7�\NO,Q�&�'i~�aq�c7$����� ��t@�o��J�����h[�$�Y�#���l>��-̹�ӑt]v���X���S^gxB&��+8"�僐��������DJ�ON��R����R#nP�.+��0�N���^)tF��e*��M�i?��w�␏^�8�ѕM��+�-�vjdI{�;�+�}a��"�Z��/7є[�[1��W���ɚ��.���4):�|vˍ�T����@��^�|���6�9�����xy܎
��QF�RD_7���!����䑮���B]��6���Hʲ��
�A�9��.����d�	xi&�tJ����6w)%��$���1��{F��e��]i:�r�LE�S���%��'7���*k�)B���Xm�g�/t�c/�ņ�v��)���5!^pi�X-�X�MҨR���4�P�sݘ<j���� . B�s�����*�T��&&_wտ�=�$��Ī�wvs߁M�1m���hQ�M h�jNz���b!'qHׇO��!�%-���XC�>�("`����p�ܑ��ٞ���u;�x���m7��W���{�v:���=M-fR����T�.��@�8$�σg�H���\A:��@@���\��5Nq>�\� [�>��6�G%G��
���������nH��}b-(K����a�e��;�u$�����g	[2UAke�٩�W@�uMi�F7��C�I>���~w:����'�nz5|oe)YT,N��w. `��bF�ef`�@��C�k*��
?s_�;�cҾWY�����/�~�ܑ����R0�hS$���Ēb \>����Pk�n�e��ө�H�0Y�3�rDr����5���3oGD�ִ��$�*L^�^$�"�ψ��P�u�V���Q��[�_a����'5��d\'�7΋Tn₷r�����>�T�3�z�F��$�[�$$�PF1T�.C�0;���H�LYA��ʫ�D_�o]~�Y��L��!�`o�3h�,4�ʳ�.�B�*����7��g���dh��)Ji�`��ձ�|:X��J���jTĘ��� ��z	x'�l^�c�'h���
���j#!�K��μ$z��}~��'u%�E�L.����Ve��`A$>	'�g7V��yQ�`��.�"���EP�}�G���܉(���?{IKP���(6��;i��HB}��@%z��}O)n,� ф�+��VQvIh�T�K����}�UN�Cf6�U����Y����[����4����uΛe>�J��$C��xj,�nB�R,v�`������u��wHt�bZí�z;/��I���b*S���K5��O����a$�#	��^�rIa�C�N�}h��^M!�}uX�P�!5�V�593^���<�������Ŋ˯�ǲ��ʗ��/D��?�g�������	K|_�� 1K�82�����e*� s�+�2��CUl2/���1�Ǹ�4���������%��(�s�X�:���x�'�#�m_��_Gv'�����MrG*uU*����d�t[^���r�E��g@SMa�!֟��c���<�ߔ��*+�G1��),�}`^��!��ʎ��?
-O�1zZ!�3�Ȗ
����``J�����,�9+�s]_�7�����C
�~�5�3�r�J(xp�o�T�Z���rF�F��/ڢ��'�N4=�~�0.�뇷J�]DU	]�v����#�j�i���RP\���w�F���_+Ǆ���ꖞl����e
�)�0Q����e��	�j�"�!l(U�ř����)¸�Q#.�'�z�c���6����ǱF�����]_\���������AG).���C��(��1?Hzـ����i˗b�\6$2z�Q�s������>