use work.CoarseAlignment_pack.all;

architecture Rtl of CoarseAlignment is

begin


end architecture;