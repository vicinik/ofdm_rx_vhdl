��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X�D�(lQ9e-.?������������!F���O�ZU"�������Bu>�sa��Ҁ� ��uɸ���p}0�~]��è>Aܝ��i��|D"����1<l4�3	V�-(#���%��;=��p��;�BJ���W�8^/Z�0�8�#��9���QSK^oh0�x�$���\�1�E�J��H+Ds5n��:�bW:����:FNd^B����{df/O�����zcs���e�v�Nݮ`��\2xf�A�{��H�~ZѮ�ُ�,q���4'h����:�f�J�I���iC�]��P��`�4YG���̊�aYw�2����x�k��0���m���=|:��3���2|�y@�U��Q��/����eoԌ����v��3�����#��<Qa����A����'��\�(�Վ�5�P�� ���~үcQ-�op�������=��g��w�̽��t�#�p���T���+��(�_���R��.{%Z\PH���*���v�!��11��.@�@�'�{�Ķb�\�����D����]
�$�F�����!�A�Z>�4A�L.	�c��R�4�/9�:��ou������jc�t������v� c��	�5�FR���]\g���6�A���%�K;�?qS>v��A�x������IF��9�'a�F%�a�2Q�	���Ama��� e6���E��x�Q��>��z|n����חp�w�<P����v�h5h���h�g#8�sb�cߪ�8���}>��PnM/��³8S��h�ftѼ�B
�"�$�����?��8�k��*E�'���_�>j���\�)�)a��"�6ɖe�~�����`h�D��f�K�C`o��f��9�H�V�w���c��*����+-���痭CNlSK�_�#�W�� �'�n���O���1���H �s��+5{=]�jg��k��2��y2��wq,�V鳎ψ��x��m��H��w�{MH�
O�մ1����z�<�����:�[����^yK^� Z�����[(�ؖ� UI����֣���<D��7�~!=���L,�R�Ox�n�'�,�r�n$8��|�v~j+�:�^�:M�E�D�z�|�l,^Of�V)'���sXc%��迓���+|�:n�mR��y;���%9��`8��ͥ!�W|!�A�ŐR�7�W�@'��i�;ǻ �=&�F������
����b����hp��#���k<ʯ����9mB�{�������>hY�`��0���T6�� ��J�qˊ]&��;�AK�D��'D1K�",c�P�b�s�}�Z3��8�i�Q>�0�K��iф���B]�5p�|ns���<��3���i�")�{ n�����R�=�#5qFTd���Y�����6��E�Ky���tq1��Y5~�Mn���{�G�ɠn��eb���2����j���}��샩�W�"��B��!���Hn9k�L�D�����/�s�7̽�q	����o��U��q~1��p]|��ЙG/�"�(nK�B�伒��di,H?�u���aJ�n���.~J�o\���	�"P��жĈ_߲��{S�w��0�$}�VWVZ�����^�&��'��^s~四M硂Ɓw�g��ƷG�OH9������	�{B�|�j�.R�~��2��P-3ޅYc���कֻ��p�����/������#�iG�b��a�ˀw�齝�Wp����{C�D���k �Om�Vc1C<�l��s���'�`�VG�����<����K����CTHN�?��[bo��łߙb��Il=�,A��$I��[\`'�#�(�5-��ƅ0&�(P�^F�;FRZ�n/,);�`�'&P������h�����_~�Z��S��`S��U/B�qt~G�ݮ�UYۭ�/|&T~��-Ѝ��}�a�JY�\��hr���V���L�I��US�l�,f	áo�W�BCP �{���ۯVщu�2��U�;�>;���	�� ��je~��{.E1�����W]6�3�մ_J�g��L�A����$V�[ 4�y�2�,�| Aj$���o6-�z����a��-��ՅJM%�H.�A��c�p� Ʊ'&���s��j@��[^�vAuϣ�(*S���܉�t�U6��{5�a�	�;;jBрO��F�J���<F\e;���Ξ��-X��P�^�K1EB�p����A�Wh�UŰ	TґYE,35�t�O�5�0)d�{��$����ᮺ���� 0q��N��/Q;s9zo/�/�{ו�<��ꪶ+sQyR�6Tb���Ͱ���pP]l��Uڵ�vW��-	��'&��?�6?����H���:���ҵ�Z.{��U���% Nw_L�-�1Ӆ��.z��P5Dխtv����	3���<��E9��8(Vn
LU��	�@؈N�._>����q��!�P��Ŵ4�E<\Ƶ�zP���F�$Ne�2�y�Oў=.���B��Ƭ:�.��J����R6&`E
����UMm����j��O��]�腁�	k�g�Q��B�T.��f����Jw��v�5��P`�7RK����V"Q�1�v4���Kz
K?Ru�4���O�<6��*�v-�a�K= ɋ�x/ �Í��n�_���6�g�qXKX�ʖ�1]?_	5�bBd%�Z�l����4g�����#6.�=��:�G��ՀD���:[.7T��a�R`�e���9��X叼�{P�&'�t��B^��r�)�FPe�Qwr�~xި���G0d��k�� �4rp@Eo�*a����{�0/|;�O�ap��b���_ɪ7D1ޒ/��k�xh�H|���!~����?��3]��t�9C/^�v��1��}��27�J��t��W�'�E�-q�g�t��4���Ke]ۼZT�iϕ���ւ%����n�H3�\��Lڡs�#U��6��B>^���m��l��W� ���܇N"��%��րB�F��Ν�r�/�0D���h<㠪B�ӄlE�g\/������H�2/HG�s��w|.��96��(!�"0��T���ɩ�6/����-��3����7�\��+~:�+���!��=I�$�T�/.�?Ѓ:HW�ӽ�����9���A�@[�'���#� ����BC��4wn\4�y�����!�zٜ�Ɇ� ��P����wdn&9���=`�x�Ȩ�����[�N}���JؠH����6� X}���d"F����XE�j�P��%�\W�ׁc��.�&E_w���TУ�:
�ݩ?,�CD:�$���k"��MV�^�q�[z�ъ'eֳ��oqı��IQC�����w 
��>�@�wX�(��r4�z�Z�ę�:
��|�J¾AXH��'������c�����t�!�/��6��U�]>,G�1�f�2�C���	��1輻�s���A6a��.{�w��>v�/�a����? ;9�/r�2�/z�I`���^o8�����|�~���aO=}�RZ�=�E�vM-6�l�֊��>-"A$Kl������g�(� �S?��m���.�k�G(s|m/�ƨ+�K�W=w=f�<O>�="Жk���'4�-i���@�|l�ƍU{�D�B+���qTΕf�t�G��ؼ�#C�zafrh�8~���:�?�@���W���z��?��F��eV�P��~���( ��c�|9�؊.�^$�>��k�S�O���@��������ڦX�����E`��[1��,g� �	i�$�$ĴH-���D缿ț$�A�M<p�ғ�S ,W���T��ޛ
2��M!�����s0W��fΈ�;��9��溨�c�R)!�5�O��V^ޭ�-��]+Sz��E�T�/�����d�	��O�d�t�!��lL�3Oe�jn��Q&ϛ30��۩[)�z1���BvW�>gx\��K�}��<��Ų]+�@���_�(΄��Y��q�;нi���� �9E؄��--O�Oz+�W�F�;b�tIԯ$Df[O�i�'
*:Ŗ��-�(�8�eJl}s9���j�K�=�����1I�b���U����}�t�Ek;�̖�4{���ˌ���j�_��]I��i��%<�C�k�q������e�-3�%E�� *KB��=m�h�8�aW�H|�:ãD�<V�W��O��E����fV�	�>����.���B�v�dWBB9��WoLN��A�|n&��@s"Yg��J���#*����b������Á&�(�7��M��3:Dd�$EB�� 7}R�s�inj�x���ݗD	[�Y��K���t�Mќ|ǉ��3Ȗ�˨�t�gC�e�=1�&�����ֻ������Q��r�u�$ܫ �4b���3�'���-a�����_�5���"�(�&N�HM�xL�2#�O��R)�a="g�6�R�޿��ל1fCm�V-�n�Ԭ��<5*�.�9
����%/'�����А���?��>m[i����쌪V�������҅���պ�������$�ȴ��Xo�d�^�	�]W:�bC�n��H�����nw����\��,XM� �]�Ҧ�?<�l��N�	�;��ZK��܋�w���*,����(*��(�s D�؋�O��S�����U�����Z%j�>�<'������ىDޯ�~��FNr3J8��-rЫ5(O��S���N����{Ԩ�j��Ei�+��t�
p�s���at��*���_M��Is�<������\I�]��A��G��$H�@	�IC�������	3g�6�U��f���"j;,,6J���,�'#*C]ʜP���������Q�M���AOK���Y��Fe@w���=-kf+���]�I�+LN���y4K#�1_�	������1k���-�M�Q�]RƦ�D�Z�>j���ǅ�t<Wq��x�b����֞�c�oDL��4� ,j����cR�:�h�M�Jf��J�~�`��+l7��Ѿ/�{�L�����=Qu.ޮH���Rą�r?�b,}�m�w��a�	���ı!m	�֬_�w/�0��xa�b:Y Pr�NV�s/���r��R@�SLD�6�R_}-�{�)2j|��@:>|�I����ńIm8<ӱ(��
l�F1D���PÃ��t@ɼ	^��a��!�S(���J�m����oa���](X��lI�Ҝ!	�V�q��
V�������pƺ�w9I�dM�%w�����Ha�'�?�رI���lc>��F�y��g�ћ3��F�<�m��Fت绻TE�C��p샆�"X��0�e2��w*��ė� ׽��(�T$����Cf�����8�QFG�{0��!Ӳy�����[�h�����_{�!�$��-��o\Dgg��E�L��P2U-0��}��&m����� �7BV$����aͪY���B+#� ��JGu�������ۇͼ�I��;?)�Mp9�@`7����Dˊ܁��,�1�2�O�o����%z�g��H>KӖn���?�`��6����q3X�<_�� �p�(�x�:�������1��i`�`�"E屟�������g���b��"|�]�' ێ3W ������S�@Nm.F+/�"$|�g���E���|�-Bhd���h0��uvؤJ�S�A��Nʦ	��U���@�ݢ�X��+���l�n�ʢ��s��4&r6V~#&}�̙t�t���/��W�'[.��
qƖ�*K�"uS����Ω9Ƶ�Y�<8�"�W�14L0��*[ԚF�-tnh};6���RN[�>9�5���Z��I����A9	�\�4�^$��\��vӶ� F�Eӊ�� q��K�-�	$ǣ��f>�|e�]��6X����!�^���U�42���y�LYD���������8�Oܴ%$ZAk��u����+/��$��<�6��
.����^����؃m�NF�Ó�"��?(q�O���aF<V��?�p�U� ������q"��Y�����+�\�Wr١n\J������\�	�~�'�J��s��^�������!b&S����Sb*چm,Nv՘U�T��ݾj"��dƒPL܅��h��;�4^�[r�NC��K���Kv͎��q]���~��6��+��7�v2�.��w������]п����Fw6�m#���u*Q�{ ���k�3�5H���+��S�; E
\�S~��6O�g ���q[�2СE����Q'�Z	\�*���UV��YϦ/d�g�j�~��ĩ3WFSd��sڌ`����l7���m�&��4��˲���k
V {�X�rZ�|��ޜ�UhG�XW!+�υ7��B���f{=9W�(P�N@[& ����юOJ2���q�����Gu�	<�x[���C�3Ru��?��#�ϙCWU30��I�L s�B���'Q�L�9@��gH�XB��an�3E�7�����RP�"38n6*�/��ʤD�oy��quѽ�ز������\�ǡ95K��3xQ�� D��8�HG�x����1#�()A�|���t�ekS��|�\�b�{�Y5?P{^�bbd�ْj��?P�SZ��H��A� �!�	��)D�������bg���%��
��er��Z��Ml:���oi��
�j���^�\j�-��)�k�a=�.1����]��r2xa��N�}`#O��m	bP����X=�@E�	 �P*�%�f��hᯓ�N7�O9��XLi�:�	R�Ʋ�4z:�[�Uy�{�؟��I��#V5���^`���;$�:L=/�g(��=�y+��wa���a����i���{N��(�g2�A �l�8�o����ρ�=y�:�(>_"=��QVa��C�}����
,�IEQ�k㺼C=�����1�>̏�#���+��DJ�����f{����c�2*�Z�W�.L�»Ꙭ��o��� �S=�����YF�߼k�P�@*P�G���+%�\On1��B[ W�21\c����<���d;λߧp;�Ǽ_���|��{���0.��39�*EGg]_��M(P#�����V��^h
�/��N9'ѷ,QL뀉��en��L���W*���ª��z5���̒��0�����H1���7��9���B4�r�Z�[}�� d��t�%TR���І)8�f�Tz�UVn��s�R��9���偲�,�8�]�e�)<�3[<%�S�w�92�A�~踸�K��|��zV(��"�yF�
��w�j�~�g3{��*P��:ABDh�P��C�X1�h���U/GJ���JD�������u7M\�q}{�[#���I�&��hf�=g��(�J��]�=��jA=6�s��
nS4{z�9rq��_��T�D�o%���lU,�VY�{nyđ��f9���y$_����n0W�.�X�{	9	�tz��5�j�_(��4w�4�n��_�����E�7�`������g*MJΐ��f��L)C�y��C:��ä�?�d�i+:%H�q��w�y�5B��UVM�
���z��A��װ-6	O�I���Eٶ�O?2?���=9�nw-������{�kJ�I������r�&ə�B��fr!���
�����H+d7E�{�۸���m�Fy�ݵ%5��2��2�\\Ӷ|i���u������J@v}�[�P)�#_�u:��mD*!��5˟���P�D���BF	z6����~cDc�:Q���m���ZNa�+���W����'?��x��Z:,l������~��?�g�;�R"�jB���������D4v��#:�">�RF������Rz�<2�?����l�9��A�ָ�$Iz�l�q|{ֵ�M�*]nt�^Y�P>9k���%�a`U��3�ɘ5�x�~l.��{�xG���T<��-Bz~�>� ��Z���\ ��~Ν0��;[�w�o��mPj���[�=��qi��^�'3E�C���&ڇ��4ۄ��2�,���[`������i�i"8Y��P��0U�W=t�Y[`�@_7� �G��N�]���]T�J��3%x&��m���W�z���ɢ���,��	�;OX�ωd?=��L�br�j��J�������,��T�Z�"��ѝ�O��z{��AݻzE֗��0\���a�����t7iU�b�J[d{ު�F��GZ��E[��I�5�[zzQ��� u�y3�*@aa�:M�7�g���RI��:}�0�>�{�JU�
Drq����w'4��%ηr�Y'��F�MW=x�"��H!k����Q(]��1���F�����[EeV1�zK�X-\�o��]�d�E���T�vf��ϸ�X�g_� Z�iu�r�Q��HN�}���`]ǹ�9���(<�����)��5�=X�W�6VS��Dլ�*�b-���tr���eB������l~-��t�8��6�F�xlNw��JO
l�k�0�!+�؍�p�76�Z��0���B9Gϊ��Z�������������d�Fn�R
w���w>����A���c���G!��}ԑ>��ŋ�SOU�$4��s*��|���o.��[&5x��j���mT�h(��W�0�I�kK\��G�}�?j��Y���]+U�3Y�����ʬuY�+��!�9�X���:�t��͕h���z�X?'��4/�
���*�)�9!�ڮ� �mE�����}�KC<zE�;�9۪�)�B�8(�r�H�4�O%���2�	(D���Gq� Op���i���:m�2D���?������YXj;����մ�Pw�����/zu1烉D���n���
^�KOW;��^J-Ŭ��5CK�6���bO��y��D%��>O�#��%�(� �����~��L򮙂,
�-���y�o�GH�r�F9b��ɽNVqŰՍ�YN���H�(Ju(<j�s��Y�N�˞n��{���xk��SN��/�2��e����u��,�Z���a��P�n�-n�m��{���7���X5�����E�[,d�xW��%��w�	?x5���On�-�i�nC��Ľ��,A�5�2[1���aTh�5�Ѹ���1y��^V��Z.m��8��i{=���$X���t�]���p%�*�|���S�N$�(@X�e�~��1];`o�z���*йC?j�s��./Wn���p����6����)}�R~�[ԑ��.X�������q����$����3��K�O:���c���
�gR�k�����V���
�dV�S��aSQ%/t틢�
�/�uLb:�:�#R��kQ.�Hu�����h��ȉ2i��<�c�ճ�±l[����V{C]̈�H�:N�}�	��چN�]a��5���Ⳏgx�=���f��2җM�]
�x?e_��c��zBH�V��&���`�%��/
��,R����c��P��<���ս~�R,��2�H&Ub�<�e��J�&�)>��)��$���~���猕{�K
��K6PBF�6�C\�Zpϣ��}�}��{*�BiXC\K�1*V��X�yʨ����P�5Ѫ|��䝏�`w>KȪ����p^��q �,d�%��gU��m�{cK_�#y"�GG�!��;�Hsk��ќ�P*�"�����RÄ�1	:Ј� +Rjd�d��z�1`{/�J����T$1�Fϓ �M�(VJ|�/���q@�zW6�B�VƓ���W(��Y�W}@:9p�R�,���L��9��- '�	��&sF�C�c\g�a�� ښ��!3�n�&�\ڇɌ+9g�ḥ�4����u6����y���sEp=��_8�UcS�ض2�w�[��d����Vw�Q�,6��]�Sr��S?lLn�l�I�:��v�Nd�`yS_|VU-���*�]�h���:�X�`�l��o��1�����L�.bdF���N�܅��y _��P���X��źj�*���K� ��LZfM�K<XvX���G<w�kos��
V�(�s]HM.Q���d7j8��D��')1 oQ�i�ld@��Z~$d\��R���Zk~ǿ�<'Ze���Wm`s���,j��I�+Bb��y�O��l�����S�\�{�,�8�͠�\6�/�F�;d��9��T��`8��k`��q�����1vھ�R�*�p�1?�-'������xkV���T ^a����7�X����/G=��rtD	}��}���Ђ[3�V+C����,�ؓ�DҶ��?��CǷìS�^qk�����.T�OE���ɏ���e�p��la:�C���s�ol��B�82�����!���u�h9�%�ެ\x�%���B�@�<(,���]W�[��D����6��ͧ��W���mA}e�LtU����Z79`���Vi���9�F��im��SV������_r�=�	��-h�U3���|,l�g{1u�󷁦��@dݐ��<����3Z�2�A{t�A�L	�����ݛ��j��`�b�n:�6�
��:z��$3�`��H�Hَ��޻�����v3]�z���o�c�Nܔ!�Z��8���d�;-�1|j|%��I�-��%s�*�$U���y�\�2��M0���T��*�N����LA�Ν��8�z�t��@�c�L��7������~�-znsS#9&iv�m��:	��8�}�ő�"�OL�#��z�[b���>�w'�+���HO���
,r�}��*���R�'���s�zj䱹P1�� ���:4^���D�k��y����~��Sܭ.���"�%���m��R�-��֏ ��֛J������ѪĞ��U����wY�m���R����a��ƅ��Y�LY��4u?8� ����~���T�� -:Y,���r[m�Z5���+���������ڝɊ ��D��!)�BZ#	A�0��#�g�a�"oL�:�da�J?�W�hw�ԝ^(я#-���W%6X�y���ܓ��0oyo�H�lu'Ǫ<�������1X�9��,���RJ��XXԝu�#��v���'�������~޹��
DRrH�v��L�7�%��������D߉^)���k�dd���g�/�X�7G�ԯ�$�u����~/�\ ��<�C#)��ے���%�A�:�J�ĺ�r����/(����/���`aI�$��a���&�n�5d�4��̔�<P�Qn�ײ��5��)�DH���� ������Q�4�]@�e:�ow#CRx3��~�&j�.�:�o���2��44Y]�T��v�?�{N�v������66�Tu2�7�7�.O��r�J�D�O����"։���b�0?`� UR.�m�#�E����rcp} >l��A�HA�$Bc>6�"/O<�����b��б15Щ�#`Tg���r�+?��w�Gz�ϝa�Gq�1~VsS.0��v�`�}9�ʼ�O�&a+��!��
�4����{sVA���b�L����V���H5�7G.O�8J3C[��)$�p�ĪJ��^|��A�p�J�(�e#��t�J�Xk���v�������Mf�hl_3zM���
HP氽�Lj��mDS�\�#dqvx�ӌ=�1�2����jLԕ�$CK�P�&���\�U����R��U���݁�|��ze?	
/-�%T;<�0�pC�X�n�����s��3������D�`>'�r��ZUQM�oD��uơ����3�/;{/� ��&��6�?�Nîc�~r��:���E�Gl�9 P=��I�!Z�X�%�l�ao	���m����&�A�?�ү6)�����`���zy�w�������n�
XA�a��M�,
��`�3�;�Y�$�]n;�I]���V[�`���
2��t ieLV�]���a��n�G�zp��&��2� �nY�V�uvw��g���'@���N{��
0QU7��i�k����m��������"|.{p�
a�B��~������Jw\Q�1+{QH�ҩ��l�h�Zbr�v2��z�׬�O�m_�&��v��T�_�,e�!A���e��b_��N\��_D�n���x�������8����	�C5�A�!�  �g��v�&r�v��ݔ��)��tV$���=A�eH�9k�4��/+,�2����ޗ�z�����^Ei�� f	|�q�X�:�I�tLpe��>����m;ćK+������K���aN6�`)���6#�sS7���Hk��"62^���"6�#�[;-��B�@v;�����\h7P��Kf(���5��A���^�y�J�%�� ���@�!u�yh/}�bl����-���L�h���]O;L��I���Q-	YSֽ��%Jg-%i��Ǎq'���ʫ�E��?��4��(��}�(V���^>$ҫ���(��f�b�e���'��՜2wR�ȫ���� I*˥��"(�\��U���
�M�I���Hhq"�����c�_��Z�y'o| �D7\��03���!�"���qZ���ݸh�q���1 ��B�N�6��He���o;��B����[��t��(e���8y��(���g�ܮ�ظ��z�'A=�Ϥ��~��N'�KW��'���?�y���bT���N�6lI�#�%6ѿ�^����բ��#}��%����;�4����,��S0��G*ӵ�%(��+���p�	ࠧ��6{��#�Tt��*3Ӎ2e���9ǳv�5����^]��M�c���2�Wy�U=i;W�H�Q9m�x��d4	�U_��Jr80�,hȟ�.��e`'>i��#�����l}^q�3`�^�W|J�ux�B��6]w�%��<P?�*�6�{O%�����*�x',�Q�H���`Rg*�h�kT�`-$�ܾϝx�l@視V�>
=����||X~5�[$��Ղ��ѡ}�s�u�,����((
�Ё�f�-�n5��1��2C�N���|�ƒ�]xw�� ׭pn�g��u����;իMF{x@!
ⷸv�J<�P_k��G~(m7�,(����/���rԁ���'�L�hϏ���O���&1�2gfK	��
N��e%�W����V[���#��	�[�:ەjd\^
dY?�fYJ��	�I�R��������8H'd�
�0����ɽh*�]�֙�bR�=��~X�2��erF���'�S��7��m*f�+h?g�*uwz܅m�G�ܣ����ʧ��ő�*4�ww���w3 �(K%�N�Q��P���m����O�%X;��������ZJUn��#�`S3�/\�e�ꄮ^9S��&�HѺ����O�%��ȦJvL��F3Y�/tzO��9@��U���f��^��6rOu镲l�qH��PJ�D�Dv(�92L ��^�q���6�:dt�l�	t�_|՚��7���T6�4$�Xp�y���3�]�zM��d�喫�Hkv�"��%[��o��1�$�]���k�>f�sz����9<���8�M�W���C2�)[����;OCr�]���d/�Ⱦ��h����Eڜ���݀i�+jS9c(��qĠ��>�O�.��<�[��)@R����X�������� ��C�*=*���u|u���6�"���WY��� 5�-E��h%�ͼ��@��@`�뮌?�_���|����{N0{��f^�#��aYZd��uAJ��#�q����oF|i�,6�l�Ԑ���w��`!Wp&X�H����M��,t\1ͧ��p�RȞ�Z�<� ۓ��x5����V�.)Imcz���t~y�2�Q}��?%.9~;v�r�"�/��`NrV�~ݝ��ݪ��5Ź��_uB_��yi>�F=�U�p49�(}� A�D.�s�Ɔ�T�r �h᷻���B���F?���d	Z�}�����S9��M�u3�HU�Y��7ϳS-l��2��S�Y:q>��h���ݥ�tuC,|��R�r�8���Vtf���kF�� k,��Vބڛ�Z��3���M�� ��
�ч�V��Z�Pz.򔜰�ϣ�q�g�Ώ��6�Eg�i��;�$�^G�v%x_���eK��UO���g5�vYVS4�Q<�Ml�2Yk��(uؚ�w��3Ң�;R�g=�� /S�XS=�]��j ��315lۏ/���ė��~g�1��cӛ�Euٶ�k�e�qR,����1�A%�C7W�;8�IT��v����_ͻ|�P�0���r�	6� ih�t;�v0\*3�Q_��!s�}Q�C�YoВ,Oध��T�G+��2��?�t�$y,�5$+S}��8j��N���VЕ_�t6d��Z���	^�޻ڹ�g�k�~@2��DF�	1��`�i�>{���Uڢ��I�g�s[�Z!��T����8[y��\�Y�YH�6>��=6�s���������m\�,8��w.q��ޘx�/�:�{�%����"[:W���bh��!��_��C���9>�?��1ܱ�=eX�%
A9��Ӵ�
��>��d=n��-�~`�E��헍�wG�i���I.�)��/C� 3�����!��bx ��S�Ay=��KXqH����`2*� �E����Fn��6�:+\����DQd��V��)��M���nQF�f����lژY���9��d��#2S��2^�(��to�~�7�Mbj%��i�N�I��lx������E$μR�4��$F�-rZ�R��"%�.��
�^N�4z�)߱���@�_�[`�LGB&,%�A38�%������믵����uv��Cp۬W�"EuZ-��+�b	�}������`��hG�٪�|��Ǘl2t�����S�uL�˟��^4Kmr|�F�b�vk)�H���9�������Vk5�:I��@�6o=��������L�y�?�h�y�<��5-�b�j�X-���]ꖟ�>
2*ع���A �=�"�nL8�9{F"��;���ulH�� 00uH�g�Do8��p��c�8�H��ށ[�"l��3�_��[B��_d�~d�|It"8n�nr��,�l{Po� �`�ծ$�ԩ����lf��H;���u��]���$�է��3}��n�c�g(լ��@�:ku��Y�VF>�M��T$ъ-H���s�U�+����l��Zl+�),��)�-Yep2�� �j��ԣ�]��D��Wd&�y��qo�E��U��裫#�HsW��Y� �+���.�c
aJ��-v���v���9Τw�Q�L�uQ�ZJw�䣍I������prɨ�'t�@~�6ϕ϶7��9�]b�p}����ELu ��8I�3Em�����VH���;I"k��?n�ߣ����m��S5f7
��y$e�!\_|t|��r�E�W��O��rA�w�!��=��yA��o[���J��E���bv<#��t��n"��4?�De;��o*�7y��!]!M����D^+�d�/�Υ����v,U��'��|D�8�J"�$5kA�i}*���7�k$U�M���Hp����F��*8�O�/���q9�4�	( 8�00Ocl���Eo؊�
2���O����/�p����q�
�y D�y�6��f��0>��G�W���.��)_�6G�!�􄭍��#ڱ#�(�#�#�z��l ����-������oV�]E��u�j���@�V����Q�j7�/�Gڝ��z�B��e�[�$�vˈ��0u
b1p�Z��|d��]V�c��c�I��s8\�n9�j�2O��Z�5M��ˍ���Pn�|�8��~�*U<I]�����u�&����#��4X^p��t�1v��t	�]8{�C����W�n^.�H��o���w�=�*\�Xf�U�>w'�'�&+~�&Ͽ�z�W�,���Гp�Y���G}�C� S�ٖ�|�E`�L�c�� �C����{8����Cַ����NX��w�K	�
c��݉�#`ށ�1����9��*O���ř{�Έ�yy71�O<hO7Y�\/i��?O�{�rr��=z�\G���Y@N��� 5�B�Vi�v�;z�0��ؒɚ{��Il���\p�����K K��(Ē3�DI�9|>�#��;1�و�t��E�o(�|�dy�9�ჴ~��@!�U�j��`�cD9�=���z�Hp��������]�r�=�??h*9�#tCA�.&��	��Կ�X@��eS�9V�}��)�e��rd��x%>�1��\�%l��%�(�E5U��54e�îzMh��rϯ%�x(%���p�z ֛b��0.֒J�'zț/:���D�Ktիv	I�k�6�t,��H�����6������7,T�!�:�lu�suh������L�� M� ��7�ə���Tgi��(�"ʍ��$&��FD�ף�F3��;O��ev��S�:����a��&:~a�u�*��o�a�/����Rm2���b�GC���Ef�m���_�ZB?q��Y�@����q��*���rX��zPW�mS{��|tk���.y���)��h��O��U�j�������ƀ贷7�/"ǌ���4҉0�?�#~Z`u���YcI�C�}�)�/�[��x8>h�'>��Bvy��|6*3s��&}6%�'�`E�fi�W��Ѷ�K�[*'�]�§��������������ER������)]�uC�� �L*i爚
r����Fσ�:Ȗ�Z:�Qe�kZ�T�T�`���/f���� ��Y�b>�A�%�aL� �U��
H����0���N`_ֆ=�F���Le�}�sѻP���#�?���x'���+&Z0���e&�!Z�Y����x�PT۵rڶ7�X���8(�u�)t��p�����*�83�V��{(|q�{��zZ"���-s ���.�/�.�cs��r�l1	�f�^q����)��Y�3��Ƭ'�'��w���,�Op��Q*�B��w��BaX�e�+�a��yeM�׌�8����Xr�Q�}�)p�%���F���B�:`�9{��.�h�#B��;M���-o���	�⩎�a�d��l]ָ��_��WY�<?�<�9Y�(�r�l{tƬ҇ �&�$+^�3߱Yt狂P������^�����p;�{e�͖%���������Z=b ��ѝ�$�X:�J�}�4�U*$���z����ޏ*�����k��x=�A˹!)w�oRn6�mM\6]��J3����a]�"ot�����nO=��s��b\/���a �]Q�~��ր\�<}�Q(�ׄ�l�j侦Q�>]e2��v���z�� �?-z�-%�'�ٸ���Gm�Mǉ� 3�
Υ����ǈ���Պ��ʣ�nb��`ת�����vt�|�����Qk���
�m�4�`Q�c�������n���Oy�Mǭ�]_���A���������
�������rJ�2��K����q�!zC�q�e\�� �\p��_�E[�[E;�jm���gs�d�3D����ɽ��8^\x�A��Q��1��z����]��V ��A)"��E��8ߟ���� ���r�}�J~p沌�v��1���9}�E��(��
��q�	`�x(Rn��9�\\!o"Rխ �9��E��� �ۙ���1^]�g�k�)�� ��9���9���wKn����a	�� �O�0q%��T u��[+}�[��̓���L�7^x��$&�����1r�AX[�� ���,��;p�}j�vI�����&6g�FUy=�h�W�,���rf��b�3��h�SR�FR�CS?��.����k�j֮~���RH)���S\W�҉,
��m��W�9��S�;uvȇ�� t��;���l|©U�:��c�v�|&���0u�(���g$X�[����b	����$�e06W��{Y� �%�;�<��ی�dw��j2Z/.�J���&�M�����ѭP=b��U7tC�3�Lj�!�ل�rt��f�=�<��b������+?��@��L�ԣ�n\M]`l�_T��RO!�#`b�%U�Q���ưrul�U�R�5�gb��č�`�E97�+����.�+Ρ��}Br>3�4��%�B亟c��LU@��a"���0,�6�	�,bI�N�0��E±e���y�*�&|;H����]��6�S�g�(���BV�)�h��_y�-�2��V�m�NЩ�!7�Ȅ��!ID.̈*�������M�Z�2��SͳO��Ka�PC4Ɩ����g�R�Zv�"4գI�1H6\\|�G�Hܢ}�3��z�}�m -o�K����8���-yEkQ���z��+�����̀9u���^Ls� :�B�����)mf��<��jD�3�0����/��g�i��e؁n$Ty6��0Y`��9��;����O;/Q0y D�>ejy�Ӆ(�-��`��.���5�`f��`SK +�T�R7��ZZ�YnX�5���1���c�4b�L"r|3<S%����C�ff9h`���� �w^�Vt�Z�����J׽�a>�jJ~+2T�At�V�H������ښ��I]��@���с�.R�;u�,�E��f�Hr`��� |�9v[;���g+��YSr��`��p���,�&L0+ e&�rYJ�^b^h���<ʏm9��k�}� ��L�k͘W��:>�2؛���W��P� ��d-��9�EY}%p��Ϣ�ܗ*Y�(pR,KT*�$a7��d��/WU�h��{��Q4b�B�8�r����=õgx���.�NZ���7؊p �{���'i��ͭCX^����E6�4Ax���'
�+;��=2�00��%��+��g$�la{���-lDz�f�߿�WWv�n� ������h�6xF��FI��W/;���wl����MG,��iȬ��2���6���z�gE�z��'+���89T�X�9�ޕ��������ˉ�#N�H��>�O5���K�K���DKe��䪎u��t4��!ʕ����C�L@�GQ	���D��J�����emݝT��7u��x7ʲ�ZZ��kA[�/	<,rg��@ ���e���Y�6�*V�BK��?ٛ9 �_�!{a�
I���3���ݧ� d�Wf@�F)�^�ԥ_x��t9�Y��
�m���j�=~���5,�
qnh"�&����b�z=*p����3����9 4{
#�Q�ػ6��%�����m.�AG����ژ�e�f��3R�"T�!�2���_/��ii��~��xT�W�!+ݤ�Q���kP��˂�~��FԳ. 7�O	�d�5&��|F�_��p"�g�:jQ��bgȬ�#㽳�	�/ٺ�,�˄���Ж�����������[��QY ���wL�XJk�B��@LM�=�9\��M���IH��i��z�'%�a�w�����ۻ��W;h���G�G�����2�K��f���v�^N�g��E���C�^��~�aOIg4�!��N���5J���@��i�X���^[��IU��\�l�*�9�J(�>=�K|��p�"��S�����x���B�Wr���͸?�ؿT���A��P�L�YDD]>3�����)��CJ�m��-\*�E�� �T��YH.YT�0T����;,z;ÿ+�&��m5o
Pa��*�I1z�߹�%$���4ljE:ܗz^�Ѵ�6d�L97�*N�<���|�>��־Y���^Uj7ʜFi�$t�P�I*�Ӑh�3�9Cيoȟ_O�7	7�D�����{��B�;&a.w5s髳���3F�'$;tE�m�/�6�:�����������ɝ,�b�S�����Os֦r��bE*��ðoP�p(։�,+ʎ0[iYI�����.�����T�e�]�8hM�a��Ҡ[
5���7�M��|���}��c��a�޶ ���h��pLL�Ir�c�s�c;�ti��] T6̱��+D�U	�����c)��nH[j��y�t�*$��>aYj�[T�y�A˧o�1�f�uc^��X&��Vk$��Y��ݻ��C�f�Yvo7��B�݉��e�
d�l�	1H��b���
��=Ģ��sΊ/��e���n�2y�c�b�/c��p
>��%)储{�Y�Y��R�~�s��2 �&��]�~э^��R��Z�x���4;�7�!����g����Eh�q:��u������P��?��O��"I[��1����[s �֞%vob����/'�C�����+���X�����[�X�
j���b���|�#������ﭠk�����*"�����)d�q�S!�B"|�		���/�pD�B��D^���)K�Kc�2P�B��)��i�Ft�	��l�'lC����c@z�JӾeclXJVa">7�ukqc[Oo#Ȑ2�m�"��3��j��)x�k� k��<L���Kދ<���^��;��s�����{%�`lܼA+��s�����,A����FT,j��rX1�һ�Vre(�4,��g-��,h2Gu�(��d��>�8f��7��=Y1�{x��˵�B'����@���r�H~�ؐ�yě��z��vJv%�a,�*���E��� Y(-o4�\�M(x���T��"���')+Ќ9��VV��62Q����{$�
�{���d�VN� X���$�˽_��e��{J^)�7{G�.8D���5=��q�>�����;(Rr���~3��~��=��AS�`�p�~d�T��Zc*���#��7��'�@������
z#R��5�����̃~�������8��[*��\��x����-͵�����A�g'/n@��<ǭ}vz�^=ϸH��WƲB�n(=I�J��؜�D�ei����Չh��Y��bo�m<H��,Qd�!�ƚ��G�Q����F����ȹ��ڟ�6��"��X,%	���O�P�����3c3D/&�����̓��3<s�֧M. �/ b���黍�X��6��ޭ�L��F������oq-�������˲�{��mW��5�{���w�3.��Z=i�8$��(�0�(���.�F��[@�bDZՎ�>u�~��$��'n��6kdS�U9E�}Y�: �Xk��c�q�Ƕ\���o�#�?ЃhG��L����v�6���sd\F����%�B[R`��;���=�{w}R�
ow�BdV��f(����-�8��Ճ�(�ȇ��$S4�����m���k�Z���z��˶�]ujWB�1�˄����^�����Ӭ4�9���e���q�ZOfs�3�p4RR����IA��K�O��4�����y�ܶ�E��sC�.����v$�߸�V��_��x��SFWQ��Q���lb�4��Z� P����7Pb�w?c�0��y/�V"r�j=t8NZ1�ƶ��X�ɽE�F�s
UG))|�W^޶b�-��N�Wk�ȡ	�.Z�>-�ř��I��!LkxB�5(�{{���X%������o�����d�G��0+��b�O�ݑӰ���o_!˃�!����++h�r"E�	��~w0Z��U��8�T���˳�?�+|fv ���i�$s�B��|E�=Y��C������i���l7�H���6f�Z����>�`�4.Um���<o%�#A�;��ΙK��1ɥ�_LJU��YW��7 n?R��.��S��ė��<����?�6�,�ֻn@�l����v~����fl
��p��v|��5T8�,�����*�)��ǜ���[$�"��(O�����䤫DiS����OUB'�d�R��e˳PjśhR�4�P^��
�Y�"�V�?�:l=�C/��z�|�VVІt����\����*=�n�]�z�sK;WJ� +PVv9�S^>AF��iI3��Hi�H��u��O���Y옲�M�_Y��|�Qp�1n<��o�j�HJ� �"-�i�
��u���Y �]/-r��,�1o��w�����1�Ъ�\�����l�F̪+_�p�O�RݫƶR>|Db8`��f��g"�w�ƾI��d�]H}aQ,02��oW9�5/XF{,l�?�,j\IP�+;�$ĤŤV�.ֶ'���q��ԃ���-�̹�ؠ���B�Nb���g��=X��'ȿ�&�q��Qb�����_�7'���bJ)�87J| ݗq)�(�%=���r����ݠ��9��
ޑ%뒊�qE�z����d+�U��\T�5\}y�+��kf�Q��Dxo�WO"8�˺���h�a;{r�1�p9��M����v�K
k�˙K#)+�JǑ��}:��D��)�Rj��+^n��ˣ�.i��}�6��֏�
a;�0}�Z�OK�]"���>��&�窐���������m�#�2��T,�rK�{	�Ϸ���+���%
�$�ϟ�`�f���_)ûH�p�M�SP/�5=vw5U���P��F��9+�ut5��ּ�98��[����Fa���2]�adS\F�BEO�4�(e:�_t�q�o銮\^�r�6�M�Ŋ�^~��1����NAǊ���aze� @��fh��E+.�xb�wf%_���xL1�JEEeb]��e�A��[���A�����=������S�\
��s�)�^ؾ����[�gg}1������ g3�=��2K�L�þ0�w��9f:s;V�ք�/<��)H�w舌�J��^߲��{>..D3(?��_�i�M*�}�C�F��I���U�Ъ�d����j���nE�B�*���Vj4�r㦇k�U|��� �/��{ +����P���0.-Y��2E��/�����k�8���ю�'���Do��&��8m���E��Ƃ�#�XSg������"Z}%��E �k�
`{R�ڴ� �Ė�,~���J�h 2��5ok������S�h�gN��ۧ_������vI�z���-I�{I�l�!~T��P�5)���/��J��OWy� -G�Ä́��n�q�R�B�0��ո�;\��F-p�;����AMi7q�
�t�|�z��seO���0��u�Dr/�����z	������-�����(�)@�V@h�柛2�죠���aU�xw��{R�qV|f����H�<)�G�Cj/���מ��B����C���
�sU�|ǩ����Ƿ9 ��*�����c����n������H�ɸ�*o���݈����ڰ�&j��P����6sњP���Iu�Os�0A:�b�B��:nl�W����8G�r��kH�+#�QI�3�pX!6ـ��!�RH�h`?��nkmh�hR�D��I�_���O�MX�"L�j[(K����ȇ���sѝ��`j�R�K�Y��V�Y��$�[@,�z;����uh;�@l�GEi�Q��,������b9ٸ�R��Db�K��c9va�.�L��9�[
J������a�w�`-[�������!�f,�Ld��3�b�M�󫋱j)���y�T|��#�z
/�a��E��g���pa��K���=�:��)���τoJn:ʡ����1����A]�¬mU"N��
��;=���i�a'K��m�2M�b{TJia^�֯n�#�%�v��;���k�.e�ϒ9���:�q��V��j�ӣd�p��CW�RGSj�U�M���_$?���\�y=q�.*98ke��e�%�m4^��'�k��/�] �<)w�����J, \��EJj�o�~<�6�nO2�*��*�g�ШQF�Ljk�tO�.wmYCz3�ҁ�ێf���Ҥ�W2�_��]�L|EHϨ?��\�u��4�a
ǤW{�sY ��Ű��ia�c���B�V7���=�(P����l,^���w&,^W�M�T�P̰��- �L�Crʕ�-n����RW��x��֓ٞ~���������+��J�))������7l*��\n�NH^�1^�4���yT�N�x5=��Z��k̍��+�d��<�(�N�F[ j����T��򻷌o��w��S�|���%�^P
��Hf�#�<�4�R��\�j��G�FXo�����@�t ��d�]��r��d��1$o�h�~+aD�����G��嬽�z��-@�����L�RA1�~�YE�F
��C��3Rdt��_�؟��V���j��d\��J��8�����E�Q�F�59�oݖTd��!K��D��]Eͩ�3F�0�<+0L�|�&'?����S�64cL�m+A�ޚ5�����Z���[&���@�F���+�+ع��U�ۂ�����Fq&���_�.�Z����]�v��&u�d�wӪ.8%��q�d�voZ:�ń���R�R�^�8�� A�����ބW��y|^����H)����X�\���D�u�s��!ޗW�c�S3E�M�}���Pi��wG� 6�3�i�xl�O��+��x�?�ڡU�?�=��^��X�ex� rw(����%�M��2zhP��DO��4r�7�t`zU�se�͏n@[p繑�&g�@����9�U֑,�8/��n���ǽ��
60ɕz3�����0b��e�̲� g���đ�>Ko�I�g�.{4��x6�X{i�N+�>a�>��/	O�*��i[���6- h�.�g�_�Wω��$9Y0JJ��
�ܒ����Zk�z�����N�ˆ�0�V(z��)jG/(��TG/��g����|(�NS>�1'�p~!�@7���Z�����)��e�������s�4]��헚� ���kX;�"F>ʩ~���Ϫ5���-R��] 4��VՍ�^�����q�V[�}=J�w ��w�N\D���ŻT����R]csֹ�,����~͂�d20Wl��"�*q�q �7���[(��I(��#��搉p�����Jꐧ����Q}��C�#�g���9�]TX�*xUU��x��S8�ט�u;�'ka���R�۝�=~�D�`0>a��p�n>��N�H�u��I�����yEo)"��z�śccV�B����`L��v�:X�S`��'>���Зq���	�hgH�-YH�W��}P��~��at���M^��S���������y���cR�W��%E��&�Z��0K δv�"�{� ��VJjc��ے�T8�aMF��i
�b��˚!��'9&s�*�3�9L����DN������=bP�� .�[hܐY�+,$��ޓt�jA�❂C��Sσ[���y�`��_/k1d�����<|g��0������O�<�,k V���0?ćuȈ��?�L�PU�υ��U���/���h���A��d�(<��y!��Ӝ��̕zY6�dY
*P��`�9=�Z��W���l�B���6������t�C���Q�Gn�#���ȭ�9���W����$gzVn�X���+z�@H����k��w�M�<D�Z�WLH��F7"'�uـy
�E�.%�I��_��`N��u�5�7�J�	���.Tx��f]���S�ԍp�ߞ��
�!�j���mW-�]�Ϸ��O]�|�@�SBE%C#.'���4�p�?I�&Z&0˒���qE�ȂC��\��_�XC^��6����x/am�F� �ߘOx��7'�f'.w����07,_S�/���lK/�\�l}>����OxX��oX���?���F �y�ӥ�	&~NC��9����	(gCE�L*��v�Mp#sH�''h��F��g��R/J���W>E[�{$�z*�1����-�#��r�d��{վ�ǅ[����~���n���*����J�n�vj�"S��=��%+�n��Э9*�&g��_�z�e��'�+���t-� >�*zȚ=���^��I5Jֱ�)�V)�r��m�	���pϣ�O�4p���Un�S9�_F�	X�J���Pm���-�>�^��!(�U��3��A�#��	ѡ�n�XD�f"1�#��ӃN�)y��'4�T�Ev�W+����+UĜ"�/�-�7�1�"J��@�:b<���L�ՙ�O�G�fI�ob�q��R[�$��ཤ��6�$�v>̇8�O5��:2p�2vgP�i�_���~��̉]��C�z�^\���<��'���)�AO�����k�rnp�;4��ސ�w�&��2��?�KCC���$����ԫ��^�|��eI��D�ӊY�~�O��4$Ċߑ�7v��R�n��aW�������ݾ��G�f8it�"����u�`=r"����ލrX���d����hr��ן)�
*3�-�d/�=#�\.u��{�K�\����b��b�,����y8t�C<{�=<N](,���?�3^����2��y��cE����#_��l#�t<f�j��Y#g����Zr��BEI%ĸK�W&�p 0�0�I��AGӷ�o��1mv�.�M�������h!H;'~�Md_���w>ӗ5����C:��X� ��-ag�qOJ5x)s��1���5�_J�r*�qјs��L��]�S�Vhn�H��")>�&۳M˔�I�DZ�x4�B�i'�W�F3��zB�<E�,�Y�a��i$��a�і��~g?�\��{���~_�ޮX%�ɋ+&���G�B��Z�l�����i<'�L�e�d��Q)�^�H�W�W�&x)-C�o�Oqb8�`����� ��6,˖{���E+f#��R���/U��	�߷N^����Cd5t]�\�����Y�jGg���ݺ�?5����b{j?�4OCğ|���t�������@�M^��`-mp���@ �{s����Pg�G=�f��\�߫�0��E��������XT��`�1��5Hى��PE֐&lC6662�1̾�苲9�(����2�f�ڢ�iu���
qg~�vu����k�0QI��`3T�q����R�'q�HЅ���u��N�s1m���*�N�>^dD{J��������"6rKT� ���Mˌ�WZa���ӑC�'��ME���E�
��VAV��-!2삗L��c�
��V�u��š_�x��I')h��^���|�W��H"U.X��Z@H+��W���q��y3�:������]��\��0��0�./i�ۄ	�fA��_�)��Q)`�)��Ϭ(h@2�=D�wz���md�Z52�����$إC5#)c�fӽFa�7PT/CM����ƫ�p���;/\�eB�7Kn�k�3%����E6��tl+��������#0V�]ǧ��/,�W$����}D�¥�����Y7D�Dg��@\�95��h2�k�(����'������dh��N��4����6��{w<�>�zQ�����3�\e��ґhIL4�h�j�Pwj�O.�bێ�uhJ�ca;?!O�+@"[�ؐ9�������L�V���v��҆*�D$�~����Cmn&������뎂!�.'Z�ix9�2�ڽ��9�rYH�6���Px����w�������dSsb���y,̰���;����w��}���9�O�h�"=�����X�km�lʚ���ٴ�����`D9�Zx�cx���H��n4��>���x�ȥm�7D%����D:(�_�E��u����H��O7��(� ��v%�ޙ���((�|^��:N69�+x��=��Dx�á6Mk�ИA�
� x����,���V(P����:������&r0������
�� @���A��z2Z�@$���JC��+8�u5�QV�D2=@���3��z��v�[տ��i1��l":-һ'�ݩ#��'������S�o�*۪��N�JPVG�̰��סw�s���i�"a��.����p�3����a�a���Vc5%t�Q>3C�t��;�����Z�S>�/|0v^�|���¾���)|��DH���Av\�3Ý�f-�u��,~�Od׆�n	�Hɟ�*.cW���>ؚAtu�P���(,��l�;��V..#B����~6�+�B�5p��5!$�L�����k]��۠��;������`�M���ro]�d~&���	R͹u�ld���fE����'�(!br��>(~��ނuY*IDByڨ�",��+4�vA��9��z�*�,�y�H�[6�l��e���v�^C����d�f�}��ѩ޴Q���x�Jm�1ϒ�nA!��8��oUFe&���#��~M�a>@��\���]3O��±QK;6)e�g��Y�S�|�kJ����`�V�VL��'E����AbZrK�4���Ӧ�����?�"���\����F7� C�P74)�i�9��<��;��Y��,]�1�ʏ�T �%�񡻨bk�/�#�j��R���ry�]�i�.�Fd�P،@���]���CوG0)��%�a��U��G ��2Q
KY�7|��`�whq8���5mqP���;_���<�	`F�B!�h��a�#aT��-�eb�����<�	������ض6^��)����˯��