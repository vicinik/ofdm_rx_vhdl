-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
X8O99sVX/ARYcbUmxFF2FvSes/jobXv/zIzi1e3deLgxqECF8ew1h/g5aBPeHnZV7+RWJBGMv7yt
niRQbplkhfJBOA22pK3gnGj2AzU74ssclTbBdESjMXGEtMXEUynQ0dMJlCX/Zck2bTj/Rv/42hjY
ygkp7nPVe0euEp0wqjKUDKDA5ZIFv+Ss6su/cjEDTxt17TXaBfLZoVeRNMDq8KZhzRdIldiOiLBY
dLwBweT8lvhXaayRqGbF/0CmOqKtFfkDJs2jfBcj+BBJRnp0dXOmHLurh+v5WLxJaRhF55PgDe/X
DMVHq5EvWNYCZKxt3ucQvJbohxZtSCHafpG0Kw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6256)
`protect data_block
b1VtdTlz6OdR6aLNFMZBUFcCAUjvcjxiVXYjdWLhyiPjSf+C04aqJ4vJ4W6vprmP7vQ9+ZwpwC3b
pVjUD0cXplyVTqsKWe4xMI0ejAdyybfootctXYj1vMpb7yJP5c0Wy6NO6rQOEv2HMjWXBnIJCsL3
H+2Ku3YGwR/Ip7MFTzbLdBWKqd/c8sRwmmxa3Vq3A4RShfgRMVQcbC83nt5g5KLDe5SfJD1RgY/k
tGT9P0Uq8eYxRg05UhkCdn575Ueja/jqnmUp04TpU6Xxlt0oXJA+lyZqT+0hnaR45LsRaHtiera7
9TPU8kbv6uhjP1Rhag7ESL8U6v6/AmmAObyjm5Q+ipHyH70j0y368DL4nDQusKfWR9RMCs0feVK/
1kRV/bAhevqWYKzVagYWLJtW9XeGVKXAq0fqS/ML5+owGnunTF2GGM6094AqdkhiGEem8s0oRn4N
RI0MGk++QMH2V9r7wRgO4P94V6s4QT/IHWHaAP994SP1t7XWVh+7enmHq96T3slbLMBnqW7kKs2r
qTdZ2ELioP/1vn3zV+lFFqGtrqzMlDpt0kRrcnKW5SqxjPlg3FIkme00Lp4OiGNKjKqBDRRh4W+A
4EN/hC3hrcQ1+zHGA8m8F12VoDT0reCEYEDc52gjDL3SwmGLhpZfORwLSXkT9gEGTGqiYShx/dEu
4i8PUDhU87jSKhFDPmdyZ4cZg7ZQuVhPY70bgfbbBlXI0canx4b5r4+LuRt3iqTDOnJhokkfYU3d
ksJb6ZMA7M4QUj/IR1X9D95gAlorWQcJcbavwdsJ0SpDB0UyLc9us2dKCKd8TY7RO40NO8bk1UXe
MsamUsM30WefP1uTnkzh1L9wj2EpuNHRYLSPyr/Opf4DVOv4R0YEcbjvj9laYC+NvyGgAWMrbHko
cppuIoNZ3px7J3tLe4l9oAyhvcHf8slXajxakh3XitxqxayAE0aqe4/J6m1ir7tzEwhFLaXuSdXP
G7Y1y547UKKFt8MtqYhyIOmpbBshLvSvepwDl01Py8kiMI6gJsusa0JmSUhOVSAKEOAC3hbhIyyA
juwZDArIcCFmFt+BZISI1Dcf1p6dC+/zt/SahTzmjY9sLj0086r1v0B6gR+BlWrCEQbP0c9Hy24b
tZtNB3rtl/RbOVa7EIeGmg/PSfW39fPMdTM1pMUy5nHbHX+5uOQjHHzw2jKu2WF6w4eQ5rVv32He
Y4WyaBYG6O50pmQbY8ysdwhj+rhLQJ7xJ5bD7MtpQw/JUFr6dA2Leih+duGqHP+tOfzw25CKUwma
tnnvoZLMJEqGSKTHUgpD1IdyKVwdBaacOuZsa9WvC1f7S4VfbC2dIGVa0ZHlBruJzlkOUWDEmkah
qHKmET87lEOE5tbzcuKFx/zBMjfd/5KsAQYlWWMZ1U2ecmoJ9YydNiKF6qIQE673lXx3WzcXAgzk
MpSwzjtma4FoRu827BndN98nd5c+fWvZWUFha6fPJUX0/SbYRobKq+Fh0UYZAXhejfOioi9IfsQ4
tzigtcwx5dLn3yDpEPpENdzysl86x3Z7DYLhaYagNeHP1LumaUCJhMDVK0hOZt6T3btXzIc7hKWh
xAZjXGVikNy68CBvGSvUmufYm+fUtIVwthTL5Bmr509jvxIed8aRbEDU6AiixBtqCwyfazcGKgay
9zqZ7edh0PeXJr/HK3VFT5vmIb5VKz+uccMKv7YiWdZTfv8nqeOyasK1ZTBrs1/Fi5Bp4NWv2Lx2
NlIt+ObGpXmITG1sGvf/dE4kUWVfBdWEDuUWU1NA5J2KGKp1zvwsID957N6nJObFocDO9oYUBKYp
LLSWpcYw6nYoV/9E8zBNETYWjVf56HfBX3XU67dGp3eY1P959lCw7uKCFjkg7W1FZV8+yE7TOL+Z
GG9LtJiCBqNFxMiBsF/fxMJVOMzuO8raiAYwkY8ry8CDegnOdILKG1Ua2sBBexdM8XIeqBc8HJnJ
WwJmeMgRhcFbi+HjkZs7/onSZxAkytvbwhM7KiC4hMkbmyLgvOk5viQlp0gpn1ExnB4HZtKnMXfo
EwSSF3Da9D3B5TxTFrU1/i2DvfnZ/OAtk4bUvk+8Plsky0QbGylEVfoFKQwa5/rlk3OiA7ckaQAU
b7AaFVnQcuE8QglvVLQFKe/lk6n8kG+hWIljOa6yj7+A0oVZr/qNmmky+w6RXt17D67KjnN9f6iJ
O+E13g5Kx62Fvt0lr4iJTnbo9bhf/TTOVkMr7uWxSpoPbuTV2apn+GL732CPt46u3bDBVaIq9o8v
ZVdV5j8VigwOzxsd26BJaWOtujY/lxRHmwiJOmEVqTjpIA/lRQlIrUVNzL7+dqwr09uJBCcB5dkv
lSYCjnSi7RHADbsluY78t8vKvRjUlKzjVO+J5mxDoontkO39ZSaYymykxS+RirP6beB/BGpEHwx7
3hY+RdpXMiVODCocp63xuh5Zcoi5SY9rsTiFnQjwhhBV9dFdwmZVdIqEr3qgLJBN/xxWYI6/+poe
8hI0Ba8VCt+m9iKe1yD63izocZXExiLwjQP4KN9JPxAcskSWOnyzzgqzNxnR6XTtyZRKpsPFlFyF
hclcRtrmsKyFOUEoOa6nWB6xRU3Y/Lw2G/u2aesOxzuMnWSJVmDxQcTH2zSF3Il3jL9l1pnyV3/U
TvptbTtT43Qatopo0UPZTqVzPghgzTjsWIP0oeqE2jW6a02ktDiqW/CpxPHE5Cqx6g++ecmmlJC+
3bwML1BZBbDj0pTGrP4iRjITQ+OisA/HWt2Efa/Qxbbhi8YuL+9Ru1/ibaoeFXN4F5pQ4BcY9OyW
89UIpYvrSBopJhgJaGN3XkNrGjRp/P2V/4OEoigxSWNdsp0mFDZL5ZOHuiQksBZHQFzBEgluCQWO
wihfCxHgGMrKCa4d/nVznQLKjMe0EfUDS/+U7v+UzhjfygQ9gqqA0EfJlYF4D9zehW2BgaRHDg15
8a2hPKEraQkuaFBS4hWYT1dfGkX8Lrz25JRJfuBSsA4hOgh2+KaKKmSi+UM9zzHVkLnOifoB02IU
btuRYZn20xF/+oJkDygcpYeziXzz+HgArSR0Oypbdg4lqeOj7uooVAPTTtKXlqIPt8BJiVLjFjxX
gZ9qY4kUyyr98oxTuu6XbTNSK3ADb3mkcmr6DfHxzXpwHxtNmfQAwjJS6VJXMJcV/i2ck+dUNcyw
Pr+Dr7YePWEm46rL24O+3S/+jNT0dcSFVaCRdnfffHQsGdgnPbLjzlSlBDwl7GTd+pzev1cUmQnh
c+W816n7m3Ktizk960eMvNFyQqUa/ObhcaYxhTRzkOMXjiNmZsJ43FnAqL8toDRAGFWz0dQKNEF1
0ria5QZiXImOanh5RaqCsW1PR9JutBBrscKNBtpjjfcEXAm5tbRqc1aE4NjboMx6pF8XmaIaRGMG
8DewFy72TIWl26hPFAoiLdTdHvMdvHxSt3IxaiJ+hulQ9TeDm2lKVp6vuQvVU1GeaWDpJLfUOyas
HkLWsnTXBYQl33l2uDuWiqfd4VUomoPSrEssnA42cin2AvsYXZMlhnLQJHIRLzGl26z46c/Xn61c
SSQcL5w9O2M1j5++nyjgrQGCL4UFZM297kKUJCB7XKW/NTXMrr8eT1WWn3x+MUURq48yXGH9UXoQ
kEahsvauvvHI+WhRRG7idp4GtDdWo6+LOr3W8DwbcgOrtcuNT//9+czxznAomS2T0cYkznUYAM4D
3ZeFCZGy4iODEyjCS2Z3aLkHa8jQjDAeDbVUBlxESLX8wezvKS4hW07m1OHegL4BsbDZwB6Xe7zI
ILtQcRHJeBJCzVkUADgYjNH2BcFCoQoWwyA91Bt887b3SSyZchc+lXV4yCwPtcnpaWbvuuTPcff/
Intdu17YOAnfmATrH4MnIt8BMfwGnHKDDZ/xE52PfPl3yF2kt8elx2bGAZ38PRUZsyzRW7n9ERwQ
r4maaOZnoKBYGMxLmunVhjvZFhqBtDGA4VAbgG9hVke2tx+3PJwZMq+bqOZ93wVpk93CSl/AXqrG
aLB+4EoWtqzaqtEaVD1J21ZFOVXLJOKfX2laBG9MYloG056Ai75LTOuy+ADhLYFLvKN99a94z8cH
VYOFJPj7pwmbyd6I85o8KU6JZLFI/UmhAwZ/3WCB4VnhFCj40ZMckYvgDkL+2S2VIOrkAbpzXdBR
PDmghiMp2hON08Y8sgPULdpi0eHAGmgWHUBE+jd0LBeTlZsXg5tifiRelrNtMQJqBS4gcY/p+0X6
yyti4YydG1QKwKZmXkUNEBjg1BixMV4LWRE2BadPYq6s9k5P05Svi0hzIpGe6L3IWeEemHIepSx7
HdsSg9vFhhWn9ipAy20OH8B4hUd86l8Px7QvQDnwtzi2lCCiYH6XhELb9xJvdcZr+wX5bmA/ZxGL
Np7tGu/bwNTlSuumSYeh9Gt9JwcvZnRDUKa8aYhTGJlw1o42NRMwPEKsR/bMdRnrEQa8EZuAqmen
Zj7Nv+m2TWqZUFmg4YZLxwI/VjXIVnwX35tL6RwDFaRBqOabc/TXXfTJY/mOi5X85tbLTM/+Kzze
2+IsClHEXR5oVi0pxfW3mGrCl8Rv56WkvQeA+/LkkW3raMPKpSVoFP52qIDJUKOSfw+bCKsJH9OL
ZXpGQhIgY75T5jjQ90b4fsQ299A5Bl56G7JfIhzXzCpB9VluGXGYTE66XXHWYlnU8xNVMy/HIfjC
TTgbfyhm5mtdbheHKqxJCa5XkfIF2dzG402UYIaHG1pQlCm3gijTOf64s3h+Qdzkt0BrBfwaDFxp
tiI81PA8UWOogXaYn6Tj/eJPAURdPLOqArlxFQcHuQDsu6KcTyXd7iQHhtFPzV2cSPzSNH4/4CIk
QyQj0DmRanAOIvKLHJHkti/z9AD+0VrsqbsJnLwhSyIYjcrtKh5s6QKj88YZOvMNOEpML3Gq075z
EK6/47xdQGibesuiQYZhQ1sqn3/aQ+atidapnT2aU6TZYwQMsP4p4Fc0ms2eT4PdZh4H/CB375z9
3kN3uAIoJJBwg0BFmEZQV1PXVsbO/KF0EkeHUf4k0qo/56D6w/to8f67G/3oUhGwJ7GOuPHrtZhm
WYchk0mSNeY6P19uPX6DZDAHcQ2u7izJSgHQ7fQKVRMVEPdegiVR7Sf5Jr5hF4usY9PTcX7WP9cP
vO0N2rjem7GIDOeX9shWDRzdnTAYkX8bdHFWD9GmPA9PmTro4Z9igFENWvOBhY3LG2aQiSWlFLzl
YtiPc+usXQcMJr6D1kyQeQg33TEnfpRinz0ISWCyThkYV/44jh+bJPCXsWvU7lnN5vtFIpWdQ76c
WWPphnkRwtdXZ5LWJZqhMSeuLRsMpB/Ie1WEB9/IObAy7tEjfHo8BlZeLrMlTveBuglrSt+kxVhU
eqHur0LqxVW74V6cl7asRZMP1trPZBRYSiOvfv5t1COMUXD7Veb+9vgZbXy6NRYM5RKfmFFLmetV
Xj1PrQ/Kg91PDmkUNFQ4Oq/wu/AMT1PhN/p28QQlmzc7An5bX6rPH4Re5EPild312uxYo0kbGEuq
JiBzAxbKtJKwrN7HTunyE+hNzdmZXq6cpUrCyG+b/h7n8XE35iSyXTHQ0fQBRHRg1YbDLw+6I21E
h8rY93fHYRyExpQExE2UP23EYSWgGsUF8AyKHoF1qsHwLO3OhR/kXZyTvDcciTyjrIyO1dvjUm9w
qooN0PowxunY3FhxKB3f1QbIolCu4G5eNvz0Z/YwWA3NQmw7GNCWGpq4oYAhIHgxXDqDfVurt/m7
iGuiSvzd4pDuzsACqeJiIP+rkbE4FKbrq052uPhEd6Oovrd7sFqMC8XqBX9XSn1vZR+nHPLRnNAX
PyLBRUzyU2TAZxZubVKt1PCk8U87F9vlvNZutH1C5IgzoC5CEeoosETbF2crLba54ElLffhjAcw9
kzPOEmdQfruqFfRRlPkWPVr/JBWznPpfb9y9X8FhFesS2OmFUyz2qbfXUMxUOumE0B5uzDQ8jIzZ
v+8GVKDffNclq67R2eUboBXiwq/XCv10BmxhHIcN9h9hkuTvwI1crLIWvavsr/ePanWHZO/wjqH8
kYGeQYs4nsRO903X4ylfznQkvnTitlPKtgASRmgjZtNuaeHec9RyZnU28xI4ClIJ6+MRsImbBgAs
bQzT09HzGwN5g1pz6oWizl/NPc/nvE+WCi+/RQCNbm+pVxinYcY93UT58O+jj4zkWSKiVl35fNNo
qNXr2/V+nA5yaMob33kLzgefxSW+hlTGaCb4+1kdWw2Dgjlu+n9wYI2VSMPaKqtYp7c2soNGbMSg
TfpaPcmu0Y6/b+6ANp5eoUJ9YMwqKxURQlCyGzs1ePBvdTDOrVTuelxmnMa8hl9v/Qp9MsQL5tVk
GMno7yPGV+Zt/yP/ObWXyamGQKSq0oVYExeRjJB1lOtwfakHeuOJ6F8LAPzmMYdbXDg69qDj+Ch2
Aj49Lj5JcdckhIbLfGdT/PTme0ofp74OFWl8nH+rXusXocAFNDye1pLFcxVUvlOAyydqnyZELl+d
aTZqxxb9b48PnowRViAjGDvxNuUCSLbw0B9F6BDpcDIOmmZw84ogfJz6qnnxLjAyaxQDg4wUtUUs
QJB+oX5cmu0AP6MAZhwDHQ1yEGftToB41X/K6+xtUtSxEO0rukLD3gHXaPJEDGqD8Z7mojS8bywZ
DIvP57N79dmCanG4RfQhuNF3BZ1rW6DbbovACddA1x4z+y2+1nf1XmUdX3VmO0MtKdEogISgRfcA
/Z59CUcuCsFP9JUP2sNswIvRSGdsYNxY2XhiODju4kNz10yCAFPFd40hvtdTBM0MbvelDFq8bcAZ
U8PrSHC1nteH83KohqRt7JFWOy87yagx1bNWvCR+T9rSl9oIKq2HjPV22QPRfQsrYEnm7dqjHYZY
rQwGwvsnec/tl+rMP8cWP05ga9BhipTfguY0svtKx46QfQYGJgmVZAR+A9ZFtSXBKZDJzHB0JJC8
bIqte+9m6UuH4uhHSc+I2V/vOmU5UIke/yUWjX0dz93W4AyeRne6/fKmGXRYeusQG9u2+WQy8iv8
YUXIlLcoSyAYwnY4Kfb4YFczW1rzEdA1IlEwrVktAxMr5U4qsgJs6aE6sCGlpAV/O9SmZLO77GsM
b8c+R/BmZTp6RI+gkzLD3wlHe6AbolkuaK9fjDtwXPdfeG03WmNGl8/CS3ledNan8FaG+Ik1l7U7
Alfj4IYbv1YsBjWEe/lXfso9ruJQXUGltDq0J8iEvnNxNWdJDOcny20QbRm8tF41g6bp4eDeoGKQ
81zDPKlZ0J62+y/V6al2eD2jki79YZu5A9SfqADSc2tZFVVMOs6ktw41Fuj8IcG8mmSEvEX58BYE
99EKccwD8mxezKvsQrq+NJJe5A53R4nr6hCaGo4WJ8pmb2nLz1KhsjSgNa0+Ek6W5bVFg0kkqSQU
kChmP9sLpgGmzjO0D1z9pinUYy5dbMAIwtctp5ABIdtp//UyAHKhi7VVSAuqKiY4//L1v9e2hT+j
0x+JZMguhte8dQsXav4ZgBlyzGwhOqjwCxz+UyQhS73ADL49bcYpjPP3dDpcyd1f1V6Q8W1VYGqv
tJIJTMW+QMfTgRa/sMxyeTi2zHmYMS4x6Id7x7EYVqdPPmvatRlX3ef+Xnm8FmY594UTu/WKVG/Z
GsPcKLTHIW2TNecv2muPfJ+2esCX06/8faFWVmSRLPXlVBO+OyFc+kx5YznYt786U0MKE+hfZxqe
tiVCd90lv5BOkLAdC8Ob7Wz+q3c7aDbZgV1JejpZPomR4blY4yn0TXyv+CU0p44/IC+F44c2isJ+
XXxGZEyZI5d3a/ndqTtmr6toZKaV6zF5zJUn7y5k1yH8FlFrym1kwOVBr+n2WccRK2B568eYWtdJ
nk4wEL+4vxh//Bg2EHHXUR85mIoZG/zaQ5oQNxCL52BQLP4VaqnO21gPn0wwIJ2DTbx9eGskaEQt
ze31B4m77i8sr2z/FsPbQLAGXmWdq9uW08rz1/3dK/p4k7MmK2KgFzIhj5pRqZ6bXis72PV6nnlY
3wKG7+zqJ84krJ03OFOwdz9I8+j00A156ulHrmPs5Rjh7pSSHGKqvJtTqQtyKcrIEVOWwu5ZwTRh
rI7xUIb/TyZsKxjlJYS2BEcPSMAeezdYTVUfoclz+0oPfj/X8pwtZBH5R3aVnQfvhSk7RuU8TxGm
eUEwqkAFa/j70ekfieAwAgOUwFs0q+bdkJvZCzE+SOgStPWgUHybHkDtjmhg/mN1G5LNF50p12YO
P9YmyuReKONWbLfJh91As6L/Yto5UBpBcuiZDbIddUdy0nBcAanRdqt5iA==
`protect end_protected
