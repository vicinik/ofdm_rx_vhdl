-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
f37M6dJsk4bTWy1it/lVXZ2JL/sZyjQYn2+Ti8NSI0voKvlKPvWNcq4m7sF5r911BFEPOXuJA/Pt
u9NHTq8AVnzM+nZGei2bZEGZ1CA4xlRhsMdRwPjeXyHhE1fGyW65C4Tq00mbgJWbwGzFF4Nh7xAf
fH20XDEnaAzXittzte7MN0UflRp+rwOLCa/S9/DKKeDgXTEEmvejMzaERkZZEEgxzz1zsSsvdFN9
F0jkma3OzT4PckEeSyUec1fOfD5XjN8iXJHCtSOA7gbiQY22yaeG7IoI29saNxNWNhmhnkj/g0k/
BAFxpmworDyWjZCvMnXUUBLyDcKxqiJcWcQWZA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 86768)
`protect data_block
GAZ1+4d/7zrTuVSchba+E2gsZCJ0RYAwNaC+NCJQF5w1q8VIG8nYnk21Q5/2oyBkX9i33YY3IdLY
rgQ9todwS95aqOEa+VvpEdtywIloTw/R6kkOrwitvGg4eKtZHKP0Q6d0GXjCfHLanxuD54y4yyEW
EMCzkPXvC09xgOgYwKaZIt/fudtIMxvjC1uNHWQ6Uy6Ggt9u9vvnjh1DhgPm45Gs7ljhOGiwaQiz
+DWRiov074NrB5TGU44fQmWhyzKNgRHcWCwTs94PZrhbZR103t3J3RyKxPlxX55VzsLek3AugPt2
idmlPLrKBPN52sP9n129JKfYypiyZwmORV1d97evA/vKSH5dHed8mfca7NBX3vHwsrJ+qUDG7XMP
OggbqiFdNKfigr/u1pK7NsabmTAZ/hNmO62FHSaKsZYmKDc1lNmaj6Bqc9PvUh2blmekcbm7+4+i
MsJoG7Dn5ZWdVvswXX7S3IYdiAwHGIw+Sa5icN4BC5hcG5rXWB5IOI+UBAe8xromer70CCbtSoI2
74AJPVhUx0m4TUduQeJlxszt6lXD0Pn8nVoxPzeDo5lh4//9G0xeL8XXFNuJaP68q6qLaS4lVfp+
FuOfNbD/sOZ3gfofflC3c2gvWRvDKDP5+ZWYnX+otrunwtbHU4FKQFJPA/Fo7sAY7PhFhzBg2jBy
innFHinaEjo05xpZf7IhVYcMskTfW1f6vVGJU7jkbQSETS4VjIt0SioIWRS6HD1NwRK+44Hrvxne
VUOX5r0xKXeE4zqCDtkbgokooJEnNJW6l6Dk1lgb4Badcmx4hQs1FGG1DpV/ErY/xiH1eH07ByzR
AjK023bLa7ETKcNMbbtCZqc8/EeaOieuKM6yDLbNoFCuYrz9B+5PDMAsR31hxE0PxU/Q/4kIxGja
E1AD3dJXH1z9ZuHnqVolIN3YfKbwb6OaYKS3tEhErGCcnv+bdxFSrCv36CfdM2AKddOLDG7Ck6hr
ZbRO4IQOyB65xvTJrARj+ZQBfPTe9RjFIuDpuYotoyb/blxk4DWRAjLtmesg3aSRCCpySMa6WtPL
2bGiDsjv7uWRmurmZIqYzxMYBBQU4Q4HzV4PhEkXkJuYzu3YMJl2qVbgH6Qx6XaZAc4mxf+HaC9L
F9djdrHuiHNkSIpsl23LTIV4EXWfkoPyKB1bEi8TpdTuDpdC5kKrr5YkE5clL25yqfHDZ6sUWNgz
PPFxS77C4jKxOnoPoq+H8YqyiP7HcGzLfmsueMdSaIAD12Yp2KsfthSB6/tUpqUa+cRqh4otkc1g
eRZjtVbYZZTYQN7NAWlrXIpxeDa1nbN4hhTxvkyswncFfC49vNe43h3xlAzlbzBYaV9Bx44BHvxL
wUUWCd5VOk0l63tpIVp3Rcj12qvnXhaBOsVmuWnfKWmN3K/QkqUkD8pCO0tBWZDuOfIQJE0srFlt
Lo8LRNehVEJcoeVKx9SdW5FyS16f2EHeP+AzGjnr8gi/Zl0WbeM8MdMjFXN6NJd2yl7LM4h16u8p
Y/u1Kte76vrufzfBaexW0F36eT3JBdS9ZKhKps3HkdYTNbz7YlcRd4bvbmjHzK9kjyRPlPRGhLT7
U/Vyc9Av+Gpu8aXzdSKh05UXFNQ5EhzazOj08fp34WdaooSRC1dNq5U1V5GnxTU6UMDVBDGgYCKV
f2o9OPbzkX/PblsSVLLF0pMp05/1EICQVODwR+LA2GiS2uaQl0BBkRz27kDCMa0k1nSynynNX8gN
c6990poUvEWv591WiyD/qscE/UM32A1FUX66z957b+ujyS56L/AKllfuYK59P9j+7tDmr10bdn3q
8XOqIuNfAIoxMglAaMiEoUCZWrTC0dN1mEukz27lqVGTRgHbyKdnrXAl0PXwfKqGwTK8hps6Ohzh
ls3dOpdtNfZFyeuc3uau1v+qY8K7kxUfBcPFZdyPQptK5ix0bA++MDqcGRv/0wzdkjENYG3Ez8lP
/sGIqy3Z+6mg/QEknoDIQvk6MHJcvpRI3T5odOMEAjw3Juz7mbdi+6DykOIVjuDoNo00kWHwxkIl
c0g5qlHxQ4nY2a38+1G3iN8U/mps69Q3/MrLURGsyBI1lGiknODAM7lpVj2nWp6oYTcsEXAaApio
ZdEtfTGc6isAR+0IjwffwrgOQQGZg+qziZ2pJOaVNaO2Mlk3xoWJdo9G9nzfkaWjQV7LsgP41fwv
1qnKWoPhrQUBDXsYbWXG1XILnGDGRjqA6o2HJukFwVZoI/t7RKqq53q1lbwfT0oOPVwV6zn539Cl
7CQiHWYadfiQ10u/e4BrtnQBKxmf1VQhodUuQX0EA7qwRpKAFmPzm0iBZ22GblRvurCZGk7vNdHy
UeaWG7ys1IB3N71vpRwgjLzAEm59iPk+2xPNnJz+Xrv+e+Ee4Vik28WiOq4mR4DEBWRZdvGNxo18
mqX3s+zRZCpxEiYXk/KcN/qnmSw0Qbfrv8AuMjOp+0xmx/VrrZhHpUDgBfxp2y8cCuWerA8Uo4kf
eu1rYxfgXzVhpRhOaUrUmrNBR2zUZg8gVAGvafgDYUXn45LStZ3r9IdtF4fzocmqYYiXixEZO7DC
aa74CBStpSG57PeIPCbV5byyGzpWhzBojkZBKDaSf5zd7xhpmbUkgBNv9CW9qhwZoy9wXrADDudY
CCT8UfnDiJ20bJ1M9xcW/MdugnLtSUwGK8NwDgqmUJthS7y8jfK8cMnmzDkeiz6pso6Wu7rq/i4c
m7seJxwFnZWQeq0Box0jIHOggG6F1bRZJ03Bdat3j4IfRIaA9xChV+EabCa3hPRWrT1WpAzzEtWr
lLFkF2FT9ZlNWhHcF5GfA7afpXMN6Rm9MdznTojrAmwvtJQnJZwzZqXHW42GA8eLw7b0dpAcm2Oy
NHkdEPJFVMouGoYayZFtX0IVkNM56DW3jKGsIXn32rFVCQH4vcIenpvgJC9xJY2PPv3irfln3D2w
He3xBNixvFZ3NxVc5pySbPo/O2mrZcyAKkKd0aMOh1EDT9Jq8E30GFuaGYAW79Lyz50LFjYvNMKz
FXRIpph3Z9bFBd1u7jBDyVJAR7GvJ8Bw65RwiDnWRaN66/bmQmQDFz0KcB/bursz2sdlDsoSiRj1
DZqmc+rEMW2ZNHc4/gFs9LL2Eu6ejjvQxV+2HGGM5yghL+qYlrQqD8dA0BWgtY2vTt6R7F0Ml7e7
CXxf59eI6G/QY9de7BWkz3HE6GgG+tG8s2aOOTjmHZ8GxCAe9NlMnrNkAlpkfBgeQJT/SrkJYLmF
FELoovtIqlZ8ltflhEfkgycv0LT78xP44otWwWIT7ShI9EWPgis8ju9fewYE8TPcCw7I8KBhCX/N
IBaNn4XUkduYAAI1E05El13iZ6L97ErW0QVcc05c6EFaFtYif/knItxnTsnY7aHOW2i/qBjtPk0p
orurPdDPXG3Wcd4nqT1oO1nXfPyWDtqCaANDikCR4Jsy0gbGA4bcqdjnL/DYrUaDwBMMC7WPFakU
m8skuxdDBCkNw0cNQniS+xvopWSOSuzIcai8Qq1ug66Rax31VxmcB7/8MrpRgravoW9F8R0lrwta
RqPXYme9jh1o83mWDdGeZDdVNca04HDfVzwira/SdiWWdEWTlFFl/nOsJ1K9nqNsn4fspvxmhCeJ
gu1jR1/UV7hYUhr/RIhIvLGXitZZau1914VVhXFDqX5K6IuHFlvXkUJgWgtY6/Bujv25aC27hXJH
rRwyqr3VMpWfFXrlhRWe8CIzruX0/ykDEHI/COAHfCiYVEdNa/gs5zCd/A4ABVfV0VM6vj1x5gLk
oQBWy9ST/zXqaQ/ui8dkB5CGXDVVZOwV7dQEJ5avfHzNiKqMwd6/0+7h8rBjOy/x6Y4wZlEKDgkz
zt+WHymdju//H/nPVExfRbXqEDSsZfTe7uBsb8jFkNXDYeNhQSWHTT6olaeIun6xVlFqSKXbbQfx
DljsRkCwXnPd8ZXkIj73ffVshB62g2KdD4ObquiShkHGuqV9KFAQ3ylzsLwz+J4Fkaaxlz1G76zr
52E6v1XzeG1qW9pGVEkOt5NulRfX0pBI9K3eWY3RwZ+R+nyR8IumoJ9Kvi+x/4RKYJjWaV4Hq0BQ
O/IFwBWfhou59ibz02Uup95KAjLGPILaCE6Tb6OGnK8ny+Y6dKMPQJxVdJiqdDnlqucgXfuqtG76
rFIEDfTGhh+GW2s0gnseAiUTgB/imT7HJw1oBNqD/YVipJzBVwv09p/70G2pKHnlWpCMuC2qbaOU
JfO8mhizADc6NUcVY5kuaLkn0wb+fo0VNNbBYMwfsKzcPufdt8SmoV3JtYuBQjODudaj5vPhnxaI
bmYPN05wHDZP7KK0CWYYsiycYbfMYcdOSpUJi7UVSf5eVOdOQcI0AxpCOs5fl4dAKsbiv4/W4MZG
jaT0ZpjSuTaRge0xM4LquBpgISppUe6F4K8s///NhWd0iwjHCz6LwPr26REi2MidOow75GXITyba
ihe9dgePGbPRIunuzJ7k2QyM5kqDPfMwauGwrKxSjCqj+q6lMntTeZfFJDoWPoiGIb4OsA8MUI45
LxTgwPwISzcAXPB3DsbaMN3dJrAoW3nOiptXidIy1/Ubr4z3LD+/5jS2ZV2tvrAA8kCgrxgxXGtq
V0uAJzEanAIznPzfshNvXhT/WIiuEqyQmtiLv6runTkru6V3amo5vXsC7Frrvu6wpuEFBVqOSmwY
aAikCm7H0O6WEmtYCyLSJzf/5Zei1LdAGZBIQ/3NsnPUAuujU2yBOi+WECdBrSPfXyyrGa1QZ42A
DgRrQR+NEY4UHsoCr9DPHP8JCR0U6jbGk6vo1xNzPXUo5BXHWd8Tl/63eqJxy89KEyaOx/eiAeP5
NWpGs4QydDqLYRAy3ALFFtb2mxZBtOPQWRCWOcWlid9TNQDhuyKnzvLYLS8kjfNnQkv/oUCzjUgR
l/T5vQAx2Xoawr8FCbmfXqTu8L3pmZr23wnhzXE35ujvDBIP+5SGaDzoRSLoI+elZhf21++E2ALB
yCns0/6n32uUfhddgQX5CS2hgPjRrrhXbb6UsuMksZPRKRspT/dKIEz2wckzwjUo0k3gsFd4ym0y
sh/0/gqPc8L9LmIcm9js2/8urg3TFwnhNCNkohUC7g17SIpcL6PnF6dTGND3VU2iSF1VaeQKeABK
Isy9L3YcTNDMGKIf+RWZFuQDBRBQqLLpDFEd4ZFs7/lXRxGuYvpvM7yV1QloWnm9KUEtq9pNQLta
whD5iup5aDQxvKTIqRrE/sy2s6EXzcQknPKYWv4bqCWfu9idW40zPucluOxfp24IDad5hgVzYgDw
Usxlh1Qn+CsKEEhTTMAGd3cMX0JqoUjKUwmJd/s8lN+iqtGyvte3tqCjHn/TAxOAM2KOcP3w6T+4
FjiOQxgk/F76L5uYaL/tglIiRW6Kf0K2FL1T5hYxnPOM4YuKExAAs4hvAvbeF1kOiLJ1f5HpCfdq
v88bghcAe3Yw487/6Rdx1sxKus6yXduTTACrc7M64AIFnzlyii2AqzBpQQKoK9Rh7QMRsuEYcgtn
NxWS3CLCMl/EbQ3fMiMbF3Wy/oZLq2l9dCIQDwreKuvPK9QFfwIX8QHE3mJx5gzVDfOkrLJDJng/
sEQxHd89udwdTaLfRpWxmvTPOr47khsvrmi2IeslO1f6al9afszUWNi/qmzkgnY9+FqWWmbd/lAx
HZRcc5xdg8tS9dDt6MHENBO2k0pZzafoFaWgBK7NMfdmmibI+v0nrummi1MLFYQS/sso7cmbgnEZ
pF5lnRNMHGAZ06/XjwypCF2C0xfvQi2c4fJL+tyG9A0txujO8zZK+SpeO5koSS5vcjuQvPx410OG
j66YZj3q96cLR5/cBE3vbfbf7ziT/vGcEyZpQjQGDMewKwsTTgdPvzVipReoDeC7Cc4hwlCRGTN9
khHSNzjM0cardrMEHEqfpyhgUqDqreFLV592Wpxs9Rhy4OFhW+LBmEpMtXumblBNjXqqxFN4PzB4
+TXo/wL83ijJWWUhSR5t3tfUo6QanSPnJpBrd5loWYkFSNQYnhx2LhpePv+a9XKfENKrdI6c9CTW
vdKrd6WGNHtQ1WCEjEEpc7tjh8qg5An8edHPXfmV5aE5LH7qqk0oukx2U7IUpeOM0TOGseAiUC9S
HNil+s1j9cBOKqlP8eMoQfA1sBQVn5rrWHsQ4GJNSmLBF9sxQ8k1YZkQA9zKML7qvofs0nZTef50
OOdXUnnB/N05FgM6iVAarAZVQpQO5yH4Mdj56lfHUVe6N9JTpwzyTeMOmjjrDtKSE6pkL8mziLKG
K9/EVanyZO5TvymzrP3i7GISQuKx1NJdoLuvNtFP3r6ECg64CgUIrz41mOsvT7I39wsS9nBj/T6V
msqhLGf1rJKJlRXVpvU+d1Srvf+uaHQX/vSN6nS0ySzoA0niEHYoUrOZMPB5MfLSAjxUAe06rPfx
V7Ot5W+Zn5P1j1Wm14o6T28UkeVBnSv1b+4fSGSWcV/MFXt/o34z1Qf5Mk6bQyujxdB+9PefQ4sP
qNbHdRmwDFjKvOUW7NcJF0ai/58wk4opYNkvxJLDXFnLX+DUWhqn9sNTDKi82J1s2C/8DoDm1CUw
78cdrLpt+TfzAPwkOA8eh8USanGRs8/5qgI7hXFuBBt65xGnAMPUGOIX5nYvQvFlEp7NIdjDvjqu
HBDUemWH2iM8MTgzBE11a/QNNi4OoSwSYrx5p+nkP6HOmhWngLrtIPU7gu93T6sh4w30Et//uUgv
AMadY/7in04RhXwsNQl6BNsEgdJYb/vXRjpv+5/EduKFlWjx/K+EnnIE+rWFFusKxvH4ruOJKz6F
CW9BmGhh0PUcJL3lwKGUj1zbrOTpGVZuArsFZotD63oDC0ieYzCeoKns1mLOgKiCtvRZIoJJ8mk4
/z75Z4sFFJ2L5X2z254VOnP8cUg25OOyEAptkRz3hXalafyPbxOqc4qnsofUJSAqaoD3FCdRE3U4
keJl/7QGkPJsp01/axh6fks8VdgbIYf8mld24MLYomUoUNsatDyCLImbqcEW5+NgbwigDfVP9CwC
VcG68cuFL1i2ggn15i9hoptY9TfZR9L+6fAsO2IG/KONFofU8itnD0Zt+qIuWEXwBqgkT3pHp+EI
20QXdT5aKsG8pO/B7CgT+PVNZVtO1YrOk41DU2jggukreHMoOEAT+gu/FyKpMXuT6gi9r8KYx7IE
xbqD6tqG+6ahM/SKfzrZpGQxPwonOrONxG0u6EaxG6Ogk/6XBz4caEtfK0E43xq27nNA9mhHiFVG
A35JQAYRYcYWugHW4QFJKm2pvvCJ19mqfBNHClA4ND4i7EZOl6HUrz/j16ZdzGFtZ6ZAdSc3qD1S
MQW2wv0OgERGRx6gQPusRFH+/X+LOPjHJo4PdemRSz3bPijquvunvjcwGlz/cEz9z4diSlTpb4c3
8ajvxAoElj+zVzmPrIB1oy9L3m2BCOtLuETJhJ2pWKiG++sMen/5kjq891TP5YeGypiIYoREWCfs
HSJLE38F/S5LNBkAOrFCaHU2aM7omowPgOL+f9k2RWAl3LaNTWqH3eJQNK66c6DwpItJbO60ed2H
xz+XUfJao9ApX272KKOA3tqM9xmYgMfC83hyMvlpLV+a8SEmrO6IegQZ+RxP0Qx9Yxz69XHtEmzA
yVHDFhsc+ZgND3Nhx0SZVGLHGGdxnJ/9ebiCqapMMm5HgNm26+1ubqdjJ/9sYKBFtHFHrFVcANU9
Ms/IPYgHmfXMy7Mwr2LLNXX+GIRBGF2zapg2+rdDK1mKfuzjcxcD0u+jjbtO17aFTVnQFl40Kimb
WpwTLfproWZmfBs/0d/oBZyOgfy9uLY2bLSsfTvESRzQUpW46Yt8f6PLpyujEdkBmmOr2uv2UXlR
o//EbS8EqXH48wfXB8ZQ4STYlKSCLkugDvEwKgy2MqPxZ6nUIBfhLwa3MfTo7I5Bt9rUddiXXR5n
PGAtkhRhU6SMR8bFqKHrD7IPi614yT+fUwXIzlgjch/UQ1uWOKMFmAFTXDKYt2ly/moPXJ7bq3Gk
0v8D1RhHEECu2xIJBtgcqHXJt2TntwFclY8EpoHQSEktEtY4GC6JdiAixoKHMJ1ZvEII3SRQwbwf
Spei4x2rKHwOPxhFy2ZireHABuBhZmk60r+GxOh7ffuHlUWA8JwcjEh6cW5lezuEnkHnHjyzJ6Fz
kBxlQFdro76mG3kDPNVbzCJR2PLuS/KsNEsWKsp5WVlcE9NPvH/LSkjUzaONMo+tW8UnXXhWQ1gU
wb2ah3suqd7Tr5YiGwsZP7IVRYzNzgr3VJPxN3GWWvklFoyveJlxzUxzTAAGZQwfkq7z/Sjo8u5c
QEIyzUFEpJBJIJ/H7I5AMoYRoC0rAax+j4qywkCauD1WFRKQMSkwvg3o9Dy/GUB+IaJ98K7XnS/w
1qqwuu2cYKL7yL22c/YQRXz19XdedMGtQVV86/+Bb+sTzzMk3bro9m42ahkJO8l0/Q9VtCEMVUok
hQj78rLNkXoD4KQkJG0TvBzaaQmiPYLfRZjw81tfhesr2GLmfSyAcliHm6WXS+AlXEVGsEzOnUgk
LW04B6gGVbRza1UpJTxUtNOqZr4eslefXU9DDuyjOL1tiE7o4iDAocvU3sbuT23eEuaMKCsAnvTF
HlXBYC7qEYjyFygKU15P5SdqvIOqAIhITm4O8WHgYWbLpeooTQW8HleKePRPlm3tkgHQJkOWp1CR
tJVGeVzD2nImFyiQ/j/ThnhJoa4UKNyz/UwcjvpauCc1gWKj+uK6zMINv4IiqZxUSvESB7Efok8J
DAJ0J4oBdQanGKKuvG1YdTgc5b4FEwm4O7bFjGzYoXyW3abJIfQcBuIYunbFUnZzQcGBQObWMBvs
JZ5oEnovPPoMaGO9VvMxRuPlpCr/3JRCLL8lFKQkWGq8+GC5N/BH/61kTZp84WT2DikGqfsDYz5I
FgeHY7hmVsWptntl5eA5uuklJbc8jAIAEDtTfI+wpPCKNtgXVxja3hjLyJxEb/PKHnVEW5zgSaD/
FkaArIXK19lO/YWI9hNI6KbcVmhx6nRbPn5+5dGu75xSTyn2fmuWAod6WgDjOqzUllhNiTSBS2Fn
GXaMu+QjEbI8O+2FeeNRaVRs8FLPmxl+G/y3MFVl4Ht2u1u389R4JAk5GkAQ9/+bnMVj7ODnxOIM
pqeRbwhIHuJjYix8e6HaYYFPzoeu8XTb0+R8oW+tImJqzz13frj0QZ8V+cKG9+jT2Pc0F/SWLThZ
Ulp0dPIPRcE6BkF2ApZaAkTFK1NgmPLazxR8er1qMRTQuoph9Edwx8ZD0ALPpxtohkO2s1lg4gw4
UfwtDiB+41Yk5RJ3gVHP+ymZm8u3kgOyN4tmFwV7e6OGBz0M2/EKQ5ZDdc8Ms8D7Qxmg9MuRaBV6
ysbx3c/W840hMF4ChoSqdIR02YKgZPMOY0+EnnzrU4Wcke2oze320FpHo8ZFQIYhTxm1QhelwqYV
4Zs6gONc7CYa5IypaRSrursQSo5sa6FHKt02Tmdo6d5ScFPUK2DS+/MZ1TOqyKPX6fI6lS753d0Y
gL4lCWS4QCX6hoiVfW5If3n5x56Jsp8DQDeOV550queCdRHHTV7ug+KXh4dLnXZM+8K5PkxWGUMw
q6D6dOocXpOumXRvjPIqNNBo8ptBy/lA2V7ir7rQV5PEAOW+O7vouKAPU3HbPQAsIZhhcuYuMb5S
0/io9GwVoghHxvPZIlOlbJxbmV8nWanbzi8UX3sWy8cHKuAKHloakhA+WRthVkJXM3jreBHxyaR+
i+P54zKCpGBP1ci7xjdxENYCVZ5FRau0xffteZ5IPEG7N3A+/ZkYwEWLDVHL3mAA4vpGZd2p7Lva
Pb1CozKbkmikVI8URuWzvtVvGhiCKJioN1RC8IsCI6tuG0eYKoYNP6g6VvStyq9peZBUrIIdLqyo
6RyNJh5GaKI/8vCJ2f7naZwohmi+2O/NiYAtto1Q0rEcEowtwF7js66GPwMte6XmLm2jl95I+z1h
PsUWhpghkTF+yiSE/jyaPcZne82Nb1wUhrixq9Wx+vOTf6QJ+SW8orYUiTVqFBBbs7izNjS+abXZ
d9lcXd1i9oc5MBBsH/l4tIsSf6f+kgqVtZMME+eICbecxsw2KT95TTZa42Z0dYVKob2tytpaz5OX
uh1Vnca+TyYv17moptdlKhtwYcKsWoXVGL8OIfE/C6EKygw5VwaXszXGJXdS3UEkKgH9zDmNxC3j
KBW4SIH5G66AfUgGuEJ0pNR4cjyJZbNePGn870lnXnuJqwfm6Lhag8VY70qAjlzNoeaA2zH+5iJx
k53XTI+Z5zOyhc3JEMKiWcY1EJ5+BxsZB0Xi77cZOwkkdjxznoExLgFB0suA5f4kz7aKFpQRQ7GL
fLq1M7dYVLBkiTV2L4VbYFqWCq4ELdQcSIyhvCGnidIhUrcP1hvmSl6nYXs89jw4z1fmhz7akJLC
K8vgKhmm69zsjj6aaQOlgitk/zHkpkmbafiY5keBRZWxQj8OFYV4CmHLdMKaV8Md2EmG0KaE9X00
hEA0e09ToNoCEs5kURFUvWEeVcWUAPa33mSyKMRGFkHXaAjD06KCzaqqAbrxOWOk7LhIQezpraxb
uDBIwKCzzeVijNu6JU4c0RDfv/la6hC+r8r1EfSudRxkgERlFCBwh20J4rAFHbY3K/oeao7mm2ju
IfSJkCRdPhMXCFR3RYXXqojCcYXxBuOoyTZdrn8ISdrbJnNmfG1Er8lEQXEAWNs4jz4mQPYNUEYH
JWuoAKzHDUJFdtgMW/C/uGVyT9Dc4Z0FgxgSJK8x+wjMkuP6sT6+WRnYmhLm38zEdmqGffzXf9N3
mpNselL/sWYKchApKdECbYdgmBf9iraGqptme55wIN+F3tW2/higfBQ0TsdmC25tQsnU9Cf9FKNZ
QtzcIp+gUhtuu9urYYn9CfHRhyT7LJS9MiFnApAuTWKkastOSSgD6FaN2bMg1ooUIEULB9DywQRU
0d9ILV8lGhcGfivOVWZY4WTngNdkxicvePBU4X/F1DCD8lg7e/g5aLw2yD/xH5/bWLzpNTj8ctRc
0E+tqW5Lj82PnUyd4kSONPzYDH6WdJubjk5uZlWFlmH0ov5zK0dhOASsmViNrejXRtL7sc2RJ1xb
x9go4K0TizqJuyr3WVPAW79nKK3CqQ61ON32DBolQ9I/rZCnh1MtavqV3k84nzffatftbKiFlqBE
6ymygvcwPyEn0vrgYgMcrUoyHuu2ViPM/QnQaSqQbTUSJuEq1ZCiFZsXqXwINCq6lQfe6ractV/M
sBo9HkR9+hJbsJAzes4nOtF2IjhjX7qRLdwbobIG0oFyBtfXjjIOFh0swyIb/FM0E/Z1nyrPcmZQ
lSkiMTu6X9aSNFJzUVkMsRuN2sv+9CAim1kRh5M2KaEPhB5ZsNoTyloWHOVAxtqx3h1WgMDzVZQK
05rXDpZI3pVV7wNp2/RBY4CzW4m4Qg2tNTp4DQDSrf6mENyYa1el6F8uodgrHw56wTtHMOQ3bGp1
i8oCueUWkTIERrtwRS2ESsXlYTp+umIoo8CnaLXv6ixlhXgoUymqwfiswL407PgDjNCnn22WBXuU
QLtpf8zAh+1fXvQT1dGBSZ6QbCxcRmLWFSrVYMRl8hzzfh906XkLtKCjZrFDV2ibu6y1tjtPLpMK
zDS8bEplWnVp+lWlNkqgKuvM7gnJuHX5JOXX24p8FAtaCbw0jAlU6+gK/y3i5kC2CAc6k8cKIBHD
GVHC6U2Uz16FvZ0X3aLVWMbHRgYYt79yCGj84tDGvEzyA/LK08KSDkGIvrGcW484ULlx3xol7VWM
Fq+f6GVjq47eI9DP0zuMB95SDHaY777dH7HIzCb6kZKTIOrTYgL6nirXS+omWYZeUeqYbHTm3ruj
VRswbds6a6e2ai8f05/71u63eEWsqVSAfj22xmHWEBBSEjqGDio3tLyH7p2Pp7rJi2qJUzo9qkps
YBKze6rviVUehgTuwH4NNTNmcKpAVDrq9eTrX2PKQrIfXOSJSBmRUQNUzGZyjkQ53Lm/MX94GdzI
bv+teL2a17yAax6p/4qICdnMDJiFl3KeRqCIaSan20e1W0P1KQFPYsQt5lUB6BR9KskSBKUFauGY
O7KGabbM+GIkKM+Qfw4flfg70hGmwBvTJfTPDdx6uhap6h0YWPi7dxmbSfdVoZpVX08PIV6ZT+F4
tQWB6JEajfeIX3DA99BiDhWo3eBeDkNHSjGChhA7ReFgTYYPKlisNVl+vswxvik30tsqfHQjjVOw
eDZmQPIEGCTmFLcb3oxanLtiWdcWk5MAKi/zQ2IPW3jFz50bYLJatGAi03oQ4YJ8m1zqWcTwZMGQ
X+rJbtlUUXbSaXU3gx5Ofhk75em07gbDlru7hQrJQnb1f6jMEGxeGneVwprSkFmuFL7tWlJIMY22
Cp8JKEHxDIBondo7fewD7KwqjP0xxniQhQTXop9HbUtyla6zwvLv+rl5MvRP1CwmMuqoErr2tl7A
x4t0ZBz+Y3lEo7aT1j63H83T2gqDJzdm0/fGykwbHYNhigNs+je6VduixhtZGrzMqf960OJaYtf5
RD5cPCrOhnXBodCHu9iK4Bwm0ZyKX2vtmWsu7uyZZMFhUCBbGsDJ7jfOxH82fmOl7TVBcw/0oQHU
MF8d24bbrhHvT0FqxFIsdTF/EmcUrEIKdJZp8EcToQAZsbrz57lBJVdEsWZmCZmWi7pfHtcTtVNE
n/iCFDa/dV7zR0GHmeb0NRE5JoLRZBYZ6U00bCoCrV5QlA7qDrea8ws2ob3wGz4fci3VQQp4w0Cs
1JJ9EbROwqRH/s78zQnZNaklautcCC4xbEepPvAdqgfCQ2AjDJLv/6pYWE35DTNx18IQuNn9azDR
/3y4w/3LJ6cZr7mvR1OiciWkhq6TxlMeWLd9QMiGnh3gXT2oS1JC/UIFC4WHbDcVbBDBA9pFZnK4
3NrrrZWmwiAokcmJg/5ou6lg6fXo/f6BHoPCmy2+EEjQRbi6guzPuo3VQx9FdzoFhFV8dM/6Ow3p
Ebz5uNav7Lfaj9REfCf0xzpLZMNCcmfOAEbbDMPp0xodTpSFCqf+t0CpNtXv04li48TM7bIrXqkf
thJNPJDBWm4Lq2SjhE2+VU/eOzmxdgnG1HM46m8imKX37104XZCXIP51tChYOQy/0WynU5GFnDJs
oihdF+vGUvEbauuAuabilt+wbPXZNjpoEZbXygoZIV3cGnlsYfp2UFNcp48RU2xoEN/e8rlKxE0k
lYl8StryW7BkezQ5Uy+iQzF5+b1+qhiU2R+AI3e89t7+TU2Fh9IUWIizErgwBvf2XSv4WaHW0FxL
efEGXrs0htKYN2Qi5/K5cPdrYpupYNGOZWdhef5NQYSfTgXUZq8jnEiaSsSfZx/zqhjXhSPcUFGE
nPnJYblQ9O2uma+FbDKMrOj4BnN67sFKy+og80LUufzkd/U7uFzJcD0UtAtrcgaTUfgunZnzKdpS
XeMKhG0I22aigP298y8QM6sB+MjJvbXulyjWDddtMqrPaMLQubekd+mm/C/xeKbf9FUdv79G/GGw
nY0DDRf/D0PuVv1Bl9Xs1yxDfxywv9jmlolK1ljF/3xMRZKriltfahDcjh/NF86fT2+NZfHfGXEy
v0kfCpaXbjKJW7lY1tNreb0q51/0a88bI4oKwSI+hyMDkyz8f94vo/AmLke3ayyDe2aLKsAUVtu8
fNMgcsmAFjBL737SgiH79QCUouOf6O1ko9cQg7S2NvOsFi68sO+kTLK4hXbZmrvcw1eb1DBr+Urf
fP5iiBFqYpBIwgER85VPi6Nx9h9/UrsbDrkJPQ+FN7FqnjmICNws5tbenU7H8kwTfsDX6UReN1Bw
5tQ+Sc7UjSQhhuiTqc2xdKb3n7oSd5Pt8EONjYpr0becXDF3iLxDYwdM+4/zYkLqbsqNNZ6JWYFK
rhF68eMifXhaerhWZJO2WY12TKeuTG4v6FV2DCoiGJ/BZJk///j7B4vlYow58/ELOs3lvHM40r+y
JJd0HyJXOlLF2mEbYKNfsqa6aV6awLgH7645v7kly6Ujc/L4WM8h16isa9513o3p+vEobB5C9Q7X
bOFb0LhBKIZmdaCdLqA6jyJzlI8V9ZE0unmTcM1usPvghRjvgBw578upP+d8XSADio8XYqtohioO
EoenzF25T32US9JKEhtR1m6iLCcV2+pD67S1gzDMosXsVK6VYwVLTk3vNkKpkDZATTvQ28LXK06X
0A0sutUxD6fN2hop6okNVD8dBibNETVD2j4U9XDrZ/8SDYQvVxT39GHVFHwzBc+y++Vrrn9+fJmS
rEnA9apXvkCZVi4wjBaPmbsmVhkIovBEe7ZVMCsu8aUy4NDtXe6bBKnk0q+oXR6F7DwJrG0W90Xw
5fSUI5e+lx7Xm6+nURV7qC2V569I8voXYhYpWfxrw6cvSVU3r830m4CkBYkSlokhf4ppb/UlCqPL
kaMhE+1g7/uGXmkNXHibTOP+Bpky80C9i60IlIitAvTIgVtZn5hpqnCASPISAegXT6jQQHBZI8hO
mcCRzj6kOO02vA2YoeivcqQmvl5FRJtzjcp+PZZ6JiaWotbjgnLwu1WFssMgkIQE8WL/iMHtzVJm
J2yYtef2MhK1IxCUMYR2p+LyWmyssN0+FX3uYimxSx/0RK69L1gCZmhG2rQg+qsJ03oWhSTYHg0e
IB2O0EcA29AqaLrvo1VotBRPTVxIjy5rtNN1ue+/bX98TpWEeXWE+MpXSxYbRn+ivmM/h4OWfrAe
qnFnXYNwLJzBymRh2dVpppnhASV4Njptt9E3lUjEW8gytwp4ceBKEzGhlz7muzGDOjn00kIzWOWS
jBdgMx3RmkvMAZ1y1oyaAj0zJ3nvurVv71HnZL6nKrBG2N3m84K0XMJmetg9TdyDIStYf/+I+QCw
r2JrrOqBV4Nuzy6lSFzsWFNl6h/8+9BOmV1AuwROl93+Rq5Y0pBks20dMU/seP18ZgGGeVUIakhO
h9Q4PFBn/ZNTh9a0cl72yPQ8ru9tone3TB5rrXuBRI6f8jdG/kZVF7lneX8WrmP/OXp9GDdtIPWr
/o3zTJYMCzfweAgFv5m0VjmnGnbpaJekcawgWwh2xLjPLrBpeP5oyTfDd+L1r+KY53S1GbFziylO
j4oQpN+X/cerfJwh7BxrlcH4TblmgpVB1F2+0B2EHCELV0zIcQ4wMJJz5vo3JfP8oyZD9nBrlbgf
04TY9JQ9STED4S6G94WZ0UANPflovODBxCZssetc8SeIMPE3Ow4CWg1sWlN4KiL/aJ3UwDtR9zs9
SIbhMJORAKd5QsPgVvI+wQWHHCf2QhuU8c5KibSgXNKP25zGo+M3nQjgPj8IdHBawE8/HUUtwKbk
ef6MzbTBNhx6JzTUvUdYsEgp22tD8W5szJR55vdbAPc4/v+BmpCkFXm8ep3oykxpssZHoKIidocc
tT0rB9xrY8WzR8S0ArmecX9FikCL52WrsEWti1a0x71HIHdqIJwXQTEgDtp8+B0GQVlNcdxhbNLH
yxiv2iU2L6/Jgd12qnt+epzvHGR30j9/c/8bLJ5q7Ht6Pqn6mcUTrZCrF7lgEoQmSBnjAcqrhyfz
kOSysmP9w9CTP861t/Qbtu2Ugi4CvrfHlnbEv+/SfHNwlIbJWPpVs38TJRypramgkFqnmYnFh5mC
UIiFRd7okc+QQCvf5DC/+8VtHThsvGqyX+ehwL77WqW9GX7GGA2691ABzNz3XQ554Ohj06eCxV/r
LLOxbHVvJm260QIH87gjBapayofjQADfFw4kQ7FWv9AVycm7le323k9DGS+slZZeqtgENblFytp5
fJZ3Fr24QNDWvo0lfaIkCamydIqgxCUta4/Bo2250CEZ4il0QmQFx1E1oFXeQKS5+OhMU7eDQS2+
BZXUph4TSfshCOaqEmx9C6mJNOhXJkTLQzKq+S0JV5S0Ux80/yd+0uEDSDQ+pdtkxaGxif9E34wo
fpkfBCmbaTlFvY7mIA4q6Q8sOc01LyhL3EdpG3YLfSMJVtxrAnlj87SMwTrD6oMOWPyn2MVmTPUK
iHIp904oHsVW7KUvucIfyRgfOvmBYS2ewieW3oUzIPnDyleIBLU/eksSSo/U7ikxBJTHFueCBeOy
+CDBkPPZPZtAKa32WevCqB3mflSwHzk0RVsjxheidkxrT6LlXDSxPZKjYpGZbMl2sHls325n/sIw
n/Dw50BCNzN7lFoZStSgORtudfkFlw5ZRNbcHF3/P76+Xp8wMfcV3LPWlZmTaSPMTR66awlhiryg
3dTYGG9uk+VTBplDKxvjbCCAQADLTSntuKUErbhROWbi5jips5+47BeUBIjB5YiihY5QBEhAVdrt
hbbo4Tr3jmgwkNiMcNTGDLkfR3hLUzTGRAATpUZH+2zkFlyJhJqHZmVXzvpIL6A/YBcOGPzeGOjK
KTjZnF6OvSLbskXmGkX2C64uriIR2O2iqgwhTDZcSD0AUcEAUmS+7INpDMfYNpWyBOojXIllKhZc
EUFePg9C5/ZuS6J2pV9m7y1VmcQmxvY4tFKgaNvoZCbCNSwV19d78+xo8WtVLwpG9/2b6O4hHjR1
8vrm1Pj/TILXsMKhIN2tKm0vwmmVM6o7WZ4Ngo0eJb3yQVnVAufnxhKNes2wlMmyJHl0nUb9BojI
eE71hs6RRKPrgtW0vT42ta3oHLmHYt/Kwssi8j/aVbZSyDjVTwXDl2ZNFva3VcopRNfbcSdREFJM
QYzTwA3ZXDdg6ez9A55ZgENEuCUHBH8YkCXQt/UnkEfnEogBCsq6yDsryBIjT0bLTTvrfo5f3cEx
/uD39b9OwCoHmDmzflrQOFt0thx2LABJQxBtnMOIIA6+LkeKutWwwIC5UQ32Wf3AdayI1rzHPWIf
/WJPYu2GCHhYIeCj9smblzcXCfbxfjUC1mbKY2hjgp0kmvyw0GPt3We9S6PdZ1rfLxSXmtod8/CK
drzPJWg6s4ExyghmGl44E0achplT6gjkGISBtItwBpeYuFa8oVSi/N8cC59YLiciblG4kd6wryFc
DUDx1Aaga7aHB2+bWpub2Ih3eJ7IPY034+Ehha6O0DQ8SiuF/RNUaRK1l8wWo0J7K+MF08pUqYFS
0FM2gSd4Eu30EJQtm6DG/gMdXDKM+2M3hBTBV2BN7d8pdsTTttX3fWvXFASPjZzcM/ehBM8mEx3x
iSXCbEGWxUXAWeZkHov4d91Tc+f71BwcKXL6aY80FKtXyG+Z7tfy5I+WXcNrLsK4SO69wJcyT+Uz
NNk2XOmDrfqo4SBhzswzPB4r2FxCQUPUFgoCPhSaHfQ0gzmCjia/9Ck56KCCAwmjGBoP0C90wfXa
noHvtsMpNQ+Utf1ydnxGEWM8OOF47kYI9hvkzv+ESgUNSyTxuGIw+coghaFaeTspkFUmBrzfphYR
90edyMTXldlcUaWkhuYSvXLYmC/8uyewEYLMtiNtvyAXTGSm+/ywtBBuDLnXVr2eDF8G0exWhIJl
/NuzeUpoQOx3+1Eis3onYwnVlq3YDYo8dUZhs6PQhEeR55/kA8KlqeHGDo5GLJCunuj7EqSu96Ut
BFQ1cgdoBDMs9xU2tgk98eXm5sYdK1ggH+VBq/N3YmhmXFVj9MVjY700onrznawPr36E96wdkmXD
tCCT/9Ve2FgGbiNTjxQid1f6/gNENdMR7RuGW6pwwKVam3jcfKLPXjs/+q+YQXOskNpO2QwG3+dy
hNt+ebq3OfD/VIZ3Ln79kYBFwLIij9u9hPSILLIwmirUNyG1tZPPkeDGgJaUwMI9rGo/hRpWwKKS
8YMEb+an3Ou9JJUEPOXEevzYDJKRJ2S3dt6wed+6wne2vfoXWlcsrUkiqIJu7XbnWDwT4YdC5q6x
sZ5WoqtUgV6t7gXikdH/5Vfym9NZC+n06PGhq0qEPaYZJe/IWAQU46pLgIDKkXj8eGvCjHzUdXbN
UOyvvC4XECi7X92NbtqCRvOz4yElVoqC9PnwFwUSVtDHmzDDL+eVlVIrmiMw6geA9X6raL3EIAU4
LtQ/QiorXqyfA7ooTaj/XUWs5dwKjS9LL4qgnaEdsQQzjlAXYq37bSv8kH1vjBPXNwe6u1rj7Jth
Ue6JNXVaNJctFhAHsOIMmcW9C5ljLKpI3gZW25p3dlBe4H3UnRAN30ps3qOt29ZzXLAoIgQHPyW1
Sij2t0aWV8+2ZKwrXnzHZLjhn1WwKPvuT7u/CJ90NfBHlKFavlCTnqnSQXiS7hynw4ge8J9zZEJL
LkJYVQM7uqjBk6Em+RZQAFVzqh5KKzCXDCkNvpmPQLYhEkjtZ1CqQ8QhITA2Zau7/P5QY4jdNDkd
Y2IE87wAzh12Rys//SofWRljsJecUFtJvrANXQGNG1RPglKsXV4pBMn9EspOyaBicznOLc6rH9V/
0kv3ESTgoAGAnA9x6b8P8NHC66Dgnj7/qbtdrOnFF5qEhWgzplODE4dFiGiymxq1d+YPUpE4FKAu
9KQeDUtSWsR0e8PcepllIVnmcudYv8lWxwVxPsebw/r8Ar4f4WxIRCNjGy2lOrkYtCNaZeU0QYq7
YGPBGqb4aSMjsoiWSzNIwaScQ/dT/yxXh7TqlE1TuBv8agT2yG1cdk2eJmfB0H0abVmraZPHmGav
l2QaiLaDQ0nF6msQUKsOwriYTsM6TIAl1hEWsY7MYof7PIOhOTUudN/oxGSSDq20o5koCbETkxUN
P8aWRkujkv3/zlGowfnCOu2cIsa9BoIzNbUqQWJ/h45JiSS/IaouoaGGZlp+xnmza5a7lxFg63d2
fogAwsa5yvJ/TJYgZvMVPhn/mMGA+Tsb+l9t5MZTuTmKjYCeyrw3nvH02fmB9fBeHpPvLcQS1Ks8
m8qyHfGEIC5MSBALnsFtkgsltQ+diF+4ziTr+bhkyKfK0nrtckHwr3iTuzOcd/wbvBv9tLauFBHN
rvCWVS0VhWITIkjHsqeVHY88keY0PXo3e6xFSV0hVTzGItTAo8aIG2SQ2gWtTQC8nfdhtQ4plgoS
/eRHNd/45z18bEYJEXx6iFhwtk753dQ2er79BGY89YVC479u6oXWbZK+5zlXHkUwl2W+ujqiqsZ/
J1gCJh+I0DtpuM6HSlLir58G90wRDh0UcwPby/r4dZTVgDpVg34dFebub2Z+dMFdtZKfrM5qpd+d
zdizDHE+Jh5dN0Rl4XFk8/z3EKDshOD0JK7sEzRl6WH2bKJVqCaORMq17YrJPzfY4jKai3Z/gm7S
vtimpOBbdRfZbPYHJy8fh3Ne5uwLm5HCJCZRGpSOZhMyQNUZhFkpVWBNsPQVM+tdMTLvX7+0uMfM
FRqNhDG0WTxg9mcny52OZBvmABOmgmW588RtECBeGZkY9U2Ol4/aJRBOmvXb/DBPx/4Nerqlxd7X
Qt4JQNQSRvbElR1D4jQ0A4VfuprpXbj6baU6Ax/EoFODZgZJz9BjDvH3nb7q7Uk8MgpHuuybyE9c
0czdOdL9CBOsDrzq5jdS+hICMPtxGMgMSHmvoaldRLUccvPPxPFFWZ4F9DmDtfLHTh8bdIWptqUx
6S3FvEAtxSZk5/VYriDandsk8YSFduzbm0NkEGtFoiHyPfyCWb8XnPoTt1ZJYs41vIOPXv2EVN3W
Q3jUo90N8Wqqz7sYg5c8alym6uF/T8Kd4mjQvdRXJ/CWV6NXphHzcunu8rtl1rYbv6MVEJboxk64
JXdDtCzTSOkdjmepj7FnkFoBhanTDd6MmZ88ALZQTd+wNL9e6bGan2SGWCIP4qHAGniJHkHv6bw/
g6K8gRqVvoiZWYOWXFYeqe+uDhkNQ24MO8C7NY3mIMd3y8Om4fcR1pjPjDqfEvP0hae9lNcuZAAq
zaUWD9nhTZxEtFJokgFbx9o1nmqYYphciekzuj4sTD6/K/N/AmBt77Xy8+ATii/wjLsyhuczIMpJ
x94IeSYTvtmOr4m2w2hSygnW/jwzyQ3ZxSUMhkeOG9pk6yLBatQZo3Xu1DE9aDR0Lk6HKNNnXXP2
L+tucyPuxIov4ti5uch7C/Q5s879EH4UVjmKb3llJ2+OyyJA5nXXCXgZz4FL5gQHN3n1ZQLHx4BZ
mUquEIBK2PunODIjuftywnwUT1KoTsIEvQrbgYEFe2TMeXNOwF21kGRUXipeUJB6VITf7OZF7uN1
u+nvq9x5HhkD13rZesmrnap4KBKUVnGW2gqkIpthDc+N/SKVs8sa5glXOVP/hJw0U4+35Py7qcHy
I4+8Sia6K7fWu3gLaZP+qiUF/kAk+qVHPyWNo6w9lOaHRTBHzhBY0mwK9Zo38d6H7gRuooHywVSR
6D5y3SIqUycsf5gELiduJbHX43vcMZ3bgvf/qZlbL0nIBps/dpw5rfMlhh51jO0MhWMbf4kPETmq
OZKnKzlO6KsBPGeHzVbx4ZdNZWysNdQmhMdS1CxFW9OYrg+gtJh6npIAmCkiydLpZ/gtHnHUihSX
gRCqIIooweDnfSiHUl4KNWrx6X5t55YmrzC6xvrPfQVjTpLNIYM0a0Y1uqUAboJ96Kx24edS8+eO
ntaU8rJnoIECUwFPvjZSw8macgZQlIMxAzNt10AKdsqODq4ATfe9lR+EkvdqK/n2+zO8KLvh0RzH
I6BJ9iG2OJQ7tW1Cg2sy7ssePKpLIWY30vzPgV89myb0NTPCoEvTLBfK52uWqcEsp/+ValWrF/Ex
SIeBPgFcbqvMRVBrdcb24ALzwJLx/UShPVutWsHA4yx8DO3AZQB64yw/qiggJAzFYdG4dp6WMxV/
a+34c44aqrYGCyURb0XwpuqgZVYJWBp031K1Ts2WVa8aMNwEzGTC1YFIUXzzNyqet/kDkv4mbOiU
xqrBTFhKybc5Zb8BzvcDxPWfIcHih071nu241xHPaLqPRtLD844wpejL8yFsNjsXRxPucw5HM+GL
YVvbRq5XXPN2rr/t8Gvzi4P8YCDqRmoy2nYQtTfgTQ7c9y8Zn8lwnsXPyg1/HjYGv3jZS/eqNlSW
kb3zxuz97X1hvMfEfrYJaVvXK52xSXfuG8vQYck94K7a4NXMU6YGG0SI7y4dMEQB+CXclq1JOHiR
6LrjIVKiJYTGoJKYISL9vVrAf3woXehVRAaErSVFUmC1d764gc3R68daXpLgzAPsnB7l4DM/gS0Q
dOSwjt5MTiIeos+5zsXUQ5zzEmWPl/ykomum1PBvANvP8+ZPQQxO9UQJ9PeuDXLzQ/SF5KqdqQM8
547w5aJKHjI2Sx4wB6eGsxEHMec/OMs76ohFTOArg/ubDt172DNNwPQnI8gtfIuLy/sHF2ugwA27
SyCacA0YZ0cNCS0SQ3sLaqrPzoIAto+VpaiLf8cF5se4p6vRVZeqAuzEXTd6hk3+jndgRIJXA2vT
r9UAevd9jPX6glTdj+8ubihIDuIAJKnoA0nkFsem37cz1LbptIxkCddzDQvH7cymer+5W66VTe11
YXqTs3jrNdnloriKfiiwfb7CgXp6Sqsnj4+OnF65uV0WE47jzdwyiDM4mYmXAvc+/RFjzKZD0ocG
hriKFrlxGbtU9mhQKOL2zX96sLdlgFAD9nxbQldOhXT4dSnoXFWyq150WmlmuGRVrzk7baNDkJOu
24yif9oEh+lq1RXSG74/Tc5oRnd19A1oXm3339Sw0OpPRTHWlCyn5FMYGDWpqwbwCzGrKeva97T0
/qyxXuqWM4B7H+nMLDjBp35SxMg02m4CPaFO/eTnJvaULS9bqMA4Umz98qlpTfirJY4l8G+COrng
E5qQCOKMEh9zhK/eVzy9yzAxrPmKOUEH71eS1coIYUDOOFzeBtY7sKiQpWKARjKr7vnlcThAwxXp
drLuXnUVqVC/tPKLWVVTymTnuemHLOPwiCi0Mv8itV8UbgvtqFrrS2ykSuQYBeLUnvhSxj2sk74M
Gi9qfztOuF5MJEIl5wovTu1iB+kqRF7gKAG7k04V6MRgqBHepyj6yhykpYKnssLwWvt8LdIL73If
d8GDt52BhpzKmtvPyvJaaPju6hHDVs+WToACA/y2Z4xLQjm7xOl8xuodf5BPHDQ8+8K1YI6BbPyQ
M4/D40mkS4p82BSnabY/C9KMviaMtmL5PRg3eKoI00C8f2F6NMp/s9WorNKuCkaFj/0pW6QK/o0b
1W8VyYoxclwTvvkIVxzHqb/qw2YoAYjoGD3LWLXthozIgZdszVEZiaiVFuIi//KUQ4mcfQz9ycoi
qlIWrXcpEOFgXEJx63ZGOS9fa5CNC5lExic83+LeqnOSlR9n3ieEyws+S6A95b7sYmI+2ka1NXVg
SUcQfuptW4lEVOlasWr3d5fUvEGttEPsmgD3kSWGKeUzqCwJaMQEcAJWqxqeuW2nTuWXpy0OXwIp
RRNn/ueKY2HFvpaPwjYgw3TQzFBq4Z/vf3IqdNvaci94yYUu1s775eeEMbuyomfqh106SIKSJjm2
NC3sIjB5heuSUUViZvGJbikxY3nUECiUTQzySN0HWb2FygNkC+W+wDI2W5kCHPAJpECM4fJ5UxY4
8FCp6fh1vWAWpfc3yLTzUVXsXLu/Tv9o5DE94XCC6spse39kYGhFUDqZP26qHPvdJTCoLigLAqO9
kwHbZfezJm9tSDJJzYDhmsiNlAoCQvQiQ2Wo0WRyUGD02F8aT+5aCpGRQ7QxIgAxW8//A41KcQ+c
tlU0cOGfu4N4JqV/+6F65FRWjkqrHsGQkRyUTuWiPCZ5IllCJhZkRzNL+j2lEWtCV66MSsNveYX2
I6vXXF+E7j2LNPnB5Mg+7O7mDVn8dLe0JB0UCuFdJCICU9Yufn6y26Ho0q78GuIff08qtoblvttF
tWL4UpiJoL8EHcrEXBaEICEwRJdzxndrMbfmxIAP2Gk5ZCxRiYrmcBS5fD83fdhJO5TcTN8aUJ+X
MU8UP9WMST9FKTmGJ8TC6zjDuURDaLwpxBMcIE4lBgz2b1U0dRm8Kslfr4Zh9WXVqKL3WhDytLXl
HWCDWyBCnqkZCgPkmsq9xqOXR+aIBbHpXYI5rHzjGx/6IuQGh7zPifkRjUDkE/sIAchgtcjwjSzC
Zi4oVCinBdIZvqIkOGK1tt9ZG4P3cit7js3wKJ11fp9HFgxtT1Rqyhniu7Cg3BTn/J5Rc291nNnn
0uGh62mFvEkuJ9uuRv2AOZk+UmzChOjsVtxRTJs/ZABb3b8QEvNM0uxRmlUzo93LwaR0OeGptNjl
wNrUVnFzAFow7wBLFfMjx8GrmoRFsRFpA/Dsxh0fsxV4o7s0qBnHSd3+SM5i2xy+ozrxvjCLgBUN
F4olzjK1Rq2YQheARbw3EO5cjFAU5JbGTYx8/05Yt8sggzjfZD47UJo1MXAnGEJuUjvLptfINy3U
IB3JVZcSHI9ZV3hOF8ovQZE+DgW0b1qTr1fCLsLQ9dB6+PdYStm7OmGnzfHle0OkP60BoVWgVZV5
QD4Wm4yOu+aNAfQFd2FAmMLKVFmC6H7Zf5aENmokeJ7BBDIdvchxsPlAU6vkzs3b25emkWLNuZX8
uUf6cAEsa9P1B1pOnHscsvLaz226gxMws63GmSVCfK9TsMRY24iDc/uL46DA5DlYdT0h5mbLqHTK
QFd6X5ihRkl0e5bssKbMm8sByL6WmKIDkToO6Ld5VYuC6lNU4BsWT9F1aHX1R3KEZdAJRqpjnVT4
8sD71nSE3Hlq8xFi4fKWvA7LAJq4sz/wylf1QtETyo+OpYMm2OJe5YeZ8OOd0jttD81UCrVCTv34
fpdrzxBh/YUTb5CI4cbEyMnrWUIWdvgrGfc2vFSiDHohByDzpPdlwDIdecoHsS/i49F10fSVos3E
RL9g8XC2UfhzsDye/CopVwiva19UB+G+3gfgOuwIGUiqpC5+PUptjSBVhOzWrr76/PLfFVlMTFWL
GuL6YANl3vHP6ExhKcq5TyaA/M7oziKL43Mx1Y6b8obfORhA+YmE80ZFtrD6bRqiaAEy+hsqgYBq
lDoBS5+6Cb8O0heMowrTxHPJBfBXllbMPmJYQ0R2Snc4K0ppcFs/ZjdqeXDrbY+bwrz0NyTPVI6g
/1JUI38jk54ipoDs+/eaIyLSC19kerg8qmGk1sMKlbPEtVxC+JoUDjL1Mh8pGrEIn9l7CXDe94DN
GGu0S3u818ceHExeWADNHz8fYgdpS0fXY+zLXc1v9kxmtFzWzzvvpu/lNb3PoEdYsZKqZIDRdZI/
kpe7OVjN7wNYGPn3UHJ5BnuBXR8QJSps7FYyZBNCr7d2Q6VbOosbyHJuHoqa4x6d//AEM6WAIl2N
G9T/zfet1rk9zRhjNgfPf1hTHbUxDiZ3OY5lvOtqaI7kfSdY3Gnx0G/mVA4BAPsU22KJ+R2KBv1L
W7l2B7vsTEFbE2hJJlQ5+m5mnkiG6IT6mJt3BmltkzbpkWcJnB5Phy+cn5qPUiBr49LkRwL+TJUY
hsMv3jirtwf1pZ4bW5pjYOPnLWabUe2OGEx4eI5PfSVtGY/YpmSayPhhXbmc08O6LYmSq6IB00Td
iTqzAKt3/sRq4OuNzY3xCgm2jen0KyiAeGH7uKyKHTNyhXhIWFS0YBml30iS2EoDcw7I2Yx/VZyC
YqwvE1radRfm6o1cVeSB/bj2hFGODpjV/coFnrHHKdzz2grDJriMPD0SGkqsuBf0C0HXl0jWU6Lz
b3dUKkCGzV+oZ/Te6xY+XerCe2T6TMKEeiAKZdi3ZBbLEX55c0NmvXNVnX/moBYeaAoK8tWH/A7x
DhEhdNI3th63qZM6DmGMJpQA7iHxDhCjfeod35GXEnvRuR2kaeSP+4JHx0rIGLYAzsih4E1rheJ1
rjs9qCoRQTsxt8q2rr/cntwwFomUtNPVjQegKS1Ubitwo1vZXC0oD4lbdedcRKrRZNGDGVCy169X
6BpLEPjRihmsWBhFzRny+XBqE7Ow8BcKM4b7n1VgWccuN8exT5ylu5hQ3LObk0fPGn5M/dY1PK7+
al+eI9+iWzd/PTZNWwvnJzI591esnCo39RzTa8iUBKLToybdo4EiQCDW9+N5sKQ6rijhUT0xsmRe
2xC5nbG/d1poZAKbtU4mAoQbwTS7UQjKA7jG5HFtFfMOZFZF8oMaIdpIaXFgpfWmkEKOx16V3jqQ
SsEY8g/zQUG004Z3WtHgfgsD7BiXsQc6M6y4BqlzwXVutVqaqrAu2IqGdz1CvzlScE6DaYlb/uQO
R37suDLiGQUm21XJ9y7PtYZD0s3UxQ0F9ptHJkmORvrz+6EXYj4DVaz0ZEhg1nokodDltKuVG4Sd
TWqhfOHWq/L3ALE1P7sLTN9+X6NREd0D0UbgdULJkIqqYg5fpjMyHh43F0a3XvwoYE6ZWlg6D16L
s9y3MSSCJGuc6ljzXs+jip5gPaxa372+LB7GmGgPh1CEWcqMJcwoh6+2Er4FBFoNPbKUzcXPdogT
Qio08xFOdYhLAnTsR3cPzk/pDlNP8qwWVegzeQBz46QMtdjmMqVGEQXRBYFji2kMkqP/Ar0vLH2K
XZTrzI79ASgK0JELDbbinn6C1CaBUhdQL8DnIXGcN4rDBVfc3/53v6QHv+MfWT89i7WBEzvHbtSr
xUcaSTUheW1fWC1K5bDBJPMf9sVQYnLXb9JXEI3r/rpv69w9GLWlwfgsaQNhY1wIumKKTDCcm+C3
cp+zNYH56KRQWDxKIG7IbbSae/rbv9hGTOuRlaApqKaTqiXo9N/jq7TmLik6nAhgkO9OGos3t2CL
S3uGsjoRcemppy9WzS1TgPUgaGIX4jWNFgI5YADfrqXQ/S+Fuq1v4CQHwXM6g6cjMfJMZznyxv1S
ipBC7CZ3wEokIgtA2Q9CmmW9v9PW0Lj5tHxzxRETU17erH3EH/ScOcJZ/2YUIa+UnqZBVNNGVNuD
5mYmAALTa05t+/VCfF1/jZXZSJHiKrJJW3u+EkDwVpb8qWiClqF5NdkhAtJioEVAfhOuFMBI9Cuq
CLX1WUXxCOXrl8sIy9CSR+HZH53SzvdlebVdE9gsuZOux+8pk9p8aP4uWiHvQ+jLVDvh+CC0pqTo
Q2hipTLAntrXRd8jQcbFMOvaaxhxMVXUycQlhEnbSYZlPX2MYCyuOaWMSISQBNIl4bjPnRMySFxS
85QVHoQQDp3Ee9eMIhZndNOQ0Rp0GRLwk1cLM0xv/h/wPuhEKOGaIcNHFrWYVS+wO5zfd4muFqP8
+QPAbx/I+xvWpxmluYYYhoMh6AI4omV8/yWK36DR3AoEJX0fJQVFqtT3+LsN4oIZBgaxThqdxY5r
CE+zUpWl4ZxM2Nh7R4Gzizb2RpkYP06XQ2+pRa6IJGZ3J2iAVBT2Av7xrYBtP3RWuirW6M8JE4hP
kXYquZH6oAT3ON5mkOHdDGATi1QZdvdR1gETim9WopbkuOae52uadM1DkpECJdxI2eMYEzwk9bTo
o9vcbgexs0mNFMc61xTLjWSHiBO9PAyTW8kac07pvbmf4qRQhc3NAuhWVCG32+C5YT7+Gqcd/b5L
mRff4CdJH2MSucRgbS2BCJH9FFcFBgl6AYE4iFxSD7iGPDyKGcXyO+mvsvMZ2gcnkGMKcQFt1UKQ
Z+0Xhkx+J729myOXLOEgg74gyMbSLaTY1pLqK0m/UqUuX8ViAj34zsPhkGg/blTEYKsesbQ5wXrC
q4zhs7UVCpgpNRRR/5FeYkfGMs0o61ePJI8oME33B1ZN2SboMartnaCNvzlQcKiskjKuMkUmukdu
PLaBordiWuPBZ2ENkUJ9NufT/+9by5qIQ5FomHH3U0DjePHzw3I/nIeOyfBHH9Zm7vhfoCl2CGvC
y7Es/9bTBXEqg+A5tcxuCDNjLzxFvL4lmX3X5RbLKHEIhlZu/S+iEaqnsLCi0eY7Na0iPa0NSDVo
NY65Vx3cXkIMIsXg6mnJidUWpWYkyFQycamXXWNDsOrSYaKdpKFDbxX45QE99PIMaudnK3tAv8ph
lR9teEbhODdJ6DIQRFTfdx22RKAtQb5iqgyXd9HyrTqCi4dGcrAJFdDb/Ye3Dg2Z2a/brweHk6cf
sKuXmEyJ27/otNrwH9u8V7Qdj7srBBcYx5nN+tpuso8y90q3iJwQyOUmhaSsmFHFvl3z2RbCv1XB
F0G59HVEKiTvRCrnfb0lMgk7zVp0+uhreg+UM59qp2K2ct3GqctODwMkm2fUiqKMNvx9x0NY1+fa
/cyR42HU1YOCg3YwdE9QzLmVZVmYqPkxXIydsdQWyfK8aToagpr+RtbpQcxGhyyhCXAu6znm+6mr
Nu/V0elFc4NWXfXtmB9D93/5E0uHc43OFj3uHNYSlWbeL6P/D5Lfp7Qv6rskesF1um8caMOfRxVz
hNYmz87mNBDkA6Yhabq1EuBZQun+aJZjZ7l/5BwxaaWl6QEziZYEln/tSG9//xTBxqZfxAElt84f
FjRCrKebvCXLdoBh5AnLxVhJLGMVzLKMam5NhUVyu6zGGCAS7SxGkiA2ehUQCpZZqLdkSvfHLWxz
ajBcOURqpjbBhiTHolNEQch0pb2DsK4mqBbMWv0ls3N8bErn8SUt3EsIU2uUgXoPESxlciEyTErG
yNyg0GLouIC3ZkubknNNwQMHz0C4DlYtpijjJt57dYp4Cc9pyg49MKlp0f6bg88HcRCghSsZn8ZZ
Bj1Q8lRCCTeJtuP1NTf5GYWk88IOR+zkkKKheJdP8tuJRRGKK1ouvHvTPFTTA7P5uIwESUuCtH8z
OiOqh3/TVyZ64Coj76ca/wkKwhlJRCrmxyDh+xy5+vIW7RcXFBxUzQAlw/jJf9xEK6G/PD5jtE41
N0JjNoLuKVG6M/i2F8cKmQf9IRP8YbFVsrs1An/w0selVl9sfV6WhmxqaBIZdBVS9PX4291m1S1G
TiBLdcW5tY9i1xaYsmVhj/MOfNkajFmenYy6XvjAA14uSOVZK+mBzD2IsVDo+mc3i8FH2T0kMuTG
nN4/kk8sb1wVsJ6qbDyNyEIPNR/o+SXkfnKUZhMpJwZWnKtHL4Jb/1wVPC0AssW+a74N/EZVuK+b
GdrhthUIbhtvflbb/Hmww7oLwvK36Xr1ie96ZjWQosr1hpywtBEOR2I1EkdNxetdHkorAg5lbAX4
bP766/Ggj9IP0n5wUdyds8gIt3i3mcn5PcxqEpZvcTxUJKYojte+eSgtGnHXMCtJUS2jLaHagfwX
GqzSGpaTV+2D8djaVXjEU5MscX3rgrNNrBc+9HW40oN7JDipBgzXedC2muLPn4bsqGksOxJXT8uR
Liwzpp1jWaCBpRtXkzWetCC67AKqdAwheJozkV2Lywoh6NSUTdsYTpKYFBdmWSXRv9cg9lla1wZZ
LS8QqvHNbSm7UtViz0Krya7kBNb8/xecr+1SNPr/QgBSuYTL0aK+7sQna0lINxm4TIAE3EtqOvlh
PVXNAEXdpn9q6WFQTbAOyPdxlOS6euB9W9jv2ENsPCyKZ5LwX7bVXrgjqJjLdBpRW+Ba9ugZYxfI
G8KV7/rOSStpMaL/sZ6nBbYDggiBRDCy258b0QqciRgwt5yX/SE5Mgo5HZLJBOEyqT7Nu58tMrN/
4MEaLvjFU4IvKWZvU3YCuK0XDUWNH5u3dNYKLgeP5Wxf3qC+CDBQVGRDTgn+aFjabobkSh/g4suq
08SC3cWgd6XK7YDU1lW3Bi1mJLog6sNl6oidhkeUS3fCLFFVZyqLdZchk9Yi+Ag2zyb3d02Cta5+
1Hlqa7d0MXMdGoqtCSqO/ndGsQ83nfyqmSeNOlM7VYKh5W1y1s2aPura2T8b5bDzfZo5dntpPjwL
/6/sD1HkiOPazFJrOgIcx8+7s0aIeQBsIddshX7xVKVYmmY0Q13E8EVlZ70Esfv3BWKqnwALDEg/
Fqjcf9XjwW4iA/njkn/eP9zTtE02WaKy/aGMOJhRb8dr8RxUUjBYXsvZ9hj5EseIfNZ+KS5VI1B9
cuNCIgOD29BwrORQvt5tavR3ohoXyzN4KcNskqcWkybnzso1/NJlyV6mWUfhOodkPNDL96PTbrDM
1FpzLAK39VISeDT3j1/cCgqOjnOURc7Xk3dwiCVZqmRrn7e7JzW4IT60DCXBNoVpSqEU/c5Hj4tu
FEjdzXVRvztTEtrovY4VDKCto+BCvEH/WMH0CetRw7UE14o19PMK4C8igbL6pOv0czV+960NH9B+
6mFhEarnQWQQXu62mvXffi88CIsbHGQZOiwBq5+0/r0pT+9RfTWdEOwtlt1y38LSf9Ez3/zrhVOo
umdh0aTXOvn9DXw+nqeZ5ur/UQlclXCBvin+rmDil6MvCVIHZEJKGLJSvX56wN65q5/na9WwWNZx
JVhCQfTiRkRgtHTmLM+5DtXaVjXmUf3kwaiSrYZf11pAOkpYEpJ6Bww+D+cRf43nfOFoPh6vdg9Z
lPQwd/vNPn+QKujj/J3W63oB6NO5wjwiagC4axKzQPGIKJ2sB/OU8L2/axRRtQTwoE2iIF/E8beh
ksKEUl2/1xYuNbxBGderuxdYXCNfbEL67wKjGW7MSvPq8JjELH4BWaS80BnfZgy3+Hk04aHFgidM
Bm/Msf3zIpcIXjWFRW87kTffs1EADFt6i3bxxz2qKV0ogLEesNmvHN47soKetFWjz16GzTGd4AHE
fRIXPxHJFGr+K3IZricScPn1w/GxDNX22QALeeTZi3FFpWQoadWjmlXoky6rPCByh0QBZx1TZkYt
MRUHHL+Qq5GaHakaxiEdUtkBcRGpzhOqbmJewuzGsdlLgDoyVgv+h5SIihMHJ2rtfnNhpsFlRufe
zGDbmnvsFYmrlL1Ao+ssgG+5u4gNNZg1yZ2DpDK0oOScpSMikrNQ+VBwvjTp79hdkF3ilSqpggKr
hUCzH+KoV/cxmnsdjYXJnL3EohhfNMdRQdIO2tS3o8Ajt3H5K/9zryqTDsHzOelElKQGrTAHCgZw
TqZHFNhsSFfTzjAiEyu4Sf+Hm87y5TpqHEN18OYfDyvrrZzJ7WxrIlU7JQBrTg1tmtzcOcgFzbS7
6L8GY6Fam5KRcTfVTuV1Po2nqVvp3C+GED1l2tVQMOjEBa8I0sidGiqpr8XQARC3wt0IxmOFcLsv
2MRRi6TgufLVJEhvbZ0NZm9vdBMSNB5d1No9ts+BL+tXqPmRE5NE2fQ+SJBsNF6oGBSCF5LdbOdN
JME9T02qffbTw2JkGSJXrfv5mbYKqdYOSU4dmsFL2cXS0RFtqnwQ2Vw7cAmiE5fJ2QRCDN0RS7X8
LzdPC9V4teDya3C3nmsy9DgX2H775HNH+g7dbvlvScrTfar9+vH5d9sv+tUYudd0h5L7/366LDxZ
DsL74WM06ujqlrXD0wy8wr/l84C2+Sg02Cu3dYUet8k3JtVbc3ekCRBVCAg55fpG9OWe7ZVlOwEk
X32OJIPBKsptF6ZelfB64g3tTQyJ+gGUtgK8GI1D10+sfb/CH5/wSIt5j4032OC6r5XWTum+3z5u
174zdRBbDTPxhyGRX7MagvEwUzxfGDx7vS5ReRCSF10aWzyUXwFHP3YBOMnZ7dEmNkCQVb7/v45v
oELuxyKiI/uMssuo77AGeLuwQE9U8PKSdoq97yrZLxkYegUF4xM2laKGvcO8qK3IufBQRij1zluE
AShTxyngpxMXpOR/pSQc2TwQy+hWYkRpbPAL95x0/4ZF87LY7cSvzWFm2Mo83VTZhc7Ei71R9xHc
tC4vieWKPYhWqGt5KFfo9BENysxKPTpNdvQN61h/x0tRz6+QX9PaPBnwW895f3Ep2+7WVx+KR1lN
HM1/nkmSV27g0CJ7W3U6EZTu7aDyz/L0hbm7KPYedYgnS9aGZKgqW1rZAeV9bIhTPDN/rFDyN5vU
m4bbxvJulV3xX4wtcRRYJEDmRSIo9bQJFf7tHXeOwu+oPLkVCOOfk95HxKVtPTNnnu+2W6iTsQbR
oGojigHpkXC1GGI3ztacDfogkyJ/zfGYgRao42/L3sqdWfBlV4B3LE2PhM5Mqd7qtnpX78Pf1qle
IQQ0rK665jOkZY+yntTrN20JoecPXTXkCOMkbvFlw69SIFHcwkHcAq3s9Hw9e72bv1x8UxQbzxW1
Gwp1DQAn3Nd5RJfbAjBYDnS2a88T03/0ea4gzj7E67dO9VTyjlF10EDAh4ZLya//cjd2p6R8XLMv
z1oDJg7vXbTqdmUhgAlYYT+BLpgPQU9kxXmJucEQhg0BSEmv2hH/A7pPsO0QA5drkGNEtcLqroVp
r2mK35AIWbGADknKKfcgJcRATyvySz2cAfybUbnwHNcPcNp8BfhkorOBLVCfZ9apErBHj4YxrvtJ
ZLOkrN3dy+HsOca0YGDVMXHmr96P278GzUT2wlBC8iCh6vA+4ATAuFMM4TvPm9id50LTSIPlDzu6
E1f5JvHvYbBrLR/nO+Be7l+yXW+85Q9zyjKLkY1nUzVRjTUIrx/hl0PsrHmQAxNQMrrlehJj1wH8
gvTs2J7IbFTkIQYsHTLNPCu5Xfbg77DTwvmiFn5NPVvTmWx9sgPNII79xfRsZVNKhDqShuJXXVrt
auLAOOmQtkh2gKrpeHamhZ1ImzXpzyuvA/fOi6fMCvZPbqv3PiGntmLVAOKjnsIhzo7HMchbpTbg
YFXdMkJw6j/HVMcS7CocQPpTkQrIGO/dAfjHqQk+F+Qy4/zwTnjMZMRZATU1iVIy17JisBmGQ2Gr
MYINoLhnH05COnUI4IwHBdobCN89ChhrEZAyTSP6xYlTTgQDgsPBl49mKd2G9WABpoIR4CxzXsOP
eQkyFT2C0CULq5xEggL1Hm7pMg8BPlc9Y82Zpbb1OOUjk6pC2Am5CJRwxKmo5KYD1ygr4ECVqlga
mkCA7s7imw3KJT51qH7dFZi4mHV3O/1U3bThL3uJ/dhGzOhgu1BbzLlmgI78YRtwjheEaNJq/e9L
yn+ogYBa8WUw+CN+664X24/GOnu4FQx8sj+fmn5iP5YJea5AkpooZ1c565ceWMc+cy/bb3+KSlmC
cY7wkJABq3S1t0gJpXSSgRQuDP4KqaNKWDIsWa9zOpId16SsfGjmoi4k9l84aEvbi8Mw8hjgfhLj
eK2szgSNPLR/qMUWheTxWrzms3qYokfX4YjUnwcO60MuX1e98WdxoGVb19fyZtMJ7wi8B++HkPWJ
DPtjEDc9vVYHRgBChQKpoUd5USq2UrdUXGO2AkZB5azXMMoPIqCo2z84Y8ipDq94dCCwSc34J9cB
kOrzJUifzhstqIBldmQs9JXfe3/1JUoOTygykBE7BT3KApwiSkNcb+InqgUz5lMaQpASfu1NYt6W
jLvjLxPGLKrXxvgQF8jRdNGha9Yb70aNVIsqNmNbd2UJMKv4VXl1t9zYOPpGCLxUh8H0zJbB5uhP
DtXY0gD+febjdwf6gsS8poEQyDvqRowhR+LyJIixM+t6WKFRrjIUqmQD4vGNElPUXZUDp9Pk+lVb
5Pa2BhlcuP+vU9Ez84f66yfJDZyKrIgxMvcguFmHtEL0NwVZhgvVFHLW/nKRL9nLHTvbcox3FFtE
ElmrPhR8sdqnbpSL7Dj8112XQt/SuT99cSKMRhHcE6jWqz3OGfCtvhYrn4AZQa3zp2NzM/OJxdur
8Cc4zvOeiBdxHGBk2kHb4gnrCO4Wm+lT2p2zHQ0FkIIodG3xge6fzSkY6uYtsHyCloMooIcvR9/g
rrSywAr4XE59ZilqPfEsV/3NGLpgDcP0PpWWDV/TnypeTdYeUGXy7BzqgHrh22fDeRb06krZb0iL
BY9EP4wEXy0MlV4ql2bhMLrVIN04y5TuzQHY399aV7Ax7EK3/ZUKp/pQqMGQBe+U18jwIsesQ/fn
J67mPfAOWUxwD1hVnJ78R6+SFNrldKZu2b7cobVAuuIm3y3fXNQpN6vVtVN1wVgC7qMdxC2POByx
me03i9zN43ztSgT4VFmsfpRKATrgwZBAD0m18/NYi0EQtyQUL1fwzelfAd5x43e9ccpHI/Djddyz
bpHeRTvEEB9eKDijnTNBOCifwJarmDqepDrcNNWAbYAKGjQoGAj7erSXruUI7I8pI8NuH5SWQt5I
DVGZ9lsGCEGnAEeutbz+NVgWYXFtrqWxPO8fzBYFnowirIq9fSXJH0IowPHOSLy9Biwc43+Oc1If
EY4MH60D/XoF2P8eRNlTLrpwB4q4RiGBVJE5v6c+J7bvPMx+cVgH+oMCmfDLHfg0HsA1d0ukgtkD
3vcFpcqhQGQQ1WZ++3VREOleficLxUlYbUQIbOH+uG37E6dszJDxU2gfr6eNxD3l1Wl1rCKv98eJ
JS2xg3s4sQiWKz6qhFeyhrIv7J0pl0emU8CnyWF3weR5pUe8hg0z3ukYhX6efFarq0JCMMZbGYtM
Amr3RHB9oqjM2wKhMsWRU7qXWUhimKvmGMTa4SMFRWytLLXE55o+dlbEW0qIDOS2MfRMp9/lPMqt
81r81bZ7/zpvqDtiSdc27KYc0VuZhUiFUUkk4ZcVOUP0K6g9E0SEz+Df8HUXg/xeaGM4gn7TmRCx
1grCEQWfFDCQ2b5lM3ziqLSNklaKOpgOhmX7gT4yQxFO+Qgiznlv6qMTamt8+syeKjwhsfXzXy4s
+UIMfqxcB4vM9xczyHSdK8NWFgfc3LK8L5ZHG0M/5igBubU5Xr7Vr7DQpBB1nOPi5wMCCPGtNCnZ
KXxJAZf6cIKrt2LPP4hEQhBmVgGwLapywhI1frWJcfC0MY3AvTe+WyrOfrAcec9s+iMKVCYLJw1P
6bv/Ko0PuMZ5kGozteHiKaOBO/YqJA95+UyBA8PSBZQ9Ub9t3KgLXRhA7Z4jeyik6sZyjXKP3Jf0
asIoF+vLV+cejY+Ty7Lv2l9wlVCwCE0k0fodyH21ZI+CgUBuB5moi6RYAIoSov0Ey7DsC+9PFUzi
uO4rgqXO2cEYG9U+sm8QVjyPoRFiFaKcamRiBZCgaI2fQQb/OlanZM/Dqc+SlwFrleI5G0TEVOmb
pDDXMZvcxm1pBwB2zUdpiurQxPhatydhV8toow1usN6eVNs9FqMkon62R/rqlk8m5HQHJo5mWTvy
wl2+b6iJSma4dNObTtNZl0UYSUpsdG222rF1ITGftFk8owK8OoyedUJNmoFo/FKzzi6TE62I9cTI
mSlU3cQVtLWeJzm53h/zA0hK9pifu/G+gubKVSTGB814tPE9jx7RX4n4ua4QSE9e6MVCNrKOl7WA
doTdc+P/jno+1Ip1Cr3eV4fUNRnz2gwTfbBi+PySMsSQPBRlTzck96EvBqIg9v41g23Ag9rSp8KY
ZNsApIgXT8V9RBvOTusgcjiWH6efuRkGA972/HAL9lM/1JJzZr5J6MSa2XUGtit3gK6jGPIlSs0I
tA18xypIQZ3w3iE66i6ErgVgFTcblKpnURJWdks3zICateHzxhhHbIJy97VDfY4p5hNh/01jM86D
zn7+VvB7L/FmBgzBuPSCO9TlUDyN4S1lxpwdz3We1VQZZleUCA95TSPGZwYM1+pZxWgKNYYJz7PT
gBy60NbGbDO6gHe9AdOnaR/AoI23arfqHJ6r+eB9SvR9dPgm9IvoDkzuXOd/OSltIZGDxrSGU8AC
FCosVfo+DPP9iJSXjmAut/46B95SlxbZSbZbO2C/8Fv+e/5cWfbKeuz+EGjr7ugRDzEBukr4g23L
OfOIfIsiF2KO8F9xRKHE8EPtzydE0o2K1Ih4+6KRNfJz0S52ixz3fRxz42yAhTjDb5UB7KjOlNwK
0l0Yd8iQG/TXnr3+AHBS/MFU/PogVW7vwt4JGwQSPSQzm5JtziH6OMWfN61AAX8yG/ki7bWiaiM4
ZWg65j1f+CBXktnlJteYuICC/5S2XPF0bosuUermlogRtRDlBBugcD5nQa+bKbfAdTqoHU7FASUD
uP652Owz0C2o/Q1Wnyeyau6fSjF44rCKaY7XZd5VunacqyaydL6P1omf3+pQzHqKP7V1n8ta7xR9
ZKpvUGZwvQr8/4dbPbPUUFf9RvtIX64iNu0hNHsb5JUpar8A44Ll0LfQDIDO7kNRMj0kG0su8Kpm
LF8NflqB75VMbaAORqXwUnC1MOVyn3STOyXMhxi7x/7qyxvORMvKOqbJAEui9NYr7KsxuOr+3Njs
7HFRTXcQQX/0SyuC14dd/mfb9UsAUpsJoReJ42k+pjjOnldb7KijTjb+VkT36bdXvMN0XgvYEc5S
Qhe9Qa5utaH2NvI0IX+HaPPBlM8bxNZBA5ifhCwHT6gywtJ1ni3x+4pQqt4uZMIojINCbdq0XCI2
3N+Rd+79VKqqVOsTzyAaQcsBpR1UfoW5SEyZDJfI+DC/Ixctp0RIfHcZequzF48+PQx3hz7zmITN
ihf1zhUO0ohN7PE4NHT0Q0GLcz1j71gxw7rE4v7CYmbTHsw8dxnWoZ358wD3ewbQqgqUABYoJDf6
WHOJd2WCcmGv/uXcqeGEXMygvBRxUS0/89Q4ayQ9BzvZAclFWTiWPIa+owVgsTRV2LW21Cc+eA4S
Ut8TtmPo35MUDqowBSyA+ZRyYMfNIHVmNQNWFJyDRlHUlXaKjNXktcFSLeIGIMz8xXLB3pLbeGCs
7D6gZNL5GP5dEPTRfdDlTRcNn6UzwIQK4y7SXi/Be6tDNPSsam2ooOyuV4qyKTqPONc/XwR8a8x2
qUkyy1jvhzoCjJ5lgl/uWZiu/sSbLnmxLPL3TzKSTXEFk4VhhjJe+GszWYcR9TIgsFezCNJOAP93
UtaI2g1rO+DqMm7KjdMd1k3qawPcUaBkIKyzSxsPXte0B2/fWYeT910+oX9ni359/zU2ka6Fubdl
Hf629MSodpNCNZyTeNi6RbQwVPAILigEo9RwHQkVyiTg+tus6VrMrYNAt0eLx5qqwnrMNv2GalFg
oqNUfoZHPuLhF5xoagpo9dowdw89DFPSu6FW2keOKySaIUQ/7rHLNwpu0gRyK8ZLqYyLzKKtnAUo
/VJTXVOhlmUKtcMiXpWT5J2ItUhQIlVkJ7mSl91ZTqT0L2FSm84PEvqMB5bwlkPf1tntbFfXtzpy
itxOEYkWOPCAMXVAI9iEiVnjlmE4XdSgVM87vpelYeIQ78o/8CJ7JpfYpissM2YINPXgO96vwuqk
0zVbWQi3b622fqQvizAbR9MF29KkM4LpaxUJ39Xr1ta9hawC86M4F18d7hgq64fVvdQidTSVLsxZ
mcl9kRAg6cv6FJpuQEyCfuTyY8/PbpNopfzaGq7Htz79EahEB0PGO4JId0v4AipsJfURJL5gIZ7W
sLP7fWyfNSogYa/dfI/I31RpVe6AshS7fxPSQx/GouhaPhUXyXLHPW4HpatNzVHZAMV4HZ7TLqwM
jnqzHD/anDxaySFwy1cYOIHW62WyG2uJbdj8m1aUkXoAYRcvc4GkAEsiCaRL6IolOdiB4Hjtfk1+
V5bUEXqIBsMqhZbKrPIQwCN3GtZwVDjhhW503YqbV7l/eBtwGaJRmPUWKJcnPgS9ARrviax2IZXR
4a128aHf1fgCE60Bf7uCtpKCMhvP1csb+wvvg2X6lOzXor/3fCBe5g0rq/EzMCY19l4/2TIHPpFc
xEiRTBmUamMYKLajD83YGC9p9l13wZM3SWA9rr2nPYAiONw8sSfGjkhVLJi/VwEFgufXsKHU8QER
sAsY9vRbUA+9nV7vW/nervtbwDYAqdc2zYmSItheASmq/YE8UxmVw3J3ky3EVLgcDPFxA5s+xQXH
obAO1JPebbsJrcZa2bHBv3N4VVl5P3vsyv8keWdT+Zwuen4+5S9n/Nid1k/8i3p917lxR8xdY3EC
0jvfq2WIPiguAYbjeD/fbMugwbQBxLQkPuNRBM69NQ3dUt5m7s2b5rEsgk56+Y7UCc9NO9cYVYiZ
MpyKfUlx9SJScQWF6QkL/Su+ey49kHvr+yU6kI82UD8pPgp31b/nyiBgm8AHQc+7KJYpXD8GgWJT
ZzVVLeYeexGaU44hEJHZi9qxW8R7fIZjVZ4VQnbMOAJ/85yCt0o/WaThhBEkzknkL7BsAZMPyBIB
rti5mr9LqhptEwSHUteR1v+ty/5GbPRUwoWphPsakY38ZMUiHEJy/tvy6Eu8cZyOs264TUQzStHC
3K+8bYlpqtpElu6wiaC9+P85M1LS2whXeOFnWcJ4PR4OSPj4kE/HzSqNqEhwGIlVOKme9IMLeLE8
RHjHjAHwlaRhXrkIEvmHTbwXXGfTQevWISOPQ4nC4jfcgzNdjH7MyS/UTfxzFlujVbKF8C5pP1pU
OpVvpWjZgX3dfrw9uM8Ukri3BsdmSNx5p7Gqi1sIO2RLlvnAnU9Q6eUvbTme1EyduciopbA+IOdA
hxkaB1T/yrKK/MGgR4jwpDPXOIYTllg62FydDC1s2Lr6t4H4+ue0jri5eK6B8HFZinqlhyM6F/NR
9Xp9xeLAJrKU3FLvRoeSMFTR5GfLRkrjdujhBdj/+mVtjGO+PkDUrD8KLKvVVsJnAWZVN+rY4DrM
Crh9zE4ka0a96N5siu6ilvgLNYXXG27BjNTgpe4GTIEM6VRFlS9wfbwSpvZ4Za6AjcO/GDFNh5uu
VryAHQ/mqHYLwamVWfYeqEniRhHeMcXwpqUMjfOE/Ld9UgH5Lg5IOoC+EeSFH3QnpfZPrimYalTS
4/URvHKzMMipg0H97skakIxYAuOqeylh+TTbiZ5e8g4vYQuCFy53yjqLJLJ0F3+66e5fBg6K0KPP
49f0VISAiY2zr+cHkWSbPiKTdPdan9Mi+7bos+GE37IR52LkWzCpGOMSdEr0/rZojUjmwNPh3+Us
NS/6Nqz9N6EISSoK58KfrQ9y/MtsrSc56WwjccL4qP1Dec9Rd5F8QZUVyPU+G25RqEK///1XlGYs
zi11DDvZjIKr8GyKFvanx2rKYvTn53QukQutrrUMg3vrL6XpauUYl+q1LPwIifN4Xts8DENxRUVW
nMV/uM+oCSr7whk6bBTqvRNq7/AudYRgEyKkMC9/tBGPOwxMHaY/2XPFO5vEkr2oXn85fS8HufGk
2qXlZXHuSgpODqu3eOHfIr7fPKGlBsrRzeNNFwAmEARhTae40LeUpwfiHMMDYzibvLpMek5SwPd9
utO/XPX/YouyKWOCpo+VGocaJcpZm2hlzUWf3SS2kqaQPMfUq7/UF4ja5oCv/W0nkjiEZPcVwct0
+PGRvEocLagfptksnRKi0hbkKAyjIeQCnN3lF3fclOh08pZdGPxuk6enPuNC90gswWKFqghN4DQ2
IeNBNKlMzfJPR1UHtxYCzlzwHXUfbUyl3oYQfbgwgmLM8z0eUOWBKVtJmfir8IqFGsemMTaxnJV4
BfuXF/kJRvwZW2ifo/zpLnAEtMiBYPXTtkIhLet1PsQAd0Th5PZzrU1S91YvoQW1aHJi+jNZ+Tmj
gaK8OGDOmamzpufBJ689A/TbO4CNnFborbxyjsmsWv4/DfG11oWCHhcp97KUK1VYCHgTb1tiALbf
g2xbATreH0IB27m95i3UM0c/QHAUwpg9/yX4szCSFfcvh9yrFET2jt7JQ4OLeCe7HKtAiWzlO6i+
d2JdEo7BaigEiCbkGc2dxKfyPdftITqR7zPX03xnTYKYg6B96FvUV2Qiyl70Cb6VuI4q7ayAE0SM
UqWyQSluLo+OxQuMtLSs06uZ+qPcDWuoaiJskXVaD9FyfiCIO9vw/ndWtpMUYspSD8mcBY5CePAM
yF/m7ohscZXu0Pm0oV013u/kqgdfn0WkZDyN7BLvDrYMNHl3NcDiTejXtCByvGoidI+7CZKGU1oQ
K2aikloYKE8XCpnr6lNVHR5a4o6bsxmlAerZsVNPNlP4orubjIgeh5IS5511Igf86C8Bvex3GrLo
5YSXWB3cThDPuXMG9VIjh7LYog85UJBJTQSlwRW8kTBC+b8sSF5nAen0+4IF6zX10Judgmday7zK
Pa44cjLQQvrtBWFLy9ZEpO/cFBC9o9lCMXTuyKNFMViuiu6e24hpLBLo1mpVkpFmd94muK1SfDq1
pycf2w9h7rFHB3x57KDc5HBo+RoHDet6RHnci9IBYo17zN7nzmzJtb8Wxz8MCmVDvK3uM8Jx+kOk
MEtYJ3VeKHh2UQXKqIyq8Ts+y8ZZa7QCBJDUxUt13Sye1/QR2uf3/vu3guCPTX+17lGw1QqqoqV+
KxClF+esmHNjCLcf/x2xbRTstjKvkVscNnhIrOxwC6onRRgIqWvjQtZbwlek1uC2Q2FF3VANdd/2
5Thsr6OmTf5xT9i9UqTRQ1B0zLogRdD+T2RiFV1Kh6YqxjCFCpnH9t50n142p6PQ9ssn+qiQ7rOr
CXv7ZYp9EVBrIe5QddefrfRP1eURZKEWTSwKhNdafR5nrc4n/AZP1ddvu1XzMHVYDu6kdvegnbbY
gnzrnZNnqfjm+G/ALqnlm18elRazz/vgOqVst0RJ14gauvdGsGDbrOtq29VTat5MaDaJr1s9m7Tr
x2QVgPm+rh4WNZTDA8brtJ1s2EMYQUiuXwr5zHzVEGaoiIABX8nEYPH/WVwzJ2n5NPR8iW4133u5
Aoido0stWgMAoRGZAOHy8iVoTlToYSUQqMCWl09gIsAkXpix09Gy7YuAgRrTCRAblePBgTCo1EPF
2khlxt2E8MhFRZRC6xNKUs8Xe10bDJejJhxPTFdFvKcaZJYASyQtTqIEkJyFxS8meowssDuwhujI
1btv/K9zSAMzMysdhI6UcRwLBCP7Cd4M1x+43LvF+QDV5j3F8gdw4UZYCVA/xb6pgTJVRdHGFG11
zHceTBz31GzcDvz6X6J4gp9fUoGyggDwhPaT9lsFZ10GebbKsRrV33wLblPufr5vmA1d/Fmb8oNp
C901zXAcrWNStizsZz7PeCjQiHWp0YmRANAgDo6GEebuTsduPRWu/WZWtSJe9tjsAfHmeyrQRoLl
OfSYd9ULXfAn//uyKyKKlfBDSiA7xGBUPdyCUKBHGsY+fsePrZzvfXNsF2mP3g0nqhtvWbh/U1zl
74a2l7GHtKE9pbfdQSpeLK1nyjVxkf/hjIjYHPi4BZff5XXzzpXTNmg2PQQP5hNlvsyBnwE5GEyY
aPPCC92IvXEL2G5sHXMVuzZZWkrD0/JnivqEtsYuF9T8QOaezWpWHSGiVjngWRTo15gA5Uko16AI
E3HySmMU/puvWYIbG0z8nnhi5dtGdoBuEd/lHBd4HY5f4vRyGjtAmIpegUs+zNBmEwZU6C2E638x
W4SPf33QBU8+KlJxnXmByM6P0tfLYHAg6EVEpgqfjLULz22wQdGraHcHfpcdjX0IBCSQQOT2iIqN
prVAIqyhTNwg3HxVdk/cQXCDIocf58GeC2Jsabi0frKCfQKSgWEehU3/zJDzdqwGB3EOnsYgEPuG
fTbpMYaMmjWfp4FzLXmJn9M+A//QXo4CD74HelzYhcLchn9yD18R26pkGQSOa8V1sHCPFyXnyoJc
qZsFcqBsZ5i5Rrl+FOI+jiExZmhm8Gf5fkHpSmT8Jm9l0rn3zQxsnfBvVuze9FmQWK6Oo9OqW/bf
AVgUcNoOP+NyQWukLAK0qPanHhkRCbSJl8m3A7zefru41Egd5/gr00UzRXBjdCRtgbpK5prdGjXr
hocdxJel7gxaCPzAFr9EsRSxcwFntQ3JxSSDDmn1hKdOg61nTjsGHQeSe/qoP5K5xb17igpK7lV/
7xOM6hKbmQeCDfpBIu1MYBeuJU+nOMWtK4dOud7TjXHOGph3hCEQjPWNH6wO9nHkWOM/QV/lCB9N
v4LoH7ri7xvIEK5u2ww2upZIwVRQSbVJIB7bgPZXZH9bQaAl03H9qwQSpgyxlq3MJP+c56B65mSU
2/NW61uVN95FbfYvw7BRmjJwpHySTbuXhFt7oKIr9RuhC7gpx9+BpGBPJVdo2GvH1x9EHljfu1fB
StDO1oV3Q64bdoDg291H+eFc9es8BmtbowKbV7gFB3sP5pxhTjnfuTYunEoVRPARVBLHbAjBKE0n
KxS2wjpgZbJbdOvceTuVjOBvhyPV7UqUcpvaEHBTf9eZGb701Im0ljAf0fkxRaPl4JITV+06ttvg
oeuRKsykppsJ8fKu1sHxdBNlQY0/WOrrT5QHw6MMCmeuwkjMJBkj0I4zlKcmK59oss8rB75yTwCB
nqexQYSTWMGB5WY+66UEfl7OEilVha61McCkAFKOiV+arMHhZ/9owRW/43miWp53RPcK7gkhIsjd
c64uv93ZkFLTWgtbjg3XPbkJvLu7YH6cOA+CG+XCr/Ia1Cv5IT0USG2d6NBt6TYKU+PcyVLGdosP
LBmZW2mJFFNmGJd/9KTSTUi6JwsVMGbtH33sFS3H6gQH/aILkremV6gXaZ/5Pe9w6QV3hJ2EfR2i
Oz97WVLIGnzP+jCCOZ5iGy2Z+mgr4ykVL0sqkR+SRoEmY6Xre2tXfZqGwSNxKP6Pq0zfhTnrQ4gW
dgkIOuKo8mqSDf8MuU3U263GXozN4TyrLqVk/gYKLd+SNjVMFbv9WZ9/cNE7eD4Z/4WOyEcyTgdb
I8uv16mVyPt551XrB+ifyTi6Y64WvDRB8ay5pNP31hpqrwHRE/GXDnrDnZPnyJXCACS2rHKJz0cA
aXTb3PlwSkYeLFjewseR3jUQzJ4LR+Hi198444K7jqEuQnkUtYD10meSpSC01GywtY9965SMRI7w
1PSK8ze8fhvz3B3Y19moQsTxmG4hnGtPGw8/+AMnjmKnbE66Hjer13IS6GnQWF+q84+IKC81C4RD
bjbiSOarRna8GNkxS4iiRjXITkRcgHD0mJNKfvkb0acSTGm+3paOl4ner87CkfJWhffNBdOCrOld
KhRFb46yLAjkdaY6EoQCS9goRpVxW2lQapblgLUL/ln58T3CL58B4sCYiYgideLa9p9pxw6Kpotv
vlzIWIFr9BdOIVsWcRSHR5y5/lJ0LWRFaeWjAWsnN9xn5qM1fjdczgsDQu+LOx6L4KPj72+ItjjF
m0qYw/UKbM6LiX75H14q07mH7hz9aYrgEakcMBFpEQbBLbNmjg7qCJysYz8uKqSVTJPPpE5Qwqsl
V0+ggZSMcFBd82VZTuteVH5QWzWCeE4Wr0yl0um+DrY3N5EZuT1n1j63Biu1Fam5tOVsReC5ZatA
+BlwUFjneqWRA+9GHW6pzGdR/jXDybxRSMTNEV/G7bUFPGl887FUejN4wtM3kO4KHbW/i7a6FTXj
O2/bTXiu//kVn/WhQkUDq+z8/PMBmDb5Fl4dC4awL0DKrfAgrOavlnH5CSrrzznLOxEyrs1PgrRo
gIhHlmX/mvyD8iIQjS9ID/7xSuuN4xQLuHvV8Datl1ToEdn67E0UEuvJhOkjNgAJgN/aS47m0Ald
accDQ4+t14zaqrPy1Xcp0Zm8bhhWzFdCrsokzgdRNpP3cZEz+4eEESUtLZiokddjJW9aMqrjZYkk
YGMcL56dzgNzi8AapDyqG0ymHd1kKOb8rF0QuCXpJaZAjNjpMsIvqW/WzkDL9CxHqYd9ZRvKko0w
ZJ6tXaabsfdvaHToreAnNeCZSQZibJ9rZPyUY/n8rZWXK02+dA/kYcIhFON7HP3LmMRfAZsqtP1D
pGraWioJpouXDkPvEIJnOtznZNkHViQjn0QTriXqKY5d+cPRnzAeoMNWMvJZ8VTylU4ViurALnkl
4W758SK1nSnbhgj7EoqSCF8F8I563oBxI006p+gakRMb3LoU8MFgbel/6VS10bv8XcrULAt74f11
4tvl2tMTiGaTqXjtulBitKH8RfSfnktq4OjY25oYGsWsS8WI3hD59oZM6krlksVmQtvyGe491tUi
4IWxsfmAU5BqkKOj6MK4A21YtoK0kAWw22ZAo6mdGApLrCH7lqfJNATSnnBKCh51kHA139CjhYp1
0ObUGIJvhGgODFGWbafAjDBPaGqRJA6utaZNpVG6vqYko3ZsLD/piPaTi8iujws+ZwR4fcB32DLG
ivkNNbELCJiLAKO2GueK7gwCwSJRL3T0Ey2cIZvdEsH80UDWBmW+/9KiS5E7fOc7wuaJVNl2yU7H
C10rB1UizyzOPsm72fgs0TmSeRNz6UJO4tFFJa/ZMWHGvyf6qaRufrK0RViLHy/o6We5NNe1sMUf
uo/z37WW3oGZbYrZVGrXWbqcngGm8zX0goX39RRzXoD2XUCclK+7UhZD2ToaPb3O6rThjAySI3rT
BoNOqXT+XYa5ofVFgtp4b3ccd6+tkCBfJ3FLAOhAMm0ntNC+l50YJcaSEdMz3K8TWdogLldPjt/D
/RLPainK3OQM4T24QEeXmyoIvZYZaP0wBGm96U34KbSN1VT9wGVcIUy0GEu4w3NsBvIxTtu3lKDP
sDPXcLQU0FOSyHuUs9v+hkKUsGkZyZTjO3dGk/WIlUhhEAIzQNDw8BO/AasSFem2xU4jVnvvRGpF
Xu8VqW+IGlF7PlMwJZ80jmR8Pf2GpMTz6C9Is1jvShwlULTtWZUMA99mmYNU/w99QzFyml1v0flp
sdwFWuy9Ghm10+6RM5o06VAlPK1Zc5qQgYNPUNSY5F67hv9HXUgX51glIkrUtAZuDZvKRqDWGiXF
HHEv+RbGvtTWQVaxzV3cohENb4uyRGrmRHFMXwzpOAbz6vlyZb/6r+4suFYUYcMmOqHodN3VPFEP
AoLajREfSIjLclD2PtJYxuYQiwc6PCszhbmkIpUJHaOezzRBvq4MyWn/+rUxyZTkePYG0JUB4w8K
xKL1JCO82IIWxGZFWauONVx/Y/ym30VPWX0KheDSlldJzZ3QWTtB9OJSDEWYol8v14OBRR4kbiqI
N1VW4kL+EHVHfs6WwKjuyhqq4Sg+2m7R53Auoibz8WY8/S5uEFsGmSctMGDTGWwdNhLIKR0tKHQ6
Pie5qrC0fIl1QuHy1Z+dsk9HaKvf7Mgy1I2zM/I3pZICDSPLR1xQcFpk5/cp7TY1QsHNrPBFWtK6
GV4Yv7IojiPii1LmoP0O1x6E5OYeu+WFq/iMRZ++xalAfMHpdt3kaX7kyOh5A/HLgmY9iZmAaHqX
VJNulAf/jGQNJJvG7ouKd3RNT6Qzpp8spvwAW7sWm9OzM2a/t9W4lH3YdVSZNLpGNaDFWKlQi/xm
gq7SAL03q7+xDumi8ieAzPYQ3Gq9fVpa6u3l/iGFxJXLBJbPOm/nNDgfdYks7k0Bglxx30pvscUe
Ud9KEXMJYaqwuvpOQstNluV0ct15HqMHkAyvk1VW8xpskIafLnQ6YCvaOZIh3syMfT4p3VxAQkMF
0RD3d2vdQk56lEGJHylwqZdukUYWcPmF/+muf4Ts5SMoE12ajhpDRiHEHax4E7VqWo8VsmOfYjPe
jL+ahL/VZufun4QY16Wj8tnR5bUXwXf3Dr7CTMZNrb0KF4HzrEfm2Jdaj21PJ4k/9cYAWwc3U8P1
v2Hz2hx9gDr/m7zu34KUvJGXNxuvLcCmkGb74mMj+xpaFgAbArwU6QzzQ0XEv4Grv5E0jLihUiX7
eChmOeSQ2DWvhdiGidtMhM1JnR3Kj3p0GXDWoaxIZSDw2+7HyzVG/N3PlMzQcgP3Fll9V1duUdtX
CJRd0KfGhm4Vw4HZYO9BK6AxDPymq8mXShLI26Kp1e0VvSZ+Q/POSV98bG28VT/fC9JDuKayeBIL
nDqWAoTCuzUZECj2zmM0OaYWpOTIQloBu8zFG7xPDyfT4d9x4ly1QNu+vXWoT2+AygSngrUj7ZYw
ic1ooNZ0oTPVU+mhg7hcYTE1apF/3RH98XIzq0jH/EuJDIfkOv2XwMOlQ3W2GgGCgGPHWt2iJwHt
8mKNutZ+260PYPdnT0FcfVqeDAb6AtBmv1diaPzNT/4K9VoK15tSHH2haMtYv+JOo5I0jEogAN2U
Byz7a4LIZ0bgfLdPVM1K+mllqAnMuce9iIuzhMVwOzYXac3kWdTLPxJYYHdSD+mIZMIN8KT+Vo75
4ghDmWN3O/vO7e/eNLGhT+09lzp7O2prm3/EeTudMZYlJ9g63HNut6GXPx62gSC5eb1rWeSxbAbi
IHbO4zJcXA1X0esyyq7QA+OJ8IULArU4OuLwO7Pcz+uKq+gkITgbU1cJ2IIa6+pg37jpg8OAJUFk
25qJE8KP0MqcMK5VHzsyorFB2c82K9Nf/OeJFsSiRlJmdA3ikXKybnOkALIVMfTriGFJZLH2IXHa
GwIbJDkXDpQ4aXDeNfQ+flzSN+Y3kP9UTqzKLd4ojaGS8YmUneByp+9uEDSOtTtLFBrhqAc5kmGj
Qb2nQW1mrYa33NjwCHdtmxLtsbrPFQ7WSqyf2Vizk3l2QL5ZKqTN3THcLh6VT5A1lFnaoHy7KwjU
yMHaXUTVAZUoU6qNaNJQ09GMtWOGFB4jDYG3MXDt9iubOJX4QlcMV3LPtJ1psEPTgiBiFdwM51Dp
yiVPHKpUYIp1SkKogZWQP7kwAQD/6iv+KzxGV/QRqo/YV3E+AJyjoYLgiuKhWSAQH+dxDMsxUCaP
4NOYQZkiCzlG96BFOgMOlDo0Kr1Rvq230RUs8kAOKF+rRICNJxuLMhFPKqHmSMClcvKmeVSY7UCU
l5jYdG5ZdmZGncUui84w8mZSsifag2TLzjfAI4Vy1ODh3WqbkEbvZe9PyHpjG/4DaOEKZsf5fqsA
uOefhAAeWGPAHyKvFytu5vXYNikVx5K92E7p9OYRzru+32vwBTYRqcffpAJrH0QF4XNo3yGIbuBK
pvrHbexfsCq+ovILGoY92eqPDSNWp2owOyinpdAXYozXF93FX7MN2rvy2g6ZAlkwy+466H4iiXEc
UvifWyuH+3Hekv9f3hTPWjHU+3IrzCiu9ylDy38JcdOshoLQEjjZFeaOG7jcaVPMA8ni6M9Hqkdm
9uU4GzgDSWhLYnjIrwUxggZMhij2XWxwrS4r0LmX4LYQra0VZBR/XSbhbH1wIL1u7effs/oOpHdt
gsc66rZn0IAsEDngy09eg68NN6uzoaCysTiwaKZMhK5JXy1sbAkEZG01wBPyGJXjz2R9lM1QjEeE
TEDgaxo0Ik+2KspE0bLeO1F6+4uA7ncAXC2JLFOZGHET34BneWbHfqSvyNfNVGd/RNfXCA/PoDZ1
sujo3lUkUsSAbXB/6Pc/WW23xra6dqH4rBZZiigGKJ8/LOqSbyi5odshSsaVy2RS8cHV9XX9i5qt
rEK8Pqd+uCr0GwQ1N0trKtHypqi3OYy8gbkBY6Mf+jnHVsa6lOnlQCdX8n609lVNv7FmPz2lEPu/
TP3XzlzSc+QAV+mzczYT15HP2V/AIbDOJDuMV5ERS2qi+djihER7/O1qtKepMWwFkZUHVHdCzEXX
UQvgMgFC2LPVctRAwDAdNj2Q8TVEKLpwG9G+F6EG//41MlMRJKU9jsFXftHiKRDcToeovGrKCMVZ
TGU4LdbMwcPgdQK0TrVtfEzbXuXcbltSWcXD9sbeLUk3ORP+P6SHKtH3RrPwGtS+1U21afBkNrwZ
RgFShIDYAYkvpIb9rFGme7SgU1llkXqptUU7E2piiywN0MN2q5qZEo9lNezbhU6HHVurlroKyl9U
kaFLZ9qo3phtBM5eDDGNzYgeMZlOPh1g4I3laS6Mxp8wufEhSVo7xjSL5LP2SnVSp1iQjCnXiXo2
oqo7w43z+5aarnd2YAFbponR1fTGl0JNNjSAuYYrJxGNLPIf5GBYUnUkwaweIl9t4Q3UWieNSIQj
moroep3jSpRwZVwrDFWfQraJNDc3d6dFrSVSrbR4t40sqz2nSpHpdkSCOf5XfCJbWQgHO+iMPwDM
1iYnk7z/ZYtuTRc6YDW1Na8jlJtLEbwacF/w6QTdJ4u3t8ZyeauYpmJYi4NfYiF9Xhq9BCJMiA3n
gROU1/UHZQVXJzR3IcxtpJHDzGuJ13Z5rdVxzieqw9i+VwFdFyaZR9frzInHB7EPciAZV/iJr3YG
D3cjJDykrPNNOddIj4TEMmmiio6FKjLk7L3Cv1eweK2jr2UIsrpHkRhj2rTppopSQQZwdQHVLWdo
b44AC1+W4N0H78NT6gb/zdEQXd4IO13WKOVxIB0T2Yf3vKKGMwBsfPRa0elhkb9n5Lpka/Fgl3fC
idXFLlwPqSaxZMEPWeJRnKXkI+J3KQK3Xz6fI3TvD9P/mv1fuZiB4P/PBFRhpVNNUGKaHdK3E1hQ
MToYUyeqUWQJghoZD+9Fy4cALz+QKIiKAI6mS+9l7BkqmUt571pUAsRZE3F7zNK1biNRDPJTqC8g
Oe2pgEGWTeEfAjtmmY+IZ+q4AAaJfWbIvl0K1apwWYEXv606AqOtLl3JJYqFHLbcWSzpCZ25FIsV
ORQJ5Aj1qmdjICiO2ClV+7AB+1sJHFFKrx0S8XDwsly1hxvWeQwxIBAU5VpPZzKWu15IdbI7ndgw
cVVEDHQ10Fdy/Nk6Dndt3YNM/hgnB4LWWMS/9iO25Xh401KPs0XcXPOsEAbtJIZYy/YLC0gsueSt
KxRHn4y/Bu7eMvrjexNn4mlbaVXauwFyGKG+cmSs9QHfc1kYsWuT6i5VZHM++8nMl4BX6PymkNb0
fGDRmqwSjuqUDiVpVPF3LUPIxznuWkfrAWph8AvRmgsfSmZ8SsgZrg9Xk69fMGrm1XC7vMYKHDui
fczY9LkiVr/GwUb6hDaquQor27Djh4JoCgEuQsdNmqEfNVcnkRrliydUiXzhWizgeswHkJMpPsIK
tanLygBqQYLP2UCT9BifXDt7ux9bFqpTyPidGjNlWvYD98XUobiL97vD7CUkKVCF0zrVfvGSznU1
d8YU3Gdrwu/KNPN+SEztJ6J4pCpapGiIKDgmBWnBfr1U9mCW5NW+dc7pGlEmItIiV2km4AlDcxhW
42H7FPcVXrHsKhptg0RxWPMgikT4ieOpsuJoHtHMD2vj9JanYbRMABrwiutiHCV9Z9Gxmdh4azxS
IayAiarXscJ5cnJnWKRWJMspe7ZmNnQKU0uT/7016LKKfn6KxBwfPONMMfQ6WOBdlyf2IKrq/Sty
H/KehM/9IhlmR0biSkOdZB6UdGmXt1tZLPbipSeyk2PUiqS+/Ei+5879d5VXQRTbCR95dnaKXX72
9TWd0bVVSZReueg+WAo7OxvoV4gkcqHry7Dpp4Kh9FNpIfSwPEjo/kODM7PeykCSaelUOCauz9zX
N6J1PAEZC41faOY1HeDPaVn5ee0jyQfIDizffr52ea54LU73AfHChC2PgNZEqMUu/xU59/JolQ5T
ignBsI8kXEpLmWYMMJwAy/B9qbKphchmusURnSpRKlyx9HXTjCUp6spjRauXjlSUyw5H3P9U59ku
FuSpGgOZFwJGb+YS6AEdTrHSyg3XMO0zSpSH7amDcKyaJMNWLBcGOoj852BtlikozwhzbgdI+2jM
BpLxLM/T/PFvScgNWpYM+AI0lVTIUlbYBlpRhlMmgvu/IzGZsbhdcLB9C8jKBGqxfbwJgugYPa+n
SWqv1enhSuEkGcqA9ve29xDnGM1GBA7K1IsHA8aFIT4h0CIaKrZ5gGIqgN1YcZqhfzO9jIinIujP
fsgOOT4v9EJPnGda3qZq9kos7xPSWZVtJ1qkQ11aLvLFthqvHKzEYPjCzTpyOzBcJmFJt34vFhr3
8e4+k4khHnUcbbOINDMe9iKsYM3GCp0RPbdr4U54OcT3Z2g0ZOGqvK999FOVCTsWjcHi2R4HZUV3
KDc4vrpDXA0i6vr6uOdYWH+YZ3YSjdevWBwQmZk4mLjPmewUYjConqIX5J7NWEvMb5rUY0twQZMi
qqEKAZBqPveOpgO9KJUtBII4muQsorTxk3Q5UCyoDMUEELCHkRchHQX1916+ex1ml0wHmlhDe3ja
/wJ6Rd7S8Y3W/0Mxjzfh3vAH48/+l+FOqe6t8GwIUCk+u8ElG2YWsPSaZpMVPN3rAQXw86Xtp6/Q
Kt8uNZkbLsn5YdapJTRmvUY6UApEq29rhyYwWncLjgbph7hjKwrxxhz5rkXj/p94qn5ZMOxxbLSo
IorRA0VG3HV+4ZX+6VCxfR0RVHoMNriLIbqLskVarKSLJiBWyzTd/7U2Dh2kHMIApQq9wds+jWZf
CefE/D3GpKbl9DjUcnd927bHtGKuQwZJ5H8zOp6bc0WSueBgD+lUk/gF/GjE+N5p1J6cm+5cANXI
rB8TvqeS/2dTQgg+jIF7oz22aGLQRgj+1NZCABsUvfPs94nsDnQ9EXTAO8R+s4imjZ2db7yvuSHI
0ZVmP4vnrkc+dgA3ngcHatH7uAMXT5AFrUmLEgAH7a+0XDn0lB1ZM0Bf/8KpC6hdX0YKffjoHg+7
PdO5RM2LSzl8h29uUbOLsjl+WDlrjIHmyKqdCZQJcJZWbMeypPQqMErrOHoxs2syVA80okiBv4m9
UtM+O23SN/o9RpcDxGAdDzAcXnMOAfcSImkaO0CSqOF/lAkBYqH8vZSWlJawL6sFypDlEGUTPafO
pT3KHZ+tDFj5mYhxxKLu0ly8NGue1bkngh12rMxqmu+D1x3fcntjGQaMmrOLBhyry5CWyvpymiSp
3N31pnVhCGjfzAc5tZNbocVpSfiHze9EPAfPrnXlk5VEywik6qE9NPf5h+VVrPQzpcxkhPSKIApC
wmyHcHm8CT7VtlIY43Qt8ALtCyh+A+q5da9X1qJMDrfcYBHnVJXmgLFIs/Xf4TFJrbGkzNwzIHni
36i9S380nAqAQ+79WzYXsTglEqqh3iuYElIP3u7YRr6z7f4EVPR5ga7K8DqfDVNDrGolJJwkRotQ
TTw4z8sE5yovpDI8RRMnmFVPJ3harLypleffr206Utvcjsokg2oDEAwYAVasWAcfQwMHL2i75IJh
zKySctXe6a5PQLpwTv5IW2tFrgUukrtjrZ4RKU/Wd3tU8gh1W90pG44HXxtAgcZQ/8wOcFzItDSu
8ld84wkB/ZgncPuFQQ3Het9pv2Jdl89u+DiyH1Pfzrlt/nsMqEIkaw15hAuc71VJc80pk5K7sfWO
TqJzj8Wu5gMcGeD42mbwzok2YegQrEsh7+tgevOAMKn5YKPqcLujnSea6MtmINAuFdDtQgssgEct
vDLizkt5158HzQgJ6HiLzl4QVF6vBPsjvYTgCWcWFIAJUj4xkTt1X5xc5gO9HsjJnuXIqKU7LXRJ
7BxH6cDl3n2nUDUF76nZTckN64OAlQwhqas4cxuPRutuEk60OODeVIts0Z6VueC9zEJEHGPO5TP8
m4S28MAbuj3ityDIV6x2q2NSkSRoPeIXgkp7aVNX+uJq4J5xU9ZAxBoAhFIAUbr8p7SIkn5dCyX8
uofHtZmb2UyNpa6PlFafHLK7VTDrBsPDEzV6DFZe8suCbmGPxI89NJvlU6t45L3Nvoa4cpcfd//q
1Xmpm1C/W27n88tRfPxZqSLN8WO6dyCMC6x0eLReOh6RtbrrrGoY3mFUC31aE6NBzMhl4QvACV8f
poC9ayY3tEiW1ObVcV3mRtQuAUS01jBRMEYPd6ndls8nFdK9i/slJJ1o5MLsA9m8Uq3Vv+Ee4zIy
PHmxQ3xFRq6zYQmnm3VqrjVthVLkkeCHD/817eIO//tzPRbMs+5jl3YMlWzMjLNZdbGfYeRZI9DJ
G6G5JiC7oquOBlDUC2ale0f6z7P8fllumx8ii3/iRgfHZYoaiZIQ7aYIrKleueLA/rx7FVuUogVE
nlrRwpHKiXJkWIpaRonRSJldxBHWrE2wWz2OsJVrQ3joDfgFdyPsQJ27tFNuNeDLqrWK/Ksr9TEt
yp0crJfLnS3eyXmHcrXFqPlDW649T6J6MS5Dpq1YmKSKfUQPtxUlG6yqvphIXzlX4UpZ7PTDFfoE
ossiTbeiiw3TaOuumYRGqqXKtqWtdWDvg9ZX7WSYfJg3YUjv8i9uYOYxYm11iQ1NcsqYemABHYta
4mQU0DdPgHitFk+hWOD91mBM+pvTY+lrP54j/P+hD7Y5EjqgD6tAl3/ccUBCXtulEynrLqXUj586
ioDbivx/HfJW/AqI6lR01Otm3LH8bDhxmN5OZPrAOgW/MCaj6ky2xZwGNkUlxpPZHXT2w+nhIaYt
+JIFn0p6YS0Gn6og5WGBqhQZGbvuNWw/nq/dZPIcHDwbj0C4W0uUROKErL3ZNCQYvDoIe7R2vLxq
HALn7cfMfssjgU5M+9WuJOSHhYCWBznUjj0Gc+Eb3G+ud5Lw50K/C8vlm22ztZ0crwPWowAkafHp
GZ0YtK8rmZbLKTfowjqzLIYgxcNPR04N54HlifVWonAFtro3Npl7GLSXjqFSMzGUu2BaaxmCdQgC
BnGxac135CrA/Ew+ucSIuQX+JeXFpHgyIEvL8kOJoSOvGQpMaGIB/HcQeF565Z9R3SnvG0zFu/f3
CblVlJsV7M+5kEdWcHSMrj6tOmlwAx7LRSwpzJW52kLMDMxIP7JHk7b2LN+XAWb9HicQIa6dpTaI
jxI8HcyjdYuDR/xAkjyjn/In+K3FZMOHiWAprARsDKqwyLjTGltu3DQArWlMxXU/92Z7Jf95FA0Z
kDsgTp2H2XkwLcvtwUhIZpThB9I1w2QtiwehvocUxOYhBQ3GJNYJ1HDrdOzA/xGHDwERrT9156kA
GQ92h3GgSJWRLKgXMJhvl9Rd6G9VUShSeTcgjCMP7qD1NO/3bgtHGhTcJ3fdBrhj2fw3SRkJqvlC
QrxqD7DC6guelg7KWUrMoWxR/t6QvGONqW5lU5xGX7swqessrcPSoySNWmHZwbrhpmtX1LxdF2lW
vwycofAiaRbeyMvLhTPtgV6ndNi3+fZ5SeJjJBkHGiHt/ASrSVRkMprh/AXoGo5iG4/qHHZDiKXM
RHBT6irqPFun/8yl2+i1CzO1lP9/4NdfZsaW6lLNZAY5AF6VJ70RF+cEC6OtdXMqwqE9w5veFgf6
f5b/zS/PnCEEH9ZDldIHEIC9FxrNPVpy1nE1mo7xp464ztiO3CX2C4qFxSS0ZT1EnBNZyxhSZ6qj
/jp4n891Xlbz6AWNbgiR1BtVAypZxSFs0ffS4vOXovlR7ld6X0LYSXODLY+FYkd2U1KqZMwYjDiF
U2qZRaWqExfqyEa0+/uL4q7yohkflV4xna0oaHyzhWafVhEkYv2WLHfn+wQNQ3yiWoCfG2xxwok6
1Hv3eog7kjfYsXUw18RR5kG4j0V6iPIMBKvuga4DKdrZ8bnM8hC8cmAk2qSzKn7vwx/PMA42FuUm
hVF8RmaERW0I/3wt/pA6EztmjVed/Pfp+JCfpqUqRfe1L09871nsysPqqH3lT7s+roljTJMxqRlo
0G493yhd0aKlaleC9pX+FR0buwoC/g9Y+rNyO2LuJvjGyLC8geM98FqOGft5P9Bb2VtlSDpOa8eq
6UPcYPJHPjvZEJtkRrO4UNpwABjLL1jbCN0SzsrME5y6rskz4qbsSKpYGXk++yBKatrohlWqKJzj
1zRkdGc6hrt0lI2Iy+o7o0hT8WXAXuFE/mvyB1eBY/bAno2WuH1Ihgs5pqlI8QIx7k/wUdJsi+W+
oKCNN+gzGIGyn035n2OVLWarTUK2N+zvVf1rAVh/IywNcD2HjR94Lw/F+0adqP1wvvFfgWwLD+WN
OPJeLTL2eTrW3W1IUY/WEM26ZgmlmgXhPB53haCB5YC5tzmCdQSnChMX4rhqQVpELud5enCix2FZ
xScFs9J3EHjx4V7ie086FjcSbsOQhm0TSjitzpQFtRlbhYO31kb29XrTQ4f9XPQx7vGG33jMBq3V
as5lnnET573kQlNslLHyR2YjPv3ofMX6kwHShNBeyZlAetNyIyYv2wZezo5XuUHQ5O/dQcoqL7Z5
L8ffX/mB8xNX7Km6IDHUO+0e+xxP/KMVBza0mXTgOLfqM4SRJy9CUo6F+LqRQfVNx5Ygp6QKvhHP
HuzCOXkkunQRO+auOxcM2RpI0J6WKN0npt9BVax11T0McerOysaa7IxsQ4KUl5zzrIH/OGzQzRXl
dlFdA6bdXaJw5EV4Oy02ttg8+i8CvTjihwwgP+sP8YrEfRf1uk61ADTLqTpBR6lYjn+SKMjS8jqa
hA+7gz60SV0baX+edy2lGPGbvJ7clKp39uG2HT+0ZKX6WV+vV3m552aOqa4oNwgzq4g9ps018kWR
4s7E+RUygk3/TjhWV3UNuWQ/nzBP070IxN1BxUVJI10ynyJF6K+t5EgO2Fb6xxXqC9wxvS96lAXP
S2AAkBsq1hjpCaAZTP0IFdZO8dYtVemvvPRzLJ/b/3qolMH5zts7b+FFcR+IdOL6C6pDH7jtHi6l
JgE7stdEIG43JdBtim4APvm/YG8XYretCwLC2JiZmHiRlrHffQUVpB1y0bdUMyVpqlek9oxPFEfs
zdgD19v42TCGwI0ZcBBqHQz+Hxw7TUolrt7GCSg6mJ2DETm2u0FU2Gm+Y30JcEMiPyApqld9nS4S
RvC5t9SwftZYxlnSXSUoxUzxU1IbSP/CMYZ/WoaH5jMZpnh8/5kW4+6jL7b0yKuHCpbQvr3Oqloi
I6/Sp472B1CTi4sXS+sa4egrwKuqGDN+diQi8/yr0HR41dw8mbAgDdU9AjkdOdtNJEBfbr4Y+LzQ
tphKtGj/OkesUouXxU5fFk9F9KwbqT4ynImC9R7P/P9M3GF5NNUOmmxyQi7CIaAgq4HtRUAl5z1J
kyCs4wSKLyQHFmA/q++6Vm8AAcLDcV0BUns4YvkduWzYgB8tFghceu72BV9mvWA84RfR1/oWebbF
vMYsUwjnJU9hVvFLjPTFbu8QohPyLy0R+tyr7rN8eQY28xKzsy+vgnGlxp4tnd2M/yP52d8NM6gy
Uuk6adRsw7OKkf2qYvU+L9Zi6Yd7WvrhlkCK44y1NOZdvNgnrUynjRSsaQ9MxQWI7ZBTFTDp6F0+
v/f+4IMAsGTlTvkS7dEyEu3iporWU9h17IBOzJuJh9lHWDRnwfH0TdZ43a2dM+AKnE83NJyju2tv
ConACfg0X37+ywfbpoC3AaQDgt+MsPBgDUD6NvR8mh0Yy9Evawie8iF8OQNQyHZTvAM3JVKy5A38
Dq3/Po9H8tT3fTWGsDngMb53mhERrJqzklLg0svq46a5KfwxHDk9jhAFlre0HFx9VWhV9RoMCWSA
ebB4Z29D6p2UbvnDhzv5iJmheAIBDI3WOcvyjvzXbMMRyMp2UFJyqGtL7jploLELnUXzLxnAH3jz
89gPmWVp/xhySeQeOtqucxz32CCrE7i2pL7SOe0CLZyvUV/Oc9PRNo6W4ox4CdNIqmQP2BW9jGQN
Lag7AnbWcHlafhrnrOqIhEf0iyf9pBLxsRfj+RRLarvwVwEXc+mBOimvUAJEoQv7ldjUfwqD7XgJ
3BJ/oE/p9UrEt6i3Ju17KPRPh6SrD2Du0ZkgHpD+/NHTJgxN6cCyHCHhjaFslarGUzTHw/5qGoJR
+MW/12baErX01HZYcF0XAtXuk4LqksE4QSDDxltwyiITyw4FWRdBVK1j2ZkM3Ai7KJcFpF7W/1xz
uBd7XzbbgWhSuhHNlUkqU7LzIkIQvjFhaeQLGAcXpReOdsn+CdMdXHcWDj1gmCkUfwW5O3uhcyB0
FkvBvscQCu4o+S+9ImD9WmL884WBy/hGoCPRYAj6ljq9EuhoVCNFjF/D+LzRACr1n3HCzal3K08G
AwJ/lPbElynH9tIpMX5P9XOiPxnP1kebwQ0iy1oflTPrwlX920LFBr6qXW8nhEmb6Ff0bDO7Uwrk
O/rr8madzee1LXjwEK91FcSM8+jYpUPYxhgNauL5HWMhE9CA9sl8rDgG+RBnmFGDxOMOSkBjbTuj
Awc9Rx0M7VD+ExyTOHbsvKKhELzsGgjI86RincliWoPzOJyVN1+z2ADbnfilDFGvScv168mbUZmq
y1axPfnISZS+QJKfo319zsHOEgEbtPaQLGYkcfB/b2JE7oCoGlMU1hULXzj6uB39dWb6VouOnaCk
FNMT/dGfqH0VsqPYPZAn5RJ2F7G/dtwr4nbufubrPJMn4nyZNJN2etsZdPMyNJCJJpx9wxVwA9KJ
b+CjV9KQOl54IRc8pw2kePjV2SbBzUKY5Uhn+DIC/JX5NdN04JlGoa4C8uVu+0Jcr9ekYMMqUKI9
SmAncZjigEZXnxkrzYBpL7MpbsR+rGJAwnzpqnsuxuKacNW2fhpJLJHKq5RnAHSz8SA9oVo79wuV
sbRXHMb4xu7TjeVh1jrcecxR+6i/4RJKVi5kQGF9FWe2w13xtILApuStzczKsdxxV6u6FwaznJcL
h656FyHfmznDmMiZod0DV9Mf37JPqurOfAj8kxD2bZ/s+dKeiThridakWcWPP7SDMUlXH46mWcI1
5Xbef6lowG87p+KaueCp6BiElu3zZtsyL1z4NHbkYQ9gl+SQIUfQugnj8kBndcllsRGIEhZa2YFc
ZdJeqAIv7xZcy83hd7k/zAn/lHIZFVjM/8yhbCGXGQDUYSgYzQ1z9Bry4nex8WeFBUSr5qrgJ1Rq
rbwr7kJHvnkvLGWO5PwgC6pStcK7zaoUHV8J7NBvcHE9KaNkHyJLIfNb/L1PADR6MuH/k1whsDOf
gA10fUHzb7uLvXQVQ94kvgkQUfSJLYnic+O3BklG/YsHDcr0EI1Rqf6sp9t2i7qnKWmoIdV4TA8N
imkeS4KdAQvc3zzA4Zqc1JZs31XE3reWPB5JYX1O1yQn+9JGShC4P8FA284UUb0q1ImAYKzBqOr5
d8v2SdJeXo8H22acno1PvtNQVKl99PeiCZOCf21/L3RGD5q4pkaL61XXtjx52BB0L/bD7+miIyJ5
1HJmpLVS8F2/0eiQ3iqOLksNQlBZZDHk5soNUWaMhJi+OwKqU2bo6itlhenpdabJTUDLngkF8IU5
Aqu0UyTPLtgsUUiKQWV1DVY8dwGmYFITF+BmjLi+btdw2LqUVrrqx/PKNEx8+D3+P8mDldcEB9YV
X30gFvVl7B7izd+UW3cnagKOlGxv/bdcx1UKey3KVdtGZMkAhaLqxtbt2fMWrj9pvgrPWddawwVn
/Yvss3lGfAvjVzBGhrmQz7W8m68azwts009hsRlv7R2ZC4Yi3BYVHDpd8pxgl6igM5UZGtqxWEfL
KJwqS5mLNg2EzI/GvFHzF/2Gg6uEuNH4W9NJSfT5XOV1yk98Tg0wd6W8PlR0wJ9JkkxIhUmX6ZSI
8kXGvGyZoOC/cTsbsRgAb/C2D2ZneY9pgffoLRVpb7LYqzX2Z0mpsYzhtKdp7C5kpajhWYDQjMlc
NL7L+a1+0GfBeNyfD6b+dCSQc0o8SSjvynBChOZZ15OaPJorieWVFn8Iu/eUR+32DoudIu/z2xjD
gXKmni75eMFk4DYvexKS7r0mIjgYVZnjHe4kqYe5vWHlxgDAbPfRLFJ9kxRwuD9X0qNOiaMXLIyJ
X7Qc5jPp1JoLYDqsRLBWY+NrHbcOQjlHUS+YcpoP6KQ3F1MeRkb1OdVYVQJdhGqICLF4b5YupF4X
DAvVrzNukYp4ampW6/inOQtv8NhBTur6/z5pMWuNlXg82yN6H7O4dyPpssbB5LC9RDax13IlIye8
plXNWoFkfikNZdNXfHaBSJjcmzT4X9C1oPSRqoEKglw3ZqNqo+RmkVolzh/unYqwyTHJheDg/7/L
vhhGY3zgSQCKjEYQcYYGUh/Dh3t/Xnf+wNlq4fQ1SxMu+DXgyL+8jzFg+7dPqf/CqN+pYBpWvS4Q
ZmhKBk3o8D2lLOGcnqQENVqqeG/PVi0uwumgx66WaVMnK8yXwD0pysRcMOSJN1yZbX9OHdboMU5j
BwH1APCz/+5C78+JjLq64IWBHe4imOTogd9cDddTukkMb1YEwlYIudjIFygrz/3Vi4DrvtvX64VL
DG84pjcpHMpy+ofeaVYtftmFaqTf5Z6FI64+i4MegY8DFQr6z+ZSAAnHQlkM5e4X6WecKBYLlx/8
O04qio1Papl+VCUcYyRiGmGoLrcVFZDayJOqhhfrlXUO1cVkttaYOCdYcQSLNcItcdCkxSi2SG8B
fqv+Fn+o9hPCh5qHd3p2geIupI3iXcVall6rb0ymFWMGCRLLhKKCrq6WhE6avl/S4QPL7Kjzx5hf
lfZXmp+CZLBucEPLnj1H5wowszWgANota0qJxOvfbUgZLvDIBgtcT3W0T2F1YXF0itL/iSnqPqXo
8QIWBQFtzPnIk0dsuU77fKdyx9BqyhW5vTsz7WgUT6LLdkULIWl2s1X4gt/j7xhcmNY9SjX2oamh
9jzo/VOVdYwMi+moWiQ6CO1pEQVGwQfsz5kknsPYE3wi6IB2a83Ert0Gb4tkTL4L4IfyhLwJMLVU
IHRs/oYzc8lGUpW6fJLx5t16J740QYdawCDzlqX3xN3OZqZKfeD3NOrvnmaKGeFUj+dt7pV/THdF
inVNmtW87Ak+4FiEz+x+lFshga63ms/52k3m/YgCzirWu8kwuEX89H1bx6mhclEMfQHp00f1MXTl
id9O4xYOZeRlKKgnUBGF4psq1uCZ/sjNQv4IChdKz3FelJ+kDpM1bZ44JfZapGUQTGLe8P2zb7co
jFZ4FNqPnQA1TF+meX6P/VfT+CosquJ5eE4gJGJzq0xi9+JZ8xZVx9CgfMqEgDTySVLd5t5BBnyj
uhCZ7w90azm2J7G1z64scbB4HTXBvPBrg9xuDr4Kui78Zt+lDJ9A2K0lvtajoHKgNdPBqqJbyUp9
pxUrngvzSZjpzbafmZFiP+PXkKUukN9wKLvhTSQpZV8e2tPRVfiezX8ec6juVQhQzFkiVEiPlqP4
MOEeX2XZRuAKhP79AaSJZ+M03GVukApcxYoPDxwCnXi3tqWLw9lOe1Sg12SWM9ke3OgpQEHonZu3
v9oerG2YCjsoT1MNUwbPkfzR4sWCNM5+mSQwn1ZyREYLrD+qz6q4KuLjTTueIIRAH02Jzis4PIYB
cO+QDaby7CD2wE7bOZMBnmo+pexjPeIzYLc9PwWqQoA3025r4/XuhBR9GZI6/BaYKnx2mpccoGZy
OkwLhgBGB0DL7QyZaZ0xOSQ4K0Y8yB0QjRBsdkEsxhpxoTHTSoszY1hu7peCyPivcYSO9SvLQR3D
UcXytLzlG++YGUwibPuWnhz7J7dL89/+JmoEABqTStsTreMKJFiIlo7KRh7kgheBR72mIYvK0KJ6
ubM+9AFs74Sil4JYjdOWIfqd6r59DItebiLUyXBPmWMtWR40HpyVqoneM5645nWdZ6iFp9JA4enp
9QiwBky58aqEv+T9Ci/L0b/R4IG036SOCwsXh350rF1F4wd2OlzFUi0zbHo/2bnKhwRlkCszAxfz
owffbpyGTc/lQQnZ9lTud7c528H5Z+Qg/Aw3QYP+KHD0wMJn9Br2O1qoDXWybuBh80NNSY+2AGLP
CrM4B8VVyoZlxm1zeWBmgFfgSspS+nb+5lG4z26Wm0vM01W41wQGBzdxboOtcotQP3uh4/2NKNbD
vVrGxffp1hTHaG2ez5GuYbgGyPeMye+9Zm/iIMOO2fOce+z+u9BTd6D4omZpBBNVHEasqAyvlnWg
ATIlPA1SDiKGWKiOsZib/mPodD96NS5Sd+EVGt/i7WrTdUrSoBV5ctbYKKS0Y5a5/Yi9TlnO8ZgE
QPtnr8SG43gUU76V7jWpwwXMVTO32PjQUo/UiflloGfaHfIWss+nF29VvH+yuR3+L4j5PjiScXC7
Z2SQRvyvAlubVtwm/y6l2OXA3LgjhV/GOqedYUNZyv3c2Sp4msgsW5UEHAVILb3T4fgVQxJ2x9fg
mtMTFZkJQzDSnakhss0OS98tRaI1oLOnzVBy0D0sWEFaIbjDsbU304v86kKmMItxRggZ9zbOJmQs
udZUds21kfvsyH2/s6XUAORnz+kByWDryTpJSQK5JzrtwnbmJAVzD1b7nA/mBcHqrr6OJWOzcUAT
Yxy/n6vk6Jlna10ppXZKs7YpIn1NACKNPE5w9JMmIm+BROPAVykxxlISQC4jaOU3Hr5rTTgmxJ/e
XXueoOfB8wP2WTYOgP5O3+lRsCluzZh9EEF1hspc5qJ1oZwjKZ2tCG684/eL1/r4T1V7WdWzH1YV
7mBASTanuPIFQcYCNi5TncZCoAv2ELNrMx7/FHyuiGLh+dFvvqA8oqRiuS/dAlyClDVR2JlBsgQp
08ttYnpjLmBj91E5J0+Gk5/IxhC5p2ToPjyIGBUbVJcHfre8JtZYel082Nt4W39G32e6melZCGVi
23WpOADqN2xx09QUaGhm2Am4iOvr1dopaSrqGTaWY5ZN96olMHFOMRVBJgTEyjvck5iczo1VLo8M
9gw4HQ+t0PNCGfRDlFWnvQIOzQhHpqsYrTzqly/IznwItsA22SNuuUkCrXl8nogzbJ6N+15F8V63
tvJYFVMeRcJA+KIPQ6EacT74JbdXDnn0FvrUqs2dQSQN7UCDcYAPq1SdnXFM8liD6cTqWFjABrY+
5uzss9nlyMUtGgYe1H/YFG/1tDsj+JD849AF8qRpDFX12zkuW/WW3JZBMTr21Fi1xX/fY9Dqwh9b
sgtlJnlhw7Rh5xWuC7U2FRO1UO7f5QR8q1uXcvZV0INwWSNNxW2pPhwGspaDPUKWLozfm6Aay3zj
STu0TEdLF7/9f1JZRBaeYgQENd5qRzKiEYwMX4FowlObC/j2IhcWYgpIH2wGX6I5p7Rn3QGE8Gbl
jHCYzC89H13v0lurYCS7ZGTTtLKkihyi1I3D814ajygdN9cNgzOw6CgwwrxBSenyR5IX/qP3/Sf1
BN3MjFe8jX2+O0CI9vj94IjxqXG25/NJOx7HSlDfPojS46SH23XGzMkmWG6Dg8ZxwMg/kfC5SjqH
TNKDJ8IuN382F/2AeZcrNeLAOXa0TP1aMaSa6VqB6+MzOvaOq3PG/o5dZJ49y3xqL54oiFFXFa2I
crZ5B0x6XnZimV8ysKe9ZOyijFLa8DuGtLTvfUWf0v3M9tWudpz44rr8asqKfWEa7+vTCl+WyBm9
C61pG1MI29EV16ng3Z4gbsUvTudGaBgq4WSyJ5vjXAfRqaIEMBLcwn+SxLv8/zrrQLsUUoUVZg86
inQ7HkgMh85mJtA/6yHR17CNOmdV/TpHuGDsoA+LkGho/qTUz3kye/nPpIOu/UcPCcb6BF3k1Xin
j6KeX1C6Luw9Egaf+Z26gZZOyQrq8Wsa/wjPYAvPBHuXltPKuoHPe+2ZVuRnm/CHnRKkrO8i30C9
qFijlVWjXWD+IRsT5mU/LdkOF6+u+R8fMdLP0JuNReXu5KvW/7iYOmH6h7CIh4jX6ZjabPocILSv
Uubvv9g342QULUBLALCXg3FJK6zLlPz1ZqGIjMeebP+DrnLOa3Ccd38U6lQWvEvXql3LR0iW9fhk
jteJ2k3D1ObU+ZC0e7mhl0bedN5WuhN8nlC3t583F6OZv7rkeBiVdPb0aQJ95XQwTfRApIvVwVLK
yyRhimFMKre2cj9hArSpQPOgnrls6UIPfqXbhtVeH8WaPtjUXxNWi5vrw5ZOA/Mvlr+0S15cMynC
PInxGVX0dLjMCAWQsVGjiv+KSAHbze5NY9Z/2Xg/Vbir1FE9yGO5YomJkSbRlxEyx7spMWSm5Y/y
C95zvcdjlDG2EPYU/lYNrCNjhLFK2BT+ReMlYbyYHKGk2ZywNaKPuDm4UkOkIIOWrXtEbp2vQXRP
nKx1TOiJ38D7MhNNhG+eSJ0Qc2XlyKoX3Vb/GvWP5YLSKpyadq7KdiAEOtaniWL7U1P7pvL7vz2q
G0JurWUatOKrz6Oh+9H/E+gv3gdvcS9L9by/WHiccHtEbvPHlEUckgz4NoNcfjthI7AkdpeUeuHH
DNWXyaqro1YBXcPFE4X0/z4bAMOXBE7ecNfF/lnl4tD9+Rfwt0Sj0AcxMcY85BRvDea++swp1UtD
GvCX0bEjBD4vOtsJfpicI5eosugb6bGkgWGny8Zm8pEYt9x9NvFXzIVRTNxs/Vwx4JjGy31aTSsm
HaAqljJjVCnhYrK1/pR/yECPUHOi1vXdjAABHqGfCzHgusKL+tl29NWC9klDzY6IwJVzIvb8OvU/
fNZN7HkhzkuT+w5tl/2gxuJsjV45fpvnsrMAad3MjOvKcvo9ty2dY1Pbl0rBJqNVxS5AYDwQcPnJ
6AnMvMdNDeKla5z1jX8//zLkuAwmhgc9290xXO/EXyace9KW/RlHo5RQnWLxXMKDHmlQc8VfK5uW
Ngah0sV/Ze6UFRUmURM1KSuQrCyttYpVQM8ajYaVqTDxxFDeXCtZBkoUc9ZZgZmVHUGx/zRcMT7a
jcH5XbxgzbNo5aOagWxhzIk6XnVJcXAQRNY/1Qqh22SyNR90nW0CaOu2XpsdWUTAjSrn1ZVI94/L
iMECHPO/hcJTSCEPeJd0BF69qq1aEXEMTIDKWPBH7i45qr/5m66aaSx2TcEgBdc2VvPZpGLDhlGv
2HDOavDXkpUv7H7NG0BWIUXVx309Ine1VxIjbN+1XzqrqAqZAzV6NlYttA2QZ2YN3P26SI7mmH5j
IorZdG263PSpZIFFadn0CimuZlG+jLTbS7T4SpEA+fohW5LLmwPCOxJ45jKbEt2NCchxC9IDQAPz
2Dewe31LqfQdMp1XF4JT2mNxrZkcBnnK6xA4faA8VaLzfL4lNfsj95SIFd9jIqMYWcyJJ6+lLqV7
HEwolVRucfhr05Uh1KwXiSLoaXfdykkdshTjEEBPwPxpWq4p2EXR2aSk1A7cUy96D709TTx7aq2F
S/0UYyE7NxbmYRS9nTXWvd+Fim/m9V+cgPSogqLDOHmUmv8ok83fMGwhwRO35EuHRu4LsCCEOq2X
p3Xocm9Jg7auG4r88iysgLeuse6QHlbkpH+VDiLPV9fvnswjl6JdnHB5QtdD9HsC9yHrJnEiCPqu
NiBXgz/V8R4VSzqVXaF4HcZ6JPeByflkM4nc2p8d5LKQQjpnzlhrKOIlNKaQondtryQFtQCFQFvc
24D/mV/F/OdOgoeOwFXnu/u9kvqiKn8q+ZFlIPxie9Njvx3YV8zSOvXBbBUxXR9l69W7gpvoqihm
E1LE/rwSCUNneenzNEuutVqymFHIxi3UJ1cz1EgjmhXiJzsfbJL8xFfS4hLdYkVkJsyiAcqt8b27
9ng9Dt1UoCgIknuCT2Q7EN5LN4ZvmSmgKf0OX9apxztBvxaZiqBVf3GmGpeAuMIA0v+jyonzUpTs
yTwezJtnNNp7T18XVfyK+QcIu77yntFtOaHYJpi0rwd1Zu46V9YfScJ2k1OPyhLTD/uRBaGv0xyQ
lsfYfbRGtwuZvQvR4Vk7GAlzcA9Pa+V3oyCR16tvtkmxjHwolRs0lknDdOvgdnDoIUKd+KJbnmMn
G4cPBHxp3IhghywEv3RKlXXioSRbtHZQUi0ey0fJQWK+vYrXnPbCexMg8aqMUkvL3R55MxMTvg2N
omLLFPUlHGtY060ucIYEcsU9EJBFvvRdtw9HnPEWS4hQ5zTrM4FDX27Hs+ofgFyeuW8mO/yu3cqo
7ayVDi5bbIHpkxUaC7lPn1nqWwtchMB09JkiiE2eQBmc929WSTM3oCOTtuAhX0y27mu9h1yomAvn
VaxPBNs+6TlFSgPJZcMZxMhUgCfxkWGPXB1DNiDf/vELGPf0tBDxJzJ1rbSNNmYOmO/WgMdKl4uV
CvUoNIEl0errSIkoZ2RM5DLyZ/fT7Y7Qz+rFOO+C3P7MsKpK69jnBvrrKvEz76EDEMCcyvAm6RqN
UsTXm2Xd6CH00RWYhL6JbN1ea9ena2SNYfdNKPyeGt3HzYbsYftV0Z3SLUhqyBHEhFPnVlrHFqz4
EPKP2clH4Jz3LaA3VAbHd++bA5B34Cir8xPkXIdsP0e8XMovJR/0/r7y/ND587oSS7eoApX2TeDm
1n0c9mm5KOknlunJbGrs+nq5yRoT6Nlwnyvr8MuAcfwREPGwkoMghUr5tprG2uM5xtnPflDySCOc
tEWcNc37VylomKrFQu8O2IKmIbePbEw7CwAfwau1amMPVe6PNjJZsf8QjRzmGm9sQzPZmU9d6xh6
R84D1Pbs6SK5QWkV81Afq7bRyQ+OOXWXSeIF4d1q7cHpGgL5EWQDy7lpBQGhwduK8ruXioUBTKiK
OU4KmchfwtDsZD4ikUuYiORmhY7/mccSAyAdSycUbVAtIyB6E6iJY0QZ07o4kNu1/AEBUWrh8cjx
XXvv1bgkfXoyNTHRRXtAeYIdikHHj3TYvVWbFjL1WNQoIOsDIUmMZQSv2V/y8bktgR8lftb6a5TZ
qBwQ4TQuIgMcR0Ejei2UnREFM2itNTlDfGOOqz7gtDQ+LZy9wICLhYzJlH6HMRcpppDBgn0RvJ1z
NAzq6sb6Q8eDHg9lMSLqx4dlxBh5l2W4EwNY3kqqzrWm28N98t8Vzy0b2cBpDli0d8bZuCTA14PQ
cn6STNEZvTnztdTpcu74WC7N9uqqhCtVX5OS8S5MAWByWPjfsssS86K3+PvLL8jOo0FWqSMtXVQ5
TPBYpF590V7uU3z4U0kkYcc5G+EyaZbXr5hBOG2fUBwy1J5EsNwqB6Hu39XNVWLJ4bLmKis9X6uF
rk8aebU6J3M/DYpEVLdAB8kx9b7PNavMpOlYMv9LUs9C71l0l/6UPKEOlqKERPC5r9uYq5KM8gg3
CRLM7iGjmAsGuI2TN4L6CpyIH4lTyamJ/4LSoHyD3bDVGQU0aVP5Qnpe2Q31Huf3vwi/8Fv/K8Ec
a5I6pTcYzM69++vH8rzzIGZE2No831JpoTTzBBph5EKjxHrDm2F2/nB5ucPdt382M2TL0lKR/h+z
kUoBly55rKTllPW26yL0bigQ8bfuG9oqrAkJztNc+bhMipm0dTGYp9dNPyzRj0oOIPqEaWw5e9vB
HJ7pa5kyqygZMpsCpah3DfOetOd3QuvYIv5SxcaxpH/K6dYRjKUWYeViQuVC2/+YunfmDt9RGCVG
MzO/9PcieQXo1mutcp5sdoJGOgmJhKtrm2HdvqCdgnofOwX9W+Vub8ANao6AMCjP43rUJX2CFdI1
GYAj2m51q/uwrpPr0PY67pth7w/BgDNFrnFkuzLnrT8AOYsqSgl4z99Xiv/KU6okw2q77HnFhB2R
5XlmDX2dzzaTKlHGN3sV+V1InkOy83V82qDoMfVLg0/ZKE/o8cJfxriY7ZLa3Wvhb1oqUM1hm4/x
5NsuUT8SnyqkMk4i85vaAJ373oX6KoUtxAZBRk7f/7WwbpRMeaXfZ3BP+aJUuqJtRwVZIF/Zjkln
ToQv8YQXvpeu+YyE2zUBzdbLFRXx6kHR6HdC8QM7qzLqv4XmWTmhmiDzEKIWfYkIzuf8D13b6Iiw
SqBZozzSj5Em1HzPUnYxYDcozXKi8Nh7F1A1kMP61wKy0TPkQ5yS360SKcoRWtW4JbQVNaNTePTv
07G4PoN2L319hK+T3MVfsUxd4jSpNG+WND/D7Onr8K7gF/NTTR8gPqyH07sCisEKWkDtXsv4F2+R
vsxgdITkj3rmjqtrzqgZq9XhT+arOLIoG+dzHu8GrgRKqvRBvpq3jiB5cjhltzzwbcxOYTduf2F/
jNXw9tEwrikGRzqREB565JiejL1MzQYLPfIwwbGteFfi7sZWgnz+MCELVqeS6UmJWlBt5Co447YW
ttsCV5vgBi7EiYrY8yBrFjyLE9p5W+vmQF4w8eytkgLmonJ70612TYn4iMO/43EJd49Gt4xWGm0n
Xqpc8Ykj8qCx+XStCzxA5b5YoFMEDGkIVEwTIS0EbLF1EGOMWBglG0LuG07YTvdmO7FD2GZ6iUOV
x9MLZ0e//sVcCFC218bl6Yj9RRsBML9v54r5gFe1xj25lNrKGfu/tU3UVUja2MCrinwnUQ1aeKhx
abN4G9cPhfPabzEjW4cVe1gsUjVyklNhCFWovX9qpdCpU4VlDRR3w29llRuma4MMsB5ycvgALDBD
lSgcB/MsNpoYrX9k81fXvVhkCrHnnFKI006X3gqngX2LZdVdgNyl7gaL8a6SMv2d1Efp2IZ2u/DD
apKT7Tznv2+IMnlaBO1EViASCxjjH2lsLI9MpTsontsa07Lhpam2X50Rmwjk61k/9atWw4uCuqoJ
NtgX0Cnc47k4KsKGXWWJbO34StRO0JPUZ252Ep9iwopNv4Jia8U1U2eKpRWa96wJMr+ntb51RNc7
BzBShITRXciK/50Fh+V/ei2a9f8wGkRL515Y1CBkOn3a+e9n9Xt6sIwaFY7/b5iD410WBJ0hqPPQ
B5CZd2lgtXjHS6JubnjdAcFCdfU1NSmp/Tl/mQguTNTmrvsZlywp2sq6TumCi6JZznjP3jNUH7RC
zMc7B0T6Y3vTXTWpsxDbTjZc5sMWEbluKOz11FT8N45ggLVYYGePTVrFbl0H2CoGX6xh4Ojpb3e1
jWlj6RIWMDfLkVEypOhtM2fbNJcRGHsEkOt3Llg3MqRox0l6Vbx01RHgx60lfohHJxgaLeTp9OAm
tKGH6mHZkHsbJRVEi5nP60kkNzf3TjSaojgqjEuYt4+U+88yXmlfCg7xRnt/KP+ourCEXqGVNj97
ym0wWXHMmse70p4W44qd1AUUgJ8xzBAl1Z1pxI2Dniydybe2RC1FehkKwLBS0Nb/k2vdohHt19UE
u19j6iCFy+ITDYgkHRckRn4jTOyNRXMWyO/0z/vqfBD3gaxoh+WVFTiAXFohinL/WhstE0MHi+ze
brEIShu45xsxcjEM+D11WkU/9MfqYOpKNqgAiAvBn0chuzDMz22qnqadKMkckYtNFrtNBmPu5Xdb
MU40PXj7Uze8MsFQmxDoHMfp1DAIJqJBbTynLs/THHsku2zNf8QpEZPo/yhGu18Z7u9A/9H6Z4YW
uto38PrZLsbvVlO20VR3xTkxFtpHeQDX88lc+6roX2Wo7LioRMbvQ0ckPgLKjFZA9+XoAnZfirmL
Sll0WAzeamOAJaib8+EK0t6Zqc3wLe4vS7q/gG07L67BIj5kvnP7xAldTVDHEACCw0wiEEI2jmmm
yCiwuKGh+fsemema0VaPV94XoHgG+B4N51YAEjtM3mtSTHJH6pBsvCIQNpE8Z+IpNTgjn8btXK0/
Dn2/J6Koyu3O69RAlGBKEfdGI7GSFjsbST8PClZq+CpUdvCCEa7DrIIfIg9tETOpy203nLh9Ekgj
qYK3QcQ27I3H83dvBuItKJjhP6DifGCN5Dy0NzSRnkI5O8HF0h4K6oxzHVnfHVIyIW2x4bS0k2oa
tU6kWjmaekr/8I426KK3b1rd4dNw51aBJ1bSoPj+fjJstNt8tYl3iMUj5elYSHHzq2qErDl/Vcul
VIA8W/RolPsJ6hwOp4neYABSHyFPPaCPSie1kC47nnf176Vu5H4owJycJe49uu3bKtjnRYlbSSa7
EEZjX0bzTxEmpJ/BhzP9jiXOSNQq9V2SPVUPC2iI8szsUF7ilOrsCwHbBolCWNzYKOBJFwF1hxJF
871TeL53jt0ebcTqyjM0M83ms5NAZaNeOi6TZORP3XpFp7TB2deKOwj2DM0U012hvu8KISo3oULU
8wxr9SUHL7BcAH6NlX1nmgq06GxWHF69j0zwZ+ydKfiT8vJi46gc8GVJLp5StInRUZCcgv8b+zyo
76v8ThMw3WmDPxCen5HiWdM3bX4fpwzj84zgfdhzG5JEzLVJ+pm4FQuA3XXgQfb5hA8z73AOG5Ar
PR7ktD+e9yKbtIrZZgqIM2Xyxu6stPp0ayhMncALT5ZSIN/PcVbF4S76luIGz9HbI03h8wib01df
PJ2iED/qzeoCQ4hcS1nk+2DV8ymkuu6wqMauhU+lvbXyJqLuaa07+0Mq5TOED4b40t+1J2T0F0HT
lyU9TvT5mYKIDukmePLpHgcmBtG+xlOU2JK3TbAshBgW5Lc14qDPOhzrby9KX7vIfI/VC+snfYpy
91jvc5z/1cV7HBgvnIIXsmIj0NllYvXA/E0/fcJPPXEcqu+GryuT6XBiRKgO+uqaJA895fTUiUOn
VDVMOAST8hx6wWNYa4NgSgCoYH2TDeDQgOLDPXIYozMMgsBaGvGaTCvpRhF8tqrd9MRNgjSEOa4l
mgq4Wevu96rtpDUt3Erb53fhmHDCz5bK0l4YxIVKZPZUUlnPm43TNYbVfK9qcGCZpxXcXJfZVdY/
VKzLcd15w6NdRHf3kas1NxwGDUbSO//DD7yCPB/xDgqqFOiUhGZOsotl8LSnVKGlkvoDlHdiyeG8
4f03K2kOqHxAWL2czbgryX41DlzrRCDjqNED14jVCmz1OnhYQykedW1ANgNnQ3jw3mU5SjBQ6Ey0
RYH8DIeYss/Ow0Ok+rUkw3rBMe4vPZI9nx2gnRFZ577yh93vEHvdzZDSbRekSgDLB0Fo5SweIMKU
hpAaqK3GUhh/rN/q0ZwlxqMhMqNnkSP2gsqVTjESg7XneDUjqSsgjPDwsep5mKm2VtjHj4CPNSo8
mZkuHSerDniIvrSOT1x+LD574YJ2vyEpmTRIzQ17797UkDCP12atvQuvu4Rk1b871/Tc+cGqUX/D
rUzdngN/zknPnjckOvM96xP5Vr0iTfENGSSlHziQ1cd4gUvD0AhfoK3AzDWzLc+xi7HX/JKnSxCU
htl7get+GaObgeN39SbopYVzpEVhbKinbnMCdUMvYQQHIzLQKCnAC0VhbC0XzCNZz529WEW7Al84
C+6Cuix5JLAkarA1AgLrSpGPfQmBG1zrbmWW3+0OsQQ8TGy4xvU0UJYas+8OB2d67ODUTl5jsw7d
nzuGURJaSu7eRBjsTVVTD5p4TIGUHXEGAilzrwTlElAnbM3XmtVjK5iWbhW64ke4wu18VmMKvod4
hxJ22tfV4cXRUYrcZRc0aGOuN4CKZtahB6IFbhP96A1lchOSFD+0JFG0dyaH1bncO2RnWwa6Eqz4
nlVWpYvxVv9Uvu4qJmYVKItT8ZFTaQ+WPh7DQnwoPQ3TtWth9b2BnLkyF0Bo/StMtZ8qmrkHDpY7
fo5hTma3wEoxzjgzwXlnDg0xZFzJEZ/b0kkQNmZIl8SBwgxcAr/W5eeLs2aqKhV7EdJPxGaUzNHm
pSKgCWj3eOHIaaGfSjLKoeHJ5Hf6e2L3w1Plo4ylrXT/z7dkbAUJgLNbIDsAh2UnzhZUdBnPbnPn
yVwp+XLlybZOHT9GTwrUQFS121FZi/NlHgyloOJjuVoc8A42+BtpGLplrA5oy7Spp13GJaBinWs7
KG51yEKgGNuECpyb+MABBTXNbjvAMlTrnAhR4LE7b7FABxWsAhnEUA6vO0hkPlfRFktraGqrGMEe
FkH7i7wt837GhoIX0+pYQWj/Hp8lwhhipT96SVifso7cCKWqwKPRLvz1298lk8Z5VQ4/OspNEW/r
vzpTj0C6do8CPs+3OUwXgB7t8QUWUo5IOWp3oB2D1O+FLzZvHmXs3CMtqnJ0qopE0u9ya/pA+gkQ
Jou2e1DrT+dNyAbfr+FU8MRCHxpdIyWSOusCqQkWHpxHCwyKapf5uoixV8O4p3ShzmJMhTc5yJjx
Ce+lf4IaHtsgrkD24RVrjn0quw1PN+nGtTMgGcYHzHRVv9W2p5OieSbEDCpUyZ9/LW/3/b2MaNng
9gaX6xq2eWs2A4u7+Xkyjuw62BnHmM7cRVM5n6j60FAUMT1HX8d+SEUB7eoQp4OVxYdgX7AJL5Kf
uxIPgTu+ulIjdkzKDjxW92SEb+2Jxv9qN5keRR3JmTF9dhvm2TV9ah/r5uc8KC4t6HNanj2jr3wr
DGSgvNmKHoHDlfiLP5C+prX9U1j8ybDJoSzQvowYZAkCGbemaVpGZyaj9I96xHpbDJg8NIP+BawN
1+efLLT4J24nwX4bU6kpXR2lr4i18ctzoXmO7ITKN5lFiLwEQCYWQ68fTGuTvMDZK5Rs2UIJZ1jX
FoSX5ZDwYg8t/7VK7m0O+cDNY0LlHLMT4Pay+s0RKsEidiODi4j6PpP/bSo3q9a2MjS6rMMx5j4a
eRKkdnpRyy1dnXR8tt170rLywgmqv/9hOlh0XOPNyndYVVVL/GBEuzyhPNANG4h5x/Cm8oaB1Z38
Aq48Y993/49kfbxxg6MFnde1rcq7+WrcMwMiND0ia3BQLK4qwPoQ3S5/dyBkc9rQG9X5+h7x+clx
hQZ+O60oMU+mQwDm2IkgqlmWT+kln2l29fnvGEsg+HIFOtQG3JRgSef0ma0JueelHnlXoZv9eBH2
1YMTcGv/qRw4qn/mtYF/B0pbHRvOc6kw2aYQyJburGqS9G2HZJ/Z76v3yxJ7LAwZUFID/n1bv5gE
yXMonty8tI5S3UCQODOjvM0uQy0j2S1q4B9Dso4R70ACriiG1Y5abS28/rtbCNfFjo+/U5BW81Yp
LuiOdsaU3tVSWDOu91WozAD3H4zMQ1UU2dNfbCG2f8VdXP6NEvVrExKxZIXyP4B1MPNnQWVDLJ5L
c5wPB5XWq+i4WWFhu5d/In3e5Zj4bi4RnLyHriEJCdLQRGDHMeQVrxK1Ewd/qHpRO0nzKCD6Kjyu
E2SLs20Lh33iNX5n16xc7teROdsbLPcL2PVENe7tECoyfIZpInYwdIXVGkPq/gL5YtbNQerW6K+r
Oih6N62QimBUa5N9Zvvh8DygIhb4OGfJrlY+nRN3ipfe4o+S2gKiNv+9zm6P4EEWqcXlDMPw6Pfe
KKekUlaPr9l2ewqgrWqSuF1uMSgwKg3vgSTVG2FLouzBDqNjISoyIY1WMZ1mvGnvG2FLlUBSRZpi
R9nAhYTEtlpD91YPJHQW2had7KftO17iia3UfHa2DqpMewed8w/k5VumuiU7DJpidTxOlYzprMJk
S5KSbzDYRSezKrjhkeoyAerSSvy7KTzLFeUDStf5ket/aXFeouiGepi6Pn3cWJefgaQJFyeTP8iK
Xy7y09fBcyF7Ux9+rcy3gzm0SB6JzIw12/ELV+8Nl6eQJIZq4ZnkpwFdlCKeCGZPwiFP8YhHD86w
TPtkyWf8Q6+1ENzbnSuOo5hAi1Clmq3e4HkALQPBaLCUpxlcnYyOKJ5aU8Jy3K+WEdBAVXD9npyB
OwBEkmMF4iZXfYEgHDKPjzyCqmraky1oA5ZqBS+hu18ywkOQwu3MbCv87JtFYuQFS+Y0ba/QenL1
tX5qG30aQFKKOHfLRHW4IWo5qY/YdWO/iews7USx2yFtrQ68LmW6e+MWRVr31JAbDZkfObcJsf0D
uz6umfclvwaQ6VmqHBL43HEvbwMYVXiDZTmLCDVd8LcvE/mytSZ2yzWOR8madJr3mEwGNJIA3Uvj
GVpYgkBWmokPAcJ5Foy1+PbuhrPMBVn8XunS/rB1e5SKQnPXMdUnYyT+FDQMXjNU+rBIBEDmQemy
mmwpd/UZ2O5kCmuQ8MilWjHtIXQpGng3s8YMyPUfRkHx6a+Tk+8L6d15fcvhPfbDmQbcNTrDfVTv
zLPRRKsnf/HJgrR2HeErFLu/kSSX7N9CHLSqKDIxp0ZpwgK9SAKcS5XLcMZo5lHvJoetdUha+WFE
8e+6PT96ON1ZHB2dqTp4X6rELPM8cjAO9wPU2D1lATyF0QF7UuFACXOBAPpHsg0/FI3EwHqxEIjO
Hy6cVxL77gqiIAaaOccyAjlAI36Sx+ZJTcjpDpDY+8kJku762+AMavivzED7uJDT5i+hFE9R1TB/
1M3KJgOnVARisk9RwCcMVil/UVJHUmRfxIilZx5aEBP1zE3gzp+zf1RXkNe10iQgOWa2hU6oOKQN
i146Tz5EC28Gj/i0ceKnyXkUh0YjkYSAx3aJZ08E2/okXUsLYHB4oGdhcBOyD/N8EDw1i+t4T+6a
CuhErAEMQHma8ow7QptulinH7mR02ARq68nBnTiCiFtTfy+6AmJToWNd2xE/ggZvwOOGAUhdoTN2
uyh+7clGQJ/oJx6FDqCzHt1o8mUE98lC2v67JdxB135mryzwsI3+QjyHqkHvVwjoT98fVZJjmLXn
flEk5gcp0F0G1LOTaKrbBwgYPcq7PWgGkFrrqIYzKutkMBKMIqmwf3G0XfoOTJwrCKoE/ZM+R7p3
9bHzIk71YXt+Pz+12f3rRxCXEzvdNiMLpl3oz5rlMNwhw5CnL5Dxc2Ss255WZRvIXpSi3PNYtThS
cP9RZcOPkPj4trIIcMOQSKAfukFRlqbWb2jNSVyef4U0IEN5qHe8eurlbIcrqvY1T5tq58ITe8+N
feTQEVJH9UmdauoyhmwQccRPzBDHvsLcQDPqesjUq67zhBksmC5DP12EF8Ip8G7tgs4VWGSJzJoB
NooXzZGL1WIm5rSI4r2E0GMa/8EjoG0eLJR9pN7WYB5j1Kh5ziADtIyCSVEFx18mYEl+qQ+dkfHE
aMAGMb661xBLFhbbLXeby0lbzeh7L+6s8kbi4H22QzNSBzJeN6MADNQZPiI/9qbp8eA71xIEhyWb
XUcIP5M3sP7newWnPOYKHOnSrCA/IU7J/59S6eK9QN0Hfb7vB8HqjNGR8RLN0jGj4JY2fZyetkD5
FmRRREaMYz6rhd8iadPal7G16InsMCWlLWZTvSF7HbDr2FLyiDUAdQR/iNQFtNhJboE819Dm9Vwm
ABxUK5JI1Ll2KxRcTGDUxJX3LvULeGssanSII2HJ0VR+Ek9tHT97HjhoDn/AJvnixx8uJfdT+B0d
ZJwezMuw18OGVCN6QZIrlyrE1FQFqQs26qIz7k+T0ox0UPAXryGp5G8EJt/WFjigZcQfquub3r6P
AljjY1Uc//e/y+LiDkJIc0RXTvbHiWFv8Y2SNZbkWbOWtTlgq24sn46H2Ah5RKRbssWz++rt7C08
Snl5VTPg0pCjtHRlASwEIEqYGz9I8un/6Z3H+SV8K0hA7+byNLUbhtHar+5W1P/n4kVgeyie4vie
TpIDE+ijN0KsH9ssKVk/0XrHtFia9/KNENa5T+6rH7qudj1KPubTKpJmrXtR+ATtTVGvz0oF2eGi
RBauNeNQL2gKG9dVnJvFTZxe4/1pcEAG4dzfZ9tejsdRJ3vP/ABiu0yDsNoVZG2N+1YY6JEzxlDu
wuDdwaMnGI3fkSmwcJkm2jK8QOxjA22Cv3DG1Ypu1o8R4ofrMULLqFqpgSMflmHbDY7yHk8XGRk6
3Plxc2hbpvRqWlqLoRkEFL3/zkKBldyJ5p7Rwh1b0iZTe6wLZ4bgY/Xp58S4xt4NMYlgYdIRixjZ
3uNFG/0aV645hvgqTcparIR2p+ELCOI6fFIp4xgTimglGu/masYM5TPP2bVeTySwRlrbd7osOUVh
/jnEFN55+lDCZ3ic8zPbBvyoNot0pvKqFOZlUgudTZe5acw6M0YJ///XTHWD6pv3F/E5ZVf3UNyu
kzz5+jBfbQBhPgg/G4Fjd4/znWSUpkaIKHiVS5XeOqZJlLeOD6jsKjL7ERCSg+qDDvkwGda1BZUw
SZDCtXAA91m82xcgg3dIs0KRhSZUddGdudnuFAiQGliye9+bo7KeG+ZPKj6nk/+DWOosXpoofhYY
3+TCw1qfaQbY3PhSHGYCdqIQ6NPyUobRCmg9FvLe+L9vNmm9iAwPplzmhOMsuWdspWc4oLGb7l7k
83hrzw2qf8rHRKY0a2dRnXEJNJ66oZN5xGnX13rg+csn3WMwfDZYwq+TbP3NhjAn0MMVeXJK+nym
4gDPjFEpsvssOC9yNjaCocd0sm7P0wmVBRbhdZ2sGGFRaxXarA9gMlumaVLyurOabv4fISWjpLYh
6XEXn6np2Ar3WVtRczjaJQWQXvgbmC2NAG6RTrqCVF5aZ4brfFzgLY5C+igw+5KEULCxuwSrN0l3
saC9u0VUo1CisVnpIV8+MZ9GPdU+FbFPAKhlWUsyMDvlN0NjMknJFnZIhUnutJsFvt5nRg4ftxQ4
X75wlLN0qAiR2B5P3cwZcmqs0J7F3ztXbXxiH4suii86+FW2RdLWPjbCw6Qhk3fmX3SQUC/nEkr7
hJzTvG9tTzw1MNFWTSHwOBK9HslU3rMHumA8boxiku9rABMN93KBV6YdL+eicqkIuvnukzbnZN5v
HYhXbHAB3tGh5OnWdOemK6+TeLB5N3+7sLs24fxaDlJgmi+W0t6MZTQGzrcayk3xMZ875L03OdYU
v9OdWQVFmhdIlSpDC5zfrhCur3FqkkAfLgc3Jb8eaHMu6OcVH2rxXXs/wup/TpwtQvbsASLzK0Nw
NQh+zsDezhv7TQUup8wcpNePgA3ZBXxPUUYLObndqTOjJqYaQECtaSGcXuQWF6lKwvzRXGIOKyip
6GD9P1+9Z5uymJq5Vxxyta2mF191FTChelOSbWCF2JYb4dH78STeiLRYGa74i4lei+iNHM5gDfPQ
EidgQ4R20tVe7PXf3AxVLOJC9fc3CcItolcAmAzrE86jeK5dpNcGf0YfinEI0emqvx9RmsWxKCdy
Kw5TeSVml2FCqu1Z08zaIC6p9aeWpzduu3bS7lVGukOsZkFFbPwquyhXgY3yCXSVwLBdQ4uVIbw7
n2qBDKbPP8iQhJGgAGsVgdbe7s3KnjjwnTt3Vd5ZJg95k+dfKGcv2RMebFiTCC0jpbGVr77H+kMo
E8SBJXlKmFkuU6sbaZ9gzXXRo0QS1edONiL/LNF4vSCR++g7OXP8bXC8ju5EQB9THZjJ8Z36JA6M
ch1w/HchfrWOwEDsCwrk/U7U7hVTLIZoP8a2kHRhmUC6qVppcsPBUBnslOIL6CSgh4prUqrQiMdn
9LfUFdQS8+XGon/q638OnqWzDmmh0OJ+PeksoxL5WSrxav0Em9jtwIxaRtajTrp+L/sbYFmW8bSn
ziKBnQZvCSqnohCjhOjKVyCygfWsWxNSV/x5gI5++j4dM8vV8uaaYnYnpiKWMMjnSoxJA4cKzuRR
ea7J+MrFwtlkS7atCUTTyF24d4e/PDuF2OnfXXaevvqQMhrHE/K1O4aiGqF8cRqRAG46fL0U9EKl
NJv46RZMqSl3g0VCFhkiLjH2LfSRdk4ZbpHWtZxjWSghhomQhF82JN6TMVFcEWaaEOfmto8vJn/o
RmBraz26CdCnQ4mSEOo9ezCq4CcK/Mgwgl7SOur9SKFNPpVINHu7WHF3HK1CEG4c4VSIrPMGbbKc
h4LV6cBBwKIErqq9q6fg2NRUmBsOdlpCvGnBoXH9xO/Kx/4lLrqjZlcaK/yB6Q845I7+YbBTZdJj
Ug1ePoO9j6FkzT5ahXkg0m1R+invDN8URRoe5ZeeE9K0YiiVUEsT38Ok668R+5cHAUNrxbBiPLfy
DnWb3xwdCLo+jtaioh12lEuEqVZtFTUiZWIA7/HbzVytKPr0tlKBrGGA4LsUAZMLNBzQ0QOCkYfN
N+G7X3pOoDGeZShadHxebmm3/3gLgrDqiLHk1QstSeBfAVdSA407mgxO2n0a64rbBgP+A7wY3dWh
LNH0wP5e4Yi7l4W7znI0iQwEQlobNX0aDZjPdiOkxNF+gjrr6Rgfl26XXsoBs1yoGNPglpHBUF2D
6sY/Tie6IgpgNH27oqSUZROa1+tuolmWLgR2GF5+5gmFPOORFUgClaL6LjwhEzP2xvAf/NEsVF37
MYOxWX+asOMOpzBnhmRocpqfgV26r1dAejwKLxMaLr9du0KDFuyKLN9SqvgDCwMgwBZu6PhyYks2
v1pY8MOp3E3pis/6Tkrfs4APeKRYz949inugwP1p4dyidCxP0Gi24D5TF6RrQUMVtEyoYHhfmAYV
1aFiAnpEZ53mqaiysjmbFFX0IXmUfQUewVw7Laq8fQIZ8CDKM3Xoam0pwZLS2rSJvU9HQylh9qWW
UJU+/UK9s8/CAgUVveli6HTKcBwd8nRxM9eHHLS4oc2oeCz2/oNsXb8WIqPolfhcd/Bsf7UFT6pM
BsZ114qUqT65mOXwEsl6fVCiQHIqTbugVrpnHDZpIu8WRp14uyP91g637KVGsNC8Gjs6DvDD7EqQ
iRPQ22srM7IVrYkrbplowthc5qCs7wMYsCuhMorelmDPcX3ip6QmdoEPxzJma5wDifuldWE80Z3T
BCyE4/3fl34VB2i0g96SoULvoN094+jkatBk6TA2C8M5vxV73I+Uq5V72nzSewZfalO7z8z7CHKg
zXTuBOnmrA+TuY6Gwq8/4q6wR4l0YkzR1TlV0ZUB8ANCgRwUvbfMDQhGGLrtQjcsVRJmyz8MkYCx
fCnWFDJIedy97+2yKxb+h16GBYpJH6SCy3TtCeh/TPhiLPxfVibxEFN3Lw4EPNjNlHIhoSJvd5ri
2ka7gP6GaQIjdWiWzWuZgGwmFMTjYvz4kqnpp8yxwprOh3mAT2tCaNJ27PCIDYb/zvCX2it1Ft4c
rDr0CwpB75D+YDWOGLPxAeTnDSZR4jcOK2F8i3CkV9ULH+0asx/P0oPlgDfVo6oneuoDeue9uBcf
Jj+TVSJySmkSXa9VVXNpwTeqBZaj3WZJKUAwo9UbjsJvb/XNXWKKms375ku25N6T8Bu+ttWcsyWZ
ZNDFnDjoTKMjfVkOF1u1w4Lv7Yzsmkh1UkgP6uK3q/ZxgPJiDkxwNxEQ7kH2P/Z/t5F4XDHs9k8C
hPyUKzCQX8CjVHfTzKIief+Noub7bNlAj7UDMv6GafexDklAh+rKxBX1myWe0L9nWbniSt/sZZ1B
+wKOOqkoRVIGEhqpJd9NHxfS7E9X0J0RbADl4R3eC8yGGl1gaZ8sGq43znyX96OD7lVZyN0btYYT
3eL6puTZKYjv/6mP747Iu4J23k1jN9nJqupnBJl68o0IfsjEUe6vcqUy8Qqz2nKzV32jDW1gXDD3
ztmYb0EKJuzE6sYKZ796A/GQAkktVtNB5i97wVwjgmnTnu1MatGTSwXzYH6Bwct6fbmRYInGc7qi
2BEaV4ASd/CFhXZcnb55gp69Fdb6if9qjfxjhbpKLWc2BIdyxBDOcWZYQqaN4qVhLO+d/jkMxYNq
8KcJKoUu87X73Z8/fIpbRzG44aN6G7LDoGxQbjJGjLovUAOSq8CjhO4srrAob6pVDlFoYLW5pdNV
BdOOd9FOK8NRO6ISyY5hviWV983A5mp2ceRRjo1qHUtmoXDpg5sNsF4QjHY68qwreUiCfs7fMgao
jcc55Sb9Fdw1GgaOZ3LR/D6h7L+HYFRco8lI2JWmAJhrdI4tJjfYRK4GySxKAgpIJlUDFYSzbiwm
pjCRuTlIsouCfZ0a/IKvqxA+41uBDdCDMe65npkanmYur4BwMLAJUPx8z/EMlMHD14FJP5/DB/FX
hMpl4Hd6GRzEyjgNrTH13a9aktG8IQgfDR+k1+EoRjf8b+vSnwgXgAQZ5wPuVO0VSBMLa2U7Iik+
VRjVQj5WMm1M6QndwCLJ/cfvor7cA10+n92N+F2VhHo9X6EkLInEpiEUlOUE84Gp8Ui+n5MRqvm+
BGBl3TW4vMRgbAjWs+EiaH3rpv15fgSNQyg5o0mu2zXMLIxQZu13flKMlJLx5nFROhjVJlMNELE9
TifP+0Kf/WWwrTgz47d201I8u+hDreMrQOBw+KyEI1PrTyU12QmxSMDhJ+2DC/GB7D76lO2n6X2g
Vvo+xZWywe0avu6SFfH9wtNN/iMRIiD5H0yjKTv3sNDkvYHUTVSutMpfXPG0GITLsJqy/fKQ9BcT
myRr+VPiieu/6UAkQ/UYY5ZUyJNZShz1XUmuD03pqFtntru4fA/1knSgwK7NNmv++iEHhQKzaIOP
YBjokb17Ni4MfGnc8nzQDDn3GWq2rX3uWWM+fj9Lgwq4VO/9JPEiw6BeTWQSXmVEuLJ4Dyj1Ilvi
/+upZyuMRSNr5iMB6AA0ovHjBQKKRxY1zcw7EaZmJnld4FdmDMSZhUgiBGqDmR++OwwMwvw+zjMv
ADYzmA6DEQoFobNNfk9lsoRyuol7Knh5WHNmrGicT2FboKFHrGEhygbuAw4qzwHa5I9VifBV1LIk
vegi10HV1dTTSUOJEShVbXAmV/2qG1kNsELk3K1cuyqAUt1vI+9LMAxFQKAI++u1NcTXoQM7DUSt
F0FaadPse60uxKbHoJ4FmyQUbiXQboVlRROhN1kWHMKFFCV8HTLwrJizHbMVXfrOgmC8hFjucpgY
oWtPYuMh2ac8N2YS/BF6FN3yEifTV55fW3PRmKMx6by617T85WwuxRh18VLWeeXhfkNtRXebbGKl
jpPY6EsXiGCyxyp8qWJtB4/HNJVXM/yqwkAkZAQVn4Fdo1a16shYNEOfPrPROdCXNQLLtBWZPChA
PQiD2sHtaaC9Hb8T5rZ3oPXkKkno2WVIq7x5SHEFm2DXjG7KCEE6WYWMJ/52EIU8CjBBl4y1EVlA
mcT3GxKqQ69SG+M08Gv+8/HdKKgRtlRdkzrPh/AvZTRcnzySlI0ddKmonAcNx6F8jcQNR6wcflD8
e83Qi1oYBOb5thFvSo4yWWC4ci7jWSn+0/qGVFLd4azUOSxYDummdC+7638Iv82fdm+1ugmKqn45
8qSpsSXnqPPLGG5i4GcmRUoPtNgrfnKBdbrrZQTpm7yVSKQg3KBfGKvtEsmAPSszQsL42wPDkmPU
nuPspy9+1hMGboHS4VRoKbZb8H9AjtHvi+0BQ5IBxXKWC71sGL0ixbJsbAHi9IVjertnjTANy5uO
1JXKoPoyVtWFCswtr1s410e/lr11L+0uFSOLv675/yMkDiiJRz1CdVCczRe/qU7ZTakkS5wsTH4S
qA4WDMt6flWuZMn2P/QXTlWOPRUE7zD7W38iO0lrmeWta1MCy5V6dhGKy/eKSqmYLdItQovacvha
mrirsyPG7sWtbhYUpciURUeimUkHHw4NZ3LVN0hqKO2q4q/SW6WXLr9L/9nGqEaoz3Wjd6SZQaWK
/6+480pkutMls+hvKO9fmyZ4J6cwRlF9iBoIpS4qfg7nNhhBZS0qyNK5KG5+K9AaxlwT/IM3hfB6
b3Ih5FcrU+g4kSB9bWSsMqlKeMBNJ44kWChlRw/9tYLkFVCPqYcOOawmqrb9w2UEX42btL2esLsb
v6MhcfKekH6UyAMcJmBv2eH3UtL3fQAEphnhVZ9iqfvziDxkuw9LkT/gb5Zr4cJJiFHebZv8DuU8
hlFw9xRhqQtKw0xXGYJExawFcMBI8RzPhOnCP9fo/0GvlIdegLBAFdxGmwj/Txk4Rs7rQJyoCWs1
579EUGAQshIhQKgTAZKir4fxfEbC2tT2cnqTAp3GHIHwQ+LDhDfRXXE45sn6vrEfxkY1kRZ2h+If
WMSDIxUX7bHXgutXk46MtsvfFbj0UXijdR0lE1h9dR5Sazj6bUq84ozYCE5R2+50yHJCIVP5kzNh
ScWBTpI/3YcJS1RX0ASZhMJyhu5x9nMGXq85+3xJ6cRBTVbN9Ai3glbaiTIN0VIoIUu9KKpkgTQ9
S9oQzHogQ4DielflJsmazn55J5kodCEqfuCXgD0fiGDbAFIYqhI4mdqO3MgVQc0ISIhL2A8lBfBU
oPpHummOTVzk9nGp8+Xf8lGXWdYaZp9qGAohSnGwCYoADIgUcxcsW3lw6Diz/Q6G1ghRYwfGa/37
azSVx8XoYyeQVB45zjvLlnLaWJuTn33xLpJe+nDQRgHRt3v5FLZeyj8kP7+o2z80DzjzNAWDFsSP
1u5nSQbpGzbbLg0lrFqFUBh+ggRIlgg0PzDfBxdxs+XxiYy/5C9DUysEotiRaU7e5eOPM+5x/RIV
yDf6qbA7kjFujMF8h8g7miKVjL/cYs7ASsPEaQiDEcnSg4hUisucfT+gtQ//R4WlReBBhfTc39NV
5w6lJuyZfldpbumS5W7w/TGC54HZIOXylw0TvG/WuQwfex2h99G8l1Fo/RJhtyAFWzgh1mC8FPbR
IzvDNhq/m0wvW0L/uJvPvOL79SHcyI1OvdVuKWn493htq6hlxrz87skRtR1vH15pqnuM8wesgCy9
p2toDazz4ONjzcp5LvBxhsb1gqClnLz8qnSLLl7xlHKLMl2w/lPfvz0mIJob7+NftiXNB+PysQuX
JTzLIEsRZtOmsgMG7LCB7skNbJIO+87ISbyE3wa3Si+HAXHOXWzUDWO2ClT8qH5Nn0Ry0+I3FKR0
0VTGZgHRXPdDM6pBBsvCXiM429rPE38UouW+h+nbdBbVciqR6McK43spXf3ic071hr2PwpTilaRi
YCgJTR99Y/U9uXhVnkSIoJvegVioWzOOQJYed0zI3jCbwz35jnngprQ7ilm3SOs3eCzrLHkI8ImP
LeGMg1DTDlSx9slqHwFfw0kLW48Khs3w62EEnrueO77LBE5Gg65s8MbomPYBE87YaPIrIhjh9eZc
vlY30H9JPfPgfCDHFI1nO1smMNaAHdKEtVFdlnrJhOcq3QOApJ4A3UlyKj5+F1Gm5OOOYsRmUPOU
kCl4nxqtlwHNusMrdZgO1DJl+zxDb4C0YIIZ6SYAsOgpG7+757QmC78ghRJS6KCmdc/CuQRTnF8V
FuPWkUuvTXQfuEdksUoszbzYTOPzJtoSpKsNZziBqWDnuugDT9K4pAGlo8yfHAsY6xDwUFmMIx9b
ficcNmBF85KpvMbDh5TiGR0NdzdtIQcDwKIbX4DtS+C/vcRCyFvAJxoCLiD7eQ+PnlJP7U8ARyDJ
sgvkQrowgfm84yt084H/96TFSpmPkM7K5co2IiF1gf/1XFeuctXN4CuYJXrQohUse8vUyTpPU5Cq
Pz7xTM8dJXEB4XwOFcvYVdt1kYewFzgF07VTWumRhYmzL3v3LlTpgdY85Qd1/54+IOjC77ej6Z+M
Mq2SWCSwBRsi7MADErP1PCdKpfzMwtuW4SrzBmr7sYdhESIeGOh0eRmhenvdjHAHB0SrOB81Q0PI
Hm0UZ0uHBwouFrmJA96iF9E7Fg4gAOf0jdYG1anQflJSiuk4Xnvdqzpsk4SIUEeYl6Q14pTcUYdP
OJl0UPgnCpbxfJ/JD7isaVfefTgMqFEEOCK4jBqWpFkjVRhMAXsS2d4NXst/x+hHL9HkttBQg0xi
xGSxMegd6xoMgOmXmFSOcc1ah9LTcMczzQT/Ebg9KM10Xczz952H+1Euoq/SgnUzH/+caO3TC6z0
NFStzOmB9+vQMM80bke31O8YDA4OZwrnD449IwY6BPVt8O57d1a40xR7CFM4x/VyBLeulgZ2nj7Y
QEpBS4WonCoebPfsmH6BrQ5jG+SYpDrbqn12GLwDP2Ie4y5j6p1j3KwTBR3BYqtou3YnD/fqsdxh
qpKul+LHmGBpMw5EazaPGKNDKmBGj3RRgDWZ56RfVk88D5Car/MnPVqtGKDMmTp4kEDMB4GUOXyq
bpxmvPw1YhsfxqE2iauIEahl0bstOB3oX+fY9mT9vX3rFL6v3692mlFclYIHha23iK3S4HYoUVKb
xGMwoeCNSDE8RlvoB6jlD2tPDCwp9NdhZRJy793CaqBBOcmsLUffTWgYOBCZZJE+Rd5EB0IM3zWD
9WzGb+jhaBre01jgIfcXR6baoPZNIJWEoeDgMbfMuSN0f6c/X5ERvSKcZrJBI1PSsFyl48UtQqeh
v62X57w0ru0fSo0fT2Pr07gcxkdcv4ufEPCW1UAWQsh/5T2YPrXG9aF+G2xoCxPlKv3LiQWv8zQI
DbNP8j9Mh2YYElKgyir7tdR8BdjvPc5w9PlFKWmMN15rVMS3uAdZR/P8QZ5UpshVerFVDLYupNgp
VZ2HCuEC1BSge9In0Ks6hE9Ek9ak9FVZt/X4auG9CGddSRelKVTExc/Zu1V84b19qeTtxi+d4SbB
S2mw0GVe7yXziSxuYNjDGdRPzOURkuO+VGJzWfJWUwT/J+lFpMlfdIgbnsYonkmjZVIfPThJ6T60
qj09E4sIKYptbPP5WeT5KADBrjWzd5Y4LF0IL/PJmi+Utvn+ZmlVbu+mtm8N/t0RuVHeYg27mJFt
ub4u8grmYjuRCDez0J0iD/ELucxRQbeOZmrbZeZmobd9Q5NCpmPJWZ6apcLmBrWATe7IbaYE9HMK
97IsW/klodXS36X6EmIn2NtAXxofhBg8uPlfHqT+3EKqyUSqjpRidCD29YeH3P4VxGdvn0sAOEzu
vV7s+ralkTG61GfHl3EGnRgoglBS9+YCBTqKY4DhiTnMCxu7+M/f07sEqihQX0H/t6OFM1AnYNjF
MfHffR0SmSwrid4ZiE0WP5qXZSoFS/uXlQuCpLpP8CnAzdBE5IJTdeSToUeO7nFFHQikHnks5P26
Os/zsLQipNfyaPH3NlQAolIVxhzug2RfTiIgM/RseUqkM4ygaBi9+xaxE9rTL/7NzrPJ0WhEg1FN
wwNf1gHCuO55OtSF/vNR1dqZJ6FXuc4OvctJE3Hs7Noy/8CNq5gKeoHsjWnZ4uKyYKwWHzrzcH87
VNC3I4kvq2vKjwmJZ/uE5xgzXd7QznHSzDNvHKhHkYPgZqX5CsUi5ycDSrFw6IjspIwfbS3MIA4n
MQMAnOFYlPBwbHaRJi8TojWtWMeQTn1IJN7wi4bRmZgVSzDJNXQCbIllhpAiG7QLy6h+1JSbNd2F
Naprpxi6O9GqB9dEft3fNdO6DxVA3+6wHUboDq7oM0L7nbEPtIPsLGzR0KNIJ0CN6+YGlAx4h1X4
/+vex813BFZ2MvuVdRtz9LZUFx7WIU83XvqR73MAUTTD//+ybu9ZdtCk7TCDlNTl1pDMtNzKzCE2
TNDN2BlpLZL2BuXTYo6qsSTBkh63DzYD06CGZhkE4lbUtQbbQ+X6oO1gEX/sVwWQvMgTHlGu+OQV
xuZHQYHUfJgmOSPhLnpuEaFL+ZRzh6BESKbyiLmdgSQT3sjUUZRU/P1OQ4/hT4EoUgjC1HJlRSIt
+qGxM9ArPuXD0aqQibucv539XDmxPzksZ0rmjwbQrZ4eLRt2ImJRl++s3wZsRnzRYlMOoT52Fqva
4NVuCINcp+YcCnbn6GrinrB++Y7zjTfNv24wP0q36CjbuU4VktWwHLezLMb9FVN3bw81C+tYTTud
okkbaxjhjDrPXBEL9W/veA8Eapcj/oL1dG9r2j5jmeKFFXzw02PKXMNVzwtNf3zuRsSGYyNAOicK
wSpQ6PCqTdXlN2J6hDkrTVgNiWO2Bqxa4PRb6hNAa0TDe7unu3EGo6SvDizkXPeJ1pbzFwAlqkJM
vP5ApSqVoxJyoL9ukIdZC3yaFpUOa4HMalk9upAILCL6cOyK31kllxJl2Z93+uiuTeSBoHnZyVED
haEM/EkbprXw6MyfV55qnQAeuwKu9Zjrnz/iy5LSXeKL1qNoQmZEhRhXjzwh83uIW3FrtJzk/Fo9
rgCeN45U4Tsk6GwLa2kIPhBjZAsNA24mbtWt/5sWy04UN5dJwwLh0JfQB3bLqucRSTKdtTpiDIXq
9aPcX9/CsRLE/pqgTlfY24NwXwsnsdUVIKFhARYy7VpGu31KWOz/yVuEUgoT5t5QMScetVDApLgG
LZatPZdQUxsbpd6n97aoSc7PCyU+/sDBPSjD9CBH4Juxeuo515eud3QWdY2Zabk7tWJek9GnbqX/
7j50bl9yeQ7WUBdWONgUxFAO5Dg6CrxLrMDkkLv4HGNllvrv4+grgEA8ucgMs4zs4W9O8vLuqgpO
4vsa9XUHUF6Zj86f8EsGzJVNLxYoWMvijgfohQosuiLbCNwHo44rDgLflfftbW28fadJ9pzaoSvJ
tCMT3L6P/g4RtOVbyb3m1wPDs1KLLYYcjhegRt6FWxsSgf4hI5xRLF0xbK8oZOkocaPIt5wAhQwq
5/hMgXo5RMIHtjoAfYji/X8oEXviyggEprs251lGcque6u0CWd0omuaDLJSkcIi4YXlyJzMig7Ie
5jgHDI+o8+lWKJ3MSjrrvD6YJHzBRoxne0hr/Xm2B7lNQiDdckUzrlneWmIFLQtoPzsH9KDwQsNN
ZTDhlBXEVyLS5CBC/4+OA08zloZRMNRGMVxyg+/H6U3v+p6vdVnZhxrNOWKLsRlG4f99GBLuEQtE
AbTzNLq/Gly/aBfP4eBxVVEMoZiusxCL4AM/pefzdYSrJ9lR9h2VcFaCArTYKj+9EA1ZX8hOUyN9
SoSlpPYEtA4GCgqCI6y9ZFIW1o1SYGVRRiHQURENtENjuVJLNFHaC1oGgeoNy1MyobfrsXEAqGJX
InLPWW1nJxzifE0lBYklPAMfVNyuoj48FBIUZF2RliT/y2z9ztjtOajUtfHEUeTDdovMLaGVp+hN
2Ff41sL5VB3/iFlm2Ig80WD7lKa0VssyqEl2C13PRrVYwhDWZwJ8jvOQ6i2kzEH0xGnfSf8Jh/xJ
Q/jdMIeEBvpLkCOwALMjXBhCEO2f73LFfTAFc4JREWPpbf9Ia2+OhvwPUUvjo+TLexncPDhL4boZ
Q/2r04nzdn1IruD96iokSEYq+uPaNn/Cnhb6/OIxjEAdnhFbh1vf2j8RCwIxprtRnhZHcvYJTQze
vihfgTIhoYHeBctQnb/jd2qwA9MnlDGZ7la+JmIZK3X54zLr2CbfbvxVc3yQSXpcxSpdIs3QnabU
UO39O25QFkjFaGCaQdGuGqBSinlobcYw9T0S/0BR0bqUZP2NbZa2e5FEZrxK+qUrrdKIBK2VkZ1+
h0ClvenEo06yIYAHNN8l2jgswvzxIVnYlNTqJNHU49oJonxXrAVxWlVVpGTC+9eW6+nuHra/WPBJ
GHJhXK2hIeo/dBp3iwmiM5D1uvm5sXC73impA15yW+XLfGyNyGlTbFOzs8hjpnEuTOEi0u61dzdf
8D68cHQ8XtJKTJiwSjPAjWUTzj6UM4OjVP0XgLP+3fUV6g7wO5tBRxRDP+Ndy7W5xOXFEnsZkD33
avsAPGBst4AxQxkxy8MAFfCTaPpDmqjxhpAjLvWyavzV2chVvCw38supVcuxOVtssPdpGSoQI+rQ
IOaOxLeYY2x/vsfR0WQ018PI1G/a32DAd9wuv+Ii4Al+xKjca6gfbgYD6Bw1fngmpF5ZRFCKxREO
HRZTHjoVsH8SCn8e/lgSkOLy1Vu9zK3nD/AswmeUGWm2KDC4beHqf/escGloutlrV1jmpqMb2jXi
RuEIn/CWzbxrHZCTmV/S853ifqvT1Y56WvIOoNtcLdI3TZMZrWTLEvSsUnhNr5vD7UxwcA1HVKdV
mr2pIKNJpeXJ+FfcAeLfevkICgHTfD+iB13W/TRp/ww8QDZUYzfBJzPO14EQedWyqgNkwgB9zaPb
nh8HNMiGwOHDYJNcodSHAa3XuiioHBgxIdXzCr79JOL4G6eo4IdiXyhxY8Z+T0Mx79Z54Ve6kISm
DCJkm2ZX6DcrEt7ajw5SaQPMZgInp8eSc8nGWCJNu5v3T20n77ftz/OviBOlR+ksqx/pune9re3H
t5TonS+KzuHEXlL3SsWMOEK/alAauzZaLHdKNf87oSiHKc6Z61LGXt9ghRAkpP4TvUfyqKQ40xeU
bnwE3Xi9A3M5ZhjnBNoST16kNCGpMYi3FW2mlGHJU6GWE36F/VI6b7Fn3r1lTUShi2SfnVyo5MhZ
Cqyfqd8NS5LJipE8SAI1XK/6/S6HPqHNwq9Grhuc+iuawOL0wKDmGqn3VUtl+ISp65iZBnfdnGIn
26AF8BhcZM94wzAkBK64gmBLwyo7zX95lqQTqQNSQajFYBSoauwoGPCRHeR6pLypMK0A5CTdTDRF
DvluVcr27Z9NVkCYKYeXMptfQSfWJOBfapJTqV7+l7z+oaGozpnui0CprO40FUPBgDzCuSzCIH/p
dPYSfr9QJyF63XpFHHlyQia2l9vG16aJ5/JskhLn3LCp8kNMgkV+IzRlCljYuqw1rqUC6S4aPXRT
Drs4Zzd3R4X8LrYla5xqvOybkJyNSlKn/2ouCPr+yADFfjWfKMEaRY5YwvyZ45dYjSB/j1/FHPib
8AxMMr3tAO3LjaWgN6pgCy88yzAuFEAu4YRs/gUhYnZrW3Buk3iEd6w3a1GN0fTf5mDNZ0DcbYEu
bK+0k90kzrSjgyL6StfOiNAPmWnNCKNIl+3sEP7xHOmQVNr3O3XpsJFYp9v6t+LBGEkLoxEalQMw
RC3updy1Cg2ZCOdtGQYVpPf/Wq0zD9K4ItufaLhLfrlF/vBiRh7KI5fEl+8+rdIWZyIomeqPg/15
Ad9cL/EyrsYlDeVcrSQgv5xvI7ayu286MN0LVg2hfRatBtHsYuA63UtKEphdT2eYhyJQcZocBKgr
mB0qGNY5PZV8CZInOvcQ2QlrrpLBAjNsmfvwkVK+VFeRx1kh50SRwyF+LgbNKUgv7DUSDecUoam5
frsGmv9+CvhXH9qR1XAbaWB8tjwYUgLkzPZnwMW637d06gCXAjG4i+4z/ecjezRmFLp3N+Xb8i1v
9GcsgiTrbMX3BzkdXqODjaudiHptaX4F0E/fSzObTejPghNjRSA+08VOZ6Jee1wKpQLAoBj8j1K6
MXZIPeFkzxhuU5/Zij50cG9wz3e/NDCr2e8TYgAU4UBTgfo4fcbWborCFuHJZLLAYkFeHwE7kcDI
Ms66n3H0vKilcT/XQjWCvKDysMGxZ3UORNN7zR9Rd4rxBwDYdCGHxSwXAXYS89ZUAJ+XA44+rj8q
NmLC3EEiWU6F6ORtAm7wqTUEdPZWqfurHLLO4hFuNfXz6gmzGWJy7eFGgTMax4E52auvtKk85P6r
xSQBfWmivvAsf4hEsksCNQd0Rl5oSCSiGbBL29bqxmzUSpG4Jdt31Nsn/DddTMKxBg8CrbCs4k9S
olsGWmC9h9cqViQ7ATc0KtFIt+m5dSpWWIYuYvEMV8SuxF0lvihIzyTdSh1em09k9/JjPrdK5OD2
eZ4WPXEnqF9VzBrJBLEwUQtAgdiv22/j36JwlRrsigvyG2notYM1KqOtxY5RusrL6BilogUMHBZ7
UISATpNHSidX7rsVWlOdnueq2Nc9rpG3RAfBtXVDsNv4Bw9wSYdr/KF6drQh2J4dOKEy/TBY0Eb+
aEeWtAeiLDoV6P5nuTkkxvgxchhGd/ec+6bnLDyOliRqZ2WEwnewJ87MDCsxLkZIcaNuOByRSKos
R5z0ZrhvZERpyLcG3PYcboxwYj+fRw4U3EezVilphcvoNRHdPzjuOizxJ2h0yMtdNWhu+lj+Mag1
iYKGQ++0/m2ybfUCahkWMYvgfRWnSLkDRbUOssZZ21XeScXiVPvUofpojGP6vWO2yKtpkvgymnb6
MCWPSNavTTwh/e2fo/RbSkky6VyjtkIPAoZASyUM0x8d1arPtBDQyZMH6XZI8FdtSsU1RydbcHid
Krp5UNN8549f4XmmvaLmOVZ9uN1Em1vzd49k9K4prlLHdr0eXhzHDMdoYJSwNnNF6C17GntwBqL1
57rLozod5lQ1hb31NLIiQWicKXVOi4QqB00/TcAYcfzz5ips4DiQVtMYa2Kypvz4Ofrp2n6kt3/q
AnDUncpgRwjuOYhwxKxH7IGI1maoMavTBw9PxpWXcamidemo73N24cHOg+dF6ZGaS7NggplrQabO
iNZgJVpQin5sYdBWC+EWYwiscuvdLMbo9YHF4al9xQRZVcZzjw+6VodCZYlvf1oeDYqOw9rP6uAr
0m7tzuqAgxaQjX1CmL+cmgYLZ0JltF8aiL5Bs9hG8sduGBJZJnkHeK6+T3c6FRM5RBSCszFx5n0p
LYNc4tvgK/EeOwOXUyldghdHYGcjzO96qEOiw5jlcIrSV+v3ytLL5tXv98cn/QF7CUIdY0hfjGq3
7V4L2zh9sE1EYaZQLnJQ7BZG+VzLvCrU4llKeWVyi4ESzwOjYvtN04/jj1IrbKG+GnSnvLrNHPf9
HkkEehtHXk7jZTqiyeD4D2jjjzVTr90sfsrB3UKlTDyEao81F69LPzaa5m7mQTIOwj3PwhfN0OXg
9c5k3Di9Saoyc29lUI+cBSkkem9agE1PqsDvKwoCjvPU/a3eUfX5Kx5NA30wXjQk5h8p3NmIpTI7
KiUEv+tN1fUps1MEo96/mxi1Km4LqaQm+sSw1aXa743F4b+vNIVdpPWibdpZnw2YMRrK4TANkY29
5MClCoPkM7SEWasygupPZTZCZUtE4eMLYqZYGiRTRASOPjEuc5GMmXX5sXWiKMpT1k4J38hu0Qm9
5yu0LMLjZn5Mk2oRZCAAiGJ8IhZzJCj8mEzDPZTFkSfkF5yM67C/PvTBCHT01KFdreQSOc0G6/dp
T1DOoY2Gdou/ZduhYuQp9igAdGwOu7PCCcqxZteR7UkPVAinmFs7UVGUuZbrtrypSli7jKCevUyK
rS0rwreNsF9K/HZUBE2ZgquQop2me+zbt/LtlBzvSDIyiJJjaQApAmRGnCExgOc/vmHNb5p3vEbz
506j3W6HyFIg4D2VCKWBWik61kWvY0mOghPhME1L62HdIDEVkESs4h0WIEQUveBFyaVBh48LETP+
QavQP3iH6wZvITA872l8VDvQ8yJcnp/+5Iimee75cU4m2yiHaFOEDRiz+LZpNbf8a/7iV0032e1x
3m/5bVVfdc8WoGQpcsqxcsYv/2eIhBY0GiaYp92GqaLOWNtRUe2wh/kLj08yOw+vX8N3r4BfcYS2
kwjIiMYy4fvlReGEGti/Zl60Txr53gD53WJnLfrO4ZxLsVDZQLzkMnnKShYjKSao01yz/jU9g0/3
OYOlgyFKQ6HOTOzdYEJBi890frwA07Qx/inPpy8CCVyu6p1GAZ7yOmLT/Oo2tPPk+rE3KrXowNrJ
5goJEFmEZMTEaCtyiZi/EyOGAY9R9PZZ/wuIje55DfGqfO2SrPy+YSS+ls6MUNW3J6FGqpNnywJi
L//foQpe9fA6EfcRZ9xCAyTD7PHVm75/9ocEUqvweP6mP1CzQozUaKBu+RU6omwz2Im9bDuqIGYE
4q8w2QOeT/lpj4O/DZfhA2Ls/M9BSBn7SjiBuusw4/LMCAdw5dDH/rnDQmKiaWvTdeSzgljTkHvL
e9zKdMp5tM29KqeBKQO0iimUv77O9lQcK1ZkkI5rRSaVFnpTtjzIzL3lyI8aXVofLXoXN8IGNoRg
cIPciyeOPlcsOZNQlllP7NMVA98dm/lBjQg7LQTIBFTBwc3lFWMJ2kkchtX+QNrVbZLeaEnfHIjL
ZLasUohjcUMQ5jTqvREIdzYWNLTmSZF2WNPSo4QYTosG87LySEgRzihxZYkdFcyTXjI53JgHCUKN
U+LhE7THPZIFnndSje7sssjxb/tOnpxYRe37PcogOcOrylVOldV4Ei4ag7Zjgl1uH5Cw+RbUuyY7
WqF9OPeZkLH1y4cyNYUwDAjXKw5JGIA1OCE5VTpaoS45H5Ivr5DN4vqbBVe9ShamneHjkUyAf1zX
aPyHyethuHxyW4uMI/wssG7TgheipWny0eujYmF+3M+aIT6Jhxtw7RS+thdmMzY69iXntXFY5VIw
ICzkhAcW98S3BwbE7XEiwIiRunp6G4758qHUm+SuzOhyRRLes81r/3yBhsNDZP+pZzn/5Dr7i2dm
9qg2j+c8mUcku6esUqYPzQjmzDAwA55oh5albYC+BwSGM+9BsAXXZaUK18Tajt6ZB+i5Ly0vEkCb
sPnyvksKDsPWxRWExp5OyHiD2HM5V602r9LzvLqoSUUOG/Qy/JPKgp3fD9mi8DRSgY1RF2bYAimN
ggD72+1oU7oevD3vnfJV+3pGs2o3LTws57GrfQsNYnItHMckxZ9BEpQ3vWoLgm6DIwvPHj0rcc0X
nNJXW93BtsF3tGwS+fXOhcTw64BAyC9kop3cKancaDsyT12F9OSessHUByucVQKHZeV09fFeGyLP
WGkoArJ65K8qxif/ndV3ExrSoCFZT0EG4vHDa+b6FCU1p3F0uSHCp+yqIMyQhcK9O8zVslvs7gj0
KRXN4c/d4fwp0mSttANVGKcmmvY6p3mN/PWrONcc2lmTe3scS8+9Kxa6WPXkLTharkEWMwrmB9FQ
7vpjuQ183FAANi5hltOBs7HoJBa9Ykt6lX0gyBPGtAYUDRZ3RcD5qJP1V00NUvf6ak6h0sKKoEqb
jUm+9O+qA14VMOimo88fKvEu3IQq46bo9G1h7qCgRR2d84VbcSHf+W8Ki1Q1+MRL2MDbK9opRY6y
fTSfYvlaAfit0vKlig5aMdIndL6YPweFU3G/lMlmKgRTbH980F2vYDl6wXLKmY5KRi85NA1ppJat
lfPEL8ApNdw3Ue6oaGWR4AHH/cRBBgFdX+GJAZD2YynqYvDt1ep5E18cimvN/dN7yZLUNsdZ2G91
yt0FLiNKVcEw/OL//t4Bo8ALkWkyZDrDdmkgSYg2QwJ3iOpjMAVPBxq3DCEV9YWGUKfDSEAUqI0D
t47Vt2Qzn//MG07pDPYaOBHO510wvsBUXHhg0GVR2wDwXGPR3CQ+BqWlfTm7S2eQ/gxuknsQ3kPg
Q7eYyziF2Bp7rtUv13RGYDhOWz+SBXTKmjuQ5XHZld7Uo7xFA6sYSFWLPCUT9/pSY9gOWkfllQPe
fFmRjVWRTPPaI/cq/gMvCocD/C6SMyUBcw8AEOT+cnaM/AR/byz0yYg99zHgGGtH+CgKi8aZp2WI
PBUJQJucA06/1uBJ72zQJhJCV5vnQ+M5UtK9vb6kpYDJtouTRPEKuxOB76jS4CoObfu2vGSImc6i
RaOK4agWQIasYemwVs3UWQW9KTFP5ZivjjxmEDo4pOfWVOy8bU/2Sls31v3x6f5yEBR+MHmDJUqs
JkB+Uhu8rCN9Ckj/fLdPP55feOh8eBcyJ0zRLqGk8m7IID9q9j8jYZ3CZaFQTviqPKghwF+ienmy
FM+PipAZclkrpolL/tYHduNH/1jWYZJUnz7bUEvHtSxf82bIiKwwt8sxQiHQ/rKU4WxTU/gzn6/0
uJkuz6W9j0OLDp61ZjLYITbRDdJUiuVD8piHkHOR8sR68PsveucTnP5idGrmLtxajMYTkNpZlin8
YJkKNTIYXaLoagtg92JWqX/ed92sstTQYuAL290mqm8ZxKnpjuppXWTgtxDkvB4X3ZkEY2TWsh6c
02TSkd1MmfIwOvgPRX/lMnukeSIDtK4ivDxSlmB6Hs5hshQssok+Gc1psejGeBunkM2yEjvrsg1v
JPe6v4cd8aoc3BKNxyDsBcUHkoDubBnHa8TpwWVcPTlVGixynJp7LkSzw9z3lHPodD+sdIJygZdb
auPneRn1LCBweOdfPfv+zoix5ElF51JvNDVgZH7srv/BpSPoB9MtugTvQuRLVJul+iWFWh79e2/7
O+rw265Ov9cZslzOWx3iJCM5c6dWtltA8NX1xuTgvnQVPJbRmvasN02CsQW+FELCpPv5R0arRqo9
OoBBr1oz/962sUTVyvljwh8Tvlu0AfN8Mbyz76KiAcGGeV9g+9t7RPVh/AKtZL/WPnVImTn6SNue
L8Rzeg1eA/MZqT3hlcriBdfhtpp+wRbzpAWPnuypQ7OqSGMM9RUiUkpNnAVS3KNX1r1fp24e0BRE
Yzfyh1M7gHp/OL1FiIp8GtlSp9llfH43QEMY0VCT48XkmGKXzTNa4jeFrivL0CRY5WePnhzi5/qG
9poiJ7LIFXf3/PZe1VIyx5sASb6TrimPFK3Je9Ma4n//9qFxAKBe5MMVxmOpAcDlNn76g06nlyvK
ZD6qz8sg2kFlqIovWJM8eSlKa8l5d+IPKGqC78jYW2EiuvDRC800KQxorYA9yNuGEdd60N6UJmx3
NQlywVrtlodi/BwjeOEb9rNqXbyvyqlIfy6aVCiuEi13RLns5IpJaqFUoYIYp8SQO1p6G9+QzDFJ
mxrFveB0Ac+9fpqQN4E0h2XrP7bRGyyuQUtF8pPkvbDcmjrhxGNYKYac3INpnd/pqnBfrQoTT76C
MfAma9xZTxEyRR9SqNFNBE7e4ocsE79Ef2amOM/vsgmwqrRSiWkeg1SeMkSro62wosVJ4KqK3oPf
RytqVgM+95DaLXVc/1q1vIJ/69fGeCNzueeeNP44wKXAxlybjyAjFXTETGmrPBQeuR2Pi65D01h/
ZHIM781I9SZOiY2PXlgXeao3DkbkfL/c8qwu7y1dTDriVtAakpw/ZoH47z1p3R12vudKRxnac8kk
r5pBtZfYQz7Iu4VUjkiJ47CGOlX9z2aqArbqkZWiOUdwV2xMxQIKBXdJloGpudY9TVW7eTmpxYq6
FXqdzJ8nr6IL4NwzJHkiEF3v0sii2Hl51Z90uKe8+4yRRaq4XreAgTiMMNs6ysks8xocKU/JeyGa
+zjJDCn7tSiQbLbhk1io19ffETZo4Jiv1A4bjimzQnw9kfydLDO08ZZdJJbr6T/du3bXwynxZrc9
MOVyPuXJSX3nLpXXut4s8twMKghjpm56KkAMTM2OslClQJt5Y+sy/uDARSEbrD9wzIIkb8tTAsqp
KQe3a3EPjFYdjjzf2ik+AUuPniisStjTli7a/Ix2YB5Jco/dssngHjTXGg5izR+FhGWorKTlMcE+
gxSSxY6MKGRfXczBaVcdryiwI9cBxEsHKynaqO91xEYMU629J6/IoYr43exvXKH6O4pYu1n0gA7o
Y3EFH6++EBKBujdy0GTzcJoX8ykk1mKdwhdF4HiO/8rv7C3VyQvaPgYVyh2RUsZcrhGZyqE9AcXv
QaYUsdS4wu+EUW7YHfWv9lxINPxZP/9DJM4Tm0j1oQXYgM+QcvODyyhlPTUfS7SjsCWF39v3607q
Iunk1Sb3XnRskiZVHCb/STiesZDcM/M5ZelpljwmsiTUQ2YMCpzgHLhez/uSP1J+AUku1VhYH1UT
U2ugjiZyN5aUTCDQvRiqA6IAmh9WwAtZzXhRo656C/gFQG/7vEA0y9TEhia39gC9KCxpJpH+8ZIS
fzhw+xjihqksM8Vg6UdBj7ESW6YXDDtGZ4fdTgJX9FXULWLzVIC3SVV6p/+wAhG7DuGk+siRD2Tg
wv6tQSBT5se2JjJh9lY4XQYL1/5Hgw5q98CKKnQPi9gIEb/dRwHpn5LOpXXh2mhSBAGXuiyeKuvy
f+2ixEfRxyg7mRbkQOddV1fJUju3ls8KS8rMPhB4ERfvNlX518IVAf1Ir5ZPXhccBc2ScUr7DqDq
aya1r2D+b0uMPWH2wggG1tFc0DwgIvuNquLufrvw4k7OYFZ3M/jbwJz6lWxnjPupTKbr88IeLdWz
2inqROm3F37/8FxORoYtvab061YPcCNPU0CxQP+GMbz1kmpc08jlbRgF6yK7n472v7o6NZT4M0B3
PJeDeSBbtz4Xu/0tBVevLDnnO7Id/MYURE5dRaZaDdGKETFbQFRv8DH6hnoF2A40E1ANZhJgZ8O3
A8d7BnetR9CIxBv8+Krj0yk/Dsoz/OAEVJh/ECoSXsrZdVqRkCCrkUfeOF7gmmQ/UwIM0sNVN0U5
kvZtDkkQXfni3xVmBNfVCrdhvZjpC25junBPUzt6wfGOCL1MBO/Qcgd3py1bGFQWnZRRMUTSOQuz
ZeMp6ml/gRWQFbGCt7qL9NZn4ox+N70s6onDIqFMlhQmhaZutDlYZNpcJ1HQuulB0cn/42jFOJzR
EpoeTgkwGITIjZOUVNHhlTXPpiabVpjJKHmwTsoNOR+axz4VXhcPKEBDSrJhkoc/X9bhwRRrWlIv
jdci8Bkg8+BYdOt6RvyYA+IBTqeWgRcbgaXgOJDiJVQte64+uYqxm8ErmWW/QEvqE1Go1HkljkYd
tBiDVsUpySFEu8GyHJUeR3WmbJUs2S7BcOtksKUpvslfleFs0dPLOX/0Y6lg1kJKQzlayqZJWEOl
dPbapi8t1uPCgmpBOoC1zSqyQLzAe9w2g/z50eP/9xjIzp5TdNAAeO9DMsctolN+Ix6k90FQ7GWC
ntywwTaByVAXnE5wRcfScT2nXn8luvV1y2vGpSNzfUXyhhLjBVarrf7M9MbpojyJoHG96mb6p//U
R4mJXGm/1rb0KdHW+HkpJGTgvUM3nTXqvtakHaQMg+wQCZ9e4QvH8tDDMABqb8PvgWio4yjtGUjY
k6IdR6OxbqKygczR8HwIVvqS8MchGod7nXwR+wXpBFracCeudF/Y2Z7QnHf4kJ95IyNqL2yiEQlg
xZ5yL2fdbsaLWD60t3S8jGgGg+mrI1m1pXhzN1isirsjYc8CvMMT8UwNvO7Iw1Iz4UWQFGYZpRml
iSvqWODcsQmUPbw7ouLAR7S+C/QxMclBNIsjP63J3qS7SpnpSZrrCqDTOTTwPGR0CXl6COTKz/qC
6/Dr8ccWOSDYN4MbafZ8ELAfl31u3tudddP0GEn78+6tF4KmgM0oN/DVDO6HPTtml7qlVYwzCB82
/ADfOqy/kL2phtbJd2UivSowvk/PabOo6x4TrOOQ8qP5oX0xSAMFQjz9qmUjL9v+y9alN4eo4u+i
alU9LIIcJ1dI7HoNEL+XsDOiD355H7cdYBy1kUjG4CNXUF4ex1boEZ0Ths5uZe6jW12CeZuWDPRx
3GQCYKBvNyIThsBIcKuC1zrnUru9X+3RojdW9uQCwma+AL+KgOPOsJQRor0ikbUYR+oawnueKoTO
ey+FDgPH3D1PHwut3THB6L3Vu5OHsQVcFKqaeQcXoR/lO6HImAgY5aciZQKYHPIKLBN0fCLIMWbr
Kg/wRhuRzjRYvHpbe1FrMrEx5xCatxR/uPEQNis6UeFk50Kj1Jo4ZrAKFGdbTAUNQsbX9abaBWRY
oUpcD7QA9uRRhXhxR051SArqfMKpiOfuU3TlYbwm81dNY8P98dip5u7VLn/yOHv9/KJdeUQtBZBq
zKf0il718+omqGra3JQI2wGopB0xd+iXZQcmu3sUiSQvWxzZu9iRgULn2f0qGCbEirOiB8yGQjRj
P2K8SMnzUaYHZesxhAgDY1eY0WmYMMEVoDMRCLODB+lueysqJmVirKO2bFn+fIbq07JhgJzzcJfT
mXt6frDN1Wf2Ph2Yr+l3AbYPD3gIpL1hAYyVhtr/vCXG+KQrXHN7Hmu6YRldc6/JoCz5Oe5DvHFh
0zaXDZsAFtFnEAdSh/zV41h+In+V5qsGhZvxaUFkbyDbGn/rHQElhMsRYu3ZKWSwJiVDPrbEOLSF
2wYWnJhvLYIj7a8MU625wCX5AI5kKG9pwWLTwHu5UKEyzjZewahQQ82H79FhSy5tIxlhTc8aruNy
RDC7zLBcm6WUeG8+QeKkZHnpQxtxrGFshXGXaE3ZOfFd7kwfk85lYUq9B9EOq4Q8XtFiiHn6Ozaj
QOf7mBiHxhsu58J9CUWJxUTvy/fp8fThulwFz0kDIpeA1j4T9IomuSJghI+cu7YU/CNfFszRmdbw
qm6oyELkacsFWHgeKg9ZiL7V5FkFqwMd1M3bPKsu/zt+Fy9kNveR4YdqT5pCLfPgSKPNn0sSJP88
gj+jMKm//U10noCLbmJRPKQdOnIbtQMomlSfkhrh/EIypjXzzCPeiRXFuztaazTx58/LH+Mqfy5k
NyjsiOFRWXxPWeIhcn5iqRjtaDNh5HUey2MgFcINPnh/5wsiahyyJN5JQrea8BNCkikjDpFJC/nc
M+LGVsxbx8NqiBDLf3kv6skC/aVv1KbbgaJLbQnwPBN8cUk2o3vKr/0XAmATlAEwHGzUKCOe4cnj
D1C9BysiTGBNmZUx9VNC9AL4LF4B7xedovnDnZa5iybBYzSK4HMIFuVxAok8o/FGXTgsSSXCcx/J
YVPAbJlKRVSd9NsiZxM7DSQOrsFD+ZpPH2PqEBec4YUbWZXsRTDCQM/fFGUSH84IC5UT6eOk1nU6
gS5RV7V4U376QfwuBDhnEI1myycD5ruJWwn9QPsnDMxXR5Sib0/DlYtLt77Q/zmycQCte8pqqbqQ
ot+DM6bW508lbab9NPlJRANg0lIJ0ucT2yrKGnpV9aWNHJ6GkGGedOVwkSfMdtkvEdq+e54nTLNv
SnmNXC4DdSOdhg2wj9uqrx8lR9PBgAg05oLlAUYqzmZHsyHRHgivc1UqIQON8Q479fPW9EZHKvYk
wf3BcO+r6JQKErYkATIrJCXEWB+XGIhHPwxjcB/DVJgSOmTm0jn+e8V41ZOSNrZop1FDIWl+KlVm
KHRvm3xAPOvX7LEKwdHPuwam6zP0Dfc+hKt2+nT+1+/73WYRzO9QSUwnucid7Ez8Gl3nz6dsQj33
JdYXf9eobCvqj8v2uEbUdqrimRYegGXkUHIjO1eCqfQYbavJKxIZHUJc1d8sXvpn5BnV6RCJocqF
U+7bwjoztrzReENrCo+tkKBFao8ZsRRRJzxAm3QfTHUk1ORHm0ALpHjFmIDdT6twUNyg4bjkzzYL
0B3JVk+ErO1ik2Am/ywUB0yYHNL612QHRuXjM+zDsRxcgzQg3Tj2oZM6ocbMk9McyJ7tziTwbXhh
SWmH/7klIlnEPOQp11DaCBfW1gwkoQJ2gO7TDjy3osI3TnQztKRWRk1F9zrBrBl1m15gnHZ0c4DY
wqRvVD6Ge2zTWR98dQ/DHDwTK8KUbgzch62PBgfifmRmgWYAsKnGahpaI8ISyAF8jES9Q62JFvit
M8hcMXE3Gp+CMEU7BXjLd4QrC5EUz6jiefx7RMX64ahHWII8dgc4bPzGmfToLpbnYN6d1ofyWUI6
o4ptBWjOMhfFl3XWMI1Zah668Eq6aWBaDnh44cxdML0DBVpPmdkc/mE+Zw8GQ+PbDrJJZ2tqUpnp
WYiwaAMRXgSBifOOXDooVG36ktOZXMeq+C+z/jf1u/xjPzgP0UBcQbkJNq/M2mCL0k2wmte9qZLS
YD0dF6de+mBtf4ci++XaRPcOHdwwdW696fvEwjLnSVY9/gjrUxgLaY+aKK3B6M6x7418RLfYK8pV
B4YF+K9NTduOK1dbz8pHTGidbtrXB7n1Fu8i5FeLTji5XAJitm0ytzapSqRGHaIFj9q+c9Qo6pem
zDmXO7IXQzxFv2YZihW/ZObprNki9UgDs65CSxokCyZ8pxqUfH7DPBGyd5XjBMjIcoa+QZDxRdd/
kxKkbfofNz1StvZBRB/lsEWciyzYHXOe/AzkC+hV7LElGlukRK9fVzVUHso/nZCb/T+Ty7mDDExw
D8Dzltzwrmh8Z8UdywJLdhUk6LWd9qE9iOILxPL65X4z9dOGw6nkliC+GdTNgfCOX97nCitru9of
NIwAyzG2BhRcWAbnJ7UI8RWpnY06LtFDqLZ6zpT1PlB/a1ropxhcL9fv5wFfS6p790WBab8ouMY4
jBBbT8Ca7ekqEZMPNN3YJaphI4lMpWnNWCS6wk3dBN5UGhTx784zPDDzRwBxmmEQr1/E25/VPCX9
KhmeJ8o0GJju0CeIlRCcLwnMNvOe4KiqqI0wCQUDpJiz07oxrNz0D2yLUNk6Dy8sfjR3wovFsKMi
zqqL8KGmzP7KiKUqRaf8S4g08ULIHjPON/ts5AUM0t0p3JV/82fgtAs9QuH+5zNdbeG6aBdaygnE
Jn6aW8s1tC1+uYHG8E6Q49reTnKcqEx33rwwdYtsB9rJBY3rAoIg0+CZ2AFYeIIDleA1wke4Q2uo
DCpTCevuNFDKw2H+0HzrHZmZFuoYciJMy9xpAQ2nWyfvS3Xm8sxIvzzoWAD8kea4LyUvsrtnSNhT
qdDWTxeEjmkMbguHsS59hh19Frvz0Ur/1yvVWe9Ie28fbTUi2xTDOGZEbZV7vvNihyxpjigzZaH+
FunL4TY/uo40HMuRowrDZhwFHwOSbRBIbS174rK2tbzYPEI5//Bt9rABQzOM8/tq0ud6PMKzF6SC
teZo4gqF4nox0pXleY8ABYz/lqETa78p2f6e7aLN44OpTXqPepuKHd0J58lLhr8/mTpnydj69h7T
Q9zp5aE/3lXzO0B7IXEygzQZNQ8VDqWQJD/R8Uw69zS0efmHVYbb0UXyO5u/1GaMwHxDeYdpVYJI
OUi6m+qdXndcziYmUrL0tXCU/Bt7srMLUhWen3wLM+aNiZjjzD3JcTgd6psg+0CPowMcff+xs4cn
E8GwYahTp8wljYQJRhupZtdGybSKhEIFCdlQGkyuN0s8RLwRfNdAlbo42EZhBQdu533MQ/Cf+xTR
TzQggh78Cewf0xsgv9Eo8UYdnYu7MyHglfNeyJbzw4wZWIJWQNkowrm93Mi6rodHu5GppiE9gFzF
IGmnNZm87IvrMUWhb8tWvTbYRLITQSbYT1NOrhSRO0NcqSHPszEbqjNW4Rq1cybxhpXplK+2+Jyh
9KvMzpTIsc5dvGqZRrS0Bims/Yrvz5IqXWcfVy5QnQFVHNceERI9sQE0ILpKkTH4nNIgNOahigIB
CmYsh+C6ZpUaCSQx8q4XVsAtdCFx2bzV2tCgGp/zKYA3+ie39jdCLg206HFPMNczrqTyY1fgGaFj
AaMsl9s6wk4fFJhsko1mStQJ5Og5m9yl7zqHVnvNrLufm0s1D8pEynGTzAareUCSl90n1nVTNzle
l5E0scBCX+RNi2EZ0DTu/SI4JETtGXAXK/ZMvJzHJfgklbql7Wpf5lim+gPSOvX5u1DcVhdfQYcS
kvKQY52Xew/CY8iypDz6sQwn856DjtmEZljbofo0cTxZmdI4mzm6cAz4H61I9oyNA+mFWbVAvVtX
c1nBZiH53E8FgyX8PLP9p67yJzoEBQFU93EcMHxzLsOeeK1MT2L47cXSX4gPlYdrjgjV5sq2Bnul
+uI7rGgoYfwkzPhwKYMlF0LeI3NYSyVDr4djqcd+qIruNGxujXfbizB1LvXYDJlaYnQbH6I1y1C4
d5cMPcAh6bNatSqiCMbfIROVB1jazLU1gVbz/7JtFm0xp8HsVEOdqHLNxyAU39Le5BNnyerbnAuI
doNWaQK0UXHF/9zSFeWr0GZNrKwO/2R7De5HPMzoV97uBwrzeamA+Uu50K2s7RN8X+D4Fg4nJep5
+7iS1WReYZOEQuQzAFqssQnID/pFL3n/W52YLOmrr1K5+aZPs0+jwOcBKFmjaS85cdkzXFHxDU88
G+PRpAa08uCPD5BhlX8SS4wtvUHOrQl2/14t3/Pd8e6ldDNw+8oiPk4ZPWPXEm5nVEXPsJHnbZug
IOZe5beGDoWzmetaDm3IWoQPrJ/uv8jxhZg3I5r+srszYZwk+H0qc0/ZssTvt9PQixVQZFUO/aai
0Gdf2hmfPp5OFgi+RV17po5PcXAjTUIIxU/JmwspAlQhsKG2QxI6XJ7w3JIDsZEFxGlL2QvEF0Dp
Ddch9VJqAH9XOEJ/3Yuc8gNbIWHFufkeOeHXBog6BZzCl3YaVZVuQh/9xM60DMe3pQ9nwMd2MnVi
mzOlbu6ErPKxwSGty2h2JYWr5KtudzB7UOXPPaBB4FY2XFfVSfF8KMTvFmS+LMV/yPSqe/6uWGBT
AR0ppBrCvTkAcjXqQndmXnYthwlsRhN+nxbB/GL6LWiuH/xxlCQK+769GVyx5Z6PgxfY27S5K6Wn
2RR4ClaFzhddYB4cfphdGAaRe9q34zMWfv0HfxDYQ60vmWRzXgy4KHNmaozfUz6X73JaF+yYyjFy
ZI8voyMS2CO0EvISrmYLoIgA06kM6kSKyHy9v06bxtziLceBFQSeDwY73l9gOwnpc6sWU67lFPrD
LGRPhLb3LyVfn4WcuAiEKfcicfgGGDODXh7Y3lKVf6sLi6ciqCHtihUTEcalXZUewPv2ToPIPT3j
mbC0qlhSEaHgJWaGkkqIyi5qH386egZcl97RRqB9E3NWWzZ5pUY7zBTkv5h75Yf5Wan83rFzOteF
9EWiZA4QZacofNXCJ5Z0ReWUhO459KSUldpoSiUjUtBDkffOMzCfrNBusgRN9I38DXpADQcDE2k6
nIUXn3G67cXSvEbokRkI5rxXBiVX1hjpdCa/AVUtgxYeq8ykosLzM6+zuz6B4eGuBow8JWSOrR+b
M6S1i7uQKhb1A0/3ZYFVIL2PxynuQ3q9OaA11WprXPq3V7t2/niaI4PPMFtjMkWElUJVVoNskkfw
qVpBP3q8+qcAEa6Z6NNL4b30txahH2G6aLVpLfSrBjQFfU/nX7QrPT0aQneGayA8KgY/a+yCpvy+
uqr2z7ZK9yI/CnmrgreEV2DEJM4Qcy+2VS20YfQ/0KSaobWHQ3pN4vJ3m1WaRIXMcX1zIU1wuj/4
HVOi0sdD5yJicHNEq7L5EpO6/jtQ19np0rtMksPdBFJTlG4knKiswpgbcucNjbW2jCNt28tL7xMI
sD5dItYrHgEx0QkFRyQGsU/xy1pEEOYTBJ36hJga3X/RBOjD9J2tIEPpzDy1Q/pTQOja766amUkB
nAS2/9MOOCJML4hhU3kC8TBl4XBgLlC372KeRtph1u35avV3eJK4MclbtqOo+m7zO2AEL1i5bN5z
Blyb2Q8KETZPp8MDsmBJM2GGpfAEEU4+IZ8ZeUC/qadgVeiRs40yfuyv1ZpynfkJYTeRdGb1+F5M
Y65mnnDB7iRDwOyYw534BuFBirQn9dfXT9UjkrWTGWyaxHHZkVD9BvJN1HCJojAOYKSmIenKQI3a
Yu9wx7wYXjBzsDgUAYRQZrTAhlsW2zyvdnpJj3iQwRVx9zGwsimfmKCnV/6ZDafmbd1Gxhl2Uqtr
BYGIgGr4bok4WoQFkqGgIUS7TIIhhuEHnHuLLu4VZS22Tn/hfciAzvSRldZCpUsmzTWz6yWah/LN
uKZs4KE1V6gN9VIjlZ+xcS+3wxpSOEq9p6qVFu6NTcOa1uRSWnEtv+zLtWbqZdmeBuzFeVW1BMLm
/0ZXGaIvma2I9eephy40jq7eyGVky8sYaybt1RqcvLI9YA9/fe9wjU939Qms8NtHSG/lM+Ikczd1
jN38JRI1kWs7yiWgSrGCxJ/Dxk4OrflYU21shWoC0QJ42fDAjCPL32GnSmYR0rnVHfDTYjJRtKwW
+R//DH9YYDQgzczzSuWHBCE4X6ngDQm/X8ldIiYc7mlo0gzTYqjrThURhtlywF0r9z6m7ohjaY2R
l/W8wxNZVZI0JMs7L/ndH6ibgogvirU0BGlhcXTf8/Rtb4m+u88+QS/eJWp/JfG4Ez8G88oxiJNL
dVbZdHhVjaZPG46dilJwKRZwt2jW9h6Xzbp1bavsUh/+8/qyKDuRJMIFj1W6Jg0usXJ+iGriuNMQ
D6hSJ/b5o7V4UzI0AcWq5h28PbjTRfIFasT1vuc+gVaEHrynp/2UHe9jXsrss3fKDV1Y0ALJMnq4
bF5UgfpWynWVC339NodM+SEpnBEytIl7dSIT27ZPfMCMhWJIhGVBovGJN77Bn329dn/AG7ZvCVqR
yXfApPvF+iL+ASe0M7ouYe9j2O6SPthIzDkgFarYqXX/nGHT44Ms3xiDiXk8pWTDgiUQmfuQxnUB
C/Nbg2GTZPnBdI1m3fQJAMDv5mWn24jlohGkXFzkE3pIn7j5yJ8t3hD5Rf7WJcg0U9n+BsjraEKF
93RvH14b07oAA3aqSQacz+GG0U080dGiJKneU6DG13Bssa7nrm5UOCPl6kBi0ztHntpzWDz4RDiQ
Qdu+rbyE288nqVqFb+U6cuwjF+qhqFj395tQO/yHD1Aac6JdCfhmo2eBZNS3O0GD39GGh/mry147
1ptT/LQdY1w9vDh0ewlm9v7biCII3bJLwXgbe6CeZODzIQE9SpUyNZUXFDfxLYrBuw0cG4j25NfC
tUl0a3Y+q3bLpgp7maliVfbqWZL80yTZEiPjH1Fmx9+++CDpN9eOj/tP97enFAokO2WsrAAufNhB
YAxOep4Wg6+KwKNxCyqFJr/bXRa/0ATseaMVMun5JDbJKySxcx7vlzOnWi7uhxlx92YZODpy5gBg
4B4CqmmMHnLiCq5Wmb3xqtIDARqWbG19ZABS7gnsP0gcnMao7bNuext4yDiioeSSQ8XV4Xan0VlD
Xf80YiQ899iqzZ7+qX8oo58+2QmZ3gxShEra+aUp6yIadAW/pwzcTcKZes2YDBB/dUfWPzY6bKeq
e3iwnxtlDXbNozch+Ns1D95DPrf12wuZKWeGPsixl1XT7wnOoS/wWT3meOwOP0RrO3ekMNzK3ZAr
mJF+tfzn01Que4tNWXYhKsDnsi00KWG1qVI6CMEW+Kh8IKhYET7r2fyLDTFc477+6BE07ovsf04E
NXH3ysLunPHfhviAmiFwlo3WKjpEfq3CMXFUN/fCXZaLE2IxIr5ToyNZ054OUkqRpPIxEDdGXhv3
IUw95EGDWdJgOxOThm3jbeagZ8SWyMk6bgjpAh4v5jqOIBLO4mSqwLPvOIglflZRwOFDICR2sZjV
ONnTnL9HXJpzAj9C2rKSFqRfxBuO/3kwYBlaMQRVQ8tXW57vx8zBb9LB0J0PBPGknIVhZsD3Lw+T
MBM5MFYM/iGHW2xlAsWcdWvw6ZYYCZTDy15BsnbrNLsG0BXIYAsDmEoUI3Xq094asStFz6d/OzIG
+5OBDQDMmutEy/c24XI4W9sAsam7YqC+fgmAYr9PKmaqaSjEbBVcGDrwU+Ygg93juhSGB9bV4Lsq
sTWjNzzTMOqjDrB5vxmBAg6PIITmBpamCys0UraRVYI125obe38Pe+iAMs18Awdsu/cbZjLQldqn
Iz6CYhqUmyWdZ8DIpoDnKUCdCgPYgBDfNN/DP1u8InwRIaEeYF9xFefxE7etvdZ+BgmjH9PjbxEw
Yoc3+4wrVTx2RQ3CP8s2CNg1PBQrnwBlolfRvhX9W4gUSnzN2rHQ/cKuzlohV9zre1tkBSXMWCK8
nxlW4ptCiSV+kLPGCoalsjt/G3Wy8dA+cLqAVaI+a+iTWylO4Nnj0CJV8gtty/jX3iP10FQfRkDy
jydcbESGy+HQVFVqlCFjRSlYABYxhiJX1AKtmjDxUOXw072ly7SFLfA8elcMiEaw0HEWTLVTnxln
ynGjE80f/NAkpbCJ9nCh3QGfuSueHl7e5FOcbK83GedheP0+j8UazV/BcmVmL5QmfOAxFGaC04i8
ZeQHCeoNV8mU0ADKZAxn5FxjsTDnqEhGWgJcL5bTUM35pyWdLiKvJ+AV7+wckghOrA4Qg+PWcCKY
I/VfKU1osuiXdkrxpqfQMlWMmBhHndnkvOqxcLkQXV5XH2w1eUde0CxmTjefPHiEeKBh18TqgcDB
LDo4rM463Bts9U8VzTgP7ZUn1XxN4i5QfqWuN3rJyQ0xrbAV8dJ+AruPn3v7ARMg/ukdLNsIogJU
51JyHwvgiYTKLvxKJjcMmEetSuUrtcqHmX++yvd2uPMivmV1VDhmIlWUvC3KBoMt8+AS6+LDx6iy
SnekkH1SdhwAI9lkUjf3GPPdc6iyvkJaoUnfngaDa+UWTd4bFBkl4SOZI6I5opmixpAk3p65tgbA
GbT6ZHCcVO9tthEMM+CUHC/aVeSAiVWxagFjiax9UPinkoBDvL0oftRifn8YmK0H9oYoEhCp/N4p
KRarHwPzB+hQ1KJlmejvAOjF3AhwbWj2pFPASGvdMsvLpVYzWFz+eSVdMiYMFz6xZDxo9QpWz1fc
wyTwfe3Uwa4iugKCAyZkE5cytLiQnLBfi4gLlIqLd1nchHx8lUly+uUHGqczlyftvx92nm/iWcRP
+bY2ZM/8UnaC4eU6Xvvfhz16EJ0VEalO0gHsDMjPS3PCNoGHjK0JJ48Iz2EMypUIGL4B3yyWTb6R
RHlLB6AR3XMvu/iRwfAmTt9VZNh/OPXNQoGHq0z6HnTTDdPfUZKLH5mBuCHvxbzcnFUDEMq25KW6
yyX2GvV9NZwHljVuRuCnUGbb+7bylNoxiYHkL/24lbc0toO4DsNSEIwEjDsr0VDCnoji1d147VEx
F5WQIr4IPua5juyFBQ3NoUS0acj3tKZfw6gmXu8k8OPAh3uINjvLw29PYMItuQbo48tSufZu8ro/
EwewBSVkXdeoIxDYpfePWvJXt5GtASMuYNyUhpu2Gv8uPafX1h+uRDYS/lsnN7lsWb6Z1wWcyu66
GMB3z2Wi2hN5difDD+JgSH4jR+9zzyWmUyDTqVIclOt8FIK6K+h8f8Ew40lfoEPJK9bcxS/MyAYr
uuKXZKylJEvEXZzFdqYHolhDIHJIR0YyrRH/Mk0zDuNg4nQMlFbPnhsQAjkuMBY4JI6D7pFYLLsn
XV/fg9j7ROWr1/4guu8AwGHBLNm/dNgsMgr6rVQky96INnN/tQ3rCW2HaUsF5KC9kLciHfJ393XP
FoJ8BG20o+P3JM+zdIShCMRoMtv1PaFlaAV5Gg7ScDQf7ABWh0lkPLcXCSHBtDYSovVuXjqVAeTU
gJQLSBwoKT/9EukysyA72qshhz0VQ4OQZHVQnr+szGDA1x1rcD+7fP1wz42hlLgUBfq6/ySuWbk2
a6/HrdyEV6QjCct80tFNbYy59PLsBn6UpHXCvu8f4DRV+MiM/Lw/DHG9myGEd9keDCN2fa6+Fape
4/3zV8LrYCaIU3aSgF18a4wW5JoJpbHMCpVvJut8n+ubfmfQ0YNgubbPm7ur0BOl4Vhhn6Gthuq+
k+c8ncU5tEUkxMO5FBFh8rElfOIwBD/Ju6l+8Dk8otHw65eDw/nxNHzBfFt6lp7uvS+O/mqOno7+
Q6fKRzzkCl0SK8raOZjMOhxe4JxtjxC9NPj6ukaAHM3JPpIFBodfO3x23x0/a+20j44Hd2Yzl21w
3QgB7znFC49nqHmEzogqTIqctWNHujwLKA7ERmOdCW6tGi0CtGdO8bZZw8nCXBWf9ua4w1coeaFv
lspwc9ZNwv/TwnKkZy0Gudi52FKwyIJtVbQNR3YQWQfhXToYOcnnUIVy4oRly9DpHaNAsGFgtKCU
k2ctn0/MAjM6A3/idLjQIINXasJsF8llfrToekIq0kW6yn8xN9nZ2+4LP211IzLzVO1iF86qVkt8
ADF4M+WtkXUuXB2figMDDI+lUyj9ENvs+YHQWl1vRqgVHeUPD0IaFsB+oEkCIReWGJdh8FJqLoKd
0f2AKGfG14Q/obTnCPtQprR6DzMPUA1xNIwF0GlUYZR6oICx0sqpTar7LqPEU+P4X5ahTb9D3c13
+laoEYQZRSf/ApFVaZQ1q7DhuaQpdVzurAEkLVRcdZIdR8NvBJV1kyCKT1YL6RVCBKx41TBsr4+l
KQGNFEIXyocd+MslVUi/XtRqWVTV5NwN1HsuHijQvqC1RUmtpgmWgIHGwWHLKfTGs589atZ4u4DC
yE4+Rt4nFPM0gwoLCazlYVACRcga2iM37gHIUTx2iktd77g2fnGN6GfH/9MBii8fc50enlWEXlB9
ep+uYnDcHxkYtTQ9CnOP/xyvPAu6SeK8R6Agzl392oxai3NJLu3OAb+ZHZ5Pg8GhbWVuzI41vR5h
hCRdmJKOg3IXm9+b1dOmQALvkr/aN5rBrrXfFnxqHsQfRxml76n1V5m5gAztEXQRbljE0m+5B68/
RjiuRq1iWG5WOqIlkWUJhKIpYpyjKoR1cOn0vgDO7ZaNweH923lTEuT99Yks3sb/3f92c7vfBwgz
J9yfsFSdX7W86epikTqPob4LUvWk05E+Ikk1CRvuwEBBlGwfT0qnHb+BscpkQDSAWjvWyfDMqPrH
rRZu7kuHJdKl9hKpOV/NC1fBuRlYW6eFzKaAfGrT/iponIzedfteooPDVgk6Mi4bVS/qQguLx/2x
VUN9uhKXU9ilI64nldht/F7EInWugDiJ/xxQ90bmTf+DOaZJI9ZGuZnhJ9MMn4FcQvDI5tKdkA7Z
/ZnRRR8KT0og91zp1OqlB1Ko7aox38ZnBD2lHBZAMuQLJJgG/DB3uYtTeXca3LorryWcZz65sDSe
GvjO+kg6v6WLWr7ONXGrWlGJXgmSXjJ9fpttzy4HTtfOuWLJGOhVsS7WHzVg1tjkv+5Pa/4Yp9eG
d6zwbT3ig6tDWyc886tik+EbcITeHxEzM8LTwKrtghNC/dBxjvjiqaLHjMXM3qgrhZeNHOAli2YC
BJ5vXRB+9D9s4ho0gpbSGkmR3qVwktxuOyc8kVy91gpM349fjsALGQHMWtRAN9d8hoXcHmRx+6jU
C5M2wLBTwhTMa4VXtP+dV5yGohDD+c7UEsuOd2ZoYu4DHyb+yD3qqf1hVGwKahEgdRhbaSbzHHpp
3uvhS4aGxmtKOa1/ocPy8ZFTR8TbiHxChj2jyeDCYAyFgbfK2oR9NVgPJgpu2CYrpeNdeWPLXkmo
bdoP+q9uqk4W1K0KnOb+PqWVgyqfDSOE3fIK7GmEGxrQCddGhNQhE83AAmVBszNAjWpMbsPTiiup
jHXHo3jn8/6yBceyEalUujFOdyESAloRNBoUlrj2QGy6Cs2u91BiBkx9qCmXYqW39YqTswGth/G5
1tJjgQWykIwBTTlC/OY4O1WsZ29qbm44rg2tX65R9OyT86FeqVsPxxSgK/7WrzOEIxvtCc2AVuZq
mLH0xj9AQmxRd5tUxbegCuABhkPrZ8aQzVQeFmFuynBPjZ/9ehP0eepHP0vicBbmcQ1HxOB3U3cg
Mne/Q84efHoL1kovT2FwJDoDVFVhuSpzgQ/cJeY6PQneWwyWlUh0VzdEK1Xc4DqIQhfY9cNBU003
kGLDKRA+Gn2bsT+cywi1anSuCy7THbzGAjpeIT4GGxajs+vC8IzvXqz46Rn6/PVFfadA6TDYSIK6
uLxzHlaGmuzl6nRm0DXnSUdtrEgck+0og2Dlp5QY/E0yyDezwsY7vdgFmGsqB0q8rBcQStv51bB1
DC3ozx8lNqFO6gXlGxhpXWntI4hR8N54XxsY+qvJ/6/xM1wBqfhazHte1R+F8yYAqWCPdKyRki3v
9Dq3eSJlPljIr5RAfRzl0ecxpZDJG6FIRGtYXiCBHWZO0yrFieBzTuU0DcVtTJ8PuVqIN9gRDM6q
dE4WzwlseS1H7hMaWkmAveXYYF1QDOezDYoyQ5ytMn11fLqMpey3IO6vlIj/yjSDXgy9uI4vZCPq
jYVyN+hTiFXiEXDAggN/ecsg4QwsYuRtU+BpBddV9kdR3dMs0l+snTmaFmeDN9ww/Hy5HkWoq/rv
xeNlOUAEFOeoZGBKx89N0bZyUnvJRRNjYk+g2J6BvYH01H6UmLBp9kxp5k2tsRdbq6NcYcgQxlEV
ZD/x4BC+co4KqRolmZRtpY9N1WBHm6PCyBOvaVkIeQq6juTcDECBvzac29wn+2B2WH+BpHbo6DwD
sXjW78ztpyQ62EmC2n6JetDNDfkwvaNkxtfv84ZZbfqVX7PhCU0Q8EjPGhnx10ew3i/M+iQ4PhDK
wuN8009pCc2sV/+e5N+Wet9avjK1+ynGOs9WHoWGDnxw0mH5tJMbK5ksZCoHygTp5dWZXow5TpjJ
RAUQLsEiktXcI0UsNthCXJ5kTKiArLgatU65ZTlB9S+iVCYeZQImqQQYoIRSDH3r3AP8GCPc81wI
qKtbBDWMDP+WyLx3g8+3NP9pKITugRE7PKRYJGQR03Cw/H/ta5vmb9UDaoTjiTIQZEcjfrVcYW8o
Vs17oR0qzFUkNh5C1q2BKgJotpUQhm6Cb4IChHuAAhL5Do3ItT2om4hs6Xmzgb8kLVE1iuWkAYL0
JE4ofkfi9HYovcLifB1qCBl/ntplW8MkW8CHE9XAAtkrvSfo0twl9JWCkuQ3jiCiVRzBFoZ/Vy7o
uwODTj8EWUAJ9TVXpx+gLjh8L3MzXkr54rncuU7d1l0ptO3C07D9pWWOvpyTolC8SWrR7JJmPgVF
6+bi9PgMdBWzHvVL7NYrVsE/VezOYVzM0ap/8XsXe6U/mjMTFtZoeHPHQfCGEgzhPzCg9Yq6dIl9
eQDkEZ5CteCyr9KI9KKDNgwU7iyiZfK6ZUL1yzz89Qj1h2mij8eVzODI3Z7BTk7G1lUzjqP8tqjO
CbOM2RSdxeIE0razf93I+lx5/2k/cr8jOH8wpB7ZhEXCkK7DTXmUasVPlmRb3dDVX8FuoL7ibXiX
FCEjBq+SAF/ij1rIXpqlDcGUWT2emTLgzd8ev7QuHxa9147qOv+8QUd9wjlBMMTY+cEF9zynNQ2q
+1suXsWlPF6GiZOP4aE9UwwmUhpnZQC8uyohe0rOtp76r+/caIh+TARFzTi2eqNIaIDmDScUOK+/
ZsNjKbACNU/c3gHqTlNdaVP2tMAWT3RUIU9aOBCPW4s+hQruRfrBGBThqjRKD93+pWh3BS7tOffX
POvah5I75407CQnLwOBZcoXmMz3DAVEp/IpFinQ4nje7FqO+Qt9ueOAZsh6hknQ01vMJinQjnzZZ
9WlL8oFJW8zqVMHQZCjvBYTG7/C/L9fVmiTf1ig9m+So2dScwshfwQ5c/CP0Bu66H14Z1EJBkwFd
SePnnZ4dxlQtuKjjV/e+Dzqh7f/ZchFFvo16HmhM1RQpwwUDAJNFIqAU9ibaqIBOzcCaoRteW0vy
MHML3bShRRrMDMVR+HIWRSQT4eYzLJnkl4YZJ4VVr8G6s/opF1O7JnZLrZ7K4oqFaX9vmPxpdm/p
2DCwjIOxi662CJNW5f8w6NpKYizRdoRHGcWfsczfoGsUs9eRo9TXn1lEF2rPAZb3Iae9LiUMC9CO
LO9Pkf3YMN2XTQABDGKFvRpRiJUibJdZRINvs367sdtxvGrIoGXSZhVj7oZFYfwWFY1Au3Ncy2kf
17+OOFIemjH3p3skZG40CG7mLOmXU4iXZZR7+qZthTLuVTYqFOzU+jEvEPUXSmXuYdc3ZV8AHEuy
MyAMkYp86kiF7sgo+Qdn9/32I5UTL1671Q0hp+UHbvrzmBzs1ZiH70es2RJYA9CFKq+sWarm/I2I
WtMF792/EPMMq1TUOCMIjVo6O3QwYMtEOnEnM+KkBB54l4/730KxWw36vveQR9NNbb6e7SVTpktx
dp8ikCe/iG9sbnm1DhRnzIqYB2xL4lMnudTTGzExRap2Q9RgyimldTiY8zdRxtwr9TzQS2IbSq1X
t6hKJ5q1T3ky5UyIoKytlixuZ751x7fG6kPJamaejJhKWKoiBAWOY2DrJZR3XN+lDqgUkt2CYSN5
AUtqHsptPSMoIfre4BZaduSQtOpsk1zan+6rw5e7r5TMLHkCMJN6jWHziYApNAggRI02QgFpgC3Q
lEe893zjjC3NLdlBfgha/yoyepQ2Bx+YfkOIwTHIDsQ/gJtje0ntg931dkzH2Q5+chwoF5DvWwpB
mvgXQUBwI+SnEdXqysSqzN68jUFInFkuxzaS9x5LDk9JAeR9V/Oz2wnfGXzRJ36hx4ZOIq1ouFlW
k6Yzb64BkM6Axe9ZEejzYkl1QaUkl3cTUTDGnuCYYGxef19wBYfnwkcDBsjogyFGqxLNVuyHmbKp
CDtXZZXvYyFKfuo0j3i1Zhha2Ao8FYU+m7M57QliL3JZX44hq/DuGkHuFU3u2rzkB+7ETuy08rT6
NW9VTjls5Xb82d9QqMv0oQC711TgcVf2b+tXAue8vnxgq6n3XlXMi3IRbxwIUFe7t4qyklIFNRym
Lq4N474PjRfTa/kWyGrCIx3aL/DonO1VD3gDxgPcMzjJihc7MoZfbdRPvRRtMeTEXmniWLVPiNvw
UjoObVX3ksomA6n2VYD72OXTZU4U3omSY6CWB977++nEvP86fgCLrLyAQ1+m82dUP7CSWVW9JKDf
ptp2j+l95yBowQCEKwX1ita7z+CXP2CerlEbRogirCfhZ/AXTnMQxDGIEmtjsBYwqf0xjZe/7/hy
9UUxTDswNXGX+OAv8RjjgYalCnvrFovDcbA7Pgo0ZYM3HvJPn0DISvz7z417wL0HB3B5bmr9E6+c
AQBBdp1zx1GbxhfEsUn2Jvrz3WxyemMygbos8Sxg0d338RkSuXBpYbFuWU/0oaXnPzHkHgbjKVHi
EvC+U8bZ8qb41JqkG1Ts9h2DPJZnKJGNqaTS7wpm+B+TdFzya1dVkXY0q5/vH50TYaqxhlxpaqZA
KZ4UXJBOEpRUfbTaU4ysgCMd6GSbBHfXEHD6UFtho+mQdlltcPE/XuuChClk58tkDMdh0rzPyJZ6
b0NRuFQQwNbCHiaRb+TAmZtYU51XY2HBX7WpibvTi41JuHnUzCE1uVNPMjTc2VDZqmEJHbRSsk48
Z+yRisO217i6Kpiqx6ncweNDiALwhj3V9WBRCSB0vnQO9NN1YEwueyqe42l/YjpFv/OywmMfMuiE
nuetFoiF6UVRaYJU6L5yDPwmir5SRzQm2iACoiv0W8Zxvm5YNGHOBdeMlg0a9EuUPIk4o1Ad8chL
A2/8XkvEfimJtyCxScxV6R1kpQIb7zXkMgXrbJz3Y46h0uDkiY8RzLzKMJEhhPHizMmdhEDmTqqk
g3Tk5sMjYS+iBdHrF9H8eQTtscqJv5UuubmZzNB+1zYCkQOIWtmxkC/8qflThbjdM2lyrpmLPdYt
gRwWbkVtxeNjFMyIbKm2MIXCsArYI7jtY5WRJmv2inlYvdQ46qgeE596veQaawydPCIM5FzgFv+L
1xtKNNAhbrmdB3g+G0jbcDE/nR60rRWVyykxv53b94nBhst5V/a7Tm1QZOQ0f3yJzdhbx1UI1FDy
Wfmvc2u4Zu33GzlG5goaW8ZwBVOHE1X2Lq+uRVJOqPCmf+PptvN1/0NgzT+od8tJcaX8uA2Jx/v1
IgopiXqlpIjERBisfk5Wxnw8BxwfoaTABuU8vv03xadYj14IW6YDDd2vZ3WRwt0A5CE1T2gjiaFN
aO7iOY5KsAsAOgEqYg5uW8DnDoljQAaweijtZC/0Nvl88wDBELwslFkoXFBA7JeHKHyaMcmUSTVD
vMN6te1d5Q/NfzvfHwel+WJMn7f5izy+AzQuuRtPqxi1DuBgHK8saSHrW4FHV674HcUrcT1V5LFu
zp9IF2q/Yqy5tg6fc5Wdff+Xgx0G9Yc99CbOxuvYuxBvNT6/RcjQbEIu2cF0/n4Dl3NV7lFxlaDj
hUjOQoljGtShPznZZniJXiilKL6wekzpCZideL37dRAwNGbs7aBGsPEPxzh27VfKn0ckkrUW2SYv
FDLL/4lXACZVSc/QM8ocnxmFQEG4sgRetIfgKqhGrllkju9dKP6vfwQAkqzdkmxU3nelAxKE6g1o
ZylhZ+gjMrpq8wXu1MT5WnXg6Ise/Zg1nslxwAQa7FiBAU5vXAREOLj18/n/WuoQ3YRwD2zJK8R8
dvTmbzVQIMdAWK8TN/y2DSXi9qb2kQQ+vEUYX0HgXAQDIse8XaxAf1mUmVULULZxz+NfBh9gVEJ/
2uiITPeVgxeNxfJyXLnn/2r+AZGhqW3iqI2mF42uOYkyRMpxcSx74mKmvf+Ir2kDV5SwZjwRxskc
oue8pHb+J1/5LwHo4jKHvwmuALYNTAvjzSY/I/+2yhTauZK8E1X75uWCTAWHJSbek/x878mjctLc
BpVtdwpk9qqZgw9RHX96rebcJ4IX12WdfoH+wyFYF9pW9gzuhgsqxXIKoZ9LC7Qr3is64S3AkA4D
pB0r5VNb6cuVEtWXI/vSl3X1Z+EY/l9AToy7OMV4CGnPdoTYiKdroufanylXZkXFDRbxrkCeJvyz
g64w6t2GNrr1frPDg2pPkvHw8lSEzt+w9RsaHuUYyqhZzm9gZ5Mzck21vHIXktIeFjr7uihilU1V
X6F0lU7ZJGIwHdJyBvOWFV+hmxe8wScnt4j2ecryZCCiyTyMNaVbWdrkmW5EdGYA5zJv3w4Jz+23
DVw7edFrZwbBDhplrn8uGaQnXzk2K3umBAa2ykAM9FeWTKeKAnHOBs/GDaqKta+8DzJLb0Cp2e4P
fL18yZrn6HdkCpXk2Ier8i1o54FmaZ/mhCygKhaVsx0Urdog21ynKJqVMY8NvH0vmypDFPEERr5G
gdd2vDw3liuAlQZ+K0bPiOZl1bWMH000N6+FWakFwHklPO6K15HqOApvk2zBI6SU3uUzmtepYz4y
3vPYqNYQr8qv3biaHfYhsZwjbvDPKeKcjlc3NuoSdmlNR3mXna3GT3IgFSJiV90bHebMS1sXkMAc
bOMI6F52Dm6tdtL5Fuw6B7RaMOAR12jcHDEgo02Q3FZAFS9Hpp5foRzRv+Q23uz/RC6nCN0Fnd1F
Imk8V0jNJW2T0vs8qeqyEuhJI8vOcjBC1TZDeQRI4FBICT7vpOSKJzLMfHnLqKNFhfK3QnAzzu7+
K3bZbRqk3tecBvyKTovZzJnxW1V9hPC7LsoRvecN5Rcu8r2OZIhs1hNBq53TxP3V/BOP0w3gY++A
soCa9y/Xpu8RLASw+kyrpD0J/7ydOdfd5hfU/UUzwQjzsdYwjb9KAG2DjnhXYmYdaeMIB5jl42Am
h+iWLrZ47drWWNYqXx7Zyz7LVMGxMTats1rVTnsVQBFPsDwLyrTmpeqR3kQ1vc0ki4KHuGuA536S
lWhjWverePoD5jb3rcz1kmxm3aygmYcwGAUaIFT/BBe1Amsu4HAgqFp8DKjczqQCKqV6kfXVqyqG
/5kbQxmaakV+Aymh489Efng+vSlexcNh8ebu3SqhHOUZ2gsR2tlA91Uahwj0Sq4HcxynRLfm+r7j
dNh6YmQn4dEnhHZIBbSLbGxKp5Kz/Dah3u9C/tXEgHH1nnhGBWqsXDK0OKwAb1luacDVYfWtANcC
q0rLcb/lLz/cccmsyIgO6eiFlJPSQQIQMRQvqrEZ4cxDNujXK5dL1K1v0QDGvuM2LVE/hze5gqqG
RBb2j6zlch/WhywodPQWbrRtb8Up/O9znZS4p/LUbHjcgQcH1EuXkoLzK2fHnvunq7ai+zkw7dMi
E2ZYFWgc5mvg29sZKrkwRrQk7eTE4z8cs6x4pcpcmjhJzH76j3hPSjokswd31fVrxqfKaRYKzzuI
BrzYVSrut5eYX2EsPC2d+GK97SirBeUzvFh0a9vZ6YuMdY+KQAHFz9yjOpT3uoyZXyfJeXswzyGc
kyDUJ4lq2AvTbrwnQwu5qb9YnKkslcrCu15R+KWbl1T8TvPJLvy83T1n5IWtnVMpU+inEDdWuhsV
R4VeiBjk8mg0JZiRntz3vIQ+xWY8MoXOOnnEhFXEvbn2CYE+7VFCbXtLDofDQ3qRvE7XQEUNsl8q
Tb7TnWHv1ckvRL/qZ+7DoMspwo3FkjcMTYOxGmfXkWLQ5lv2HeLhQJ40fD6XvysPMU1/W3sBHKbP
pftLAgKaM0S+R1nBHEjc88nGFNalVVeTbEb6qKUXsRR/+IeJ9erd0vv9NRenbPeLYRKo0ncDOakA
+OigrYqShWVXNfj/h3rZWgcNsAU64b3U22QyBEKsTrM+KW0dMKJv4xC+ik0i9jr5jei+UYQEnvAc
pQL7yarl7EDGx3pO2+j0kei4XxB6/qAQ23Bykt4UI/Ptjr8uAH3nrTuS0gJWdiVj77IvhBMa8ZlE
KLdgrxDAeAGFD9sP5mthAjJEGMzv1qozUv079D608Saz1nCoRhdIX48DTKKJI+HbNnZD8ybk+dNz
KS4qSJKz/6eoupoHpdWF+H9HLcxBq8q/e1m+LYTjRUSElm03XAqMGPiLTnO+sgfox0+3qQpFBBmA
6AIEUUQAlgk8lFchuSDhevLVEbciHEshD50SAusJFZp516vJZuS9U7XHFynFCHgCauMh6gcGRTfp
UTpL0LKzGzDrrhzxCJFFZIhAHIk3bmRopgLIMAbZHN7r3UazwrYSfmdhRgMaXSUcfJvYJuCS+iCw
XoQX4ku/1II3aDDKT+uItE4mjNO9HlhMfESccPeAtr9EQmMx9gyG5U1x4AWFCaef+Zz8r6nqx9dD
MyQYOd1GazGogYxHfwIHgYI08E5sjjebN/wChnaBT4bGPloH3K9U/TsY2rOXoQ3E/vDEx9xE5lBe
HvRQuLOSg3t1ErU/IOKHPDbwBfz/SiKChNRZ/Qe8btJex/pkD1cQXTN8e39kYgankWnD6WS8eqoY
IlXlYNhWbpW/cn7gjnyifddmRvPf6kR2Nz0fVITpR+e/wYvmosUr5eVppOGPKsZNonQI5pIcKTtc
h0aQhwJBKRjrY+FfU5UxdKrTXtvwqR1+Ndc/CJpbYrEtygx4YVmBMjhmS4FuHwxL0T4CvSKxJTwC
DA4khctlHcwNA9qLOxOi8TLdkwQhpM0NJYCaMGClzBk6ENmqXxf48ksuwEFxyMVuT0lK6dOCleGp
7/8vikON5Wr3nwIzwPbKxltLaKJpCULG7jz2uN0c8XL1G/SvU6+Eq5YJeG0K8daxffMZnXlAMEMO
T0DB/U/wy1AlZLoM+HgE335UyGHcwUgcqGfPZHdXprojVDf2mDNabpcRuHdkJVFELZGwUucOW38X
SVLS0d8xdUvodyE9sYbaf3ELHoQwSfFuJdwE8NlZ37c8VgBrYJ5AX83nWoULhK6dUsN6HfuGI+YM
Px8FQd8mnMgGZY5cXp1WCyPnGsO68DL/D6E8l7bfKaXpU1BxTvbJ8PoRcuYlINJISpxORoYnd0D8
mfmIFK40M0+a5cVYlmGgFXO8sNqn/MR2fW4RGtAtF6IpJYSLKRyICQN+ywdFlPW989T6hu0KUNm+
ZAS1r+OiVCTqrFzZlzeDaxNfSs+DL2EEzGm5LUdomynsmBgHmlNuvl6YOOYEHC6uKrXxAElgfKiz
LuqZAuBxWHDNwlE4x/WVgqu49cYrOj4lz0pIwkxLA5BXrl0gtzacYBbXqV71AwxR/QWxo+HW0IH7
d+sIcxZMJlg7A/QbHFquj6E0iA3Ji1dJfOD+I21SjuvcbW4152buWhS15AuSahocaRfOGchmrRYm
AXB5PBSYifJTm2+fxLLuXDq2buBnl9aIpgmBMjLqEVIk4zv+maWIbjcMJkH+DxF8cSAviAG/DAYO
zOfX4ZyVmAlD3lgcgV5dTcxzYGLWG/WDrY1y1JQlSPv/rgZH6S1r2+tNGoru41S1mDbFKFlR11av
+F7gu/xC2oaAxaD1CUMLZWJ23zQC34viWiuHUTHiY4/VrAcSZI+L6y8wQOzNCCSp7GzPhnkaW7FY
bY2CXFhGOBYOCBU5CY1jL5RSq2c3PJv3Vula7njBRnnNWh1ZUW0r9nUsElwhcKiJx3LNPDRGQW++
45fgVRmKvF9/2d2Mk68u6K/pxlJp2AkxMBnsxOH1ixwPtmPZx4v5oWSlV1Qzus1Bh2QL4hYyAar2
45vt/KWguENRV9SlFSTmYeZK6PqhNMPSkmjewxfYA3LtCTSy+Gjp0vmggJItZNPmd5Rqy53H8jW7
opNzZaZN2ibdBGr1zgemWx2Yjwa5towcTQSWseUu3q7W9AI6pZQ2KTMZXqlbTqJV2a+QS+84K20B
ZeaeW/+nia0EXDcTOHOi4/xQjDV3H4mT6d65XcuZkQeyvahdnlZSRcNp3p5Cyk2izciTU239lsSx
DIccJt26mi3W8dT7W8uiGNvEwX3DOzsIes2fICGU1t6JDkgjCsJOCiY+aze5zAMjZYTY0XEt4Peg
PWscHMk+vx/4mDStovVYZul+FqGfaDYKLfg4G1Q/0bqZXNLsfToGxgYEKWS5RIdwnR+Rat2BVipt
xy1NGvtgXpld7kxNIInz5KaNxEiAFMbv4fnjpLVjudjMPNUPRIyUvFapm7MY7cOM2sFL8GTHSE9B
FZg9Nv56V6jvz09EfkU7sc0hJliHpo61rf0mcPrNDEwxB9BkCC4p5K48UU6Ct569KYRouF3nKbfa
ZtB0WWCKzLrHjjCDP4+NJaw1U2X9s8tRvu9hBO3tp3k+I2iCCJIu/CK1JP3pwL1ZmnoxBBo6hI3+
VwNSo2kVqXQxgch58iRpCZda0gozuRNIsQqvPNnNJ2tPuObQC3yevAeR0t04VZ1xp1rPvxQvu9Cz
3RkzXEftMUwziQY0xK0did0UxjO/e++rY9F3wivnCu9LlYoY3XvOGDM+JV63yS3PdcuoVmGQKSaf
hqGUqmG66+VSg2bqHXRor6UClspfc2zX6vgHvkar5zLoR9JkgnwOCfSm+XbLH7JtHAXG6UakICde
d9fjKAxkiC3ZvM8bZfyeruusST6irA2A7BduTL9av2w32QcZ6SrYfQI68tHI8xPA1lLcFIoS43T0
Ce346X+Y6UqAcc3+vcFznXJ0+ek7TG/FLvYXWfIsQw4jaZEwqtcxiWAkS+f7f0kP+9sZKIZNi5F+
bs8ge3z7gLuuVmQ2MTKBg7KqBqMmi4OgOI98Tbr7TnkWOatoBkV0EoDMtrUTaKngaqAZ7kI0sugG
WAca09nXONcB2p9Pkk1KOv5zsyCCVetqf2T+n39lO7xSfXW2zeIkY/l/nI5SJ0Ym8oqb+WGqhdGr
ESeTzd21wTAKwT91JzE6/VWh8HrXvz7onADawVWdRN2CYHp3033mJXNOO6kOEKdLIOXvG/fEJA5Q
mgtZ1MGebrERB7+XBkqVRaZy7M3/LR0fE/RA6e86tDCyRKvF3xiq9zpt1HnzFpciSv7o5Yx1I4iA
m0D0R9nqlc6skyYcmEcflBOm3gnoP1hRdf3V/gACtFt4xgoEJo0qTY1X3sShuZOMuD0dMWgbUubV
vNM8KkK6aZ4a3Cqj8faj3TcniqdoN4/+RfhEemHC+pdTXhL4TEZkRo0T6tmYHVUZt/K5Gd3KjUrr
u2mtMFZyzX+26g/THs4+pXktodUoMpWrQQkn8wPnkGHD1DJZ3PE0JJgqCzEP3wp1QjoGIjpW7FkH
Ikjq8NGJPf1Kz7Bf1Eu711slOOZLypcNaTZJVmL9mo3fUa6cWBJSsyqzyZMhFVa61DFhCZVjLWvi
gTofW1q56iDOAePryA++SLA3akGpeXWeOkPh5NA8vzGr5mWih0iZ8iEYjA3xS0WCgTDYiEQM9ylG
ne3iF4cVasqBllBfz/K5Jsraw8/PZSeX4ggWIcpHX3J6GHkGMctl8/vJRZwtXI5jhBsRJlUJFUzd
xI6c5GP584tkG+Y0TpqMTMx+aECIqP5Qw/ayfpVHNA3l6CB5icUloU1dfWByJzNMPnnULhG1R1gc
Ghnld5PbdoF4RD8yvWyT1d0jaLFjS07+9jCMU3oGV3qe5UX8kAeL3b0vFNVwpFqtGg9QtG7pPD/3
ct8UacaJL0AKDitn8vHDo2JO/oVef+H8QNehWIE2JD1V5N6BLiS2AIFSnjcjHM+f19n/JMVDYWN6
wDeBXdxDO3no8FkGzJE=
`protect end_protected
