-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Kq/OpX3BipI8BSqbDpxPyLI2kVOvc6yJsqG3MhB9iDWoXtUJP6+A1o/k4zzOxZ8+MfycufTBRneA
NFalY9mhCwEWu9AZs5EUCgy8C5AZbYlwwWfkoAIsUsmmjExJ/tPPxSxKsng2g0vb9jYKKC7wH9jk
hOV0iUhM/yvheSp9RLalMcW9li07hAL2D9FRQ3smnxkReJ7qNwUNLtBUloLYInS3X1YVgvxeTsEk
tmAbEQBvQPURpw/6emt+XZu0lUWHTyuLeNmtvJWYxkxFG/3jsuXiQNgYhSyxSUqVfEewGZTdnITa
G2eR3Del7GnoK/SW4ozKrBf554qraTLbofMZHw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14656)
`protect data_block
HhVI5Ctl7Dab0n2PzSBHs32mGzE8MlpniHQe4W0p3ZiUA2AvUAUUAPhEQy1D0CpS4eFWeQap1s+p
iC+uGKstqjiAUvUUaNlI5ImhBDDPn5emZOfrQsx3u8wOHHBrLVRf/rnJNP4VCeDT+ZUf6/STBe0f
q/39uwVU9ArIeKLJcn0kvgbhkoqpRxrwqYMoa1wRsk+0thpKcyDaYpb7W77/3KotZ3rXESupwSEO
pA1GZUECCcJVQBnyYTnAxtEiPrx1sNWWlf0IfMqkPowa9L75WPPo+eBhj5CkCq0NlOP6xd+zK3m3
Kb73JR+wW4+837VaZd7KvBnOLvf3WtR+L1qd/dVrUKrQ1u+u7BCjftszrm5mCRsqpHxHJkhgnO0G
fBqEv4NyZNKH9vUdWoWqSl/3oDGj6MN4mgu4L4xWQ5MMGx3zxvUQxXMvsKdV9p4GP+Lxwz0jpNjq
25L7CyvpGsuSBDEYN2543MqSH/Vd8h7t72Bmet9bTYgDtN5meyM4/ZbyuO2BitNlPFmjqZ93RxLp
YKMUpdE5knGUTOxyEpt2cPH/lAlYUfv/QBFyXVVT22ywW2OS8UkNWMuDtJ69BfkYmNRwdByrQ+4U
dR68tVPfhq+UCo3YtHrmB8yfiUjEvC9b9So52fdmxVSIOpWAMmJusu0Qxieytt1aVFbwvTGRo4kD
DKR+98fMpuXuZj3JWNvUiQbGLUt+Z7qZ5qjbTik1If9a94SMo+CPu+zBDdUX8bd5BkGknVWKwpBJ
s5/wpKlRdOO76d4qvSS7nxtUj5FjCQ3SMMJAJeiEunfs7ZBLmrM/FzkJIoGcaMfy5pl/f4lXWHKS
YXOjq5Va9Qa6K9jGJQLTZueOvEqMQTZorWzkRuSlHTJE+u6jE79X4HLV57b/Vu5xBwT5rfT8WFip
YdSNzbaq5ObzUXRp/8jCfnEz1wJV62/PxxtjzT0fUaJtHNDIxIp+QxNsTkakkhhB7Ez9mztjOtzW
pBqpQUT2o6+TOol6fS3PQjfIRFsDIvLlxaywaRfa3AJRxPEkbcoCm6lX9G9kSKZWU45QdaQLvHfp
e+H9jiLke6pLRYZfhPqWFJHpuCgFUqKvW6V96x7iQOX1IN2OSdulKuo1M7xES24KZ/ERhiZcDiKg
2Wxxj+BBuhWBDHV8Z1XtKjetJbb0yS1Fz4E4FD1tujpmTlyAPVNHWyXatiNcCpR8EfxlP1Xu7SiR
utIklAxo3UNsyNBHF7XLIyhGzdUVgWxXbtt8NHuo/NOoWWG/APCxyIsNmtDO+jo9iXhEz1ySu0em
Jk4Q1mhIK+La6cHTi4OukYVtKZ0OLLHmdOEOeel/rtEB1LWh3dzHga2f7PocRZbhH6h5BRrJuzSX
6KIvTsCb8zKZjjjECgO2snSCZmIE/9uJPumXxSusqB48FLQfbQczCihbwVmOfvQZbEFu6k0JsvU5
N/KyzLIvkHBDwC5Nj0SAiBTQB2Ky1JgxoyWEMFuSq9bMwBpOE9PNgHHBaQBVOxYaWVr6GyLhkirL
R4Yftauv7HIBB7EunPhbqQiGH6y/eFysMHQcqRqUlPNL1j7JDF5+mNUrgPgs50otthx15rFS8xuT
k1Of8NkinvBWyhwPydn1fxop/IBiWKYBIDVx3TNObk+CfyBhg/v8s6ZfnlD8eS8ymz2ryMYUhF6P
+licjYOLMlQuKkq76ULHUYBFoATb7Jgjdmz/QMfyk6hbJGW8xmm5xC3uMEKZvEi9iQPF/gFkR7ne
qlfjtdGK8ra6L+V7c4WSTjmMV1yc6Z1uZEdeMy+6HZFwWJZ1K8lZGXfwJH7Y1sNvSmr3Gs19m/G5
6hdNVrCx9dnCova52Ub5ZqTlysruXtzKOJUqdy67n+ShnvljrhdalZN+VMVfBHvNt6d/nabcT5NF
TM/BL3BDgIBhjr7o6qVXPiZRAJYf2RDm9zbsPWSHU8oJlSsBKsNAx64AQAr4CFlQfpBuB7o1xGcj
Iu93mwP0sLDVifAEEKwBbgnS8/GaKMXUA0NhdGD76Lf1QlNbo9nZtGIR0jGPWJRjdaD3aayuz1el
WMPh0DiEhCWqIa4RMzzXj3tUmPDKNtmgr+w0wfR6gFVmeY50TsDgmoAB9Cc9NKcEElVHTnfTnXpL
bKAeJZLlTzqFHvgSnc+sAyfKnDmxQBeibYrjULRl6qu0Vuf1xuo9vZ2EQZsM19WswvHUdrT0pRWk
y8XlL3eEVQKCKLU7xAneuAFn3gHD0JLxFrxCnTD+ezcenOFs1EkE5SOkS0NvSAYFIjzmglPFzMH8
6y9HmOiHrWLF3F2+avAX6vYchIvkBbwxNM+xEMDFgNWDjP+3YwgENEC4hQXgQrwN4G0gcfz0cO3s
PiuUdUPKI1dJ8PyjCGfdJfswl1feTPujqz3ibQ6NKA0Y2FiOa0P10PnIeK6k0NRL6Z2zbsxV5gXi
Tn47OTZf0OhWo0Saw8l+W8aila1mbkaJkGO2oqY5GZ30AefD5omc0KPZ+auehCcPzLj/PRRv0ckW
AK1wgVy80jSopZfRpeaLnJAuGR7KNojgIcPfImJ8stFW2ZG4QK9Zi7ckfY6sPTIdztQJa6NPkYSr
7mfJNzbPPlI8iU+RRbF3C7l58LlAahXTFJ5rH1SNkPEhBx0QeKbdarOW7lUKU46BayHahZtsrwxw
NLreU5P5AzKlOFzp65XIUuvacDP70m5gzt4/AZxfFJEa7DaBmEhz3liDKm1buTOU50ESO9CDLy6A
QbFZlk6IiDZUgfhzCLtzSVK9T63ZGHU049RTq7WndvdG+dwc51kENpgjvPw/JCGsUTl0QPJIrv4w
OGKuSEZsroF60pbwnxzrxa0fr5yNImu4qfxhI5yqtJ5P8RP7zP16YUGFAHRToBOk0hOerAyn+Xt+
EQaP3OhDvqSJSHDwGOZ1i+6aW1xlF/cXs3lPgetg2Bjw5qds655wclD6UKWhT1blaZp9LylKbO1N
GJO/igq6sGhvQlKhjLB8Mc0Xm9mG24M/5Wkd1ugS/Oe909TW3/eyo3KpGvYMccCapLoX+JO7HDWH
JNhLHmj/2BB4Xlv67WzkYgv+MCebgxwfzgI7qjfASkB49CHs966sY1donBLRZuijAXJTES6S+/+2
aoO5kHSwEiVZFPgoLE1sVRIFcVLaSOPU4lrtgErDsI/WF63IAyKERKWhiAAjD+HV25SyJvrTU05m
omtpSKaEtira3YQ+9O7Yp4QAFwouMFBthGEtseWBAkyuIECauzaYeyCBoAi1BvHaYKTCHyuVCKYu
cTA3LBBpiFTGpnpOVyHFzdmdbR5q9gDYLYSCxoNRyi2lO9Ca70ILMYwTDR1TWAcJsVwEskIoGSZP
hmsQuUXB5u/0B7Si0c/XySXzDLrLLMYRBtZTr/d8Kl4Qlhc60t3YSBlTxSyGFbGl5TXIoc3U2Y5Q
t7HjKM+DU0C1P39qC30Gae8FFLZWxaXeaJgNu5wL9I3pcMMyNQUMxpGAOlikB4Jhj1J9BQj3cnpm
d3f2rDMg86ZLoZw2t5OP1yntKV36aNQ5SPrZ/LgX1P+rLLBWcKmxcFhN5m0p7KPaBeHcfzTJLK/7
doQl22akWNEW1+upKPlosk/Hof0dGWBBlS8O8R/pL0zJ60AFKrJpxRyCscUJTUe4T77EalU8EWT9
0TR3fbJeuLyOYcE2y5Zo/8RaZ2zOXuHw8f7hppusF0DiuKmZZsrET96zYa97NrW0Xa6nOvxC+VJh
HepqRrw10UosczJlFvdkhsNK55UV9/O6RZi3GOPNQK0Lbo6sievgUM9QHqmRG6Vs4otI0AaR7xf0
zCOUASPJsbq4IxJlx07Dk3EjsP4+AWjRwLwpYom7z4m5bjaLo59Lxitw+hgW7eiZIM5QUQ8rlJ0b
G3UKPG95M8AMM7uQKfBqCAFmwueK1XdrmXmzRWC7dI3+PoE1pZ0zo9YBAwb8V5+jiUB9NVkr/w2R
jmv/SJOCClcCMjA/J2DuBKrKw/Z4LZxTKVb0slMh8b6gpjpEMTa6biQHUsBmf5vmlvn3vXGZfSR7
f0NBP3qBGQe6yQBbJ/RBXf0YxpqOi1jCJn6fIE74+CfTkXwPg78PU0/9nVj++NcTouoZinaTK7E1
tH+dtK/Wf2Rg8MybV0Qv7w16BqLAq0hX3YnsqgfLMaSDAc5vQVaQUJq22QY6WqzU7QkeZG+XegNQ
UYj5f0LgYMZXNw+85JhIK4stv7VTp0K9dtbDzt9Ysus53iZYUF47zS5Hc7REn9A/tE6faheMf0iu
EINDwMOzEF5TQyr/HvzqghwGu+QRNooUtnbTJMxbE2E53nbr2/N8p6Ia4oOvNhzZlK/lj2Y+jmWM
u0sLaxjqBy2ml032bgkQlM8lSvOllEYeZLvf7NHh5oa+hR7mOtZ7NGM+koGjx8Ed2EusQIbtrVDm
NOt4XpWElxyX4VKEFuNQiC5Ls5ysONdI3CaIa1BxG9wYCjjtqdiG36dj9nXpxeJDKcqbumY5LeNk
n8ke9kL4VFckJhBomRr7TicR3uq+AExrNm6mW2fqF49lMRAqSFLy5kyW6dIMWVUgG4Edgt/FcfeV
BvOPuNHYJO2Ce2BRDNOczmh1eldrKgC9vo9zcxRHOkpWd/PdYjJ1zKcveagIIkiiaPo+VzkURfxd
Byrdjmpq3nuRzZXtD/rKZrQZ9iKLahHW4KGgPICZeJgJNxhQyny62LjGD0LdGGfh3ATpypZzlTy+
5h4hRuHQhxRzuVDvb47m6Zvn7MFqvjznuiprzjQE5WUFPW9RuqzTkpx/Cr1mvLTYClHMSQ1uwg/4
yf7A/I3T+gV4hOS1B9XY6jUACQynrcUe2RXGlSbVlSevaSeqA6RBRx0YzwHSYgMh/7yNB25syy/k
iSDCnOQheZpn8dCQAClvVK6VdsV51ahcdpifdYwDqgxiGKqcE3USkeEYX/yyZddHk0znViekVHR7
RrUlCc7n1EAD7F9+N7xZMLVD3yiyq/Ad2nYk26lGChEsO06y1MqMFKbJdYAjspqfzhxdSSY99SUN
H7BxkODfxwLq06XfBGl4ZDYWYDqXtWaNL5V0qUBCfMGyKVMsZEIL53roOjbYMkDA6SPHkegVZ26S
Pkzoj+RLCrKoIItBV5SQ2oNeudmV2WUF0fRkagGmBM6KyZwrlzZ4tw5qm2pgZYjZLcb3sr70OYXr
H1cJI9niRUGe3Vz1gGOrYHkYmbwdQDGA12gmAAqzsBjOt9dz6J+5C9Uq2//fxwxj0twsIWIAGvFk
5KKcbnFC2rF8X7aJWT8MyI7s/cQK4anv64sPWCkOMMbMn84x0nLDexXYhCZNjmMJ1k3b2qaluouv
q0QG00p1wOXobaK0y+EOtY2xT2/shonFNggw9Xk5Qxbvy4hVUZggKXKGApz2RCiSw4mRLLqrt95f
8IH1VOM7m7RYJVw2ppESc87ZQBSegSatcW3UhY35HEqPGSZ/iXFrQgwTr2HK5O1bx5+3ja3NSIfr
L3regWoWGfNN5pD9xdZ0y/rJsi1falCQSlSUbMinL3Z2q/C71QDU3wXMzH/NReG6IwcNpjbPuaSh
PreqLBGAJLGkf7COQG/SyNDqqmfMoAq8/QVXHSyx0ZjjDugg0D8202qimisRNxSivhdA2QddeACy
XkJ/+xw3qvHlvUkWP+6YbAqH82ZEOuLTsBSrZbBcO8Y4YPJcuyDOz2dHPHSNleFw49Z39OqqPTMH
aZJJAfAtwluRm1pezH+jc2UGg+FLgnwdEpIWNA0JjLaoZkDpDmiEraYLLRYN1wrwtrDh0ImuRIpy
uBHXNQjragffYI7css3escBWBhpAETiXD2RpYItGv7yCelUpNS1oUNPZC3INCZy8ygmZEwfzvMOg
CPB1ue5sgFfFtFwvTK/wgdVnBxW3cgkoz5b7AslxvDnh1XjNtujf4bxrgmaVuYBUv3J6DcrORnmZ
qxxicswvR3Lapg20JfTKB5czYa019VFOmfXvYyJGeAkaKOJMPMNzaBiCwTfRyzpnfA7S5nJpF7dl
0Xhhy3CjI4meFNIb4uL8LpNbIbbavEV99Wf1KJkqdcUaFoDPkTQl9OeMIyc0P5sLDkwbXDW+4qi1
jIWhxXSblksaMvr0YyebLd+v0ThxtioXi3IjdxdRWJbaWtQmx4BPlQkcyedsdnHBXVVyeEnN0EHE
3zXpraQjEyQQlVcGR/fZbpn/0ozm3k1aeGtWKgKS4MpmZSCIPUUrTH6xDZqgpMBeB9qbY/gSV6QW
zKqq4f33i52h+77gM5y8kjYm6kO/8I+qpKrAt9TL3gcgypEpJqFwyL1y0Iy8G2m5roOQmxmzDc4p
aSFCQd742os5o6BR5SkVyCNOBHpYXgpbODpsbkQPNWE1uAji3Q3L88S61COE59B5PcOhkq7ZjCgl
6Y2ljHtKG+mxmonB6iVF+Wlbacz0GzH/ltyFuIF3ez13rYA/Wd64rDiwOW9Qbyn/WhYBFX1kj2DT
g/TbAOtUMY311D0KBF3xUY7xibRJoNLMmL4qgfubUOF9iAQyrasc7Fddt9Yz2Tp7ltNMb1nqFl/J
PQ7cbpocqz3CKK3uJvZBO7IwjrpBNJyhtA+35R89xkBl9BqWaMhvTZeQzwi/Xr5NthZs1Xbp62sj
5pAxIFjAjxRFqSP4t7gwhhQaztwYaHh7OSZpQbeMBBmKQxrh5uuE6JyY3MASM0ut3mJ9tkapKnhr
HicQ2CNWl2PJ2Qz/Yj7ZcJLU16voweNYPXW8lz4QadX+svbwhEnq+5nrXrHm8nZf/L8/qTTC0f9N
//ldRDDGp/gaETAUzRNoMNblNBjoXZiip8mBgUekmhY276kBVwTFsvXDnpJaRAoY9nQ3qpraNKST
B4vgTFPk8CLZUwPZ4CO0N4urRBF2HMOMx8edGk2zML34z5v27TCKU7FekjuvlAXXmHuaux5w2qA3
AcVWQpaxQr0/Ru88jUuiaNppRH7cvb0zlkDNdgX+2EV0FVkIwqjy81ag6eWkW+hl7yN5FEL/I49m
CNl3OBRDfCG+zeOz/5BmMzhsIqcUJRGWA2i3KW+La34qaxLx2KqJd/uDSu7bGvrVEysisGtSCerS
OGwqKcMd2PJzvYDYkjZbTlobmwBqAp3Hbt3+U1oiHwICfX/hemXFvtZEgzcu0FL+JYbh++qwHRiQ
iSYFIg3sCIkXks5rjqSNnxvgwQIlgnPqF3j21CMKw7hKTJqvSlm+UmGDf9Yt1K+Vt0d2UOd6PgqL
2rJT+fnNrapXM/RYvPjLK8Yr4Kx9cib8JsLOfuhglF4DB9UlMpM5QGvWdPhCLK9vfb5UjjgqDXvU
wSWw02aL5pVNxlxVrStBbZ+u7HftB2YqCrHGj7EJBFkaoXHFQMkL1hCHcd96k7TeVwLo5bV8YFuz
Bagh4oNOoXIVLRDpZhHrKViKmqgzRQB2CBT/KN7iY1oHx+/RkBnlJfIb4OcAMS79NSfHnKS4Al+Z
06cm9cMtWQzvsnvYT4BzRI6VBVAOJOVlg4QxGgKbiYatHDcuBQujxFVIeYI/sQQbBfZndKbbal2y
hbSeoVo9tmkGM0kq9NJA2CcIvz0WJb/62NkmTSfqaKvlFQLYya+iX2x44yGl36buj18YKYiZgJTg
buaupgWGilbLz7qEhzH3qYt9qbXqu1oKcIl1y5RP7tTKuu+y82yc8cy5zfLQ+P/U3pMkJ5Pqxnv9
TZ3+K4ZEXbIEKww/06nJE1HxssnMHUv7dhcY3bSgyowH/UrTzlRJh1Hz/FOjdhWR705nFRvrinmt
Acg6tOvmMeRsD5qodSTvDDPAqJg4EtUcXqGJ2fHlTG00CdQKq3Zx0/cQnxzs9P62SiHvrO6RofMj
xY5Pii1wVYDG5d30O1ETekNTLl51DrgAq9QwMII/NEJbdKFpB35IjDfqSOf57SPei0bdGWNLB0v5
MrBaK8xuT/p1TdJTiDmrfirLP5EI9v3KtxqwtZoqyLgSsdApCC/ptKxnp3B7G4zcHguVF3BAIIf3
zuVP937jVbHH6dDvjpGM5ULlMb6UUmIjq7roTQ5zXKUib9Y+f1NREVGx7+CiZR/Svzs+pDWkMIxI
nKYOin7C/uPYzWvszd8+hgL9NRb83lBiJRos++6MwSNjxpkNUxm4PvUFdcoxzxd1C01En68uOihu
7qHcmNTSgNsi6Q0cV0O4cRv8IZagVl7/GAr7Op8ERY7zMyEFLuXw+RjqmbWxd6pIdAOSSTjgD05d
jZVr0Q3FpQ854oKE0hPWwW/MOkL8CvXJxFnI5WjNlbtwtvJbPrLYKfc7ovUau5K9lJkYYYxjjNMb
WARbCDrDvZQzN8r0BkWAStgoMW8wN26+jlnqIKyYZU+gzmrcgkuT/S0GI+Raoxur4xI0vVWrLUzp
LaD4si2pShLX7PIUed2ooqiedao/j1ZxTYhz4atglFE3NvdcyuaJFcmyNijxNg5S0Z++NFKDb/8A
MdA+8c+NUcuYuBmzGxHQkll/KvX/325nFjgQrJb98e5Dvss5mwQFcvQTV+ryn3LJ/Vttmxn+O9kN
WNzAluEm9ijetKfV/3rIrvr3lbJWWqc1gljuX0X0ChAcnA+x0DYr4V3yDpwiSk0e98w5akY3VFAO
amLcszUEcI3DMCuwTRMzonFxCDqY6Y+bTc8+h7IPpP+r/q/Yhr1p0U00RlRUzhpGSz27r4Y0pqf8
AttUpWKnYWusY3wNtbIsepovX3V9T2V4zmoSMUNu65+WCcM9M9G3Wyu13i5vRrfkMrukBdNu3PqH
BdUu+VK6nIB+JLKLMOeb+MFe4ptNE9bYWWTwwJg/sk5FxiC2cs5x6cKpq5hnUcg66TmvaohMRvtt
ZtvHvRUE+cWRrjk/vOY8kPmCyn3gVFpfrnzt7BMmP9yMZIumpMm9E4TvB0D3LoNmulk2mcUsJE/w
5RvtVDbvvu77BBecXYxa015qwE2x6XmJv9QUJGqm6RczF7jaIvvo/TU1w500Aowrr39LdDle8OXp
maq7AFADZGBQDc/jfjoeHUgKeFB1sk2nYVhMCaiFWfHNPGFcAnX9Tna8czb0crGFk6G4WwCFww7x
cHJjosz2QhzP4Q6Sat4MDHNFBtIZJBa1zDt0b5LwYB9mh9H/uHGSzCbpp93tU8KimCtyUluMPosG
Ibp99BJiOCR5+jEqXAPdE7Xg0+8ccyez78J5qm4+aWCobLjtv25ahw1oGtCa4UgO7qi1u8qe3Hbf
E1sSqIAfVi7kf+mUJzsHSAJ7lFe1MI0cT49RyTXeXRRRSKbScazHR2mrEpF74x8CR4zSb2dZ4PAG
wbJDjGdv00hk9pSVnpTG8IKJVwELWmyiorvGzU/CpXfAYuGo1V44VHZQQM+XSBE3xvB0Vs6/K3Ve
ol2nX2ES/KHrY135TV/j//mW0GBS2ONmB6BTFsMzhhVTI8XDQV9xki0YIdaqZtNq93ziyAIfcR/S
oe/QCKszJ3Dtvs3vzmxAWde1NtjdPU5cGY4dVYsIsPYyuxrkBlSZayWQuVhmn8b5CXWk+MvsnQay
DsZQpwa1IKkBDivaxC+fYA1afEdYt/xL+z02AqqCMc8z/Mi4Cc97GZVCjUcFD/++acDGSq5pWaDo
jbyPKw+9kiFoLu6KJ50neWS1VVZII4rd33vGUB+5pKaG7djuLhKQEhL2j+UIB+z4WNjXC3xuinO3
o760nLN9TX9utSMSo4YSKtf+VWW7WMmT+yb1mRPHPcWfIkyBWEeBJPwm4BmxeSYjweGnQwj0hrlF
n41FRodi1kOBi9peVJ2ZFpIEZAIwUz4CIb58lOW+Ua48lblYigR+hJXHo4AUSGrordKEqyYVcxGy
qC1UbZo92maqPC1qZpsvQf0o+tgtVZUe9dp5OdoW80R5PWp+aVgmrXhLTWq4panbRGEBmOmnYHn3
FIjZfRJJsbRZ0w4894/4R8bswW32bJiyj6Ec8JrjFXZ+MpG0WzvsfTE1LVf66BaY5Eu8fCX185/c
omuyp475gdaAJZPPzYS5WZVaqbOKBNw8eXxlNbq/M3/41vZJygxWel020evMdHkacqpRWTE3Mpyr
DojmNIpjeItAToC6rwAB7CBe7r9xmknXk2kUGnGjHKVkC8ReQgSxcHmOcZcRoN0GoLMDzhCtgKNG
EK1CyZAESTCACBerRu4R7mxpdK2LI3l07/20YNJ60pc/AzAdbJtn4e0XcU39fAzVasjJyk3IyWw1
VCPpYF+xCqhGnJvUML4dObhVjvh9QjeSCRXr+HxYDkdwM8F7pwV6FtB9EhnRbiwVxbhoTZDdU+2+
s2U4kSKU8mO0h+8yczpGmdtfWGfiPW7x3BkHQtch6Wln8URE6HWQ7DkKxlUcQe4rEAgZ3RDdKe5s
pmFWqhQVamByrGVodUERt4WSTOVSGGrI1Dwl6jOaQrpS/3EZlV1u3g3wEADTSIqIA9nc+v5r1luY
VpDRLwaXalTBucCCXKKpQBFhm2KflHuTv602stNLQM34EpGXiEYOz0FzzOTT0eiEyrRH46A+D15t
208Rgmu8tcl9f/p1YQNXLqaHaG+wbbqoTep0KJo95l9FWPHUtMYadvInNyV+QJv+RrxGWp8qf8rd
Dfl12dXUVzTpWz614iWgmKQiWxcyPo8fkLgA19HjCreA+eu0KjxoUP6HLIya9NePB0k/a9/LdGM8
4+O6BlmPqDfDZJpU8Tz/4DuC2jIRlgKEUC4PeMzqgb3X4JTe0BpEG/bPuU87qbjMDfZT6Midqv7i
Pm5oJDRJqReO6z5f5eYZv/4QaLMbvKnsu25ue2962oDDOkPhjHg4mq8rDva5s62MIz3h0tM1u/VU
g/Od40YB4uDO7N22VgswGliAAKv7N+tF/jBZTF+/55JjytZMXHNMWgMOjGEWVfDCj5pKrYq2gM6o
npcTcG6rFEl77ddGBT0zUAU/tX2ytJzli3suqSVbfjAbW5kl2EZaK35N5jRlI5PUhJirUu+tUFgy
sQyS0MhzqOXJ4lKWlA5tpNqogkSAUXD2QgNaTBNBhmdeAdLVmr/ORerc5h4RyAIxeabrGSgT60Gs
IuoHXSPCVTqbAs2Et0XHVWytA7EdddJbOfAWZEnEyOoUPYEEhsbpo5D0JAJaekVQe8LT9XBHv/MW
rvQBmUOxEWjETm9N1qUj8ilBkG4uCVHr+JZ61VhM0dgka2b2MJjOtiEVPxu8wtX45BlbNmWjzV0M
g450eREhI7PrAINt+fdtpRPZnEpNSzTn2CLmynm42wphq0mUv8gKXR/haYpLsySuebZumCuO/yve
ze9RHetys5hibZIYOkT47DlndwIRvXGfS0wq2Kq/5AawmoG0TvphKIKkumHaNzHudGKPkowFA/wB
3q7l+K4u7eUOPHqUtGZtFjClD9foRccWawuzBzewUT5tM59OwGdv7B/LVpD6LofjxloZ8aI0rvxs
I+viw1B0DwHkZnp+gs6a+T0PbHJZ1JKVXDrCwDRqM/ZaGwxlkezNAHY6/Z8lO1iSwKr+Y8Led8dW
R4RcgQZKX0fRZPcXZZHNfYvKRg46TRXjHMFe0O6UKoGd3ZiwvHjSk5XlTmq9ZlXdMqxjlOnzWr/7
2BA13ubUFGeRHw/rFaMeZPj/alY/R/PWFNIlyH9sJQdE6vnTXmYM1GEXtEv17nJSxlowt8QcN8Xj
y0RLo9ov6MTunmFeYgKl4STnIPjhoLjlYE2mBVa4BqUYmxefG+nEztmE3zQ/bXjlSfiRTvoGVymy
eCCDq6vnGUrA1pMW58L8PW0qBdW2mkRg16Q5aV2yyR4NEojy6dFqzE8NGzIPVhG+APTHyravwa6X
0Lhq6ntBfXErQ8tys8B6zOmN3flbxNeK270+CNJUg7Ad1qYJFoEUrnj/HRVw7VY6Uk1Xn8jl3+Ba
Hjrc50LrvcPFC8qKR7H+5Fw5lv6LQPt/hc3/V7l2Py4esXmXqNdi9JUvlS+7mB2/Ax+Ul8IWY8PF
d5Qi2UH9OMLKDSiHRvvqzKIo0vMosDGW2ACgiz93Sjb9gx/XSOKuZMP1k1wMYGE2jgPAvEkkvJje
SWwunvKlwtNfzGtHqjAi56zN0PlsoIB9BN+/FIHGBZz1QtKxCD2Lx+ETpYc3lWHHaxxZcjulEckq
JUgz8eAp9Urwqjtde8loGnF9o9R+mao2gu2pcjS5IFY3GOChYxSKhcdDqAgKLWysIb4F3Qz0yxk0
W2R6hBZATRGsXUMT4H+a5XzQIWsy3dvLl4XQhaLQOxIOPTERgBKuVmQ1s02VM0XNqrsltX3x39RU
JcUJVL/iQHm9GQKVU6G1dAUU8KVmdEhnFjGryo/lMStp7AD4ZTbbJpZ90Bb0R96sZNiJFL6PsGxb
hH7yYbHTBQRuvPQmOX3IPuqTYw2p3ryit2sF7buz9lSOHjswJwUrRts3VqD2kB92PaXutDXOgYxm
Ux+bWLX5mpi0uE6679ccW4Twg9HtLVcLW+QXJ9ezDRhAz+lGb4WBr27gzRbi5YTQawJlz7ZtEKkY
u/prN4Swczi2Hwsv9gF+bcggxbPZjaN5M5R2TsnosyrfzhXRcdnSSGtAL9qVo8v0oj3zMDHjC/49
x4naybjjEHu2pymw5J2b0WnSZRR2ZvU4pcPywN/JDZmvxS4+ZD9/bvdkrfoaNnMGCeWYH5RzRlnQ
d3LBBgL8BCt/LxjayZXQdhMKnFww1TOqMQw9J2MozXZZwS8wdIkpCycFPPx9d6v/+gYDkxraXuhC
Y70FxQAAmlX2cbVPdzE/zH8MP5xiJHy/aw7ltqK58xmahCNf1/nFXB6YpLMLZ/x77DXq5hw5DvCk
6ncNACy7fhuKW6fUlTCgJZQmhhFEulCgiCzI/fbtfaJKcWJYYKEcM65NgDW/Gf4wpZmddfEDtR1U
AB1il/gRuKV6ZRKY4r1DqoD5GIbJTq19l3X9Iing96f/mY7NT4qmxVfo8LFEjHzdLXujhLs1l/N4
UaHGwQfjLpCSE/UCvOzte9GKmOxBRUP4KGqxS64Gw+nDPwmmMDeQaWAfT2gVaXcdXd0Ik3NaMR0L
Tqdd2nD/hJEK/gMqrgE0byHv6wLzVqnnf6i1G6nD6soxI3w9z2ZKZJGl24Ty4O1Wdaih7a94I1BN
/RdNBE1l0DlLCrF4cpIcyUTxDv+pV2/gkUAeeyDrOTnZGEp3q0s2B/F3zWmgyCkaBY5mS/BRovlI
reQs2p0y0gE9xSqr+KLbKM3nwQXL0Hawvcimjgl5yWLk940virD7JQL9+YesJvFKivcLUqH4rJ7C
a4bx6qfC6Lpe5Iygbp2yKZapjbUzLYzMnukZNI8JuIy3b5o3nqDATxqPV7FAXXd56+assk/MY3pq
cCU//zvzlIubr/5erSEF+aKWNidW93w25y44AkGlyvQWQXquGmGyWDOeFgqT35+qFqwAVwGZ/GQp
cfb2iK2GslJeR1iCe884ll4bWlGUwfriAK5gCZ1mbJl4cjSCYOHjWnt+fvgmMH5EVys6RrxnYIvo
3w0J+wmUi5CIglFv9UdK+8A13SB0bZFWWWjwj0p12U4XL74jj0hCaiyKWn0o90vl6Ld0Mdmoa9gO
9vKELP1fq23CNU4UY9vd9QYAJTB8gxN9mH9xucuWMaK+QcbIMoUdIc1tuDOIxrF2gM3RbySAzXhh
OsLbEfs/C5hZYx/iLsQ1+f1Lwv4XSzP91TjJjg7z28Gd9vtWxOAE3eYxnNZd0YB52L+WORF3VPEr
xmvqOE8WJT0TNLFLVPf40L4NOGCpYj127nlq2XgbCOVB1Hhk5XZhAB3OPGbVSk4+DetRFCTbn+oZ
logh+ocEwa0TPtsHSr63pjPRc0c7bGK4Ksm5nvw1ASv3HfVZ4bJC/d+ftxVFf2qJzSgV1S2oVOF4
qHq6un8v0fM3G+YIAV7whmHy2/qiYKOeQ6ZchtuqwqZ1MGMNAyhfBxlISgV+XZSd7uwpcZauVCjA
YcIEHFa80XNtNLP8SztWXMdzDpkIPr2Nm6hxAgFOXTvCHo8MPCEAbNeFrzFPBfN3V3QgwH+5cHjv
gAxcAFVUSZF535ISaRpNYLSBXloLquJPL6Bb2olc8tRO5u4LeT09OFqSW4fIO38M5GU2PILI7lK4
D0RX91Kohq0GYtT0pRKctuPuYzm2HWdsecPf348fNNu81g022EsZskR3x961NYotiORxLDOH3ioI
diU70XIggBK+6LwJiKltiYBd+WMPGEfRfzw1xSLQwDtgrxFyzeEKnSVKWhbpBi3ccIf+h+SC53Mp
Gi/WAWe4FmY/eZOZUBKpM3qY2qF/6okmf+t95IFncfvXG2vOkVR69Jn7ywjdUtW8tFyF3wx21pqs
NFFcTDZJLLIb90gktMw2JZ/UFtHkQ7waX10yv6GvViqS42DT/AM/h97Djjut8RciLcwTllhVwxhu
e1aB11l3P/fZ9zzSH8JnhtA2F51l3h/KGQGcQwhaaFuaqWRjRDWa8iMgJ5COwGnm2d02TfYALAuP
Snf/Lg5K6BqkgVy1RxSvmCzNWsodNk+hqYqXe8N6cl1M7/2KBAfprH1+f1POW+vYka0nGCz0FCH4
VubPkfTopyc2pI9i0qgyK+80oMeVrUfL578Ch4KVc/GXlCUOh6OLh/6Th7CQEoxdZqkDfhy1YmoV
voB40VV9OGNkP/GN8o1GChrW9e5/lte2ysEkCfhXybxrFkTgJR5rD+3CcpJ48H7Hnf3k+cczx3ca
k+GoMG6LX2UfGyvmXV98SD2GVhezbno1hGWELuouNbSqK7DxmyeCTmHqieGgqnxla7sAWIEaT4RZ
jfydCwJce9auKM7Bq8Hk6+K5F9Y5JYck5+Bp0ngLlOLDpCbPZ89GiKQkzQGYv7LuICHOUfttLSLF
R6THFVGp3sOQr+QahvsKEZwEo6Um5yjnhDd+PsjZV19r5ousS1nWaVPtZsvzMn2UbeQ+xT9/DJBo
69VgssqPtynSfl3LXQwhgx8406inICb0i2hLG8YI7jXjpAik03QS9vmPDSvPv4LPRvJLAFH06kvD
KtYnVt8SIvTosMYgf9MNoiSo3lbNPsKzneevBcUP0WgnbcUaDAkfENW7fkwWN7HKnZkr8aeMzbtd
WYGJFyuo2Vx40mXSVjVqd7NuWPDkeAV9uHC0Gv+jGGB/so8N68a28LQULYAMEbkLyuYb8SVH054/
UXxhgYjOoUM2k2Xu5IShTYL+g+q2e3Y7EtSiVS5LcxjUCH94jwRR1Tk9iTURBccpPRd4g7K7M55r
xkQOOvWMU/mOxMLCoB88cR3DHvAgidAbzep0ttWcik3UDydYqvH8BtaF8//ORKbQBx7X97SqGUTh
K1A7fCTSZk4r3STCXyjlSVTJt3t6cdL4tiWBU4fF19ojHmhQy1IvjV6CJvrenU0xZHm535Daz2pr
RO5Mw6Otkuqci8VT/tbTZFcxnh0UtllIfhVagH4WtfXleqOpFWe+1et/uSsS8NT6NaegGehDBWtE
u5tOzk9dbFEsX7VyfB5Uv/ZKi6Yx9kFcG6a9/1yWlDxdKu1Hyg1M/mKEoNU85dic+oMCQacun6Jd
g8Q3AxNEgGSJ70zl1dQcviYvG1U22SsWYopA3QlhhSBjjnZt6comE95BWVSzZNwVB3BYLcNySypB
d2u/Qbn/bSOwF8Y8T3eZ7Buq1IkWPDZNh+ACKZPFfX/5pW5BFp9AahkqgKSAOfTSFsqUA/SINmn9
QYEha01QojUBZKkZeSevH3ZFCPcLP/iOyWNdgJVJkHFSoVJUwLqZX6HKxPV63UIlUhXnAHbVw/n/
0bk+r6HqENb2XR5lxI2qbAJJphEeEMDfcqG/REX/gqhZupKqsWjDgxNOQPIFaL/DUwxSwWSTohsc
Gf8kGviYj4IbuIqadfWFmLkOZp3GhZ+Bm8ZQYxaSPmqoPYLFl9aNf+peT0AB6cNUxIRh5GcbkK1B
fwJjokaDEMwxr9M75WRXgz+QkKhbKevxDoaWpFjkGWggFDS1KobjOAXpjSTUWwdC8gu8ZENNnocJ
zZVdT0dVfTGgwTZlzn+DAbCiu+/VaY8W8XxEyPiO8z+mSUttDpuLpOIfDQJmqnzNYHxBqcT0xF8E
AS1Oqfx3r617A4R9TZd5cozTKcriV0Q6STHcg7srgX41eyX/+hAWLn5O+Dkw24KQPjde23PsUgN/
kLLM6Df4Unz9gJtnGRVbn0azKhegyHTnMwmqFLAbaNcgYYhkIURx8ybcpYJpE04qldYKu/uJf4Ge
d5lPn3BlGMXaMx11PG437VMASJFhITml0lVtjpFfSyj+6bqfSH9eGyVO4fUHS9Jjk/bghzP5Z5un
fs0yMXQY7rDpoKiYv8kQSsAO7k8XfU4/8kzkM90dwKUE/PBNuWcar6r2BJ284/XeDHhDB4NASMMW
Q/NqT6tkyS0Qos8ztWIJ3d0bc9aRXXQOZfkQrSVhi2KaVR+Vy17wIGvep0P2VpRZQpnIKU14caRh
0bZ62/Wo/fvS1Nsyz/txCfBb5kzWaTDdGEVjG7Lju8uhF5FmJ35k4m06ppFRWcQdBIXkQ+l1xTaO
oVSqeZQADFkKdU8V5uIhF4Y3iciZpGDf5KaOvrxgX6x8AawhZXiBb/+VIPJmb4bs0qvkHg7GUnIw
b27zCv7h0w7Yf8Bfhs6iIQINOj4Qvc8LWF+ybAzcMhUqOo8mJwAherTQEaO0weF9KfwvUYPrZ8TW
30XRxs9kU9IwN1A5YXAooZfq9rTqujZiDxKkWXBN0sc00teNJ6BCj3hLSur+Crc5+JUbPXv5CFdu
8dePhmP5ksATl70jejxWG6AoeM9hYCZyMmy8NbCoyzdRVgQQ9XSZKZ5KsxSrjlOTXJUCb7pXYfgW
XzfPiDRJunAgRI9AF7L54w66Ee8Cykl2gcNyvKNdIDiDy05Z0kXrSJsliLc3OOrL4K5R1CuWmdjA
sDr/mszLidMb6a9ZYE1WzrTdt26gML0j8pD9qAXB/DKq8SA2Dp1PMgUPpCX7mFEcAKtZywKtADvn
o0j8uNfmhhdWCV3Jiys/KvKQ9gxUHa79uSqrOY19KwvrUaxQTrkFx5kPqJoRXV60gW0twNRyd1pr
fIQYohty6ynMTeWm4+f6kozE/2STCAVtVOWRxVjXo7FGweMsmZd5kQhpWXZEEb2vGH796F/tVFVU
toMKYq9wlRu73TF5dxuHf3av+vYJHLDqucNfvsdbjKZYDV64Eno0BzvdVFn7QgKCuOFlR3stQ80z
ApfT1dbzmnJ7Nvw513Ch/5up/Bd7Ei0ialRfBNBZVE+wA7sURvrvcDLjUiOLgRFgsmnEGIZcdRyJ
FEJrAB20UFZRAJhIejI8fL3GNgRn8+Ybd4PKNmJi7848uK8PAoTzj/Lovkh0ya8rO9UZo8HuNYkF
hmrWspQ6xzbZV6znaEedwAT3lS0fION2RpSAP7d9l3kkLOyS5Ge6IC+Xe4KThGISNZikbCEWpRb4
aKLmAu9swfJkRRP8wXAGaCH7iS53q+E3R51CTogcsJTXp4yw8j6iYqImQt2Q1HOgsEBoIoWuhoca
3RtcIoSMF/al+zs0Gtg++rRvZA3JQ9uJNaungLsqcsK7Sfivkuzae/CSKf3yIvodTGauZNclWwAQ
y9aoVDmY/ipqMh86MD7bSj0LsR7STkr5aLAseLnZ7VqF55k85pGjIRkZghC2p7rrz59X319YUFnT
7lAld4x4+Y2lJ4BOUT9ShJffKfj9wHaTaH/HWuPQjNFSsQA316AtCP/H5NBu41NWvcLXPyau0AqY
Ja60QRQeXu6iAH0zqjJycj4vO8hXe8UQYktt3t9xIRY4b6k0gyAxRC+krRXrUD5Dt5cYLveadKHg
Ik52582IpsZaggm1bMuZVwJFDiIPXLVD14xMKPAQ/kkPITq/PeYL/GvZyNizPdYvFM03lO+IAoVO
ibZig/Un1Odj/dlZzvozEPhwiWs9eRuoyZe3CZNCUyub79V1SS2BfZbMRodHThqPZAe/lb4QRshg
1ECLwTraCiyc/iHn6fdlKdPU/Pe1E7UteSy/NP9sU399HxM3TP1/VroPux4/KneStkieVmfR+alz
jlQMPaJeNdSINqjoYlACpeqIFt5SwG48EHlyr28QDpXiU0PTzeojwDCt5Pmajf58khzwhUFS+nnX
7UuTFgdA4DUeAKChNAgKLiNC9Ld+zGzZU3llUDZjQv1mw9pAPRIKY9RXdF03UwcQZ5Ay7b+doRVn
5gdMstofEzoKAjsSNse7i3iquQIFYq9laPUwgaqpMAuPSVbVJoiOCvBKu/qrTKhowv4WXTTO9i/M
tGlLmAjt1v8ptDMmHv1idrDIK65dXkF6zok2aC5h//MRLxF/LbPoBK1dTanG7n6BbcxHHoQ4P7nc
4tWvFG4y4dpfeX86+KyjV6GkJxGlIgKrgGko3uoHErt1pVSyY1lauBIm9H0gx0yuo1ifS9bXoC76
qvk9t6YSU7rnuStLQACxMcZbQN52NZkSrvRvrhAwsvb+E4tZ0QeDNqxlHpFcyda4xuAoVuJ7M5ah
PMQ6ktaR7Tsf7C2HfTx85xwL+IsVOhxNe1nWjQofTFn0FhdsHI88o1tqZkEljpAtMdMLqW0Ha4BT
kpGZ20YgjvhowSxHJPHIYj4SPc8tZHcFxhKhFoGkXdS7O4EeYzh1fRG4pSixXBPAQdQr2+RqeQYE
3cYjiuo75lQCWs/kndVo9bn2P05rLzLyHZn+VXYjNCbX+G4jOSPUUkAYahaH7NOdyijMb+7aq0I1
2SJkXSXvSMF+tMcLuHWYR6IdDpCrEW9x0Y82wL4HDqTTCP8eofI5etC6oMhAM9Hn/xQU5t4CocY8
VoHbHU2V4vbqU7vYDQKqujrE3pWoq1B1HyxLcbHr1oKTYpLmvP/PCvQnghK0Sc5lokIJ4jOXxu5i
paoMxkLQRXaTWCGbnLsOd9VbPKcJP6Dr53Cu4ryYzXvJNZOWS6Zma+V5JqY9z/pHnu5FclQvEmcg
04n0B0Lm3VnIMmJOOcz3w3sTGbDpo1xB9yyThKR6vtj+Tk02IZ3kpMhRMfvZJAnS+w2tAQ1oukqB
gaYg6JwQhFpQ/ZlQLs1aBkOXeRP9PxucS4fUL3YNrh+5rnGlCyzHQN+wgqSyH6b+8woBtUZnq9DJ
D3sPrHygPB7ZeUWD04qxkhJ+Iqy3O0h0qslB381TiaTLpi3nPhnwGXfOy3PJC+7jwY80dHgEFsG4
2xVW+UGFPE2I17tVRDj0e297YBj5NT9iqK/mQyf4sDpEzVMVKij9N2B/tpIKgQI6VtErgDs6ORii
rH3Tecdpd9WApOAY6L2LPqjPCragkyaBGXsIWPqSl0fnYZhzs/999+2/73pt1TlxBKll3Cxs8xOD
Mm5NwwG0ktWW9SoaqmMAk56X2cnIYEttbdq95qxsbUOheFJDJNnDM1dKVbTnI6CEe/CVFf+Zg6dj
RiPCIjOG8X6hw5unKF3nWEPuERwhhT4PhLtIHydBNChp9sdNazXphZBXu97eukVjPH1r8DJ8OLOf
QXU9ddghcap1VHonDcgnN7oxXAwzSGL2rca0OUkUQuIZv21qZZ+X5rMvQmKyOr6MPm7TCUy+uCy2
F7+VinEhJQ==
`protect end_protected
