��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��[J���$IJ�@�� ՟��H_�$=�Bu�h��S*����A�P�?��d~�<k��KL׽f���������-�p���0 ԥS�W��3p�_�rq4j��N}�JʄY�Tcz=�	�P|� W
E`-U��������3r���#S�<Ջ7��X��e1��S�PVw�}��X�*��j2�����$�a�kf a�r_;
��.�US�i�2ʧ�M.�6��y��W�����dcu�vJ�؜
I��QrÕY�ŤK����#
zqu��==�[���w�~ӪЯD�DH�����U}m��������lRԼg�Xj�
�N�Z� B�����d���n�m�|������r�~qG�ʈ�B�I=�ʐ�8lsw9HT!�_Dn���G`w�D��h�������&�#�=8,̟���_J��Y7U�HQ�o�N\��&|[ϲ����[�Ş~s�0[���W+�t��¨�`V��}��&ץO�&9���N�eq����-��A�F�Cĝ(�; F�<M�,Va�p���3av�X�Vw�������4QB� Kz>D(�_ȧ�#�W�"�\Z�^ޘ�5 ��ֱ%��k}?���h}^��Z k�4���v�1^�ʙ��ηU��f�J *��.�^c�� {����e������8#??���m�Me}hH���[�³rk(�k~�ү������tOۅ�I�����`q��� �މ��[�%���w�������q/����` �g�i=�6�d{�������W|���u��_~q�NՐ�g0ϴ�% ��T�͌ �����"�������l,�|�t�c7�K�Ի�1.Ƞ�1 ��1��>H��9��n�&{oJ=fF�	�[��Y���R�����nc�g����.'E❹A֥@���?���E=�%���ru�la,zyRa;��<�{�/����__D��`��H1J�/F!5*�j ��~�&��\dm���5't�hN�S+�G�(֮�^^���'��� L����
�?ϥpc�Ɖª����$�-g�:�����nA�c^᲎��#���An��#�:�
��Y��?�����}T��[��%N+�<ОV����5���7���D<S��B4ϫD���6�Z(���"
bw8'W���Xs��|�D�%K�Wo6q?��)����37ܳh�w6�&Ǹ��9(��"��������C�$k��7

\7Ƀ/I|H~�%�#
��I��SM� `aG��WZ@S��kjL<"�L�X�������~���	P��ҝ���^��4A�4h����G���׽>��(�p�p��Q_�z�%�����T��筩:"�`�A�J��=�m`�� �^��!�ԮL��� #��<oË"����p�	�4����LvC�)4�LG%)�Q}�2 +�g��)ѯ���Q��/�,_�8�M�gd��".�g�6���5v�`L��3���Y��ǆ�[k+k�
 D�*�}ZC�В��v�mz����ͽ����Ѐ�D�:!�'�3�,��r�}����H诩�u��J�|��U����$��4N���k����~p�;�(�t���\q�
r����VE��z,��F��K� �x�جȨ܎�n��P�.�^	Z|֦p�H�ۺ�j'�zR�ktv]��q$���."S�A:�Z+m~h�F#`��e��P�F7
����ͼWo�fk*�� ��d^�����Ұ]�:������DÌ�zs�]H��W2vU�ya�����պ���]*�A+L���\6�P��Q/�s�^7<C��4~>�c��Q�FB�Aj�ܱ-����p$�)^�<p�:�N2pRlꡏiX$�:����%�6ː����B��á˹���1+#�e��J�6]����KA�wJ+J�[6�ױntTM�m�$u�#�M��(�T#�_FU�^;�^<�a���}���ߋ[����ٽ�{�E�� �pg���"P�F�hN�l��^2�[	�-�W�"t�A+�%0q�=Q�)!�#�odo��7BԆ�m�H��� �S��Tv#��K0�����m���c�&@O2��J^RVa�I�0{�����/L�jI��	� u+��bT&@�Q�++Fisy�^+6��V�T��jτ�[���59I� ��|:�$���V���l�4U��6n�DL��P��E�I�u'_\h���ŕz��HA	B�d
�/��<KF�B~����d(��T����P8u-}�|����+�i��;ðk�����x����L�k@�m��#Vg�/��L�bά�)+jS��q|ʿ2
}+�h�+�p��w��8/��s�{ā�/9��ʴ����nc���=�w*}D`��+�>r' ��
� (3�U<��}.z
ٌ��#R�f4!WZw��K!|���4F
2��>�m5���$9�ܔ�CRuU-_�� u9�L,MD�t�u%Q�]l�=�����;Wۮ<��m���� W��6[}i8����Fķ�h�4�ډhO2ā�L��߇	y�ф�"�&����\Si�8�P�z�3U�g�<Eênvn��tQ�F����K���>�-ڃ~颟�ܵ�<��7zP(��aӝ�0Ҩ�v%������֐�(�}HÝ�Nt� ��)�Ŧù�տGUS�g��K��J�$�6m��=Ov�ѪqRi�2�G ۩�ɕ|�P�ڿ�|�&���_f1�a������0�E��se�3���xk1H��[���:�#��� rf蒚�LEӳ��J6������^J��)�fFmG+c�'���6�`��3�X���`9���R��X�X+?L�bZ4�0I����u����ʍ�,�~��X��3.�V:2�v�[�`��ɼ�_���R$6^n�e~E�N�v,�+�MY���d��z$J9竭��e؃���|�d[;3���q�r��p#�17k���tz���1�_2ʇ�O�v�X���r�I��c4+���-&�`E�۩�#)7�(����
�-ܟ�nsQխ ?L�.۲O�*��s��ș9�� �>�E^����f�=�C&��n�w����̓�x�\X$���a��JZv�{{Y2G���0�Hv���`o��[�!�}0~��X~@��Ȣ�����$��4L�> &��p*�MA�1ZT�E�#{͜��׺/v�t�!P���0$]�)@��պqLziT!�f[`���0�9<$����q=���u�����x��I��u��:�>�=���{�'��0��WŞI��'�@S�$I����E|���V�ཌྷ�ާnX�u�r���������j>��X�� �xW�W���O�4[��	�Q� �1����58�ǯm����G?C�;�>�-H0�3����Ot�%v$�ŉ��^HT�k�U^�s�`���G	�l+&��c���ô�wSu����=�􃿠���r���R�?��5�`U0������_�d����E�~���G��՝�e���X��7�ю�xOT"�{��>�����@S��qr@iѡ�"O�9��nW�
=�����2��7�i�[y\�u�eL�w
��8ӟ��dh����+~�,hqs@/�Y�hKL4##����}�J��$ڴ{wD(�"��z�I�׭�GZVT[EH��T�-a���d�*�PJ�-�XX�����+:�@��;?��n�ײ�P�Y��sf�9�R�s刄�#�?�$����<�;���QY1EN-_B�2�sng!�˺)�FP2����\����;�y�R��_�R{��&�qu��+�u+t�Ȑ(�x$SB�qi�+T�*�2� p�;��5��X�PԒ�u��S{�J����_
�c������������RuScw��&��}G,.��v�������6VZtr�3�yBM� ���\:�%P��H9i��Y�u{Gx��Lv�|�*n �����*'(�b?���A���/���02�_aa��������,�7�+�7n�3�K�$g8�l�kr�� _�MD�L�X�	gw�b�I&��{�AV-Z6]�m;>��WU�{g������DI3�|��[��b\x&�&�;���6s^���ĩ�!��N�l�q���C�"]ky"����t��,��6���PJ!��|�DP5_,����&�F2X�:�F0>҈�s�!8��-�㚳Y[�vv�B3���}�{ϣt�z��o'�y�I�v/wڧ�]B�ġ]�!H��1<R9k2�J<�g�`U��
ƻ�//#���+����%�s�X>�פrm�.�'��e*��6��u2I��2�1�[G(�~TہN,�SD���|��`�|��W��h�H�h-��t�
#��_�O׎Hܚ`�^�F�]�r��4}���\�A�R͒Պ���"[��1�B������8�4�F6#�ȸd�.uF�N�>^��%?���e@�����+�
��X�;׆]�h��>����a�N�?�����&��w@ FM�S�?Y�	.}O�<�1��./�Gj�c1���N4~�o�a��K��1Ȝ��N8�=R/7�;7���t��s^���T���z>p
���?]((/I�^ת�<��c/������h��l����r]JD^'���� �nU'�%2s�RPᅷ���h�C�M8��˲�����w��b����!�%`ɜ,x(��|��:�*�Y��F��7Vz���o-��2c�`�Vx�����U�L������_��O�a�y���4���0l�� �/�qd
���u9��+�Jx�]��@5I�(E8ښ�92�F�&�T.�����|��a"��²��K�9Co|M�6m�3H��7��!��U��Ær�{=�R����ּ����:d�(�2N>"�!
.���>D|��t[�k`>^���|�]j��R<rx�S;z
zN�����r$%�ے5�뷏=�]xݎ63��n��C��E�T��d].��x7م�1г�F�6��L`ӬtU�6::"1\%��z@�w�f^��~Yɀ������6d�=�YQ�����r���M�YR`B0��PܒH�" �+8�p|9��o=��#-�x������� �e��qu!��Q�R����}ω�=���a���.ɍSA7��G]�/�g�y�o�*(���PF����R^N�-���Q��U�y��N��Ě@�J5]z�_93>�tr�����@M�"+l��:��#@Jg|�#t��՜��D���}$�}+'�cĩs�C0�-����㈟'��E�j��k�h�g���j}�Ne��A�;�Aʒ�T���C�l�~�?��p!vj
�VjB��|�_��1]��wQƯ��e�p�F	��mjU-�A��z[��r�e'�����B 8~��E7���������po�� ���D��|��mf�?ջ��\Ճw`�tG����$LG����-�;�4�Wj�7���B����ۑ����F�Z��"'�)���e�-.��UKcf6��ۚݼT�����|U��8l��;r]��CW,����¹"�)���7���P,O�I�@��2��L��b�;�$jZ	��0X7X^��ks�ξ@WC�l��Iك��zt@�<�1ԺdAnQ�k�+�O�-3�dDF"z0o������������qenWX~sW,}���'D��ccϓ��J��4����ɔFi�°k�}��t���
��m�p���j:?�ܕ��׷m9�:�i�nĖ��NyV���r
\�8�Qj��p��.�Tu�كj
���ߠ�S�fH����ª*P�^'Բ�S�,aw*���~�>���/���4�X=�N�X#�H?.R��dO>^�)��fFjNA+�9B��yŃ$�]i�$w���}��`���+fHTГK*_��z�/7=�N�rS��(%è�̓���]s�QU]|�l�F���z�����خ��cF� ����6��������16@�W�gU��T�Ik�Ro�Ҳ[���[�颬кk&r��n�����b"�	�}�|,p;��J`"�hR�KS�����͠8��Ȃ8�ԥ%H������z���k�5DU�Z��h�YWĕ���_f�5L�����K���_�|�3�����	
kC�Z5
�^�0 G�e�� `o����PiT�o�Cw�f]@(��3M�~�.��e)�N�'�*��J^��YOMG�8���,u:��Q�KZs���o�ɴ�?H�#?�y�� �ֳV�Y�{��,�3����U�}�=�z�����j�W���Ҏ˲u	`Л�ؘƕ'$F�����i�iLM���zP�`ma2�:6�d":i(Z�̷���i���?�c{�:���>i��`I���^�#7ؑ�(����~�8�h����{O��u�),��$0�X�������d�&�bÆ30�(�aˤ�L�R*��ӟq��`��2?����%���MXޫ��<Ɖ��)gO2��<9�(H�=�cS��v�N��#�����r���܃��eڃ�� �J��^��j��R�vJ��g�Uf�9�K��g!����0�\�i�Hl�tv��Y�_hG�|�b<�-�^�B�/�sĹ�nРV�;TW�Y�ͺ���6|�z�pTd��0y�5N=W�־��� Q�EH��+�������b��\�2�~�@H
�g�(ÏpP�1����g4��&(�Z=s&J���{S�6���ީ��l��Y��*1 IM�lv\�h�|��q�P���0r�Zd��' �n�/G־J �сv�P�8k�zwn���-�g��Q�t{�`1�^��wTj0(��6�l�igȬ�g%�E�L�3(�Q�_"PJK!R��%� `���}|m��fx0es'�_;�.�}˥�a��ί#����������6��g�LQ���9�)=� l���c�K��=0Ī�h��1�_���~��%2�X��s���6w�
e`;$�z7������r2į�:���T�Pa&1��>٫��W��Fc�7�ǿ��f�Zi3B����sx���8���U�y�Ul�b��X��/9��݉��4Z�s�5Kj���C\�����
����\�Hh��c��x�δ�	�]�ց� A����6�6Ѯ�-���gG��^�������x�Y4�`2�i����m��O��dα����q6^��Q�"�3I�&��3��PŻ��4*�
���q;�O'tO3'�h{γ�/�dj�E|�Q��|�uKR{{IŘ�%������.O�-B�F��b�Uyf����{���YD�z���:�r�U?F��d`;�������|�Σ�<�����4�r=RO�y�A�X�d@@ w�f�g��|�>m�fen��QEO,nu���������gH�_O��a�PH������܍���L���5���P7��"E=쟆M,���
ә�k9[:��+�L�y����Tǩ�B�kK.��wk.�b`6�G���9O31����ztz�����hqX	V~Һ��BD,���ڢ��2�9m�b�^�$T1J�������w�u�YK�Jl��Z��4�9@���]��ggJ����vcp�FZ���c�RV�Z��p���	[����t����6,j��'c�>QWo�1�@����>����h�^�8'	��|/
�y����~u����8�839q�b:8�9�9�+�>"���r��P��*�C�8H��Xlm�o���#|�� ��L�ެ8[�2�ћ��y+�IF���y�O��/cڏ�_�����
	�^W�Ϲ����bM�,Q+��/Y�ǧ��8C�m۽�$�:u�1�B��n�v2����l�sz����`rrU�����HX�v5�e�$"-�jŰ�[˲/����ni��Л9��D��Y���x�UH�ο�H������%/:Ri�Euue	�F�cԖ09���}לF�YC<>y|�A���p�غ�VJw � }K��t�1|+TӢ��&��Dѣ�rPm����9�#���Ӯ2tx+�58cAY��nt12 ���� ��ke��?���Fr��g	�g�aC��֋!�� s���E�F�Ъ�*�)~�d���/:���BR_��S��D�z3S^=i-�&b0��tO��5|�P�6�:1E`�&��q��cG���������Q��Դݲ�O�a��DC}��k.�.�␼������5��0�j0.Zd��!j�=��G"]�����rc�ɧx.G�.F:�~���e���u�:|������"6�<�Vݡ���c�!�$q�4���c�//����Zg��{6�c�����z6_��]يi�V��c������й��M�;�bDDC-:�[��r�̖�+�p���8Uq;T]�H.����Z+(��Xkm� }}�G.����G榁yq��|^N��`����!��T�AY~�LH��JP���
��7d�~�YSE���KŞD���������7p<s��6�b8�a
$q� �f�2k_���Ю�HD��#����(WH�?�.r�/����E
���x��Z3)�!�@��3
�*\�)蟈�P�5�_�������*�b��f�ǙC�7�l}~N��銪��,� �&Z��Ίi�kʂ=z�sHvz��KQ�Bg���1£ɟ��N�0�4�*����5���>J�#���1�I��E�)���{���I͓uMAy��Or\���Z.>b��4iB�&�9ڦͲ�cտ�H�?{F	|�z�ވ�=�[[r[�¾�I�$\���q�-}�V�{��*_� B��K��ۛHyp�01<_�Y�f�TĖ7�rp�o��k�F̟�63ZP�"5�_	���{�.�x������1F|��>ѻzgp�I#��^�i�X��TF��� s��VΈ�����+�u�s�t��ƅ�կ��݋��=1G�Ry�� ��#�����*sXO����m{:�u�|�:n���u�KԦг��E�;�W��%n�}U�����cvۻ�t�S�ii��X���b�p4�?��0��������:M`&�W����7���z���T���wDP�s.��}��J�$�WEJ!m�!*2�<	��
I�w��ߴ|~;u<��k_~SV��p�NZ�,Ӑ�f���IO �p��46��������/�L����{uW�����'dDǜ#ӏծ���f1�I_��YiH<ɨ=���$޴^�L�Л�J2֢��Լd������9��1د]d���	��SZLk퐹��X��z)ߝ�5�� ��]߶�Zcs0������`r]�T�h�6X^ގ�ة7�.]�p�ƥ�!v�������mꏑ>t�k��/h��9b�������Խ3ՕQ�r��w"�:�A�X�B6�-��O��B�����<��о_�� ��b� `�v�"/�S���0�i����j����ӟ�*���D��xd뻰����o�n�o؞�|��X�͎�i/�z�QF�!�q�@\�B���al������  S�3��$h�T���\��.�U�N5<�A �- ��ւ�*X�9�QM�TZY��s����� �9�k3�f�;���]� HiBX	�wK�A���S���nQ�p0'���1m��n!���_��5i1�=e�:v~�6l_����B��s��������%�b�f0	��*M�:�ei�����O����
n "F>�c�}��(V~KPݒ��|���-���:D�_��:9&��_5(�r��+u�"�0/̴�:aDw|�PƎ���uy^h ��,U�`kb���nč3	c�1��_&��Ԋ~���ڣ�!����<U��Ȓ�Y1+ڻ������N��^�sB�N3²E�		v@@�?�t�ԇ�8�S���\��)�:P1\�D���� �'*~��(�pzǳ�&�
�a�vHs�*�xb�k��s�����Hw�xԪs�N�?�4�G�-w� ���,B�Wqr~�&R8�1�� ��r9��~v��a:6=Y�����ROw�*Ql��x|�6>��2�\|�$F�,�]�����v�ܸ��n��&ȟ��ʀ�y6K�� �#�����\�9�ı������W��N��F��B4�]r���=L�S!��Q,�&9��m�@׃X侤ƭSN�QL	%-�q����e�Y�)���?K^
��~������_k�	�~U	2��7h3��M�{����K =�ΑQ���ilx���i�¤:��(賠]��42!"�K�N����W���T&�L�F���-����c5g�Q�����S����W�
�ⲭ�_�!��.uYo�٧��Ȧ���������r�`��)����LV�}�y����wzC��JP�E}Hq��:Ed}\Ӌ,��'_�kVQ��(�+r;��	��`���%g��^~Eh�r��l���1��m�oyҍ)i�(���f<};�v�0�щ�,�(ߢ;�Z%8���V��f�K+��P&4�F>��_ֈYd��@�P3Ut#�Jn �.Q�+nQ+]]T K�>��*ns�� �A�á z�b,0W��<unN���]V��J_ى)��`�T�1��W��\]��=oq:#�yi�W�+P���ꦂ:�6Ӥª���G	�>ʫ�����_��&b]8�( �}��=�0��^�iW/�\���w��֑e���bܲ�7�l��f/l"+�r�zտHi{�g���Kվ�@ԅz�1���f&��	��ѱz ��B�N�?1ʻ��r��YR=Jc���&����]$�^��>x" �nh�D���z�t��봄�*���RHe ��9�L&�h*��S"��ӴQ��ۄ�֩��DX⼖������(4O���]�f�^�L	����٦����Fe���Xѫ�%�W��!⼮:��˄��?�*t�g�g�X��ȒPy��_�,e��T��>�`y��꾠���\<+�>ly�y?,ҋd��S**wJ���u�v25�(�[�OhNs�o���6e;Z�}Lxs�K�ۙ~{+�B���ͬMt��J���fSq���F=�$�fSl)������C]n:yd�)��U�Fu%紻�T\<�n�9P=�l?z0z��7	m5����kz�a]�Psߧ��-&��R�����?&�.'�e�����_�ځ!���.drg�e�_�Y�q �3��fYg;�V� ��'�]��m��tn��z�+�����wat��d�;�믎�A�9<�7�Hp�\[�|5��օ���G�]��BH�u}��9�pV�z7�$Z ��<�v�l�ڧ�M�T���;��_�a�9�	Wp�Φ~��-�bbl;ӭ������#��Gk2�-��/6ᝃ�A�(7���Bjn�,J��L��өޣ����N際q���Ð�$[�5�F,WBO��c�r��k-E��?�Dm	�aA���)u���^~��^�(���ǩ<#^ځV)��H�(�Ϙ��t x�g�A�M��Y6� �s;ׂ"��m���Rp�E3T �]r�a���ܔTE�����>.�^9�c����Z�kepGc�1�C�]���KQ�|+[��E^�apf�#vn��jh��#�.�V���_L�^L�7�s?�$�s`�(�����g�D�]z��t�4#��M� ��	��AH�f�V�w����6I*5l�����|���Wq�(U�|�(�u�kRI���=�(	ui#�6)�1��Z�볦�Ҷ�~؟��x�A̗�b�d���]�L��CC9�MF&�����;* �R�F6�J�@���I���+^������́�sj���8�(��T�h�/o	�ȹ��Oļ��Z��m��Ƚ�P�$����tm�⯢ƿ��a[�lE�#��'MUH���x�f�H��
�wf*_r�]t T �5��3'z�ٯ;>9�KV�[w.W���c����sʴ��pJ���f��Q����=�-P��mzo�C�Ū�܄zǊR�go[����=(č}�~m���T[O���ĸr4�Qd	�4V��+d�/�O�{0�پ��-��)�'��t��1�}�QH��`+5��pX�Sc���-5�� �AU�)p1�kbB��H��l�y�A�0\,��"����Y��?Js�#V�>H㧳�'N�0n���/���}�dg�A��kʇXG�8�운�Zjo�$SIF＜��	[@�1�D�I�W��v$%B�Y���<�(��� �E�T7�ir�*�f�K�j��.̵3���㪓��޸iktT�y����}��d���s#�"�#�k`q�p��������}=�r����V���oq��p�\�c)L���n��2z�s~$�(�xl���9Ѽo����聬��B����_2��݊y{�L6��'�o��[�ͥ����3�Mj��E0z�^qzg�dSɋj���~ [/�!�6�c�Y"|ȾE� �ŧ���)+ݖ�-�@�Wdt7W� �9?��k.+��"d7x�����S�m���� ��%xN��2����{h8��7 F���.���D[�3��R�7i%g�u���U��lE�I��t����k�[Z8�
>���w�YZ�jS��³��2����0�[a�֖
L��p�������}eX AV�!���-����
3Np��~��s��3�o^�^��	��^j}ŕ�p%(����8t�ͬ�ւ���V��X��ށX� �7[Wv�¢`��A�~�Am�2�/@ �o��J��I�k�m2u���Sv0�6P�Q���%tл�`�k��|#k"�ԃ8=6nk6�K>>!t�c���r�e��A?�>Y�"҉a�}��מ.C�ί?:��������j=�&j�����Z�ʈ?Tf��H!"��[2
0@k���/�ŭs�;4���Ј��y6
ؓ3�y��,3�(ٵr2ӓK�]�t�1 �M��uP�*Ϟ`lMg��F�W��b��
���9X������W|>�ў-:��I����]�IV�m�e���QfA\ u���,���h��ǖa�A��@Sv�r\xz�*u��M����ϗ�@�g�5��%p�y�a>]`d���Q� �DL���#��P?�^b��	m�}�4'���T�
��WGkik�c�΄SR���}E-
�(�g�ց�/�$���6c1�&5�6��U�$�mHº���a"�v�U�̑�H���r���!En��r�趣Ĉ�<�,�uP���c�)��X B=��\�K�f�P���]2��"�CA)��s,�R1���J�\{R)����NRl��`4yEHi��H��7��'2�ƿr���uMw'�}B�D~N����)�g�:�o%��^Ƹ���N��ec�����s*@y�Mȝ���|Ixck_�TX�qD/��8p茨��b��d:����E
̃p�^Uav��N��T$>�.?z.RC����:/�p��(J���f*�b�y6&B�x�F�;a�a->�"�
O�n��E�fOP�+) ��3pnÏ�5ǬgC������J�)aU ��R��ć�K�~՗d[k��Y��,�͠Ș�.!���� �մ��@7&�Hb�dR+�?@!�ò!
s�3��&!�4d`
(Ts�N�ߚ��m�@��L����g�ö_ٲ5�OWmv%Ue^�c���ȉ`�rm� ŏ�2@+�������P���6����i�e3 lv¯^�i�[�`j��8���0O�	��_А�v��)�(�Ck ]J���y`uytOA�zw�`�Sɼ9��ި���}]������Ԑ�:+�#�_���C�]�fq+f?��W�̢�*<U1����Rg�ѯ�ު(d�EЙ ɺ���l�*���B�֢z��1���5�J�ڽ�M���^�V�4g���J�?���N�9��`rs�P쯗���x�7>�5�01H#������Q%II�q��ȑXu�k*�Y&��������v�<�G&�%q�V��R�r����9�Kn�q ~�;g�X�r�p\ �3�2O�f���5���y>h���[��V�+jpV'~{�5����t��2ǳk��0��E���C�,L	�%w�q�ti4l�ߖ�B*$-�l�	}0��~0XgM�qO����9�P�Y#Kk�ҏ�Y[�u{7���h���c9֝鿄����6�4�ţ꜂�r{�/%w\2݆���{z��,���j)'�J���j�olXxf���pQ?�q3Bk��a"�C���!�@m�5�dGC�Yf�M:������i�8�����2A8�{�Ȥ1n ��ƾI(i�����r�3�jv��+w��t�O���A�vH�Z=nb:X}�G�I�����>���="X1���տg_��J?#+0�_v�dȆ�REHx#���<?n��W�y�{0 $?.�y�9�b�]8�\bvXJ���-@�Z̅�%���=6�3]��}�l'�>βw���7(M�OA��؏3��:8@��s��5Svj����۸�&O<���^fҤ����_�x�="{�iۺ�� �����sL��[���Q���rI�/��2�KA\�!��������j�y����T�A�X��n����6�5Ofh��=l���E�~#s�и:})!_~�YQ�`�R��_'�QzVq�A�_��Z�l��%h�D)^̠�1��M����9�Jāw�)}c�e#SJ�8�tË���ܯ�X*�$NdM�a�O�|�m��m����O��G�>���P<�k0n��O��5J�#Ҫ��	��w�fC�G9��X4<r��)�<l��[��A�5�c���|� 5��h���84Z-<>V�g�{��F%���ԣ�����ȓZ��)[i�Є��b̀7����(
���:F����C��l���g�8�H�7���:<�L��ڥ~Od|���V��
�K�Uh�[�	�;�2��];,u���j��[Y��򼮰MC8��숁���~�yH~�P���4���� ;�_3+ZQ��?�U�|��Cg����h�2c1Ģ�:�'T��%fl�cd�o#Rj�{�̆�9�Fv��vax�LX�pm\�.�xB�My,p�����(Џ����ss/�ԲQ	�p�ԭ�����9e�![X\6փvB�)��v�W�c�z�`�L ���8���z��Xt�y;8���
��%�q�����y@/Q���*�w��X%�aÓ2��]�{/�7\\gVƏ�Dύz��<T�����z�'�ܝ���ZSZ���A��l�::ōL��i�y��W=)��O�)�H�� �ؔ`mj�g���I:E�_ ]��Ȝ���^���^�OJ��"���Y���Vu^t�u	���(|����ʁ�#��9��Dz0��ʾ!�]��Tʇ�R�nX��*�K���P�mG����Irr9�)X��)�>��Â��3V�.N)�`~=cG���=c��)�AP�ȵ{�ɟ\�BM.���(r��O��_�����W��N{�ٮ��k�p�(�A^/�ɉ��,RmGq�ݖ�Y��Q6�x��_��^,E͖m�����X�ڇA/c���$��z�d{��(���ɓ(�<�>�A�0;4���T2L�C��� �!Q]�뙫���TH�)2u��:#Me�H0)�Jw�3+�� ݨ�Gҗ����Md�a6�����t��0�]�sC~����.`�V�2\����<��h��>�{�s�ė�c���0��L�&�
�l&1ZeZ��|��c7�ip�Z�}K]`��/�͊��bt���W�&�Ϙ`d��ќ�i#Lh�Q��`�_AaiD,K���4�#������`;�u�i'*a��N�j����0�G�/:��^��yOK"����aذ�+��ZAe��7����he?}�gO�b�ӺTg�鈟�X�Ց����J���(�._����"�[�/���s��L��� ��K�!\��8�AH�j7��l��],/Gm�؈��I�v�)�w��1�� ���a̮�q�o yR�=���[��`�V=��Ĉ�L�H��9 v�w����5���Fw�ܡ��+C���ڦ���bomr*�J��R;��qD��DC�C��&@
0(Kc���L"ܴ���3�̡)y����i	 ���%��>��>�(�/�p=æ��#{��+��k��5_�¦#��h^�ۂ����e��z_v��m���ٵ���;����dLה�6j56�ޞm���S>�g㜯cj���$�,	=C�k�y�:�u��:�ovM��9�WI��x�me��a_�+�܉����öe�Y�&�R1�������7X%�����e�$'�f�/.�0
^�?�E]��X܂q����ݘa,7"�+^~��WوL&�eyb:J��j����ǅǣ�>��4��
����ï¿+�������z�}���7��+"-پ��Ս������(o�So��wD�x������g��"�#C̓��s)�����ƛ0�^�7b!w0Zd6���;��A��\��u�'�|bՔXCK�ז��
cF׽�	ؔ�9f(�^>0�}�\��tȴM���l�5��/���J+�@��,�=�C�,#O�0G���`ױ�����=�mkO~� 5�㌮\�a&�(E�� �c3�Z��3�N�}vDaqw����ZR�E�@����m�w��N����laBʭ��GcΖ���&���Mc"ܛ>v�Nm�Ծo/����LM┄�N������}!�Ho�zKٕβ��d�ރ�<�nlC#�A��EqPZ�:�y�ʖ+����.v҂��/��1�S�l�uQEf�1�N��+�����t���������U�Ϩ�)t-�iө���͜8�@���p��x��ݵ� 	W��S�-�``����X?</�ҫ�X�*3>�xC�ґQEqo�a�:e� �߂������t�ΐlI��{q?���m����4ä�������ZK%O���~�YC�8U@W�����_r�"������OK)�Ŵ�])��3RZ��y�K��T�"�|=^�9��%G����Ehio�7c4愑R��Oq��j.�{��6�YQ�!%�k��]�H�H�W���>t��&��T��a(�*�E��U�:�S_Y��׌�,���ي�9$� C��������<�}�MT,_DzM���6�\CL��Q-��Ɔ"P�j��`��M�Ox_�l���0:�u���g�6"��1~O��qߍ����td�?L��$��#ST���'Yo����Y��Zq��"i\�TJ"q���{X�Qh���01�B��R�N����§M���kP4%?����l�<�u����~_���W��Dȋ�%� �|�[[��Z5r��n��7��/N�6������MC�<d{�O3��Sυ`g�-�F��2�֔%�iQ�*e�����AZw�`>A�y7g+�
�r��]Q�	��U�
�`b�Q�H,kLv��:��j��oɯD�r�:�az��^E5��e)I��K1��-�נ^lN�S�zψ[����"oa�9��(�����<�E!w	��m�8y^��#��C��UL��I�4ɞ�����6b{�ha�d�f�[�H=�h�@CH��B��JoR�L�B�^eR���c�9�},�&O����� ��3�pAh��m@�k�wm§����Z^�y>�ReY.��<MH>�t휏P[�]��%�;V�i��������΃C�<,d��y�J���ND�7�����,�F�* ��Me��󻼨�R�^��Y�|�oI��f0����3b1�Cy���PM��d~��_D��tAG��QV�n��D'���ڕ��W�bl�i�V�)�0oU��J�x�ID��M��o�1�������	H��0�8+���n�w�
4�k'��e��з\-� w~���)v�O'����_�;O��/F� ��SfB��Ǿe��� h����*��r���U;�EFkP�;��*�T�c4z�ݵ�B��R�t�9���l��R/�<�Yy��@s�J��
���h���� �L��Zx�Dtr���nL��/B�mh�����fHm�����U�K2y|Q'��<�@)�s���6���	��c��EĞ��Kf�ν=�-o�#R���έ���HFJ��wR2�8�+�:h\�h����<����W���e߁��Ag�s�C�6��؜�KEW��6���]��]�'eӥ4U0����&^I��P���r'e���7��e�/�����l�Աp�X�f����ݖ�(U����<��>�I:�8�m�zΘ�AXqj���؇s�d������-M�B'�{�����U�v�ܳ���P�����U�Դ96K�!;�:<��bFA��|����G����P�A���ĐsH[�e� LCQ'�
R�=o�/��j仳<mNu��x����(����é�4�6`\�9���r�5���):�9)�{�?*�L�Y7Ύab�L�]���an�_�$�:��^�xF+R��w̝��id�����2���߶�H�3=��񚘜w�����7�5�{�\<̟�%낇K���ғ2��M[R���dX�DmX��QH��BEqj���%�0W#D5������0�O�L�����C�� p=D�y�C�qf��d�r���b�L]����C���`�O~'�m�kŸ>��9E4�_iH�F�eǁT�V��<�7N�C���MZv�߸f���T�9L�����NZ��Bn<\bu�ށ(o�߳T|-�|�_yx��O��٢~c0��$�)h��p����ƒ��=Ҥ4,gE���p��2��(�v�&�J�LN�Va3xB���94֪Ӛ�Ax��x��@x�e[M �n�!T�0GH��]�������Fِu��6�hX̷ܓ� X�������o�bQE��=�x}g�/3q����H���ȴ!�%��D�J|JV"z��<�7 2ٚ�u.;�[�6�hT��v]3�k�����f��&HN�Ņ�:J��������Y�}Hs o ��k4�H��oV<R]JLx0W6�s���VW���6��I��͢M�զC
�8i�U��OI��ܾ�8�G�o2�q��7�)4�v�#sw,�!6���֠0G�(�5���?�g�Y��ѹ[Є+Ql4t����"࣑x>��EA?$�T������	�^����~�ð̓90'+Ә���f7X�`��<k	�ޟ� �tK�?�����G$�=�)Q�3���x
B4���7��$��J���q9KؚAl�_$yH��T_��a�!���=��%}�a�p$;�,����*`q�=�f�~-�܅g��m*��W��`CJu��}�n�e�iY-I��u�ɉ`�n�㍫+)v#�۸l��&���#ܫs�D��lru
$^��ӭ���w3����[J�r�$6�r�a	ح�6��M��0z�)<e�o� P�)��K�Ԁs����(�篭Ѓf%Y����S�E�;��Gc�_�I�!��v��.z�A��nyy:@�VX�W��J��)s��1�m�����(E��t ��v�p�[+m�/��l��bJp��²!V��qM�N�Ϻ���%��01mA��8�i]�dݓ���Ҕ��Øߨ�bBK�|E&�p�1���f��:��Y��N���`�;����t�|Z�/�U�6U|&`_�����q�|��U���8�:�#	J�J�n�I���O:��}N�svA�1տ��l�[҈���ce�~bЌrh(���`g�ݏ0�����X'�di V��Z�%,PD������ ��^L�۾U�=J(qÑas�eF��L���Q�� �)�C�<E�}�ݫ4LC���~�Y�Jm$�ein���_���o�	+cl8v�K�L�������r�R��>�v �߲�M�q���X���Sg~��@n��Ժ��饟��)x���!�IkZ�<��/s�tqӴ�Ok4f�M�	"�ƚn-X5wi��.�>������"tY�}S�6Yd��&\�v�x��A /�`�fB~�]O�����oK�\��2�N4�@�gH��h��>N�]Z	zH�h�Ҩ�a�r)���I����e��,n��0�П��������?=8H?�|��t���'���C�v�xH�Vb*dZ^U?֤�ټjW�~�Η�zNnX��>O��T�K�!��*!JjQ��|�k�S��o/l�u2��Bɇ�w�LǊ[�}���Js�\s�i��V�b ����q�"�|��?"�2��!^bQ뱜)�ʺ4�3՛L�-�&ZfCb߁��ե$���e����5a�P ������C�u�$�;?�;}��.��P�8���?�.5���~H�;ɲ21��)��F4��ߔ�ܔgQ����1�.��7��Є�����~�Ou�:�{�o@I��ߚ��:�I�7�s_��w?Q�|f�D�=�xv�<���7P�YQױ�5��lOT�HO��2��2��R9eͰ*�I�L-2��n���K�����hJ�6_�u� �zqyw*@��T������C���G�A�9G����v��4!1�Mh
\w�~����B!�::��Sk�<��{J���hm4X�{�@� N+t�`'@���Ěkl����ګ4�:-�ז��]�Iʍ\��7���W��k1���4����,1�hp�T6��r���|�oi�Nӷ�k.�;��x�Y35�p3���!����jT]͐�r1�y��j�����:M7��Le�$���q���O�`X+3�\���G3h#bo���CB������3\�Rا$ �{5gd����k(�T�`�ų�S5^���������4�h�%2Q$��{w)�1��#� ��8g�h���*��L�?FkI�]�M�d���ۡo_��#)2x���B�/��╈�4m���l�	���<{���W��q�'Y�&�n͚o�`X�i+�+�`0���>{L;��hҘ5L�X!���O�
�f� (� �DX
���SmN����[�f���SG����:�N�;�2,�n4T\;B�(��p��V�M�,���F�mm�{纏`S�p\_��ʢ��"D�ͯ�d���^�
���R�v��R�St�Y �U��X?��;C���3#
F��r��ӥ�ܿ�@}u\���\=P�o9���d�"�45�Zn�veD�[������Y:z�՟���ko۔��_L��Ґ[r�2jr4v�����*�j����Y)N�B�u�#�F{5�xEʮ��%�t������Ν*�����Ksλ9�iV���-��A�к ��.\�� {�sB����1�<uC����'�>mt��5j�Z	�o��m�*?3��h5�PƲ�pO��>&�m3�|� �JN�NY5�e�M	��&6�F����(�0H���t"��ۨ��>C�r��[&㉀y� ��¬QS�ٹN۹��͹�9��$��c�����V�W���0^�F5 �q�R��L��_Z�)��2��&	j�����b�Tt�S:%JM�Yf�F���Rʚ}�T*HkI����;R��[ �s���h�|�*�	q��X?�ו�^W��UsCZp��(����L`P�-���aB�KHٌR4��{ce�LM�i2��Uq�����y�E2�E�9� ��%��̖B�����w[�gY�DU�D�U/.�+E�ϥx��R~�_�+^��H �7�|����-6X�"��Z�;&,��)$�[/������?�1��6��O�q(�IXe�Vr���ň���)�J�9�/D����%l�.M&R�f����{䬞��c�N�u�%�*������SĔ�}}K?�%+��5�gy�-���X�Cg�m	�c��p��f,���P��Rf�w�����ƚ��7d�9#r0Yn�)�#9嚳l�G�����-�!�%mU�ev�@!y���;-�]���xm�Y����F��d|0.���w֕jp�3�����S,b��uKW{��N4棉��T8<��=H��Y��_��=�v��������|o\��"ˌ�<�`u��5�Qd��&�Me_S�o�!��%��s/��mA������!5jf����zS��N�o�d䎊J�^��?��OTu����x��roavW!�p6��}�]�؟Ǯw���>�����e�ތ�:A�E�{��X�hb��Sp�� 0�4(�I5�8fK���[t�8�pE��Z�ۯ����q�ޤO1��Q�@\�1SڳQ��^�T#bp��)�h���7�
i|�Q��U>����Q	�c�	��ė�a�]����An���׵��K��Þ��m
֩���?J�����R��:i��f��tx��g�$J�9��S���i����3��B:��G[��V�xe&4&R6.p�&ě�4�Mjl����]���Ak�A�T*W��M���qة��&��#��%�-?�6��ѐ�R+�_J^|:�`7���s>A�=O�/
�5؈M��\ 㹳�K�tAx
_{_/��4W��JC�Ȫ�Ԝ}f;��Vf77�e&�� ��. ���7ʾK�in�E�2r����na��9�)������o����B��&$H�KU'�Z)6e	X���{6+�#5�aY�a
,��ΙW ������#���fzES�vTӍ�:���a
�?!��5J��w�w�ՙB@��z�����zZ��A���z3�]����L:!{�P�܂g�:
��S\	(�k�� ���;�%|Iy�$�gz�%�G-�N�G]�[�5%	�������t�U�����He��ښmY���Gf �a��jo�~O^��~=­i�母���
���1��o0}>2�&��)�aT��������s�M�9�YO�o8���Sc�9KP3S���W�Xϙↅ����]S�|R�{���Ƭ�[þ'�"!$&�}��O� �������n����_��ܮ�a��l7)?㉟�ˇ��$��ː��Ե��M�~�xJO�3�{C����|��=�4S&v���`~��qTU�O�/����ˆsHW�O򺽆��il�/��8M'JR;)�x��K��F�g7��eh� �m[�4���Rw�������J�1%i
�㌠��x�Fﰘ�N�7���(�&��1}4d���t	'�Ǚ��ڐJ�))�N�����=H�+��5��>�\�o�?G���C&i#D}���P]����[h�NT� ��׍)��q�\��=!�ߵ��4 �	�$���(�v�r�P4�?tv��]���~e��)!(j�cL<>#���{����Wo���p�+9����{�#�Kζ�f�Q�^����t��e-����M�ϲ��Ǹ�7��G՟sV4jH!c��e�_�keLR?n*	�~��e�w��< )}V�����,�ڈAX��U�t��,�V�M���X��V��� ,` $0�N}ɏ�)	�U�b����������:UW ;�h.�n�eS��R=��@K��ƃ�����O��<�[��dw��&�=��
�6s+�θ�������,=�ȷ�+���]3�F��fz�<b�/sq��ʾ��þ���ޯ_��F�g�/�̰�m���y�Yv�s���6�xy���þ��������;U��j�e��(�:�
ɒ�$����Z�w0���t]u2P ���-����Zμ�Y������l��c˿ll/��E#C�:uW'L�cF��.�G? �^_��@x�nͯl��aAB�i�������a�1k9�r7bQ����Pj,�<O�:���=���C)oI[jA�1�B��[�"�^�2��c8[���T�Y?�i����:F�5�x�D���՝�+�u�ep.G!�C3���,$]6I��U�4h�3!��0��������j.DO�y>Jr.�G�G6��-��.9U�?M����?����'�.��ErF_��	t.�w��cCDeu��M��a�?Q��=�3N{�-_*�ڐ�_��TN�T�jgyؤд�8p[�a�7&qyJ��agL����7�)	�i\�I��"����ûMJ�P�#/�vO����"{�Wrc�RQ�5�c�{rS��[�gT�����;������@y�F���8w�e��iw��Dc�myUg}��	P��J�ן�\c���r0�`����릠Whc;ol��C1��|7=2�����E
�	�a���D9ۛg⎁��]��#U|t�d�PJ�z����x�.���G���p?�j����վ(��92-�zm���6����DQ���)�ѝǙ��>�w��+Z�d|H`8�D����;�J$�_��]��H�d��f=�"����?�ɷ1�� �B*ct�OZ��������1��h�>�	��:��cO&���x�n�($�Q#�
�jؾZ�(�W�%;ߤ部#���X��"�QR���x����������Fq�	&��H0OUzr�9Iѱ�z�,�9��0,�.���fO޹2��h�;�l�#�J�n^�?u?�	��m�[�hД��Mm�WE>�k�\2��q��3f���M�u	b�w]ҷ�;#eU��*\Г9I��C�A�ގ�-�ą��@���GT�Av������$M��Ӷ��YC�q(����w{�v��n=A��d�9��^�a��VW�m�q��Md���َh��Ve��(��:-x��>B�S��J��i9�6��I��k�eE@�f�����n�p;�� �t�H�tq{h�I�ᢱ�x� �E�	Ջn�U�s'��_����o-����ʻ盬7��?J�l����ǐ�wT��]	��L�|1N����b��t�J��rGs�<0�$�䫃�}J=yKP�= ʹ�~V�M�IU���x�t&I͓��[����垯L�l6�3^q(�w�������O�p&]�#
��+�����¶�8�n�O�rlz�0"�}���	\��u�ݛ�uV��4��ѣЍ^�?��<�mON�U�tS>z�%�Ն������J�k��q�'=G����m�Q7�n���Ntw}�4��O%̓�� `�3b�@�]��#�d-
p/�{�sjv ���H��<,����d�BB�/�`};1Wz�^�ڗ+�p�{�ϧE�o��lC�K�-���杨�H���.4�X�C�L�+�n��k�r�%1y�����|4>F��p�� ���B4��hJ9�*鍨��9�U�(�������+��j6���x�jn�L�{� {�ey��ts$P��ب�y�s�����"���yU8�+�E��ޫ�[��?���!����o�WZg�`b�_"ݨ�C�D�Ai�"V�rLr�>2�g}C-����S� ��ü|�L�0dw��6{�h�J��7�6��ρI�?�T�mg,�=�z���G-hq�z��E!��5 H���f?'>�U�6��+��ntŏ���^��8�.6����V�A��xt��)q�Ǹ������1��c�U#�|���]��ׄ�@W�vok���+z�q��B�4/��uaU�� ��<D��0W1i��^�؜'�ҕ i��T ��-�^z�����N�+��Ƨ%Q��|֋;�\��h��	�ǡϹ*��`����+
�BG�j���
�` ��z��\��J��q}�40B�C2���a�9���b��@�lN�A΀�wf_���L�ZU[��B@�قہ(��U�k��L����%�x��;а��c�y�88r
fU�o��]�5.q��a�_F��Q�z�+�ğ���~�)�Ł�b�8�t@3(�������SB%��������ҀGt�&��^���lL��)�w��,��N��A��/�u�6�?����4U��3G`&�gOϩ�>"���"������r�8�'���I�3�aB�����A���g�7.�����(��J� �*��a��&uB����`�5����m�U�<]�=���@|�&eS,��Ǖ�������A�`Ky����J��f�/X�}>؁��ViD��}�
gAp,
F��Q+��Y�y#����L��L�����\�p\ģ�C���W3�tt�F{t��9(��ZVgE�v����U���]��B�H<��uuN"�_��<����W����m����#����ʒ+ͶI"fz�`��5�C��k�2�p��)'F���!̂k.M��3��4�ْ��1ߌ�e۰��Ә�w�����2��+�GD�m�k�
��^J��kB�_e򼽐����ҜKN���4���J9�TkG����Ot�V3��i�����=F0_�>�Rl�[�����Z�ΨXD�{��m(�#�Q/��K׏M�sx^�V�Gm�f5�0ZV]-v	��^%A������J�O�i)��}(D/�HO#`Ͼd&cH_�ē5P�A��jh����"�;�sP��%Ǚ��5b�֦�Oe��V�>�,z�&�ps�d�6Ǌ��s�,�j_��T5˩��0ߜ�H��5�rв�K��[g6��jW��E��c(/��~��zߋ+���;��6�6�hɚB���@j��A#��]y̰��q��g_c[��Ƭ�.�ܿ3�P@`*R�jy&ONt̠Tܓ2�f��΀k�Ro�y�X R�r���7���t_D̈'`[TB�E�����?rS@!��E�7)�_,E�x��\���9)h�8vE�B�)��!Yd+�[l��[KX�������9f�����P�����j�3WN�%�*@U;q�p��J���QF�/�C�
���W��bq#&
Frp���):�iEގ�/Qm��n��s
Tݞ�^���q�Vp!6��
�f�<�e5_�.+��ܭ\�|���*w�9i�m����UT��`�zg�� ɇ'5����ER2.e�����O� B+��XCy5�y�.�F���Yhju�~V��(U�@g�8��H�8�g%�p9`��">f4xV�y���6�G��H�ݏ�����\Dƍf���3��_��u<�Jί�[����I��[k���Y�(G�25co��N�pF�
1�r�s�P�v�*ɱ\ے�NG睏���s����z�9jk�o�%�� ��=��yO��̗���<J��'��>���{c�y�F M6��x{\��[+`zB�5�3賻
[H��,��Qa�0yr[�:�$06Y��!�Dv��3���H��N�����#$���§�c�9z�)2�YN��wA�,�0Ű06�������.L"���
���˔�N<Z+Uۛ����LR|x���.Y<�����������d60;
�R��m��͈]Ѩ�����+�ږ^L���'��W�J�|�BIQN4�B����l����#���m<�4�F�����b��<�	F~p.[c�C�<PB�/�+;�A�=3B27�js̓�OxH�,�Y�o�>\�p���gܫ�pyp��M��ꭣnY�kf[rJ�O��F�,nD�� nM��Q�Xg��ݓ��6��w&$�E^T7菆5����
�w���}�(s�+b_f���9� ^�n+kΘ�_^��B� �B����"��|�S��1����uX7�B?W	�M)�J5���;�D������+S�6��z�6]ۄ�أ��5�]�c�D�K�IT�·��
���>J�r
wæJ��[���C�m}3a��(6��2zo�g+��*T/�)M)pc4|w�Ջ�"��Ą#���0��%*�7dX~�y�lR�V��a� |
M�����۩x��V��^O��+Zv&�ۺ���O:�9�l��&�}�	�+/��9���Q%�<AV��k_9<���9}�&������R���F6ѰR������M7���&{P��/�T�|I��V�I
<S�"�hr�R?I�c3��J�N\n���WKwf������]3<U%�Q.�3]A����e�*9��0�(�B�z\`�`^	��|\ xL����8nYfL��9k!���D�d�4�e#�(��^Cwθ�G06�N�0pO䣏��}���K�䞲��%�Iw���$�S�5D��S�%�5WA]�:��L�(9��<k%F�/&7�Koo_���AoY�������
geLc�C~�y��k1}��Q��p��e}"��B�W0[��= ���k�@����c3�A{�e̒~��8�L�U�3(�Q�b	���S'�U�i���?l(���trq���D��P�*'Y��;�qs�c�9Qy����{-����t�+����X:q�J��&�X�qL���̱Re���4~Kɣ"󜅇������Y��؋
��%��qy<F��S�Tؘ��E�����O�5B�酟���+Č�����s
u�xI��]S�� �J�
\�D���I��r��]�dR�va��|3�$���8�n3W����Wf��-�> �
YE]��a�����*���\��ssUMHJ&�
����[���[�'v��sC�����7ї��@�d�D��z-��z�}`��/��{��j륋Nn�\�I\.>/�,W�mpZ�9��/��`!�1����,�����2��HVƏaR�.�4�:�`&� �S>�OD���ޯ�|n�[x��g�6V8}jh�U���ڝ��qi�0�#98-K�,c�3���U���ȠU_H1����9��H~���jP�y���K`�Q<b�&9���2�t
��	vZ��dt�Vmq�׃�W⚎$}�z?�@��FWv\�u9&YWBf�%�.���M�'.7���}P=dPb	oLUh1+�e/"V�aiw��]&{���>���.%��^4^@]��zֈRϹ��*�d�{oF~�H���h֫l�'��JG,݃�&y�ʙ+���q���������x0e�p���)H��%�,h�A���#�_/��QE�w�qOF����C���G�?w�w9t�~�*�ϡ|a�h���7� g���Nѥ�a����'\7:b�CӞ[Z�3�7H3����:}x"p�"F]ʈ���D4��������[���j=}%d����sܡ ���Ј��t��x�}����)(��3J4�Y83x���Y�"@詘SV�?xTJ��r�!.������c�?��a,['[?JWR���LὶH�V���ca�&X�
1`r7B=��l݉��%m�un<f��	+�������/�C{q�,�XIFj�g�~�A��v�����&zĚ��aS��S�=��0>��{J��}&��-X�;R�̛B�#����6�uScZ�����w�+�l�$��dr���ca�A��U���QaX������M����Jإ��Z���q{G�aS8�H�3r�-����ٚVk��XU��[Ӟ&;�f.�7�5�@���乴׮�Cn ��B�@
�߿|蝣�zv�D�41�C��̉���th�X�G3��S~�z����"
u�1S��3����ڏc�&��O\y$w�����<����/�*`���9�̋�2-�S�v�v�h�Uܚ#��`c��hǠ�������dz���|\Y�{�������m�X�G&^�T������=�t�s��w�1+Y�6��8����dz�;�mO����v���C�L蚪�pУ����4�~S�vO�4t�b�N�j�ݩ�b?�h���b�W�|�m{�Ňh�+dGf�ҥ(��lfK6����!\u����,�K��3Mj���ۣ/&C�>|<�W�	��#0�M�kYh�b��'���m��lr�b��Q��Y��u�t�d胳�d؊r�M� ��e����_!�Ѐ�\[Q,���!n'jd�Hb^<��5u��G�L-����!u�I?�6:��������&+�*w��!�x�O�P������i1E��W��8!*Z�T>�BD6�0M�4���]7����3&t�.����z��{,�P��0"��ֿ=�����d$�z��U��R�X�d��uoP�4z�{�*-1�*�˼����I���d�b
�N��K^��L�S��?ڙ�a;���1D���[����5���X�M[�4���������B=��f���a�P')�V�9Z�:�gƎ������jˬM��A���ed�_���ɘӡ� �H�)n݀_�(M�V�Ʌ0�к#�I�?����N��yWvږ��{�B>��ԃظ��tu�[h��1�N�hlP�d�訉rc��m���{� ��:ܛS*%���hEZ�a>Pʋ�BtruqCk���k�ظR �&2�aR�JRQ}0X�Ma���8I*5���5�z�z�7r*+�y+A�f8L>�c�E�Tp�������>��Z	�]������G�r�x ���mC���^��2��dC���E,٦�����\��Ģu�(�b��D�Xl��<���>��u'5��VY�yV�6�;�}�?��r՛w���� +�����3�W����l�Q+���65�[0����FS?l�*��+�ie����0eW�w棐vP*���H��O"ʃ�/= ��$�f���-{bu�]r����ͼ�8��`�i1MNJ�ŵ��d����]Ν�{_��`�>�-��\�&���I��i)EaOh|�� <x�ɏ�o��24cP�|f�S��0G�x��$
g%V��ŝ	�c�np��B���w�wv�
����_���:���0[��K>�$E��G����~H�k���E���@:���ZȎO�zYz+qc1k����

�RJ���Gw���*^�$n�Q�F.��֥�M��v
0�����$�Z��Ȇ���K�"���c[b�|W��Du�{�q������#g�x���Q΅v$�A�Vv�[w�+
��4x���
d��;�	�"��2Q�I'���zc[�t���O�J��W���=$N�4��S���_h�J�����[_�3ƕ�'
1�>�ߙľP�'��m��$f �)��m����V��%��,8�4v��ג��B� gR�[@��N��2��䥟�3/�3��L���XA�c`V�x;�5��;pl��n&����m�W1�b�f��l?��>���3'"��!)����ޗ�Z}=�P�B�P�sd�r�D��B�Y�-fy��#��%�sC�%�l�/�>�>%Gf�� ~s(ljG�Y��&�4�4��U�2a\��G�H�G����X�r���>�`"��t�C���n���
��o~!��|��n��
���:=�}�˺y�N�JL�j��C:��b9�{]��l��$t���AL�|�r�q쇆�����JM�V�w��V`d�Oۗ��m���\*CS��vM����a��S,�z�ᝓ���P"����<?w�� �{�"�Ԥ��d\�:\���M����\zB:-��2,�ը8���X9Q�/�#ߩjc��b	���,��F	��T.����d�*�8<�[����w�������#��{��O�N9��/���V�H.�w-���r�hMVԉ��N�>�y�&h�ס�$��c7�v ;]\{e?YB��)@~�E�|��|c+e��T"��J���>�)���CM�]���r�#'/�ۈށ����,��!�����yr�T��%p�6�P}��_K־ �Px�G���su?6`[�ի�n:�z�&㙃pb��X E��¦����#*(IFm����$t�#�T
o�͎H�u�����'�}%+e�_�|���SJEE�ɘQ������%2����3�E����SU�<14�\YL��pQ�O�P�\�}.d�lY�BY�:HFk�:6j����͖G��9��E�гK�IE�N�����X	�d��ܵ=\��riU�C�P���u����w20�-��h�Z�sl��`�-"&���m�=�ժ��d� *��������=��x��"̽�5�S3�Bmh�j��qcx$^o�)89���~QMH�`� Ē���z3ea���� :>̳i!�U� ��W��(��(�X��ܳ��q��sa�����0+U���:��,�����2^��U�p	1�[M�od�iZoË�&/X~��	Ar���{~�N;d+��Nƪ $(0����U�m%���x]3KZu���W���,*�����$��\�g�
H{gR{�9�>���wNE=��I�Wp3H�#y;��rqlU��U!���!q!�~u	�$6~?�UtVԬ0?��Hا���.+Nmv<�?��A����0���X�w N���6<�@ZRE(lJ�a3C��/�mR.�>�B�޴G�ȒS�NN�u�ď%�N�S��@�2�rǞ-O�l}�Mq��c�ţk�t�RHBϏ5�H��B�؍�6����p���{�v�|����i?����~NJ�h"=up_�{%��G�8��p�4"�ŎQ��2�ڑr��tEb0���|z(%.n�T��ux��'N��(؄V���<P,�y^��5�#��FB�];��Lr�;Z@G΂8~���4����Zbk�p\^k6���hsI!�<��+�}�@��)a�$�O�iu �D�$�Ĩ�?���~�T���n��� JY��X"�7V?#�E���T3��l�J@���� 8��&��A��+����?��3������Uacr<��8O���tC.z�u[
�Q�9�u��.�3�lC�^����/6e�L��k��N%QY2f�C��Pޔ�r�θ��i��,(��,U릆-x���tr8�ᶢL����e9H��Y<ԁ%��m�G�V��!'�����U��k?4�!�K����d���Ў��T_ބr��'�Ԟ���<�t�����4��Z�Ֆ4]���5��$�B�̙���Z��S���)�a`CVd�z�(����7��� ��a�
�?�.����˅��HP�͆yԜU���.'FI����G7���d������!��Á���G}V�m疋��kH�ݓ���W�f�]<�4,��+���C�Yσ?�X��=�ZZ���m�J7��d�D��qD��"��pWU�k�h1�-w�UV��O��<���Q���L.�}:�fq���ı�0l}3ݗ^����ˎԥ�z�gϔ7�����n��}BD�;��ϷT0�N��|��ܓ=�������;3�����Y�����,O4ys��;�wk����l�G�h�9�+Ꜷ�9b9a�P���D첚��K����a��s^��s�� ����p:�@N�.�@yFe����w���<ߟ�xJ���%�kET�g�0�!����gs����g<��d��U���cn�%��g\Tk,튢�3c50���}�V!�Y�d;v7�Eʡ�p����9�I6�W�
��j,�Mcp��ܒ��|���N��uE�J��][�g���_v��FP���}��՘O�k���7���z6�r�%Ƙ��[��0X�!�ut��c),�-SL�j{V�~�a������X+ܫ�I�bd��!o������%�W�����O^�Q-�&`ZU���Ss�#�R��y�����ף�l��a),(��p����
� ꗴ_����5��y���j��Vj:4��[��`��۸J��Tew��0�-����'r�!�N��ϖٺ�F��8�˂{+_,�}�L4Y�1пdw��a�_��}�M��pKQ���p�Uq�s�v$B4�z�l@�Y���8����`7�|���].��3$i��Z5	>y��v3�U������i���T�m�������@ �Кv� wFl�� �H�i�r���lm��������dr}T�u�!�*ދ��.Oh�Vz1�3�37q�,�!Ƨ�.�A�2@�\l�N�$�5�&E;D��\Ȋ�Y�r8�k��2t{;�%� ا>
�@�w���_��ƛ�h'�P
�Z�o'�� �e��t�[���k�
v�a\6{ޫ�jQ�R�zu�[J�5��A3���κ�pn��|�4?oݜFa��vրx� `����H~��_��{�XDA�:]Fe���3[y��WA��&�ډ��
<ǆ��P{� �tM��Sx]����Jq�AZ���2��4�
յK˱�� ;�M&[E���j��T���DUn�l�Bj�Ԫc�{@·���;A��-i�N)+o+�x6�*�����$��ss�eVM�z-�3���D�|��"�l��y)��ƲlF��>3LS��_����Ҿ�E��cq�10�өБ�J�BK�i�GrtJy+$v(�١��J�1�/K��N����ѫ��hG�oʕ'�4�"��`����*�C�*@&PF=A$�J5����q��o	���*�g�[=؋V�~��6V3��=_��,i0�2��r��A�?t��@b�=���UN�9�D��qЁ��b�mK-y�N%?��@�����(��ฌj[�e��j�%nV���*�Gi��� ��Ƌ�"Og�>5�}r1� �f<�����^q�k�0��� pn�us�̵㴣�����:ᒋ�q�4j������r��t,s)��"J�,M�)��W�BG�+�g�Ӣ�f;��F��G/��$��ɀ�[
?�W_��T>xrr�M�i��%;�����+�Zp<��*�,�Z*
�@�)w�0��j`��Kz㟂2.�8�I�yZ�G{�lZ�����2��8<���M�M䈧2����5TAWaz@5�[��W�p1��ڻk��êld�/R�ʂ*�.@�9~ۅJ_��-�6���x�hj�CKx.7�0�����C�U�z�zh	�F�q�y\�-ЬM=`���u��I_�����U����D
�&+H����~���:���f����(�̎�?qm�3��]y\J�0��Ȋ�t���8�J�si! ����ޜΒ��n;��;��0�o��V����ƃ�I����p"W ��2�+(�P�T��϶��kO����|��39٘O��
��c��ZOZ֖"�i?I��9�R@��2��~����o�f�������Ѩ�j�kU��X���Tw@v4��x^K�@�n?h���:�M��^n�68ߐ�����_�cW6�Φ��W��Mgku�l�~�/��‼.}N2-L�(�6��&o�⟫����*�����"�����l�
�����Y!�<﯀��O�`�rf.��FP
��c��z&��}��i�}�Yʱ�u��2�=Z�ˮ*Jأ���tz�cW�|N���a>��_��Q����}���^]��6���ϵ�V���F��B����7��k����Uڽ���F&'��$[7��ޚ�������vOy(ܒV�O^a#��G�l�l���.��N�q
l�^��J,�lk����-<��Hy�[@�L�Q�'�4���m<L�S1sʽ��Na�Q�6����nh���D�m��`Ȉξa �����E�R�I��Ψ��ͧ�� ��o?8/�z6��"��ئ�}`��m��N�J;��z�|5�,CB���e�GÜ�MY
V1',�FE<�*i9��-oe�)��cY®^�::8�Y]�A��g�|~7o��>S|���O~`׼�؄	�Þ�5�\��^Lj��]����n��"�=�/�𞪊�^B��\��n�=cܯy=�ԅ}���^+�
|
�Lׅ�}YW[ r��M�>}�W%Y��a�W��rbr�������X��N�6��gvU��(�*�����	Id���=f�rx�'=��0�8�i����=��ԉ$e�~��R��� �+8*ݔ6٧c����4|)j�
e=�g�3���k��'r��� �IP�s�%;HL�n���{h��k3→%P�5�`�ԥ'"���	w��9c�1���4�n�Ū�?W�3<�ob'P�q�r@#?B�J��(�0���NY���$��ɦ9s���I\cP��T�1HL�Y����w����MFW�ƨ��(��MD�_^�81_����9{�7r���t�y�bʾ��Гz�u<�M�čћ�w7U� \w��*�Ƭ� �M�G���f^*�N��f��\HM���evt'9[']}�[�o���SlL�����w��]����*mzdli���9�� �k�3A_nIФN���.5&[�������`���"���5���u���{����6���*:b�}� $�=����g�W{���4�uf�u����W���}1�Ia�-�n=3�܏�Bij����}%9�мa�*�z�-�KM�7�΀
Q��ƛ,�:5��gCzMP��s�8=߯��hZ_��Q���nG��"�'���l���i]�F/�GS�Wa�3c.[(wd�h3�t�L��H9��(���]w�l�vv�Qf�k�cW��[�ڮ�di�K3�������t~d.*&�&~��V��˼?��!�c��7�G�f�L)�\+���z0�hy�u��է���JN1?(��iM�ѯg9�C�Vg��@��Y$��y����KN)▧4v{u��5ށJ���Ҟ�?�ݓ��~�ؗ���>>�/G�|P��0nE���L[ݸ�k�4ӯ!����]&��0$���God(.��D�(}�;�_��n�e�����T����T#U	>Ӱ4�F`p�5X� S�ҡԓǈ5i�I�S��"���Wߗ�}��x|i��˖�\\��꿧� \��@�� ?�i�P�4+	�Ye�g��F9
m�>\���԰Kb�M��,�.���W��B��&����/5`�S�!D���Q�޹6�Ʌ�; ��b*jO�����[��r�H����8j���P�7�D^u\�nō8S��@�w�h'�]�5{�;�{�U�}�[��;!�a0Da����t�O�����Y
X�N/�L��ǚa�����1�1���2<�E� ��	J�����[C�+���Fi�̳
dkT�|ĕ����l��(�����䁤g6Q���	�$'���5w�&y��c���7�I#�Sl2���ˡ@�6��@��#连"��2M<T
Ԭ7u�^�,�`�l�A���=��<�zI���%��p�U�e�ւ���Ӻv���¦e49(v��a�w]!��G���RZ	W����3�����:�@���V��"�e}��LXq/�c�$��͊"�ҝ9��O�l�t*�L`q�GO3�Ĕ�4�_<Ľ9B�B��/�)@I���CG��OP����͓^yp!��.vG�7�&��3���e�Snw,Kj�ܣ���#�y���K�)�$}�v�RQ���ٴR�9@�m��c�a���~�OϮ�\HC�:�5i�����,�R�k�T_��k���G���]0�F���D�jA�3����qq+>pt�2�2�W�a��+Y�zE�7�����B��j��1hހ���$>۰��9䗵/�hAE�P{dp����j�g!���Q�~}���-��Q��S-g�|݀z��lz���B�A@g8Z�X��#����A���H��E${=���emE�#���� ���4)ܵ^z
Q����;��,6���s��%2�/GT���V>c�fqU>l�eEU��M@RD��8o�.�-�/D$�Ṳj@��^Z��i�G��7Ux�ԅ���U�A�X�vڌ~ۨgXJ��i��Z��+x�@@�^���J�Dh� C
�Pa��r��Yg�{�/[�m��%��g��b	J�W�ܠ{g!	
�R)��Z����>�Zl���;�Md�F�����^o�4���=J��\7cK��ֻ�1��>��ā��3/�3T�vij����=N��̨�P�g���<	g��$��X0P.�I����P�u&ROľ�Oǘ���:zݒ0�z"5�9�龓�1����9jq�z��ޚ��>�TI5�[ &"{�+� Rg.�C�#E�?OA�f
���L�켰��"��`ڻӔP'l�^� ��jPqj�Nrg]�4ғ�՟y:�vr�'��NCX_�g}�_��+�w�&�wk`�8��q���;�s���vC-aj�@x����J!O��XgFMgO����P����@T��"���'�zY�Q�rxdr���裠��8�b�A]��M]��qb0�
eM~�=�Kg~�mn���R������o5oھ�;[�T�R	��W���d�Ƀ6���X� :�v=i�nK}:b��yr1��[�]���^��@�ѥ�;.k���{�#�M�"�0�⽺h���^4gP2��^�Y u�)��g�ШF_o�{ޖ��^/&�+]�8����l��:�"0Į;�k�u���L�μǴƃ��a�ֲ!�L�D�6t3�x����w���S���mX���B�܌x�O$�����=�0�ogڲ8̩�ʬ�,�y�j��ϳU�)�
��q_��ш	y��+6��G;o��G��WM�h /&�-v�����?TF͊j�?�������Y�*5646��KڐD��J���*����Áe���[���t .�ŷ(.�&!�E1��-��$�/�!/�u�g9qz�R��|p�Q$��=�=ڹ����tX�\D�S18>9' ��e��� �/���?Ǝ��uy¿T��MX���8�r^�����+���Ӽr��1�hzM�-}��VbR����C<�5p���-�.�զ11)G�2��Î-�d�
�9��qlHU�'0��I졼 j^�#p��i%��F����
��{��P���wLM�;}�?W��L ��鬋�f�;�?��f/����u�с_K[��:T�͛t:8���U���r����'>򔰕t�E��S�&�'6fܒ����&� O��%�u?C��,L�Ov�o����UF�Zٰ�Fi�X��P�<�=P4Z�:�{�d�aT�Lt�W���zb�8�%�1�r�����H]�C꫼�:#8�*�}�D��%L粳���D�\E��-GBBXÐ����xW�Sm��k�nO/'XJC�	���mx� ܧ��1���Bڶa���_m�WWU�
�`@Os�"����.g\u�<����o���H-@�!�v-y�:�ϹL�9"�j�|�bp�WM�~�v6������Xk�:ު�����L1Q���ce6K�nĝSǩ���zE��q��i)�b���Z��!|7�O�K1�;��Ǝ$�>����� �1�U<��C/Q6�R�*M�Y|�!�	��b��7��[�͵�*�D��~h�8�n�)S!e|�����d.j>�OM���H��m�M�I���=��y
˽��.f�O�=~.��Ɂ��.V����8�<�M�F�]\�kJײ����/K��h4�!i�W�*��4�����Xx]��l�K������"(>�!���7�w�q�4Z�dxj�K�5��:zuCY���5��H��T�	xT�Щ�Jwl�j-N���_E��G��s�y���BwB�O*���cG�m���
�Pt��~ΛP0���Jt��=<7T�X0{��՟��k��=VtY8|̕���6�>���s9���/�ߡqH OnCa��l�0��ru��[1�Ӭ7���a��Ϯe��1��Z�7�� R���%�u~���߼Df��%	ڟ��'��w,���| �C<_��M�����bё<�}�nULQ��S�ms��}H�������y ��t'�x,�N�AT��'�݌�#�ӿ��<π����vv�sf"�VSDJ���:�f�'�����`q �>`'<����}e��,]�eJ���Q��� h&�;�N'�c��k��Z_D��[b!�(�Z��D@�o#����2 N;9�k���C�E7�MP��1�ɲa����1б��)�6G�N������Ja�O	�O�츇_�"m]�?�t�E�S�zM��M�s�ѩW'zS��5�s�>���^fX<P�����%AB�Z��!���}����Y�[\px�upv�%��X��;_s�.d�R��7f�ޭV����t� ��a����J7j钑mҧ���2�f�ʡ V�1T,�(n�����wfg(&h�G� qS�0�2w��<"Z�a1��47�@vme�$�IWE� �@6j�F�%�~g��c���Q?ǺT�Yp���ӿd���T�4vVx�zWàL��Q�iK뾤jp�#��O��H���s~� � Bڐ6%A���p��(ϡ�)c��j���* djf��y)��'��@����P@W�~�2����o�.��4@7�Uf[��g@C��j�U�(�D���u	��"�
�7DәR::m?�^
+0���eA�������`9�&x{�2�d����Mɂ���Օ��|�U��ƜMN�q7�E�R��y�����RE��ql���w<�����ݸȲ��m}Q��^�H���-ȍ4��q x!���f�{r���dҁ��kȭ����{$�|:�*(���0�8���W'�������0���=VR��u�NN�'[���9/��{��2_�ҺX��8̔ 悉�'6�l�|��0$���vƏ�VZٺce�#R[5H�|;6�F�OS�I��-k�~r��}
�z���l�o^5��i�3	�ɭG�O_���M��K�˭��n�18���`X��ns�-p�E��{;0��w��Ep'��=��#p�k��������Ҹ��c�H�r�z0���
;WK��o�Q�k��#���B��H� O/�k��w E0���s��ֈ�o::��ϫ�s���:�P���,���r��U�OL-�zw\�b�I��cA�%���׹�]
8�����Hj):ٽ.Y}������M����]3(D��$��B� P��Ҽ�,�C@%B�bKx"91����q�M��̢T������Hc���M(
�a
�.��-D�(5:����5��
jp �w�V�8˥�ݴ&v%q\h��u���	5`�i�M�R�Y]�x��QaTR�Y�2����3��+r[��Y�@:7����\x�8���N:x;Q��Y�%�{��YG^�����K���`�H�P}�}~�<�g��|x��q�w���]HjKK����V�W��+"��"��u����o��i�;ɠ�#�߃�*���%��hU�!zU�St��P߁ zX�_r_�# !eGz�ՠ��#��R�3�%1���_>x!�A����p:�7�	A����FШJp�Bݝ.�d��ƪ�ċ��#����0���<�]�t�敨����^g�C�K��Lr+�o!/#����E�̲a�C���	& �{�gj�נ��ǿ��Y�0�5��5+O���1\�d�#��7�U�&���K����˦�/}�awU�Ҙ=����$źЭ]�oVFCڔO�;,����4�:2�Gm1u���&_�TN+r�@�|U2M�e7��-D����4�d�C�-y�"��')�/���1����>�����'�����mv7�`Sp��ɫ9a��)z��L@{��Zf|�>4� �~*�`��4]*$B�^��lGy�^�y�v��A�{�Y��G&��m:��*`����L���Y]���\��^˪G���*Xcs��1���}�}e]�o+_6��Lsz|(����C��#I�w|�yL���i���Ȯ���WA�YP�4�|�sY���Lo���L\1}|�:�Z޹��r?��=� �Ok����mq?U9�l(�/��8� �����?&֢�NYcβ�HP��o`%�q��V�rp�
q�D���~#�wIu$�4=8��^7���b	w㞢"��f����]oj��$z�e�+�S��N����t��\��.h߽��p�=M2̓�e1���oM�:�t�ێ�x���y"�	{t����&��W�atQ2�Ҙj~�ӊ�	���>�S@�#��xM\��WN��U4P�`ݙ�R˩c��@9�Ʀf)w�s�a��{��e��Pf�X�+G��M�Ͱ1A��RϺ���̈���x�%��$&�6�^�� m���65������tf�}!#hs���HG�8.q�=	���9
[f�D�W;�� �W�([L�YMOnA������OcU}	�Fv(��Ftz�X#��f���u���������h9�њI���&�d����)�W0�+L�B�Ш���~����.��@�);rAeI�t�1�\�����בb���46��v��V��	ɛ��?�k�sx�cM��O�-����b��� q���4�rq�OKX�� ��Ԃ!���	��+7�=7c����CU�>;�ր��[<��f��Xv8��Ws�������n`3<,ݞZr(�= �ǰ��6?c2��{��Sg�e՟I��@���#��o�+
���������F�1aF���$� �2��jP�o��;,�'@<��8��0�E(�x%�d�~mt��ۺJáXNa!]�{ǀf��ٴ|e���@�ž(n�|$J�1���d!M���{��N�7�C�]j�W�>���?�:�1�V9!�����\�ib�H"bd��K�+
D���4�sY�T��4͜�.���C�H^����f��?0 7"\�գ� RD˩(k�y���8Ge��%�g��p~��δ�����	�c؀JԺ�sS�p��|��1���x�e׮�D\�Go��.`��m"��2=��b���8�+���P�hqB��F�{��i9ԑ6Q�6��F�	��Ѭ$�]���Ȧb��ysx�`	�ί�l�s�'J�"�ߢ%�S��m�S�d�V�:���"1G����^A�c%��t���
��c�@�A�dM���9�g�>�LF�'_MF��O��T{�m[�yӝ�M�8��@�GA�+��kw p���4�� E�e���i�̴4�8��X�ǃz*��F�����8C��DA�s��q����+�u)�1���AXMn*6�<h1�[�J�2�e�X�{p^�sL�Z�EaZuО!S7�$1��07��E�ݾGX!����Qn&K�Ϲ��ժ�=�N-�h���1l��"iR(L{4�%G�Y�]!_�m.�q�5`&E�B�ǥ�i7hM�H��f�4_�qB!�|�.�;9�*eS��Q/3}���#��(�=�]`f�h�5���cu/�L��%�@��K(,`opV�q�'}r�kx�I�S㦞z ��5�C��� c7)A����:H�LV,����qp��&|���q�EA$����8)jґ޷ra]t�d^���M+dƨ�)1J����{g)���BH����j�3}�k�_�Xhu�T�m�7��2xv�gL�U�T����*��L���k���qل�E�须Z;���xfI��R'o\��e��P7r�ֹ;��;v�Q�x!lk=�� �s��$R[:P`^��ڎ ���&���P��j�愽@ț}b�S�AS�3^�У��Q414�gtE9��X���oG\����~�>��#�������U4w��>�[�H��ЂiO���z�{����߃l��4%1J#�e���C��H�{��%��˺k/
jȈ�~݃�
�!'�Z���<q2	l�/|G�AV��/>��;1� Q�Z��6}���PC���evÐC�aʟ<�����k����ٴUp3������t������9�A������֊;��� �E|�wF��<55ʖ�"��B<��ߴ��0mK�#��0��.U��1���)u�X}A+h��0�Z����S�Q��W�"��ׂ�<�&�"������kL�К$�]�b�Y���%��WI3@?�b2�j|�	�\��ѪO�ԦqF!';)�3�Ar���giA9'3g���"~vaāX�]�O� �f8U��B�ǯNRI佱�Q���J?۰S�-�V�}��cM�����Ʊ�m��Я�SɎp�����C��#g�tP��y�z�|IO>S��	��4��𘕫%��<�ӆ��#�����bd:�bs��w^��)=�<]ȫ���� �ߦ���Z~7���)[g��1�||�k��<L���7�*���Α��u�Rov`h3N�EljD���s,���������������G��
YǞ�Wa��p��Q���a�`�ʨs׈P7��wc�����j`���ev�g�Y8���gԥ�tM��P�1�x�m�-�z�mh�Z�V��2PUu�1��� ����*#\:�"O�i(,f0��_�R��a�q�xkVQH� �^���9Z����O"-C�o�>e�6��2�^4>��	<sO8�UuS� �/e�s�r�9��H�tD+eY��b���Z#������E�I)�"�mD�4,�n� +9ni��OW����)zK�څ�K�,X��K��dr��x���=�j��l��p�ǵam��Vq�&��}o�x���{�i��U���}��^W�g���{Y���uv��S�����!4����6_��f?i�
H�pW	�]Dw�%}&�ƍP
��i+8Vw�8,
A�j��e@��Y�v7c����v?�ه�X5���v�~�)�O�Km;!��#3�	sġ�ޗM�Բ���kB(]�~@B�KI�t����01�5&��4�@�B&Y��a��?�NCJ�[�#��lE�3���o��"qD�� �:�l@���ݽ��FʪhW-H($�#QS��þ\r�������2�x �*��rĢS}6���%�����5�q�*��ZA�m�~Tz?$�H��I���W�_v�G,p ��LpP��������mR����<�q��;��\�^';Z�99T�������=����Z�����.h�]�YB͟�I�#!(�D��&Lo3�[�٪إ�����~�a�5[����T�ѥ\xr$���k�"ݶ�xz9���3����IWL$*��7��t�͇��5�4��M�}
ڿL?�������6aop�D��k&}��݆���#T��PMXr�^��A��Kc��;S;��,�/��t�
��f!��9G�9�ɶ�X�&�E�Z��R����hM�+�WȒ�[ùag1����d��c���k�p������O~�ω@{I����ڸ&��Q�=�м�u7Xǐ�=E|����bp�dC��������X�.����MV�w���*���6N�6��$ /�-h֦�p��ٶ���t'/�n$gp8s{���� e�T�`�*�`�L��������^�H<x�:,�:��5ى\|H-ԐR��P��m|����ϼ3�*�]��{�I��X�4z:&:F,|���RjR���! ��=˽$�<.��j�24�+N]Bt������ȩ݆9M���ą"񺂪�IB`%4�a��L���L���U�
g�@|z��xzj#�۳�=�y�z�ظ�d�����i-T?��z�u�>PA����9�"�>��1 �>��七=T�$T�`���������DsQdR	�'uU��~�g(*T¹�T�꯾p�F���-�,�E���o�ru
���b���&(rlB���ȖX ��5{��uS�������:R�^�����?"f���2���?��{O�1���2p�:c������������x��)�KG����4d��t�����"��1М���f�j�����p@���l�E��(.�S��Q��[$��&"�$�~y�Ȍ��P������q��O�$n!ԏEO˖�7H�h���rC!0T��#�ȾL)�H�-�p�F?�]k��F��J�"u����pNb^��a]�Q�����(D��.�r5�t��_'�5a�H�H8J�;>�(n��	۲,o�!�� �hӐ�b�,��:�y3���4��(��|�`wr^��r��M���t��C��1Hy
�'�- �3T4�� %�cu���L��`�WS�1������^D�����O��w���b�{�&A�CS�K�������-s��_�bS�d�ly	����(
����]�
���Ԑs�q]���1���.��3 ������f"�F����:�=��$1����HL|6l:92�����%�"V����.�>�`������>�c�g��*�"V�Σ���w�{� (Hw��A"����ͱ����1�$W4{_����O�S M7��u�g�f�|e�HEi�n6_��.f��}��#�qD�F���̖�)G��Sbt���G�Q��ǻ�l˴sU��W't�u�#vE�o��&Z�d^��&P�Kd�?�뢳+l��4���,h�G�Qed�f�p�/�6չ��F�*;�#+� ��,�*�B8�Źβr���$wJi���x�j�K:"0��ׂt���S������\T�b���+j+d�,O�1I90�`�z�u��4�BZ@<bn�(!b��f�ϵ+�i6��b_:09Ѝ� �ޙ�`���X�`�YӨZe����.���j�n/=��|!���p��px��Q�5���[a�S$z���{ ��k����E�$>�,2f��������.��ֈ8�����ߺ@�E~��'�ϳ.)H�$��n� }����!����J���UP�����Zm�<7�s�J.�s��R���LZ�TM5o[�����-����R�gz�U�h�"G>s�Ay����+�1��b����ѯ��"���p�\��C
f���_�3�a�s9�6nՍ�Wˁ���	\J�y��w����pR�����;a�j.��X ﴀL����Bf��[{L.���<9⏍V'�_�]
��z#�G�� }�C�Vn
����޾�ZEL��~�QM/
���p|��v5TD�4�5lV>)mɚf��|7Uߪ\�T��F��� ��������A�;���;N�c��6�x՛�!�{*���o>aq,��c#/�p'�#�y�K�7e�ġ�W�m�  ��[)�1�Ι76@#��<R��
cw��#�#Q"ݣ�Zr�����lq� ��+:�� ��2�gWD]��� 74�(�YZ��ƾ�dh�Ǝ싄�pw����X�	����w���p��Y&>�=K� ���P[��P�<įK[Z�dO1�s�=}(?e��F���/��9�qy[�!���&1v�2�|��-����,FC������Yh�h�F��_K��6� �"��"!"(ƒ�� ����a���[�zأy?vy5o�������̠,mBۅ�I/��dJڣ�}X���K҅�rYP-�8;��U�V�<����?�[`rzvţv���`)�m1��R9v�J2& Ǣ{@ qm�"o��~nY��6:h�HӒ9��q ��!��e�,�˱B�[PhAݴ���L�2&r��*��"��z��!T ](|�x.Z��,�"�x�d�����픨`��_����B�_�A)H�sӌ���,�3�b��F|5s�6���S���֫�5��|?��<-�9^�S��;�q���u�4u9�M�*�C� E˒qK�B|� �]�L���,}��0q�P�}�kހ3w� i��H
}��ι]Rv�WƉ���ԕHf��*���M�,� '�Um�?V�E���u{��Ӏ�%�����A�YV�)"�\�:>�;�e暂O�٘*ma�V�F_}�]�r�� �L��/Q]Bo�*�,�Oz/�$����.�Ul���X�����O�p@]֠�� Z/'�~�I���G�Dp���.��U�Ɛ��Q���Sƴ~�@n�G\?a^v��n�0.]��c�^��Tϐj�e���{�"�|>lv��2c��*���A5��u �b�/�l��n=�u�L�L���T�3�M���?�ȯ�E��6���y�\#۰��Ɩ��Iҥ��v}�D���	"5�Z��?�K>�uS[�T�X�d�FM�v���.W9�C��q��'�}q[�_1R��*��+�� �3�@ ��}	 �a/����>r$`ܧ
���e���C���t��a��I���&:A�)V���q0� �5c~�	`�)��3Z���m\��:�����A/�������o&�,d9X\�M}�����8�@/�]�����X�uZ"�vz����n` 5��#Vܩ_Y��s�r���lX%�E>.%�R���xMZJI���[���\'��`jJ�]�4�iuz�����i4|����v�}!#)��y��k%��So��� #�L���m��"�d�iߢ�@H�����
<���#��< H�j��&�������<[��W�D���Kt�.a��I\���Q���n|����"n<�gcm�E�\����`�Y�oȎm�ہ߽����&з�6-hb+�SU��M� �����	޶c��'�PYU-|��6�*Z��&J�4˭�Q
�wMfC�WȚC��3�Xn0�Mˍ4���R�ԟ�t�{x���t��e������9��c��e��Ţ�6E��.�O� ���X�FIŤ�_y����N�2 ����j�_]v(�������_���y�%|1�N���m�-#>B��V���F�]�ᄜ&��u��SЀ9Vݠ�2�S0X��	�d��.�z5Z=:�Z�N�I�7�f�ֿ�����S ���;�b-��)�.�b�vN�����4����bo����>�^���|��cI ���\�i�<兲�i�I���cM���LV��\=Z��l_������%0K���B��49���c��'ִ*Z���y�2�Z�T��<����s�GC�H�p[�a�H���)e@/��5��C�ϱA�۰�/��j4&��V�K����I]攵��;�����KNP�6$��	�!�e;L�{��^M$7���m�=yql�[�2�+�k��`�c�͊J�j�Ƹ]�(�4b�tmMB.�rFS`����>HEo�@k���#D�����@�(b�:�l���4��=~�K̨W$A^��;DR[ߥD�.��9p�#�X���v'+��(��?O�분Z�����*{���E\l">29��(|�!d'���k6��Id织6��)�"u�%f�l�fT*v�~�Y�8#�(u��b%o9�΋�C�p���>9(~W��"9da7m�w�0M�B�ʹ�2�w��*����
A|�����B�x2OkƳ�az<�::��j8D�unF�r�
�?Xh}68/�ݏ���{�y�6d�EB��	�nl�)[o�vҶo�4�5�G�ʿ�!��S[�i��T�Ź��<�܁W�|4�	�>���.�Y�Qr��f7�%�C�}:A9Mn����i�bw�_whc1��ׂƺJ�+�QEo0�8�Ɏ��R�3`}L$�@r�|��TA�U�ģWn=��>Ie�P���2��#2غwD8��V�Jevl����H���������+�4QzQ�'��'�hX����R���<@�|�$,��b��W��Ӂ��x�raB,��N r�(���H����*M�CU��l�}[�0�յrdwpM�x��w�Qm�&�JiNJ���B�Yz�Hpw%.���/@m_��I@;3��+�V�@=����+�"���ԕ�ݺ��R�/b ����.:E���_ZY��V�
?vZ��p�YR�75.����~[J��d�h�G����HfE��6����`������vqW��Ke=�=�=�P7���aG�4 ��i�B�r�u�3�T�MD_���l�J!�-��!'���g���`���s1s8cA!�-�^&3�i�0$5�H�+##|β��,���'����I{M �Z�|۲�!"��II�A^�$�N)c����AW�|v�9��`��?��w��W�,�>u�V%�߄sM��ԕ�Ѝ׻�fy׷InP��$뽌�ֺ7Wġ����T�����DJ���2{�w���k�|�#d4@xu��?�f�@d��MjrȰr������(�����/Z��A����аԧ��})&U"�~ܢ��I{�@y*)����9���(;A��i���>�q����7�����h�5K�ݐ{�.����ȶ���*Pm����D�P�Ba���x�\j}���gl;F���)�� VNLك����;�"�~��q,�����VÃ����Ő,�5J�;�kQ�L��6 �n�y�o�^߇GX3��z0��S�KgP��PbW�n�(s<�����6�O�&,�K
��Q`��sb��J�	.�����Lv �S�]��%~�Zr�R/���tA�Ww�ZeS���K��/0���D��
TƓ�߀=H��X�dꔿ+�l	���n��)8�;�0;nm��h�0VH0ܝ�� ��-�}&�J�(9s���QQ@˥)A�F5��]��eW��ѭj�f_J2S�B:��2��A����E�g�og��3	��φѾ��]�>�5����`;.O���W�C䁔����2�m�+����)$=��ގ�q�&,&�z�Ó4����il�F
���W@��M��_����xS[��,�q�[�ZBM $�s��~]L�hO��9`#p���`���a�(V`v^q�wn:5�L!6�V�Y��q�XZ�2��@�Aw� �9�5���Ѥ���nCx�汿��J���K�1J�l��T��u��%8��	F/l�JD�w����T�QÝ�}�gˈ�~+UX�iT
���,NM���R���ϮT�����Ɣ��� ��u'dRu��Ka�Q���;J��^��">Q�}�����H�J�&�r4��a`12������y��ꄑ?��E4�z,UVn�Cm�漏�\�`��>ۻ�H4�чxX�Li���C 8+�O%��Zzc:^���}��aC�&�����@鳧/&V���@�We�f��/�	A�f���Y�-�BQ�s�ԩ���ˏR��dO�cV�੅�����!��κ�ջ����	�=������o�#E�B��8��U����>�ɲ��c�$��ʗngq(R� �,�K���c^"&����{�lb�%�.u[M_��+1%NnM.�]�o�K�@mk� T%b�O��RG>!TzJ65զ!��J�sІ�m	-������\��]X�����S0U�IZ��'�|p�Su�����
�F�y��Jw��#�mؖӭ
>eN}K�G~Y���E!6kS�dߒ�ϫ�Uϓ[y�;���qi_��8�pJ�'k%s����,\f��K��-%�XP�z����<�"�?���v��Y�9%_|�d(ŵrlQH?ʏ��g,>{�P�����a�A��3��D�x��IG.	�.6��L�	!bmQ���r�(nҷ���)��,����ݘO��n��V"(S����EI���Xd�<zF���BR�o�tz����-z� �/�T)�
���dBl�'����q��dbu1��ƾ�78����id �X����a���<R�]ɿ\�g��U�<:�����'�;O��.&,�
�?���P��7�����d
� c$�z�����JM��o�.��@�|�G5^�-Rj�r�[Vh<,U�y��A�71n���W�"YP���\K����s�����wޗˢ��q�`B���B�)��Ĥj�7����Q�f��`=�:�ˡΠ�S|`��
� �l��<'x�$�z���D�]	�	Zݤ{4d4nh�ب�����QH�����q���Uy�ޢ?��^��|��]"��۟����-ee{ �d_[؝�ÿ[A�����X�k��DJ{0Z]t�,P�O���6��/���3w���ba��.+��.�,���*L�{�ם7
r�U�	A^υV��g#���K��~���Ϟ���T�b�"�Y��L��t_J���[2�����k��J�
mw����ji^������(D�ҏ�ڇm,e�W�S�������������?e�@� uaX�gf&J��(��9������kF�pUb�v?��,�1̒c��cP���~������w%����?$�J�  m�L�D�*72�@��҃(�C�f��5v~����b�	�qD)\z�):�"�M�e=��Oh�m]��_$^㛜������l��}-�0 J���T��������vN��]���W~�)A�C!z�&~\J��@��2��_t��涳'`u>uF�����sw�h;�}�^(?��m��A���p�=��)�+�����?ᶪ����:�Z���q�%@�����=84;�֞����$[.��7zS�{SB3��1&;��;�rZ���e�9�~y�A
U]_�g��ƣF.+��f=�f��:�Ѿ�)���3w�Z��>bSY�]a�-?P��g��"�+�?"�@�������岟�P��X#���v3��6�/�cq�,ꀮO��|�Q��D}K�~I�R<"8�+y�Xw��	�������z�_H�̸����Ê���
�9S/9E�t1��>��{T3y�u��I�V~�@�?D��?�teP:B�'����ߋ,�LSF�M�����|E���T�F½K`G�wq /s>keҟ!MJg,���+N���L
o8^�詡bCrdf��{�+ᛴT)�K�~`e4��F�n��ZpՇ�%J9o��D�6F5�������<������R���Kŏt�X�)�V5�MG��X�^�)��w��j�u�X�y��'�V�.�
��s�[u�;;���'@����r0��j-��m��a�@�ٗ���|�g�G<DU�Eh�o�̆�W�b��By�K�:w0Tr1;����5�+�\��E�7�tJ�h�K�O�g�!�~�*Hd������Z,���a�li���������.�f$>�|1�cL2�g\�D�c�2��M�jŮ'&-�(�1��$C%����2��R�.�)qT�����w9wc´��
����}��#䑐�����Ѓ%j�Fx�\��!S����s�w�����J�W�9x�r��`�?�t�V�r�fSλ8:3Ri��[|�6*YUZ�UA	�E��ɤ���K��a"���~F��� ������V��ʏɸ�M8�Ya�0�����C��wXh�\���[e���%���F@�~�m"V�x�O�Zj`�̠�X9�%eFa�p���_|&LQ쏟N���P���K�pr��'Zz񗘫&4�M��U�̖�U� ����<q<O"F3Z�
��'�U=������	j3cΐ�����d��-u%h.#=�:1K��P�^��񤳹zkO�z
\�O6Ք�N���^5�!���[ � ���1�u����VЃ������H��t�ƅ�E��+V[��fi\�ٟ��(�hbw0��ynd�i�l�\�Ky�8�Qݵ+*��.�k�Q�+��g���/uW~Q�2?7ܥ�R���|q�L��]}y.2���t�6�W&9F��Gqp�]��A�M��	�0E�hV�!Q.
��B���K����T.Iy���<SNb�s�@k��>����^u�������ģ[�0$����AvMZ,8��cY� ����4hT�C
:�"�7�����o��sAa7!R���W�m�eA}��h�Ec�u��
���L����&��وt@+�'�U���,�.��$%%��'/�q��JBne�a֊z����&aO�6Gnp	�jd1���e%�+~>��:��#���5��ĺI�٫��J0π�/T'�/�BQ�Z��8�p����IZXT�o�O���Y�J��������ӏh7��H,��@KC���tާ��ˠڎ�)iw�H�����H`m�,+�/�d��-r���l�'|a�&*!�!0�4��}�p
�덌�	w�8�	o�t)��e[�B��ܺ|�ot�DҾM��by�2��B�<�n�$�$��j��օ�Iu��[�C_��'�|�B�ᇺ�4n�=L��/���4���Q��Ap���F�G����h!.8��S��ٖm�U�
���RkÛ��Ra��������/D��3ы��"	z@�,�}'̛���1=�(J�Ү��A����Xv E��_�4j6N��cԲ��>�!p�O�'O���XY�OY���Q}a�nrnf.��_*�.[� *�g#�u�tsf]'E�Z���+����K2�2������N�'�m����t�4�t|����!�7蠂ة�?[���Qb=��_��s*:�����q��pL��i$z�-�o��$�.�����H�*Ux)��ۈ��}b	b/P����0�U07�3�G��h����Cۇ�5Y����f�/���3�g/c��Y��կO��?i�.�0/���Q|�<���0���e8�s�����U}J�݂r���M&�x>��>�0����U���I�)��;G��X�)bn6m g8��n�����A�L����o�՜�@��V�e�q5�Qz�-�N���J�,��#��\�`�,{��B�IgB�����D��B6�*�4]��GI�G�����]�Э	v�<]�89�2L��xE�Lq�vl[{T�|��>`\�N_Rba�����z���&�eU���zI�c^��:���w�͑�3��W�#��f����m��M�z�c����k2i�)�/G���q�q�8?�۵z�1�@y�b����WZY�4��+�`ۍ���[�0(^X���%]�bߓ�5��C��
�����_����2mOU��!���ZI�V�h�����-��pH� :Ź%̪@߬�rL��ᖳ���*��E��̋㿒I.M�(���l�r���!�x����A�;���k�jv��҈��h���$��C�tJU�	zĚ��5�bN3����)؀��}�3 �MƧ�@���?ㇲ�d�e��B�P�ԯ�YW$X�J[<�5�)�F���U��Չ/�:@mg�K�Y��V=Z6ɓ�^+�v@j.�F7p���#�.��эPd�`���8b���n���1��~�aBZ��,hk�C��m��ʐ�}7�æ��%R��3���N?���A��0�*�ƢX9�$ҍ��k��u��#�7�e�͵ZL�<�O�Ęa36� ӂl��i)��P40'M�@�&��R�怵����:]�8��m�^;uP��n0�b|�m�r,�6�&�H�evyݡ8�N�������%�$7�������/c� ӂŮ���O_�W���Dq��!DDUG�m�$ǡXȴ���c��n�}��V
@����OW�Nܡ�H`�\]��j��bQ[��]	o���A��þ9TN���.��F��| �uk@%>ĺ��?K��.����{���އ�X����siL��41h��D��U��hqm�=R3�=�:i��x@�dUsV��Y��k�����3Mr�h�z+5� �c�&Ҥ(Ʀ�S�QF���RV˕�T~��T'C��α�Wp}3����<��	:�Q3́�Gj�R'{�/�����h%��I�jDTT�
Yt����hz��� ��d�c�j�rq&Yoy�Ɏ��.#[�h��a~ߣQ��̲*LL íܒb�6�&�w��-|h�L���]0(�0_u����T�t����`�_��xn-�ID��&*��:���Qw��s��ZTߋGh��
����e.��d���.�2�4B5D	H�]j=Ҧ[�0s�Ǫ2)���* ���������SHx� �
����8Y0��|��np�ihd����x�1��׺)�N�+J��fH������]XY�����c��;�;�T����?[����ERzU(�k���	j�uEZd��OMG�Q�tп���${~q21�E��b��g5��f�!�i��b�u(��z�ɮ��UsI��r���p�e�f��sǝRh�0Nx%w �GH�vg@�o�s�ɕ���7��}�H�Զp�PiKp�c]�.,�o�HM@w"7+,k%N�!�X'Ε��oG{��`�.m/z}&������+5��~���D8�* �kh���s�b�K�������7�+5�zf΁ ��QU5�̕{�x �B?�ůs�PF���d��d��u���9�^���*m���VW�p�m����Y����
�����U8�>�	`��,�~�����"��h{�R�-Qy����fBVB-/����!�g��s�����t{j��QMDm�(��WO��x�oo*���� �_�<��wAߖ}�U��.Z�	Z��8F��R��{Dﰊ"d/��_ߙQ(���$�lt0J@�J�O��0�O��~́��+�)H�rK��G��Q1��,�xH"/�����G��7�XBݿh����
tZ��'h���Ȑ����ʭ����_O�O�eC�H@[ͷ^7���K�i��EH���G��=��*�\0�L�|��iK��:�װ�I� ���p�7���2�p�#n�%��L�{
Ov����_3�Q*�r�9ǯ�X��/��z�~A� `'E^5���\������_w�+�Q��/xM�N +R�(!Z�i��ř･rL.Z��
ؤ��~R��ډY��2�~3�nx��z5�t3f�Nĺ�#v��CJ��PGܝ�ˢL\�$xn R�Q\[��R�>�.&�����o��(��֧�*�0��}��#!E���@����_��6����]V�-���vd�4���ˍ�Jbx��l(9��Jaz�C��2�(�>�%2�쬯���GiQ�ɑj�v��H>�����.�	�2��*( }�H$�D�7�~�`����C� >�uj~p���T��֋5|'A�G�_�N̦��C��Fzeuw����4)�w�t��M��jf�}V���H�VkP��?9���ǹ̴��*L%:0�s$/�.�E�"2e7�Pe��:.��P'��#א��,ӂe�x8�x�P ���0��&8������`xz��cY�L���,����J�)K� �$]*��u����-� ���E"[�/��l-X§����z\g�н�Ɓ;������uՉK	Wh��#Iw"[��~	#��Yu9�O�p\��'����'ـB��,+a�T�I�9�V���.`�G���&b�ͼ�i��6Ec3������,˸�2}�?ZB5$���g�� 
�~ω����h�F��~��e��`>�=� p�:� Y{�����)�43.��^
�İCM��@4M_u?��)�DB֠&\�y�<R��7�ל	4��5@~��+�Y�ߔ��"������(�E�L� �J�H'�Ej+���:ɢ8y83�V1,�^�P2}��)�lฯ�\���U�sUm�;?��f�����e�+{�&�	E�Ʉ����.QJ��h����;ސ^'�ɭ��e��I~���ݩ�G�+���l�������b�cї��ۃ��P���o���)?)�D�RBm63�d��!��8k��=����(���9�YeD1�HT��o`[�)Q�Ś�{��gw<9�uW�w:$[$�7�����kjR\V�^��u�M��Z���z�=ſ	�M�ۙ���;�{�oy����B3�^1�v�]P����f[|z��U�ٶ� �k���j���z���dh��˅���p��M6`�޶"7pԹh�+D�=��OF��^]���Q#yc��/�H�O���M�s ,N��,�_h�`�҂ P�<`����ƞI�l#Ɖ�jȉ/���1c�o7c01�u�u�s�[���|��?�o��C��k�y
3�Ӝ�ȗ���d᝿�_d�Q��QCǴd��w�Eu(�L���0X�7�R��㘸nJ�Y� )r@�蠚�eL�$Ex�������G��h��Ƥ�"����f��׺H°#�?�^�t���^g������H�?��5���[�}�#���÷j�Mz�_{���Ȉ�Z�
��ݎ�S���X�;��fnM���
 <�)[�%=�V�.�9��]y�BM��a�P��Э��l�1Op�����gC#���9�1�V�'A/KK�}�C!=�W�j�(Z�'¸R��u�v���w=�N�Čh�\p�jƵ���$p�^��@|4܄�N��)^R�|�%�W8BB����.(�~Upϱ"Ü���'A����V�UN��\
�	��#!��?�2�,&���L��.������O�_H�ٯ��A�>T��٠P�릉o�tu}-�X�y�J�{O������Zw�'&Ε¥���ҧ��#E�!-�u��Ѝ*�D��?(3����c�Ҧ��*��(��?'R�(|W��|�9y��y�9�8�}�&�O�7iRJ��Ƣ��Qx�"u�5��zj:}pֶ�`���BN�����?�H���"ta��S{��/6-|�S��w�8@R#�5�T팳�>|���m�-��z`������-�PR��=��^YzOVݴl]!��b6 ��QZ�0Yk���^��MX�F�U���g��$���^p#m�k��LK�y$�"��ye�OH�o����
�qS
��3��u��Y���T�s�l4?��X���Nv�7� j��Q���H_K� 0`�4<��X����c��Z��6@I@��F����>sm�	L��b��D�?,R~�-A4�����8*����b��Ybl�i��'�4�� �,�ذ�nU�D[���8Bc��+F$P�r�l�rЇ�x>X�6}�!�_��3��P�u%9A|_�OY�F�:c����\A�1�
���l17��t�m������wS�!�u$AEJMض�k_l��΁��`��N�&�	rϛ�Y�i!�����n礕<�w�i��;��y�B�-^y��K�`����-��R5��4x��])��\;�oW����}���n��3�fՉU�L\-q�P5�!�L���&2����1��la�5��s,X�SGf��hv�ŎR�tYJ��`��7,}neW��ڽ�XCǆrq�t���k��S�y�
v����w̓Z{�3�|ͭCk�L���Ak3�Ɣ	��o��z�`���Xo���K��zt�vT�>O�^��I�2����at����G�oq�N��g��(7R��G���w*�Zz��tK� �~�q��v�=I�H�,��g��p  ��䰳s�����57g�72Y6w��B8CF�!�1�E��,�˓r��HAybHP��O�9�A�����d4}.�~_������	Q%�,�so�'�k��6��XEQ�#��,:��^��01T?���u_[N�{��-��<ow�:�#3�9��L:��gKP������T8%�p_A�z�j_�%m�C�\B��`yiv+v�w��T*-�@f���l��[��B�d��&�Q<m��j����½���ʒ�_S^�G�pU ���ď2G&t�R���w���cj��UN��
��:���.k���/`[5&0�����5]�.�ՠ��\c"_��4Vm��Ơ��[R�s%K��%�ޮ�}�J���k��������_�U p��*�R�������I�>l�U�4@`�d�	��_�@�V���s"Zj�k�~��e�u��*���5n��`bo@�~Պ0�;�h�֔��H�M���O#ޝ3]�Tlm���y��S�h�Eꎩq�?Ȩ�Χ6`�_^���\�b˩�͸7��r<CΜ�7�f?B`١27ݏ�v+fw+�����f��M�}/dgO%�$ДJ�\��KAW�(�״�͵>I�
u�¤�"��Q=r�tʳ��$~(y���e�`�1��Q�Nv6���U�p�@]��aI��`��ꭙH�{&���{h�7YxM�q���"j��o�ܨ���Xڡ�Ǚ;���w�@�RJ��h ���f�l�H��� �deK�s�p$j���'Ĉd0-ŀ)�9�zpu#n�S�C���]Z�XU&�ǯ�����Oj��b���z!�>9����p���0��5����9n-�{؟��do����^�Ÿ!��o�wB�|wI?��V�x(V}�Co3��Z�"��6�0F�bK��g���|��J��Ǝ+|��?��Z��z��J0��LϤ��
Oo?�����2�ь��K��(QC^�@�ǭ�Vl04�m��j�w�ƒh_4���]�'E0�~!m|3�j�ǅ'k����S����F����RT����Gf�;���6qO��_��'�����R'5�^9��R�� ��J+�"�
�d�0ڃ߇c<ҭE�;FB���]���I�5j�Z���JaVT������d�x

"��3ri�
�Y���2a3����"/w��,�j��t�p��Fr�`�z�E+���!��+�o��BS�����Ó{�1EG���iM%������b���V�&
:�/�]V�!�������#|%����U�D��>v"����ộ+'���0�0�\l	�𬮺�	`��V�k��ڄ�w��׮/Job�6y���Z%t�<�L`�2lZS�_V?!��J:�������E�(�����S!��e�.pc������2��m�����I�t�c$��~i1׳����Ⱦ�GH�]7���%��O\��ٓ������fB�z{>��i�	s�?�I��r_�yYYXʰ�
cc���PÌ�����A��g[�6\C9S��=(Bz��<��lNI�M����a��ʽ��2*�#6*υ��.4����k@ ��ɋ�N��ݽ6������'c��]c���'g�
;d�w>1���zM��<���͈tۥG�K?�'�.
����Kkz�=�6}��=���'A�� ��CFHԴot�,ݒd��m��8u�=*�FDk���V��Lpɝ=����p�t�y kcQ�o��F���*g�2l������k�����ior�13R,}������7�)v�bm{@�'&���MP
�
 S�dնp,)������E�S��Ц���o���۸����+ml9���W���d��H�����G���`U>�V�S	"(�4�q��\�
��g7��hr<f�i��g���.H	�m4��x��%{̴`2��\�-���$HY V�c��q�/ny����0������:^5�t���Tgr�J�./e��X ��iH�����g�;Ƨ>���·��N�N�ːԃ+h�Ǩu8A8��������|��d��E��S��2�t�������r`oD������]���1��1CϏ�gu���P�."r���B�o�����!�(����f�[�-�%g���s�-�Iv`g�Έ/\� �M��FTi	k�e\�d��o9O�
�݆�@s�DL@���)%�oҍ}���Ӗn��cC��P9!�� �"�8hMx�$��W�=wy�yֱ��?�cz�2R���8�2���@4���~<����]�����hFc���!!5�U�:��E�ON���k��J�����A�^+F}g��LidO|�s���0����,2W.?���6����L�ن�V�
��M��Ŷ��Ι
�_�F�y<�:�\m���H������NLҋϰ��e�(cxC�� ˋ���լ���-���ol4��������{Nz�Ԟ8%]N�,��� |>�e{�{�;00��Cj�Rr|R��)�8X��@�JG� CkH�V���H�crׄ��¢u2�� �H>�P��%��dk#�/��:S����!n5�6���e��ͫ}�'d �j�3BT�]^�r�׫���yk�W�;�lrw��)H�^t}�uyƴ ~�^J�i�c���(��ݍ�^K4�bh[���ɺ��mr�������dA�z���R�O���;�ON��CoY���d�#2>��2�ڨ�U��h�	��&�5���v��a|����$�^Tq�al�;�W��Qf'���m"\�{�lK��b�X��j$:S��� �W�|b�b���M���5ҭ���:K<_��t�~qȲ�$�77Ҝ��/5��͝��>:-�l�|��.a�3J���k|�A^��O\0Q�x���YF7��,u�v�m:H��/�c�߉��ߚ"l�{l�h_�jmw4��N�5�X}�x��6A4�z)���i�
����W�����~r��� U�BT��3:x��(J��>��uZLoP{'��t�J!x��6�o*����fO*+��nbˠ�R(/���-�RX�镭C&,o�7͉kod�$hiۡa󋄏*5�~�l�R��sh<r��,qL���c�@�̍�w�"m����]�ٗ� ��ɉj�+�F(���D0N�	 �����ܐ߀�KCTE��g�<�ߝϹ����"u}���%Pps��=*6���u�_�t1�*b�͗�)�� j�GҰ��� 5zCk���;�[ȊpY"�h�i$��Ԅ���/�2Ci���
���)��Fb=��m�ic�Pg�5�$7�����m!�����<f4ʨ���y}�C��f�LL1�`��ހ���ows+76� kO����rYq��T#�?��rY7���ș���o&�,r����5����&/إ~��o��/I@t"5b ��/@��������맗ee9�"���B=��2@��w�F���#��_�S0a�6!�y���Bf�5���[}Ɔ9�/�p�Yb��|s���Ν0W�c[q�WV����g3p&���uԹ�l��;��%�O�0�<2�=4�`��+�ף(J�M�н�Q �컖�ע|K᧻������ot#c�K�r7���j�jR�������P\.A>�
��zTY�	���V�m��d#��1K��/��>*��jt��p��g� *�I����\�Z���|)h�U��%lN� �(ea��Bؚ�k�z�N���[D����`�\d�V5��� ��ab2�o9�	�-��Oj�M����8��0C�_?߽�	��T���%�����5��yG����3�\[� WD�<��� �{���h�6h�C���or����[�=Kp���@i2~��G��䏐�B��&⥷��1Z���g'*O��*�C> �$���#��"J���I/2��4��M�S��}~���,�q#q�#���E���o���![�"ƽ�xڍ˧��<f��mVo,��d�J"�S$WO9�%�,��s8�&COB\0RU���|��;1�N��\�d<q�����-���Y\e��a���K�/�'s�!�}���6�ʅ.lM�K��!4��\�F�=��$�o��?
+Ό=f�^��/�#�b�� � ��ΫިG�q��w�3��`�-��6�4�&�=C�z ��ʬr���Z��emøa]6��͞�<Z�v�'�*%�GG�������w�&��PTU��Yi��w�4kn`.*L��S]�䗥�ӓ���g	�|�j��s��+�-������ ��ZbLB�D���}���^�#�6���3�5�z�*�XQ|���E�����(N6�1����R��ś�7�4�)�e��KE�}F*Vm�1�����PT���p2���d��j�'�v��\����2	$=�m�?�'6�&o�zR�N5řwX��W$G:�Z��h6bG�$%���3˪�Ѭ�\��B���jś&�?�q4?[C?�y\�h�z�5���$��#�:qh�ÕKS�\���	!����k/�bp��g�6^|���]&��U�?J�  o��5��C[�+����T��U4������~}���],H0@�c�g�@'�(��]�h�bP/2T�b�L�9708�0k��7��A�u!�'�;���!�E�=�w�}]�7-Gѵ���D�7�7>��'zd�.�c�D��Qu`5�r*v��>�6����X��_�/��&Di�~�k�U�}˻�D#ѻ�ID7��[�կD9���d�*�Fk�?���!��9e���f�K�_}���Z_���6�4'{�b�P���w]s"���s0��m&{oZ��C
95e��+q���G�UZ�SW݊��d�j��2����W��.�#����Ml�B�� ��ΰ�Sω��(:�8 ��r�A���H��q���ѠUz����In��Sx𮥹�
���yأţ�-z�9�{ϥā��/0���޼jS�71��pТ�y���&�UemC3Ǜ�)�R�=�"�TP�Jz�����>]���Ӭ��p��;���V��a�d�H��3dO3�/Xg	�0z��5�w��G�ѿ�D�f,���'#�<�*���]ňu����Qe��_�r�-ah:*��R��'v�]�x�t
�a)�m���0T�	�dXvPd���&l�R��m`�//���
,<YK6d,>_����R���4��}y��O��ZU��{T���ƶ�����8 ���O��k�o��t�I� 5FE(y������|,D"
ms�R�@�-��}��K���MvA�ݴ�O_UY)yo����n�����3J�-3m7ؐb�N�d-mas��`��m��@7���s���HY�m�]uQ@^���(����-��Mri�<\m�t��Ӵ�¾R~�:t�*t��������D)��h����z���஽��f�DIu�p�<^�I��7�y���<ْ�0�D<��gp f�?h7�{�Dnׅ����Lp����l�TM�ep �k��*��B�������XQf�TͿ�i�v�8���y��Z���Bf�!��R؝:ȯ���@v�Sۉ��89�M���P�3���)7�N�LW�� �3��/<$+�悐�k�C\n��� %z.Ca�oK��-vth���]kٴ�
�O��D�Z�aX�E���!�*kav�-/*ˣ�)��e�x⃘"eD�<E��K<���oL+�P4C��*:���&e�� i�dZ��(2�{O��'�T�A��<�URg<�蛓��9ɪ�zK��H�!�����C�;�7S�j?F͎'�8i$WÜQ�<wV�}c�+gk�e1���=~�ߜ+�zT~k��(�n�Cؔ�3��aU]��#�V�8������3���#T�s�z��T�d9��m��m��e��q����1r����E��M�L������.V�ܟ�ZN��F��Fiy9Ie6"+��ErH�E��`�+Q0ѥ�ۃ���I�\�3�92��8���#��b�>�Rګ�%<�;�ګ���;��ܤe9������&��"!��QØ�\�F��"rf�c{J��Wr�a�51O�9h }͸F���I0&�����ص��;�=��e�Y��ɻȝ�C��mE����\���g����1"ňq��qKɞ�����<���`=m8��VF�mus1�B"�}��p�x/�]7|�^������5xX���}e��y�݉�|�ѺG��f�������F���7Ő:a*R�cd}��՛�����|pمt�N׉�se�5�4�+D��
`�. /o��C���S�RA~ю��,�a|���5(>I_D�?AQM�!<���Κ�[��)=�@1+�+15��YM9=\+��վ�Z�BdEf6n��/�1�@Վ�6؀Y�����dc�B:�شI��R�Oռ!���(�t�8X��Pc�7��R	~-���^b�>b��\J�K����l�T��~�H���J��\�vu�"��gi�!���6X�ebc�?a��;2סk5ﺎ�z�� ��e6���f �����:b���穀-F�L?ܲ	�X��?+��{6�iOt���>�>�'�i����oR�����z�w�#���cXL�,�Z�����o�A����6 4dJ���"E��e\ kFM
W��v/�p�c;��ڏ�_=n�)E��ˌA�Id#�/, ���C:�Q��"�D5Oߗ��mH1xH.�1m�	�i>�n;�NM�=)���=�]�p�5<ͽ�o�{i=�?�3r�^H�Ӎ>��0.P�9�g,Bi�S¯�O��Oc�䔠�R$Qt�������{�t���|/�-��5��`ĩ���:E{(����qc�6�����ڃ��"�O:�\��������p�*+�,�d#�m����x�P*���'@��Ԗ���>�O��y�NKk��]��Ʋ���L��M����R�\���'�n����·W~��b�UK��O��.����-M�@�*��B�;�~��T�ڗp�L�=х��R�v8Q�����[�s�$+��RE�r9��k�|��@V�H��V"�"i��+ьBn5 ���A��@�	�hp¤'�-��}@=M�R lg��mL�>��	ڸ.�GI$=�h�=��0�"D;�F}J�ե�q��̸A:�x�T<>��%β�"3��=ᰱ�>,+f(gc������J�� '�t�E� �RL&%B5ZՉn4��$�-0�f����R�8Ib�iAP�f���������rWJt�́O��A�HQ�����R�}�l�h�������>=�y���O�/_�d�@`���i�O?�`ؚo�8�*� ���Ν�#�\'�w�Tɻ-}}�\�M�r��gwVq���k0(0�Z
���GS�{��>��vf�x�w�B�Ň�H{ ��+�0�d>#X���R2Q#}ǀ���C�6CV4�h��%Z9c�����R�p������(���מT��. ǵց�|\'���Hl `�ʎZ�gþ��Oz�mS��e���^wJ���!جT���1�ZQ���#}���%m޾��U&�#���q#RD�+|w�����E�ڒ���6�w�͊�����X��6v��{������N%=㐲�O�R�ڍ��i��`����� �Bݦ
�8��έ�8��I���7��B�"r/W����*`�����-���R<Ŀ��.��A7a{�w��h�>��
�������]���l��6�	����,�]=��ƺ�S6�y��ۮ�x��*���hE������⳾�����+��ax��[�ף#�����w��$^!��FBe��ԀB�y�l���*�U�ղ	��2��<"���=�k��M� �;�T3��sE���?g5�ۅ�E6��}��̬
I �u7�.��S
@��t^w�b��X<$�n���Ғ�q�������7Ƌ=2T;@F�>��<f��4�s�(�}Sh��3��F�u�یʫ���$�h6�Ϧ	b	%ĳ�F��|BV$��5M�N$߻��$G�Rm)���[�ݴ�K��;����gM$�D��]z�{�y�s��Q�zX]S�*�}L�����V�]@��'L����!`#ne>L_s�ڼ��CH n;�]f�'�7x`⧖Nx3A�z��e�u%�iAJ���}W�r�Ώd�$��N�g8xh��8��"���Ϡ����<�	�l(�
zi`u_��񙜴Z�xE�����JL�.2��w�8�jD[	\P�خ�3�J�~?�S�(b hq��Ia���|����w��˚��z��Y3��nj�����C�S�v��ﮰ D�v݋�1�c���z���H�ta��E��闉1���r�TE�	<C� �Q�S�Q�)˱ ��v*���C�����ɒ� ��8�}�Dz��?�5��]��r�H!�3<���_�IZpV'�0�<r���3��~-��F�|��OR^p��4�|ڑ�jԿMZ�W�L$	@js��QT0UJph[ɟ�Gq,�����B�]����L��nr%$hdv"�zT�x��ی�yV庈c�Ϛ~n��O�&�_���Ҭ-�y�!�K�������^]Hu0� A�n[�/%Z3RE��-'�mo�3)N�>������IJќ�_��ύ�}�l�IV��VZ�ݧ@��ү��n�Y�ܲyH��6��e��*і)��DD���g�+��W]���"�pB^�c�.q]�CpK���vU�Lh3��W����jz���8#��]9U�4��nKH�Q��ݲX��M�M޸�M��b��j���Ìm�A������l��1��cJp'JF:��]�:)�����e� lR�/�2��R����S������w�H���.��s�ÄM�P�g�F��ȿ��Ֆ��������~�'l0~rY�DG�(�\M�mzc�+b6�/�W3"��:�-q�J�XwIE\e�����W���Kܴ��@-7+m��jU8�6WPJ���fs��~�3�4�Ƶ���Z�&8Ho�g�lňKEo���5vn`tD͓+�������������.G�Xc�@9��,4�����d
�R�i�6��E<��{9d�r�@W�:�)cf�qa�\nO��
tj�r�5pP�=�m��m3u"�~B���]�Mz&;�]��<�㞻��"��L
b�^�����R!�sQs�޻F�ّ�X�K�����D��@��Z���Σ.�	1���-6������^�߰�Z��R�F	*��0��[v���b���jUh�/��a$S�C�d�����~0��V�Mn`�O�t��i�5�j���4��ͻ)��apW;�.��R��<�Lf��Z�z[��֕�.6�7_o2��\A���c�bu�"^��jJ�U���g8̼��r~_E��s�ʘ�ۆfm(54M���\�ڤ��6;#盨��=�N�VD�Bì�-�����=7G�e�:���i3�k@x������Y.��í�	5��W�'�n9�� >9Kָ2���Ez(	����ќ�Զ��0��y@�"�Q�w�@4��ѓ8�vY5=t��C�g���^B�3�d+ӟ�ګ%�c�.L��h�y{���Á�_�IL�o��N
�6�<'��2�q];-j�>w�[�.�ݷX�e!@Ƃl�A�VIP@d���y�r�s#]v�3�MR~�E��h��gfB`��g5��@0�<"�H}��$��B@l�d�ںRO}�e��-��b|\�ӑ��$/B���{��@6������\����-d!{��nӹ�IT�GnWl܋U7ڀ���e�j{k�# ��X"�Ţ8T7��H��؄%y{S��\8X�Hϒ�jfU�maz��@���v�Ń00O�����f��V��������|]�g�*�LU�m�7m���ԩ�F�-�g�(����4J"�o}L?�@Z!��Q)���g��L�{e���׮f�AY�3�C��^�؟�>=E5ir;vT �R"���c��,A�:Bt��Uގ)�Z���*��l��,��U#+<��Q�03�����{��xa+���:�s�s9o��sQ&��5��Y�B��EwK���-q���}E��H�/�c��v�[ۯ4�;w��~��W�;��euJb��6^��^����2����a��2�ރ��8�6��T=v���-�zbʧ��Y�+�������y�fȝ�S �I�q�z��@�DQX�'M|�@}��{�W��[켣��iW�c�2iV���ѐ~�6�&$��F�^�q���}$B���Е�ֳ�\���:s��ˀ��D�A��M[�g�0���?��OSK`��
G�H?p��>�h�(/��m��H�6~gO���0��f���d��2� L�:?�����h���G�)�jw�3�.�>�o�	jհ��k��cS��>y!�j ��l�{�[���O�˲�p��`��p>TZM2J��lpX�;$��Ĳ^ʗ��"��nZt��QCq����T�}+��s�}٨��7 �8�`��rc�qXb��V��Ц\�8�9�"���u2�䈼 ��2�Z�}4k�!�rP���� p���b�wfS#H���k��"1.�[d}"�����?H���q�D�pW�Α�����|n�H\b0�a�K��6D�VØBz��|�$/M�+|-�Q�܄\�n�@�H�6|�����x�{G'`8��8�9�Y0�D����J4�>��XP;'��F]%&���T[9���2�6om�PK��4x.������|/�F���n���]��O�N����.�$��n�����H��%����Xg��$��{rB��
'p��&O%��x8Uĥ��cb�O[uxiv_cO�ꟷyXY4��F��,���kڜ�#����d҈��ή��(�j�bp���H�|�Y�E����Gj�`VN)O�	�ə9c�2e!y&�`�	�Q��y��7�����M���!|goc�{��2Q R`͏�v��kz��� ��q��o-�`�W������j�s}{1��HWs�]��@5�a�ȷ�ĳ �����*#�.�-�����Mr}�������z�̪��N��?�w�:�Q�k��|��.,D8 j!����Jlԍ��o��08<7���Oj9��Z
��sJ��ѪzΠwz��p&c�n̟��ӫ	��!�u\�LT�=W�2Cvi�s�����p�s`�Qĭb�Z�e�ۏ�&�c��(aV�������w���;�ߏ׫4��a�(VOG�ϳ��꘳G���C~h��E�\�����& 3�f�ofo�� L�r>G���.0��v�a�f��1��z��=қ���z� �
�δdnE��'ab$��e_j���qC�m���M+Z{V��u4Ơ�>�]��u�Fq�٢�ХOl3�=�!v��,"ˍQ/�A1���/W�miJw���Џ뀦�Ay}�s%���3�o'�@�7(*�/���H���r�P4��QJ�]�a��'ZT�c�����8i��8Dޒ�uH��x�̯@����e��wN���s�w���������8�3��T���f~q���Z&'Rz\�A�u�@>�� ]�Bj��	A�D���u�P���ffg�v-�T��x�z
j����Y=�Ҹ�[v�ߪo�S�
���n��oO Ҿ�����+�����a��9�:yq�����wؾ���*�K-)����K��Wm�o��5�L�Z�1+�IK����#�_���E���Q�9����1��ٛ�hf�L��"�JG�|�|ѯk�m �k��X~�`46G���o�p]0���WN���C1p��*���A�X�(te/���J:W2���;��\�P���Z��ˍ��r_m�\΃��~2�w&-�h	��A�Mka�W�D��+���?|�K�B�X��X��D�87M�p�w�� �x���+gu������M��Fġ�'�?2U>�t^8���V^�(+�{ !)(e��|�$e��ڨ��
b�^�k��*��#�d�2L���4�MK���v�6� jC���Þ%��Y��Si5�8����yH�%������s�ѕ���D�@j�Pk=�N|�LΛ��>��J���@{�{;
�$~�4���֑e{Oi�ڃ�j�uYI.8�P�n:�}����+���Ve�3�5p�;O�d:�+jڮ�4�{v+��H2%{r���%j��99�(���D����/�{���f��"�( ��hI�	��逗q�I���ƹ��O	i6'���dܗ�E:&]|lQ� ����6yO����T1�BY�Rؐ�/�o�
z�7$+�rhW&*��Ed� )*�~�+5��qH@���*v�e��}��Q��e�G|r���m93�qO���.���`ajk�����2��.3p�|7����4Y��������3|3J�/F�L4�qb��!�悪�v�[u�Kjm�c�� �8��9�ua
��"I� ��M	1�[�$�m҅��V�e��]����"&��R&���?^af��|���O&��&��!4{�VU��V	��K�u��fۿ1�P�����E�����-ޙ��~�V]A�%|��5u_jvH���i�>�{f?��7�Z_:�P��h=��:�s�u(�w�/��ҝ:��$���F=z��ė}Ƌ�HE"U��݊����a5�/l�[�w����	�R����Xi3;��v�d�f测�B�Bƹ2���2vf��a��-&^p�ٔv���}V�[��C��2`L�p���W�1tJڰ�Vx�H�Z���[�ov�S�\=�	��M�=�{�Ͼ��P�PN�0O�Zک	��j��v�;�MҒo�}+	��KR��~�f2e�jmp�Β5�t�L�h�1\`x�bdҊ�U��R�!mO��G"$t,���fH�-o�6[������8
^|叠L���lz�tݦ@�S��\j7ؗ1?��9R@i��
?�Y�Ȉ�|�r���]��:���3D��8˰��a�+{��9O	NF���ǰEL�fS��A�\�{���B�V��;�`����WC׮:.f�-�W~$r�"d�s�dy��5mb����P��\Ra^֘�Q^�7Κ����f ��{n�F��f�wl&��@�d����k�YԩP�S�xȎ��W&C�9%��U�E��Q�p�]���=LcumE��{���/w��2�j.\���IM�L��D~�����q@�Ͼ̼<z��y�|�X�@��*�k�w��vY��g_).�͏���A�Md�0��#�����$�S�b�Pn_,N���R�b0������� �DB��tC� .Hwk��F8r� 6mOa�+Ѽ c'��H�ɤv�`H���":fw�Gpy��%��+S�튖j8m�"�ͩsVOS�ar�fG�{���L�x���B�nnh[l+����Ӱ�'��P�z�6�P6u;�'�u7΄�z�n{]�eR���MI�&�.P��X�������d�I�2���!�"�g�s�q�M; #��'o5��ԯDW@1��
-R^��4����vl��C�Sh�����jY�v��W^�g�й,�G���[6�w"sԜ6���B��'�� $�C�&}������Ǻ.�r�.Ay����J1~��f���3Z`Bb+�aG�3@��?o�W%	X2�'��r;�ơ�k�<@�&�VKy�3��3D+�𐂲y0�z,IL�1�MQU���aZ�x���&�d�F�ėU�L��
)G�l��*�-
z��տ�͢|@�nSt���s[�N��wD]h8[���ܫc �����=0�_��լR��\����>�W�$Q�!���Î�%-�U(�T��{��xv�����Ϸx�Gu�Y�.�x��#���	d�d��q�S��;�>Fݥ�|��x s�sa��~���$N7a�`�#$��&<�E��<	v�����hσPwH9�R?�.������y����'���P����Z.�H��`'�N���Id�{ r�N�g�Z��>m��Z�T��j��3�q%9
�/pMQP޸�q���(\��vr|���F��G�C�p]rq���C	<wdX1�B�7y&����ElKvKZq i�t[#���8��W����OV�����B�&�R��`Zl��ůA��]�������k�;	�p3E��ʋ��64H'^_>�Ξ��8�q&Fp�	�`C�x�@��]����˭3[b�,qVS��+N!D2#UO@�>޲@�4Y$c�����-R�g�r�"�D(��i\�v�{,��9&RY����B��k-�0>��0��ZC~�:��@�[����'@$[��e������A��l�T�����JY@zV8B���	�)�~��w���$�����Z/6�̖���ǒ��?������_.��P����ꤩ��{�8Ⱦ1�=��̐:&�[���+�\l�e�b�&�3ٞ�E�����l6��N��B���
�n�/J������%)�2�%��H(����t���e3��k��[�p������½|G��]�F3��1�y9ץmgj?#����=������~��rbd��q,m�\�+:�_X�xM��"��ѥ%���p�?�u����� �@�	 �04^x�1���e�0�7�f�G�x���A��G���QQ0����W$��%�ӵ '�N$Ċ[�ha{L���Qvz>�I^�d]�p2��+��PU��h��J�z`��=���9��L�xN:������kP{7�6
����[�!Az0�	x�S��#�	N!Y]��[��>I���ץ�K�x�:N�\���.�R�0^X���p
�S�̓Z�9��Bz�&��k�M��1$��nl��g4Dʪm��xy�6Ճ�In z�E
�ဗ����}Wf�\ĀS�論?jAA��CY.�RҰ۫�1�7��gf-����q�lJ��0��4���	u(� '���w�tD2�:NC��*RQB����ټۓ/6�re��a�lz_V���J�i�?��>�t�Z�+�L���t5<BVO�)�+8ӐQ��mzo�bI��HZ��Z����DE����m��0��(`��K�0n1<�U�ޛ�H,�S�gz�������;U���d�/R��;�B|�����k���^&1D>3t�>9$�YЛ2�HG�g!j+�K
���JM��C�3"� 5�BTltð���옶����0]q�R=G�d�uj�2F�3�rcl���h���"��kr��C]���7���x��:*�QBT���$��.#."�ԛ�$����)|��X�&QN��m%�F��F�r.U'��hX�|��bA�>�Rf����9��7��@���HT���;�`-l0�]Ѵ~�ψ����x�*�u�M�`�,�@��h_]!wݟ���Ό��(�]�c8�ܗK���q"^F&?�`�Ϩ��l�nl�D��(.X�h\�aY}��b�be�O�� /��hL��l*���@_�Δ�a��g̾����e҆-��t3�L
bs��)���#�+4.N~,֘����}�~o�'�u�Z�w�a;�u��`ٶ0��������EvK0kh��ړ��_�������$y�s~�	O�}J�������E�X#��{�)��9J�v�}Y{����x���#�h�<,������`��&�u�"mS��w�5�A��ނ��_�����}��& g7�N����h�|�~������5��X�5�A}�}���Jn���@r�̃wͶ[
�'��cA�KH'J�#$'�y��?���q t᮸v⋨2#שE'�g����� �	!��/�|��on�h�����RS��0�#�Re1c�� ǆb�d�+��a0ZipS(��Z���Xk���J�ܙ���
<�^�Ē��|���/զ��)7VIKl�8�K`d��}����
�0ס��&���S>���u *X��cUR�I4�m=�ž���L���v�M�Qta�����aT�q|�����o�z��/�t�E*�Yƍ�����_��nH+(�&)�p��ff�m, �Ӫ9o�ד�[R�G�ە�Jp��2�)��G�	 �B?L��q��T Q���:j?c�}���^?%{5�ɛz~�~6���6+魸��p{�$�3=)���r�zq���}���>���Kc>���}�*p��h`&�B`&����K�ckR_+ik�Y����/�Pm�Jd��u�3ȑ]ۂ���]f��g�S�:]�H�	I�� >K1��G�
NE>\�5t���{�"�ǈZ埉9jP�� �A��^�æ�W���C�%�.��l�f�1�IA����>#D�~�<?��@�X|����4���z����S Y�`Μf���D�>�[�C�RM����TAmhtұ���ܰPy���d�+��7�a'��n��$�'�?��IMkb�KW�V|9�M/um{
��yS�b�y ��K&:F�[үǛ�q�*��R\�[ <	Ťb���R�t:�b�5| >z��Qvf*�#�@m)f;=tH2C�ϤR�1���e���i�����.ˡ��A�(��Y�����2�s������̧t{T1��Gp��G�+y�P����fyQmZ�CƮ_�D@�K�p���o���1@�"�Tg7��,�6Ū�@�J`_g��^''�w9�>1��A�������ne��G_��TAW`����iT���=�r/gz�s�_c^��/�eB�njY�	���u�e��������"�*��
7j����ʉ@Pw���)�Z&clA����#���.)�^��� F˷.?�$�pP�6���n!�H�U��0(T)xy�{��u�W3��W}�6��{��:6�ZKu�En9�_FV`�|Oʌ-��������� ������>��"���?�����DJ`��J�n5N�A��t��q�O�{S�����.���zV7�}����@�Ո�$�\��q O �P��ߚө���t�f��c�����Ѷv���j6[�GP����W��+�kЅ�S;rv�5L�D��鬞�1ZG�^V��ԡR������߾!�hN�EO{6G3�[�3{?6�)���/O��v3;�zd��_V�"(X�/h]b�	Ibv]�u)~TR艜e��a�*B�N��ɱU��(�#Y�S2ӊ��j�F|���b�,n��	��icv�]\Q��c��9�j��U�_��O@�>�fZBWí�J��9;�2۞& P{��GU"������f�ǯL�r��;Ո�0U���=���(|����2����NC~R��^Mqٻ�4]ӕ����T���uv�Nl_V���*<#�`��<�I��Z�p'��&��1�8jX喈��L̯�}U��~����.����0Wv�����X�d���r��L&�k��Cj�����̮}*������ ��ҥ��ݤ ME\M�;�<]��8�L?�.��矧�)���:T ���\��E#��8��Fƹ��ҿm�}�7�I�^0�MBH�{G��6MaVD���|��ʨN��'B�:>�u����mH�����6��:VOn*�Q5��(Q����!;�_JNl殚�[X��i��=JR���)�?!��}�63����`�.�ȷx�FVw���~����C2_*�M����T	���b ��0I�[ew�����k�/��(�&��ĦZ�!��	|O��ٶ�I�M�q�4{ӕ�Tե�#?J�2�haՃ�*f �W�-զ.i��_��7�oǫ��T��TS�ƧQ]�Lr sc��Y��yï�2mY��Ґ��x%[�FVzm��I�ƄK�'J��;��L��'�I
y��p��!�2��#�G�;�͖�J��g�+��´���b��K�0�Q�
\l8Y���2_�:i��͸=+�W�͓���%��t��j�ZNf��bNZ]ҕ�m3��z�Vo9N��2�L��wGH)sf�o�]K0�*�'#�~�7�0D���� �$h{	^�6�;Y�V3��� `��VLF����E�a�W�uV�ٙ*�'{p&H�(�$�戌�M*��w�qѸ�^ ��<٥��3�#�$���D �f�c.�w��Ӯ��\��8�r�<�
Y�� WM�0/ZmdZR�*�����!���� C�M8?|R$�j�XyM:�Mg����꤫��k�|�_}U���� L��i c�5vXe2��!'��3��h�`Od{�ި Yտ[m4�R��E@/��� �`�=7aћ�ڤ����s ��Z������ɥ�\��~��C��X��,�&���	�>�Ͽ�+ǓiUS_�AƗ��P�J@+.T��Ɲ�(���J��Gh@n#f<��6�3�B�:�6Ra���O�|���B1j��.}����H���3�����W�����lr��?wi�1p�2}���:��X���E�w��gl�V8z9.�7��K-p�_�1fJIkУ��z���Ox���G��e3�e[�����LV���Dr@ҫ��;w{�",�ڥb��8%�]�}�[��d m����	Ƃ�z�C��V�����?y�!faO��T$-&s_�]t��^��d���:sp]R�>��^�ҼV#wc���GZ��$���a�2��I��|M�H�[V3�e�X4;�m��@x��7�K�T+�z1˞Xa!|Ll�k_,��x��JÝ��@��T�}���#�4�L*�P�ʩ2u��RQ��t�P>�u�Y�+����3س;��ɹ��I�z e����S�*�h�F�T���%���&��;�a �$Յ�W��mRz���X��)�G�r>)�֨'�Fa↏�����v�.�4gB����*����r�F'��?�#�}��B�G��Q8R`���С�و@;>��/�L�yY�J�~z� @���'5�����O"��[���4�uCЬ/�@�'1a��?*�V ����g:�9�FD"��9}F�4Ա�*g��vsv�ߊB���c��H��6�&�G�j�:?`�	tZ����+�YjMB�;�U4�Ū�>�d����3�7s�`2��=��e_�BP��h����RT.�z�C�)9}1����o����{�9��O8s��g������Zo�����hP�~�sH�k��8�o��	��;h�H�V�7P�ٓ�~r&����=�&�9��|x�Y/D��A���$�/���P�_D��k���@���d��G�KKN����st{d���8��-D杫�I���Z�\�WNWf�usX���\��1���͵F#*�c9�t*h#0@XO�U�Zݳ��#�rط!ӥ ����"��b���?�<a� H�/�g]�L��%?T����3h�b4�ٗμU��>��]�ӷ�߲��0��b��u��?�S�������<`�D|]Z�ArP�[R3�)j�~"R�Pz��T�᯷@*��-�MW�xpj7��� <�Dq@�����˺lk����.(:���azd����8�Lk�%�~"j��:BǦg�۶�7~7L\]�匨���i�]�A\�zh�.<,٦��pN��� �4]"�*z(/>�7C  �6�ܰ�/�Ԣ��C��I1�R����n0�3�;"���}�F������DӜ��~C3�6:�;jv����n�`�� ����q㖎�o��D�7���"{%��PT�&���G��Ќ/Z܎��ɬF����{9����nl�N�||d^�����i�MR'�;�a�#�S)�ߓ]2��ʟ��Ƞ�W��B�7�Q4;Hs�ԐI����R'�4J�Ë��F`#��Z+�Q)�'��B6`��SS���2����Ҵ��� ��r���W���{�H��A`�����V�*W7����s2���EmN�n���B��>��(�5�ay���wc���V�"���%��`��}%���9����5I�����v��_�����y _r�r�؂Cn��>�����@�?�b~df���k�%�D<{�q�D��.��O�5�}e\᠎)�o���q$��p�8>˵~OF:��u�F�v@W��֛��d�oX�b��P�$�7��m��͖����4�#��f�R�G!E���FI:p̙��*Hp&�E�Ċ�J���^'	Qb���C�u�TE���%u�F8�>;�Ye� O�rN���R 6��'W�_�TV>�, y�֙ �kQ�7YGk��r>X�r$Zߚ��P��Ճqӧ�l���\��m�l@|�:}S(�Qc`7��~�Ղ�2��d°{.0l'$^K��1���M���%����"H-=�Ŷ0%^[�< �ޓ �X��9�9�qXΣ<�	�t�W�LT�tح��3x�92f�#�k���6�
��6W۹�p�YCI�뒏d<N�z��������qK����h,�O���C�
sH�g�Σ��� 5�	J�>�j�/�~�A8ډ:�A��������"�p�j�0|�c9\���ΐ��G��@����}��7�������!p��)F��-�Q�+�=�F�+�*��J}�:(�x+I5�ct~��Cmv��7R��/�qg�f�i 69N�:k%���Y�r��]�.:c�)ac�ɬP&����qnjTg뀨��90�xk@t$�P.�K��ې�H2�~�����_y(�\Y��g�z�)#��ǁw�%	'���<�~E�i֓�1��1�Zp�c
6��H,eV�d$����c����Y�[��(��J�#�s[b����:����#53<`�MB9�,jh)�f7*r��
-ך��u��(7F�6ɾR1[�+��= ��]�'����M^��Pph�F�������"p=Fo\�)5}��:�li]�PbO�ގ����q���I=L�JY8��AT+%')��j� ��0f1PU?TCS-"*�����^7g��B�Y�G�5rIt��8�p�,)���H����p$��i�r�xk�_�$=��q���Tz{9���y�~R���\�FW����/G}ż]h8%�&Bq�E���q�v~��p�g1y��$s�IO��J��	��;Ъ�T��#�\������3���k�P ����w��/wd�uo��~��x�r�R��k� �B��z�b��i�(~^�w����i��7�
�F,g`sٟ�b�c9�u�0Hb�U��u�}-���b�LT
��M��
�~N)h�n�o#����V�+�J�Y.�fb�E��&\�3v;�òO�$R~�(��e�'�)n�>��x$��3�_�Y�@ԙ�'	,I:���EkACZ���D0!� o!�#��U��uXc)g�hD��'0�6$�]$������<ReA�����J���I&�;ɭ��6F;e�M�.��[�~���>�sxr�E��a�2�
<-��P�ޠ��P�����q��F�2y�y�%/p~�ʄh��#��n4`��K�gA��q���Rt�R�v��U�1h;���As�8���2Rײ� �Gn=)l%�ʔp��{���!gJ�:�.)sӹ��$'�3a��=Ee?U��j��)D�ud4�C��f�(&c�V�9�d�JJ;/�:J�#V����챓��z��݉�˱���ĚMh�DȨ�Sc`���uwo�3�}hz~`OE.���Sw��"��=9h��"��^l�Ve��/��^�tT�}R� �JǷX���|,��{��Z��d�1t.ao���E�Hz��T淜�H�U��4�x�r%;MZ���[�_h�q~o���" _�Ҕ�� �G���׆�I�(�z�=3�c���}/�>S��r����I$-6�,G�����۾����7e�������c���X�F�8P�Q�Z9� ΊA2|O� ��V�A��K%�s2U!YÓ�j��\�W��N�ç����o�`~�c�dT0�W���'�
��_�o2�����~`���%H�a�K�ވ���j�G�5K���r������ar˪�s���ݣ����t9��3ik_"$��	!gZ�,�,"���v�!=�f2���.�0�v�eS\�7��B��#���T�x��j.t�g�@���ށ\I��vpW�A���dO���pC��ʚ؉l銷��S7T���3�ӝR��]�V;:����c���Z�ᆜ��8f���.��+����ƪ���#1���KJ��5��̏�W�ƽ6]E*�K�ᢴMl�)����@Nr�4	�y�ڛ�AO��лz>v`m)��ʂ��y�Y�Sl����ѰP��i����Q����ﭺdB��(i2�$j���Ml��E!a�O�;ߦ��F��u�䱣Ok�_*/~Ͳ[��� %�^�}����2:�C�=�\���-�b����f%�c��s�: "S�Z���X�`�z�iU�r"=��[�:<$kªa(�M�fʣA&^`�����'B��#pH��O�1�F'}�zy�6�󞤻�=�V
J�T�����#�s�Ɓ��y)!a�s�d��Е��26�3ߤ
����N��{]�6��$����f~���\���H��jyO4�H4&�0po�ۭ()��q����*iM���<GҐ�Y;$��d�@�T��{5��!V�����EIR15����/O���L7��B	�L��<���Ó�?p�U�����_��.T�"�vO�X���3d	4jT��|p��X��?��/�ؒ%�ԟ<�&��B���4�M{h2k�_�zt��J�Qh$Hvu�r}c.ܷ��ȒF"��$Ԅ&ػ����,G_[K6j�����$�@�6h7��P�m�8��}�oy_����Y��.����9V�1  �;���f�Fi��n���{3����_�fE �L�vy|7��_�����ǭ<P�HT͒��R��7T��C0��
�͂�na�|����hڃ*���1Cb���2D����L�㊊��σ⅊������71�s�ˬY"C{�pT���
����W�bn� ���1�"MN���ܽ����w��׊ �^�	�3�h�FXWq����EP* F�?�꺨�\��C�=8���0?����+�w:��x�%T|h�0�� ��Z�����V�N�x�p~	����v�>9z���W����ƞ�Rswl��`��x�TԜ?�2�{��S�͑z��g�+��'�8���۹�0��ra��ܥ����0Қv��Fm�{K��TR\4����nOz`�ל�;�8G�M���r���$@�Jc���>:/�JĚ/ǫ)z�4�m�OM���Ebl	�"^SP~���ڈ�ɐ;@����x^AūjʹA���4s�;RH��a2���F͉ %�t$f���������(�\	�1"�e,�[����l�O����+sY�G gX�3�$��^����š���,
���.G��1ߚTa�R�[�fG[7c�GI�>��+��+�f��$kO�P\f�1��;3�S%n�������qW%���Uw=q�K�4��v7���mS	� ySV:�y��ʴ��h�Rz�snΣg����{'��VOf�H�U"�}� kn��4<�������T��]L�K�7����jK�M����,8S�R��l�g4t=��,E�\�$BM��%�ug9(�*-[#�w��<`����]\y�����ԋ����;��^��8�4Pq�(������זּ�2�f�?-lA�#�%I�k�L=�`�{#R�7 ��`��D[5�JU�j@�JnMg�<�=�Щ,ޥb���o�/��9�j�^���(uiFc�;�`��P.����Y�xl�e�g� R��`�܃O3?�y�{7td���CE����6��cxn�hg�v%�l�c��PO��ky^Wf��u�p���dsi�)�-�,�G���W�v��e��Q �5!t�Ԏmnu�Wo�9��Dm���~��Zҿ�o�h���֌jDN�m~_sC�_�=F�}E�ߎ����=7�z1!B5��"��F�D s�ټ�����*�n��k'�d��ܮ����=��A�i�ɣ�ۿ��o!E�V�ꈖ�l��dԲ��V�1'�9���47$Z�H5���Z�hH���A[v$�!�:p�s*r���TD�$N>ܦ���U��=�C���&�)յ��� q>���p9���%���)��|��q�\�A�G?Uj��B��D���j&�˒��L{w�N�e�=xy���������|~S%<Д��̐α/���:�&���41�m�Xjo�3�A�7`z}���>���������~fJhEd��1d�c�&ؖ��x�O�e�Θg���|�1����,/���3���~�_MmM� ��sh�x	|*�<�b	Q�����g��\�鸏����c3MщG�ȗd���|F�K?&�PA#��n�Wc��Y�r��%��� ��e��Ǥ���ҭ�߽�|]0ť��6��b _�h�Z�mS�"N���^�T*m�ul\[�xo�Gn����Y����1�\�N��0�&�W�������ڌ�����^�	�������[d�Τre��X77���-�Z��j�[�Z��7�i�s�.L�%&��(�@�o�p�+�e�S9&]y��J���;"׌/vM����]^P�f���O����/�6_ nhJ+�؆p�+������2üm�w�FS!'��m&��ߕ-�M�%\=��Y�V|�/}��4M�(�ig(jJ�AU��Ҝ���>�R0���7�OH�hF뵼��O'��f�3Xx�`�m�al��ɦ�	�z�I��S�؛��+e�S$��i�#�E�0њ�oS��+�0�%�A�a�*�E���C�}IA9#dG6�%���������MP�.�,��ʆd%AV�>�2#�쁁X��0A��w����h-���"���5�!�G��;��Ug�J�>�ĽMn!ؒ������E���������M����^i@�F<:��q>���N��@Ev�f\�F��`*�ﭭ�;j����6>�>���z
��Z�^I�r	�M��@��=�~P� 4�/�.Mx�I��n�:�#�w%��V��J)"�l�{ڮN'k]6LI��S��4c�w���eS樃}��N�	=E�%�������L�Q9vL!-�e�9�Ӫ����	�S�{�O?��Е&ݽ�C�Eݷ��9�"W����Q
�5�kCo[__~&HQ=��j��e�
$ޙ�d䔚�m��, ]��/���ӎ@�	� nyP[�mIћ���zm�AN";�q�|;�3\%���Txq��4���[3U�A�����:��m͇8������.Lk2���x���?Ā��X!}1�k�0B���46�5�Tp�F�H�^�B5�ːe{0Zƾb9`�P�W�P3��;���u�09iSj;`� �7}.?Y��l�{��C&��o��@	t_����p3R?����D�&�������L�l�s���5y؄�=���Ƒ���6kFv`ζ*�_f@Jj�l�>����SM��I���:��xŷ��*�$N����D�F�*ena�j��gة��}��,�Hc����$��7`N�+�Yg��
G2u�G�	��+������k��֠
T��}f9G5��Ci}����oZ?�M��[9�����T�� �Ap@u��nr�`��'!:�΀"��M{xm�veqqiI��e��Z"�W��6�Ѝ��>�V��b�
��wYU�B��ʤ��7�=@��Y����P���o�`�\3��$�(*M:�<���*x�Dg]��]���ͼ���$e�J�T�}�Y[e��_�c���7�R��ӭ��g�\�^)o�6��+�{2v �T!�W��tI�c�ژ72��k3�u�g�����8؉���J|CN�����|�,�XTa�3r��t���8P��F[��1 ��O�WVb6p �<�8�/��.Nԝ�&���YӁ�'�.3�
+=���кQTj;'��P3A\Cȣ"�E3��i�^�O��T���۹��褜LmT9*Q�sc���AЕ�����i���J��7
;	vHS��9����*m�^��;�^�m��w:ƽ�Y�N-^� 0@��v��:��K�W� 0=�T>�^����e�)T�<vF����>���n;�����-ǔ�dLA$=���=>/�$+�_t����t^3_�+G_�l53�p{@�o�\�'�قF����7T <��к�I���L��)	x;Uދ���d��
,����8��;d��;Z@���AW��lP��-�m+H)K���(���g��1��V�:8#�Q��%�I��o�׸@Rc�An��6D�e���D纑>vC����L�ݺ:Iy��q�k����SWN��ĮܳQ�[���ի���vhZhj�{`�]Tvڱ"w�oIFșя��U������s���2&s`I�
(�'luqG.��"�z������6�����}�ԪK�S��r���/~��yVA�}���Ĵ�bӑ��6b��ʈw��|����i����wA���^����(:�r�T	�� alW%��7��[�j����G�p��,<�"9Z�����@O.��"Q���:�^�����܌���aCnRL��<��T�2ҭ�N8WJ���_H�H�����\ʵr�ڈQQ��o�Ն���,ڎ`���Ś���	j暇�^�(g�[{q�c��o@Г��Y�2��v�0��'0Ev�!��3���6�W��׵���c7P������?�f�.mxdi�e��3:Nt�i���H��u���;��_EtX��n���&pr\V����h���4��X�N!Ӥߡn���sZs<�a�C$����s��p����o�"�[�pV�XK�2&���,-Z�6�/���'6G������u��0��Դ�1�F���m�6u���𚓷��i��������+r��|��i<(�N Oר�������9�.ڼs6`����b�[U!;߆5���:���M�M
�:Z�1RAI�T�\j���2Jq�?B�WIh;���ǰ,v��m�mq=bq���AC���oL�849)��e3���4��3)��$ɅD,7�ٚzZo���	�]T�+���[��Rc�[�'�j�ίb�Đο�� ��[ݥ�h~^#_;�� ��~�C�x���*��v�R�ly�07;<����OVa���d��ʢۊ��ڶ�-K�y+m�)�a#{^<��R(�]ZKj{��f����.;Tƴ<���� +�N��	�?�O��g!��P��,/g80�od�3�ؠ���kI�*�ǌ�ȭ��C(���ס@���7z�/C��I�Ñ�G�N�/J�/hO�������i*$/��V���3��+�Q��9���ڛ�Cқ �ـ�/��թ^�o��F�/�ޓ�{M�?��`�����c�T�y�Mt�_3��J,8����z�%�Jr�{.>ƽ��4���`�)ҡ��m��ʯ=�� @�w?����I@����4Ng]N�W��2��T�P�Q\l�q�?��Z	��������z������ƀ�N��W^̵�;hfMo��VNb��/e ��Q��a�Uݲy��_K>5W�4�������|�0��=!�D��D7Pُ��v@)�4&ǿ�p��0%�����[���''�8��>��:Ik���=�>�W����@]/|c�@���F*ل����{@2%��N�yW�۝��B싴���Ui������5��R���K����.i���z�(�q]��K���d�}r]s=���}A�Oǔ4�@���\�n,��'`�Zfd�C��;u�ftB�2�����\bX��܀�����X����!����D��f�h��9d�F��8`-c�F�����YB�.ⶆض�(�*q7�[T�<X�Y��-w c��{�ŰS��� /4g�����P.\y�i���2�H�`�BvS�h��}��A�Q�;��r��]�%֎��OSr�J/��"&6�x��UR������b��N/aF�#/�Z��mr:zuVd�}�����ˇ4�[OF�=�a�ڡ{�o��xs�&H���t��Y�c��g���ꖥk��.����q�yq�nIUVZ;�o"�}A�{Ah�w ���K��[��^�{�rB1��Ҏ髀��`&A���������I� /�8|���i�h�!�S��|4X#F�Ō>��O�~���֟�l��/e� ��ɐ�U�/�Ο���D8�t�:E�7��T�JS��l�:�=yLsTMU�H�|�5W��	�k�Y�&Y?!j� (�����F��0�k�m��3Vd~na��d�[�ФW�<Z2�B�@���3'�䄠۫�E��Jt�\�X⺳�Xf74�GOsb�F�K)�4�T$D)�Tqu�U
��-�ub��"����j"r�����.?4�`"y�L�f�\#�9G���+b.�qϮx-�*j>w�0!�C�*�'��-XSX��W^R5Uc, �$g������[w,th���U������7d]}�����-]�%q=-���6��oN�c���P�������������8�e�ܲN��&i�9aY;��L?
qJ��2Lӷ�	�@:|�S��S�?��{�[���-����<j����5�]A�2>2 U��0?��f�N���1�����O�bTdG9u4���>��9�[��vY =��ݯ�_sCAq��z��9�I�o�O��uKܣ�hՅ��b�	)�3�e��2n�7J�_y��ASe��j˨|��G�Z�א>�w�Q%a���q�qf��M8�w�7~�V�xA��{騛uï/�Z�J���z����d��܋L�*��ҌЈ�:�"�m���{ٚ�`:��kX�=�+��/�^����ޏt��c�cF�}Օ,��oA�z��?1g4���[P~@���ê���V�Z��3�����5CE�ДII����<���r��7��kj�CvOiM��(�=�4ETip�P�P3:���=<�=��L)ģ�C�N�	҃$�Fp��_�;��dl�ɰ�?����Σt�8`�Q��c���Ylfx��~�����;�$/iu�y����j`	U��Vж����vvKl笈�B�[�|��.�e�l���Jݙv�4x�,��|+[X�Т��W�O;��nW�Gmb����o��H6��u=��LR2��D�uR�P!��~2+a��;���J�s�֓�Na3�a��1���Z���WT�ڝ�A>��ȴZ��#��S%�D�]�ߙО�ж�����/^u�����#b�Q��Խ��Fzժs��$�*%Ţ�N9k�)ɮ���D�.�U�@������|(n��TpEWw?��{bN��+�
�p>ʗ!���Q	��`���A�r�)�f�+�ϭ�(�����ۧ�eF݉�\�ln�O������TxZ�A��H��#kMm�jr�ݍ�z�2����4��L����Q��zug�:�����aTM~�r�Y8{�t��;e}���ł�������q
W�LB��Dv�=6Z��qn���(� ����8��GRG�B����E�I����l�U�~:��M/йW���1�aIY�'�V�DB�v��8r�4��N�����[�n�0rv30�^������������Ua�oX-��(�:Lڕ�M�G8W^y!��B.��ݓ���-�x���NHVA/�O2Z�])�`U��H8����K��=���H�͘�r�-�����d�~�T�����b���74�wq!�hR�N��y���zQ�6~}< :�C0FS�"����*ܚe���N��Hf����������R�(}��u�֎�1���*m�J�2�X[<����lAc��g��c��_Mو�9����|y��/W��B�NbI�u��Ɩ��d����\���|�Q�4�'�?��b���U�Qw������e��p���fpe���E�͸�C_�,�x��=&��ؖ?b�yt�X1P|̭kA�I>�C]���fxp�0����C>P�O[���>�J��6M��T>go< 2x�G����2ˢ�I�VA�rē߃�����9��tS��݀Y���qE��Z9W�\���o���^�40�.{`a+B��C Fu2)�7�W���\��C�r2�y܏��)��k� m���-��[��ؑg���/[��e�mF�����>2Em��|��� �*�����b��s�����?2���MoHMw,�5���h2Q�O5�U|M���%2���D���M������;t6�OD���C\6��4 ǴXK�G��<��.
`�kw]�����(��2S����<vE%E��}�a�)g�� c�?������ݕ�����\�p)�/��	_ȡ���h��u(Y^��l�qā���!5[C�~
�Rzq�80+�:ވ���6�o�C����3��$`��'�mt�H��B�Wщ��abGG�a˩�؈,���G�c���a���RK�R}���HXи����@���h���CmjI��+Ѯ���y�H�M����:�^��Q�;��&�JF0QmH͉� ȋP�U���N!�6�;c� mh����~���1`d:�F�	���z^�y�T�h3�۱񻰬(|&1r������r�C��°�1��x'@���cPFh��}?����ԫ�ơ3b4R��_S��QqD���B��4L6�&ƙ]�ő�T�k7:��LsTP�'���z�������t�'�'���;�����5���e2>�Ms��`��[V	�Ho�|�c��f�~��!o���C�ɔ(&ǝ�_���?RD:I����9g}pL��0���Lf�^�I�1��)g"�=BB�UY̞9+4�=w����Z�͖S�Ρ�n��O�NP2c0��e�mO�9���ǋ�9��{��R�U�E����P��IE�u�o�+?���/����L2�Cd%���(:��P��Q�am�C���:P��mYk��f�~��
��B�������P��aF���&R	�;�q:�D�h�� v9��%Hx+��@gE&l�������gy�s�P�6��+-)h���g���D�ݗ(B�&���@y�||��I&��o�|T�?X��6�ʜ+��s|���[7��BV�~G�?%w۞�2'�{�Z��%$�f[_��6�2B7e������fy����c5����Q;Դ�IF�qR�p�ΦY���9a3N��\æ{[�0&d��H�/�(v��j�7MJ���!	�Ͳ!�D��_�D�a=>�`$�<�J-��;��W�	l�ќ�^1���*]f#.�+(N��Rf�Xw���a�����NB�u�MIߕ�S��%�2�@��cXZ�-a)�İHJ�Tt��{nW^�+F��*p��O�1!mT.<C�mK�6)Ŝ���Z�%E�{:�$�j��ސկ>6k��9eSi�s_� fXY�3��_���B.�R͙�~vL�	��ǉo�Sl�c�ޔ˸����I0��|#�嚿t�gq�s=8���>�Ce�k�6��+���n��&߳c�]��zy�X��"Hj�\������>�Ў�Ž��bծ T4msD������֖	����W��'In����p�⊟!yU*˅~J:��Y�aD��4��(3��f�$�����;dHL�x��?_:�UE�$�����h �2֩g�͆�_�:����YU���b)�&+YP]�F�|��/%/-��q֪�f���e�B|�'�����듂�3���F7#N�z+�w���Q��ͺ@�l���R���Y�>�9�#�v�ptd�ߊ+�51`o[����2�$���Ӻ��,/��,�!��!�d�gc�OޑP�2Y(^�`�&��}wՒJ�%��e����tig8��[�=���p_6�1;�xS�go�I���8�I��8�FE��K�=�6.~X�^W|^6����� ���b�\]R[&N��Îk"�Ԉ�&V�|�M�ւɦ9�g��<�i&�z�@��7'��዇��j����JG��:Q�o�`�ᑥW:ٳ�)n���չ�,,�zd�,��!��o�1�+�w��׋,2� ��������^U��as��,��b,)6,�ԅ�H���z����i�x	-R�V]J.(��p#�1������Ƙ��E:��˓����)�O�Qq�����2hf�v5��-�v!��f�M|7����T�b^Cl#i��V>�m֠�?:yA�����r�q�^>��Qڨ���IK �ývI���;Vt���dTx҂�$<oz��G?�<�>,A��	��wU������-��By^RNKc�m�V�Bb6u���[��Z�x'k��{��k���oUCǏ5r"Jϲa�
!��;O�����,j?~�$h��)_S_�Y�C8�Xr��p��Z��Ƃ����νTml�f���=l�2��94�'Gǩ=.�8ة�J��#��X�;��e��&fA��z�æ�Ӽ�X��;kǎn�f�#x��3%��ZD�)5�3�7a�p�G���*FAv���P����< �c7�U�m�sE{��ՇS��o����|-V�g���*$-�8ڊRv��9����X�f�����_Zy�ɽ_�5 5����LFu��Tr5o�Բ&��`�>�E�C��B^<mʌ �vW.l�]����+���,�F/�Hte�[:���T����r�nN�y��D�A���z`b����4�������wήO���2T� ���2G�vǉnX���_Ѯ]��B�EȎ͜�D�'RVi����u��O�3YulYM�]ovsM�I�c�JQ�;�?�<�&��Z�g)*e5��Tu0Їv�,�R����
�j^���J�۰��+<�<��I�-n��DΑ�������9���P�9ːE���Q�-h��Ȯ��
�*i�ހޯ����%�� ��F��<.Λk#[�5}�?�oD�&�z	�i4�g'���a�ӗ	�[B�+p�f��VB`~�1�a�P=,�,�m����sH�r��`v)q�-��!C�7��,&i��&���c� O9 ����D'˞�s�cX�y���ȯ�*���,�:����+PM>� {͸C��``2�;*=oV�U3��5(�M�r�߿(hŠ3�����&�(()�����ˑ����3�l&�F;��K��GX��ڜdp�v����@�����3;�DC��׹�O�e�����Ģ�OZwX����.$��5s���� #0���V������H膉fA}���<��_'�I��{�qK�c�k�?�.�x�(���݁�Rșna�F�l��������Y�L�o�FA	�i&g���
b�i����3�6`�s�UA�}f<� J!l������Ꭸ� -��[rx��#�����T�+��!�j����TL��n�&h(0<�v
��ĩ�!��*!��CO���9�D ��B�@1�fs�E�+XP+H(���H$ӤB�@�Ic��^�YZN��쾨��m@��4�mn��)r5�u�e��
G����^�(�$�ZWspk�Q��:���Ƒ�<��A�Ԭ�����羱ֳ�=;�����\^��Z(|�w��^w��3���$a7?�̄�B�����\"��YO+d��n>��żwKd4$4����ã��Q�#���� ����u(N�~x�3��2�|���<޴?�VOx����-?��� h{�%��+X,�T@��_r�G�s���J�=�ކ�#J 	2���8~��?�ݖl�Il/E��9׍:�]*x��������i����������V�sZGM0[�Y�6 ��k��qTvUa�T�0�zh� ��_�5L����~q/lX�C�$�����(w'ؖ=�3�9�f�[^�xo��4*��{"�e1��9YQ��Om̃�Hc��;�?�����/Wѐ��i���eJ#���:�d	Yyb�>a�Jh���3R�z��Q�m�a���)H~�r�J̳�����9�x;*��q�S�v~��-g~z]��U��nd$B��C���D�~�6��|�ߍE�5�-���d!��������6���.��L�O겓��q��B��iE\KO;�sŬf�pJa�X� ��ysؔ�F���;�������V[�������a)�1_��o{|H�S��5�)M$��"�2���B�=В;x��w�q	U�2X�mN�S�_�W�'����ׅvj���R����4���{~ �'&�Ōrj�v�!��	�Mo�*��NuRl�4\kk�7�s�
Q�>jR�J�8���=��(JZ�EF^��e��"Lk���EPg�1�seC�;߀*a6,Qjj�9w]���$� �F�HG.���6G��X8{FԞ���J��TI��F��e�{(���btj"�
-�q�Mp,�z-?��[����*,q��R��͂�d~������L��O,�]�)$SM:�m�yt��H��l�r����b�[l:�k�.R�i��δW�Ļ?�l����W7�"uI�����w�E_rd�NEy!|�̫ ҒKȓ.�p�s~q�#�YF�̶8ܴ�_�gQF��?�V��g[��}S��С��kTP��TT�d��d�[�Ի-Y�_L�H�LC�IQ��|f���	����$Vu���r�c]�wLa�ݒz����O�}-꺙�a$��2�˴f�Y�/�&�� 9M.|��yl`|
R��P��	�S���.6��$�W=n��"��LB0�<^���و���<�A��ެ�I�}��������	����՝�y�ҾJu{R�yUw����S�Ǩ�O�e�q�����^��CY��� �YW��+|E��LH��ϟ�l�[��xO�]ޜ�P�Fz��Y����ᾍ��i�n�/w��<nr>��n��9gL��,?�D6<	�#�7w� �������>����^�����l[m��e�$��1{�V5�ԛ��~�ɷ��)+�{�1�W;���L�exB��PX˘��z�/T�!��ǈ�-�V�OO}K���ъ����9���lPO�6�ZQ�,�w@�g��@tY��u����Tib�{���XMQ
��RZ.X�V�!�7�����'�){��% T񥐗�l�˃ ��#Ɗ6��Q���{-��X|����s����������7w��Ac�L������ɲ������63�ᷧ�틮x����T�:vR��{�l���||�I�r��� �^�;�S{@)�':���PPso�[�A����Z)�z?Q���'ZI]6�2Ȇ�nr����S!U�oR�	A��6ηx�F�>��<�	4f�iቁ֞��g�B�&�Z�Q�z����!a�z���Cd���M���n�+�����;�9t�$�=:�0�E��ù�8G��m5�sqYs��-�p!�v ˨#�!�9*��%dH���n�g$	���dv��{��H�K�b�X@t��Z���l�e坙���<����K�[J�4e�G)�������Cd_�ƞVۯ5���㚋Wqg"��Eb���K�J�/�n���Ր��([���$oc��р��1��;(~U�Z�ۺ�%O��^�G{��2��A��kR�
a>���-�\���qr�l�`���X�E�g���GL�R�Y�V���7 ]2&'�s�M�[Q�mY%@f���[7w̠���X�,����������A)�{��<�����.I-P�P�����=�b� oF���q���S'.9�-�
���Ë�V��h��w�%0򿕟U�ro����P�W%����S��Xm𭥹'�h�W��Q���L(����{��vy6���nz���X�&�lS����Y��T�P���.2�??n�R`!���n�� ��H�bi���L�%$���"#-|(S7:w�>�ag��#&P2^�j��>vS��1@��E���0�x�)��h�jDў�
�c�g-`�tU��T�6�tA�g�ĢםP+|�)���U9� �2�����<eU����rWŎ��g�'v�w��G%d��!@��D�����|��ӡ60�`�iFN���Ƭ^��r�F�����z07�Gѡ�2�U��t��G�6��5�`?&9���&��S.σƮ��`�Գˀ�Ds.�C��[���Z���B�L.�V��?��� h�C)3�����;�;����/{�s�3e���Y!���7O
��@�@��KA��
_�7�./�z+�l��]}��o$d
h�Ji�V�l������5���&�7>@�࿅y@	��fݠڰ���Ou/v�,+�V���]^~�J㴯�R9�ڹ�7����QJ�6�^?��e�%(y���H�)4�����Ģ�4I}�~���MBm|ut���1 �y�`�xq#	�fuV�ZD�����%��_���K�k#5�@��uuM&V^!@R��o?sat���{�J�ۭ'aE�������}����c�Zǚ��r<�w����������he�l'�����3�uj�z[,��G�"�L��H��&�Pv>��❁|v���*�,]��(99�u��qT�z����?C>L-ڟ8Y�8��]�A�_W�;&d���� E�ny�(G�+8h\�4Ns�|�lI\bd�=��'�
�P�x�^ů'���zwp��>� �?��-�>��!����}��"ѫ)�谴������U�(��Q�/JF,߰3h��B
> �R$�x,�n�d�j��_�i-�P��*w_��� ��ce"��^����L(H&��8v�rC�w��0������|KZݯ�wg;Tc_ۯO�?I6Fc�l"\3�-=qg�#u��B܆*�c�L���w?�ov���M�,G� .�9�<%[���|���l���Va70�ʮx1^-�֔��w�~l���h�~p�c\��m9�GUv�X���]m+�N{m����M �K�S�bkO�����D�hc�+ѹ<�:F}x�~��`�}Yݝ	g6��D�7�T�����2���	l.�w�I#�������ޔ�G��Ȏp����[�x6t��D�.�W�VMM�|��U?J�$��KP����`xu\o,���g��dD u1����&[����?챶����Z@�p�����L�f˾
+�So{�?���1i#X3ڼ�r���]�5_t��>��,x���h���+bRYn>e	�nZ������VU�6m��Ҹ(��K/�I�HZ�4~�b��qM�,	N����	�qA-R�:�)�>���$��]r������U�S`�@ga���Յc���c�[����jq8-S�tH�*x�=Ss^S���3���;�-_�w�f���y�ȳ�i+N�z�+$C���A��D� �a���{�_%�^h` dy&I���%_��TL㮊�8�$Ǟp1+0Q+��W��`�T���+��b��n����7��K�^9�xwΤ݀ ���t��B��b�ol��or�ԝ���U��f�(��N}w�t8�|�ʁ��+���a�^�Tg*��y)0w`�wm+@�k}�����e��G�<�� �J�v�d��=}���ġ����c��C��Xr�p$Ӆh:�"�L�*VH���p׬���J\ː������Z��s�/��V�J�-�~��e�hA�l���k��q����1�B�9��aq�v:���c�VU(#dnO:��Y^�hRv�jo�8Ս[`�N�
�� j�aV�u6����Z�w��ϱr��sW0ǨRL�
 �U�oQXςtN؂�e��:J��Q�Z������[���x�^��$��J�_�ӴØ�v��e�[�^��~l�f[��'���H�3�[�]B��z[C�F8ڱ2`=C����=���]���Jp��K��l�.d�D�@�\Vn�+��K.I*l���vX�"�N��)fJo�V�Q��KF�|�E�>��� ���n~�$�j-�%���_6�T�)s��۩3q<��pP��	~N$lw'���;��L����pw=A؅Y�)�Mه#�<��b4�

u4#�����C�4Rw�	X� ��U��6͊��t�� ���*��@����^�g
��կ�����2��(W���:9���U�09�Ŀ�������C`��sn.�m���8j��g�M���B���<�VD�s���"���dHJtԛǏ������c~8��+}社�U��B�B���Ie�5�*�؜$I���V�uo�0�0�L����g����t�g���
©�g�K�9��W_,�[.����(sO1��,?�
�'�H7ْ୵*y��&�6`�H|.�w����%��q�g����g��΃A·ۘ�wOQ
4>�*i���>���]0fG�ؽ:�2���������%�z�i���CE����9�x��%�۪h��g�V��Ҕ�ϔ�}���
f���,��	42?�����|����2����1������)���+1�pS}�{��1���4�{v�.C�����-��[-����5�6�w���G��cn�
핲�f8�=�̶�71-|Gĕ��F��Y_w�0/��@�/�p�^�N2�wm�^�����?�̴�-|AТP��b��*C�
�~�w {�!�}��ފ�C=���zx�}��{uI�F�>sn����ǡf����2��U�����\��t
���0򝥑�Zo����2C�v�B�FJ隱IO`V�$���D�W����η)2�����y���*w�ѵM���*�������~�����Lㄍ��%��Mz�������/�u-��c�dm�IAb�8������$�?kZ ���ަL�g����z���m�C�:�)w�<00���&����&��g�ǝk6pg2���왛�mh̽ͽ m���p���W�;m�orD�J�_�R���1��ib��ug�{5Y���	��6�����qtlͭq��iLW���<!so�Fw���n�]��[k�W7g�[�ҟȘnG��p���/��W���,Vڞ��_|ܧN_�!�����v�|�;��!ϖJ�#������ƀ'j��|d=m���ﮱk��X#�.�ϙ�K1OL*BX�td���)$2��7�y�pn\ƕ��}^�6�_��ǭ� 'j�5y(���g�t�ղJۣu��ۊ�}��p���`�*Z��F>*�}����o�2 ���}���k�$7d��n�v�N�(��,����^\���m/�!7���fi$ ���
�$�b8�	�<�[Z�7�\���S�Lm\I΀,�$yy�g�/�����V��1.�\�@ Q�nE-��fi�6ʻ��R�Q��F�¯,�C!NO�0y����q,@\�H�MQ+���p�®	��9e��������%eȖ�8e�Z)�A�o�-���2K���L���geYՇm"��;U�Hj�W�0���d���Kˢ!��;�6#��.���0p�*�B��8�/'�i2��x��U��˗k��1�A=��y
t;�Ң���6|�S�'���0aG�I�q�f���p�S9
�N{달=���u�Q���'�z�a�w���/�̀<K� ��K���be�y�K+�{�4���s�	�m�%�*=�
�A�5��T��#�F-tEލ��%�Կ�-������i�-�w�5,�IMF|!��0��^Wiwf~�8�`�I�k{�ۻp��EdJ�������[�ܟ*��s��N6�p/�� ���
�<p�����V�ܬ}ȅ�J�d��#��f'�	���1��ua�T����g�pa�>h@*LTU�ʅR�m�Y �k�/Z��[�CbåQd�6\	ī�(��Lp�`I�eݢb�M�Ȍ|�y���)Y��]�G��X郏��ⱈ�E.�6H�b����L���ь�;����qxE�P��@� ��}�+�
��h�-U�J�!2�*Aj��T��0_G�[�z�+n�����K ���5x�1C봔�f����f
�J�Οnϲ����!�.4/yy�up�<�L`�c%BXk��a�5/�]��{'}��Z�H��A�ҍ,�IpCS��"_0@���Zq���m�#�-Zw40$/K�L`�Q40�K�wD�~X�F*�(�ξ�i�-i[&��I��e#�S��rT}T8�&�\�����,�zˬQ�Ok\������N�3t�;h���^S�����f@4�E�Op���T�S@�:�95��}M�u�Y2ݥRۜ��ǩ�ъ���&����_zs������]������B!�8eX�c5Y���Y�����%�b�[Rr��)�^��5����Օ"��t/���.�d~���X�V-��"F򲭷��d��q���԰��5�3�tp���Tq_L`���W�O��y2�����tRka�U7���˙t�d�}�Z�r���։�ҹ ��yO��䚆�_=�^<�ci��]%���J���DcT����.��kU�O���ݥ>K=���G���?������] ]<r�2\#�W��M.&�9{��ڸ��a_�Cijqװ�̴t�
�l%���)�ɵ`Q}s�8�:E���e]�&�N�q�}�f�}�5d�/#�fi�+J"�c����#,�VF����"�@��1�:��Ÿ`yB�@M�lF
L�͒���+�v �/��	�Z� �Mx���ہ��Q�(�1tZ=���w�ɂ<�D.T+�&쫊e?�K�r�[�__Q�u��� �1�i#\}�����~��B.�T@��{�o��ע�r�栬X)�����w���ك��rӞs�#�Ō�}���"U�`����6�����G
��k3ağ�`��D[���7Z|o#$�b�S,H4����T`r���đ5~�0�id��ӚG:����x���

jW{�g:�ɩI���䭷�E�ek ��k��Jx�-R���
�C�'�W��	������ F�c���i6����6����9���=8?�Ų>��� ���ݴG�pt��-	^�$鐾��5p9���f��v�_877l��ߛ��U,�Q�*��;����Z���Zi�@iR�.T9sΞR�]�t��Y+�J)|�9f�O���Zq`i�n�4t���e��  `9¸�,�\5Գy��'�_��g�?��yO�_BB#��������PhΎzo-����
a�դ�y�}Am+�2L\5�\�2��?��]����%�qgX24��^k,�W�?��!�VJ0�s!�ff�U�%����]�Y�Կ�Y  ��<��I|��Az���5�IN�c��i0���U���0;܍"�f���K���
%X������{&��24�D &qvMY�uf��n�Bp���&�h�v�\h��#c�ز� �Q�+������¡����[�Y�ĜD<yӝ�g�^W~����)d�{<p~ۀiY ^.1Q]����-4�jZ�?��<���� X*ݡ�j�o�c�@Jp(i5����_�d�R�{��t�5���п��M`jɑ'�`��i�C�G�x�?�TV?�-��w:C�ܭ�h�4��^����1�6���9;%��QB+��I�V��W2�!e��M�D��g��r�T�X��G�[��רع
U��o����>����]B�MP8r����@Е~\�r {k�>��=���-�b_ ���]@ƹ:K3ѻ�'G�'!+�hH�ht��}0o�"�ă�X�m��	��V��6L���@+���週�9���lF�bG|��Ij.vK�0�{;�ҺtO�h7] ��)c���f@�e�����C�&:H��z͎uJ'��ԓ=�^��Ջ�3w)7���,��b^�����p�i�'��U����┎g��4!ԫ�H�1�{�+kg���3�j�CZs��3�S(Q[��('�̕���O0�Ӧ���D�� _ÿa�� 6p�k��P��A�Y���z����U�k�T�M!���56�w��h�����RT��6n����q���kl��l��ծ_�����x8�}ŷ&-1{m0�9�c�l�Pwѽ�g��t�6�-{��?�c'
WPF�Nt�V��,!����)F>��0��NF[�ݪ���l!��o���-zg��^�G	j��#�P��]���ꏓk�����%˛����UM��d3o4���q���]鬛��\B�騡�h�VXU�Щ�7I��������uZ!�}�9N5�;կ��sT+"m�_�L�ɳ�t�����\$���z��ІeY�ǻ|�c�^�X��7��絅�g�PyN|�����^��G���b�ƿV(�zP}� ZA���X���#x�nD���H'sR����3�9@��L=��G/�Ό��(��?%]����z��4�5z�q<�C�
���9Q�=����*�����1mf�m��
U>����������TD�^,��`ŅRRj���s\D���d��j2È^%jo���9�Za�ɻ�� 7\H�eԵo�� ,�Qǔ��N��4��{}@>�'hTr�{j���0=x�2	ޛ��2��ëH�h�Lu�0��@Qc���jcTڅ�Nn�΍�%y6��bHv9�B�Eܶ��0������.��-.Ծ�]($iutbU�]�}q�D�r�z�B����z*��Kh�d���*��]r�^��� ���g�����=�UQ����	H��QlF��lE�����L��y��Rr ��n��\;�����������SJ檵{�e�3�˖(��MUƥ|��e¼r�u,�6Y|���H`24Q-�o��yu�DC�F�~ov�:j��D��i�Obˇ���ݙȂ����fS�+��K��^��ɉ��6ob�����6Y�d���<�a��r��+��u��n�hwԍV���7��B��ܮKr���^Cl��b-K���?)���Pn��������Sb�$���XN_v��<�ѦO����Iv�����!�[={��� �����S�5JR��vq�e�fF�qV)�����ZB��W��j\��9C���+�� t2l�11Aa"?���k9�t��׆����=�[�h�4ԖTM_����5� Ӄ��>L�a�� �>�~���vh;Z֞��G*�*z<�
B�6`P��AIsߦ��B�ڂ��n*)=uq[�]��OQӭr��
�hw?0,�L��`�~X�bj���>��/������|�N.Y=i@\ M�<��fRY�a��/�� �͂\+u��o����܀�&ߑN�)i��:`П1����\v�-�U��DN�����8X��Ț�kPe+/9j�gآ@����X��p�>�]�2,Q@f\t�ݳb��V-�[���jt�ɛ"�(rQҥx|�A#Rs���q��3��>Bct�y�k����*>��F��b�~As3�H��i�?"J��k����4�	�>@��Ě�%�!¨�}�7�X�\��
{��h��{{L�=3,+_���C�2b���d�5�զSM]u*�(��r)[:�Z^
���S�h�xu��.���/�ɻ��<�c<K<�c.EA����y����@I�j�}�v��W�D��#�����~���9�8���'�'M/����vZ�֬4����#\�_"q��#j���L��Td4 �b����
L5^��Ԓ��|��W�2���"Qjׂd!��3Y�4*p��+���:,"{^���p�O�p �͌�f8���x��*����i��BG\A�:�����D�e�ec@�j0���1V5�(`��2�l� �I��PT�����Ǆs��r��8������'M��Z ��(z�t|Bqu���K�O�IX���n+��(2"ӕ%C΂e�Y��f����H:�O��iϠ�6��"��?�xU�Xꀦ��vmq�?_^�-aR������GLx	��.�eQ�����<�c��E�jν��/��'����a�ܓ���?C��o��o�ߑLk�9'\�����i�X�ku�ƽ�Ѻ�9S�wg��ծ���\wT�-o��z)hߗ�?0��-X��e-�+�4\؊<�W^�S5f�?Vlφ})���ׄP���Sp����pf.���Y)Lo�5&��;�����i�1�z쾭y����s�Q�Vk�"�0�b1���sf�����F����3�����f���g,����U22�%��8����nl�;Ⱦ@���Ʃ�����xS0�u��oE���h�v�F?*IL�9Z{t �.�\�À��O����ߖɰ���?���q��0'2�O�Wp,V	g�|�O�h��m��?P�CU�)��sܢi&��+���݆%��O칵f��k!Y���q��)��!7�:���#�{:>��RH��TR�O�Nhl%Q�;֞Z5i�fW��}�Кo�ܿ'E�=<�֪�$��Q�����;�`�fpv�����C3��IY@��? +-}S�l� �3��	�ݚXf�J�<�rhY���E'J��������M�W�|����p�SD� �}&�Uo��%��0(�SѼd���/'�1M'��E���>!���R����4_'���H�X��>���Fs��n�P�/v��_2�j���	�j8�42{���	q
H�	o ��swZ�������~����(r�$����B�C_��X���r ���P�G6�G�`�PE���gw�Q�T���_�ޮ?����1q|3��������I��>���ԉ\Zi�Ѱ@B{>�qV�.�[̜��ԏ␊I�[�~ݏ�& � �=�J� "�"ü�v�(�}o%D�1�����M#f��.�9��_лQ�|W�k\��u�-��jº[���%��Oe�3F���ٱ�p;I��g`Гٶc�mы{�����z��3�P`�E1�L{����5Jȹ|[1��-\*��fC?�����0)fv�үZn��E�$*Y,��c>E��Б��ԦD-H}q{��ʫ䗘v�k�!�������qn���Y�/�Ӡ�3�P�ύ��!	�x�sf��S\�WYLmʻ5��%��k�'�y@6j#�#���2XW_t�Mj����QB�G��^�>n� H�~�\O��&��A%I����Qj�r_u�_�n��/�0��.dr0���?ۥAO�Pq�2?G�vA�M�#q��N&����C��-��ߙzƩ]�<�`��}	i��46%��Y���yp��:A��&��Vώ�{r�����x�����~�󝂠HX^��c�`����@����ނ����7R� P|崫�5�	ܰ�/Ӑ���d�I 
���n�I�kӅ��1%����ۏ�{�l����2��q�;c���b�4 c1L���4�%Te_�UQ�z��g�F=�Cd)}(������Ə�m��lgn	�>��y����D�E��6���z�X��=�.n�ގ�����f��y1F�>*mtB6�Qa@:��:D5M&��-�{m�6Q�ߚ� ]���U����$�a�e�Y�P�Y.z����_��ن�\�ibD;��Wrm�J��W����|%v{]?@l�aѱBě?���ךM���7��\����h9,��s�è�>����v�����^�	�]Ó��ϾJk���EK�U�o>���5�3A�!9��y�����*�4�l�0�nz�}���v�V�N$$��x7h$"u~�h����E<�ځ#4#K^�Y0+�}�Ӯ�g�RV|�>x����3�X˷R�N$q08%�B�+�D�eBB�0�7��	;冔��e@��>oi����;���M�2���q�D1�Z쌲���o�V*~�-K���D����k$�n=�yI���ǂ�+W�k���(��Ji��S/iݗ�Q��Vx�S�V��a��1M%;�&��,���u��=�<�M#����B}-�A��pr[k�z{���@������B������.
9����木ݰ��E!�+I�U6�J�"m�����S58�+�����Z��h�Չ��U�4��Vi�cYQ}�?�ܦ|f̉o�v#�i¿���k7����ն�L{�,��w/�Z��G�O���>ln�q���K���:	�����g _@�x�B��T�
ʱf|BIs�}�kƫx[r�°���^>�M��'*PnEsa�S-�b����a捣�`��t�=�?,�Ƥr�.�L�\�/㾄\�bw���!^%�U��I���L������M9��x�Q�����[�,x�w7}�DԷ�)~�ɷUrqs"�ё�P:F��NM5�1�X��V�P�Pt�8vbT��k�Ч���~k�RZ���z�5Hp�x�K`,W1j��te������E�Fu
��RF+��U��%��ی8'��*� VF�Fן���b@Lb���Ԩk��F�"E�>�c���P8�Y��R;b�&�r��(�\(}��䷿������UyM\*�
�31M[������>C9I��w�	+��WIQ��a\gI;!����� ņ�r�As括 1�G�Jnz<)��gD�u�|�չQ�*����I�f��L�nu��-��=����w
 �E�vף}��6$�TBp�M��;���Z`�ֈX2��d\��}�5���h:�i鹣ʁ��ޓ�uuIϟ�aݞ;�!������dI��ԅf��p@A��-[��>�o����1�F������ <l��1cЉ�\R�+PS���Pm{���@j2,��zJ�4~5�6�"���)�7rfE��g�O�za���AK���>��}Q�#��* ��HJ�"=��,�w�'�-����#�܎��؄�Zy ���?��2��Z�w��*��gE%����W`�d�K I��r�jڞ*��aI���'�췊��p�5���19�:�-�_�(��˟��O��1�a����5	��?�U�a*􀈽�R�_�a�J$	��P7�v��Q5	��)��񯪄�6,�ħ+��Fh9��xEE���g�sQ�����N��Č��B��QC^_�a�4��r��g�X)�YV��S"��#�ҙ���ա�ᡵ�B�`H��:�o��z[�;���ܘ��-kO��>㜡�6g�LA�h(t):ރ����ށ	�.]�+�ˇ�͝����� ��)��n��ciOs�*2'��dS �W@�C�{A���;�p6�o�f̅~�~}�[[�h[O�}Y%�o�zg�US�~�_�y����`q/��Y��}ΐ�𣙒�5!2�^�����G�,,S��CVM�#6�G��Z�)��#�A�zR�o�_�K"�lɧ1�\��,��[4O�fY��*��2��m�:O�6b=7ӣ k�|�T�V�:����A8Ђx��� ��k�qY�QM�S��5�w�@/���z�@�P�*󯰉�����v��۽����g���}��6��@����"e���J]�|��ƉHl��2gK�SH`�-�g�2d6c��Tz/d�9��z���,�����f���=<�BC�{�-tSaG#�R�A��5%��ӻwe=�g���f��RMG�c�j���_��@K�aj�T=rc���]�"US7*�*�W�7����6���=�o`�xY��2kuvl��`ݽ�4�,Y9�K F���
벣a��
�!@��1p���k(��s��Y�&�d�?>�QK��H]�-N�k�$P����*�4����D�����F��ocf�A,���?ݪ�LH�~��4J^�����x6���GB�!���.
�NٽٴO%usE��S�Q}fj���l���	���U�ZT�
�T���t����� ��AF���D���d�� lm!M��f���hY�օ�x֕��u+�ڥ@��[8Xa�^�) Q+����ވ֥[52�jAm���~q]M��~��2���������n�2tU\!G����� ��a����0��� ��o��X.��*��qbpS����=b����X�++U�2C���-n��n͸tx�ĭ��QWPit���^���-��?����ېol����Cjn�~�*>hPB2�\��x��W��Ÿ����$���6�>�94W�ًɚ�AֳX��O�[��� 3@ױ@�8�@Iکؽ�CB)y�*|�o��j߼Q�"u��a�r����<s��p3����5O����R@0������{���*huA��� U��N?7A��_sM$��}%p|	`Ҭ�-��vo��.��!
b��Qn�r}���t�-�m�����ڳ˽�M�����&VvY1zF>ڏ��4��z����SK�5���E���>�F��[ɞy��d�:�Q~
{��]�9�	Zy煮�q�U�	��{ɵȶ����d�(&�u/�����b^��,���2?Ls!��8# �Q>h_�<��'��޶x��u��Թa�W���X�#�����j����U5�a�����_��"k:nJ��7>�%�>��Q�"�섻���i�h-;O�W���b]�
���L,�i�̬�]ꈙ�"�鈢m�?���R0vzz�3��'[㞃>�N~�ǟ�N*���u�����U�m]�R�.u��:i�<rƤ�4�3�tQz߈yu�|$eg����C��%f�Nb�z��5�o�|=�4�Od7������S0e=��=
��TZi#E�z�Q6~;���a�6����TCR9Z���$h+:p����;�l����#?�s����,��2ė�%�B�H$�[�����T�A�u$b����i�S�W��T��S
�������;3�.�c8/:EЁ��:��nO�͓�a�s�襈�^.�x�ǽN� 4�8�~A\c\ޑ�?�����N�gu�n-�@[�|��Q�	�d��:N��A
�3��v�8e�[o�I$�Xa+'	��py�kBU�����?>A�1�Ym�@i|!��h�������m>)�=�6�]�L�[$�
'[4��y��9G����-� C���"�A��݋�8�Չq��t1k6�w��	�����.�vp;��3-�k���A۾��
]GKN� FR����u�;uQ���n�%h��ԋ0��y��@t��Vyh��
��Ν�d+�r�I��b�������h���3�ê���Ә:� ;���л0��,���'��C�r�� �M��k0;a˧�]������$-&� ��&�OY<I��e���� *�m\��\'	�C��1$�8b�Y;C١g�(�S�^an
iV�Lݵ��@l��n3�?�߷E7E���07��q�U��8Zs�|���P�^��� K�d kّ���H$��uE�ѱ쑢X�z�'�)X�	S�b�+n35�7]��1�~�7�������� ��&.h)s���8�_%�DR�nE����A��Ll
R\[��b�.ꂆ��ˡ���?|�y��p[��[1�S7,2k1����'b�I���H�����#2Y��z�{ر���5����Ll�0�����!���[��Q�gO6�yt{��!I힯ܑ�!`���1 ���Ƚ�'?-�ҟ[���i${q�a΀4�y��'�>�LV(��K'ds�B�y#w������j67mCU1�����ڙ���"��_��hT�}w*�f�lZ��W:`����1G3�F�{����\����߾]D/�����M\w�Nڍ6��]%���"'ś<�?�%�}��z>�V��x6�A���Z�E���+�;���M��J5��%�+z��YbZ� �ė��ت+���A��*/Y}������4@�H��-᧾�)8�h�
��+�^? ������ OQ�e�r�s��'j�q����^E)��{O�!����m_R]�+�I���B~:z;V	R 