��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i��͌c�iv����'ό1_��A�����G���H��8���ř��wJ�S��U���A�,�{��k��2�Og�L�@�_=�s�d8�7?:�&�ȁ�꧕��׉�F�d���	\�J	�q/|U��Kt�'���%l)���~��M�	4��ٗ����ɸK���g˟h;&ύd��G��H.[E��THg��e��ʢ奷]�_��/�ː��)�d�ܣ�`���̔�צS���N#����E����)������y��X���w&0�&Y���7�j��Kݹ};i"���V?ƃ!n����N��I���E۷��`LtŢ�\�S��`����Zc���<N���<nq��t�,kX��_��#�"ǲ�z��$:yj����ra�9�Bu�b��
Q޲�tgN�9�2���7%��o�WO�\q�+2d�_���r�z�rW08$�k��C*�ق��m�]Ğ� n�ܺ�ش�D�(�_�ɏ~��P���7��i�L� �\��nu+��,X.��2e�=�!����/�RC�d��{e�`C��s`��O���>�7�>�|��}�����k�'
G�/Jy�����Ҟ��X�x�f}"�a��*uE_[�F��1�`� [ 6� ����dM!W���.��� �5���JLq4�=�;����Źj�&?%�%U��\�1 "��
Pz�ܫ�U��=޹&�[*ͯ��
l�Ӵ�Fv�)�D?�&�0��%g�۹������v��}	jj���S�f[ȟ�=X��V.��]�`���Ty,4\sqw&�)zlH��X�--3/��7� �D$\�֬68�,��[����m��!�	I���  �vr����H��M���w�H뛰���i���l�ѵ�	G��z��|Gp*�5�L�|�v�6u�[�u�p�խ��BQl?�2ܗ_"�ֻe�Wz�I��y�!pw{��pC��se�W��,��hJ��/�_%��_p;jߗ'���V�tyc��X�8'�jY��C]�=>	��q��%�W��n�ߘ�pW�?8�5ъIߜ������=��FϗL��ްc!q8P��枅-n3^k�`~K�.+X�S~)	aM�L\+�c*м�D_�ʕA�d<�&�g��G��''�m��ĉ�w �D,_��<x+?�fn��L��W�O�i�B}��#�{Y0�v��y�B��a�3�`n��_3�gt=��T�T�������>u�������=K_����Ņ�FW�����:\�g��MC4�o�{M�τ�[;e�C\� 1�R����*T�����|��s�?���^k��������TQcHy���E�e���%~8h��҉?��3�('8h��F���d��e��p|[�3�<�c۟o�[����EO�d."�Y"��[�*����R�����N�����+!���8��(o�j�B\7u�0kP7!ݤ�vN悋q��U��� ډ�&ǛD�065��y-qt�R�E��}Q�6���0b;��R�C��* ,��I}I%�ϵ���V�ka���xtP�{}W���3��e+�۸B��O�}~%Yʫ��m�Ws
2Ɛ�D�?�X6�X��Ql+�-1N���p[��,��>�W�����c q�z:�S�,[�9��Ayv.����/~�
���:]#�)����2wA�G,η\��PD-w̝��ɳ���L�߻x���t���l'�ۈ��}�S���a��!��a�k�)!�E
���5d`��A\�ݿֳt��pK���LB�`���$��!���-��m����-g�Z��X��T�.aF�U<���`���7�f�?R�H�/^2cE��ʧ�d�$!�8���|�A�O���X�����Z 4�^~YcݕY�����VI鹹���uI^����lL!
|׊Ll�*{bQ�ʎ	���ҽ�v�h'{r��EV��u���gč1����4�!뻞� �Q!�=?�-�/(C:l����%�������i�X/-A�>���U�Ȓ|��{�L��\�G�)ahmw�����p"���2���DtAmJ�w��|��Z�q�C��Q�F+�n2~P���؍�����QYi$ m�8��P���E� �(���g*E�K{�{p�7�8y�$O���ᆘh��/"f�	,7�)���U��F>�Z�`&�D�LU��R�_A`�Ԛ+��OSr��r��|���^`�F��t~�P&��	����R_5�:�+���S|���X/+�r��B:��	�_�2o����'�]a�೺���f�}�`6z �#��5ƦC1	U �{�Ԛcö�����M��aб!&�⣉�>#>\@��.�}��ȼ�q�"����1�t:�:�,�O��x$`������i�,�akN��#�?�̺�ȡ�-JD̑��d4���qY:ܖ�>1�S�v͊Bÿ��^+Q�� �5D��nT��ϱ����Ŵ�>��c��]�Y�����n�Q7M�������,<�4%	���l��4���=�v ��'5�LTm�D%ٿ��C��+Zl5�"�.��:��&d2���n�fb��K�ķ���oZr�^N"Eإ�Q%ts�&}��*U�-�N�k?��"ɦ+�,����q��Dw]��P�}Y�6�Oi���+��I���LQ�C�P>\��
�E�>��GTɌ����3����-�~ĺ�?�5���#G�rt��m�d����I/mw� k��%���=�-ถ+0(>�)��c�lM,�Y0�z3�(��d%�eќ�
�����H�����j+~uC̀e?���э#󑗯�1���)�X�?.r�m4�Ͷ��wq�c��eI�9���1��WȾ�NOA$��Զ6P*S����_�;?WSڣ)�������	�.�]k'V�eY��~t�"��?���eU�� ���	4�nz�Y�L�GG�G\�f��7ƹpKw~FC�
�	Mͺ�9e�9���ϵj]�-<i�Q7���)��>w�d��cߓ(�=n��3�S�D�SΞ�X�&ȅկy�T�nE�r��	x�2i�O�n�~7˸�*m��O��w�^��7��P"X~��8&�Hd��!?6����S�G� �v���W����tۄ)Y��[�G�q=	!5�9a����@�};�S��g���g~o�������K*�%�(������E��,Q���]�Р"�����%��f>���1�7�����t<�]@�=�`�J�h���߯�`1���IǇx�A^-�F����_&���vE.�!�k�{SMp9�����@ьm 2�O]�pPRha��"k
��աvЗ��5�[fu��