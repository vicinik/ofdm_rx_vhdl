-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MWKaoTj22VTgGXqfHxjiEQIclw1FqIWTuHEIad+PZE2Oco7ghg697Lez5wC2FHZnxrnwP7Ygf9nU
RNsuBIBb5VPaRCeQ0sAPLThnXGVRqIys+LGvfDHt4MUkk8hv8pAUDh6t5XUVzl85xFDxRrKuLI5Z
nnLsDRqt5Y9bO9kb8XFYe9Jq4HGbO0A4u7JsnU/fWW1d56YTKBr9uHekAV5BCoNVxQhRRbfeTef9
qgoLNaXYKUmn08Xl1kSae3Kjpea2aLYOKBjyk0AmxV0H7gbRQimeK8K0vHd8ZDsfgE+zR7cpuU03
HYKCFnT7SuAaFnbtd7qabbUBDg+P+LPeumy1Bg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 40224)
`protect data_block
xQ2ESigWAo0q69rGYPKW8u3uElislQ01lq6/7YHi49rSzfQJdwMd2dorr85EQ+R5CjiDVTdX/GHt
3xvakANYLGSa7jXU1/CPgLyHe5C7tP7BJiLU8SdxZfgxlvO+we9/J1deyiclASWPhGhuS2RTX592
Nqeg+cpvtgsDXW+JOsNNVKz3/JvGTI8ogvfTxYZTw2eJi85OYolZAY7XuBpM3S+LVEJ2qmKTmLlu
TgOMucbKUPTbwReM6I9tCVyds3t9LToEo11yd+ngtDAFZZRZo9K723KmNPDpjKSStl4x1oqeScI7
vQgI4/Sgg97cAqw8qvQoPqZbyz0MdY71Zh4zOA3XSplx0MStFnt7dbY3EMIoa9ymbFcBBvlnfkjK
I8rViZCBkpiU7JEwksxXemb7/8PlQBl1wdcIycs/zbg7cAwU/x6Rklaopp3t40D6pEo1tQZtKSGV
ZSkGq00tXlSgFFCow0zV+RiTTWZdGJ3ipYGte6zcntI1+ggrt01egIsITyEw1ZeXczuHtCOZN6+9
v+6O3pc73QD2PGGaY0MG2IjEupI13uQJdKLMAYlGNBKaifTmNtKDtz5xDuhQZ5YwDaq2J1Ojzdag
9ey9TRMZcoGEQbR7EUsmRcaud8fe29jpoeSNq9ud8+bL+LyBI4BZidcrgiyMMgm31VrEQbmD3XHC
vhEqLt8X+3TbGaLrcOtNpzHb5Dfznl2V2WVkU7qj+Xpc+dlHamYEtNQPzkInIdyCvOnksDYZ8sdX
ZbhEYEfdw1s97N4JkpSrRnUoFMusv2N7pLX13H5MqmxH3whESIqg9Q3RyajVEkbR2U2xhDvMZTxe
Ftpf4fZzo0CKjax+tatLHN9Su9lMMclU30Cjd7Hy1hTXcbzafN+l+AzMHWWfKWAy2cojTswOtzHH
VJrxMBu7stPc/UHGmcDp0P5ISzrY/3i0LeZD60ON01e5vVA9vpLlBQcXjZoe/YQu42ouyr4BmX9K
TENwFBl7u9RTvEMI6BUajsQbQkgOVhlD9cDnJWlmFIE9gcjFWR5I50qpAdib0pBeNGcldQ0IASVS
T3z8By9ZiOL1GdLVRZH1iSKvc3nLH1ddpPRXvyO+EhM/QIo6Gu1reWU0fW6oMT2rQjUGic3M26ck
MCvtumK2Uy9K2n/tFPqRz7mNwfsTgmZO7n++4K/FpQncYWhiyDBQIwPvsliCNvVAGfrWD9BSSp7U
U5kMNGy9DFNqaCCbSDd+0BrHephoQI7gtRwbCi4lgHqySCdVxl8D4Y9nHS6FhGCFoY1apuAw+LmU
M44EZn11lu9LEoSA27fqVcvK/JN7MAC/4S528dtl58TRUYnB8qjluaY0TKiltLXO6ws6v3t6Qbq0
2A3t4E7PT5iejoInTeI/QZoNUSoKmwn+rqqIm2R9G423GqJxaiKrz33/A/KdE0sTZxuGTNwKCpv9
OVaswmIsXDUY6zte+K9HpmNoWQC2cMtui6JReme4OGzPesA3TIlbkp/k8P/8wAINkoDDgACD0HGJ
M7xVQZgXDi+583aTQe8pWo1U5iwFvUfVhp3M0j9m5ziVXpYQg5h6Dh7Rc1ZndHyrTZ4cJIWnHja/
95xCrSiCr1W8/dpWyUQAWBxwUxjWpQpNWfg89zD2AY/eYigWOr3tdgeCP1rxvFtvsll1MHl8OSMI
6NKRqypKTgNNNyDdD9VU/YFlE4cV+euU/OW4axg5xhNTsymKslylkVCWLpIfuDeggobkYeVUAL+p
76wSzVgmcwUm2rKhRbjfpQ25IsVvLvDpHftYi5YLMUlWz78KkiW8/WX/STsNun6KRId1r6aK9PaA
gjMHlUmZ0gLMpAcNKOlof395wQsd5UTuWBTIfKUDkdNgpWgHWhK1AvFz/+iAygcDwhgXGt5YU6GU
znInf+YjkHlTQdOTfcKyw4PrOZPkjmEU2oS0lBBQPkzli14AUDTXLUhmM6FmJxYRZuys02BSfuO7
WhP/KkRWYZYyEDdZTutAqtvw5JkVKETZ47IDf3s7lenUNNH3/1HyQcpkAnnF7GnCPcACCNASQ1ah
+aQ/OgJjlT4VBucupCdabkpj0uHyuxjshV0V5RvxJ/uuS23cARXhz1ZuFDm5RyKgcCi7FYZGtIea
1AA5RaTIHpZQdanPDFMVe863VOuphITDpVMNSrOkhH5Nh5CEi+SzRCtp2C907A2k/7IqhWYdvjsx
LzD3USsfzy/WceU5D/Hi+lxsTQPFGtq062c2spiXvEYPt2XR8x8RSthdTkUtG8VXwPH5Nrl+NYaK
KjOr+NELvazWour+X5amra/ExM9PO2+cyukwbl6a8Z6AqFj4SIhFthZO/CeWKlsPMt+G9cftMiY4
ntjG4AW9uiCncPTYFAOipq4OCKao2TO41ES0E927rQ5parVEBW4gPg+lj69XJ2Hzgf9T6MzfjGDZ
HcMmgzRZYZysT1BGrPixSx/vJSPLsx6k0pQGOH2JPXdYE1EtdBZIpjhYpmRwy5bMNfNCieS94z2m
J0K3QKHU5DmFRuggVIQWS1g03OCI+Ro4fXy8e7N0OPQWh4qke6sJ3OBHf/YpoYYK1+uTibjlE27a
9cV1ACofeu3XQToTQBsLttuKMenUxCUZ/miLq7OW3ahPHqJU22tlUS+5r+uG9HrzWjlEKO1sa515
uGUnBnjgMC9zgurtvWVUpcL3HjIF+Hw//Qx3mAfnh6tEK//SrScDOtXL+JH8JFjgd1M+2e8uhOvT
giuTp/Bjwps6SzsNttDDLq1bkaspz0oPfihGQMG85q/w49D/yZ9AeT/oUdNQg8Et7K6TsPnX7AFs
Ioxjit4FyOK0pSqJua08cxhQ+VqWz3YaZHLl9p4DUmxGb1X0XOG5EpxV8IB81Pk/puebdrda7zqU
/FDfkJaXApYeBG+2ilXnK0U8Tf+lqvq7UwohtOZwdZaK7btbtuq7pIOH7A3hJaKA9Qc3x7DIKWiR
rZv2ywYDomjKARNXNnKfwcpkA6mKsx4faoZjWU8tA+bcjdWOKXgzgRN9aY4q6cBYyAvJQFhua1Uq
SzO7go5Tsk6H4ewjx3TJJKBM7tIz0f1inc8k/jLwX81gvEcnPXYbBTnZZKwhouoffqOCTrwFrTqe
a0x7UNMZsxNgnZikTt+OAntDCCyoWuuOl2W/wlAsEhRjFhtXWn78VjsDasbBcxPp09GlPJzh9ALs
nZZjm1Bp4Ii39giJ5xIC6YSQgU6M4EEhnvvOkLzl9ifyWQhJcFMrEl5L97/18PLpDqP+Bnpk/uAi
cdPHdfBVVKRaojToAXHukUq4mUjPX9dQU6IBJM77ed/q/sFoHSOBlUurkJ9h2hvDaMvf4gsrwRig
VM/EBXXAOrGaNOOBK3I5xTksQqRhPXV1SvkXgrt8bqPAaKuNsbWlrkoBAv18EM7hyiA5+sXPpAhu
tqwQPxOGv4izfePfOX5ja8SRnFyiAwAIuB1455QGVTIlNy1gOdNnCoMyfpWmSO5nTCXwZ/ZUq+DI
v95+OWfXp456B4tUW9yPFuwaryVNT4niJD2jEM+bEpVjSuMUAL8fGd/iEs1K3foj70LwNoT8Gqdj
0tf7IdQFJNEBdDvowid121ZCLLvfmd65GPtIybQMvOMD1WvRcjS6vXhNxUosB1nmJSvYZQznd/4W
GvYtqJkGpkzb4len55350LSBoPQxpTb7Ade2/UJa8rBKOu84Uexdhb/cVmuKdrCC1hVcC0B4IqJ4
8KWJuaj4lhMVcHhGT/ZGpwLv05TvZI8+dmBREpSZFvFFVPfyM5xOjoaRENLiGR36tHWtGd7sBdDq
F+9k+TSZNjJqj2h1KA30vaEa1YDF2kJM03xMJ4hBaPKXcVo67gEWEKsUBMSKExdPa0clAAosMLFl
FZwFfPP6etNoChTshnKL/rM0gsCaubZgcRVN1WpNpI8kr4V/3Wrg97fCeTdsow2Fxxyn2XI3wB7q
V0aloJ6d+cjtKE0dtHB5i7UelOwASgb5/88R9oizxp+y92xMQ12YqMHiSMF3V5hP1EoiqCD2azoT
orIXc0lrvjiCwqY2B1VBygEUBgIztrLRU9flekuT11houhwWmsfwn5r6jHo1FUF537gkoFtWjXcd
ArxjuOwqdLyOUI7kSY/VKHD/+WnLKbLui8uNjn9ULyYyTU7zUhoSJ7tfJFj7rXSU4XdYazYRXtri
8DTVSSmDWRVDNAnnTd56UEXa6qzSaD3MfmDw4OJbpH4LTzXhI+yqV4zv4l2HS9JWTWRoJTZaLmCF
BkeF//QQmpvOSJa1bh77aNsmjbz/WscJ/q/qrtk8pR/+1HyRMOlxfxpYiW/4648JllLxmjfAlYMf
scut3KKE6BLP1KLipGO8WEoVtJCYC4CB5H59SuOyEXfSfz9cVZDh3hpJ9trrv9Yi7afTqmQcEWHC
kOtvZtMIBY8hLVf8NnP1C++oxggoLU+jFaQwhvB/52LDBH0BWC275lDW068G69/c7ejiLgYXXFlK
jc/3QJtJa/6ik3msS2PQpc+bk9D6huUqNBsNPex/FEse/GdYDUcyS2b5Kbz8X40IsvpT5J89CIAU
zSSdYXFyAeTaLRMho5sIX+HINdDV0v2vhoHJSLwWhiRiLbpgya7118Qimhrt1CFkvYedlkVp0yhO
ySbukscb5AinZ8fdgnnerC9569xAEAPhA2pUe2y8HlYPI09no3hsd62xs/KVyBXtvIL3A2W+9Hxh
63+4xdNGV1+KcdwZxuU1JT3oASejQ1/TXgUtbDRxy4N+nWu4UO3KmPHLhkGW/sR/CBJtWudVE949
CHnyW9t0Anp48hIoW8QVhnCrqI9vqyW1JEaFoJ3yTvLTPpLVESZtWsNp0VUEfsLgMaFqlNpzv90r
Vemo17Hr7zas0qPnvPak9Oddg5wePkAGLBEH88+qqMys+0QYqZDOAhgIxtqHGg+IBcMvsFYML5tO
baHidYZRiYod57/DAkQrlJEpsIpfqgQa8QT3LqLiWDaMLL1T35QtU2ssrVXLPzD0JwNOhP2/XU/F
0MFmoKEtpZq/gyAySxJJaJj7kMtzRFbxy5asx/KMCSJirlAvA0jDMp+L7rcYCCnHOsAuFZxBGfT6
xIvRqyVHph1T/wduxUEKOcPunyQoz2EXsT2/5Vqm3gykxvGAzZWF4W7LRipmNrPC9ii7daFkqzdm
AYsVCa5Cp6JlHJktKcXIZr27SbayhFj11/o/kMATjzp2uYoGR4LtTAqC8MZD1Lx/bdqKdHjcPXYE
Kzhu3xA4iHVUGbX/kFmmCGr3riq5oI8BtMYkv2JjoFCcYu2J41Q/Cemtcos6M4dIrUCKMHhJ/d3F
o4+FkgrOxtZNFfVOBIO7OWGQQ0aGslWnThPtgN8L5UOyrruradbbC1U+dyolwdWuWfg6C5m0AbDp
v27cY0bgU3Za5G1OxygtpPLFw6NN2wm9cVZmMc2jjOaUzlpcC+qZ15oo2QxDYnTr3Oj5h0nK+9Of
LtZVGZniNJIH2P0DLT/BKq0sivMZMeHC7A0/FfhGHcZRwgVq6QwQO5jVKEM0hLEcE6+7Yu6ueOvo
Jnla2UHEZRKbMyOvg9l7vPBrU7gSXvj7xtW021EW3ejSzTg9fpnNHGOO9Je9tSXbo6jKzv2yrbpD
MbObP2FgklmE5nt6durHXluqtew/F58tb2dGSXf+TjTqffQ4p4jXXF5mYeskomzwWiBGrqr5BKFn
rQS0ei9LeSYM3YFqlVeOlFSgyDxR9cRpeCSw6/mLiNm6TTsCDGr/cfBKQY3+EG+5ag1mM45rMLFE
cZQCvUgJ31WylR/QG+//BuyraVC4BWq5oiAtFHpL2nssa/Iq78tPmQJTJNHOQjPhqTMoGQEkp9D1
IXu1IbtCs//6gWnkjb9kl+FujiGxLqETveP3wF7s1Hsw7IgdF6f28vXYYd4W5SL5VJplnChZylFq
C3lrvzEdCKYhqVf9KarCZdk7CS8LI2eT+08OaM1oCFhLPRhf5aeYiUWS4fndkgOB0qiJD2VIc2Hr
g5e0V7oE+HDu9CGJ1r43n4TpYHWC5ZwP2Oi4x1W/z0WrJw0HAgMyE/TF0SaPfezQ3rFGuYY0pHtS
DoFXcRbavcMc1MgDUqCI8w/my0W8ovPItJe1W58w1RgPhJ5Nhtrjz9XImScqyF3vln2DeA0ymoFM
Ocfmsql0K3EYaCzY9YINuftZ4mKixSwRAPgTg6ATJkcjPfwERgTbQUjimTRdzv3slevVDhpp6KR3
o23vM3fvCDPW8SM+t947if5fcZ5u9kfZMY0BgbajcNoXo9SIfxw6IrZsyCjc0huUIb0xu+wMmucO
CY5lBvqYaho88G+BhBYoHZNxBxfJic6vFqScf5ceIr0nNZ64wm7d/ojNlhLNCyTZ+jl3+IeieFMQ
BULdx0DPuG91RxSWqakEat1UKodHK9qOR4BcuJb150p4HwmvjeiFHSsMFRdQoomazDe+hg6GJSsS
xgpuoccrm5I9zuH3TB7do5KGi/0u3Xe8fxPot3Rxgtv2x3zFLytA7R6Fa+a0RTh31NeNDBKM8UIq
aj8huIdcksjlj1J/XXA1TRot2bxWDvJ4U+NkXj6DmKkFuQkU5eXyaHkuyR9DjoNuwRtwPh6lIGQ3
IH4qHwcBdt/WEaFSRyWHckGgVaXhOEUv56h4YTu28YJ6PNiJ+pdHb3+Pk52vYSWmNAHDun1bsKGb
jAgWGLoEOTQKdKjV1rcYGEAfW3PDI1YJssM4sxqsGoa06RlU07xxx2psZC/Ezm5pudY/MZiqbOci
19xOWne7ajG+EYggke+8+axpa/azMSlG3JhN4eHB8wNTozFx/6OTxjOz3px2prnqZKRgw5lYH4RM
/7EJ4TwHA10RyVrRQJacmCKXQ9Rk71WqVK4x73CogLx/D/RVALw2olKBej3Lmah8Sfu2YfbMHJpB
CXnYI22A3XuQF2oqA9X6b8eRO+Vl1PIl6YzKjTjEFfqvpeB9ErB1ehONUeaVwzLA2W2/1UTSL3DF
a0lyaktU5k/UOZEpT9/SuuYdyZRVNb9ymcNttNTGHrMqtiYyVh4F5b5PTMwc4G2Vr9NIQh3IG40s
dyPZu6lxnnr4UwISfR3yb0+Di/tsMRuOPSknR8o+7uXivrQt+FtLzhBEjHZLH1resdXbF0M8H7Lw
rJEcMaLfAF9vxLUv/7iENPM4OfDYVyIW+qSwZ8Q9gT/E54YBxPEywc+zrokuE7WUZht51vNUkzFf
uQ0w6BC2f6fititGzdEyvqremeshJG9JBDrx9zRYWf63b2zXwqF0emj7At/uYhMSBSdlvEQiEKHd
VFvMwxtXnKToxtcjJsWMtiJtdGKutVJ/NpksU2yzbuJqmEInUrT4atq1BAkZs1G99MNG4vXE9b72
sf8vD08biGVoQSbimiNRN/VMINscuF3on5lx4DSGw2fO2lKpRmXK4i4T8ciaTJJ4N5EJjZ+qT6pj
UPcCZUVG4n0CUCgLsgiZgVu4iAjHKpDj3jP/Esbw+sTy6P22Aej66PhvvHDqTJAeS85/ty2KyA28
y31GylIdfZeYSV4lc8BuAIG1khKnANJoOfdh37IxYhB+s2FTwAkN4y7o5dQpeyp0KMDvjr1TWBGl
YYxNlfksHPqiwfhlzv0DBLgWMZi0CX359gPSXcOrkVhzQnum+SUqqZEkQkCD0Rnb0+njbenbYYZC
G8YFSzm6teZx3+x2/63GW6yc5IP65e6mSQLK3abbmzJVAxO9QUe5YSmUqXWuRhgz/FblJfFkSaJm
5Orjj4B0E/OSYIzhycH0dCFpr2fRpNaCyS2kITwV7O3Cqq8DGbw1Axaw2l4msFW7zv0E7l+nVmyX
TowNHWV1BfiiEnBqnvu0iSZaIGyt3zvPUcABpzH0OQ3qsBofykE+arUPS2DQgHoDl8eFQED/fd8q
UriHAqGN/dp4q+NV0eHhezJr3+uIVIkbLuVrt5qKyFXlyZeUn2ngXar9rAV2XuGNjQDKff9AD2a1
tVsf+Sdw6mBWbDgxAt7g/C0U4eFleGUUUvoIXRXw/6D04i0C7tBZVtaH6wZzx9lg8TDfzWIRSN6F
D4xE62gRujrxcRS6E8sVI4Iws3+t8Kwq1S43pZtIlgpVrJ/2BvJj7Hpy2ng1oCA0JWweWYSYcRgk
SF92nOsNXElA6LzmKyQZR5ZAUWnwOZ2TFKcz5Y4Jxox0LhAITpEi7rmvhQIasH7zBiZy3G7CmMXe
zUD+UMfwfTHYjSxGVMvKl1SK3BxebeCJUjfu1CwLRERkLqV9u1ILf3tgNK8Wtu6XQgzvq076ZFxs
AHRBfGz0O63xWzRgY1hPHAaKxLLWdsfzzLoBDgm+ibnL5H/qLszhaFmaiH5g+MrgIGemOiE2bbSo
HqcF3LzklcIGZvr+s/+D7OIW8aQ3ep6AZ9FI+l65IeEtYg1TcyX7Lood8fgomYkv8TwwH5lIszg8
LC4gINXHQzqkh2YWd4fnzxSL7Rdf4ScdPADgjn0hf6odYGLJ5eHCDabsT8p4+/yWE/6QH7DOhh+9
9GeP8dk/bzsmhFvEqTNPcwZ6ckKQcyIStri/UoqfGjJFc1l40uBs/77hGZa5GOti/aZF5JLyc9zJ
yxh2tUp5mfWIBaAJ5OM6+dZgUc+k/OLHHfZYTNZHj2cwDBrwKat2A7JxAkPqLdQPCDg8TCaPtn9W
9LBcChDHrWlX6Zh9sdJXarQ/f6D4uQ4yC4wyQydsrwPFJh9SlTm/5rCspWqjnL/s4qHnr98UW9A7
VxJQLyAfTobZ+dM5L32eTxczAL8BjpUBX0PWEPKsgX0ALj57pSxnrvOsRqHs7Q4UG59jJwv/5S3Z
yeyvE2kQx93TXj7/G4/BVW1iGTNbSUjCRJD/Lw3WAmk5FLUiAwqVSgOvx6FdUppoxpF7oysjCSiY
2EjhvV35jEMYAonVhbQvhuCoHUSgZqmVKB1fQXET3rzVk4gVriKzRIUaWUFkCLrHdwYlezutVADa
zwQt3yj6EW68rKSGh7MeGdyOXfwps2PpOcMguXLdeib/aY2/aw1OaDddnqhcHhlQbgPZLubgPzTb
9UD8oKviIayD6TsnKk54CTe3xsQhjKCmceXKF/UIeyU+v3//ij5hIEB+zBwoRu8Xt6hTBoHb0Q7H
94AT6YQ9rZGDMFJfB83XLgDhK7ANK16lWM7bvLJ53xBQ4G7WGrKGIwXLzSnglLikxAVWmYBNF0RJ
LzxcDR1jrbRWLmKG0Ey9CMAMYm3uYP48ecPgk2032mr2exsQoXk0W3e7or3l7MteONWVPF6Q1ZDK
rxk4GGa3Sdxw/QueLGCQwhcQmLK35Zzn7FQI5pD7klDzInVYbswhrixwmwaPWUnDva8Jlp305jnQ
EvNtuzsg6x4UfXV/atPJKYUaxjteNSUpuJan6VprJwJFE/7ARV1PZh+OFDuB0X9TwUsJKLkjZSlT
mXi7PsxbIYx8UZ2tm7WAhBfgWhcOtZ0mNSC2531aXWnC6MaO1PD9jy/sGjyVDAnmrNEje730YUxY
5KiEvPjAdR3WXnA0bucvV+OS/dbMEwpOhZ+bU380xNXmJM93fXzKhZazPvX/CXs6QKzdNohEPudh
E/3DAhjKMigIBuA1miLI79tEz0PkxC0UJTmGiOmjhTbnqfTA+W38qXBXeL1JmxD7wu3NMCgSID0k
W2H3ZvodGY6GAsH3zuo0TOd6nEEqcatr/ghogwyLqRS/dF1dLU8JZF3WkSL7pYrm4ZNwqSBynSkQ
0Lws1sbqsVFfVS9xMW6Z4YJROokjr6MuSBrLikYiO94m1iundbKg7okejdFYCDJv+6qwemQg7EiI
hLDKmhJF+89I9Zr+knYarmc8R5Mmx9YSbUn3kFjjiPaYcQdbEs1makBkuGtiyLQxh8cb6rcx7LAE
rwPbOb7lQXKyTqD5uu1FUaoGGeDV4FsoEJAmyMGBi/8gDC73qc1mi5cGnsqR6SjAAgBdsyKUHKfa
ALbRx/BKNs8sW00xTRRQj22IC51gE9empUky9n2E7KRe9XV9kKMEppwnfmv7ymNsCCXQFrwwiaHX
A6qMz3EMmfGAnB6x6CNVBrC4YtjVW4vydv29v7jMRk2pCfbQYm3zbMlHR2lL7AGETUphMb/Lbc1f
yHsIgrOKSdKEbt2ZjvkDEioyUtTmzVR8ld1HAGFhXVVK7+1/r9qHCssTy4iXZ0YZdLcVhIJR0Zj/
NUMrjXgaKESosElVqldMXZCT/rpINsNJZybSxKVr2gCHBCT4Hvfl8tCHK+/Yqv+hoi82q56pOUZ/
JCxSVker9plY1iaiIyzoe/wpkga7sbRh2DgvACTLJpv8tn9q2AAX5Pq/GSD1/rBQgcVtAhQlgbsX
dCw5c1yIbiGCXknePhXwoEY/ACaIL2nD1G28h50pxuR2Nuqccs0ztZi5t+ThD+7Jwjp1SaE0nJWz
6jy9Nuz1hA4INGZW5MhyDdt5E9CnC7PQOFfV/34liPXilUACgKJ+SKbbIAKMtjORWn+WwRiyl83Y
MeS01HLaTCCP3B3ELtMjgAYLRlYim8lCSylb93j57GaQlSYuuqgFo1gcflh1l/vsGat+4Q8s0gHy
y1EfBCNl13yHnVsoVKtYc02JBXV58dARZ2pjm682azxNPRqHk10gNiMJbATHr+goXHiqm8rRXXJS
IPzqJhVaA2e9UuSu7cWseLmDbT4MPIliC9d+OQFTNwLBnNtcfZ8TN02kRZnxxqsJT92VHYYNVzC7
xTTXYQDmKU8NffElmmL/4MXnXKU+qpHwJx52ybpZ7fPxPVgnA6iwqooUmjZnOWah/xKECuk4bs8Z
KHxe1YwP7uf/FeXgOXTaWQMP/ctw5IDEsQl6520UXZt0YViZ7rgLayXpIl5SvGbRCGU38CY9kyPT
JwqaXpE0V8/beeZbzJ1Hvazw6b0yoLNXsiZWZHQ/gwsNoHXCvEUEX26C5+3pv6A/NdfV2emH5RMd
CTlZxq11oK3+BS7Zn03gMh0jR7uU5sIc7RvoLpD3eAOlm4G3VIoQBxXdS31gweXK22lR/9N0JO9R
RZI/0i4tFA0OXcKcv6HKNuu1QMbEhJdCjP7UAQXgAhBRmHlmiKkafZW/jErJo+2gOleM998YhKrf
cs6P623IBeOd9esupFukXrkNKYDXSApysBms30Oad/c8BQ9ZInPDZDiirNQpsYkYpjdfyxWxjdzQ
LnAeSyAw3US2EQAwMExKnz/nV3fr70R+sjwqxcHwFMun4+5HCh904OgmutEKktkHiWNFVU4BkFAP
xSliZaZWd1EJRl8alwp/ApBeE8q4aomcRmXMgeBuebDnNZ44/PlHJPOBA3L3JMPx46jdAZaKaNFy
EqKc0ro3dXo+S3jRQlJpSedhwWyFU/lEN3zIfZJYmnkuY0dQ/MhBHayxOwZvWvMFP+LmipqiXZ0W
0byTwg+mcbJfFtKi9/k6rh8vEEAVXLHvD5byyMrH+pWpqvcZ6et0caESdanzeIM7PnFE/0vMOvM6
ZfRoIV4A7v1H3bCVdLngCRiOcB5X9qZkR+5w8d4K+J6k5bgH3pUeG0a4YcDmRj9DdH09KBO4+ymr
Qhhy+IeFRdTUqU6AhCYA2pOFqWrddSVaVBjlOCeDl0QddE7odlrlRYtBCHSRJ0eSXdnzyTWDeKOR
UG/G/esWlKnvrhQ/mhKfMcs/umJ+hGJHo4sZ03qN1ptQEmMcZ5c1S06EFou1BpyYHfxTJpd9WfgT
1lKk1M74tiQd3NubgHNq+YOIOzntnglx5Y+gQ3p8+4xcug+cuUjx83caIBYgxQc4ryVjUoONLGxL
h3/xmR5iDmJD9Lmx4sRPHQLLLSmQwZOUkmFeCEAVnp8/QrhPdtf8VuAlo7nz7zBn/U9CA7TgJgB4
4p3NpL/MrksWUEi7znzlaCBD8fyGSSFQEqSgWH10yYp2TzyQAXHUxaQkUIBkkkCKWUoK58tJdNps
vPm6NF2bJokij6PZfr84pCDfMwwc3xvsJU9HXPEzuj4bYuLL/5CzLr0mVTtGm7q6RwnKC/VJ/N9v
CdUIdcvWley2mVJlrBG2VMX2QBjn7lgY5YyEZGb9fe5KjiDYNDeKD11sNZKzlSvUM0TxU7gn1KEz
vp3u5oJ7UkU5u61pPGj2YuD+SdjjknNyzy4UKM9dspBR2bjhHm8QHUiCaa8B+Ah+ji7JmCfAw7he
OZk6Te2KgxTLd1xIlO8K6+MxcS0qR3o+IsrhHV8aKTaPfZcROBeD86AeqaHl0SO1CrlLBeWen0Em
R8oX0LdT2U8ZcWV4Xr7ZihzBGmlxJ0Blztm0HtHfd86RJ4gK0118m9WJ84pAxW7KYFD++Wnj6uOq
kpNxPzTYvHdxx6PL5bTLeFJchS5h7uzSs6cqPocu8OeAHDoJ9UoiEMz0OQXI5lFw03D9BxbtMIQT
odz2zgER5dHLODPYeLljB2JDh7Uuo8zCkK3kF1Hi4zZsp5gNjesiPxup4pXLRaHvBOi5LldagAlJ
SeVeGCrpTdAl2Hyq7Pbr/G7cwLKdZSgUvzKfMumCE+ruOeJAeZerM5N439Qnn4ZlpiOzDZSm5smx
bjUiJZOITaLAIkk09dIiSKG6O4ZUhVIBpsSqt98HWL6q8sD1vOj1i2GI3SvnreBEiCAb3nXsWP5B
pe3vgI/jXQJpnSdcGtCSMHpIxInIH3MQaSWtytujYmSUKtSd9N3jueP8WW6EEwkjXG187ARwIPfv
ZrsFsFykf2+CrBG0NT/PhMrPIkQFCdA5ZAJO7udRR8HHgBGogLf+6D5YDLc/PcqpqGkcp9Nz0FcE
xdK2l+DtjhR6tJJLdKw6UGihny/rZc379KeOKNYNSZS5XXhlA5dTV1ylupL53vARwjvSiBOjYys0
zWPfWWCRkLXkYDFeW8NGK5yDxkt5MN6AVe5euesluX0PsmovYkKq3LW1xetPcqd86Pv8FZDJzLMt
EpaULJz6irmUmDRjSVrYOICHP4Gc7vwF664J1aR2Hz8QI6Bg6ePME9a4I8AvgTNdt5k7lCsRKHnz
HbC3V07HS1KrmR/ypHClSdUuc2r2F5FqbMJUY5Ft/0R8iAqCPfxRsPqYrCnJM5Do0EFDpWqccoP6
F+g0WSLJW9X+tq25SUHbCae4BZyX6MxrSYlxryfGfSWjBpZS4ccGATyEfUh++ivTticQxSQqlPw6
HwrYT/xh71PEthOCtXuRSTAfVg7k5r8UvcE2hQ3KF93m5dZ7ZYxgEgtn+dHyAIV5bxivPUFD/rv6
rzXfTFIKgJr84hw0wpdFwIpftQggXmd3A7y7h4jbmogPavmTktwP9ckopv8fAlKSb/PDr92igS0p
9h6BrDsDiZvWr6NXlOl2H0qJ4qwqYHBql08bq2ZLuCNQdj+Cd7CZbHUfIFmiYz1v9jFxpy/1Ywcg
GOOLP4j/9Z5c8IdPOhfDda06noKMOApy9yf5r6wuSyU5rZEXyg7m8zjxgxbgmSkbzEVE9FbAmUV3
iZdJblvGeQS+dmreK1gNJ5wQPnrX2guu/AcUjHVivuRqiG4GUSC1djXem2JfOk5tpjIqNK7DY9/u
JfZgt5GyID4jn17sHsskykXONUJiO4tM7LaXfEnMuXGuvons05YdX9lqrWGcJCnzgODBgC3krtx2
jDDgB/dLvZ/D067vRoMcxnyuJTNKVTAEDoyKvQASWRinRVsw/3GajfvZ14FGoIpPB406acHu0/Ur
myQuwGUUxxRBT6176FJft2V/vgVWCEPH/DvPzFvEDZnE2BsHbMJYMIBx7FMqlFxsh5HFDlQR0YPT
n6PGbuOdWDJ8CgIBmSjVO4+qH2200Rt/OdSeh2YSuUyuMYYK4kwWufuMpu9a2tu6SVQaxjlpSGYs
zxb0rwBjREkX2ax7645qPOfvLpAtI/iqsHckAkVQB0Qg2dB57PzAfaGT0ygE5wcqjxEPQ6N9/gtn
O7aW1RHuSdly1ewDRVHe+GHSOtvOC4t4y8OlDycOsQkipvQEyx4NPyewi3UYPH4NgabiSTiIgv/G
fWbdhAJIB8l2XTZ7bd6k9EtbRWvHQPl0L4KTey7AoYcuA6ohtpjyJtHivVFD+K6U5Ll0bU7BjU69
VCrvkH8MU7juI6qHaMb1y7uu1vN6RN7nViGEbj3vJAo2fPiIoqJcUBjTbn7AsTna7+VPqkVwaxUL
11qezBxAY6CozXW4pgXD74U6Qi5zQTxElZTDTOZXXaw0HMTnQ0fQMzivjIehCVyQeF3J85yHS8D7
P3e0V4qz4Pg9jEQUHV0hxW7R0ptHmXJmYw/MUlkDz6LpCK/y7ZdF+7NF4AmEKFjQnCwyOGpgpSiF
hUXYbZeDZnCW9jilROI9BhP1gWAUGnphWcQopf7DuITp+JD0mXzDMgw/dQlrOoluKeocy960J/Rf
uTBR9+CGcBWvbzHrR32knnYFrC+q0XA4XK+xWS6RxgX+TvJKDsiCLARVZxdDyJ8w5pz5LZCN61zc
XxtGDeS0xTGJ4C+dgu95VfCEEd3WH2f7NTkSI4ptFR3wTCJaprdZ7ssFb1NI7Haynv1NjQODSJpK
d6qo+IO2MLWm+DqU1OwSrhmuNlCTdUK+Gai11UC8NWG4e1hr0MQxJnqk5fLIDYebKSFvFMxDk/GQ
6G9QVQZibGY0AyQzpYp/lYQz1+q9dHcSiuv+VR3VzQPZuYXUWkBmMjQSfjDcqqVJKOdJO0GKaX4n
b+R/ZA6LpWoxiZKBIgmeAxsL6qCLXYWZ2ilKVvWCzMImNrSb/6mGbWK542i9UiUhyV/2I7yTqHqs
Tso1NTJAxOfPP9yZL6wbJ/JqE3+QabaGmiVfbW3hFP9vLPS3Ud2m8oezLIByYm1NDCjojX5haNz/
Gxi1O7IfJifkMSveRqFY07dMQ/WGxiG4D9Ho5RMP/Gm7pgAtNQ8iA0zKG/IP4tscXiIIDiKtFVOo
CISRHtefScSGURj5a5lXFr4JvJ+96eN3QUqsGyIOlSBOqFvG14T7VfLGpvDAxjzT/1WbthiIKEbV
x+VcWpf49J+MDm2zstA2gMM/jiP996ch0nilKkrRUMRscF1GA1Sa8FK8LGfOKR9xH16lftdYJZsq
5QO05geapvAGODRUpUoFXAZ7Sr41ioVSYxPCJ4MDT/nRpJd3RMHnxe6pzerE3xAwCleHX7YaFKJO
TABpT2W1T4q/B+IxTXOmZSYQ+4xiV+bTiE7zPjOFPp0kY5QxbZA3E0+BwyH+vigi28todifG/RpX
VVM6alTXsRspjiy5ePliAurhumr5M+aUadYfChafonqvjvP8S6z3KpuhF/t/Gh3wiqpn8TM3wZIY
P1koN/pDWuvEFXPoYSRlSzbeXxp+GhbMOwe/OsqnkESJIofA/MJzfAwznjjiOh6qUbS7ksEO1V9c
88djfu+qOdTipb6GX+iDfX/nOalyQt2lxjxDlNFceNzIJ0zpD9AK/VXfDtPO3Kds2Q8V/1iJ3P/b
pUVqQrKArM/kwQ2TzL1uts79Hz4DWFssEglys/yEmdbrAQ+XPc1BMC9zrNvHdQu/Oy3UjvrlzjT7
Yf65dAhf0sIt1tduR1lRWkAJ5znwECS/xW28whSoi4NzSdiIBSXi1Yov2+5HR5Mq2J1WHsJVo9pV
lQzhHDtsL7Oo+wyRbZHvBA1cKgmTzGjb++p0ezmmtKJUHMgfRYOLdm3NqVRRjWVHa8kB1Unj9A5A
/FSKzgTBzlwco0SJtrzNY0uE8ArrCmuVtJPx6k0XbEA0WGvz8JllQ0gJC2NpW9ZTp/bFSy1zJJP5
OlEz+jJeCGKXJ4tlOAGHWWlMw118Ax8YA96agnznAoydHTcDmIGykk3fuo98ytwoqBpuqRpWaokH
6iM9KxRChil6wmZwKWn7KtMPHAKZOT4KRC8NCb+JnTxxnOQe3dwp5Yzh+PQmf38x1dpC5eX7Seiy
7Xe106bIAYJNJIz89NjGKkJKl9WCvNxbGpBIVDWdiTLfnoumS469YBGY9js3epcnuKNPY8CNBb6n
ykW+NlqwIC5POKHjtYtfB/WNaQ7Sj3o3CsC2QE2dS6i3N5y947xaDDeHCzimVxHae7jD8MrdDcOw
icedJC6ZP6HBpfO3/C+L4PcJFrSHfhEHz4vRV2PFoDrmcdaoJN1n2b6rS7BTEhPQ37OqPkreShJ/
WqjnXP0d58rc1pkCfB/VIhA/RP3I2Sid5bYziHblLvCP4P2lGot2xN32Iha+WrW622VrWhM3B549
OnC8c1R22MDe+S6JPN/Bf9R67BRgSZ93dfdq6z1acj4Po0rUCChBm15Nvpv5v4ZBIPTKGk/K0ZJn
NnhEdmARE1t+T4iuC5yLYcdV/CC2QifLLTmmK8ruS+CM/PihW1mazYquKiJrHF5jL6RXf+X31enx
IB/jKHcXF0eiSqBCJMWCnnJZrVyMcbdYyWb6ty9eaFb1bTMlpHjX8KOTrKTLsudw7uyPcDgrDwaX
w4zVysWG2tn4wzahgfmXywD0V9NOEXOBCxnm8aeVKKkQt4CSvjwDO0tv/Hpo4C3Nez6BkPkdNlTu
l7vbevLEjXreazTv4fuPS+tmRiBxZp3MblO8OjbL7auq9MSBgVdVfFZz15VLmVcJ+foiyadayfNi
PHKix3Vgh/ZdxzpLhxRf4L/EhcSYOj/QWcGQyG12mDofvKUg6vy5VbS79ty+SFkJrMJs0dOQOaA+
1S24X2Gz/3FikGONIke9BLZKRs8CTWxLnMwc9DnchF58UAnzzb5aHntl2GXxOsOZlYRBJ8AzXvWH
E4MfhGTnxLicckNd0CxKFUVv54xO+pez/QvotfWlVi1eyaTVGCEzX48ojhCLDsfmu7r3gMBO+xiX
+uDnz16NvUl1gBKGsFyEPCnEfep8Vo/PqLA7tZaLB0ChZQVACf9NZ0JNDesENbJDYs513jDX1lfV
dUMNkm52YUWzf1Zw6ddpc5r9qXjmfNqNNW+VRRWBMK0J0cZyg5yK0dYR5ZVgxjK6dNwDO9DoTvFN
iBm+qkAbCLblc70WVf/uDSb11JWmgTFGmcWnCpQOYkLBfLIKaaXfk6zkhooHU1aubtaI9bRvmHJz
JV7dlRQ8SPndJG0GWKJzkxpHqbEkhrJ/ZuJ1k+bpzqZDDir+4lRo8jyJ9Tac5UH7K1z6XlFCMGqC
6KgbkFJYX2S/pjno4ceYB0hhfJj0dYnqRc4ToDZ4wfcswCAiOgl9D8iLV9++7rsQ8whD0PbfJrQi
YZFjUIhC58FnRiQtSLaazXWTpRMBolpO6MqXAGdmhEGp06eI5l48GeN8kO+kQp9WBbyxV70Ng1OI
v7dAa3SpyO65KZja6nFlKINh9pYgN5xMgwZ7TZq8r6Xv9lL3aCOu7bstPdUvPQpXBj0rpCWLIWac
gu8fkJ81pVWIzzWmSXypV5uGmz73V6nrg22kMgbrMGlRPVz8ZqC1Z1xtn5NJDXFnXXq2bOqea+hb
dL4Tf74vW4ZPkNkF1DtUsb0N6ssNBKmIOjGQjbDyuG49PbrD1AIBlj9CAL0vQD7ktT6erbIjKNPK
SJmUntkOikMQAMSHtSWrlDNSiDOf62XwI6UAREHFDF/oy/ZJsh6zpIV4i7A0LPsSuFWtIKiiVQvj
G0+kOk3yctETLITJtgFBGEfYnnhfynYfMDC7QXux5jkiTyKkiP1RWxUVFbdicApu8HZW64drhXhQ
s9toZ5WLOMt5lXgvQVSeAGbRS83pHamM1rfkjxxKBaCpuKSKVJ2cO/95OjkF1vDS5h0ZOfylKpBb
GpH+0kfd55rvcN0DrkZ+4SgZbTsRga6wWCefqrIixQTtFWzi39SudSkPY+CsqaaELKxxSr91PKOq
n0P9a4HTxqkIESwH6y6Lwm3zZz/SAmuOP7OnAZXHL5Bx2lqPPsISlPSUS9rLIh78wqQNNBqopRZT
2IzRLrf9eZgPhUH3yEwr7D+gYzsE+PLhDFXqnKpapDeS8ZSdfy0gxZxhmPiCeZz6eQkmnfnsau5x
/UdM2Gloyo2JuCRNKlwqmmSc+UkUmSowlhLMRZ2hjtCrKjfW1u/PHaRWyQbxP+0J+yJqI5NOL+bJ
F0CjwSgQxP4JnSW0ynfj6y65zJIStIPLx3H9RXjO5zMJDq+/s/nwUD9/ctxLeImlOBoTSyneiaRY
bufPl4eEYooJRdgelQwjh4TeMaiDYofCvubGwqCN5Sldl5ZyYW/LjbKm3bOMnlpMh4l15SM+y4yo
S+o0+iIiwHU24JRAq/VOupuM+gAviCfW+KexQTrLVCFIq1hOxAb9wC0/sYH6h+erOrIDE5+qP8DS
79OVLbhyvTWw3aeJ6VG/ai/Y1GL/c17KxgVlgN2xDu7yw4HwtjrpYdCrUHFARPUiMqnGqFrSe7vO
sL2W4dYGA3snqc+G7mivnvniIZ3eitKdsj3tFzHbqw1uiGM7O7CgvxpXF0A2jC+4sPNZgtnRybx4
C6F6kOCUmRAccWWu4ubph9wcty95m8L7Bq1Q/fNQA8yET9kwFazWO1NTx8P8NpCfruVI2WbV11iX
qhBxlhG2iTzn8ao1nz/aAnmkira6Vgpx154g5GCt7V54PcNIXiQYpZfDT6U/+6dvJzSo/EiogO2P
bPdUCD/qE5sYopFi7TEZitMuMvIP/Jt9c1+Hqb1WI65dd4l03hAlA6HgDIfKiZ5r4+DnjXrhMjNL
BTQfTLh/HNqL8/isUSz3JIB+8OT7BcVlNORCJ2lwRiWOT96zuUnKGE1qIqZU3E+47XHWmGyw+VjB
9RtFnSTtrOEa1bUk9ZSrz+/b3J4VI78rfWzyCDNPtNftd2keFUzV9ofoFbT4BgNG4mPc1cOYugks
98PXNBYNgfx5Y16K+6FhxNMjeUkQYNYADz7iDTVhRABH3bWdcStv8EwkuqahAcv7mDe8isVeQwc5
8IsDG+jWQ9OpIifuLgekIHl3mbnqrskhcuZu6IiuIE5C3Ao749JM70hO5fSUmFE+rdl5mi9ij30u
1vJj3x/Afhy9sKNlynabsiUTxL+djj6MFoNf50dp2o4B8FLDrg/mCQaovER+33g6P8nNdhZsdny9
juAdo6x4IgwL4WajiRsrCmApqrzc6CeOP857qB1Bnl/0RenHBjgNRfpY2Ut7GXpw8YF2nJ7HDxwO
DlQmz+p5e+4fiLGIExNKfUR9aVE1wjj3fPsftggLFNwENNdRf/PVLrRBRZC8sTYfDLbEDbjljDLB
SdCmWUGQjHrhD6FGveMZoKxsxoShW0gcwU8tBjq/PhXRqD7zVUKxnBxygJ3p65StUo5g9QVxgr2O
nhun1n9XHQ0NFnf8PyZ2PSV++rc2oJko0w6fjLvlrFgdKVDTAj46oKxHfrLbwiAYyF7gt2BWMD/+
NXgO1JM0jqdWdEQylh8hNLXGvStZlJi3yBLBdHj/8ewI8o+uMfm4IRqwRrBeymq6e9bPyo9rYuzb
DGowzilW/6EqxOYPdam+AQ1GCNtulFtqoSt4MW3lqlst4Xlnexh8I+SPMdDaxL9zro/MPDOOwqc4
6k7B7039TCzPHYQgDSMOiLON8Y3fDTqFfh+Is2/WTaXt+ENwXCl7+B2YpU3Ns087fc9b3s71y5Wa
OCeOoUWBuq+NF0omrKBRr6RPQx2fxFzbEplCLMbWwERAAC6iqd92cQ6LI7ymM4Ya8exfaOCzgC5O
bC700iEyfoShncNR0sPPwA967F/OlX40GzyDoXo4tfc5womGrBaYLUkN7bXUxVZD+kaM1iFFpQzc
m8kGWCNSmzYfgMEVg6Zs7QMYhR/pWl5VVGjsbpEWJ0Lx1nToeGdeVAvY/8a9ZdCD80qRPFe+NZMB
pTjAdXaFX8RHRJmWgogoh7pUpeE3xbO/Mmycsl8pK0Ev35Y2HoNPZI6jXUwkvldCVWmKWhvjpUry
hgpPIqQUb6utVq8MMoVMhNSGpS5xlZPJ5DtR2/MtpISTC62qC3fIutCNrFh8Ar1wzY8pdJSzpA6p
SZYX9sx4Pe9OCfRF3j40K9hszwVwSje8eZyHXBdHehsWWio7gN4hKVfAVM5dH/r9NTBVJa7wjksI
Cul3dmPCQ0UcUWfb5RNctusG0dLkgwfothpfRMO4tkdB+J20QdGWshSgGqMyeIbalN+fWh51al4B
LqHUkSxPn/Ik9K1o4zVvRMzur46Lo9gWbLyUacnSMiSNygbSeDkbmQqvpGS9Ycx2VAcukdbW4ETg
7VEiBk7LOHTXbfGbxJd1jrxlQEVcHbzJRR0hu3j7NPl6GKmOSxT/+tgOM5YTMaVubN4/BnNOuqdK
waEmv2fSP36ATtG4Uv4sbOuWuJA6oB9PwNJymp9nP4E3S6M4N6symcE8T6B5L8mOMhvrrzbA+DIx
WgVG9lFzo8lDmy05+a77/o5AJrCOqfgW+ZYzMghaeCS/FjxYW3sVIlZEcFBpthdZMDQEMideql5q
brjaV92dJ8a6h0rModB+sRxfaCORyBY95nNVoY/7rtN98KBE8gkuMxz3dnUSe+9TS3k1DtngQuoF
TMZbVNDy4o41aYruAthuQ6DRb85PZiPiFYSbrnV9Uq7p+HMiCCBEOpPlshKMBCNgLkyOR10F+sUf
+xNy8Uuky5nBo9ZJLBHUySmeSwDiM1nicSfN3qCR33bbH6TF6piucHKYkC84y4gDo28Ulsq5kDDx
X+NAnfdp+IhipGfUKnC2bZS+HMJDsIWkFsr+eAFIuh/W/kkK7t/4tMypw1cBTPIIHLibg+BzwVL3
o7F9MJHAGUGqewErhfpncYheyMY7+ZuohuPM08MHQDWAtw3snINpMsGE0zh9vIoMofOWHOCoPI9f
5u4gVY+llDrIuN7Dwdf0U75yFMoP5tMI4wAWaRJGkFX6XbHScYL8yHpDPMfeQM8IOegytIPD3+8D
mL5nPKC61qzIVVw0x9JT8oO+mB7mvcxLWtoWQQaADg2Ek2mc/hOFcTiCeAeqbXBVtJc6q3V66wBO
ZmSRB6BhZkmd4lso1KXVzN9vwAMFidMndiiCwhtCisrR1t51wzcM80xsLMaatQBM5QH/NhxoB19y
De6VjqOok/C/W1ZdDxfLok8TKFjVGtYZ40K1kATQ/nBbehl9PHPXAFoczLU0Ft/CNGbe019UMGZu
9l/MMIzlpyr/Lcr9/mKfCv+ybBqgJNGbKwfW4oSjgVnnv4ud/zLKItRp1DJO1Jz7UoG+0MvvpO/F
DmojLEmJQPrzXUgaVUyRQ6DzuGBAL2hvLoPURFzByWoN/U01xhcHRMYjldYIDWidrIVn4truL/Ej
596U6XuyLbKjxKhK2cz6g7xjZNnWuDUXYeOy8SHTxIa8lnM28z146sbVLVRbkVPbyeZIJ7eXKRkR
1h2GpsJRODBhQzTecSEw5rt76YNnO/Xrws7xX/Levxbn4x1ApyYluUlgeVtQKUf7QFMDzcxP5jtM
aZsQKGevgzRtaGKwZ1tp47nxYw+2zMZSkOD6zGjaCK2lxsY6wrdVP8zhKodDkpYkl68hBR+9Y6Ee
A3aX+CzxQrdJvkuGogrdc9/ENQ/si5AB37r8Balnh+qD7Jb0Ln1FJnD+iy0wM4ieB/h7C9F8gwnS
K/6a+co1IYSqxpyTy2sElE7vuCKRIlpVWNJV8riTn6mhIhTDAl5nfSMrRRTON1xWQ0SDkM/rt6YY
OwIfstroVvrBUBq+qPgpYAkfb0awbSf6B7uDitxPOyKHOyx37ZujuzVFAuxTUokRMt1ThxYZV8Kx
t7HJIk7+E1PsIkkQaNyj81yAA9eVmn1itkQcjjW9+hNYdX6adGN2TarJx0bPu5qM0fLzEwtPYyDS
eVyNAAfDNzthc96FaekrtgE7PCDcqKH327Yg/lR3Y5lT2KQECJi89jBp7Q+LWVIKoZ5e8l3NxTGE
mjnMYB7gA1Tyq2zOMbtbirY221BsIFMiuhTNz+1I+MLrG72nGs2esXDMfb66F+TeHKoStOKVvJMk
A2ssdIkuqYMdhQL4smKrXUmxpzDsR/cNiN1Dvn4RUn6OwkIO0na3wibe5fezHzrf2qH95sRwrA4P
ZaO8P0CVtQdP6qZk9f22tgC6HfO3Ngx1YilBf2rbg7ZQM6I5fbnPwAWbVwi8aEwAKJ0pb2VX/2K2
b/2Ru/Q7IpivzN+oxaogR+rvJ0KhBGtLyYf6EUQ3kOJNH2gK0nmFYQs1PELWmqtPC99M0DXUgAVM
wj7C+k9Ti0N9/O3GL2SCYKQJ0KYc8PizKvQXpbNCMp9HfGF17ldJ9NUlIZ2tlWKtk42Wf/7M6/CD
LtcBVRmGXB6Ogk4CjvPZ8GuAQGqPWeRlBKh7DCc0pCUzMHkSiq+5BLVnw+7AkpDr3LXFEDbbhvzG
yziXHtJzDPWNU1HnfP0I3deeCwrHrwkpwRoRzuFiizQfDONo+ohC6f0tC3qAtoZJQmE+DrDJiVtj
/jgYazJk1O60U6BnO0eWsz851+aHOyy8vUv6darAyNq337AyXYGh363ZDlU/2q24+ILjEto1Sydi
Ou/7rUceR71gPtcD/o5XiE9L6KmOMAsl6WGNLDNL8sPCjo7BWMdRwhHt0xwj0U1OyeFGCIG7ZfAD
w20WPC+0o6NXCFWFpQ+8vRG8mSiRX+blUBifdazTGWjsAJWwPy6u85OYzXa4sz23VImWtlYAHQlS
IUjgt1Iru4RbIXvEnJAoClB0dRRRFeYxHJ8Pbv+AnIUyRERzYdMI7vv0ys2SpvdcXY3h6vXFxPO/
XRdGobVSpJZrzHtlE9BmSaeWlH2eKNYwyexZ0zWF6INXTqcMBsSi3gzem3rnZFcB4OwNYTBBBpLW
0W+cUNCc2EaFRibbXQGe9odsC3MerdqcaqVqiNxS2yQzhO+pDEYRJZDDjSDj18A1P50V/VxwlPkj
7j5CfLhKHSRlE0lcAFSSyeRmT7REYWBwe9gCwMQv8JwNhd4tpBhTs2w/6jVgkY0hj+BYRzmE2CGm
HmHuwZPkjMZVYjHkuQ6DY7n8i2juglu3tYRri/VRNasdGMV88kPZpLWf1AmpMIUi4CbGiIqlFAlj
pD7x7W5EsgPzL90HkNn0Q3R6KnFsCO7a1eXdpz/4P2VH5ybNUEjx5yAqwxA1p49KQEaNjoYbXwoH
a0FsW9IeS+Ys2TWxvWREgRh51cHkoIv3ej0dNrRytwhaXe6rMqfqvhqkJ/alDCHfzcFCWiJCuDfY
u45zEbnqGUVhPfGPhEF40DTK+OZyuxfdHuQ1msipEGa8Z/4/OcOkUPSc29skChop8q30WgEuxymD
uUr8tLnojyvmsqk+Up/pOJL7/hii2ZeEaa+D+4a2j+0XjFZRIiLh4pdr+bHa/xaEU9bqQNQXWELk
Df+c9RJNvYijqKobsI41lLaLbSSNSIGZb9WnjzG/dbNGbTMEYPorDMn4pjuz7HgacKJ86wQN6U5G
bhWUp7DDPf9oRtUyqy7TbnNQ865jAIH/jeRK27HYcLreaNFy9VHsDhSHuWcB1vValWVArnm+hwRU
NrRcoASZLE2XroDEp0TdWAR2JybymtH5pH1SYjcYR/Y/vIPxoFCNPjV+nH6OIJp75GiytovT6JY3
iUEx1pvbakq2hbqmlzTjCzNVanr6KSO3HgwjDA4gO3GKPcctr8UYgFadGboHZopQtUkHL0wIBzum
VqXKossN3VBL7ntLSBR8XV9LsquFAU0XPdBpHKzIqoRN00PWUJD4cdO4xn7hAwWRF/jBV5lQlTRx
xkahnLNuY64vIcvmCu7WD2tvJLTd0fdDNKFsh9fVlCRFwQBVwoXKHS3jY3X25/R1N2HHRrtfmEyo
b+XsW+hWIEMOwVtECD4ocwH5LBXTxTDY+0bVeVAez3D7zOQdxkw7JYjJfXGNQvc/gWs0CYBC6fC4
ZA/s+16PzRRfMGXk5iFhZIK1+XOjRlQgEiBHWgiDbQoIhKBNJqF2j0tOsaU+wdftdW2qoD7RbH7m
sjwkpGOMgvP9VNiKFYPmy51Mt8BImtg5WnYpc2arvrkXu+NTkaxgQXl6MrV79vDb4gZpmf26bHdc
qSUG1XorjlHTrvfU/JTSS3JblHCBWk/v9xyJIk46U6TKPIynuLIEJzF+TlnBqBqWVoC/VLxV4uff
12UlGHkDFtetg5FybAHgjYTzjW9duJiKD2m7HnA7+S5Iab7agmfkrga1+fJHHeNl+dRYFuVaDzeM
Zfu69DQt76yxDYbAVKIXmc0t53+CR0s+DFasYFbC5oFh3f5+9az1qmPL/bt5WVRPAfNnw8IpzdsV
t9PpOpygLwxhGcSmRS/GpqPpCiEHccqM6aC7XslJgGGz1QOGTEkg9MHl45NYvotjQV/1TVh5wk3K
2T2oMN+TngRYEBabSe+t9qW7iolngi2cGZ9EFHwdlGDGRrPwqCc4ZM9uAQFlJQFlyku7HGrGGoLU
wEqlU0o9paaTauxMqhCbMN/IKetIrTTYvBxozywuhC9/uC/CK+jZ8E55TlkpScrTMmR4m9PNe6Og
WLrOlqWk3LNCR1yyCqJ4GJFLP7c5OaQa86V49lpEcI0N+VxggnbDd2/460uwbJRuU0/JSTDOz4gg
sisPkblMZxNRndodf6t2XtKIhuRBLgC5VGGlIQ1iI4DF8xyazUwRLIBjJwQFY0eZmQqydfwD6Fwv
nNoZjsBMGTNcpWsCK1lPJGlnLklhqwnG/NEJTGsuu3EVwjsqHjD75YDkpM/i1OO7ubz7UX0WlWWM
e7yaQL5vT9j3sELTnawb+TSkkr+n8sB9+ZmdSsAuF+JGuuyPdVXV/kqVilocC2hdEEmIZDFSs/t2
yVhO5qhlEpoci9KhWguc1tC6obAbJdg1/2Bg0ax16L1iu/BvX66L9TO84QhUrYyaJ04fnELC51fH
w8cdkoytnDqbW0271MWb+kl3sLJEjilJt6prRDP03w+er0gP9NrEdTVUkMkL7LYCwQMPSuMyYRLm
Z6dlbyrLmV0M7erESsJPDkGOKjRj18pcD58ZHOy1DnCk1q4gYpfZerlGLGSxlbD0iPxIuGARXhEp
b+Po/eR18nLRJhcU5bQsoblHqHaPepW2hfwqexFT+J7gZgLX3N4wDYgX7xHoz8Rm42abWVC4kdPX
9my1pQatFWr1hk0+GXmYl1106nZbehHEKa3G7lBF4uVE1hcxqsfGrajcGL9SbQGcv1nlv9g9z+6y
HMNzp2vq+RaXlOfbTyQOX9LRFtst8hCyA8ehwUUkaXXVcKLk05ikqbbaGjyBC5ivsd4J9HrR5nqP
qQ7wQ6IOkJxG41wHXPDcJ5Spbndx+alvioTb0EK9Dka6nhs3mgXcTzHXjpHlVFSuT2IgNbuXIah9
O9VwI0Tvsps2iXEk/UXJqJLeiTgcZX7A7xcarMIxARhPlA6pCYIM8OKGdJ0M3tsBHLNBhPrtyn+f
NoC3wVcWLSeZ1ETC4Nv7/gQT0QeWaBRCaL2rh7ut5GCFvOiDBLfFlZ6yW25UuIaTq+eU5T/b+i68
FUEDs6jS3VhkMzBfCHceaviEmllY7dwYCZwGwiGUEEzJVGbYqDTVQRJo/Q4AFFdSqNxRi9bpSlOK
/zJtSAsCrbDcI95pK2+ELCHvH2Tpr5KHdkAmB0yshdbB7iLTcZZ+8sSh1m40mUEt7aTu/1XSh6rv
jMcRQ4J+fsdWXqhm+7EzHl/ud7zUdYgHKJSBiv4+S0kdL/WK6x3wgtzjM+HkheNfMyuAg2Rgt7Nf
DCXlWSIgpaOmv6J+roBFwoNAztCmf6ctbc6HFRwKiJdWzmSAtMJQ6GEsHVpZaF7G4BXnM8do/tqe
AoxucBgLF4X6Kz4OKRkyLNjwld0qgEGvfEtxZdz/DwExMp2XOfQzvIbY5cO8jfGfHRDROepacxLE
hQS/QwzmcN4eimKQ2mJxBZwsn35VvfjdLGJfk7OpnkWlEboM4IrT5Y1mKIXzfgJVFiZ/sajwBlvP
V9+9sxPjVhfflS0CCfirE2NNk9D6UUX7a4QVBKlK3Un4QuzMjIrfxwBazY75NchbkXgcStkCxUvI
6k3bXmNnyE4ajZm4/Sa+T+IsqB7QVN9lV29gj5Ozc3OKH/HRJwFLKNyALh4lIFpLLTfd0BoJzF5k
KODyvlzHQfD1tEoEkCm/4IxRtUKNG4cxSKKGND5x82Zrseex8Oc1LFaiN1VmOGfHb2S0O4Djjy/x
qXAIy0ENXvMHCIuAm9aGasuX5moPK2XEag4Ypy4t2SZd1lW1jULA3uj0UEw73is+MaOCol47k73V
S37zBUCS9inHA/lYjtQORvuzezPMj5L108EtpLv002vlEbMBY8QCQ9tTN6d4dM/eq8+dhb52nT29
fWf3sLDYhO15ard01Tvia9WSlA3nDfeu705jMVD/devPXOZbCos9If9zqaqaxYok3eZFBHGJPtvh
RaNCJKkyetK5w+l2ZxmHgedP249sS/thEMO3Zdvt/Kn1MWcXMtcFL5xTs1xa3Ee2i/qO2O8OoZ6i
H37WK6ubwf0HskYsCnn4UZn1lHXXtuPpeYfrLptj/1oAUQ5gorkKUzBWtqozZZ1vjhkb/29ojwv0
53KTxiJJmYTZvRr/E/0VRcwdx54G33gFRBtYPdR7JPwlUl+Od8nMbyfmf1t2fS2Ll9Uh03qLAM+F
YFLFC9z5CP1PiX5inQYEM8kHPV2jKoia3BkjpWUJB95qvoEaT9dy4wd5/7/1M4gcTOa1oEDu17V6
5y6Tcxzl60YZZa0zQEkn1v0CQCcuUdWxhNOUIBgMseyLgPXJL5ZBnWIyKJioT0viG3w9+sGtwKxI
jrY9XQjStfNXNHzNE8gijjAYSLhFN78OBWeZz0P0RvINjHdZjSOeiLYh1+V+PYWbfr59QeSNM9S+
kFr/Citgv8hiuwofrQMcs28jThzek06FGz142VTOQgpAOm+Xd1a+FgKoy7fWAUt1PLHinTwkBtyw
ug79Aw8NA3N82ghP5kJekNgS0mB74I6doeDfmjxM7tnu1H10vqSMXhTSA2rDq28JY7XIlVKKPbZW
O0tfjNKzogYLaM6w/h/xVPg7i7csrCgXvkn23i0Ax2N2/jHnx/SJh6BdBd9UBKL5wlUjp4HQh6+M
abpZmgtgV3LDjCgQW5UMhAknWp/5XAknuSfxYfRuqdS/9UtQ9qsaLYQxnqK5zMO9il4SILLwQ7qT
waG6izfa1V8qKHCedxkJm0VfYtDKpEducrpUXkpCILmmzSIgtpvnyP7m0wpuDwYrcw6HuQ4Ohutb
2QJiN3nN26BTR3Q5D9VYk53s339KH/J2WWXLUTZVMfMCBTpru2E0FkgToeP6iqDX1fBk8ceb3vjP
tJSDqkhnHcEphbTZyC6KfO053cJZK133oX3xY7HgDNecPSy10sV95rUkIn28qe/2XFs2Gy264kL8
qkC4pNZdadfJf1E18D8DM1tvwxmwLHUBtXI9akgmWPmr5c3noH4GQdoRwp3soWBG3O+XP1uLcQmq
xiFagw8DbodU/BI6HNOxxd87HqnppcEhWKgqdvjIj4UQzTPQzQEXzKBJUm9ux3QYE4ABmJSCKyQP
hDCPG3M10Q84nxfDqAHtodPvaloJ1VAdHZfTGZd5nsrr8exP799AIsejxZYdsTP/LCM7tz8u5ech
Rpo3vqgR8PMLiaAZrcK2oVQNa6P4bmAHPhy04+iOsai6AozK7R2LsZzk38vUEYcpNxsDw//NdPBM
x6XKAELOOEUVGr6V73IfVTu6g5l/l5WB9VxrZS+ZsGQmdJbDsZUtW5G9ms3qHeahhV1qWmIBdExE
Ox7/q1XcYDkTsfRG2+WvfIsNbe2HnFRq4SA3v1lbqfA9VdNE95AqkMKAw9UVwEDg5uO3T29U8EBz
Jt/S9AdkoUIyIV9UlLOcIqu29NCLOsPYt8fOmGwiGc8+ETuBuGDTWkr8nFytMki26AYkNTNeZcjl
xu7R/Hq4yiLHk5qp0eNlAng3sQGdh5hgjhlupOP2nblfHn5nw3MG3oP6Li7ZQO/wZUdD81Qifr1L
QY+AqeUB2zqy+sd4Yb7XjqSfmoLctSOZVOzpQJYKhxcHPSl97wVyc6IyPda5yg+dIPrLbpl1SeZ/
qgKhPWjJnJS4Khv7E/hjig+Z/5aNTUzTXhANrFrKCD1rl/KiOiQcN9YzxBraVm7O3vW8bG62Oq6C
NtZz2lFmBgGyUoEXTFnvezwXDbYLT1PtwVuNJ6MTkKU56FpdaE/d49BwfBC4lBaQ/umO5YME74dW
j7iVP07N4wPqnQ9ANv5zAve2Fv0deGfgjuI40rtSkLzL6w/RxDqbSyYb9gdh/W7V/Ya5aZpqmAa2
XtwLMcztD97lXC5r4UXCSVXiLG6WoputspHJIim8MQDpHqpuVcbgYPVgCcKVyQ2HC73pVno44zv2
6ceN0PGqQkajLwrsEu2btAa/QCbOWCIIdfjOd1lfgtlXw9TMFCVk9v9xB3lenaMdxWJRnp/2Qlgv
k2LXpTFe3uHkc0Mc5J6Tb5cJUUhM+BIgpzgIlRy16BDOekecsvrrV+m1WCL5OttLJawrFDbg/Ozw
0DWewaZvfRGRE0/bCn0bdKjMxDkT9gol6aZuaKT6/v66aeYM7cgFcJRLuh6j8N8k9SuR3zreGIJD
PRJDjCUCG2di1QnncPIABlGka5jKo8fAkjV8JnzqYvZnLRSOyDtN44L1IKysXwHAtc6g41wRm07Y
cowPXgvQCIeVGZk9HLhU2SROjvdTCnUyIUxaswq7QYa6GO542X1HcLPD4SCoXrGSYJ/XEM2I/Nup
9J39MxyNjwgIZrLbbbKwoG9kc6/tYLAiL+ybti2tRVvlGG1zVWOJLTpDNhDgnETSYdxpCkF5Fehr
ofqocIqZHzaNVtzcSKnIDRaCpPQQDbKXHJ9dAdn+lPcOAO+ffNSLOIePdGg2ZJjZjO8fQLFir0mS
onEBxiP8qEO4gbwp3Ch+oQldmZa2BmYG5lYV0U2lqfguXimraXApzXJCLDF0O0d1jRO07S4pWKgm
cQC1vzSJUrr2oT6g6I0TUzCHvPvo45ErQemudPK7oeJPm2KbPCJ/mxaEG0nE+9hMxAWoK3G1ImDs
8pxzFUDFg4SHERW5h7MkJjOQbEv8Nl8zSIQLWt+rUj8cKI9AtpXw4B6Gh9KVaTPGmJzq/C6ENtCc
4eG5RlRfbo4o1VDqMS7uPOg+E+XWW2hoHfq1WzrwGcGTvN3MDK5tkgs+Px4y0om0jVit+W0dS8IV
w+JYio22UZyvL8jz2kbH4MSvGM/WKudF2DqRG077IpjlxzSSzgrKMGPdNW4tbkO7SznJfPU/k13M
UX1wt9OudadZcHJHwslMlxtMc5o10HoZdE3Rpq/tKUaUijolY3wrPak7utbcZHXaz934DEgcdd3N
g1yOmjTGqdpfgcj0tYZT6ujxEIjPcC5HacNJIAcbxGBW3DUX4MqWF9poAiKzrT9E0VTd6cx7dfOT
8vnzC9RCvlfbK5Wukar017T0Xf6g/uG/GaOCLvq64X6mZA+RN1850tSLgiAJJxo5sCDNkVhUTfGu
OD+XJqanJc4rAZLScHoRRSSSTFI71zV2o1s5vXkn2wvtO08fb6mig5YyjDPo4Vp9OU/rkk0aGpoG
wiTKZqvR44Km9zFqWokFcVEte8LkB5SHMQiXVv6v/20diChl7jWd4QV6IEuZW9ecJ7FtJxUstg+4
obSNVaS1flZ8q7aVW90sLw01CXo/Rr8C4Y+q35hOx78wqCFNoaV8fdV/VV3YnCdR7mS3M4MKZCIZ
ON9ngjYq9kRPNHqfIiWtNK/lIRulUa4QVcq3ik590nfCYyLJxCtApLRJuUTqZiz5tz1OBk2q1QoK
gZC9mC3U4iESUPxmdYL5i76mR/Jpy6ngjhJ2R+Qpm7SGQzuQgYfNZOeC9ppqeZ/ecKzwBXiELS2r
kktTpXWvmHlxy0s3w3jhqCb6efjYWR/xbb1lYXBgQwwgsfe6PsXCSKpoRljDuKWceBn3660P3F6n
ji6r8oiC3Sw8H+lw3EHrZZt/FAdkwPZ+R1okF3pZn6T9aT7UFJyIwtk3OuYTRvJI4ET7m9A2Yro2
VrFF3tJspENkw7itC2x2kGB+Uy6MY8ZFlKwXqWPksHw2rvI3qkpTfSsERrwlQzgyS3QXTSGZKRPL
cIBbaIFMi0fUV0yBldfVR3Pllk56UC7OW0PbcMPX5A8JtodZndPCQqE1pIc+aEWKlp1unEAClYp3
jmc1oBZYWWkgxSXUcbE4fYGxLXukTj/+Y7tvWPU+cKK2o1WjZ2CdjioH3Dot4BHJFDW175VLt2O5
q7z5tVUc/O8nmYkLDrYqBb20ZcOIMcFX+PsTV38W7HfzstQLRC1IE8/i9wHeRiaOkvLuYaAHbzQd
MAlAkYQrpd4US17Zz5J+fofsCANhMlMv8JpoPfTo/hy9M78R8i2hzBiExJktlj1wde+sU/VJ17uH
BRXnhTh/Qd0DTRktAQsTPZamP+50mHUIoMLznEaNVGvHVp9hrTtJw7mdrjHC4EWLf0NxcAHhTUyh
/cyYElk5TQZe+uBA3bTAqO5VzZjWe/uH8RfOSsc7cCxOWDO4tSZQkyM+xCupfVVlIBkjhy2iVd/6
3p2DsyaLQZXaf8MPb+y4grR2RwdKqzsusFvffmtmrb9JfeB4LtFSJgvz81g0iMJS1mwAh+OKIVuq
sAyVnVTTK87PF6FuoQIMb7oHOAl+CwJvHUI5KhomjsC5kk/HZSakHer4IKvaRWRip4qZaaF98onH
yj1GMBHtPZiXH24YNfB+ar9Ry5b8yh/otV9FC17XHAz0DNs3T+8zUlx7jNO34nzdNtbvIzv6o/0d
iSM3JVMjMy3tRGfSFsjWk7evsXdd6tiN3QbobF3sXn3vHzmx31vc0ds6N81fJzW/pWtFwMKb44RS
qiJkDhAuYjPlKy3VenYHT9EY5TBPxgmdU6FPDmo62/jl0NnltIP4EPhqaJkQyUJS96x3oMV7Y2yF
JE6k3HSzFsXwDzFtJ4e7BS/mCrWwFfdUgx3msRhUCFcMoHbFQVeMbr/Haf1yzpuTTamNDuBBfOyT
nNWti3xQGxzt0QAWcVacHgnWL097qQq8g+14Dykcg7vgC4x+KOghmMaIlKThRvzWg+dULj7DhdV1
FAVA76aMMt5PYi7Oe0CXQ8+oBHUyYZ060WpSFd3YfNknBgu3fRLbN6e/2pzcxXdL5cPAQthtChLV
3bNvscTfuY+KHkY3e53RYtxdGMSO+cM/N7QA2RclQN5TCNHRrzasRC8xp3K1++Wq0gJoF/ILXkDs
tdUCFs51qxSxLRrhQ83CiJAom6+VQYhX5RHt2+71G/yEePYiCqNrc3CSJ6EOfqa/928Nwzql79pq
eBPE+vQUiZ2mbC20LJ/gXCVhH6JCzz/5sAlQ16/BAxSiAATGHnryR4PPBnLVkxI6TiGdFKfh8gbE
pvpN9nbIuY5/ziGR4hEgiQWEuu9JrnKMmH/DGGnje46rya0Y/FsWQYgTar8vMv/Q4nuae2BZ1zMt
n0ubbuKYn/Oj7MS9gbqpl5SpcrwtH3nLtcdrtN3bqzFFO3owR9D4m6kqlMMwUcoampEK60SSovEs
AVCHWd3go0QN34fAJ41S8EjEkCpqpEOkfBSemdYGZzI2epnLyCAufGg1wCXwFvNUgd2qCv8uNzYB
oTFeaKuuqN15refqEzUxqtd64y1en/X3MUE+zmrUGMAe7WZOogZb0s+4IOBIrWPi5qtehv2YyFTp
Geq/rcszC+Bf9DrtGbXSaUJ0tlbmC71gz8PbrJ/vQDgE7RTvGtHfoagwoQQwf9F+52tOqKI/qLMn
0P0rnW/lYvwVa+uJ66nrtSDnEAFdEgCzXJOZKqrW6jPz/XOnQRF53xWNjooZpM6DR3K0+bfuAnWR
LRhPvMRmqAXp0WzWWwlcBmcGVwxygAP6868SE3N6ZOniPPM4z9xZpaSNFJxNYz+ZqSYhOI8Nw/bO
5cQW6eOMapiCJgkfTxsv3Qz+rMaFf8yOXF2KIw/pPr0CKne8Od7DTIHVm+/RF3aOS1vdbwkpGo4p
VuctgxTaAvURu6gKscp9IufT5R48myeoduXjQ0l/qaOmL13udB+ZmxTtNloBDIxBzP9DcEk0SWTN
6u3OFhdx0+zMDPlHAO7L6/TPUGoZvnZSkk4LAqOZRAcGb7804XWo6u9YKRQgDNVCCkGrrQIueyvo
x6r9rfSj5V7quMi0f8Da14/14oIOZGNZja/i0Yg5p1+zYo2W/MuCbffUVkCNesTiRyEO2Oo/xKQF
nS2X8o3bloMIMPXpKttDmH5zWWT/BxazjyayGvnbKlF4fc2mEqw64fqanSF7YfbTaBQyEvYbiIc0
39Q09Zfso5HOGQJLze6WrsRR+O6gvogxvNFcJrbSdooVp0ylds6aqbmF+82bo//zT3XB/U6wX/GO
7dgw+v5OvjF5CDXU6L3H7cfaTa813s0LO9oefwjDaY1yMRF9MiSsnHDtQ0SvJorLAvhYvg2CLlE7
cWjMYUcj8v/0sXSvDzQzD3663W1SEy5hnZ4Egfk/pWAfo74vo6nC7f+gd9//v3Rv43e/KaovXazm
QHCFHawTeZefBKCsnpC9npN+oKS0fCBuAKnBg2ynjtWTkHHqI159sAe0eVoaYP5B5Ni9vUhMQ5X/
5x02NCD9Gjh9noPlU1R74Fjsz1aL6zSfhYnzcncHnoXfE12TyqA1KP/dYY8kS8YQsWyb/8oUWCO3
mjAD868zfKWlGeHfs87LJQU+7zuND6CquicQ7ULjhMlTHxNljECOhYJrKKYLxb+WU8xlLgcN8s/T
SOBcMJ3Nc/l1q/trLnQ9/T6k8i0mbximtJnK9ZvtAvRhaOm736Gb4H+0rbif+5lUopvkbXkvZdlr
10vbqls2VexWi8XzlFFz1AmeZgT3m/D/sl8Qa0Tz665qY4PwOXi0Fbu6wBOem0ONBcfr72uuwYU8
i556zNp3ZPRUoeSbte9ODSR4aqUcXd6llKuxpH8CAuk5qX9HJ+fb8ILz9IvHLsPfjLPRYUfzhH4H
5fpqHAF0QdjNEPGwLi39vQUQCyGIn/+OQs5xNe/UiyYK4A2U9aHOPeeEKO09FS8Wb83hsnm7C1oe
p6O8GtayWpwaO9t0bFPAs69801kWJfx4Uzv/ht71jd2VXOMQ8gT/1q7KRvOA4+iDuNGcfB3WXlsb
bFKiFN8yUO0SkJtE3qtWjDj9rSmWWaXE5MKmYridE6LkFVhWWIN9fLsYoY5laGD3vjYZu9dpWjV6
usMVGd0lII4PsgJxBSWNUyDz2BQo0dLS2v3RnB4NRBiV7jm2u4XyvPeSscZZuR0h8VkvpeoJEars
o4YVwLKZP8awFinLQy7ulnGZyBPcw7cK/a272v2jZ/WDcKWZiXekeq1o/3U+HcbQuj8nDNzC7QW4
4OZf7+spPCvbjymUao/YS7yAPKMjOaVUdDtaYQlTUuhCogboA407OQLoh02LvqD0GB4gc9S8c0iN
RPrxJjfKGszMBDFIMlmSU5xoYAL2UjhDfIpREiPHILvekH5oYnn25YpFIaPKviVwIjqSWBpuj+Kf
kdwOstFUVbN1GHfTyAXDVKHnsOxGAoAMnqIKRU+YzkvzHi1cPpnQIS4i0m53cE3g9cE83eilNfTI
RP39h69UaiQBwuoBYRbyc4REOksGqvAt/aXqmyMNPOwIEPgpzZPQTgz2CXGeAj5TQB5n0GLabs/n
C5IRE/V+pGzFG02f9OERfBaVCZlFHAoeRjAS4fI70VjZFo2dBLdH+9aeuz+UbWScC41sboMMflS/
odvSq0eVWN/8ElBV9zZR4KCNj8iQG1RzzJGZlYkkU3/ZAz/FHBtQYIg2Wsh2kzJvkVQFQh71yK/E
qbRcnxCz2OiPTkT9TP4doxoi7THHbnkxjm/D/fSHxmvK1ukTyWSsb1KN4MxZKlskEPwya7FIWDHv
Rse1Mb2FksXOf8iN2/M2+o0TZyzohutSyoTRX68EGeZOWMj/1VycUCeDUJgpuSCSofhnfhn47+6U
g7dvbF0qG93fZeZQN28tc0ANXBLJ4KI7pAfHLUTZuaZMiG2z9O+3KT55JQ7hlTvzobJ96jrRoTwU
HwQL0VoqmcJFsc9pPxRPYZH5aQVkbnz23OGp5EkzEqWmX2l9zOpMg18ecCs79g3AJx6SksIAH0XZ
zaIoGIgfWiQ2qcGrCTx/dNGCwGDzCjGNlTmk0967/iW0FXJsgG5l9igIm6pCbiASdLjOSXUgi2Py
vSRZ/rv5Ok8iSJRbJ2ZkrJpFDAKFFovKEEeVvU1oee4++MNXlamEQe0DFnckePita82eD1BhiNAR
MFftTZN7qfQW4S5RCFvTzuKy6uXqGOCTpdN1+GSuBlka6oDiL89Z5+OcZHfDi+4SrDWfogwIX/Ib
+WLTsVDTDSz8N/ovniPHw8iNRgcFlmTHtiTBGB1QDCcN4pPZJUTouLuD066h2cQ5oOSDVb1Qg3vt
So5ez7yLxzPWbb4An+j4AVruyiF0Bvt+wb2jb0DSDJgTa145gpkJ+5jimg2hktApX9HAUpO/Geac
ZzyUJipPJF/dcFZxUwveJvpy4g3uef98J8vMDK2wraOH8uCHOla0RUUt0M/C8uWMiS45WpY/RM10
Z1JVs0Zpwt22bcCty4PkfBqTIh0mEjrR5Vy1I7WRVtOjvDJmV3tmbdVUCg0/yG7qSO4e4KJoq3vC
Zh7SNiZRs3LdalW0jNodTbQE8MiOLwkS9PbH4V5jLzA58az5pyYHo/NZNlV+4o6Y9tpZtudQw5ik
6sx+uwlyu20q9FW3Df6tkSLX5Lq5jThrBWcI9cF6FkICjQLCkmEaWsnC016sBmkblEiHnZ9YOD05
u5NY05X1gm9EyvHIb/38HgbllZpMElwkMYW86r7AKrvr44BB1s8Sih022bABi3lD1DEiXZNOMbgA
vmUBDmfSJVdHvdvccFXHdrtAGbMFx7wT4HFc4uViPtoBAfUyT5rxMBNsgC9ypXGI/lQ01zYexQ2A
l1oBI+Mhq6tIe62AAxWIbxyPUVXn6mPrPtCyLagd0g4B1WN9m+ysWrGz6axUni4OWONbUCs5jZ1w
ZH2fBEq1lbioDZW4RhGCNW2K8DKKneSE4oSzgB6qI+GacbzEWULlJ7071lvufB90CSmO+ENeMZwu
N0YCj3IcG8iRmM/pNXVEi27TeOtkDk4VV9WrmgGkM+JK9k+YZCZiRwCcaiULSJLyG6rgqWP57cPo
0aqG6IyT8haPpVqG+OFGlMOnka0eNvs60tvbg+0c2HaVB6KKaA6i6hO20t/wytxp70bkZ3NW9pA9
EuKNYkQnIjxAkleRMlbxhg+b4ABRwNXu3E1BFLvENd2qcgAJKN1EkgDOdvH4YVITz6UvLdQMILT1
GpxZbErf2nzRrs6aS67Br2PrIAc7wqSiHElUW2OUuWzHKUnhTZ4ETTCVdPQJ4cvpYxTqNFNaudJ2
nDrDCWEnn7PcZ8NTT/7iKBLvCxNtehGwssHporcpwBtKERvujVjdqc8hhref8w3Kt3LxwN8PQqqB
eS2vc+gpTopeXHW8neUyTr3K3ENE8YsqW7y40mH/xUZpTYfpf19geaWz9EtC9DMlMIPm90UCNLv+
6bfcRGFZDagU58qNo0L/qS2XSHS54KHl/PVvzezYDxfLubjg9L+zUZ2H52oFdsue4EK8BZvNPXgp
mlstg7/Vw+Uq0sEgwCflDw1BCXUzzi9gqUiFaf8195UBYg9XtUXX5YoKhNuZtOyw3TrP4DVB2evA
nBbLNWsgey1IjVEYkJYhaSNtq2UX2BbTkcJSg6JSJs9E0ba24vHFdGMdI1vGXIlrxi/Av3DWsuHJ
1P257Gu9hWrqWKBcuvCfKG/7av+BmF5nQ+aD3m5Utjv2aDr3/WkMxA23Esw8GBKaMN8wQ3Ppd+Ol
swSQiFixy+tgdJ4T/+pS0kb3uSvVNgHTVv4NrqNVkOsOIE3Uya1Ci52J1LXEK3rdXKIuw3Ern3xJ
q8l6wBCEMuE9i1gYKmuITKDHpfuHMdjFT+Hh9FwNa7WY6XXSUJDSwTZwUsZydHIzVAWhvAK7snmI
5Hs41axpz0UO82JgL7Hr4+Nntq01gsb6Iv54Dmh6FQTTWmwFyo/PUx6p5W6/JU6NohEO2hmCNDC3
hIqxP2RAZSN33m13N/bSshY5kB9fTJ6/N2dT7/U54T8mCpYn9bTtcJX7qAXrrW0aO3ee7hDRo1ik
y1WqY3gRuttz11R7zhTvYZb181L3kCPUTbFx3DoZoXK/NC3AsRMDbWaeseM+1API9Skx3ZXTdL+v
9sYzEL7xApcknS/FrICCXYrRAuztdFUBurUya5yNjB1bW9WSmqciounkxSOnnIGttHuK493ld7Oy
xd21rjk95sBMrLpOVScOE1lyEZ8qgswLii85MTf9x0bTU+0d+44SJVg6qiZyB1dPfgvHYNngZQDF
JMYP7sspFcPksRJxlZABj+xkIm5sx78grrrlBY3k/+J5GiGqNDFb3bp/etWbyu8vaQZyC6RluFwB
un0D3IFkSDiMDPco14f/MTU2pjAbmHpSgqlD241VtAKCdU6fVw8JBdHh+fCBJyKzIDXDrDPr3AAY
pXFoVoWfAZX9ZR70i3O2ALG2dOxMuQxn2IZS8X4R4xljqUg5xgg40Ru7bmnOTgXpe6yPp0HmWdVF
UyECXXV+B0/vLu1Lq3+hRWcRuj6XOT3ogRcB/Rq8CmAkz6vBJBgk//KmWy2nQo468EsnefcH41VB
Cl19YK9xWtfQhGMz61bB/KP8lzVGaJ4V7oUZPdNhiVC3kgiiAJH4UI529zKt7JykuhwRtU0LavgH
LGFweDom7pJk0L+z0G8iWzLpSB8IO8tPwU/1mhuL4bgi6b+yMP6LiIzQSl2WUAiD3m86Z91+rsvh
KsXOUNzazdvX2kdPVTRVSnaPM7vkjuT90qw3bTLjNewxciv3Reh1Jhr5gqZvpG4cO2bW/7Y2107V
+VhoVney8F56EdLqTOgwet8c8HWAGjyuHpkPLoi2TBwh3gRRXbh7ZgH1goyxCP55Bfd4KNMDyWvC
rV4nVVID6uAxlvuMGg9AHR/Kf+8+HKQJtiyewKhe0UEz5xG/qjNcArrKHPvY0fzXEr7joNRL+Gg9
wy/TO/zyzwR112BDC3Fd7xVU/cZ7qN2ITPuCkEVrZURzTeOnMzv4ev9/wh1kVeej/F9J7qW5pUFN
1AOeuijwf9RF91q8Kl/4HjhI9dqvCtXdZFmYpCo7Pu6yWGnIoz6DEsT8SPJth4pLoChBV6Mg83dy
/vtEzeogUEgMdKa6kKi6fvgu5jBDXv7+TIeM2z33VRipxcDD+p83s4lVREMsjV6uGvRlcs5qGzBk
gRfd8CWX3XUsfDHKWpHsK9vKmFBqIThUN0LofSMhUOgO770er2tc0omO3Skir2zZj34yUA+GjlR6
34kEughqthaptN9sFrCvUe8nBWd2FUkfdkFEBFIqVbcsndqdmkfnP6Pjkux/VlY2xf8K9m5segkN
txsTwGnIN54b6W2ZH0Y2cmmVbrV0u8jg1BmfuroLJjoa4aW+1rwAuId6TMUgpvkphPbpqUz9MD6I
BzmzJo3c2DdafjbFGuUo9L8zudp2UhAUXqg4TjyRXs20AFAN1B0rs3ECnEc8xhKE0CCHNLCo1X8K
waG4+8iwOYbz6/EYoDUJfYS7o5HotAi9JtrM0aou0ahoAKFpYOdNAktfIT3J0gei1SWZEEqTBips
DuAgYMAN0ahN9q/AIJC7EfdTXqkCNIZ4GIDul1s+gojV88Z8HzJuYzhVjYMaWatvpSbG0aM7BOhl
jRRMu8dwG5YzMXnQG98xEHvN0hy0O5U7oqvzf/fU7vCtDE39DRgNHQYzQeKxwqVzrsYVJXyTJsU6
zPKQnRBh+WNVBh3A+5cElIbulvXK1amzUswOwfnupUf0sS47iwfNsKS0Yk7V5Qxpi3sojrGikzZ6
nX5CIbGOqU/f4Ia5NB8M+FVVElh9tNLJJHP6u9rgxRizGZ4pjRMrz/BAXoltcPQXS4sfeTFcUAFL
r3UAYn1Y0QkD2e+e8xbBGydqWYpr28MykuVPF8GXqbtnj7K7v/dReI+jPklbdFwr4fHKIWeN/Vf+
UAEbaCv81Mf3YK+J7GIHYahO7Ft2VDKgY+56WwmalssQTOzTDn95okMxbIr+dW0/FiKQHxpE+Rro
3LQfQvPWvRRQDyOGbCkEDYd/WpBBUwBg/VH8uRIcPRohFddY8q/p6daKsYhGiM7WXaphPZuk2NdD
OieZhbLfkXTGXWzzebztV49+f2FesJxliIFkupt6USOOqqUiiutj1rVnCReHCWMx5JoNPnjSzuf8
jSQCrQeduM2h4xMN3ELmnoh0OqjyINAjJSM3Y0G2Rq9F9A2IET9RI0cXMOAThpeQWlZISSHpg2VW
pVEObYcozZ+mrvv8F9bk1hw57AWoy7rI/kdSnhorC0dDk83m9fXVeF8S/PjMH0eTXDFmxpxlWfpO
+GabRG9dmGuRIGVl3pz1amP8/OTVTJa40ou0vHxbvoko8u7abm7yLngWHMQPQPESFSU1cAjF798t
WkbrYoxTgNh/eu1SqiR1TLP3DmIp2KPH+KBAlMk3tP0mupWWxeb50q/Rrw48D7mrcxB0BJqs211l
Gn98nMqgyJb6X4AgM9FYTv0PcvRv7n/F6hIODGuDUvuvZwEsXH6f/AY1yglfg+Wj++maMIsrwN17
xyqXICWfnl6cugdk/xsCWgSEHyvaXimqOAXYDvlnQ38yFkgZkisxJCEcw8O9OxCG5gd7giiS3MfE
/nua4eXyey2dHqenHe40BYOoRZmhp/FZnRqkoPnDhD+Z8SzNnxYF0vbsYTaC/rCrkGxDEnL9OIIU
vbC9uyViXflQnLgWTpWEbnbjEdB3zKPlyWvNatKPmSsO/dU+RehjWY3CUewz7LhGGZC4ypVPMXaU
01Fgn9xxaMuCYcDqB+EqOVPPPIzIqphRihWsDsRDouQA70tBHPN5s41bpB2cwRX9aKAQucxk/dmN
RNobqOvpDg4Jz4p9H0H/8BDrJfudnoojPsuyL0UVmwwLP9vm/bVw/vFdTLpfVueBpzvhovy7Vm83
I9sjlGKHSdoqAlfV/Iui4W2acC9hNu4l+JTLWaqA8HcmAuJ0M/VhNqv5nFUmfs6Ob+gojG2CQsaR
ZMqNAgwbiYPvEbiwSkPSp0+C/Mr48Jhj+Yd7ym0/FyVNRIg/7UiHHL6mSEWtjjz9klu+WoCMkWsC
qvTiQ28aEvkeCqW6lKWkjS6jy23/5/buw9oFvD5TbCfh+KfX8ybsapqiwVDBW4kwMO7UeINHpgh3
cbmdIBB5wVXWZjJ6yNeVvP+Pz5kSVaJu3eEoC3+Rrlu70D77RAHLxDO40IuN6EqZaBBoPklN1+w1
GocDKcHjNliHlo6k7Yzc8wLYFMgWF6YVrWqYpH/bUXiMs8n7arDQpoPd9lGbKVhaa67CVHGSqbQz
Y+Y+5yh1i+vLBKBgdrgXR8dGmUub0dTmosAoUzCHTJjUfToyrbi/rmSQq2uVloM2IFClyiaPJTAS
cc6Zk1SgnKoauoWlYkzqB965bB4L9i7o3o2A3X/lO7ssD2CQKmt5T4A9zPEmOwwPtiWM6xLawBw7
wa/RdQrwm3bPKXmHUWMqUVAXDqfff5HSwAWlLQukeEtOexscHY3xbTRAsoHEHD8UgoiPh100Uu7K
RC3xcsL5UzoqdlXW5AM86TfbP97bZ5klqhHyzebY7aVVHd3YYCiHRP9f1SIsHAluaJUb5T8X8zWn
+INpWLNfGb5/JoPfn4xDh9AeP+mdZj2taTarZqc2MEbHV6x0P9asPY3zrygRdFOjf5TZg2GH3yZg
JYKs6VLx4EGe8mXMJ9i+FSgy2AgEt6gz/8JvoOiIq5D8AI80DyeOArKngDR9fGF5BMi8ytQypfed
7joCZbCmNXJWok6Wc1E8ylcwYV+tCVF4uExV+cpCG4ERGDEBiBQjRkag1GqLunWMPUd1sSxALv+/
Sv9Wz1nv8D5wMEywnls0j8ahOWILNmTO8cpUAo4qE6i4loqkfh57ExF9j1m5ZcPiY7Ko4NQQDmI/
EtMeuRjr+qNpG/BrhC1cLfaFAohXRrj0VfY7RaFyYXz/xTsZqq6ZU4896K0UYd3mSUNG093rY1DH
/0oxUFNXmfwChQryzq2ZiOWaed64IExQ9aJSMhRymSODwCVe9+cB7kNqgfBpYYHd2vV33kkesb+K
gkaUQYBf9USifGOk4KehZNTAy/LNzgDqp5Iktmc02cMWieqEA88Tepyki3urrumZ2NXQdXHk4suZ
zMT6zVQClGUMhVM1oFd7n5yC0Pj1WR9y/KCgnPKyvNROwINjw1XuOPGw81XAasr+qjke0dGoMMBV
gwvy8PFPbtx3fB/6TGyvupSrHrMP6QY9Df9INWGIBSXjDfnCT52anAm+VBSmCtablxGoUoPfAIFK
DQvASDLLoizdqrPD6y3XkRXdo/lvhOJym2SLG43BDOhTX8qUSl48+sztGtFQibfWQHdXTCUW5Vud
61Q8SewiumoVTwnFDHTqdtAa6ypvoOIffwp/MMdgiIuWTh6HIwQdVSNLbgEBLOX2uMEkCWtrCahh
UtVsM/tKYrPFEJNoSBmvvwU007EKc9gIHao06+2CApCAgISDMkpVpSK2/XHyY7dS3XuBq37BEy7D
5WV//iEmgfLDo7ZqWpbn6J1ZAR7KNRjvIYlTvhR1ebLnG2i8yzPMkW6NFXzHNmW4wrTdRt7+jUG1
gF2cEtKIwQKVQZAj6/nUt791TfkWp95n6CKNG2ktBFm8McmcB4JFURk5kPlpfS3dcIuQNtMfn4nQ
MwQw+TQnYHv4SvoBS4PxcxJ3cWNdCkz0rd5LoppA2ev/eIvGJzJiTd+n2SS7i5hpZDPDcrDTtgGH
UuFdSSihFj6VMG6hImE/QX/zxUR3F3D+vyEJwbqYKYx3n7XLtB7teTHiawWwNDkHK1Gru/qN7vwU
ru416tgrdespX45aFuvskpppYm+FEOShMMI0NG+10m6hg2S361fRCXQBN5bP+vS++I/kcIY0Zai3
ScDtGeFUIZbk0GKG9cpiEK5hxkMYYCp5AtHvVpxH0IevcC+ibq7FY6A00wZs1G3lEBQ6ReqOs2wm
9fFVuG65R3m2O9y5fNb+bt0GAtTM/S3aFIOqgo1zZJS2C6EkJyqCDtTxH058N2aFpz2CaZnbZJ0p
WL4PBV6YkVguhTMetAJM4nWI9zx3Eq91XYPplemIL7ohA8dFOuEb7weswDuYLWZYIlLY9NR82hQv
RSWelEv44i4l9hEJVuKQCQhoLCSiahmcVHpCy64JtlAJc7gD94kYNRKcCo82GZPFHSD/QmtnW6Zc
aE/1h3dMbNaEWzdIHhaCP3QJUG/0P9r3UoeJ8celw/WtMI4tr68nhzVBoLxAFeVMXQ/L93mR7xHm
wf2cwOEgCEMDYYtrZWEJGzl0j8zATWt7LKpHSj0eItr0ngagpRBJ+2frjVNd9UNcgWKa1E/llxJR
QHSQnG9PLZNcMwjLs6ucwDdElkEJiGRtoN7NnKSoOLu2Czpi7WfTB/A/3eEyRCeffVQhCPVtZt3f
PKDcFL382x8losWZqWVgKKuFtPoKq6Z3rqyur6fEzVIYDr0JEHMIptcZ4fBvi02L7ziSmDQ8aptq
rmPDETPuQvY/6btf7OTggJP/KYHsw5nsQGlG1lIbmf5Cgt+jytZRBEnBKC2jlg3RPc5djJI0BINz
oD9VbgstDrtWabg1S7uGM62JVoPf2zAhYMkMDqrKRJNyAzGatEoaCzayRZAL9hbjhtINsK81gXLH
jD4dxuw+gtQv0MGyawOVlqQrszAoISaIaI3rLYJJszCgwYMllzZujAHi2NuDpS9o+tclNwGSpkUS
TbNk1qlUEbwHQt3VpE9DBD7v3l+OQKnZuusbS5VraOVCpMvOgmfQADoCopTAVTu0/gJ64VPPFZKk
Zo526wwwJp3OEvNXPXzecOCMOYZan3rjKjwub1Njb3Ykk9OLcFrNdHRGOHXtnFGCUv1uS9jn8obW
IIvQGWk7NNAQbwH0jMSMDJZKABy0/yA6yOREHT1FYGEJzTFpZlKhHNCh9FD+JvIfU4t+kA/2Y66k
fRXtSJ6yWSX1NPumkFbB0/GAB0Rt+4XaFe1VgW5yNNEk6zat1th80HGjZAti4U1rrJkoJpszPX0C
pco1h1rN1AdB/e/X6JdLZSiW8RmM5f00nsAQ5UJNSb7J9A5r2g46BiUGBL+oC1nBtyltIFkUImzw
Zt0t/+sJaO1exT289Ue3vAEAB7rVICH5nGYiLCieg+ttiJGTtNdjUzbgRXLoSB8L/eUF22OcnQWy
AkEEfsiJLfhiTv3Z43TpkDvaRGo1QLdGZqd4brLL/+xOYGAk9swFH78PobKsGhzFx6uVCOk0Oa9/
+4H+qa1+mepRa1r5FSbpDM4B/JK5JHc7kjHU9symwKJ/Zg+hiXEKBZkn6XAiR5CwZVn66nXEsOx+
UIP4kr8h5lEg6VFze1rnLmSeKcq/E+tVL/Kz3uEGu11ANRzqow/oJmlMvkRP/Q0PhzdPMVde7yS+
kx6IVHsdA3CcB/pW3PVV43XqvI0io9ZvcvtFiSk7/cWop6oUilvrfiz3HFOqCW/ZgRAbuDV2ZM3X
D46EFmAxDpUGY7ra4e+xmGbWo3o6M4vlHFez798aCYULlXjlnCphFG2cgcukkOAf0esgKJYSzgx4
V1pF0nBTGcHKkoPlXkmBlxDkKefsnDtkYJ5w8ZV5dr5indNknVFywKxs7xieR8cGnjCMK88LIkTS
KADi99Qj8MV28eipTYPSiRtx1Yt7IExoWQGpjFHcT2Lu6ordt078ro4gaWdMAO2SGnuHrmZdZ4M0
oFtgl65dRvdaKzUf3YqfknhtrUVWFtFkWG7juTGSkF4V2UqIkga4bpHQjqKYZsMC8n8ManRKQ1Tf
A4cqHMRApkOjZGMT5e84hynxD4kqtj2A1yUcNE+RzscZ+ZsqZY16iQwCMWSMcJFem4iMrQuWJ9RK
TYsm+ai+FEh0Mc3yrfmNuXbgSA4Q092DknyfCpWLfcP62k3qRyoOaqQXSLs1KoMzl5YK/rhBsK0z
ZCM/cpNi46og5aAvsUGQ63EEeYJYqNHdbu0N3Lb4uUgDqwg0IvtdDNFWBGDKzxAniTF5Xxr2BtGA
aAyu/sseKe3cfRZoAQ7/f9hXkTQqobBsJ+u5ZyRrckgsnA40P7Vhp2pebyh34l6lj3Ok+ZSHFyIt
aEI1oYi83eyZgvSKgoMJGh3+YO5RWMZkVSGY5Fw68nXCHEwW+Ark5inH92IVKDwoF/RllJczAxMW
DfdUAciWilgmYSuuE1yZlPW0XeKlHpF8HHFkMXctTzCWXapMUZxffKVvGZI0CEE0aMzdHIMquNl3
VYylc08cfRObqR80ElHnBdnZqUkia7a9+g774/0YnGmZbd83UKZ700At4cHX1D/UYCdtklVxR/oV
tgXkOgiKOw0k5u63Z1PbJEjNZq/EqkbEJ4qPNY0RBKph4yP+LLEuulqShcywK/Ct5NQkdKur2wWK
By2An28UomX9dU04tVWSEzX50DnBIZUn8hsaaIOuRYwOmiDUcs5AIhEe1X0AhgfawUjn0MTdjf0V
Zd7m4Ye1OGJYfS8dREpH50iPAHjWuTbKHLBb2NldufcywOzb0LDLyM1+zs7OYC1DwUjiOp5Fg5bu
BimeRJZxXUFIeGEfN3rW6m+onOzO0XitDX9I1zSd93yRgIlEZbuEu4dmc/PpBH4BfntAVyomodnv
ClWuR3d8F2DLGb6/zHDon2i7yjnYse73Jd459034lpn+9fwRM2xGENqUdyqyeKKCH+QBN14OPPAX
FFcpGgwASRaULAwKoUljkAFWr4tjkkjq/SwMIxIvQQ9iZ+knXYEivks09tXAIEvhj4WWlHfV3NnJ
aYGX1HxB4T7iMNFsEe4s53JYH2lgiznJU4u5x0+hM0rxmnSgqx2Flnswq9q3h5WZCxN28enUdO3W
8ByPG99C15u2YX++puU06L0yJ2eP5HnwOZfC/TTNhtJ50HUiRxg8LdDzp5klAFW6TVR7KIYKDrYs
tcbj3rz/SoKezH7sof57r/RULNFiTBHQDvcB0zMAKof7bUQTb5AZZLH+azFWxK8usOagrKTVnr6G
63nQgvui4ETU88JRuEQan0rjuLdjcpP0crtErMNY69KUmNy7fjNegVt27KaHah3SB8zgT4wiF6MH
k5xRslplg4hwFGIyzCDowTaLWD0Tt3RjnHNWVGsDwbSQ2JTXkoLJ4I5+aC4sR03TjGhZ6A2GYgzd
c2UEBczKzOfOE6CcdtVh34LnRpAe23KZGjnz594vMOinSC2n/1/fXTwVNPdBqX+dV2WQPwFi13XI
IELHVQn+uq+Vo2aOWUzRgrYfn894uRT7vUKFThrXBtnCZulxDr/CS4d7LhsEJ3F8PZ4M79UG8jEv
kXNHuDryxFhVg5LJx5CXnJ5cAmMBrLCOhE/XDx77L5G706bIemQnF0rqlv9fPxqv/ZswVK4zP++N
ck+dZEYwmvnvcMlIL+DxKBjC+ZsQYegklhEqiH7B5e8m9nwrxtsb5IumZzwyORJzyplCRD4Ll4CI
zXHNCokbEzlmT6PCXu8HRUSa7zml7IAKhVeeoNfD+8znQr8nqBmPX98z3qEOpDbgAKvA9LuZ6Zog
ycfL3AfbXrVlSTRtx+TJr39VRxo3Sp12mj7ilD7hmKvk5ZlFkas+cTb8Ia6e6uFjckzg3zeCMPg+
jfVcQSQaD7lYEHS+kHOvOmGg3IMsIgwYzFPSC0A6y3AOUhyF24/bta5xgTp3S/Nkunmnw3gmIYyO
IKQeW1quShMXf8nA4bHDddnEO98LiV2my/JAbgWm2b86dDwRFdpez87RE6beilIck/44p66VlTmj
WV2892pnHc84WrHhswisP/IZLCTENStMu4Abq315nFWYGQCqRnEjAWq/zJDizL9v1OxCfw8O8aTk
MN1R/BcIbT4cy7WfMYWUfdEKScYD2dqxMfWYU0QorltPvXhBCr6vUEyrhDzYm8VDUVbEiMiJz9fi
wbl7scjOpY3FWcG9LWl1y6pE57Yn+fYW4HEFZ5txxUxSpyAaJznf5eU9EhwrUwdOLD0xtL7/SXFX
M5FC6ZrFNOBRCMxztywRaJqloGwEla8S28rleenVPWQ0qmcW9vlon3DGphHxtKBncMfyeCiB0Tiy
ENNQQnGY6RJ7nHLCEFxqsrddOQ3ZS9Uxf+ahgD5iybwcB/pKdo8AdaAE5CZFUGW+X2+3PPi7vrDC
7PZU46LZxVPohz5fGq/PlUowfnjpGMjSKif3p66Hi9xnUXORLtO6ThpNaWrdSn+FhzD3xbKeW51E
1G78CNLXbX8iXanC1nUnYM6dE2y/W2QYG+GEeeXFcLHMf6AsSE/yfF88xo3GQkqKhla0Ks7N7B2D
aZvLwFZpjSRnUXxBuGqtASbLFpMM1FdvSyMVI13fRKfBPYHAFPJCCVkqWlBvIrTcm5V2tiEWmhR6
50qWHC6oIY4o5HhxBsHQe4Kh3BBhSf5+17S9SKWmaHmRqSL5/zVapCAsEPBlMWMfLqpFcyx9vZuq
giXRy3gO8vXMIdFq6E0r3bruOgcM/QE/ozYUiRv06+yaQHdEwljndUgf0+Psp+Bq5BycdncUgREX
R66f5DnfzUSJWqJkQnTb3lEV0A56ScFvFiI1AdKY4nu91PGg1WEhl1KnElju/DD0KArNt17+5yyq
zw8leFBhClHGzJ5iVGREwVWOEBgaLskpPWJGLlEPTLG28UdsOKQznyVl6nmD4dIm09U2FPGwNh1l
oOIShqnpEVNkvcnu2ainHPfJyjwgiA68fQoNZnJN+I3Vo86Ja4/J/cAvkw2JAc8XTMUW5BSJbH0X
UWc3LI3tOB4ybanvUjj+B3+Fk3Q1cSp0D8A8SH9deZBpeUk3sPJiCEoJetr5v1MmHrsC4ABZ1jlP
DhNSmiWHbpre7vINfyM/Lo4CoVRON6slzognZYAe7V0K+epO7DOc0nEPDX9RBvRf34EuZdUUSsXu
wAaBb5+VPicbmVmWrHxhkVvHMZlI/E/+20O4SsGWeMUbXC2UzZVH8WMDR2uiIEFyI09ZBxI/zSD8
iLbaUpwO+mRv0TNCLlLwxC4LvRELqVnrMpi1mpMlygX6zGedheHRCtAG/nPBLtJGVu5PAnitvU/0
ylbZpNAb9y3TNaX5oqJy6NRrolLl+ibVY+QhV1DBG8/Ec88/kKVWseMCtsvw13nj37MZ/GF+6edl
dZs17GyhnGBAsxSJXzJc34mSYiUjNtKf4y9Ah+AERgvBOHR2uWSLQO1fCtkLJwiMWXLCQ4qa4Iq6
cvtsMU/OiFuMIVZEDc/fQoVBLf042ksWdD92jhuFqBg/uCZNfGfv/5lwMlru/KfO+tAxiXoCWg6y
dEufmZFNHLTj4E9suEAIWK0vcjbWWALrBa0JE7rDHzDN518mgpE0CAtBQbw8Z5C63m+6VJJJhwnZ
Yv1dgB3gGjr6CjuRFhvOT1UeDTyrwgDU7XWySjqlwRnKGzsmMJZ1buOGELVhRgCafEi5URPPIvd1
o+P6YKcw8LCCPPmDwtJeTkfSY5zGroxc8QbOZnHrgIvEMduK8rYNS6jpk6qPbR124Dz2zzK264bQ
fAKOOjCJZOvMP7zBwstKwmHL6fXm+IZ7yOpXpifmoxs6J3f86QOdTM6UrS91YSgH2hrJlClGEogc
cL2f40qb3bOmkzfOk8B+QIOtktJp1Q6xziLBdkWkjp5PHHfXG8mvRa+QUtgBAGbgjyqf/cRtGRZI
Zg0ZND9IuFEc8wbYRz4MwWlPBhDUHkoD1i4QoP1Cm6eK34tA7ouMMaxTcqDe7r+0Vl0u2tS+B93C
UkKhhoGXeYZivX/Wbt0qgfcYbTsTJcNjRpGJ93fbJ1lqytTPSELRdn4v1c5JCFkXApxeekFGz/Sm
6IAqCjJq/EcVEACki83rd02BAwKN2Nzaeqc7ILhxuVzhOHfbHG95m0UKfnKqF+M6QDgfWzGq7b+9
4o690w8H1vHEeTInUsMHtr5pWlIpdNJGdqtbaLrkEenc5+zBScT0crhuGqCA+Kqez8zhN4hVvBLs
1oFijkAsGOo3+ojpACsCHLWx9aDivRZTFzOsKuJji7XYaEkYw7Rg5Ldcx9mu6r1KSzK4j7AkpxZb
agohTgUASQ/kAMQM2JrjsWrEmrWNH2Mx2NzduCN73q4dU8XOcI8b119ScklqdM2TLBXw0Kfb3A3B
fqD4Fuz6XIZgRuurFruyPfyy+mIxDeLVotp975FwGo4ZtjKAw5van6lBKgllX3wl4k8BL0oio0lJ
ycSYk7JEAH/R0y2/auvo+n1vSnV2YDIEP56cTvPFASullTXagQPIBtJEza1vQthQ4ZgVv1xX35fS
ehWYulypZZ4IYm+QywFMNa0c7gBLU2Sb1EifjnliKPe0lhBjtBkIJHo+GeV16vt09n6g3dn+/5QT
e0DZxFDkUZSJqFOAfVtQSLXuwkgaNe/oKTWZfncnbzGQtbtD2iPSXrO6Yp645s7KpPPJ1EmzXwWu
8+LCxL+cv28c0jXQdqxFlHTOuL4P95fv3J+r4uNKAg5SfKXJCe/LzVYidMewQXqXDoEeNqenbCRD
J11yuzsBfS+D8JJz/rzjk/3v1PXA12Nj8AG8p9Li734hjBGjk6GJzMW2ZGJV8x4xrgTj5DPW4Gsc
Kj0rWnYxsHe5vy5Xdup1/1g90dsxnPXtB3Eq+s4Y5+TgbU63FuKUVYkhznaHDZMhWRsk07ttVkIg
7yPeV51EP3jgVs92g6wJUOL+St8FsphVbsMEFbVjPMnNsjWmJeNGLRLiAJvXoDso2pKXjckE33px
2JVUU73esRktgx/A7p2LpIgyZ+/rVjiJvHS8lnwXR01jexaFtd4OrlFNRUAQf5yUQbrAPHFUuGIX
TPP6dG/1rAuXXWDM8OqXHp/Opn1tcNZPIhVRb+TVlid0SYUU2tpK4ZlQQasGLJ65qQ5/M0zIQgYs
G59ZFIMDs79qKSz8GbypKSc+eE5K/Z2TlBAeqDr9nDmUVw57uNPSehhivcBOnRa9mjFjRAPhrpt/
vw8jj6PO6iNvsfA+cL7yqniKhan1Qxy/NQJ9xvis0we5+CwE0jK40r9N6SfhmN7e2wC0z1KTmZxo
dmH9MN0tTUAEIqvSGUwhYTExxVQYq9zvdiCIN0mXiA0l98vXaxf1GEyxrP/SeJsZDL9Ux3B/ZBmN
V+HgvXFnHRWsDaitZ9nJHl4S5pP4eak8EkFR9wL9PeJukLqnBmZ69FM2sAym/dTUa351rZh4bRU6
70QXu0ui9OVB18Mo3cDJ1Fy86wdsjERLS1DUyNBXdETU4Wc1dARvUDsmhagyayzJNKaDciD6nJyq
n0sFbvQBy7nZ1jrz+dcOetgx5s4WOgiHgWgYsJKyfG2LVL7S2CsmHZjchlgOrjGqNf9Pv5A/4/iD
n+n5ArEGdu85JRdLvqsBV6EA/paDPMNs5iP8xSk/3SflhtzU5vjrwqFWFhkYBaauFm0+e1IGNLNk
GaKTV45cqS9uWH3wxz5TPuVsonB3vVyDj6kGG9hMAVIGkS5Cksr3QQ7jilLpQkxuDyJZ2iXDK18r
vfAoFUaV417fjRdFZHEcoOL9vdnin5p4ubbYJjohYATyF0Q2QyAZS1B2651hakqoJsWxOwnbtCcM
HhRoKu6n23vN2YrHCPQsi0M7rT6ggX51lYXYkSdrewZIw0TTGSP4mIyghNUYBpOZu1KZqG7y7cKU
ZIrSfOR0XdTz0POKLnJoNyDmcAJUpgmFziCwQ//W45FurHEXbjjEwmpi1F4d0F3pWXmzb1dNgCWe
gntbkMHsNTIyda2zBL78WCEn3N0mbSRMtSGw7qEzhuTV4vnGAzdfuj+TDSE8t1cMaVudDvQKUrKz
2eRrCvRqThA1zv3gNBxCiv1f99rRRmxdfF61tX8+a3IMvTHonMTQnjXqGgaOq8amp0mPi8OaPhqC
nsNvT72Ec4XVKjrq+p0eMT9+33I+qaFaB8u/wK2FK7z/FnLtOSruVVD7WF+9oZhXFWpIpmYla0rL
X16h7iwrPcktace2EUGshnLEx63qtdJ74+RKCwbFlDhzj6y3gAtQkV3CEIRKaqcXvUk/EqPcV3VG
SlCb/0JmvgQDuxhvDdbh2P4Dau7S/GqM6JFABEwpLtIgrqoXWzcgJFTbBoToZpnbUda8VG9Cf/D2
gPGTD+PuHU06JLdI+YA4PWQ5o7AOfNaPYjwgX0ACWiql/vhY0U1cY7aR9MQ861ADBlsdx6An+6R8
Cv2/nTC0A+BJqxU39tIXTQCzXy3beUZBE0xhQ9PXMBPBq8V1FOa21/WhRV+mACQlJMgonOzg52Xg
VsSIA/4P+9ADlY/rsyiLdXP0zGRSv6AiafHWwz4ohaC8tnx5obFHwz9H/FnESJy9wv716KeCDD1+
mZnE/aO9ZmoXkFJv2+l9BHwPtnfVlhnnldmy37pVUifO6FydSUINltq3gaB6DfUy8YcK+9tyy9BC
KozOUUia1B15VX5MrDOKacF5QZygG7EACxsnXyi89VERo2yG3m+xgE1bxlAlLm7MNqOkM5wTN/G9
gtQSYFxG2oyKuk4fnBl3gULXJAc7g6TfAE028ZQqffjtLEiG0DNqKjxRRezu4atZvZA1zBWkKJD6
Hc858deOosHQLX9JsIHMeSc9R4jOYg2GzU9Nxqe5iUoxznRh9YD4UzJmt/NHWb0t7ixjzX6aROlY
TyiqafMM9bq/vJla70jMViGooExePW5RE2jbzx5Fuv1pg2Z3ccGB+e281mjqdPkzNscPOPzpwyTq
JfyXcDZLOP5T7W79zGAzIz4PBnjJpwf8Cd2Ziq7HV18cBEingfH/nxvVClPNEfMwbTEHTcELZnDI
nvS05+eQ4rdFCSieiwBaQOBDeGFLALWGjZNBL8agNSsLSHayM3bqK8a5gUbUYYCg0reYbWP/peCG
hEEJsynzfai2JoMuNl3fnc2sYMWWVT1W73NdnEWgEWZjnqq1j0jtYXGb8KjjZq/a2bTl5cfjrUpR
vuTp3k/rCZ2FZqFmw3mRJ4OGFVLGuYKNp1/fEdxl4lZkUKec117y0/mbb+BFkwILbFaQ8S4VkBoD
5a2B2jOU9KdW2KgzWHwHzTCFqAEQa+WKaYjBUIXgBTTySekahNlyZskavVsV6dPXwF34Yi9C7Xnh
vWNb67b/6J1/d+BbrM/Am7d/y0fv8ZOfL/F+bEob1jfJSZnf2gcdli5KC4cO/YIO10MQnxRNAG/u
GG2byUoEhwba6YbcDqFfnu2p8QAAszfdHNm6x+ITP1QU9SUru7Epdccw2ISL3JGVS6xrTdVJVm4p
1TLm+Jilz0U+g9z5frGjfX9uYsl6822CyZTCme1YKEByrDDK06k4lX7Z7RF2YZ8LT9LZ7gB7Q3Ol
P6pd2t/ae+nrO6vV6mTSlL9eHxgmlLW3Hl2N72Lo7q6RtuyX/la1q+rYGXKiq/9Dhv3yDEdHIP5g
+u7tBLC9l1jDQkunO/uo1DLc73t+p573J925cEaJMSEx+LMwMDWCsF9TUKJPo0Pqlgnz7nJ3a/Gh
AkRIDalofbdqkGj1HWHiLdbE4KA6yiBlPtKuGlHQRAlkB46MkD++wjGVfd7J6icKzPBoUfYup1no
05/GCTqrzXxepQHYYZAIo/P+VPsELXgdtDjDhozw29g4Lnz/WYbmKURt0VVDzXwD3QfbgwTk1twc
mPiUDPac4PJJMSOmWO5KVqeA3yuPC1dJ3fSRdDe2t9ldf5mJTaCU0yluIFlr4mTHmUfQBhp5I5TU
MmBIWuLMB8xCA4/9LJF8Yx0BvxlHbHWRPMbxUzDOEnE1Wd6x+IUj150/x6Fz1maRuvIXtiiFG1nS
BeuFqqobqo7dIbKyE8ClWiDBOXGuIYyYZ19O2VzvUselWLiB1gb/6sayiEfYwNAHCr4GNkah8H6C
agHgf2iyhwSrfSpRRBJfUTyokCUOF6goemyt0p5s5YCSrkXkQrTZqFDzFIfIWO3LpBxw0PwOsTTo
m9m0Sl9W/vT/oA3vHsCyGjyX3+TaEpa6gR40g7qubzS1Z4d2YNGd61s7RcgNQRC14cCSQGiuRs1r
M5ysDD3pUNfB7oviGV/tYAspVTWadDsGotCMgGKPHOsxEUKIIukmpCcIr2CdDh18eLzf8Uy9kMng
sR5A5fW+5GuNcCyZ4AHrGAgNO3MzN3LYYtsxGmyCDgtxpnWTy0hNr65tjVfTmsifyQtQa81k7SHu
K8QECzjWHYB8MfcEm40Np4AHmIuXG3aVrOebUF7rbBLW88/t5gUnXV/CKWgvXXgNj8ClLXXyECNf
0djiMblxTtuVtK/CpN7Nu0GIuAdYwiqI3sC9esMbDcvMHjqX/5S3yHsoBBTofbR41MWW8cBkPB25
AHJu3FnZDinmfTLP8aDh1sMV6vRmpWE/5i3AKDAga4SlSP7Rdb341De3X8kdDZtBFovCbf6i46cp
sM+9tddUDFTScrWjlDu+hQb4U48VKGbNk8LqtWozb+TCpYtzfzgLCZiavHC8grtgC6XSyeRH0ljh
yBmDSYr9LHEJUrp//TY9MCo29HEVBtPTo9elTMxEkpFYbNMY74ra9dHCxx3Rf0IFCknOQYtz3abe
03gOyZ6lBq515gSkqgPSQzFg6CoIWLDBsyku1ePdNmVeXZyIeoYoJwgkvldtx97/wauZICeyYNgp
YGIHPWTXVyGhCdNqS+H//43beVM5gAm6PC5hTAa0zsP6oyQYG0iOPJaXfuJFMSwzF8fKf85EParI
J6lSsQZZrVjtEfM/as8zla5rfkvBX21eypDqHSyMRqp6h0PQcy4AZIPj6tV34soMvlero+B989sL
n08yRdDfUNLJJNMiO7HEixTUnOfvwi12KPL2OTKLyamSaiYhrpTOV70CqmD5+a83CnJtjlu2bHDE
J8+l9Nw5l7bS8AePqIUHF5goPsbiQNVhxpcGN78VnISsYH9bCsRNCkxe706e9Ubdw2QKJPI1vkBj
VOv6ZSCc/UB++oUcnEfdWh6Y/OSb0bUWlafCXDAvEdQY+RQGhYFhyljW42F0PLVPlwuLbPuUbGbe
h5UvcNNoJFwmtjNgTjyo9J28HDXNA7X1NyeeWhC4mxKTZlY8gtzJIYj+TEYvO9/2j2Um1c7DkTva
G3Su0Jt99WgnIMkEGZ2ShrvLDHAOhDawiVBT1z8l3hbmqzPOpDnX+PJql2l17xGzYQTaDUdbrYpT
xMmaJe2KxcnZcUZTp7cVCQDVOSvdqB4/yEO5kqUaqu2TEQSbYBSBDBAjXAKAYnWZefPdtvNaKDbU
s9nLV6nUvk0aIXgQ5FBHrOptcaPIIBr1TYfnAjf4OhKUwdVn3KAvG2XOE0tfGRNwTAv52VkXRNFa
2D/Ib1rONT00F4Vry1SIZhLceoRxE3jiNkeQhLk1ztPNIUqvbA5OL/CRr9bjp4YKOTOZ409ZFtUL
RohM6sk1ZjgAsAnvi3CXuTmAHQoCD8s+1JSDqjNIkB0IzA1emSrGMdhBB6YyYK1SZ5McKd5hta5p
a497pyhWgFGs76vYtpzdLkSpQOuA6UzFcq4womkrPpfme+seUIr/DgQP3mZOu9fb9zRuzDdOKkl0
IMJUyaVuT/zyxamCNmDEUZc3sL14Ug1aFccrBk7+cBNYdhu/yp8Bo8HCs+43RX8YHswr42EGQ/IQ
Ja18lfwUhBOxs/dsyJeV+Od6mLBUiD9UoV/hxuyP9rvW3x5iUa1ZE+xg9twjz2J+jyLeTAh3m2Zp
dB3OwsFXAKPnU+Jw+tnE9GOV6fq9iUb7qCLjN9k+HlFH/pSrQ/S9wG4biAJk0fLyqCd2sGBdR0l5
EkRPyKI8rWJ278O36yXkk7pWYvA4DnKhsCmBm4SAgPHNznFUMYGyKtxYz/oOTGU5BNYw/O6pK6KH
we1UNu5QlJb+8WZ7OeHFNQkK9GCpNH0N3c7/V2fxiXLMbIl161/TpXtf+IIgyM5pRJedFNBIs5eT
kgj8ArIlkF1j2Fxwiwm/f9YK+TjYri2JLD0RG8z7ZNjzURRejZozhad9WLH+bjGgSgH1Z/k4eN5S
D6CdQe2B4uH1rTTZdHm0Cy/HbocMJ68GvAxJdaaoLs7zKRGPvzX91irFMD651hMQFt9xJo+YJtCG
l2uVXatI7ob8CX2ygbUav3cEBb9OITMKdIZs71/ehUZjy12qsS+lJohBSrzcEhKRQIPOCHG2bd0j
5W6PEevCZt/swRuJDrKJkMpM53ZdgRAW5O9Zxy7zFCaP3QsMJrAU3QaHVvlSDiLV/W0DRRAxWzOc
+lBsQRHTm6IqS/bVAO7LPXsF2SqHtHQUlYplQzifnlwp+6VCVByzKP0z/X7qYEjDBCj49CtpxlaE
5nPTf00Dtx7dMtP5s8febcJzebT5/OniHAdUwDyvlOT+fxOPKk3zIEa2tRlSAEavg90ysTVT6+hi
lxMCy4hPBs0YDa1mJAJUFhQnKHg2edVcT0lHdLj6oGCi8BGPafxTuZ8qSj3piNuZES6xacqfiBkd
LtQDcKKOW8yFNDbKDYh2NNdODqIG/wRSs3Ps6io7UmzJM30LXYeC+GRRFK2+2/dL3U93UzpEF++4
YtdNcwkLuVfofJtkH6i711ncl/jDiq9GbWwMLFM+/J3XUr2GmUJZ
`protect end_protected
