��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��[J���DV<���Y1?�s��A�.O��	b����F���0O��(XjX;�rf}�%�����(oq���7.k0-�HA��d���ox�q�P?!��^	9�\�44��_j㜰yo��P��H�$A��Bz�)��Z�s��Oa�,��o�l��FH�{����ZAF[�v����{^�p>����z��m�l�B:6�Fͳ	�,9}? �v�(�7(��I����[�!Mo�������8��Ik�y����D�h+�y�0������C�憪F��.��6�]{���\�fY	^�n��-��&5�Pj�^�%��5�\�(A�;�v�7���.�;\!'�_�.9}.��H�#I�NDP����Y�i-��R���U�[�Ya)5���~�zXH����)�JF�Ru@�����$��[�2\�dA�w�: 5	��������o����#3���qߕi
H[�xԲ����:R�#�	���	����Mh��s�n�]E�q�G�����[��+���_kn���@�ٗ%[,M8���}�����:��j@�p��Q�k���>���!��"FW���Q(Ueo���^�������Q숔�OM��g�DAx���;���4���K[��I6�q,Ô��"�0�DP�}�ሒ��b��?���cE\���#i�u�1x���&*y�̜K�.FČ�9)E���E[!���?k�{�� ��&`>��Ef��ph=�=1^�����t���P��=Z9��Y�j�v�N�A�|���-��'�Y7k��甔r+�!�j����4W&3�Q�d�8�>k5���Q����H�i(��t����ze��~���c���F\���y`jK-)s��毃��ŉdf��?Q��n&�Ǜ�#��O\�{���rG�j�X��"��>��NFxܓ(�^*t;��퀆$B�?W��{(:JI�n4�5<�� �UpV`lV���7�#�P'N#q���<B���f���me���Y9s�cL��,pF�r�b��7L��49��_�(ucWRՆT�}ѹ�\���PR��@0a��A�uF�s:�n$&1_������ye|�o���h�P�t�x���#�")a���$����,'�)��.���Ɏ\�꛶���ڂ+���ޤ�>�R*����6�ԋ8�_�r��L/[��&��LѦ8-_�������y�+�/�,�:�����I<��j�u���<p����T?c׀���S�7��K��w������I{=���!��c��8Qv<�����mI<\|�.�#�["�M�m^l2�x'�q���qJՔ�rv6�+*����1�=��b��Y�v����nL*^tc�Ԓ5\��:�/p�����i	�����Z�����̮�S?��b�ퟳ�A��e)���TJ#���/���էp�_`s=�<13b���v����V ��Z��3�̹���ۤW��hk#���t"�-D��n�S����a�`H~�\��d�`W?)#�Q/����^*0L�z9������*N��4�T#y���,\��a�P�N�*��Q�Y��i�ߛ��������!��m��CKN���E�Ѥ��楖:��!����q.#��.��S\�}��ު�O?�����>��*=����V�1;�r���<���_�.f�B�
*�Es�`"o����Q�	��E5�ɤ�����&�Kr/�el>�`'�������}yP�]���V��,!7E�B�o�yGa ��F�������U�����Nʻڽ_1 ���h����QW��y��̴UA8ld�
���[Xq���aܲ�gl�3�Fڃ�Œ.O�M����X�9�E;�ǐBIP_�ڝ^�H��p�z۵D\�[KOϩ˛��4�1/�W���)���0�����$�V����������pDօ�a<�3��G��+2kD��E�ݧ)����Z&�0,A�hx�p�F͕0A�	�e�Z�U��|h�ER�^�C���5F�ӗ��D��U%�t9�Z�R���*lÛ���>�2�����r�N'�B!�q�gL��ZA(�����|V��!��<�6Cӌ�@at�V�z0G]���Vh3R]�l�b��CI�39��r�m?�xQ6��x����5fxp�b�J��]�rD�n��:�(�O�z�� 0[ ��#�8s��t�O��c���u������ f��}��jL�V�x��`�$%d���o���KpXYь;MO([��s��׉��NS��j��E@; �DC�;��ᶞ���Y�z���U�H��[�[*ְǓ��'�Wv�ӯ�ɮ+�MJ��$y%"���4��Y7��J�����|�]?-�^QD������e	��g�aV�!Y��A�N��f�B��C�jX�c�%n�����Ì�gȁ.��zh���z�@�j�arx�]@�/f�')�)��k���dl΀�6)��7�>��L\D�Ef�k�� 1���v!�� Q��KͶ���ZO�t�REY
	l��xe�:f��2��e˴M�>by^�,%��䜻Kz!wd4���b�Q�L��X��@�
d�	��{|q���M��޴�]�M��>5ܵ5y4��u2�N����U�ިep���0c��޺!WI0�.O�V��9��w�C�ⶫ�|Qi�>��"8z���[
g-%�vrm�#[����K�Q��@ľ �1�Ŏ����i�7b+J��<~M�k4WzE��n�9�$�
�b��@$%���>�����z �@,�[o��al��[P�^�˵�y���&2f�܌!�Ns/�L歶W��`���];xZW�[pe�|>�����A�-��C��uߔ���C��ݖ�|�����7�0}j}���kű2\������}��L��.b
g�݂�WP�AR�ӣ�٧`8��,�d�?�l�v��PK�M�6'�>g�e
Ø-���t��?���s�HRo���e��P�+b�SD�p�y�x��n,���Q��p3$Z7}�T�Օ�U��@���B��U���&T���5��y������`��*~6�)����D{����������nyEr;��Y�0*ɝN���S�q��`�#A#H�O��b՞�3P�E� �Ѧ� W)6_��m"(F[O'�|fm��=�o����k
�gȍ�`2�`"�J����K��pcaB�K�<�n����pg�L3��b�[����%��cS�yr�m��~�5��
x�[WŶ�R?|�m|�FJ=}R4z��ar�mΪ^�#����0m<;��i��z��
�Q`���e��=q10Uv4!��mY�e>��ȣ�@m-ۃ�稐��y�˚�M�&-�R���0��ȧs��o��9����j7�̪��펜�5���B�����wXʕ��ǤB��I���҉s�����eT��;�&����v�2O���DY�,�"��0Hl`�T�����T�[nxt%�F��EpXMO�flQB�%�������E��H���MR(Q~ԍ������4z��g�7w`�+pU�H� �;fOn�$�B"l�\�����7���Θ�<�z�b8��Oc�ksK��d~�U/јz�0T����R�Ȱv�J�A��;%$��ʚE���Ã�Jm��'n+=�;����̼h��Ŋv�)t�����Zǰ�ٷ��*ɠ�k'������~HvC-DJ>�VM��UmM�~�n�v�w�j�>L�wL��ǿ:V����Ss�9#q|}��*�n���P�����8��gg\o3,�$j��G�,
ʙ�H��sv�C�вr`zĆ%����>�I�Q����3BA{���G����5@' �\n���xs��5�>�*�f�� ��R�L{	��i>PA%n� G�2^�PZ��W�����S9ab��gA�γ? ����H['�1����K��$��F�*g<X�PW��Q#}|=�9c�C���*�Ři�~}
ѓ����1�/�g�����h�`f�c�d�w��{��k��Rd�Wl���'��FK:����*~�E-��*��n�`���J�'��Z�d�V�5��|Ut�x�
�!̾�×��E6u7��N��%�%y<�΂�ح8�aB��h]���X�^;:0�z��#�A��/#G��������I��fC5�c`�YX	�B[z�	�ZL��E�ȁޅ�e�ҩu먍����s��Jt�4�N��O�T~��a�Lk���½,X<�"u�K*�J�Dd��ٿ���1H&���h�V���@��0����~q�6)�'Z��o��������j�0d�q?�����K�Go_EE��C�]�=���]_Q��ɰ�[B���N����g��HJ�ِ�u?���B&
l,�*�!7IT$C����>��1��)�b�����Ba7I��Lײ��.Ԇ޿(��UF��Z�k��B:�"��l�e���&�:fZ;lm��(.�zk��:ˮ8Ql�
e��3��[A�x�V>[�i�L�h��P�
�C���� �txن�'�0[v)�;������[�u�EX,e��o����g)�l��q��N�l�Q!�m������hqYs�r6���%-��s��_B��@s̶��_{3�/��:���~����gA�P��̂gk�dG-�Hur�J�ם�5��\��e~�KG�����q���7+�vmh�SMgn�J��xd�Z�w���H�t%l=L��>�_��X����c�o㨰w��,l�%w�th��{.�ٍfv�*��?��|}w��~��[�>ɣ��6����K�f5N!� <8�����ڞ�����s� A���6�6�ii�VO�
i!T�g�$�nq\`��d�E	��w��S��%I gm��|���-&���.C'�>�
��� Ⱦ`�{'e��+���	��9"c��>j�-:% [��O�yA[>��h��A���Ԭ�M�U��2mЀ�C�q]�/�sN���r�./~`�Sag�(�;�&�;��:dD)mc7#�����;޺9�yچ!�9)�4S�ON�{��PwE$�>�+�j��uFDR�Fh�[#���S�C`���ASf��ʖ,=��llĺ�*�ڶtᨾ��|&xMgOo!7SR� =Șs�ܣ��!�摾�w��mm_�_E����k���(|6+�JXB���~��t�?�� �=8!�c��8�oߵ��RW)��
I\�������1�T�|�� �[�a�Dd��_b	����zK!Tzz���B}ͺ�.	Ȅ"TL���J_��bq$}R9�2&� K��L^'��\e��x�a 9h/o�Jd����mI7������xߪ�����h�w�׿"�QM#�����wٿ^ڜk\�y+섢��ڕe���m]V�q�>�vwZًv��@ �(���+E�Dl�p�����[7o��4I��:�F#�U5��)�x�4ϒ��\��}�֢��;J�1 �j�ي�N4���("pX�OÏ��l����Rm�1�T�U:$Y]"��F����L�2<m��֚�$�z��-	O�x5o�s��Q}���Z�Y��\ou�N���C0��ŵ_�X�1��q�o,���f��j��O�j)����~�hP6��B�\���1ۤ��~��#�}�aRL������pH��!�"��Hn��g�\p+B����Է�>����¯Nm�ǔ�Ԕ�Gb|C����W�=B]X�,5�W�fn�����Œ�\�X����0�ʂ�ח٘�YE�X��;X�*�����ܾܣ3u�.o&;J�<�ǘwL�rP�K�ш��uZ��(�~�?8�z)+]N����i�Cʹ�f����?3�Е���,f��J��y��7�e����}����_�ǕBd}���N+���q7,S�yoh{ۄA���`�TP?tq�pMV,I�/	NQ��՛�ܓ^�?Jy��RL�t����qΩ���P�'b�1B;�6�pd�^��P�����B�KM%�M�0��g�笨�dn)�m����n�*q��`�#,?Il��}�v�$��J�k��&�uN��PtbՊ
T��<���Y�Ս,�)�;xm�_B�N��D2��1Z#_���.̑��;�2�-ȅ�G����d��_��{�3	(5��i�R��?�HТp��1�D'�ݪ���Ֆ�|��������|^`Իc	Ү����"̒:��پL��:�Q]��ܸ��N�>[���ٵI��cRL<iV��������.ԥ�W�sU�b�*��m<i����2J��v�:#�S���k�_�l�.TuO�j�c.�����Y��C�&O�a�':;�S+P;��"���S���b��:�n�l�6�qŢG�s1�<�����%<���	�[?��Ǜ�S���[��j���P4n�g[���
ݚ�b��}�(
�1�?@�����o^$��W��(�Rt�m�r�"���<�Hj�M��r;h;LȆ�����=�:��^Kly�K�ʪ�1̗^m��G J��H�G&���
�V��k��[�S֔ށ���q�ǩ.�X��Rm���
�g�<��(�tÃ���s{_�G��&�iS& �[;�5^���0�.��p��w����9+��D�.�{�))���P�]��ʳ��6ڂ�ŽT�R;2`�*�c���?��2v`#g ����R/�?��s���������UF�m$]�YV�S+�~��p�4���M�{*�(aI1 U)��[�ȨR���3>����s3��8�c��o��yK_@���D�RG�[R��r�eȁ�����.@�������6��Ġ:b!\4?���H��d����U��O�����>U��(�����q�{韲饥��Ҁ�>}�;?E̴���3y|Ѧ�n�/�૭�C�;=@_��+�X%�V��v�2�tja���Խ�u�E�s]�ku�6\��_l{e��c��(?iE� ��f@cj
E��72�Q砞=V4�8ĵ��S�F�v�� �D���ɨ�׉7˰�~b�2��I�l�
��Rl���~S�_�h�$�-C�9�KO4e��c�q��[���J�5mwW=��W֘	�+f6X����9{�ߤ �-a�����B��Ң�j��˖��֩�g�y�:Ln��|TWhk��F
`	�XrD^�*-Ġ�w���)��4 ���|�ZH�u��~B%7H��̢1M�Eޣ�_���UT�l�Yŏ�)��]LLxr�S����'{8�9����BA⪿�
�8�ɣ����Ј�F��g�0�9�%�z�F=Bӡ�r}hj0�G������u��r����Ya"+�n���	�τ;�uғA$�}��יBO�$��J`߹�!vB����Ӂ�)���(i�^C���e�\�V %���j��Mp��
Il���l�(X3�y� JOL@�AV�^M�z�Gn���N�VJ�����i��2�|��Z������X�det`���T��I�ӥ�4�]��.��%.�_Ӣ����Shf'�^_Vo�ŲZMuJ}V#�E����L�DY��_+ lK�ȫ�\�x07��on��ܹk�"�H�B�@�9k_�m�%.g����.Ypj��嶱��#�����.�Y����:XR�6�k�w�71����ˡ�Z�-���48�&�^A�3��![��.J���F.ӭ9���ԅ �
�7������;�@���'by(�ȫJx�Iyw ����کi�o\�=/�=ۮ0�Mj0�U���z���(�=���ʶh	�����'�)��*o�����v;∍Â��o��O�)r@|�'g���θ��E�-�_�O��p��/�=G��� *�?ΚRe���L_=FAD$�R�)��+���H�Z� �(�q�3���6M�sYD
W*���;���6]�&�
�]G�t��ӢE�U���<���`�;�f�q�kc�'��6G6�2�F�3���s�7ܣ���7p��&�nPm�u��z��^���n�ܫ��T�i���y:����a3���G�+�&d��f��ˈ��ԏ]�'��	<�i�,�;��ېS����=��e4rmK��i�I�C}Δ������
�3�OyؙBݚUF�խ���}@�o�F��p$xO6���Q��k5���_>_�������\BS�hM���/M}�XW*� �y���'�Z�7���0M8���E(��yf_�	e�(YΧ�L�(~�%���y�o���{	���0����x`O}QFk������ܗ~whk�R�|a��-��:�����@]��p����۳c�3��T��.�.�^�OWU)n�=��<�]H�S�f�� �;C#��/x�U� <�ք�>{O���Ԝ�J�eRdMi��+�7xW��I%]R��vC��v��??Xg�IV䵺g��2A�M�N$z����:J�#Q:!�W�����YBds�O���p� o�����m��4w�>�����Oj���[�#m7B�[➆�����}�%��AK����SHoK �j:8"�uD��r�?/A�m����&�W:	�c���3�j��7ۀ��9bz�J!5�=6Iw��-6|8S���O񈪰�xcz9���M�d��dmٞ#z�d#s�r�� Cg3�ǔ�����0jW�OC�Fcg'w��F�]�=��<O�`�]���g����$�jO�9��s�0v�l�A��N��4���;��q��ǅ��W�ٴW�Ҟ�=���8o���mR�Ĝ�٧	R��E�}�b��z�W�q��5|nN����?t;3BXw�|��""Ə*�2���x�,)ξ�K�|�r=u��f,���������
�"�RǓg���a�,]�F��'�!�څ�%BoNﶡr+4E��g��=���(��'��y���~�T$�hC�"���J�:�3����E=�����u	��^��Bb!)��ї����Q�Hu�`
����}Y���]�z$�bf�K��l�u��f�tX�*
��~)g�7��d{l��Q��r�����+>�B�$0 �T\.kp���8���5�.����YA��`�uH��|��d6���
�zX|Y%���2Z�*p�R��݊sK�U��3�g�)��+w�e4���(ڦ��,�I���%��2H5�c,��Sa�e*����Zj�H�����ڴ��9x,�y�w���j��6"JI�^�J���?�ʼP�	x�yj�;U>@�a'���V�젼E�-�M^�	�֒{�y{�W1��^��,�]������Q� 4���e�@Rh�S��zh<~Q��=@H/t0�N[��Fx!su�x��1:���µ��e�����_u�n�4|�Q���?�ZEO��i�G=�k�
�3�@n�É���I{�����3j�fbMl4^�W��gb�f�fs��_��<�� ��F���go��Sѐ�� �� �.��1���{+�@�̋�([�Pk�ql��(��ݽPk;]��.�*jN��{���"�'\�5~��Kk�+��!�;�Δr!�L��C�Q^���=�����Z�����	��f�
���6�ͳj�Q�jA*¡�2~.�~���O�e5��QOM+SU�ԁF��&�O2�U����s���r��4-��e��Y#GqB�ZG<�e�8��2�{�W�F5�*j�B�3b���K������@f	>[��:d�@�MB��3)�V��霢�T�B��'�@; '��U�I����%r ���� *2�Ƿ��,��.D��ٝ���*�S����T{�C��#a���z��A���Ї�Q�9B�G�4���.�������[`?����e����Q��i)� �\��l)�%8���E�/`4��r���7���ͱD[�����,���ތ�>�/�ĪȰ��U�p�?��h�C�R����X�;�~Č�v6[<W�+�v=|}�|�G����Њ�����ķ�"��{w� 7W��Y���j #�D���ud�"�T�-T7	��7N����t���Ր�7�Qɯu?fz����^C�X�5D��A:X4��V�X�o� 8W/МE�J���XL.�,��뒒Kǎ���{*t��Z��&nݍ� ��m0&ɬl�����DR^�S�}Qo�D�1�9� ��F����� ������L�߽�Z�>ٕ��J'N�"���3���w9��Xx��\�;i�*���
�+�0��E��cP��A�I9jM��Ŕk��҈��L�d�b�{�.�PQ��Yc�Y&XC+)��_ ��!�JI���6�\�غ��]�OmwH/Tj��_4����\��O���Bҭ�0�	-%4o�����$�kZ��MÌ�������T�O,�}M��;3Z ؒ[6�����)�M��HI�^T�k�A})z�MԇH�2T�e�%_�8�n�P�E)�>ͱ��%�=5�`P� f�l� l�f�|�o���ZL�|ɲE�̌�Ѫ'R�T3��<_��I)�"�o�ǦȚ���#�i��'��K�Y|̸���躭sɴ���D�$���\�4K��V�;ڎ��oZ��;er�nS֥��
��F���O1�/6��.p˺��8	g��ʑKsQE��yYR���mXx�D�?���P��L0������O5��^���n���oYs(R`�]LT8�D}��?##u /���H�"�7�,)A&�}�PzQ���1]S%�;��d9� �0�n��)Џ0u�f�M�g��)�U5�C� ��)�c�L��W�d���0�y�U������EO�*#ALݤ�]_k9\�u�	�:�A�²�AD�]�mX�GS�_��'bN�*���;�e�<�-��Yк�,'�~�P�Jj��� N��'�$JpٿQ���H:�+v϶��M��z��0�l�g�	�GY���/M�GS���,w�[r�įڥ*���D֮j�ߠ���#Ix׶�f$���d��Y�	�vVZ������H��y�m!#�k���a�X�5�pκ4&CD�K�]���	ncG킅XmTl�D҅,�'�+��<�������zl��pC�A��!}��9��7{��b��0�8�UV�QI �[��,�tۑ���� �VR��HQ����>"��UbF)���%Ia+ �2���p��z�Rȷ�Hk�X�'�{�F}���"���wZEs*����C*�_��2R:}�N��﮶����0��� n���TP	NA���j��K���^W��T��X	=������f � Ȗ�/��-T�e5��:*/p�̭͜(T=��]cv����E��ht!ړ�z��K�����,�z�⠗���!�Z���]e�ʳ�������'�Y���~���+�%���"�]�m�������Λũ�=���xݴ�gJ��(�2T4\���ϭ<i��mTe�}-������-�5�Ƭ?�Zd��]�������>�.�c�n335/�2�M,�������ܕR6y�4���qŤM\����������b�����6�f����.$#��^~ }י0È=\1JS��������Hh KX?��S�?��9�0��1 �Z:�b��	�˖#l�{5�.��+|�uĦ��C��D攼���B�^�9�`��Z�����nCp�0?�߬�X䛈N����]��R��X9߫%�0ƚ�@�LO��O׮�����D>h����Bڭ!��% �]����)a�_��w��h�dI^MI^�X��f����R��5��aˢ����=�YGUO�(+q�� ,t��t�I+e�s�j}[=z">t�C=Ϭ���8Æ�!8w�ɬ?�4bՁ�.S2��ѣ��l]
ר�TL|Qr���6L�j5�,�k�RU��ˏ��ܶ��q5��Ī �pb d�� l|�!zm�������Ob�0-�T���0f���T�Ĉ���`�E�)lg>���Ĭ,<�����\���g��a�d�6�#ˮ#0����dY;vŕs�*^�	
��wb�P����N����S���TS���#�>���PV����Ђ�g��	���J�:s�A�ލ�k��� {�P�1�E�[�����Yk���� �j�mP�����̤&���>�g���ܙ�4j-&eE�e]ԢA��桪E'Ģ��,H��^2j��{����4�J[X��"�
C��;���.:�sm68� ���8��FH�d���Uyf�$�(�"C�C�8����L)>�xZ{7"��े�h;���nV��Z��5���mK2�`�ں�3<�Y�<�bC{OH�ԓ�ؘ7�RF!��%�f:#�ID<9K��/�h3ռ��9��N�=��a��2�gf� YƄ��_;:C,J�Y2���r�h��ڼ ��)`����(��ҡF�u M�'N(��z��@�1U|[�Οc�)ʅÝd��/���xSS^���r���nb/v|��9b%XKF����Dt��H��d�F��P��NY�C�p&*et<?ٌ�O�f��E(���\�� U�"������筪�lR�I���ȍ'�0�ˇ�ܲ�f�Oe�жZ��y@�ãO�/��<�Py1m3*���fu�R�+e�㞒l�����-�[�f���'����9C\�]�)c>��l�-�T�A�	�H|��U5#^�r��� mƶ\�f`�� ���6/gr�Ӵr����z�s���!H�Q}$KZ�J��}�J?t����m���?z�];��A·J}��#����t7e�4�$2m�UQ48�W��$����H�$�������R�� >K�q��5L���QӞo�;�@���F�JZ�`�߶�}9yN��p����E�+���7@#��&��g���hd0����l*�5�<�!�N��H�qGOZrP����5ֲC�|��*�S])�GT�ecv�JZ쁊xנ�䕨���goѼ��v�^>c�9�-5 I��2���*�7���t֬�`n�3����*��$7�7Ω�qT�
8�y�)�9�t�[���eI�R��Z�k�j��3�*s,\#�V�DSR�]b/����E�����oϨ�x�V9WHC�ǭq�> �7��P�Xj���cDm࣡���de��~���,���@���ã��7֔� ����j
(c9��܂)d��N���;��P����Yc��5 �]����o��~��S| �����Wy38�ymO���J�i�U��Ss��!9�3�M瑋����&����k�����+��8XdΖ��mih����5�H�]kq0�7�������A]�k�RK]��W�9�t�I��:<�]�@�K�柄�"2G��?o}�|�{�Àl�:Us�'p�CFNo�9�h~���GB���%Z���˖f�x�O8Q`3��:�sL�1�D�	�k�eF(�����[��6cL���[�*��Pfr	m�E�H~h��k9��ѓ��^?�<ԛ�g��]�R�F9Q�U8��T�-�� x��L3JH�w>u�����dy�ol�Q�Lג�����4l��[����\~SǶ����$����m��Z4ׅ�s����97!wbr���Q��Fe%R m�e�jA_"��JG%�OiC�_*�=E�:�j���	u��
<�kG���/���y��j�@8/�9$��Z���h���I,���B?X��.�9����n�S*>�#���c�'�F��M�4���Y�����>ZC�c�hX��:xSM��U�n @6Qu(�^�[(�\;��zo+[%(ëqz�G�&�_�X��'M��u�àEd��l`�;t��6L�=L�=���7�(�`�0K�[�m܎�b{|'fϸ�n\���]���V�����Ե���l)ةP���C����s��t务���s��W�t��&q�E&���zeDS���El�!8��(G�x�Kٌ�%W���C�D�O(P2b��q$DNEq��{ZdH�=Yo}�2R9O�OT�(">a9�6@�[�m>@��p�(O�����E����	I)�J�$Y��	�j�*��it#,�9ff��V����&e�N��
`._9�7S6�A��r�,QD�)��)�*_!OJ�g�#����g����j���v���� 6�G��<��f�t�4x$sо�PP�l��Ϋ$�WsLg��r�GB	u�8����
��榅��	[�p\C�%Z��	H�K[͐�����A�v�g,Z�mֈJ{#�:\��i�}s�fl�T-�%[Vi��8,�:��p�!����υ߬
ƨ�u�	��<k8��n��3>K��;��=*F�ڸ{Ol�>G���+�ec�P�tR4�+?��PO@�a���b������+jHe�I���_A��hj�ZX��H�����J�iB�/Ke�d�MQ��eu�Z��*,ɚ?����B|lͪ�>�{�4$1��~���s�E��f4(mO`����U"�A���\���J��eި�m��q�%��~��S����&yߋZ��\g���ְ%�|c�����òpX�Q�S�G�+:�[v���Ν{�̢"7b��j�Q�k3�����^�V�&�C\��s4RYZ\Iͳٹ���@�=�<���:�<l;�Д���ĺ����s3<}�Z���1k�=$�^35�'��{���j�\e��g�I�&B���:~���A _'qKՖ�B�Že���[�(���<��l����p�Pp��PSj�<���`ks�<��_@��z�y�0�w5��W��W(��K�&���b{Xf�S�7�6������wp�� �f�hMl+�M���Bu�]��I�5Mڻd ��7&�D�w��P��O�^}�Af�#����V֎zU��0hj�޸�I�vg�%�r/B?���!^h<#���S�O���'U���yT}8��h~�49ze ���`����9NX
WR1�y.Ps�[��f~�13�K����x��i���%� -�b�hiwgϏtt���O�{,���d�B�7M��^�	�r2L��Y�6�$%S��������2z)H���!י���u�;O ?����ϔ�D���N5����0g	��:�v�����n�
�r@��G1��|� y����{4��. Ns���1�*�l���ާ(��	�f��� ���e��ʅ.�a��(�{*�c2"�	d3�K߰<�,�^	�tm����x9��]��"��Kf�]�ͥ��M|��8�������B����T���g᱖#j��Y���+�+�_ ��,��|$�V7X+�#��;�?Z�6�ENEΨP��E�������3��͎iY�T'�Vpr�dy8�Ly�@#�ȱ��lT���o9+8�[Py�wV���4��;�8A��A�b%ҝ��A�)~���4��
�IՐ�����
T����޼�)�r��Fd3�9�x�����J~J�`���P�LK��"Pn���ad�D�E�!%-L���|�:�wU9<�q:��aq2���泩��Vq��mϝ���oW˰c�)����G����d+��8�sp\��R��5�7b!r{��JhL�>=��9-4�4��c���G�oЮ���U���5��ժ����%�$���c��JC��s�	�]��Y�k�����ɱ9$kg@
Á����[� 3ō䘾�B�=s�D�D38~�������,�,�.�]��䆁ɡ�Q���=��-)Fi.$��6�cb��m�~�&�&����oc`#��Mcx����9�*a��l�j�$6����"����\M�ͨt�-���鋐ytL��<*�6ţ���6���و^�/,^y�pޜ��r�d��ҫ>�M����ꕠ�PA���P-����=�ǡ��S��ƥD�Hz���N��$|Of�$&����&�U��B��<����7��Ի]*�*.s���0�[7��p�����q(B.YƧdX]�GQazu�����U���N}�={�
ש�^���#ف��S�Nu�^�����2v�SO��&A6���܁��/��S�h�`�A��=&]]D��&���o���{�!`�� �5�7�{؋eFR�Sկ��P�D7���呬µE'� ���YK\"}�$ć�艋�pk;:�}q�5ܓ9�pD��>%ot$�_.�F���R�S܎MG�O�&.I��n3��""��/u�\��k�6�2%<j�q�?���Ax?g��R���~������	�m�6�H�`�>X���'�U?yG�+ȝ�n��΋�r��k{� }�Z�fjz�l4)��7e,X/��(�i�y��^s����ɉ���R��p,���R~�����H
ί)��}l�����Gsq�4�3`�t�:'��L�� ���Z*H���a\����m��׫��(�~��	(I��@��P�3)��ΣP?�yQ˫��^�4��|��P��I����5�`��|�bf�dQma8������:%���5��R����cj����m7�" ʔ�t� V�Ej}!#��5��Ѣ�#��O��n
�.�hV�gzHɯq,���7��a<T䢇��Y�+J"uf�-\D�au�H�EBZ=4$��j�yu�Ϛ�Z�F�QI�_�'wC0�^y�0�=��AMn�ZH���k��M�2L�E�/`��(�1t�u�'~8�"�K��>���8H�`!��&\�#]�/X8��|Θ�ڙ���ŀ����r�k#ݨZ�����f�E���eǏ��%2��*�Eu���{b{㸟8Li�Xl#ڙ�S��gZ�۝w�s{Trq�^}���SI�!s�PZ-�jj�N�����﷦vi�ѽ�VZ>��[��Ve#�Wx��4A�	�����ꭱp}�G tx���0�k B��e[�ÆNt�����J�}=�������PXo�g��y������UǰŇ ��CJMG���'�JX��Oh�P��ޘ��˼�>�ݴu%Ÿ?G)����xE(��l;�8NK@Xכ�T4L���T$s�����s�X����O^f�[��n�
�^z?��
�HY���h�Žc�}n|�l��e�lM��aW�n�Ȼ�����b,q~>�@�HJVj!ަ9�����!wJl��+�;u!��Q�����Z
� &V�pZ�A�RsT����)%TlAF0!"Ua��>�ԑt�K��hԦ� Ϫ;�C�'�B����`�:#oܫ��E�s��ޡC� 1|"	㍧�� �g�K���u�7׉�OW�k���ʿ�R�bJ	����x�5K���V��#&�6ɑ�'v~^��բ�TY��{��k)��Ł�4`ډ��\#�7?�7����{�8�\���%��ey!BpCl�$s��v�N4�5��8���w+^�hX^o)�y����%��葠�gJ����\)3�4>k�������i���y�"���B�x�o4�Ը��1Xk����y[K`���>�A�����5�k-#.�`@�sH0~�䉐{,��ʅ�\�Q�v���ޟ$?����J,]�Y�4�J���o�U��M����������\�f����Mr�B�f�A>�($?���y
I��E HT�p_~�)�+S�7�2�bk����4����dF떘�C�zWU�$���k���@�f����7n��� �HtA���	�դ�eE7�{=�s���f�^��h������F��Iy���W,E�OjѠ��'�}Ԛ�����g�9��_�)^WJ;���޿�F0�ic��c�M��D@p/��QN�e��<O��+���{��*�J N?K.�	�˭H�=��1�cc�I@��R���<����j�>s~�mڭ�� ��*�)�t]�� 	ʜ?�g@�W������X��ꣷ�ش��S�<��F�����ʍ�։Z�TZ�e�������ܕ��rWL���%��3C���Au�"ť�3�n��
Lp�I�����	�W�� ���,}��Bf�繙�"����J���te�����M8�)�� ]�0�9`$���u�ִ+b&.M$t��H���I,cTX*�0�i=|%�¬*������&xj�����y���2b�͒(� ��ۼ��V���=˵�
���Y���2D�Mۘ�X���%�jx�ӓ]r呤7\9�(��}�ى���cpp�;�p���i�l�:L�0�u�b׬���H�A��tasf�>$��TƸ�?��r����P/�+�Ė�(�욒=a�C�m��Q��n� r9n{j�r��W�sn���+�Uy8�q�"Z"�Yf����Q�~�'��V͋fT>'���j�Q�	�������`�[�ي�@�XI�|��$���NKH
m����� ߾S�p�n�(��ɚS�C˺��CP �J����HW��a�z�T��R�w�=�G�I�m޳�����[k���y�m94"��B,d]����{��g���?,P�R 涣�v�K6�*&�G���k{1ߌY{m�{��/���Z��+o�W��[�)��:�G��Ѩ�z�W�ꅭ��r�jZlӪ���r,�� ��U��X�&�H���sc��k3$�j+����i(-��|i�jk��s�V7�B�H���F��\*g��_���3g�����3����B�7y��B�����9�5�'�5x�XI�;��㨽�1x�!�v��Z��ە��#�����g���K�@�.�-��%C���|e)�l_����}j��e!�#�����H=Я�9W�$b�/ �^�[��p�\��S�YS��ԘV��&O�Z���l��@���{M�h���C�^�ղ�p�f�W����b�%���_[A��� M-��'L�L���:ߴ��Fr��p�2��Q� օ���S�n�����ė���^eӒ�..}�F�#�}C7�k�?�ū^ J��%�9z�Zό|�U2 ӣK0G��jڣ&������� �#����v��x�@@LG��3�K�ʺ�O���bf
}!�[9X7�i�$�%��`���ْ�	feE>��䘻վ��0>"��/Z�AM��akO�� �S�c;;�x�h�T(+�k�y6k'�h�6Jg�f
�;;�4�;�N�d?�WGC�j���N؇ڍ-�/��4�:	I�"�G�|dc1ik�0$���$r�� �F��˗���A��݂-< p�%��j�W�C1Y������{�{��,���(S �\�eq��4k�������A����#�*�[yOs&Wb��g��B�DR�7`m��A�KϿ�S<iS�!<�m�cc� ,$:����|l�'�~��������G�X���&{Ii	���vO��L!��uA��8t?}�d4��h�>�7X�W��F~�6M�t`"X	����B�~����<u��s�>E���#��)�ҮX�i�'W�߾�����h!0�W��-Q���t΅������X8���Ag}~�z"�Ht`Ð�3����I��^8O�Z���ޢ�%�8�j|��zh.pe����1.V����������C�"�	���RH1�hx��j�~i�ZS����D�|��6Y�҇�4�tR��+-��������R�I��?�wEAh�X	Lq%��!q�>���8	4��Ph�b���#L��D�ׄw#Յ\K���I��H�4(]L�;huR�v���^4���v�B���.�QU�U�:�f7eI �ă��ۊ9K?�k;X:Vq8�L�Sn"��JaT���]h�w�E��-�H��Q�#-�����S�%��mԬ���.=�<MӋs��9Hc-�τP�?B�#w\���@�����S��yO꘲���.��rޑ���,"gZ�����-||��K'�$���`��K�4f�/�a�۴���b��sP2����V�q��O�J��#�Th$űYA�g_h�e3^�s��e��3`kp����:~>�L�>w*��g��A���)�����Xa/�	_,���Ν���֯ \J���(㽮�/q��&��pP�\z���/�X�T!�/�;ڲUc|4��$' �%z�&��2����N\n�W���,��1�x��t���:�'t�} @�4�+
T?��:S��oNq}+��%���j�
�cު]<��}L��@7먖?!I�	̕��[ߏ�_�5(��^�,��5
�'�g�hc˺g@��h���FW7�q@�a����R
�6Rp����V �_)0�����aDHO�i��̓�txש:�αʹ/�E�6� �#��2"�D$7�9�_���n'�����h[�I�T�m�
?��_`�<�=R*�X:�n=�P����B���H�ٻ���k���M�ok��чZgLJ؆�	�����ה����>W<TV��w���F�[CZU
��9�y�,P��F�y�ML|�B�X�t2�T�E)?g�����;٢5)�z��YRero��P��^6�-��*t�?!	�&�y��̵)�Q��]�L�+�y$YS��� �.���%��mX�VjY�eHڊ�}�x�|��UB[ع���q��4uZǉ��6}@�S侰zCr��'���/#0D��G"xH��<ݙ �~ �G��z�t�������>0?wI��$F��� ��x*U�}�5�u<�ҁB��&gJ���+F2�q�~\��K]����p'|�G���%�,7F�Y."�@���"4e��]"A��}K����O���w��\\WA�j	G�33�?@}ۄ���N�g��]r�\ʔ`��g\H��ؘ�r��A�˰��[�����f0�t�;�̝C�1&��F��d�U��n'9���y�-=�4Ojؐ�ϓ+��6�����2�L�/y����R��ы�«f+MtpU��˓����A_��	��t�P�@-�q�V&���+�ޟ���͠)v����L��&�K%�O������#�MS:��GD�,1+�J�߼�z޶6�i]H%Q����s�ïh"Ϩ�r+Oq�)�EJUeO$��+-t�5�����^}�Õ(77:�'��?���pn�_����}]:Ss�v�kZ�#aZ�CzfN��l���i�����B���G���%�!7؜]���6�D
�>C��Z�X�����Q��'_��T�Ń��a��]o�+��g��D��� 9���1A��_�()[p��%��}V>��ڛX�/�� �Rz$1U'�]��֑\���F�#50PXୡ��Q!�;��t�!��41��O���X�RJe�Uf��Vo"����	F��(J���EN���}����'��#;o�2�e�>Z�̓�ϲ_��k$l�@P�s֜�*����//��*�7'���8��h<nM���w�:�426>�c�$�ѝ�jr�G����^����z���k����͜A�R���PK�t�zک,��K�ؖQM�*lG�3tc�N��З,,7�]��U�)�Q�)�il��du�p=��`&[��h8QV@��8��0�]E��;t���������:��J��~܁<��P����[ߓɮ=�}k^��ǐ�/G�δd��r��RX\d��U|�8��L�M�g	�>�UrJ*?}4�P�]A):�q)�3���}AX38��n�������/7��x��f���A4��iA^li�~Vg�g���cw���XN��3%����Q�
�
�Cá��[�)��>R���4ƣwPѧ���E!L}���`l���dh�=b�h�kw1�^<�j�n@�O��q� ����P�B��+*[�qC���,�6N�?ݒ
b0�<)����F�˸�nYoaU�h�v�/=@GN�g����d�cZ�vKb#�e�YC�ifG���
z5��d6�p�V�ƥXh�^�-P����X��u�����fB_���-7������i�H��Tn�3G�u�\c���O��ys�}n��P����s���U)�=|�%3	8ʺ����7a��g(��Lq,Aa_I�/��$��DR���#���Z��ҷ���@��e�BZ����pɘ�ip���Z�ň\�1,4��U�=�H�U(#R�27O�`���K�"�b���>�V�f��ӂ�{��c��f��73�m�e��<Z�g����<�#�������^�_n�:y�'w���g
��|K��X�0���I�O=J��������q��p*y��̉P�����}>4=*@��\	�C�*	�XF�0�.�x�;ݏ�h�C��^(�����C��a��p��y����R|�㲷�yA"��'BtJ4Xy�	�ɱt�r� -�,�u��	�� ��۲5lyg��짿/�Y\y�en���Z�mV#N�I^ĤE�L��I=�`��\�M)7�ϫ��+'p�;��e^��VT�*ͻh��8J1>]p�������W��=`��N��$�b)w_"�:ɶ�-�cD;ZN�}�6�m��'��ƒ!* � �B��q��e��D걘���KE���I��x�}-ūDk1;�V]P^����.rl�c�*I��{I�@�����r)^����VsO2�n<�����Q��s~!��@������+M$�s-(��]��B�۫.n�O���C/����`>E���޶�E��,���P�K�%���a
��X6�I��i�`�7̙�v�f��8��+�Z@�D�I��&�m��g�Â14���ԧ�Q���6�+�4�I�d&ށ�2��vpi���r�S���5��@P�;�*9�GyI�����6���N��4�c�����#�t�QñEv�䂠���i|�1=G����x8rz�]��g1�� �&}g� ������vmo!	Љ���کZ=������]`�Iu�<�0:�5=�m;��"���vj��p)��7u4�4��Y�B?�P�tH�~�ӵ��2`��30�11�=���L�| �n�$�d'�_n��/򍝭5
漑���Y"���?#�؎�4��v�� ���ryLN3���pA ��$�q�,�eA��Cy��\Z��~� <�R?�!�)�B�{�+o������K�T*�&/;��Rb]����"�R�Y	+����p����oE3��+
�G0���w\���0������������,��;�C�m����L+�v[�δ��sJMq�1Iy{���:�P�:�5i��\^��dSH~"w�c��x�^��
���YY�Q!�k��맧zc�:`����+�5pL�z�~��!��ꆄ��Bb�9ڱ-U�/�y��7a�B��J4�QHA����E/�j�)��ț-Ⱦ�<u6���<t~C����.�<�;
[N{2��.�R<�e�~}�zs�u4%�V9,L�-�JD�V���KA�!eѝ�5?��R6���A�9�鷹�$�4�P�#�Lb-I�S��({�%u�_*��<�dp˴*N @�&�4,q��T�&h�<,V�����v��v �@�����	�:Z�RYe�d{[���i@<�M`��z�PJ�X5$��l�Ia��,1d����>N����E�܇���=�=D�V`��w:��rn�J�n{v�^��	:����<��*oU"l��HkP���S�;��m�� ��<>��P��R7�@�:~���Z/b���vJT���:5:;��0abP�V��c����&!�ڨL�l����9��գ�>�gFw����bG�*��əhA?UZ�(�XH'�Է���wV%+�
�?c��/ v0b�ͽs �D�۾OR����.��]���\�&�9���wa�2x��@d!¨%��ӟ32v��mL�o���;�r����D��/}��=)Ɣ��@�B
&����佲����]�,r&��"F�U�^e�]����
�09����@�y�d�7B��2O�SO5�D��9fS	�Tr���������4܇�,Hr�]G��˗�L���l��� ��8u��L�z��6�]��$��������+M��nA�T����o|)AC�����'����(��z�����t�:�4�*�@���2t���ќ���7��J|�s0�l�?�I�8��a� c$�Br�՝V�p.xbh�L�I�Ĭi�@��֣yb���sgq���T��d��r�i9=%���/4������a��醢�����Af��_��Q�ɀ�q��pfC��n8��`����i[�Z�4���zO�$��ܒlK���߁��,�ֺ?�������k�p9E�Vꗖ060�����-u����Q2��Z�����C ,�57��#Z9�׉H�B�9M5�E9���n�q
���|0&sl�$�c�݀�6��\�G��&��
6V�ϟ�;���!�����x
#$E"TR�{��RM��nv��ӯ�6g��ө�4?�I_!�a�����PE�DO�KN��ւ�b4V9��5xS`�ٌ�V8%
�ݺr�R�"��ˢ�^����f��#��:Q�A��^��B^�Y/�za���rG�	�Cr�����l���yh�b:!�0uM�t_Pv��fM�wx���M�p"� ���+���֒u8���|(o+�3懓����ت�v�v�(V(j��-�T/Wg�K����|" @*��G�o
��gn{�:GQ&&"�""�r�a��E�"�ze/Й>_΂�5�A�57�Í�Y/���y��Y>�0!QgԊ�[죺��o��59j��G�T�~�Н͛j$��T��x�Ԯ	��H�S�t���({V���J�g�Cl6��lH�Z>�!�7�`zTAE?�^�)p���4w\%�̟����K�g�Ω'!�
!��j�"������߽���m;�h�g�M���k�B���Ź"�?&U&���}P)d_�y��>��(��A�Q4Oo�3v��*8|��uE�D�N� ��w��8^ۻ�aQa��͍`�x�����K����(:(΃+ia��z�R�=|�I���r�Vec�'䋙A��e4�}*cH�����m 6��W�&�x��q��Mē-�;�,wv��3M}blz~��^b��lbn�8Nd�O�X�9v���h�����A��M��p��D���s)�'�=zU�8�����=�9	E�q����Y��2l�}�إ2���b�b�><��%Ә�
�@�W=��1�A�̤'�[�<˔�_�����A+�{�c�<�y�ϩ�S�ur��ӽ��4y g��Ԑ�� �.f-��Nj��1W>��b�Ώd�?��V.^O��_Ï�Y���{��e��wz�|,�ߖ.��Iu.�n঄Dٲv�&	Up`��e0{�����W*��:�j�	"���z�t�O���D���^����̟���4c��nT:�j�b���}/h-̫{��)�g�j4Ad�
�L�0�g��C$	F��ߘ�l`��0�le�Jڇ�,R���������MW+����[4���#^_����!4�;�|e���Hd;#"@��>w/��F��0a��,#c�H:�����~B%�����U����q&�kϛmh���f~�o��O�[E Iټ�f����C&%V��fh��k�?ݦ1�ݺ�}�w>��ky}hu<���>-��@�{	�j�\NsZB��'FP�D�������?� �
_�$��z�=�le�R��'���i9����5�����i��Q�M���2޶7*�SC#Kﲥ�tWw�G�/���e9^g%��~�1s'����RSꓛ+U��OT��
��BV�غ]��D�E�:�i�"��b�bǌ �>@1uq��a&��7��%ay�B����$O��^SF+�DƷg{'�k����	����|w�x��z7h��@���~���nҗ0���o����{Ze�.:�%�,�>�H����{����v� Ecj�~�~ћ�Ip��φ�p�4G:�C�kG�.#ث�=hs�̧�ꃍ�b���5M��X=1���s��D�&�w,�����1�-�{�EF���ǫ���#��m���JRh~]SR�N\a�s��$~���Ԧ�*%V��Z�"��Z�xi��W��WCR^�oU�u�>�]*>�*�؁'	T��;�mi��\iJ���er�a�ރL���X���goN`+	(�7��Lu�,
и���>.��\M=o=�E[��A��P�8��l:�$_j�5��	Sȧ�ְ-o{���^�,��B�`P���I����;q��hR)j%�-�N�,�`���\}�!�ʳv;,|c]�9��
<2�+,F�t������*'.?nd�����=8��L��\�� ��p��臏�0�
��i��j��O(���Ð��(��4���&g��xO~H�=~e�9¿���86)i�`jI*����q3��^ !|s���P�$핺�	������vw)N�ˑ-�R7TȘ���a��N0]!&��M�Hu,q�RYFFT7���8��_�E]ی �wct���?ȵf���$�R���	�i�>��/J����{Sl�}v���9l�mtII��hU�Kv=C�R��	�Ήܲ�w��竐|�H
G�+�>316~�@knU�H�D��`�#�X	�%,sd���Ť .
x�S�Z�Y�"di���]�[����$�*��x�����Jaů�Tm�ij��4q�FWcP�Q��_.Cm� ����o�8 Z B�B� f+����ѻ���W���H7�n1Gk�@�Xٳc���w���f�G/'Û� ^���Fڬ|���̠j�<����a�~�[���h����Wd9L�	&�{��ڂX�����\N绵��f���Fl��)Z+��$�����\��g�:����S�A�6����zg:RW��J ����V.�*Ab�[�ln+4g0��O�m�n�<��B�w�3b��<'��4��!����GHO���r�<-��g��o�֮ҩ�W �Rs����>Έ[c�:EG\�=T�uSD�[����1_��yCCi�8��]�OL�7rA����E2�q�V�n��C�A��'o�,�y��{\����Qc���~cS�3�M��%h�i�L������"��S����|���q?a�O;O�^Th�5F�d�L;�����Q��ӧ����P�<͜-N ҏ�A1�dj��Hf���E���=%"���U�
�[����	9-��29Cb]�#t0rlF�ѧ4�O��e�ΞO��8����+O ��Z�����
9����5��U��?�Aq��O�)&P�Ś�9���6����(�%���z(̖;q������T�����r���+v4N�sA�W��'����19~)���y��=��8R1^-�6�d�>V)ݙ���m_b����V$2.sўu-�8��C�g/h�}�!ٻK_��k��&U�t�%¹���P��1��jc/�Dkt7C����Kq�h�O\Zo�\E���`���1}�Fn�P�cr8���݇���o�Pkܲ/���?p(�5�e�$�|+쏖^a'�ȉ�����d�F���]&��:v#b����l�ɠ��Jgr��\�Cd�7MfO8ƊN�x鋩GeR�'AN�����0���0�z���c�wĎ~D�вZ3F(��E^�0�s�� ����F"5V��b�B�c,�$�9(�+�-�����
��C�
��c�}CX5�2?���
%�U�$32�v>��13$�v��f8����~��`Іf|�}���Z|�z�g5ć�����Qa��AQ����Z3V��FL����8"��;��ӱ�<%FB�֓VJJ��ދ�l�́]������2���ctT�lBP��ai�('º��n��2�����~KȐ��q�"lc����M�u9���{��q����������N�m���V��<3�V�ߵT*���^�@PC�z����6�g����G���b�a�4��ݬ�|���w�sô�l�ڟ��J$55ы1X5@9Еj��L\X�N��Ŏ��ja���:������)|�:�}����X�L�
fR�dů؋r|��~�\��.3C!B�6T;(�5'���<�=�"��:kjt*�%/� �5�)q=��o��C�+�ڮ�q);��F�No���X�[����2H��ܯO"8VL�gRjs/Fe Ρ�&c�TP��_䰀w��v3&o�W�����$��|?L�^g5j{|����5���R����n7[�Z�(5��a@P�����'�a�n�lr;=�3S[=��i�3�	�k(���E���mY������Ģ��h��E?Ϸㇻ~��"c��į$��#�q	�+F��~]d�=�;fd�^���]^���<8ۼ�����v�^G�P
QƚƵU���q�T��%��R��6+n�,7�]̓q;U���>X�)�CV�y���T�9\5�PQ���ׂc�UfU����}-���O�-�/�S��?�u�p�b��>aͱ���Yz~���R�b����e3�՘�G��@侲�j��D��܁}�$y�Ɇ�#kH:��9�m��D~�v6FV�f�;G�w��s`�c��[�0��ɇ�?�V/��y)(�D2�兯	3�ń��	+�<��[��)�d(ғ����L<#��9Y�s]u�v�\��M�?�g��� �9]@�*�F�#
�TMᔼ���^����D4 �%dʫ�5ӡ�����`;�~��6}��T\�h��R�5d�;oˡ�x[}�BF�e�.R������o�[̛�|�?|�2�����{�S�;���%�=�7I�� a���Ǳ(�rt�c��2lX����⦵��W)z�S��j���A��L�bPO�Jax�8�UY]j��O��5�oYfL<I"b��[Y�AE��$��K�qaN\��u��Q��� "5�Y�6x��٦�� ��ddw�M�w�Il&=�]�T�eeزF8���x�Ҡ*q�p�,>X��"Ҥ=|n=S�6���V���;��r���цm]N����7\�� ���Ú4z܁b�g�N�#Sy�>��]��5�������/�(�Z.(�� ��:4t ;ղiq1zr����=?��}U���0m"0�ab���Vgwg=/#t��QA���r=\kQp�QM٣��@W��鬅S����̵��o�Xv����6��
���IC8�2�'����N%�E�Z�RAJ�w�&|��&%%��*�8M+l�v�( N�p��qޯ�*�,��1}��oέ�6f?uD� >~Wes��fMr�j�I~��A��c���j��_3vl֐Ӽ�'�0����7��f�De�D '����j��	�RpGC�6�zd=ͷ���D��*�{\���v���a��Q�D./y�rƌ�\�Xs���&B���v~ń��m�M�"]��ч���#"���I�~S	�	�~�l�Hu3���E�t��E�g�}���\T��l��a�r��x(�o�
Be�n�3Y��a�0P�M0�f���P�|�~�ɒ����f¶+�U��{�~�C:�3� 7�Ff�8Yx�\�R�֬�8��bb@�Ӏ��N�B-��$Gb�������e��:.�n ��ꓦ{T.�R���ՔQX��uz�k����<uG�zF�������L�݉O�"`�bJ�p:D�&I�j�^�TL�ێ* �=1�����iG3�8�*���A�p�{^M�T$�u>����,}Jz��VH"���<�=�rs�Qd9�˖ 1�z�;�����o:��^H_�{C[�ߝ����#id�P��MEU��^�q��C"��ڭ�F+�.�<���%}��+��1�uM�]�!��W�Nխ|�	�v���f��/���,�ot�P�]���? �"��[w�%3��x_��4c@2���L�Ӑ���g�k�#��3L�sb���U�����i`�����UQeS��ۉ��?���hS�j�@Z��bY8���Z�_5�`	�����"ռ�Ut��W+!P�R�y�̒0�:�W彆���E�լ�N�u,�߀����<�{yK�-yo�y���>.�,E�od���h{m�$�����vS3�H�(ϐf@+6�~������v|ܫ���LmMkް�����j�<�=>5��Hfd| C� 1n ���2���q|�.�&��k��ώdf�4F�ӡ��f�9x()�zb�w)�>�xe�$�x����>�.dG~'њ����u��l�)����6h�Rz W�x��@!�	x�Ĵ6"�L����X����ߪ� ���Ks%MJ�`]QZq��mll�C�W���u����+1@N�8j�O�W��(��FZ�;�#�1���fJ)�}����q��Xݫ�VD��P)J�5�s�T�ُ �G������uH��9����̓Z|4C̠��,��N'��>v
Y��"W鍆}n��L�����2]X	Ԙ=�+h�w+�M0T����U��w^>e���{,-�5�Ј��L��:��=�d��x< 0�]�s��F��K�����>�{)����}���l���p��o�H�Wƣ�b��%8w�C2e�zh5Ap��Sya�RPR�G-)�Ґ��8��g;��[t$��.$7�lqgk[>ʸ�S�L'4A���\��n�TO`�k;'=���c1����ȂaVm5fW��ڂ������?
T���b��R���p����4h�+2,�a����pz�����:q���h�6���Z��dׂ͹�1!�5X���>fp���U?��9|�vٰ�^�,���7w�o�mJ+!��ȶ̉�w�y��vT8�rETi��ªӚ
oZ�~lf#j��7ec�LH���p;�36����t�Ll�w�#TM�]Jr���Z�n͚2��<�� L��uu{d�F� D���H�"���V[đ�(�p�'qe���Y�P��W�d��!>da���gr΁���娘�<(�Y�L�4��hG�KN�%��J��6���SS�p�I}v���@�eY�QLJ-v���A_8=,i�;n���PE�.;t�1!���,����������_G�;4�����2u�uh �ga�^~����~5'���NuI2����Cg�W���'��	�΍�P�;a��Z\��a��pE��t����~����5���e���"rM��;
	ˉ�1������U��~d$�I��H%��B��f�Q���2V�SS�;�4����6 �jd6�2�-�W.7/"��ju�#˝_�B{�}���nn�Q,���h��p#B���[����U�~��s357�jgƤ��C�
D���M�۾��+5S��HM����U��7�"(���s���*��O&��i�Ē�en9�섇H�����\x�ꉿ��Ho�m����J�.��wU�F�]���/���G��yN�0���e�SB��S�v�Ja�.Q5_�@!�s�7��?n�j����O��z��cr49�h���χ؄��vcԇË���`Q^(`��Q�{Ckmf��
<L�^��'){�|�-g�X���=�;��ܔ��d~#(f��k͠��2؜��As���F�A!��޺n���ʙ%�34�>�Ú�du�	3�6�vΓ�q}�H�Q������ř`�4h��&��Y���3�3~!��wG�=ՂAh�S �j���]
{�ݝ�:���U	9[��05��:�m7�-��bĢ��D>��³������\�����>>�}L����b'ޣ^����$*��<�j�Qr��|.gB�X�y�����0�͌��}{���8�(�`�Q�y��@?�As���!l�'B諁p����������Za��x�Z����@�唊�У|��l:��T���	W�40t�8���I{x���|��C���ȃR)��F�FR��2�9�b���9dg��, %��؈�F�fT�TiC�>�B�,m��VO�Z���)�Q95��1�/�$�@��t�)��ˤ�H��P�t�����9/=�!���o�e߱�g�2a�� �����p��d����I�V����8�Y��2�=D_eS�*ϡ�S�	�����]W��?ju�o�`���p JN�^��-���آ�Eu��o�_�3�Il�^?��r�n�r�V�w �z��9�)��HTb��������G����_#��&�ܖ;��;��}FL�{"�},L=�ݮ�������1Ū����ީ	�/�@�ȫ��+�%"N� \]}����a5pX�~pKي�����Ȍ1:�&�z9�e��7 ����}�<5o��x��{d�z>���>�]U����$l ��[�ܡ:XbW��.:gEI��ub����8H��к�*<T��!�h��ȳ3��!N�m\ɕ�rnq/`�Q?Z�� �$3�Ed��69�^ �ѧ�b��_��&��:���5TA|�!�2�Ȅ�7��}���|!�n<w��߰�����K����3FL�$#��T���*]Oz��%�pu�+y��1�k9�A-۸'�@9��B��֟įG��_��3iu:�"� =@W�Aeմ�9&@����OXp��A�--/�V��@j�p(,�P֏{nI�z��Q��iT�)�L2l<e����Jϔ!�F���7Դ�j�8�����Ը�ިI ��4��s����U��o�i;�����f;�r @9�^,�����唹%��B9z�J���E4Ȁ���L�S�D�,���1�(W3��\.����yc�o0�+����{�f<!.�Ck����g��sc��ن��~ ׶d��A��]��o�A�}�.�ٔ��!Ds5�|��k��3e�5�.iU�1�9M%Ȗ�! ��]P�� �/�-��O�~��P����Σ=Sy\����y���_T�E([��1P�O�fT��0��ȁ��a�-$�x���D������Q�f$i����G�}0���������gÒ��bչO2�f��@�D9�� O��1��lPjj74�S[;0h�n�ct��s3�\ll��6�(�%4B��,0����d���?���PAxK��)�"�8���?�chO\����K�{R���_uT5ۮ)�b�f5��	��"���]����_RKp? �}^3��?�_�ڰ㔡a��+ٛ
'��=�(�f@t�T�l�_��
&6������+������"#��@c�V	�c=���l��L��]��$�f���ɷ�ɖv�i�����K��(�����6O�t³#kb�7�p�E�+��V��Bt3������u.����p/�z���{ۑM��߂"��?S�w&GX拵�%<���k��+���T�:0@�<Xzm�A��u>
�V&�n[�X�2jf���D/}���_D��C��]��#�

�8�l��
�	��:�|�a���%K�`{����E]�-S���gE��L�Btͨ ��E7:�{E?w��2�Rts�[rfJ�J�<�S��@��$.r0�b`��(7l��}���]��AT(Ij�飏>(B�Apހ~u�����D]a�@KԂ���AȪ��K&�)�%����+_?�����3�����R�02Ē�>d�җ�'�
�<CV�BL���$�u��\ ����T�*�������N�����X�VKY��Uax�[����H�rf����Z��-�2�����n�=�|u^�P��E4�yC߅E�JV]GF=�s�U$��F�t�f5�����:��;�d�6�q�2�JA�8�2��LB\�tmJF!��H�?�{���dViOR����v5��sj'������������p/iA"���mN9���`K�5�r�K�ܤ�es��,�{FT��	@tFD�⧪�db?���8(6���D	�_���Ґ)�
�Ryv�1�,[��W�z�&1F��k�nC�m�ݦ��&���̍�e�3r�������na'#F���ד:u@��6�����`�M�ډ��9	O]��f���x�g	]B,@�;�Q�+���@{��]��rR�dIc��;i-�Å�p�R�'��`|�ym������q��q@f����a��q�Đ�Ua��Nq�� �� θ�Q�^�uڡg�Z����3��X`Q��������	_f1��KQ�g�O�ZG(i�sP����H2��2�l;���o��Z�ۏ�b4��^r)a��D;��&a��X�>����Qpfک����)�^�*i����� �_b?;o�Ь
���ƾ�a.�}m��杹���)�R��
��Ҽ����5��p�lyq�0�`J��2�Jᾑ����51X
��
���7Mi�ߚI1@��jy�5 m�=9 �����,-a��o;u��WL���1oQz(w�({�6�x=G�-��*�F�ل�(� 0[D�ݴ�0ԭ�*���wf7�i�}�~o֐�l���vVS�b�&���f�2�.���.��u�W��� �K·�E��i�kP��Z��Hr>�G�1vY`��:�+5N�CE�����Ȱ.܆������-'?�2;��='�ǟ�V��f�;jCS�:TW�P_)�zb޴1@d�C<i(�l#@w,eBP}M���/T�+����a@O;w�Qsb�q��
:�d)� �^��xg��\��à\E�
&
�Xz3�Z���m�<W�2'�o��k�`'���{�g�fc[� ��dڍM�o4�=�[�������(v�5ۧ�>M9��|�Z�Vk0��J53P#�I�&�����wRd7P���v5!:5�������xS#G�gkʂ=L���)n�Ip�J~��Wrk��X�;��Wo�8c�(,�6�sA�K8ۑ����_���b����~�`"��My����K5RcŜF^�xV��jV����l�-u,�E+n��I����*3BHi�x�uEZ����%�A$������oyG���J�:I���B�$e��|�x�H���Μ�E���IzO����Ի/A�rم-�D��{��a���7�݁4H�B��ނ����= ��X~���xhFI︄H�{q���{�AT�p��m�Z-�߈�{�|��e*sh(�d�Ь�x-I���g�Sj�튢A�8�D05l�۵s�[����c��*�.+�n!h����Y��� ��	q��^�AR��u��s��iI��eNr_��U���E�q<b�_��LYH}��י%�����?/�Y��Ȣ�鍲u���)�>��q=�n��:$�v�|���\H��̙�;O-�t]�fyx:K1k��W�Ne�qy�F}lO:����S���Pa��,��g��Oa	��,��|��ߏ����`|�.~��/)_�rez��1|�}
'sw�,kس����	���BN�x-YI���E�V�l&ނ����+ߍD'=�Mq��.l~�և�!�)T�w���3���`Ł#�՚�r,�ݼi�(�I�9+i�%�	���Aw�J��j��\��4�*l|��hZ���C�?o��*ţo�T��h�Gxf����k��E�=f��ˡ�膘|GO��+A��?���Q&>b��F�q͖y��G����PV�[z����bwvgk�ÿb06��>��������́���	yͬ��E���{ؔ� �ߢ�"vz��H����~����l� �������r!W�J�Bƴ�IR�?%}�M�C�ѩ��8��. �$3�s�������h1Y�?yk���ކ=�L%��&�x����b���=���\�j�=cw�%G��i%�|���l;V�Ue[pېc5����Yz�ܜQ�i�!|ן�!��霫��<�pn0�l�c�����,��Q�&�'~5G��V���߮�P-��Q{���!t��G���������Wp*�8"���dzqT��ϛ
R
,l�YN>%5�8|����n���Q�~��X)t��r|����E��/9���˳g�&�]Z��Z��]�)�!5�GNF��LE��w��5+"���m�x?��y�"��r�-�~ ��݊g�U�n��L+F)�����s��ٰ���W1�4���\|t>
ve.��UvA�T��}Hkȭ�����u4��Z��Lz@ǲr��'V5U�.��K+L��{�p
ku�w#�(�7{�lk�*p7
��/K+Y���e�y�##��H/�6 �v%��v�~��ck��s=F�ѫ���s������ۓ-���u��ա��8^����>P�TrJ=$C��o�	��_�����TC�V	.D�T�ة�Yv(���v����Ll��K�QՆH&m�E"7l����{ ���`],��[}�&�u����чM|�N��GK��Չ�ni�g�Т&���&� .M|1Z�%!��8����pAю�	Do��-@ܚ��ג�EZ����D�	��{d8Zq����o����KV̚CI�.?2��"4.c�sZ���-��&~J6�C�+P̃}�L�d�G���Ը��݄�3�~Y��9$���		���K z �C�/��������"w��%.�*�F�B��w�Fu���W��P/���\�\/��I�uuR%?���n�W�G>�U1_�(��i(��i$��\f�j��I���u�W���:?`!�A��@���.=�u\����@���5�ǒ�6���#�����&l	���la��4d�i{������2d4j���z���^�� �X��n�/�w���9�8��G]����|�{�0SA�l]qSC�U���FR�/#��=VK7i�
0`��k�XShC�ey�o�k��8���
��_3S�R=��Pm�<��7��5����4;P^��8J�)�-j���H�c�kx��:� �l��be#�<��!oy=�M�vr��� �4��G��MȺ�T|�b��Ek����ć�(,�M�zJh�Ěf	MN�^[�N��"��^Q"-��zE�A�Z5��ú�S��ň��\���C��(���.U�Rо�w�|_<dt����R�F������PY��M	�jEx/�:���Z.�Xͩ3��΢��J�	��t��!LE.��6����,7�Pc�>v2
*j�C����j�$lc[���Y��9�����O�����
���Nb�\*�+ȵ���.Hhu\��M~�jG�s�u�r�r�{�wVAE�.w��q�]S�N�ݎ���z*��H�:�l��؍�t��s2_~ĉ?8�5�|N5b��:s�bg�q���4��y�q���$�qփx�v"4u��j�g?u���<Zp�9qQ2G7w*��ݕf]7������D,CU�-����s߿�`���r��?�_��A� ��!��Z�g}I/��i ���У���m�>8:k~�ȩ�5[���	����L�y���q!���溹��cL2
�*]�[($Z�Y"=�]�ɜbi��6uQh�y�Cs�
���0��Ш����#� E���ۍ�e�e�Z�Ԓc<��*N�E&ahF������^�����i}��ws^�����]t��Y��V����詛��W��b�g��JIJX��E����]$(�UsenS����FK�!�[o�� �F9W=u�J��çe}SM����Z՚e$K�Q�*0k�i�`�q6�4�Z<��jX��5��F�����a}�E�΄l��rkk�(�.�a)���~m ���Q��M��6��%D+�(Ƀ[n`����1Y�4�4R��Y3��jp���c߫JD�ē��A�f,������x��'n�8P%���j͇�����؆g�8��ك0��Ju+�QH�6߽r��A`�2����!�ؤ��kϪ=3�s���ҫ�FF�S���l�˻8TD=���n�tR��3�b�f�y�Hۭ�%E���Sw���-�x�����G��������E��K30��񀎉"���)��v&`��xO�i�O�t�U��m��a���X�C���~\����HL���b��oi���Lܛ�z�����'� _����Ci�A4�6aaw4Z��$Q��N9/q(�UlNyi�i���o��k2�w��-Q�g�����|��Nm:g���_��Y#l݀���̖��ϼ�|��ozܸ�2��T%g�}.4!5���2��a������a��Gw�1z�/��Y��n�n��obK��n�yX�b�d�#���A#�D3]ԺI�#[���3_.mY�݆ �M?U̫`Qf�%%{��k��L��튵�=?S09S��i������D��Y�]���V�KP�\'�E��fH�3���,Ū3�WtL+��a�ǀ{�[���-��lz����Dp�Ƭ�h��>!@���'��lW֖p��k��7���t��H�t��VE�|v�[���*.$��!�	�շ�cݼOO6�B�QP�֯c0�P5]]W��5�
p�p��ؗ��p���ur/��(���7��?�jv��G4}�7mܨ��W�r�C3���5�ty�-瓻Ms���l�fPr��=�Q�+�sp���̝�Н�mG"�6��2�``0���[�:�������ѹ$Q}��~�����[Љ���j%�Hp�lO�q�mS�|�u4(P���j�V�i�6D�l���")x^��l�1���]~h���-3����F��/uw��I5���*LE/''|���KqO\q\Da�0����y��f0@7
Bլ�~��8�C�ig���3R�%�3d�)��p/r�Q$J��
���NX��y~����쑮c��(���bN=Be��Է`?X����s�� �Z�6�
�RZZ� ���y�ރ�.YB������� m�ҵЃ�c������f>n|�51��K�݋���C�����GV�JF��U�'V<�!+��a��m�hx�q���@%8�
]C�A}��>���M���D�/�@�s� y3�7��t�mޠ�����GET^�`�����Bf-)<���,]J����|������%��/%�Q�w'�wăxybR3����k![�D��b���x�υm�� �{��lL��������I����
(�����d@i,8bك!�%N�y�m��H�x����:f���S�WsoQ�tc���V[��đ���R����1AB��6P��ET�F֗�F�5`��X��	
�����]��G�j���a����:ھ���)��u��u��1˛�.{�Kb@���:D�w/I�L����ӭ���z�ؔ���k/��%%� ��#��zՂA�í�_�j�h�g��WD�5��s�V)5۶mix�cZ ��ѯDu��)�\�����˹0����*���[���������<=�'���3��fՆw�;�$�s����v!Q�Ϸ����xk6��P��H�R����e����<;}�!T$DbDXq88w���N��ENB�Ƹ���R��Bߺ)Ǩ��qf3JC�s�x��V�����cu�~��j?=�%�$Dʖ��Z�Q�?:\��p��Uc�}}��U��Z�N}[�n��aÇO�%H#,R9��
�IH���I���T�1�e�{b�(HFPYer�M�^d����ӝ��{eN�a�Z�,T%�1 �l��?����i��;F�I:�{��gBR����4j��V�â��Fxd�h>A�ꍫ�q���?�Ficx�%I@��<ڼE��F�������0Z�	�?f���}j�:]C�b��3d[W:��y�t
����	]ab��I�;�B��I�R	�5[�8�U�8H�D
X�+�8�I�T`w��-�iv�#��1��J-D�V��$��M~Rh:��Ftg�,j��
�n��њ�?�w%�UI��	��
U�\@���p<�.�5�I��,�X��\�d����7�]�
tɨr�a��f��"��
j)�4�[v'�M��V���ړ��J~�(�*"�t ��1~Zg:vrH�}��5cHBrI�CJ,����˹��36����Xs0�	 �e�v6*XH�/�\  k��@�γ����ر5��tؙ ۪���C1H�u�L��X�ֱ���v�,�S�b��o��QI~��#FuӃ���1�_߂�T��9$8�2�≮q�o��ȳƥІhN�s�Y������+u/\���ۭXj	��`=P}�j��z�U+���5y����ߓ/��8*չ�`� ��D  4%�0�Qf0~SsZ+��r�:�Q�sd	KB9��=y�
*=��[!*5�!A2Q���8߀b`�'����祲-�+�B��{�??����������� Z�����Xw8�ö�鼓H�&���k_�W�gF���o�M��1��v����'�h'P���C����$��
[J�������2µ�(�?W�Yb���מҤ֯�0��O�l��&���E��ZG>���o�ߴO�j��7����{FTG���}"j8�^b��J�MJd4:�3ϻJm����{�^B|D��E�;8 �?�'w�Ν��qh{��(��\��J�l7��/����w�9sѢV-�����e�V�)W���Q��=�W�0rkX�}U̞�`�g�<|c����)o����c�#�'*Ҟ6|U�@?'NW���J~��bQz[אb�������"k�=�[{ ���(���yD��j�M5u��=lL���o��u�U�(���hD��kƄ�J�9�g�m�v�	� &��� *T�=�u��!�����?u�� �}O��$ �Gn��4�d5h	��{��ܒ9W��'D���c8x�"�^�뻧E�w�*ob9B~^�j0v�wuw
�L�h�r�?���4㭤8:3C���0��4�$�0`f�zxD8+�o��<�KҒb�Y
A��ت_����E�KPQQ��g�$�^� �
��S]G&?5�ȱ�u}!x��������w�W���ɸ\V�RO�K�۳�%���X��;gVx�owW�>[�]-J��h{�!�ak�n��gZ�*Z�w^��.yD
�: qu��?���P#�m�N�v�<�I�C���42������x��L�e���=p���.ʳ게#� ��u ʡ�%-[3�7ş^k�����@���P�+�++t�z�y��9:}���/q"�N�l�	�Z��f"Ȗ�@0� �O�R�H#��,����`�"�C`����s�r<�8��R�U}�	1�Ȃ�P��f��v���l���!�K��>@�.��� �ܡ>?E
��Ky��.Cǋ`�	�GAʘ��Ո����1&yB�_zW����g��9kVb�Zߞ�M�(��������֝���f������+�=�'�-	L�Ag�jo�jh�7�F���t�z,��{���� �SP��j�n໴���h�Ld�e���u!��^�(�}�\➐��h� ���:Z:b94"{T���g��S�J�������;D�F��on_�%��
q�"�5/>���w��U^eR~܆P3�	Uf���D��0	�:��Ex�m/��Q���F�db@�"�������5?�����Wa�U\�d|o�  ����Ϯ��	$��9��A�l��uF�����
��x��_�c^����i	�~9����vL�4�ѳ_ߊkԠ��w%^O:�m-_�5p���7_F
M�d)�/~�3�>w7*��n�pJ���))	�/A|>Ƥ�\���F�BE�Sܡ�z(H~�{����tT=b�ŋ����=�G���`�	�̌_�� ța���F���{��Q���S��;�]z�]����4'�3�2����� ��UP���7k{RXh�4���0y���o�V��Pz�|f�դ��p{Gv�\NX\%�T@�M�!`�q���$�j] ���9��d�&��jzɌRo�ƌ	�<�8Sa����Ǫ�8l �Ê�;�������9�)!Mk(=Ж���{�I�T�Xן��:ɨ�i0�-ڼoƛwJ4"���w��[=8ҩ�k��r����TD����]/Ɖ��Yn��归�L�BX��迒�ә���Mtk�.y��n�������X7yCL&q�]a��>����b:���$l��]X���� p]I��$h�_M,�V�b6h�[�	�U"P:��22wˉ܏�{���%�>�XHW�`�I}�2�VR�=�Pj�PqR��(����}��!F�Cޡ�^e��`Mò�j���7]�,._7��!.qR_L#�_�1n:�����ʣP-���,����>Dc�Y�/[kM�t����'Q?�%b�%(RS�q�Ws�Ax`�E�_�$���X\��ò�>���~\οM�����5;Mtμ)aTR�}�KY7�$��m��~(�١����Iy�7wqg�s��r1F�|�i�<y��&D�ME�ԋ}�����fc]>áb�߰D9gd�6�O�z�BAH�qOP
��&���+����s�޺?�Lc����J�RbK|N����J��9j��o�6�����^s(��4��q�QʄV�>tP��!�I�\�x���F,�`^�-D�V\��)F���p.�"����/���&|]9�7k�)�����_����o8~(%a�1�d�X;"�:L)��e���J|�ތ�À��>$�������c����`n-?3����/�˘�?�>V�m+�Y	'���A���N��:�T�6�-���e��V�2Y Z�ԙ{\�\3.�G�ld�X�s�Z-1,��E.����,��"'�����2�ԍ���F}�{��d�pKa��͊���Q%'#i����FX+9�T#�YQc>FG'*r���[��������z��Đ�cܜ��p��:W�ܶ/�������Yx����
5�N���jP���&*&Rj�w�S� ������%0 �w�mcߏ�׮�Y4O���I�$�� �y%E���-<�V'��f{�!�/���[� ��PT{�������	 +�I��e���X�qv3�+4�-�͒�싁eYu?�O����#')����E�Q,����.<��Ǒ��&h��(V0��P�q�A��Qx�[xP�kY�H�*��)�!������;m�v�k;2�-���P���f�\�fL�8�e��#��}��B�	&~�__U[-4)�(�U~���׈���[�rI���I��jAx"��0�&�&ę;A]���T�0��Q�u#~��e�b���G"���cF�c�����,�,N�W�A�F	?г@��A���$\�� �M���õ6a�d����K���~5�����a�W�k�j�<�t���I}����ݲiAO!�|�x����r��7��la(#��>P{�C���Ft�Qo�����u������o!}lh���=�,�
A��$��3�;�ɮ�d���w�]��2�]`�.��Q���c����-�KTf�^��6�B�7�_j��1�%#�y! ���$^��?�z��������t���P1��.͆R�R�w�����3%'�2�Q�i+`�1%����k�;�sʩ��8��?�����K[@0����/�'tE�a|D��Y�����$mTd}�c��&6�ֵ�Jt)�Z=%A3���CRZvW4#Gn
rQFO���2�HБ��3)��Ҁ�$��,H��c�}q�QZIS�����"N���n�ɚh�P�s�_ ����6����!�>Ob�����g0�d~.���QN�u�4\�S��NrIr!e8��; �nԼ0�U$-A���zmI��tܗ�k�ͨ���-5���Ӿ��m�lȍ��y�9[A/�t��ۊ�;���w)�Q�����<В!9���`6-�IE��J��iu�~��\�T�h��7裒�7�X�mM6��L�)C��Z� �~�^'�X��U��P�֊���@-2�A�U���B�K7��r�U���9"�m�H�@������j�����~�Ai� ���O��E5�F̰�D�R@m\z�ʾ�WJI6��@���9[�D=���V�W���άGj�P>��7{i���[��ab���+3�k�&��ˍ�&�Ir��)��,��>�	P��s���~��SȮ�ю4(�L"�s[۬�=Ec�1֋����O�˰R��c@����T�~l)�DE������Q��X#��\el��2��d�5t���rM��B~��1Ixؼ5�P��r��ZR����^�F� �ow��#p�W�m�+���s�~:�55� 8f'^�_�����-iX�����~��@�����U�ϑ���	U�&��~�7u�::G�+��c�[!���f�_D;zR��s�����HIOD���i+�e:���m A����4���{'fl������N�ʮ���k�(��$T�/v���h�W +��5Ͽ�?+��Ͽ�Sg{}Q= ��;~pVqǑ�lX�,���NX���g�Hva�ΨQQ�u���|�����F�ȁ�?茓���yy,)>2K��9�WA=n�cz���(�X�VM��+�'���I���'�:IP�vQ.Ј�u��V�4��j�A3{�[�.'���%B5��
��fK+9q#���O@?�o� t��3��]x	A�f��8��R�����-��B��x�sL~��z�(���Z�e��.�j:��h�R��!/�Y������#'���Q)����.���;|]z(�B?$Z��V�R�v���!��$쾳޴3`ǂ�v�G�(H�/K����lו�>E��;Ek�,�꼁Q�W����D�Fe�����Ӷ��;5��Y�k�(�� dgO��@o~Յ�`3��sQ�������NB��߫YU�`%�+N�l���e�Zh���H2��yV�'~+��b�W�$�lП��	�n;�d�#斸%"?�,"��t:%�`����"�y�7�t�;.Ȼ��c}�\���ܜ�[��_C��Q�P)�XϘ��D+����0O��:�~�K��_� ��nT����s��e�Q��}��!x�����8w.S��y����v�Ƶ�I>)$�6U+�`z�.� 8Y��g5F�Ӝ����g�o��UJ�zƐ�����+weuK֊���	����d�,
��� ��,�����;�.N��F�R:(�I�$*��D��<����r�Y�h��Ql&y�{��)�5u
w�����,b���_��>��l,�h��DL�6mH��
|�P��h�G��w��}ݾ����P� $�>���<{f�CjMtpv�^��Bg��v":�y���H���.�Gg�eg�2m��L�8Yi_�<p�r�#���7��s�����=��i��GƁU�_9:Y��Q���Ispj̬�ް�r<�2 ����G���˭$Zz�b�Jsu�WO{whh���S����YjU���i�6����ws�J�s���
����$1��0�?Ը�Q�Y%Is �>�\aa�SȌ<6���:	�v���H�ʧ��������O����FWy�U�7?�y@C�qJ��㰬�������i��y��=;D��B�aè�$�Cţ;)h�Bŀ����6%Z��2���ӧfX4o�j�dFr�s�a 9+X@�dPc�潈j(1e��g2��S�g��ڊӜ�ܲLR����hR#�foF���D�5l�;�ۃ��A�7jv���s�f+�#B���B�:�ַ�֙�6��MRg�)��!�~��_�u�5�"��ðð�F�<�{T��(~�Aq�G[��Ӥ3,b̘�i�YY�)���&��T��]�~M'��_�0f��[�V�MKQ�����7�$"�=��v���V��z�'�)�ⶒ���"�a߱�t���m�xֻ_��� =v�>�����wF���=�!2�����p�5`=~D��>�fA;�B���8���:��7�RwE�0�Ms%�E]`w�^e~7�ܷ���ڬ�}���5�u%�]����0�ү�f���?��/|��ڕx���k��,i�,��B�"�D�����O���g�
��Ϻ�V�"]���k��i�&f����m�O��Fº�^o*����p9����|xS�} ���5��m[�WU*}d���V�/�L�5�A�t��#�$�y��̈́,ulC�@���P�G�np8)!���=�,R$��#�����,13>%1MC�bk�@fWÛUcY����^��1c�+���l/�a�SWC2e h�[Q� ,�����si���u#}�^z�c��Rk��7,�t%�5H1=�V3	��]����Z�`铖��Ü[�%��B�p�c��"�7.�s>��!;�+X�M��&CriZ��̼zW���L;�?����<i�����z]�.Z���=����5&v)@�q�ÕyJ��!Pv��;5���(��:���(����jYa�9 �Q�U���V�JU}����{��@M����k�hЛ�al��m�9�KO,���+	��ıp���#Hы]���bД�4 �#,�۶�����?��1�!��� �#*�gm��E�ʅѳ���"��������U+�uwH�U�M�����m5o��G�ԏ~�� ���Z���L�Oڥ���s�I�$D��\_�<���x�Y�:8�E
�p�7�f^3�+�\d�WY��e�п#׊7!���&���nޤ�㡻[������ӳ�Lv�r&J�Vxǈ)�ב<a)a�]O5���j>�m,��Lt����t_ۿz�B�.s.��ğ>���������NOr��^.�鋎��!�=6�3� ��B�6 �E�qX|��a����"Dq��1�d���c���d5u=�!�{�H�g����(����H�Ʌ��K� wn�K�<�oPV���nD��K��l��_߁���l�`��m��\�rU�����9��ˢ��^j����j���qcO1��Wd��Js�0��F��sZ�/��>[d�ey�E��%�c)������ؚ��"�OrM��q �*���a!+�'8�b�d&�	�Zg���4�9�c��� ���� ZBl�H�:�&�yB�!���?�L�*M`eA1���G�I�2��Z�r���f��R$���)�C��j`i��Gm��uF�|�>-߿��%��fT��&���YJ���I�0�G�'�%:����7�/%wd�@�ܘ��XUz��.���ںd���7�-Jĩ�������yo��-�KΚ��PW��P���t���HT�dEԂ���
{���ˑaF�����}~�����B��n�ؚ�gQ�u�1ib�8(y�,t&!Jش����n��}7�g��:�Gh��v@�����x ʦh�CUK�W�u<�AgT'�b������:A����w�%�	�s�֥"�Վ tfe�E���@h��-H���K-/�D�'��d�zP:;!Sk���"A��_�3�!76�L��wx��x�p���莅���~�<A�k>}�(J�g��J����'9X�N�Nl(�:=�(��Y�+��ʗO٣��m��Yf�p/��vk|�FPqs�Ny�X
�f�/ �������s��)�ƣ�l�Zʲ��㴆$��'[P���L���J\�V���+C5���Ѩ^�<���t�O_����%d͠n��|H9=�X�Wߕ�{L� 9���W�E�z�/��w���[>�l��H�Pl4X3f��K���:8˻xq�c����e��*��N�AN��=՛T~���Xr��v�kQ6#��Z7�.���=�ʵ���#���pf����o|�|�l}�bc[ZJ��1�m�z�Ͻ���N h�t`تc9n"jDu�9�,<H���+T
3�?ϕ|5��#<�S.�n�����9J!D+�B7+��B�[��^3o�LsB�#��@�"�.����j�M�EI��"����2�pI�`����0�%��VA�������ӓP�&�CiP�@���}�/�s����7�v��\�+|M�^VKn�\cBQs���@�tڝ
Eg����[��;��wO�r���`��R�'Ei �H��T�u^i߫q<�C"�N��;���)�_�W����N�,���C�.\�['���'S�ق9����iVI��J���}Z��?h�z���ʇ��� Ǖ'7!W���&d_r.o���lf���#�k�H���?�cVW�L��u�,T}��|>K@h>����e;�P�9�ڢ�Dx?����ѧ��cVq�N�l��7� k�!��AlT�����6˶쐻Y?�VjrT�A6sW�wV�F_'�U����x�<Z1�^J�b��I�;�8|C$[�d��Z^�e&^�<4�ȇ�ᶩi8���*M���\�Ym�y|&q8$�nnpH<�?>E���+69ha��H�/�/���*�ך�$�3�Eoh��w�8h56�^�-dF|&!��G}ֶz�
mpd �XG.�Q��dI��v�ޜ�@������p�JfA<zl��aF"�9���!��I6�V����z���<���Q#i~H��(w�D��)�h����;䔒BW&E�I�jѕ�0 )��ܢ�z�/3�����w��_���uϘN8������s����{o�?���n�{0�.��a9�_���T����	��R4d&]������� ����{��e����q�3N����	{�"��-���ƚN5P���~�e,��%��s&D`g�[�n���"eIM���kՕ�;*�\�) a0��m����;�G�f��	���.o�m݂m���h�x�� �Y}����ka>�M�EB쉴ǭ��2�7���7��g�B[���0_O�I?�	�<p*�bwK.SL`�ݓbf݅s2�ސ��i�p�-ay&�L�<أ�80�ˇo�i8j �o{�Q���͐	o�7��<��-��%Q��~{|����a)��R��h�Cap�F�#��
�k�573ƭo}{]��M1���Fӹ�ǈ/J[���E�C'�+b��4
i���6X�ҿ�+5��7��F�ρT���a�r@��z���rv���_9�Wlz֮����5�G�OJiNT�}?$d�y�\��VunزT�o�-��Jda�{����nDC
�Yn-<�~���,�v�f+�������o�/�����f���eY}߰�3G^jIRGvw�~O��O"�'�Ő��{������z?s�ц<�n%�%�:,�{a����b3As����36��^?}&[&ՕN�?�wS��7��T��w�O_�s&&6z;G!?S��qy�E��R��\R�l�~S�T���)iҗN'�2�{0�i`��X˄w �@f�a�	�)��@�b_�ܐ�N�}�Q�/�PIdK�wa���=}Q�%q��k�+O�ѣ0���L�5 S�H?��XoZ�Ttu"��;����k��^� �,���䫈��Uێ��[k��GɃvK)6K+{/��آ���a������������:ٗ݄2ZD�S��o0�c+�Xo�9�U(��1��\[�oty1�z
D�~�)t�,��]8o�cw�-E�z�������s�{�ݓR��_�^�mkk2�S����+�aD��P"3���n�u����H#4�.^W�j,b�+�V]�X���L}v񾯭?S�����+i�,�bb��Pm@W�Z����BH��h���-E��M8\�w�-l[�Yz���{�>�Y�Rab��鵁-�f+gl*t�d��C�G1��R�S���;TK��ݽ5۱�?���:������E>ݘ����!b�E>b)I�&�R����k��u?ߗz:����j�x�fU�Z��<,��k���#���i�Am?�n]>�Ë>��y/�b��-��oJO���_��F�f�����?4L||��¿O��ԉެ&�gu���8�옙w��&�?�At�1�N�~�·�[��@��j� A$�}�����iK�����%�8�@SV��8L~��"�q�$�Ȏ��7�.�"=_��sl��.53KJ�U�WS�(���Aٟ��_GB�Xw�v+=x�	�l�����H �^�e��Җ;�߼�R��Iꃍ�K+9kY��������`�s� �ߏu�Jɜ� d�ey�Qt���s�~�h]nU��@�U{2K�/Ƿ��}����a�ca��Za8��ȝ��5?���l}�;��d�\��y���Sݐ5ق�8�G")ko'&=f4so�����:�i���<�Q�	\'�G͖iDC|.�&V��`����1vӌ�{����V�t���'R��a30�T'J�������޶��1|��3_�M�]ۈ$���L�{g@���o$9��'��|�����r���y,<U��T�g��D#��u�-�&��Qc��ᄤU��3����jYP�~e9�i�jn��kd�����,v��� ��&��L��3H,qi��U ى8z�1ʛ��(vD��N�~��d�a�n	�h'�xX`���Ή(�w�![�3���'�=O�df[�W(D���G���$�E#�����K��d�a}��7<���A��I7|i�(pi9j�k��=�B֫G�յl�Ѻ�n�m� E�y���p;��a
uD"����@�R �~�g%^[�{pp`�^����7Y�;�DSaN,���T��]КS�gU47��@�X�wԡڿ��l%��]/�L�����;l�7�C�� u�E�Z�+�-*7©U�"FQf�$���!��a�25�.,Ԃ=�B���d7o,��E�NЌ���!�c��?�{T,]���e߯�i�P��"^W�q����\��M��Y9�����h~��SaxG�~���o&��˪?W*ۗ0רk�3,�%Ԏ�Y���� �\O�"(h��� �J(�V� J��;7-��(��4Y����K��9Y����<�� B0���N:A�eN��hM�v��VT����^P�Jb��Z��'d=��h�Hl�-��p�<�bZ�=)x&����}֖��Ѽ�+�2��Ź^���8mYb�֗w:m�sR�Ncyr�{z1*�x��OF?� (F��(����0p�j���Jl�^5/���}�����O�����E��=�p�+�dX%sWnO����S맅�b��~�^28����CD��;b=	dO��8����)�]Nۉ;V�$4F��A�ó��7����7iA�}����7%�
r�T�cc1&�rҴ�g_�͢ct�!�%�v�n�(���?ЊPmQ��>Д�t�v�d�kV�&�.�^���v��$����>�*�NZ[l09�#6(��r�s��4H�U��G(��p��C�p��8�w� Z�>#( .j^�^"@I9�>�k����MI.���J��PዹR_���r���=څ3}j�t�\�(UY`v�L݄5��?
����ˎ��X(�.Z��z��E��,��Ē��J���� !��N_�4<^��GAM����J�uu.�l56X%���è_c�g�U?&v�Sxӊ���B�{*�V�ί��3�'�LuU4�;
}
�'!���A i��_Kw���C2wf�!t{S�>�.@x`+P�3��Y�|7n��}� �`����ʙ+B�|{���f�T���{�|�HQm�;2�]C7�N�āT���5H����ER��;s��Z��E��(6]g뱥�?O�o<��W�0Wx>��z)�m�X�"{|͊��+��Ѿ^ф
�O7�*�x�2P�֧�M�~��|=�dI5��нA)�+'�x'�R��@��!y�0U��$`a��nKu?��+}�ܒ�\�S��YS�m���J�G���䆭��g�m'��ŗ��0q�Ո@mhj:���(�^;_��,v�.ߵf���5����@ȓ�i�`rM��A"#��_��e�7 ��CrG�½��n��QGiR��ף_Y&;s����f0�Y�>��H�9��G:Pxz��� ���ֵ����K&�]9�_|.��?�y�=O�-���h�y�}�֟ɨ�N�:�?9�;@�r�go4K�\ء_���y��[�k���+��Lˊ+_���_��d�;�"��־l���@�'�
��h���c�,��%q��Kw2���BI7z�I��	���iO������s��,Gä5�6�T�la0`��3��k�v�60S1����]� q��/>Bj���m+�N��!i��WAhtY�!|���:�c�{u8�m���"�r���� _��8����ze� �\rv�T8���b2�ySܛ-ci^/^�|��������g7��W~��='��;��7vjh� �ӑ�c0�_��mV�
f�\�����'cxO�:��^����C�I��(OpRq���AZ��c�:�҆����>��G"�Xe
19�E���qj'w��;�ĐD������ [�*�S�V�5ue��2�.����,�h�.Dwpk���1!�#_vC����@�|	���f�,�He�nS��?J)ܲ��0,D�x�Nd�� ��'v�zb��G�8kL��b)�����������R�_z�r�ġ^����1?=�VN���u�v���S~̼�S`��d��QC����'���I����ˮGki��f),����@P�֎�$����=;ak_6b��?���g, �.��kڙ�Y��Q^W	�������"�b�,�@ҥ�,RQỎ�<�T2�"�>�
�A���v���=�a�U"�$�UuU���K|�>��<6�٫~c�*߄�_���=-��;M2�mk��W������)��3W^�1/䨹8u���<�O�ri-chP�K�hV��~-�A����`f��s��k��-��Tv���^�1�H��N��i&�D���� �$�ZQI����N���в�c��7�#�(`�uN�H���]$}t�)k�Zh,<(>��f��T���)\y��z���Z*�"�<�j0��!%NrM��c �7q��j����ʛ�mА�6
�%0W�����<�J�����nQ��W�r�����|�\��S� �4s���צ\7�1�2��=�q�+�8O�,��f��WK�����Q5��?bӱ6��BDzo��*� u+�3Ʈj"�s�Bzp�Y֌�@�A�Vy�جH�)�_���r��=��+�/݉i�[��x�ޱlW9�a���<@x:+c�x�A��]���^Zx�{ԟ�P]m1��������K�桨Z��b	��6��4��5(zR)a�X	3-�X J��]������6[ ��gT����+�{��:���R�Hd�9��"��w�r�0ILv*zw��3���s^��sY���S�%ȳ�a$�FY����B��1v���I2�s|6���=V��ip���پ�Y�;���� �t�h��ȳ�#�fx�sV��{��<k·�?�~m��Bw����(���~�l1g�0�R	?F�:��ѻO�	���a��So<�<�����؋�)�z�`�I_��]�x�����,���p,h�я�Zx���J�2����SQ>YŢ�+������%��buo@������Bt{�Rϳ9�9�>�(4[wB�쪺%�J�d�t�m��gA7����G�LO-����işM��y}��ON���ݐ��]���Qz�Z&�{��q�'�FJ��, o�{3���0��%��EU�͎�)bs =%��!���e� ����4|����Tx�ɚ�_�9 	 8}�ϠT������b�P�S�S"pA�X�q{�Yy����xCӻR5c�����.MoB�;/�\�m}b8ʷ�����S��)u���Պ�-�n�TM���Yjl_���t�����S��>�@e��VT�v;\z��S�^{&�,��̙�$���+�v�l���hU�=Dq��7�����i 
�Z����-o�Q(�o����N^u�|?:�f�$�C�[��B;���������Py�7�����Pܡ�g�^�8�m󳋱��d�h%��n�y�<��=�ޓ�g	:�=�ڀgg�t���%�K*�L@1K��D(��'��y֙[�F�@Vr�d?��B��a��O"�Ղw��&b!�����zFܾ���;Zf�p:{�������\���rm��6o�g�M������ 9�f$?���>�c�q�l�U�f��%E
s �H�E�I��xoβ�J���8=��a�ER33��9#eS2!u�}o������J����:x>����(2&�Mm�Q��Oφ�`�da,�(U;��y���$�/Dn����1�Ӟ�����^�*���މ)}�8�����#vx�=������;=h���&y|;���Y��3�"�����&�iP�ߺ�[��GRx���EKb��8�f%�M�'�k�a�Æ��8���pa�2�Ġ��z�,�
j�-?��-$�4VD�&z�^e�a�f��`MC=;c�P�y���G����`L�^���|�}zV��^٥Y�)�ۓ���m��Nh
���������iG5 �� 2���ý��1���kܘIUZ����mx��1Y�r����!�k��?�cB^�g�_Ԉ3Sq��v���Wq8� �����P��67vYt��1�A$����;v�7;%|�9�J3��җr�.�y֣�%�Ḝ�/��𨂈�VA&���k��d������-C�Ak���ѡ����]Ŀ�$s"�4��eU(C;�]��dQ��"��L�E��y�~y�ϗV�
���M��_*�!��˾�Ϟu`�f�]z�@l�m���p`�������}L���S�҄�a�A�����!�a�@��њ^���1c'����~��y܀�n烌�n/�u�ˡ���9]r/}lo4C����|�����]��NG�,�6�痔Z-�u.���xB�6�My21�ڼY��K?�����(S���<�J�2g�] � :-��b|�v��F9��=��;8�I�%/o��I�Շ���Uh�3a��ܯ�E�u'�E�Y��n5N23�f%;��I4�
�����5n`��
�4�Hӷ.�,�qN�t�25�+o�{�5�.��U�n���7�J^�C��#���ϖ��i��4�lk���=O]UO��	��	�ࡉ��ʘF����Xc�ڿ���W���G���X�rU\ �Y9hA۝;+_{��N�CM)�����:x�T;���J����ژ�6_č�/�fP�*H^�H>nQ7�vLxr�eE5���.U̔�+Q_��V5N}޻�&���4��o<���<=R�ٝZ�i�G���j/σ��P��oŒ�ID�@�+�y�����:�=�f��i�"��o�(�t��X�?��g��v�Y6�'�-X̘��A��d�%��X�hw��C"�Y*L�\T����� �`��eQ8	9�Kd�p�)a���YdF�;�f��sw��~�a�@@`Z7#	
�I���Ee�,��+�xbP�PE�`��B"4Fٽa��گH>�rİ�-�ewZ��d�n��Յ��=y-��[C/O���O�4b7H�|�⎃���:w�O$Og�C�κ1��I�kZ�I���^vs��G�ФB���ְ��/�@���Ru ��sR�[�_1�ڸ���*=���%�%�"���ۛTQB�OW3�NJ���(��Χ�����jZ�jZ���C$��,Y����@�U�:�6��ed����AE�>�C��28�&���}ssx�=!ٚ'O�������ob=���Q[�N���З{{�X9��O͓����zU���P5�@A|)��%�{�b��l�|4�7iWQ+�.\ϟuI�ȭ�XɄ^���T`�ޭ,����=���IQzDH���N�kȆ���̉�0��;�� M�Y������p�5���>��
ԭ���POK��F�|����V�n3*켹��Y��G��I���k}� An5R�"3z��FL/��r�E�O�3!�P�3*��Y��90\)�u����Xy�T~�|������$)_x��5��(�d9X�@���S�7�<	+��F�(������FDM��p��|��㯥pc<@j�_/�:��7�4C�~"�b�C���k�ƥ�Z+���iX�5J��}��q��,w���X=H+�-/h��6`�Ω���%I��"���C<�����&bgz��R&�5�a#�3K��DPK�9������
�P��;qg�n��0��iA%:�wns���U�尼�H !�m���S�j�0F5I�Fy����n�(����&�=�\Ϯ���}�k������`������N�ʶ!��F\ӏ�-�)�.�D�V�6��va^������b��+�X��^������4�6�B�e��|E'M3��� �͔P��K�tE�ǆ�܍L�V٘�%��F�;�y��n�l������$�dDvUr�1|�v���M��Z�?ۇk��C�I/�KU��d֧#�ť��j�:�%v3H�>`M�˛<�;�c�bVܗ��X����z-� G�/3����&�s�R�|�	;LL��W�/�����Y%o�����[
A�>@ f��B�W��'Wˤ\��gZm��Rh�To�~�Z퀎eX�}ׇ�����l,ĩO�1��H���K���b��|K09��y]7 xY2�T�����k�*.���٠#�����L `�B����W/8?���"C���������`�Y��p>7�Te��HV�ݔ�%�ѡA�l�Ď�h�ӵ���f*�	uu��%&���L�@�a�H��$�el��x�ܩ 
:m˒�k�IX�7Gl�f�����9C�K�~�D��<ե��i3�T��N��5�����qZ�͟<�e�t�{�YZ$�ͥ"���*�E���,����Ixh4߻I>�5 ޯ��$�ΰ;�k`��|t��3��X1��!��j�bo?�B�n�S&XT�_$�c}Z7� ]������D��$�ǯ�a>9M`�> ���4v�8h�Ҳ󸦞�W�et�O�L*~GJ-:��؄pi������\����I/�W�G;xK[� ut�G|�t��f�fꭜOܛY����������E��Ժ��QHs�\���8��5�<�c[�4�d�F�+�̰(lz���b��"kFS��@�ɕ�3�o����-�m��F�vH#�+Z;���\�D�,J�9�X`��9-��דwШ<���(��*��D	��r���L����8���V,�����n^��.%Dn� �Ba[�E�4�}n5&�m�P�W��G�9 �GZ+Ǹ��mR54Y�g�苈/��y�c�"0�ND����.��t�����V�	!f�X'0���2�.��N�n���G����9��i8�[�� 2�� Db���k�J9�̮�@R�����9 ���W J.[qr
�a�c����,�����aǆ�xc�v��ET�|�.r�ﯺW9�a�3�5�t�GcXK+}
1�W8�F�RJ\�&A7�p�s��G�yG���4�鋸e�T��<Q�ڴ�CX��@*~�>�f�/�w�^�_~nͫK����*�:~�T���L�J�2�$b�P�V���$8Ulk�5�^��A�[��Dq�0wF�K#e�Q������6�/|��T�w��"e|rE+oD�ނ"������ �k_	2�ag{ic�R�[zek �\��Ӆ����6��H��G.Ʒ���0dq�Z�Zj������/�� ��de����8u0�E�W��}�
�1%�^2�R�<Vf�x��x;�Ֆ�6�����*�t�.�$���vZj�B��^�D)A�*M�z5�t�Lq12�:˻ďPsO�5�P�࣡ɵ\��ri�.qU�1mJ��ﯞ���r��������\~]iG���lY�dY��� �go����#�/X/���̙8��[jVC��JUL-o
��um���Nf���N����v Y��3^���[�m9��E[���au��p��Ӯ1Zj&R�����O��c'�G�m�������O;?�%��g0�ˠ���ļG9 �]�N ]?���I��FQ�����"O �ۢ�|�����>���B�r:EiuS�%��Ndwg
kJ{���EL�#��{֡R�SX��)�+�p3<���(.AXB�O$���8��A��v.a�����>��>�1��A�`D/w�(ݘ�h�Vti�4��z��n�3���n▙q��3�	��֋���~��-��ɼt\��G���F�n���{�X����=s����t���R�9.�	r�}�'0���D�m P�I�N�ێL+�0hJ�	fhk�V�ɇ��+OX;.�13D�I��H�s���=�Phh#%׶�Ak`R{��M�Y���K�n��(�mR8$,�>������<ͫ��S��tiB�<*��
����=x�=Z������P'x��Y.���*)��lT����;����n�%3�̓4�x;<lp�)~d���5��qz����st���*s��=�K)��Qk���]ny����Pϗ�mz��l8�xK � ��@0�G�G.�P���͚�i͕�ޝC��#��-寒rk4%뗈kU�0�i�BВ�b�gZ/��rPs�s}1*����� �y�D�J�>H4�p-�9�[��w�� ����|j L�hV��#��G��B�<�QE|U���͉C��J���T"�RμJB� ̣O^R��H�B��\�K��d�:����ޞ4-�d�|��"���V�:��Mۑ�g�h�������guޯ�zǉ2I�BC�8�0eۉ�����ʊgq:ٌ���wCj�Q����J��
?� �bd����14���:�:�i}c�_3���,�6����r�Ԗ�+U�QԜ���8�ѕ�L-�W8���R �sD�x	�E�ڽ�P{��*��Y6���YV���C��C7a�P���F�m@����)V+��_C�jp/x\
� HM�V6HD��kJ˫<o��/��J"��"�6Z?�J�%Y]x�YYiF���$b��#�Z$J#�6��󣌲EoY�@;r!�� O�g8��sy�Ӻ 5�7�m�Rh��Vn�J�_1�.t&�s��*�:B}J��<��	!x�(Cs
􏔷,�~n�(�n�?�M�as���'�Dp*q�%�DPՏ(�[_m��GS��a0������5��q��e�/M�,1�ʵ�� N��ʹ,�}+^qY��5�a7ovvV�	�՛%@�%���k>V���B:����>�Jo�p��M�~����	��J[8po:W��a�]��:�~���"58��c.�$3p]W���ϭp�<��&[�ZQ(;��9&��h4�W=�{��H���E_$m�c�`~���Z���md�uG�e��iJh~�%������bd�K���LRY��Â8��������c��`��ڊYat�R�/��ˢ��P��Mģ��~S6���K`a�_�?�ߠ}��/XV�v��.V��]�>���@l5��Μ�+#�C�Z�s���V�~��"u}��%?�g�}�{���WN�E�����l�C�Up��=�Ϥ����s��-gxG���fMUb���
F�|-�:N�@�}WW��S��+E�
����g4(N��H@��q[�6�QM�ɉ�'���o�}
���<�=�7ǝ+�u�u�X��k�u��V�o�S�<�����.���Eͻ#�w<� UG�)Lo�9��M��1��1��͙3������	9�q����zR.f��GT�@��3�������N�/N�,}�f��VB0W=n2�>�U��#�T	+��uZ*:���q7�0�1��Ydu���vD��7Ұ�bGv�A�9Ż`���]ӈ���ʉߌk��L�!T��"H�Xp��7�iC�QA�d�;�3���TK�f5�İ8z�;w�*�rr�wM�P�"x̙JQ�/S2r�՟C*�l:�{����ͻ��<����dp=nl�4ZS@�:�j2���|�E�@��qi��'bLs���v3E;J�CS�\\H����_��$��0v��.���N-�~v13JT�0��)b��z����A'~B6Ug������H�����+�9% �=��:��>5]X�(oB�-Zd�ݢP��S�csR�����p��Ee�i�~#K:��U����ڪ"�{���o�{_=s"�W�H�)���Z$��/��f�	��t��ej��N��
�<�a�s��)��ϩ�?����L>�ۓ�J�����p��&�fdn�#�|'GZ�#N{Q�a1;���7=�F�8~I
�X|�� �0X��]�p�P�J��G���%���Cj�rG�@BK��V`�"���v-A#nK��E'��B�%K�桪�5��Ju�c���V-��CZ�0���IA�ޅ	U_C��]Q"Q�*����4���U�#���*�{�2��������T�ߋtknP�R�yڰq�����˄&�(ʀB �x�=�5.�z�hc����e!�$����	A�3��؜fD�@ß
���	_i�r%�o����]��Rᛩ���U4;�(&>B;{1�7�s}�2P@$�q�[����7�/C��('1Efb/��-����3� �(h��[r�Ma\�D��m&����^�����t̎@vN�r�`ib�����E&[w�DDʜy|�z�4���Zѝ|�-/:�+߭Φ-�BTT�-��Y�+2�t��i$cq,=Q=��w���x�� ���k�%A� ���u���\��}��Ye{�Cz��R���6�� S׃��әVB��k��&}�o:�_R�䩦�x����+W�C�ƻ�:*��9�qX�f�I��M��� ����L�W9���M(���@�;t�,6����P\pm�z�l&<�5�R���{�0�ru] \��)��"�ϡ�:�ɔ[4�ώ�S��,��-V]Q֙3�S�Y�k�H�]$Qo0Om^�/��rv��X~��rb ;�ֈ�[�ۖշ��O��Hf��"�Q3���
s�P�5�o��$�s���E�� q�3�5�{:��@�n:�G�j�o���N�7�V��g-�A��W�E�y7�a^G�+n?�	t`��R�h8���>�]ӐJU����a���}� 梖��R=d@ut��H���Yl+���6t�6���mf=�V�/G���
b��m�R��E.3N�]������{�{f��5҇Q��;�s~Tv��@S���"kAA��(11�a}�q&|1_�Wwpb7d\��ǂ��dXK�o5�Y�����)�A<������%������*��ҾD����N�d�-a��y�e��^K4�i���,qfY�x��,;{��*{;I��M�y�Z�Y�s� ����h<���G���@�mA��6��K���~Zs1����O�(8�����5��In�Ϗ�f)�:,��u9آN�L���M��X����p��x�o��Q����Z��m3���f�M�-�B��3G��ts���Q^*�]p���
�쑃n�B|��dy�8_��Ot-��
2zMk0�-� G@�tw0��o�)?��5��Bd������=ᴫi����󽍡�ֈ�w4�ْ$�~_���j}�[���c�(A(���0C��G����c1s����,���u��9�dڟ�	dZ8S��M�~���R��\R�����I������T{������^y��Π��+,8��Ҍ$DX�
I����+2vJw���z����l5M�X���������*`�h�!�z�7���<8�I����
�����(K���f��Ġ�wE�n�ASN�$^h ��D��_�-!Dh%�� IӮ8����,D�9�_21�^	v��"���Yݐ2�IQ��R�r��� 4L�n����չX��(�CFTp��g�L�s+8�ʖv����?�rwj{D�C~�� 3x��	�pnH�~C�Se�V�/��E6�C;=Nб�"'�.Z:�i{� GM�q0���*��%�p;�'�/h�)Dd�����5��͘m� �M��;�~uD�nv^!�q/�4ҍ�*˃8�B�|V�&+�s��`��r%���u���[�Gp��?�A�� �*�%�� ,AW.� 7�>�^s��7��+�g��;Et�LS����M�� B6XZDc�N|p�
#kJ!P���"���풞78+ B$�-�C�bo��8��|p���4_���lj9�9�M��R�Kث�	�lP`=�
T�|�h<W�k�kI�=��(�Pz��7Sa���״��i�v�/�%l���[rPJ>T7$(�Зut|�juyu�YNl�,prCHǢm�y�����#��+MJ(�����2�rH��:ܗo�;�	��9��p�2�4��GZ3�Cw�`2�Ɇ*�>���d�:�;3w�����M�*��^dgr8��9DA�	�ؚ#{�ݧj����L��9:��5۸U�h3�Եd��5���ӡ�(���4r3h���oH�m�w��aH�6��(��$"P���f��K.��ÿ�Zg��=M0���M�D&���b�HA�n�
��I�.>9h��1Pj���T."���Bd�[B {&-J��/�x�Њo��|~��Sɇ"�pc�남 ��*{�^÷�+a���=�	�4��uJ
7���/k
�p��;�\����?�4��q��o�Q�4K2$����5G�=Za�N�Y�_�bq����D�_t������V"�c�׎���?M���f��ǂ�5rƖc�u�ZP"���� �aT�R��-� f&�QÚ�fǵ#����Y�"���k�tG�[�/��<}�e=��6��iXQ`M�h�:��$�XZ�4�MN�*��/Д����X�Ba�/:Z��&�v6ܫ�L�V�:D�z��3�e�Y���9�6����6����wJ�q����,�`g�5c��u�sF���k#��3���I����s9��D���%(o�a2FB���Hl��Ɉ8���Qi���+����y��~[��8�/Y����: �6Ba����)>�}�'߿=�ӷ�1X}�^;گ�Gfj��A4<"Y���`��8��b �8Tcՠ)��+%J�����p��h3���r�Lj�jr	���Щ՘ʺ�ünx���D��#j�����Ԭ�SK���]�r/��0yFj���&!������.����cN���$X%��zg��� 2���,u�?b0���9�#V @'��V���X��"�0Cn�	�xSiEoe���">�����b�$�MUڌ���p��T[��JR�Y�Mx%�U��yK�*,��V��mFr/Duf��,4믳r҈'��w�� }WKIB �)xX튭�)�(cSnI�wL:����-<��;��]JOUm� �N��7��P�����6o\��J�>]�z!3eR��r�`%S���i��8�>R$���8�v\",w@xǑ�22�'$��-%��ӣ�r6HD����&s@�a~��x�t#W����o�i=��m������Y�ٟ�˥`K�l�f��y�͙�f���"���"�ݷ�zN	�>�0��E�PV�p�" :��̃O��a��r�bˍh {00O�)���@y�q2��x���U�a� �8���]��k�%j��&�c!�i�-�_�C�x�.�exs[�2��g#�~R�e��������BbW1�gPHb�����~�kȟ�x�?�a.HznN���� �'؟2o����n��",!��3n����hC��`vL#&O� I�;Eh�"�&(�xe��&��Mt���jr��QtB	v%����XW�.�B1Ήᬫ�5��y0i��*���ܳu@�"-�3��pZ�NQ���L���5��u')��EG�WEַ�4�d�Ӄ��ۍ�7+��3hS���㶼7��;���w�- �N��s�i~m�w㯎��W�Ò��d����f��J����s���d��[%$����sy��R9G�
a\1x�!���=����L�/&	Gd�Z��1B���9 ����X��]60��%ʠ��̤�I��Z�ed9@տO3����O�ñE䆂�%�q�cݴ/Rп�KN��zo�F4GG�l4���;�Q���AFqCl;���S  �������u\sDf�U�Z�$��(&����L�sH�������GF�@@	�e�ra/ I���L�N�uO��S�\��4H'����B���eބ�P'0�k�v�D���:fw;�l���$�p��;�72a�T��o��bc�A�����}��	��aNIGG�?�����
L��t�ˬq���vs��LUG�)g�q�d�q$t�5.`-0�p�t~�	~�ףBPɍx�+yy�y��U�����a/���1�8���8�^�����ž\��?��r󚆂.�]?���g�Q��x1���z����wD~G%�S�y?;ݑ�XG���7۸�������O�	���f�z���ZN1��t�{X]���p׌�g}Z>��V`��6�P�䟨ll�N�{PN�3���j�)�P�k�A���\������P`��U�5��0��[=���������]���Y? oB;�2�u)�(
�q<d����[e��1���� ��� ���8��>��x��wW�@��N������C-^<�d�tJWks��x�?�$���P�>�ۮ��������J#��	T��s���d�E/�^��=~φ��(iƪH�AY#�����+[�x�_/��`��k�J4sZj*�|�$�N(�pyͦ��z���pS�ݜ{h��|�j"nUµ�s���&�Ǯ��1-�;��z��Q4�"�Z&5�i!�V���BZ�h�F�������)��	3��G\	��}�z�Ω��W�0Z�+ч�~�S�|��^/������Q��p|��}�}ه5�tw��P�s�}h��A����C����r�f�C6�t%.u��x�����v�����*�'�Y#2?��Ρ�|�PB=� ��tqyBNz�[�=�QTQQ{���lN+�/��%����\W>	o�AaK�_7�d�=kǜM͉�#��xZ��>���A"4�rR��	����ٵVab�~��v*�x��)��v�a�-�љ2��37�D&B%d���j�"arؔthm�!��j�`�oSp`jZ�FF�r{�nn���L5c�Z���{s�{�m�X3ZZ9x�f@c�@�s2���})Q�	�����$�$����ބ����p�%������j���k����F/��Ks#��� ��=� *Y�Σ�h���>�~#�k�o�W�f�A"�`��W�(=�J������q{�>�dp�7v+�?걖Gk�v�nrgz�vdfhj�`pk�9΋`jE�lg˿�VI4�V��ّ��Go
U���/�;��7�E�;�A:�n�)��s%�B�Y�� ��A�g�?N�%�W,���3����b/�s���MT��3`3�ݩnN���`���q5򩘯�3f�F�Jѿ���[9�A��;Bp;��*�#�;=	�C�<a��$_�F��w��9�J�[$ߵ��#��6ґ�n��P� H�U@�V�mN��I�K���LK I-%l\��_U,\������i�Ec)�O����ז��r��	Ec��A��Mڂ��X�DA7���=0�a"�a2k��rf�F���S���F��V����O����л�[�8yOr�}����Dr���
��E mvI�w3Oҹ���$xTY�7�X��t� ��d�0p9Ǎ�xڡbaDO,�XA*!��|WEU���Z��N�u����7,�I������Y/�I*� isj��-a�Q���h�E��K��[�n�M-D� �	��z���/�o�^�`���nO
4OM�
5�k!�&�-�u1k)<ۥ2�CX�D�E��Tv�O3[���()�Pˉ�b�@��"���jq%�� M�3x64�G�f��$G�{\3D4��ŗE�s��BD�qC�h��1Q���1D���1�x�ZE���.�MH�M���L8����"�p�g��`T�S����<Ӣ���#)Y���u�H�1����
�E|�$����ΏܞUAXf��/:��O�v4c!��r��8�J�� %b�����"����+�S�Jn��?��x��9s%6�� �y����K�&5Jl6���d��9��w%���l�6�e����0l�.]fC���r�A���p�Ҳ�/������)�`&I��`Z<~��������O��Z��	C��^�h]^�.m�I��̻p�	q>���r�Ҏ7���O��4r� �=I�����Ɩ?�M�4���v�*]��CU�Y�/��9X�ѣ�{ǌD7Z��\1.w6T�Y���h-�� ����8֋�L��#����/�����@%��x�c�����"47�㬋~� �<��p�&cy�2��g\7��s��⢳�6���?3�-��R�S=D)�ޤ�1��}��\�8����E�GE�+N��M�uT��y��}w��'a�hf"��*B5?�܆��[��V3� T�����Y&� �}�Gٸ�V���*��m$����q2��P��k��w�.<��G����89�%e1:%���h~9��!���
~}�&�KuP�c3��>Dl[1�������8|A�偷34��n�F�ۖH��_��*��כ&��e�J���}�T������m�y�(SM����U�s#/W��9&��C�7��j�O>��H�����|4'���#)W�4���n�An֠��c+q�:�Ё���a�'�,L�z�H���P峳(8 �d��:
Q�؁Z�^�'0i��hRظ�ױ�,-�u������i�'�,�Hd%�Ed&bl2n� N�٧����mh��1�&��$)eފZn�!�"?1�!��nvBp|9�w�x�o������d����3��{je6�J��l�N�Q_����j�,��ȈNO�T���kCdc��|��B�N�t�)�gc����dHղ9�k���Wfn�>��&�c�����	�bp�b��NBuz~k5�ҤZ�������Z���r ���0��Q�tb����1_I� ��J��K�e��,�J%��Ǆ�p�\�O�C�����ءZ�e�o��\00�hv�S-����U?M�&��.Y��B6�D� ��s��l�Cb
ܘ~YG�r�7ɻK�_�t�[��V�S���X��C��/놡��U^AHFEP�l�Z{a�����Fd֎����-@ң�{�$m�,~�w���L���p=�{�]Z�ɤCu��#?R/�;9"����5�����(J	��V'/�-9c��{�Є��-}��Z��(A�q�.�����+��f�8+8դd]i��︥(Rna ��SΑ�����9U�t��zo��I"��r)k�}�W�t��}FM��`�!tq�4З9R<��)�-�Ӳ��7��|��[��:�m����ޑ%}Éϕ(���=��H)�l�1d��6nXnsSXk�����P������l$�tM%�W�~/���0�m��A��X��!���b܌r���B����Iooāj��2���)8W�VO�ʽ	��R%ܱ�\�������w~���d�j:�?��tLvR�Ǟ�d݀�9����3�t�I7w=��Lv��W�Sp�?�T��.F�FF::�(��N�hu �b���>�����G0]Z�nN�Z��Ԕa<F<�JBY\�`O|d��Jn��<�_3��1�� s_F�����\��.d��=&�I��_��U�p�&���� ������k�R��ӧ�)�\01��}�f&u�X��4�z���A}n��m�𡛎��b�P��m\*�L��Ù:���ߟKR�蘉Y)38��qW{�X��7�w����m1��]� @H�eD���5���<_.��?ߠZQ��חH���M����&����C���g��Cn��g-��E�-���D)q�@�.�������
2� ����P��x=p��8[�jԚ�w1��ف�.��M��`��А9�e���fŵ�ў�p�p�v����E%J��W�����z��+񎗕�����7��Y��9e��7ձ+���c��~DB@�-0]�����Om�J|��TKc��p
B?����Y�wk�w�_�NT�vO��@$��.sR�k��*FV,	 z��+jn Nws��t�ٲ��!��}�+��|E�%�X��h��\fJ��B�fDC�$ �&X���W�P��
ے �6�	���Qո��^la|w�Y��d%y4���B���F��d��B��u���˦�6 6�D�^����*&}bZ��%v`����S!��Y�LE�=��`��1����Mq�o��a1�U�3��t�
Fw�
�=��'��"�.e�Q�k��������FyM/��پ5�����aD[FHL�f�tJj�9���C�jL\L��
�`T�<�vS#��ԥt�AJ����sM�|�yU�.��F���f��><�L��5��V����8-�8�L��N�E���U�YQ�w��'��Mz�����L�/i� ���<��H��� ��@<��T�Y�*G{_���rM�4W���D���b�=A��u7��5m��'�Yf��*;�#�A�NPXg�h��I� ��#M��� �!+�TK��ŶL�/�E�p�	��ĉ!�z'm��⩶f��kN�n5d�jB�Y�#R^}���%]�/ǭ�}���B����S0�Ҧ�]ĕ[Z@�Ej������])�_��ߠ��z����!H�"�^�����i�l[>V퓹��=��g����Qq���0��e)�7Yk��L�v�<�R��5@d���1f��/�f�����Y?��w���gͨ�C`S���ʣvc�S�0���,�3WIWr�hAw�_���]6��RV��u�)����?)�/YO��ViM����r$T�ޔ^|�5�R+�lb!��:�Ī��2;� 9L��>v������m�9�*��%#-�0�P�D���E�_��0),}h]�=��q�����[��Gc=��[YH`����Rc����4W��r�H�hʍ� !%4Ǹq@d�hu����U�Y�!�!���5��/�>�[䑺{��m]���
�`�%��&=i-d���j7<^&vm�3�f��9�)ٗav|J���9z���W]˸n�~`�tt��Q8=5�%�BCi����hk��B2F�2��8	b�%%.},�x��b��&c$� ׬�F���B������Zd�P�[��l��T�b~Q�ą`�"NCn��"�������JX�#!��������W�>#XO"�c�o0yhvN����'JDP�yӫ��x���0|����zQi�s{��L�jEh��͂��^9�I�tW(uOH�G0�jz.H]R����v<8^�,E�{J��V\Y#�Пrj�g�r���Sef`H7�Z���"�0�2�m��[�g3�,����q��7�jM7�<���=U�P�@�#oWc돴y��ȩ��E.�0[����&% N]�ʥ���"��r�2h��
�6U�c����tx����<��T	6�s~Pl�u�v�(�;˯�����s`�5D���J��\+�g���M�����ci����Ig&m�-inS{�=�R6L��Wg�s��C�|{i��2����+�M-������ae��u�Uc�3��M� �Pt���Q������aٱ������yH���Z��'{���N����V����A�<����*,����^E�;ȘbZ�<�_�{�lo��i�9xAe�|]JA�jgf����t��C�b���
�L.�̭'�����紾~֦�4�i_��8�!��p2��c�\�~��ݤn�&q'�@9@�s���=�������*[�F���"��V���ߒfaSM��]�����^;Ç��/�U�V���tS��I҈��ͥ�jH�o�23�5K�7�Ew@�:�,N3���B$?��͓�����ԷH�R�*���׫J� uB�qs��V�x�B�3�J˴"DL\Tf�d��},O�J�;N�~o�\D�XGfzO�(Jw�0p�\l����U����?b�"��Φ�~�� �.c��l�R��&��c�KX 5[
�Jn�cT�`2o24����Y��@��"�Tګ�q������	\@=C��#�X�s��
�A��E���.��.W���[o������h|�sO(�2�å�RW�>�[��68g{�,�ԑ���ݮ^�k��/�1�Į��@E�ID��K?�Q�.
��.ش ���b�#?Y�1*�W���~¾%��yF�j�Z�A���`���;��Ƿ�k��,|.A�S��Aho]/2���V�OKY��@0n1�����˳ޢ����3ا�m���X4�&�.����j�Жn˹��(�oV �ǆ#�?�7�	�r�6z�G�$��D���s�����6)��潎EZ�+���_S�)Wu��h��i-�-�s;��v�<5x�w��n/{�6�j�	�l��A�����xc �Z�u������l�'�Z�`��Q�ъn�J�����!�nEj�T1��J�p!�j�+BmhD�n=�!�H���qĮb��O��E�5X F<%��w(b
�ֈ{|N]�{�ycW� |˔`���H�1�a Bn��k������}B�^�����H�P}s����]@���1Q��2�D�z#�0�)��y�tt)Pl����[OɎ�0�j��v/��̝|�y\�Pu�+p��}Y�nG�.�D��S8ya�D�Q{������a��GW�����c��P�iP���O��~�C.��<�#���%C�YXqN�M����"F���Γ���ѧL� �CgY9�Ոf�j|C�P���=�{���O���@�����h�����x�U�`W�u�� �kQ��ɤ���^��O��N#@�mE0�/�C�e�~j�
[������Үo�ɭ�]�	C^�!�v�8SK�cN!�P=4�{��8���M��й�*�xy+Wѿ��Oփ�����+ԁ���fR��M+�AI	_��Q�:��E�)4�"v�G0ڬ�V_1ً>ݮ�4Z��ah�W0Vz1��>cv�0�f�w����x�n�t8���
Q(Q�v8��B�#�N�������0�@m��N�yR^T�թσ\�q��Á�9X�U�܆\[s��_�2&i�~xE�P�aX��bW.��,�N���J�yl��G>c#�=ի�:��⁨�h ��%RXXe�q���r��1<G��G\�
���sqDr��k�3��c��/ˆ��A3������1��O��WMFC6w6ƬL{u6������˚�I�T�<=Ϫ�/N��Z��iR�	���|��gY�l�0�k�B�|�k-c��đ�-��mD�Sq�ށ)�����̓X���.�*�4<5LWw�v5f���B�i`9�K�̽�� ������?o�$��L|^�:��&ή��gĂ.�	��t����9�0�5߯^��#x��e�MF����<�{Tx��ʎ��/��H���Do��R�+�Ĭ�&�}!K0JS'w�K��� @:[XJ�`\��>�P�b�8{<l�p��-����:a��l��ʈy�O5�Ή��&�9��s�I�Y�[M6�nR9�i!�{4�� %	�����I,!=�a;�:y��~�[��9|�-�gv�AܾH�y�֨���0���{:���X���+F�#�#]r����Z�0��'��$$fK�ͣ���'���ON�&i���Aȯ��!]���(�{F�� ��T����p��rZl[��>|`�W�x����1�ޠ;��g3K�7EL�H̏?�N�)�怂��榫�{d�ӳI@�ĵ��w��}����K{��y-�h�k���>�Z&��֟e��-�Tc/�K�h�bIO.�;��uB��(�	��Lb<�~>6���kU�w��bA�3��ji����.�6�7 +���~k�9�h9����E��rR��<��_'꺍&B˱}d�Q全;�T�4�`�L?�@�ԪME	��U�*|���|G}T���u�s����BHe5�/j�D;>Q��2���������qm�o�}�=�ą�]�O>8�vT����@�&���4��Τ�ɓǘ�f�/9מ3����Q�*��?N�N���pF�!�������f�)�S����O�6:��y&$}4i >�<����t1~�i�G��X�/t[a�����a@U�����|�ɹ�a��"g��~�*c��TCG_�SW�LW�=�Z0:���s� V.��<�o�^�����1�,�6 9�|�f�9�`f�E���[<ДY��l�#���4�>C����t�@��`�5Ci�<�n��x�J+)���J���Yz7%i�۫���N<�����?���`���ys77��[Q�(��ȒS��	����`L0sbB3�נ���0��ި �J��vO.�+�y�������?�Q���h���d[����CV��Ե2��:���}�3��Y�� �������0��sUL��Ȍ"p�A#�L^.~O�oac�bRu�G�^xM��E8�٢a��ۭ'�T>g�aķ���HQ�_m4�z:�q�Ar�o���2"���MR���Ҿ�Yf΃>s|�.Gv�;�%D �)�����؇�V��%\�%}�@��~!�`^)��zY�=x�	>	���FF�xإ�&>�(E��ވ;N��V����Q��u¦	Zp�} ��k8Q�c%E��p��	� �E]I�����8��Sʛ�j�c��Q��%������7����h},���C�q=1�ܹq���� �2��]rU��'��=hř�SF�^GV�/x�����.�s����c
�{ɉ5�]\��JoQ&Z勌�<E ��B��=ݾ:c(�/���ʸ�Ƀ���\���G�i�o����=D���@J29���4�.��T�GF�E����,����xë5�o��eɬ�喃K�u������uZ�̩�<e�=b�|�7S���-9?��Mޜ��}k�{�2lYϨ���g�C�c�q�GF�p��nA'�$��-U�-Q�k&�������qZ��D�O	9�V���^>�!�s%�$+3ڌb��u��Ls!f����6٧ß�괒x8����&{�|M8�A����<��)xu���SKIcN�ַ,��]3O��O_�(��\i��Πm
Xk0��v�bw��E �4���Ԭwd�| b���s�`;I/�i�ᠩў����� ��3ӀU�yg{�iH&�\�x6�����dv8�}���~�Iy��	��e�\r`�9��d��A"v|��!3�ՎBrc�[�����U�`�x�*�?�����#֥��ج��|����U�a\��c�-�?wz��Ǯ��
��^�����w�n��+C3�3��%:D�z��q�?r
�E�[U)���(���$� ���
&�Ğ��"d/����,����#�v����-�t�3��B�R�ؠy�g���l��2�cAK X.y������O�ڻ�����ʻw��y���ؖ���#U��!IŃ;�`�V"�`�5r��k��P"�Mb��$;f��H��֜2��Hce�E1�_����R$6���8K&Y��o�(h�ΖX����I��?���e=I؈K��I�0�:��7�U���.��s��Htͪ��EڎB4����A���9m���f�}}�$yS���L0D�����+�B�>��2�g�h]���~�����1r�����h%z��i��0�|�db.i�r��ŷ"����ۗzd������Ye�֨�q���Ht7��J�k�9���}�c&@?q�^m+��$���}[a�����Q�e�i?" �|�bo�a�����ί�l�p3i��WSL����Δ���<����$Eg���B�3�-1�}�g��y8�~����W�.3,.�,Ih�!UE�d�1���4�������Gٗ��cc��S�(ZL�d���༾��}��Q�9���7���}�v+4&�B�W��B��I��L�Ug��ZTe�we�FiC]�}U��Mg���<���� OA���0�{UG[�B�WٝI����L{Z?�
��ʏ��:f� ="d����'����,�]�ܮ'/�E[[��T�q��׷��%y}�R^�SK6�xpi�E��hm�'��b���O4���]c�"��ǀ���+�ގW�kY��`���?O�s�@fJV��������]��`�?��|��]�#8�NE'�Y�}��ky���8�7�9V���'��Fؑf5�Qv�v��	@a?��D�3N�O�� @Q���]9 ��� �-W�K���R<܆"���b��N��e��.cF@���%6Q�u�����3s�ztʷ����%(�3o�`Ҕy������Q%zyoq�+�k<��L�x��`l�֩!�`�Er[��Ռ��4��L�cm��LZ���êͯor�ђ5.>z;:�7^r@'�mK���	u���G��n3��H����t�.:	����]J\�~2��:��"ә���J�0X"h�������=x/}H�����h<D�S/Vz����sA����D%��m\�g��.����,��G�d�@�\�4�)�.z8�����!���wղ��:0Z���:�*^u��p�kWo
=Uõ�m�bǀ�Y?�E���(��>ҍzb`��Z@v-����̴�"1O]z|Hil��;Z���8�ׯ�2���=Ԍ��W����"�\�5�ar�{>{�)�C���S��H$�U��y�mU��r�b%��:�`��bB�+Hx�&֨^���[��&�q�]?P%��z%��ڪ��3��I�"Ðr����ؽS/�̫r/V39��'��4C����n ���m/��1w	����ȜA�Fa���2J ��@�71�����"��h
�!4;�Fw�?��X���	�	45VP��x�ɭM�T�=ʁ�2r1A�̄����q<U��J�Q�Ա�9T�S�OZ����E	��G�e�M��w&2Bv�֧�sd����-���O�w��A�n��SA�^~6`���� ����2G��czK��9���
�
�P2�5��0W��z����h��h-s	-�$��Ɛ�_�
�j���)�95J��R<��2*��hyb�B3p��빲�J�˭[Cx�l�1�J�����6뮓�T��3	��^�$"�.i౥�zط�d������Jp$U�Qx�۟� 0�H	�U6W�Ab>d��;��^��|t�~�{[:�~��9���+��	֌X���a΅2�L�0푋�tL,;V���V�A���PS� C��R�Dfx�A�po�Ҵm0�I��M}&-�|��-Vw�w׸�x�
B��������ꅤ����S/�%y���t9=R��2����H�%[su�/,7!mr��������
K�ZǛ&��KU��e�
�[��oqc�d�%�_����-�6e����-Y.V�G�1���H:�_�+�~�_�n����ӷ�a�1�k��3�~=�$�>��("��bɝ�<�:��fK�>�z��j��?uیL�y�ɏ����c?g�ޚ� ��t�h�z��ԟ(�I�x��K\h��0g�k�X���͒@M��mٯ�o�\�M+�Ԙ��'y����z��N�ƂfX@�ca�|��Є#�PXԍ�ػc�����s_�#�j{~ã��ۊa%5�M�Ȳ@E2A�׿��1~�ţ[�]c�g��up�҂�B-o֤�@�4�2�Y�rJhP��BL�� Ezm{t$�m�j�g��2SG�j��a?�q�o�Y��3�YR%<��n�o��ԒoO�<;(�؏s{y�������PE�?�]��74G����٥Qई<����w��ƃ �/13�OG�q����Us-�����[f����r�� 
�v�7��Z{%��-�n���8@X��D������|�1����LgVL'Aҁ���z�{���˳}���3�u��ϖ�!yѲИk���*}�M΋�N�J����i"�Wh�>�0>�V�Ex� ���$ʇ�0�'HG~A��喛Z0��;r̲/��L�t�Fl���NU-eC�|�b��p�X��~�R�r��5�OˑPjG TǹM�s�HK}%�B%	�Z�z�(�6��d�X��o�1mZ���k�c�*Iq=�֣��f
�e��np���9;�vqk�=q�?�H�d����_��z���5O!�(wQ��Y�3)����<TG��Ȁ�X�"_+oŌ�$NX��T<���4�7�Լ��[������e �%�+�n�����/��ٳr@��(����/�`�xdA���\U���3��4����Z�����b<-���-/��ͥNm�_��N��:	���-t�g����k�ASq�Sx�D��T����,�(����MuRN6[�\2,��4�a���0d�S��No7W3�b���X0G�X(En�bf��%��𒌖�ƣ�B�n��a��ї-�,���� j=&�X��/��Qg��(g>U8U�
�����Ǒ�nZ��;�	,��*YK�{[|�m��sw��h���\|�� 3�Q�B�;nQ��n�1�r���Y�ա��9q�1��J�u)0W���Ηs�.Y���P��f�Fj�&^|Xwa�(
��2��M��G�w����V���6�7{�8\���U��F�U�0���s�������rwbW]�q!G���#(���K��*˔f��������*"O�}/Ϥ�{4�1?�	"���K T�dH�z��
�m����t�P�DO�W�4d��A�����Y�v��z�/���$�E�<�I�6�+��T#����ȫ><�U�I��]��0�Z���Q�!����m�qZ�P��'�o@���vs~]]�-^L<bQ�n!�O��o��X�N��(�\�U������17����Z;2yOn%b���.[�1K������dF)����v�@5^����1����w	T��|����ȃ��YrrlJ��Ӻ$���q���~�
��qv�\�FTvױC�Nn�6�w��u�Jy�H�Є70�`/�2�@�9F5ez�>}uRx������T�mVO��T�V�\�y넭�*�ⷑmr	i�z/|S���ɏ4�j0��O� zQ��B��;�x��-Y��8v_��r��QJ�2`����fg�lpVKO��D)8Q�Њ������V�?ג#NJ��#���Ġ�v�u��i���ol�P[V�J4<�v��c5�=n3�S�ś�,��Iϻ/���23�&����g�W�{y8��̛pL�7hˮ�{�\y���M�:F�8.S�Zcu�^�8�>���{I��.�"'�	a?�+	�T0���u�Xֱ���Z!�Qi�A