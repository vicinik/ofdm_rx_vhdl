-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ac3uSy8KQj4XsoUBVg30MWa1uQTCQo+Of8GsPUo4IA/Lu7l2HR5E7o/MPOFg7I2Phpml2GwhYIDt
h0P2ap0AtHUFWCeIBz9n7xZm3OfzJhX2jt2d2JkgEtARgE4/POkuAqFPhxov6ZnFZOwoBLPwzBzk
G+hVNr7bhGZxGdDG6JTUWGXoJmvBg+iDOWsyq46lgHY9dw13NAy05rbScckGvjve5s8nRWJ/C5Wt
VfLaa2iYjcVg9CiaLT7ktVLJzXqDG3iUeemoECRR2QWWFgF2Le3ANLiELm/+FwSv+b5NTEFDTFOE
GrFWiULMlts+i89YoOjmwHcoSQAgCtexRxcK3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6656)
`protect data_block
FR3vHcpr4ag8VvEOhItsoFAKFjzKPlTIsbADfPVnKyx/Ejtk2DMDfc9xzdDTTPbMyrU5g9ROWHpg
rK8xVeMt2m7y+jNUAot77kKB5qa8zyibJbkCbSRJOmPtw3hongEXKcgV1O00CRmxpz+ZOzDEnnYz
T3pu4PqRByFUOTbSSePEfEpOBhhTA8tjWEH66j+hsR7az5MWKcfdpn8o3yjG0gwFbuvoTE6t9Jhm
aFJR7ABzc21MniCS6IOc0Knq3c5V5D351LFndoG9dkmkH/sZ5KhWE/ISrseBCotKUoZgo6lW5Qb6
IRTRnNlc/lLHrS+pioGXIyPFZ6aoXFwfjCYTnqqujWetxQDBrI9AHQFly57pDkGJ5q1EUop3VjZy
Er1f2h8GUoeS991NOwfV+L7yb66Ml38UDEPG7VQ0eoCYUPVHm/4nzuibxE7hjzS/gCGW0xq4dEut
3ne05oOx1Fx4xvr+LzEhF02x2DT7iClbWohMOo639hc4tETA9VNKo8AjSOTOIu6MzLRHWnPyyjTB
tEWGjsxHSITtnOP0QZLSKUCuSoRw12OfGgj7455DnRaFDD9DLb2XK1TCS5zsYcMZArqz5jVvumoF
Gg8HaWAofnTGpNtdmCyHYjNZFW56dj3ZOR9rddRQjpoTIIHwhdfoNyFKedcB40Mocv9+S7iVRTXn
89XuZBUQT/ELmBpDvsi1sOVaCQUUcmxpRoNty7vFEU3lTRwQywObC2aYilN4yBM/8FgHaJmX7HmA
0PINAWknEJfcLn0MEBFJFdeyBfJf22icSAUjA6nqlQWPwziCbugKJcMbyfCeI2l3VV8moiJyreKe
LP5hl7NX8t37l+gmum5X4c/QhJcYOwdCP3Z5BU2+KA353XymCw7UW78VUu06ZD9D1irVKB4qCtOv
lK+yJHO4Fn8t1Pl+IkICAr2/exFkwBswiSoPNDVapJ/b5UzvMmNdgf3/nfoHnyHQ729jYCHFY1Iz
DpDIxGPVw4YZxXlx0HfqQSS5I7dynjfOyoIix7u2QztEOwq80+V4IYG1OodQpRpe9ugrx9pblCG0
AfVpwFYRaxi8CgKE5WwJRYYl6/FgY5DUB3+2AiNe4PhQATxJqFf6joyklk2LbxGdfgXRyBXd+q9M
MXVvPB/6++ZsEJwT6R6uOloZHypMerkj3UoMGyLnc1hPV1vssSLlC3S9Fl7t6OrRjC5dupVIhmuL
OPcS++QUSUbiECWUSpFkNrO4WYhD0KJLTc049VyJ9sl7o09kqoZF4+Yz1LCGZ9fSfIUwD0myktLm
/t4Y4laF41tBO/RozWZ/RYs8r1y4IphzksgPOwRpgaO8QpymgZfXHyWpwweuHDOcP6SlAowXDVJD
DK5nw9vila3hmy8IDKPejpoBoLZ4Ua6ZO1nHQEPnSWVuTOs8NHxtQTwpeKfkiQvHEI52yKI3R49f
Bcu5fDEt32ENn2estpPVEfJF08yvJn6m8/1NZ9CtMorqsQlAXV9hED5YryRTsvQUPzy6q5g0KRvR
euVsXIFJUf56df1t4yWVH8zGwrWEnTcFqJeHe/EhsupYfgQMSqD0quwv41xHWjz1V9M62pmhu89C
bqxy1pB1UJeQOEr2xgUkiYpC71GGxLwpJhR2UtArCwI+3bKW1YXgzJMNrVsv6eWo9APkcrEYmg2u
eP/xruSabvoHYiO905trlYRwPHAQxYk5jcvgvOMM3fmhaT1EXJOwj29YmgNlsiofURPyMeW9BcWl
g1lutA9eJ3ahiGfFiEnY1fPaY63mw+XKElHt2pAUCSVzzuxbcX7kT4DHEAnQfLjIrDnEQ3+p533M
9YGHuRrFJJv6cKOMRHUwzunYRvDMbJkPbHF2ppNVjJGa0COZN1YzGjcBssyzOUNkg9/7vKXSTiEa
OL3/nFGeM3wL1wgJ/WdN4OCvrqADaDmdWYRsbUFSjQIH04PXMboU1Uj+SbCI5ySC8+15CxmuaeoB
CeREV4VZ8pQZoNxH8S5U5iekrKQ4thOnA0LEMG/Hg00Flfg8e9JTSDFTKpJcE1AWV2e+g8j/3kYH
jzgNG9DlBUx700CrM/dWM8ghvPaZDfN3XCtVQt9sk/ii6DmP5KUp91CpAvHij2edEHCiIQCFTTCt
2YYDfDlDqc0YtZ6OVh1oMUXhcFFJb8Oo8I1MDWtt2OVo2zHHHcbSnuQaXrcZjiN/q1fNuit9MDzw
B0Cul898RDUAy3oA7R5rlMvLx7qWsNkdasPlBRPscf8Va4Np3/6drAEgxwxN742ethmmUDT9rXhH
r/CntAn/RyU8a9+NK2U1OKeqkzcsWl0+1H5bRvk97mcOK4ATYvqOMzjBGqScCwnco18fs+ywvVrJ
LYoqVf4EN72fjOLglKCByZDQRBUpHcGs7r33Ez+TwarsQF+2CYUnqJRlgfPRxJiSuY4Q0ibVkTdC
S0+Gpc7opSzDKJxUSZb6k8sedBekUv/8YVextyRJp5im2rpe4T98ucqL9f0CVEXFyDj1+MxmngJg
/MVWaZuuKg3vAP78d0iITXNBIVVnoL2GkWuNbl8m4fqdP0C920n28P4w0llYxcvCeoA8uRVs4ftp
bN2shIz//PDXyr9B5REO1AplseGQIG+jVAcIL1j9JUZfdh4R+ONVUBOGFKBoggxpDgdvxJ14/kaG
yVhBOtQQV1+Sb/0N+BhbBzhykWBJuBq0AlW1Oup7oDq7iQX/EjegcWKxWIWBgjuVD/n4PKvvKzHF
ovlt28ikx6zIxHUu6kcn1qZAv5rjRg9iSW0iJ4wgJC+//4fpdG8IzrOCfmKDkja+dG2hwibqmp0M
yjQI65gT7K4k1Q+2RTum4pepEjQGxNlHmUCPeHwjaKxGRXwwlBsMBCzuWb7/q09c9zKpkQEw86Dq
D1r62FbbwVbaMy2CJvQD6Kzv0juARQtk0/8iO5mzs9Ms6paIWOoqHRENRfYE38tfiS/I4JBFcxbg
ki/vutglUw38A02fSWiIqhq/Qk3d9//D0dtEemmLGPBgass3ALUZmOx4iy32KDUYKiX6smg4ejNs
doYAmWoJ/915MtUk225aIllIcHLQvJMS7kWuQRKOXXQxZUpzaYCvoxlmoHc4SwvwYSbO6wb5Rgg3
vi7fl3j8vSRZJi/mgYcZKNyxoMV80WFMPF9TywxcjvjCMvbsGfHq31nvKxtIOY3IsGhOmdqsQpX0
m63CObCYD6HmG2IRe0/d0P+SrDjAfhRcp8ajqFZxMyWojZJgfvxJInCbuqok371aTXEscEQXw1og
wqrXbJIrQ+malpl+kJHsBkfnxKfXMK3XBqbBXaHfEFNkpK8WkcPwMBoNl8I0Ce1euhgriRde4YDB
pn+KzWAGa4eBlHEz0Ybs3xGIl9Yeo5sjJXryihWyZt8cIHpgtfUmsbNqcOv8Bho9j2VWPB/5M4TX
0mhGZY1MKIbUo879Qj+4aAe3Zl5hN58+hAqC0+J5saeXcn6BOMLXowdl3+aYItr9fsr3cIvaFaHg
mJwc0Ejs2ixxa+Kw33c7Bf4uya6mytNP/os6x9R3YpeYzy8UuvTxgvQ6W0RLweG3a5PH+e3MrRg7
1xJtnkm41mcnkfAKuTFMSRbEQ2JB4mNi4jVht6NDjHeMUAcvsd5mHLx2HLs6E7OvcYHgn4Gy3ZSl
DTChQX8oUHVP4LSG/6qY2dYBehvqjfPkInucOPBEodzLGX+ZVdOvfFIR5uQq+9jA67aJMu2Hw3Jy
8Pad1lqfVCvbM2RwJtuV1g1O6ujK/qSv55olBpkMy7sHSuhyHXeRWQF9PN0YYMDy3JsfBz6ar630
DRROUQ48OR3pR9KVEBfMb8Zoum1zaSK6sk2L6TA3J3l5BA9NTNpz+Ozd0owaEEH8+SCngKYHQKaw
Ww70Qwj0qeiXqSKGPTziqTELGU6LEAKOOCrgDTAuWnw6UBmKCebYS7EKnaDpTrS85MIiTZo8/tmo
6VsK7CTTeyGZK1i09rjEMwwsCIAnBksHNjpl3YINx0h21fmml35mIBxPUzMvwsDRMt6O1RnoYMtr
XNQT3UIA46whguDb16ODOC44IaA+OXW0QUqCvzA+o4T6wTJNQRlh5T5MxHJnbCa4XZXwiEHP75Ur
JAkrJLDqhZdApyozAgzepqOx/kbvX9PMrpCe3oUWTQEKcgJHYR+aXUAWEOoeBp1f7W+mkRgT/0uw
TKx5nxWCPbGZ++1qm4skIjMjS4DiR7K4q5z0f35dxMetSlG6mVSx78t5pDO/Ni5pMOmf3EgPOOPZ
gS81whoF0MP4wr7gEsPLb4wmJDm+OE33jtQH3OFx31e2SAnDBrVO7zgopsDWzJAYXuSDSimBvT8X
bkMc1W2rkWyUHD2YFYnMn/3gukwidpkdOLBIs6h7tRiliiG50KlVW+sZN2G1t7/mMFvQ4qBDt22w
mAMJ65yIsPcwLfinIg7JlsL9jw5cjFoVAIAN/j2bfkWZTBriIpfuu1QpSlDnNFHV2bSe5B4cjyn9
vLRYcphchvFA2Mo/m/atN8aL320AVf8F/bkUvNcHtiMnpiefznWpeDUmnO6vMX1kFq7NY0jaV+1O
eyvSrq92FXg42Hifpdd4E1PiK5E/9amxEmkXImFVuyzRCT24D/vqFtRJ9lsFyEtEQaQ5ZuYdr4me
Hzc43C9f1AdYWcQ9raPus6myfKOGHLS/Qam+mLWAfEKk9p+9Dr1TWDqUwkWPrnAzSgj3QGf4huoh
wAnAHmcXNHpHPyqbcd7KrrePqcWrgl8NpWlMp75aziAgne85hufznYwExZO/mWKWeY4qgfoWteQ+
zO3WZlDl4/pXAZznECSK5KZ444v+5Cqby+u20J/8pW3xTnUPphjK5XzXvMIzHzQRlMtIuUPznhZ4
696J3e16esVyI7ahL3n4GlogCE+DnJKC42Ktngq4ITli55SCydsvCCOqA7laDrY2nfSZyXUVKWzs
8U9Pvlggaszb4G3795szA+cP9o1j8P6QJZqbbpSvQVc0YTdHwjvtI/+rr7n17YCejEB6T4WsQX6T
PKDPTeHoQWMt0kyhIL3gUx14XixYOeLv6o/MfSgAl6z0gXa+H1B9PvalaCdKGeTc3yudPesJDc/1
KA05FF0AKMOlZ1t76N5PB9zcpB7Q/WRCuKc04Qbwg4RB8Iey6neCdAwYLhNDgroEWAnhAZU4cKkC
Fzhbz1eKNq+gRLxmRm+FeS7t44xnpkI8F9hMUv7TxHIsOT56jHV4UFFbaajSh1eDTc6uaWYZDK7e
m5JTWT5oOsfhDyY22dmSO5W0Pe/p3wGVFYXyQyN3VIDiu+ci7qoAy2kIeHSZ5/0HIwloM8TpaR7M
XsGQ7dY1ZmSp1F+r9GDN7/4E8UKPiJRq5PzO57wyEy6r/Q7tj+qt6w/xUhMkV+4JAUSnLL8+FlLX
sjVLoxitJw8rfmg41/IYhHip5WmJQakBgKWAmzAeP6URciJ0tl71QdmZfkQCu3ckz3t67kYtrAZR
eRcJfKfIdnj/sIby18xKpNZB+zIIcgKMAkSWa29uIZqBcpDSIVszU2AHjtsvs/Hrw0TDaxD5FF+h
3LZNPk5XjWJ2YnI618h0OYgHTFU+qujLUTfpAtzyGeypvP04PN6OEDig5l41D65AmBMi0KZZZp05
xcupxkYedKFYj5cRjYV0nNLjZ3atTn2wFYq1uvc5qiuGJBKesrvpKsj2Me/RwZFsWG39OJ5m9zv2
c8zUzetmXQR/pEARTyd6R3M2yqubmdRbtfX96eup3ZlOSf6VdQAGQPxViLQ1fexWgJJsvwD9IgPO
pxxwpby633yyHRUXEEiEHe0X4Xh/C+YksCd49fU/OZRZZEUhyXRowqkXlGrVodIQwzJ4PpVb7oTH
VWgsoj7Am+pD+rbeOcn93rtYHRxj8jJV1ecMwiapmo20H8hb8HsvFvvk1MHM+aqHvmuMJbYzrscm
+k9YqpePhzfCtIE7jxgfGzKWjOyaLZLOUCOvh1NuH4gWiF0nEHB63r6/AlHAQyOE2/hnAfvnYG6l
1rBYDMnnMRSG1BfeG6UUqWkWadv31gZM2k9ueMGBi54z1QgFG3LO6wf/9BmXWL77njx6YjafKRmT
MisRW731EZCEYwOyslD7E7LEjoYSdCxz8K3zEWBwWRdRvC/fYfXI8QoJskuU7Z/M8BR5PieTV3RQ
DyqXmU+MEHS7MaXJzfkbN2kUBM6vkM3q1oL7Mg80t2urgvC4sWFDfzwzPgaXVJUPEXBIaibAmWnE
cBcqBC7fZBeEY7RF3a/jyAB7RaJgdkEGSKZZ2G9801/GvZXNR66mAMTBNzLlPOw67zo3w7i8aPWv
z/Nl+xBTc6mG0iY39S/rm9TWd2VmSZ9geCZJgZOEMqH5xirrAnSwvvtkf7KxSdSlvIFiuc2atAjl
jgySuhtWQp7xw6IJVpzLZV8pQq2SFi6T9Xdn58yuyovUooUZgXuu2vGGI4j1q9VT+Jthc7cr0R+O
/GRT3TjQca2nTW1qUYR7VIuMi2MaKPoykweAdrCOQVhBrbcoNgDov3Gt88QJOz+WiuDgVZScm9+4
oXpNeWMzK0fJp0462BvEeBahEyja43dteD2kObgut3quJKyr87bPKAC9604v6faIuEq73MEe7i9H
8RZpy+VjORM5xN8M0k4mXuJI1Y91ryg+bwE8GR56nYonZMCZJ2HvNJNQJWQY4aNnbQukF8YZUJIO
ZY0fq2uScO13KETV4wSvYvkwBEj1b1lCtZfDwWStf83yF6JOeZ+DQRJIp++Jj745Iiri6PmEof0B
NXtZxeMfTdiHOfBQhpfsYqbizXOSLF2Y4yWtagZAJDqUbMq+tGvQZIyVWqyrrT/hxfTt1jhLJ6KC
iwkqGlctjQTj0D5V2PdX561CQwaHVrFWZAb0jdv0h9wcFDHnpDXSub9Fk82+eksg8Rzsjk4/Xnvz
k+4eP2WmQVdUlW0H49WOIBXviJfi4I83yn0Chmwa8wYkGFlpx0RFKLQqnMCFt15wWgqdqJsXb8u4
bWNkgRQgf4pdN8d8st9EWGI8GSBG9S5UF1eAqopd0ZaHi/FL6sbKocKj/USE1CIrBwsUFK97BNoD
pHmvqtBcZ9d2fVF2dNqNbuPKFbKET3Bw2HPPBa5KFXMOyU6mO8tUsc8OjPs7nt7oppqxvVNAgkPo
P2fOoPKOUmFsSqgcBjBFRgksTM37dquRX1QTfkx+Up75lTKx63NZzLwjahE5gIIJJWd0qKKNrzjY
bWYuEafoa/iyqL2qjdQFPYa5Dfrpkhp+nn/bJm68sENZ/ENQkLXvc/d8+slAN95EpqL+6fWmEzbe
INoRrRQroGbRt6mJbp55s419x4at8gZuz4uZkSsGmb/5/IpkJBXlgBvHKae2HX+/opN3NOs4G5L/
6XeBfqo7mdv/fMG9LI2C/nZaIQo44UAH496cdXc8fdFvjk2mGnXZmIEOW6CioyuP6lWoLRDguSii
uW4JQa+iaDZwTKy745ow+3v/OvEy6bhy8n3sV214Vf5st7sjw8gpSyDXvjMrpTjW2xCqRuey3azY
EYXQS7pxGnFqFY3FPAksyxEOUvLgIQ13w3DdU0mwncAwRJuugdHG/DstMVS8qNtPjTJ5OzcFAIN2
V/CvPf6wznq6jETTp4BYP4wfti4L4fj9+KxMSr5Qyhgo+AXnn2jdHiAK2W7a8PMVizzl+SOvBfbT
ig16yxuwJKu7fDFmGUYsIqGHHXjjZ37wle9MXDNQf7WIKgGupc2dp8neJyIc1HHDd8ADi9CtpYF9
9TOwUVsKk1ksh25hYa5uDF471megl8jkxFIump9P/tEkqLAMnja10/MH4g1MXz8GEjjPhxosDoxS
akdlLReWNA7MjhH6thaP2Vb1xWhGDxzQB4AZRvJkAAqO4EmCYouGI7fAXm5C795BqN1vBv8JfxZb
52ATqsr9kmsJ166z1FUqe7yF/KPKmcMD7uMgoELPjQeIeOQjlhP2i5LytmwQ1iW99yQFeGRrIFoz
HsGloLhAkCSlyOX5oI6UcHK9nT91ZAiMLfCA8TGNo/Jw6WFnGe5MQs6jrEoLa1SCfkOndI7B3f/R
c37ugZ34TX/R/owFz7/YNQA75NYgfvXzhMDwWBIthHBDebECmBBjBX9CL+94acDph1WuKiPzlU7S
w3JLdGAi+AQC7EHLUv+eiDPAKL6A1dGnwVrFVwKspB9wJfzS4IU4pGAiBWldmT2tg7UUzYMYWDU2
/eM0gu53oXgKyJNi4TJ8s81TPalsKOqROYZ76Mx67dOJabVwDzPCRvRWLRux8tE4Jscy000vqZJB
YNnTDN3mctuAuFmzpaMuVpJMYgn95uEV/eAKWs9wf6Wxh824YkhRL1Com6tbRHmZH63ctwosc5zP
iX7rNMLflNPUb66hOzxNVeuSVLBK70P6I8T/vq7q/Jxo3S1vcH4ffe6u/VKH5efkN4WMHUE6eYu9
bp9aJWjZZUVVouzKR+oRVYCuyTdcBQqwOwgvN0M8Rv6BD4Qr/L8WXgDTXHh1OBZElPI5mKfaV+ik
cnB2BuyuGUpb9YZ8mT9k+bpqJCIynSsqJBsgE5jtLliYc5rOKJBo3YTcT9b/bGH4Q9JAuVUJH/9a
OKeLh6CoTQQ7NAZYghwqZLmcD+D3t93u5riw3LVgDOoP5y0l/Bl+9poeYxPdv06r6hzkANE0Zf2A
GL+2Nb5gO0kWVZhgjzJU7cDdnnhoZ4Fticlh28qC6wyb3KiB0tg0nb+LQr7S/R0JxtdiS0BsacWo
V/p5ITANe7e3iYgd0bCSx/fAAUdm4e3RFeY36kvsuHhSnLhyOJioHCDF40mgSTB/Lg4tybWy1S8k
bf08gIZaPoGOa90/SGrtGSx8PJzMhtKuX3RhqbKzof7A3Oieq3teNmPPM34=
`protect end_protected
