��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��Ȭ�SWC
�^�a#�yu�b�+˒���62^���f1?Z�b��tUԑc�~��ĻyC-���<M��B�rN����M~�VG�����u�������+���Iъ[uIJi���E�8��s�m��x��Um�7$�q�� Үtj|·��:B#{|1�֠TE������,�δ`�5z��L��T:r���2O>UQ`�Ng|E�Y�(v�U��O��|(_%&o���Ⴈ��<ĩ�|�F��N�T��*ib�=��,nZ96tt��pt���8N"p?p^�/)v�@�wgH��O��{W��h7�vF�ʾPT9����?V���U@� ohx�z)��2���{��kE���ŜP�B�^L�y0��3=���ɱvbzXv��6�T�hD��u�K,ZTcj�,��!Pa���ATQ����a��!�FBn��[E���)�,��"�z���	��@_?6�g�6��A�nj���b6-
���:�Q)��J؈t�YU\�������?K�F��W#�8+���uP�[x�+� ��7b��p���
�Y?tp���H���{�S})��e��f�,�21��V�B��)Xj�c>q�U谨�XȱQ���Գ�7Z��0Rg���
�GD��tr��S���x�D��j�\�;����(9��X��|���"�k��{������M�.��{V�=9)E��T%+���>v��A53d�ĳS���f�Re�'���p�e���K�����Y`���sZ�nw]��x�U�L��P,����ݧ��:
���iL�
;6������qR�N�\��) G'\=���5��n#�y���J���t*�[�1g��U�#i�}�vO������ =�8�'W�����m%���a�W�5����ֹ<[ӧ}B/1��s�tM?+D,R@�^_�����k<��l����	��n.TB*l9ta��Ƀ�����a&2�v�Բ2	���?	�XΎ[K�@�����ʡ����uy36�{0B�w�݂|KN|�6�{��^�P@.8��d�G(m+����dFP��V���b�O+�3(��;��ч͂��G�]:�&.����"��������7?�-����ueݝe��o�:0CZ�5��l��I'�Y��&�w\�NTb��E���b�R���RM�E���>�>.��x��/�.���2��Ș]yx)��������4��*S>��W*5§'��J�T���]�C*�6���� g<:���1�e��}����}�r��%�SZ`�wGx&Ǭ\��$���x� �P����^gт��0�'�v�>�	���WE{�n��9rש�:S6nS�����T��M����i�c7%Cti�v����rk�4�V�;́�g���4L%�mD_��&+i�	E�ғ@+�G�5%=����̀��Y����p~�(S^���y��D�ZY��ĉ�0] u�2�N|v��ْ�5M�x�3�d��3�_�c�wJ��B(n�yq�-���X���E`)-��Ӳc�:ڨ���$���2�3��м�'b��+���}T�I�0�il���(>J����eUe��M��Z�kU½�������y��=���HY(�ɻ��d�d �w8��~:l��B�m]�ݺ�|�N���{����G������+���&Fb3�"IqE�z�L9�K�吗{C�W�OI��|�8�y�n����D�6�J�!ʂ�$��Y��~�ʭ= f�}��6 ���O�K���)OW~2�`������YϑĊ�U�gFH��)��H����Ɨs��vU*ؽha;��yw�~�� A�`��?5�"J���{-��SimA�!������ҽݾ��g��2�>o9�"!�APKP���
8���_P�l�)���(W�n �^i�%�E�m'"���~I�x$�_Y������Ma�NK���/�5Mf(`׶��Cė퐃>�xH(�����|r�D�X����84?Y��˸���>�H~9�^�l�������$��;� �����}��b`���[ �.���W��� ��QI����}�*�%L(�G�	n�/B@I�U�ٻ�Մ�r� �~/��i�p�Q(�~�<����K@��Sr70yn�`#�\�~y�����ᕿ�%寬�M1�y�@��+�]��%�h�'�jP0,��q���_�L�T�2���Jl
����1N�+P�L���І�uܵXn��&��	��_h�ߒkE~Yc5��i�3<�����b�u}x3�B�����բ}�Mm�QngxU 용�U[c���s���uδ��4L�2\�,���Z���[+���3��OP�߅N��S�c�D���D����.�vb=���MqHZ�����������n��»{�ېk�R6KJ��~�Xظùi� S���ͅ���;���J�r/q�
!VU����vh��Y�.���r4�2��N��M� )��;��ۆ��E�I�e*W4bܦV�2n	+�i����B�P�iU�[��f�(:�5�6��������i�S鰳���B�A�G�Aj�KB���G�!zVh�$�cnU�Ve#��֞(-�&(����8~K����������7H6�ӶV?���	�2�F)ŧ@V>}�i~*_T���)d�Ksɯ֧eM����o��}�2}R?�_�>����|bE݋n�i$i�h�dҰ���߂��0��}Q��Q��z�Q�7��L��iP(w�qtq>��͈�],� {�5�2�jj-ܙ ��;߼N�[�ӵQy#��Uے�ﷇ'J�c�j�=jh�EJ=Tt�%;�U������a(.��J�����0k��mp&k�?���_�Jܒtɟ������٦��4�n�����@;:�i��*BcZ�ۙ��j$����9ͨ\RI�hor�hI�FID�1�$/����4r5'uA�.���h�l�_5%hQ�Q�^����ҧ�4��͞�k�l����:w%�'ߨ�ܸ2�;��⁑1�-t��Yۗ��BDr�y1�J�f0<���8����7�è(��W)��
�`5}B�֪�Tx�
��-���=�L|=�%����>�{�&�U����%;��BPEe��g��ü���D���H",��������PG:�Ѯ����E�*�kʷN�j>L�}�uc���IW���p�x��?zՅ>����4�9~F�1#�҄g�� U���F´�O�v�C~jσm��8�]��x����C�Ckn8��`u$��C#.�,
po�݅��.
ŚKbh�w�Nb��u\ E���wސ=s-}��qE�P7�Bs��Q��h��l� f��Aj���w������8�������t͛������m硚lZA�ꠢDD"�,b�%��/��4�K.�?l�f~�T���!am.Ɠ^ri5�h�\r!b��8���{��OV�~!Uk��%�$�bm��e��W����2W[<�^�p��MV�W����c�T�6��)�y����2P4A�~i�:\DI�/�K��UDPWp�W�釠Y*�@Њ����>��x�2���BR������f㦢?�(�d6��_�y�тx�D�|E/<>_mWA�����O����4sέ ķ��+(����{EZ��t�t����cܪ��Cz|,�����.\���1в�Y�훊w�-)r\8m���h8�֏&�f��N��k�zt�}uԍ��ׯ�H"&��C�9@?�k���_���Z}|�[�dy;d1�Q�E�՞��K�6����p���K� �7	0wГ�ç��i�n�}��%)4�"6Y��_�fN���W��mHZv�a�H����A�Չ�ݞ��#�I�)C�HzR9>�5kv�yj��h���zZcL�:��"�����=,��hx��b��#
4o�j��!&�l�MȻ|�T֒s��;�$�=~a���~��?#@%��e��\�ĞGt����[w/}X-��i�sMYu�A�/��KB�꺴���l��v�6��|>�e**���}zsD!���f�:㞋V���+��NHCy�D���D.J������Z��� �e�E�9,���D��:�Q����R���]����\q$�J��C^�3MNٛ'~��Ky�_Ǧ�P�����҆>8b��sڍ�J!��M�Z�?tQ�]0_���ۻh���$���Θ���Z��~Kshx�`�j����*�%,,�������&ˇ]n�z�՛��Q(��B��1��1}��ۻj �+�t+Ƕ���,C^��X.i>�����}Zㄯ�F���w���u��� ��Q����e�_��vG�/��&����;8W	#W���
'�"}�������3g�:�5��8n�.�+�7�r�y����P+̞k����O��!�%����r�^���#n��8Zy��l.۽��UsC���Ӊ��2R��t5���'W0X�R�K��m<����6xЦ���h~��+"�9��:̮�cⰢ�n�68`0f���x>@�eb�{��7��tar�p�Ej}ww04D@�w��� ��E�*�$,�� �B҅��jM�*D���g����S�G�K�����#_�� Yπ/X捧��8n���!�Ȭ����uPN�`��@|���j��_a�ק��F���6s�ޱ\�P �R�n��>��8�+�ͦ�ߋ��o��4��ꝟ�n�+K�4�����D��8�:R�hʚwds��vL����`���&���2l8����=�	�'��`	nMIwZj'��5w�N<�ښ.bA�j��<D�jXAж�Ai��"i9'�;}"e�2CBLmE@�8��K^��*.Mh�e$�^�>�%��[T�i�u鵥��~k�a悙VG�����N�e��|�0iLL_&�� O��[�q�oS�T��W�~��']I�y����ge���*����ڦ;�N�"M�(�y�`|I՞m�\�hF2�!"����Q#��XY���4�5�?֌TI|�r�5�F�mk'�ԸAxю!D6Et�j�+���u�E����fX����0(.<�S�)a6ܻQ���b�|i?a�0--��4)$$���zc���^8�M�;{��6WBe_�lhM������Mcν�ѷ�ϋe��t&=2qlHe��M҄'	��w#jy!�~��T@�I�e�ü��Z�C�?OHjZ`\��@��$AF��<`7�%QU6����V���[�N�Y@��?~�h���[�b�	��L���kI��3��O���<����N�g�Uu
>T��>>��͛����tk���D����[��c;^�Z��Q����#G�����.N�SE�l6�՞s���|��*��]��4ki���������������7���� ��6� ���FP�����2b��`��oj��\��8�)�l���쏺���V��gf��E�O�o���׍A�E窀�����y�]�G���5��ɨ_�����y�����pͫh�ʻPt/�wԨ%��Q��r�\�^p��o�b���X�3�=� �v���VkԌ3�+i*9��L�x]���h���N�����U��WG� �7�պ�7W��ͅm�į2���� =`��BA=t��w�Lc�̻�mRp.��*=�����2�� ��O�,�psP�RI6	�N�Q
�V<�}(�=��`�����g�7	2r����d��S��v������9�n�?����	Ss�]�_�*CZ�~����i�]4�\�'�������\��𿩠v��ً��ՐBAɛ|��T����6��@�E�d;]�1t��gpHr��S��t)x��w�޷�аH�ۅ�9Zv檮�wp��iO�Zg�a
�
��8{��.3��v��Ořl����-R��TB���3P_z6VS����R�ude�}'����S7�Q��y�s0��(�On��7�w��u��aNU��������z���O���qeLĬ6�~Ս�,t,�a�l��hzY�C���Y>׏�#T�&���@�^%��d��e�.�c��$�8��g����S��c-y���J�/~6��+U]E��>��E�̑������ɕ� �xO<�nx�����B���������cw�г��2-�pC���Vh�X��&�)ey�zE~_!:_�Pp�
I��oY �gXa ���ۯ���{3z{Ms�c���EN'*���|5|,8n8	z�QAi���rNpy�R�u3�s������Q���)�;�9Lz.f��?�:VJ��Zl��*u?��{s�k�#K�G��.;������+�<X���`�A�@�u�0�a�1T��&C�gkB��Н�� D���� dZ�NG�=��d�4�c&���ZA*5��6����"Q�(�8͎Y�c��aR�vx�y��4�=�t��{5ī�n��کm 䟍��ڑ��ܸ�'���cX��
��:KqA|ޥA*�5�E��U/�(�О�Zļ���K�8�� I��@�g��Ny+0����kl��X���N,&$/l78��ǌG�%"R�?1DyvB2�M��A��/�Sy�Du�p��dh�@�5�Cx"���N�_SU:���9D�0J�r�슃�=Zq�.���M��1�Ar�X���iPV؉e�
�w��l�*�w�F�)LJ����a����"s,�@"� ���:t(�)ZUc�N��N�n��YD��i>D�$όk�2O����S��yK���Y=CP�Et�H�ᴎ�[���)Y,{�q�������	wv�:$ǹ8�P[��8��L;��|/y�أ�m���.�7�� 0��:¼�Z�t�*��8��wi�V��Z@|f�I�d�n��B�b�f|H�kςh(�Mk'�VH��,Gf`�(����U�d�\6��:��cS��nE~S�7Ί��"rܯ`��5'�I��ZI{E��T�(�O��������t�-g����=Gq[>*s��m\�S{�Zl]�c}�wZ��rʊ�O��q�A�1E\M�@�&$�o��<P&�Ur'�v(��U�`c���A��S}$���vǈ�s=��c�R�d����Er����`��_w+S��Ɋ4�ź��Z༳|3[�[�e@�0���J�]����G�����S`�6y���!Rv�1����E��01UK�.���L [ӱ���?�zݼ5���K�މ�����sٜK��0�R�l�]{�
|�^O�sKh��Dbں1$�S�mJo��#
��(�la�i,��>��C����#~.�'�Ќ���UX�^?���F�N���l���)��6~_)��I5v��W�=
��m��$�rs���ԋ@�[�Re�"	�`.�c['��4LpĮ=���K��-��À�r��$���C�D&Rr�t�JV�"��M���MP#��f�/�$��u*5���.�������f��~��u��|a[�^FTj��u�?�j���2��B=����c�d���]6D�y�8����!�"�\#6����Zв� v#IMff��h����<I���=*�g��/�����.�l�F��/�o�k��<��w�V&I'�б=��YHv����x�1���[;�Fۣn>ZТ���/-	[-ݸIq�KQ��q�x����4W�!.���#��<��˹[>�z�f�O+�f����#C�1����N��ۯ����s����l�-.��}M���k�/</�>��i�6�r��
F��ъ�V�O�;��*�����RL�8D���'I�$a�q[LE�L�"q���a���;7L	zW2��\໚���^x<q��YD#^<�q�L
⶞��k
�@S�����ے��o�@�_E�n��V1E�95����6����OT+Um�|�Tdݘ�?�|^p�?�3�ي����c%w��p�X~�������°9%���e�����9���BYT潋�J�8��5�d㓓�n�1>�\D!U����%��kU��H
�}�sA���H�g�b�+�l���[C��ry	���7��-{��$�mv���Ǻ�����1
�ja�
�0���aCkw�<�����H{�x���i~��]�ۉu��6k�ux�ֱ1�t�`���x���U7�J�ʯ�ĵeˎg��u�������+����l�3��䦼���T\0��l�7���L��������O��֌Ώ

�[��֞>(y��m&������>
��H����C(�2�q��W+���u��b�슟=�������3#@��8����3��a���E������R��6:�t���e�|M�&R����X̄]Yʶ��q}A�"�)�s��}�� �}�N�ϳ^�zrb�3��-�*���lE����	����� ��)^�u�(��O�1���1��V��N����f��
��ۈWfO@��`M�A����M�ڨ�E�n	��P��,,��#��5-dȜ?��~�I �hp�=c8<M����v^��X�^������tQ�s
�;T�w�T�:�͊����!�5{���l�*���e���"%�D6�7��}���8�}��gc�