-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ABhl5hr5a3DHLZcOsKav2Y/NP+SKQltUpwD1n++p6MkPG9bAES8Zc2aalCzZU+ntPaLvEyldl7qe
ptOR3ow8H2DYiKvBrVFnrO4/pR9imh9XVozZ6XIQ7SJrwRxqdupMRstfmS/rKv/Ef3nmn4Qj+d3Y
1/y/AqmwuWlH4/4Iev+UQ+jY21Qw3BzdztNsrZM0LN1FROkJNGVRPEUPZf6U3ehMBrHGQc5QTgsY
lyaEcAv8Ujn7HT+PkZEu/x4qkRxB0OTdX90/OA/d7Nhndp4zNw9Vdfs+h1J/j4fgpXnemwCTfnps
81t/oaNPOIFyn+gjOVty6ziTQP3xkiPKdy70Jg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35184)
`protect data_block
QOGeF9wxC7zZdf44yly1WSSCocbRLXdAqcz79BTaS9V44JTh1ZSFZc3e/zBjr5MrEf/ie0rc4JUg
1NXsdvMX4Xe4rxYLsnUod9Hb66LkdbD6PezZiNbA1rUm2MbqdbFYS4ldyFHoLqFZRwJQer435nC1
t3XZbboLqTg8TLW4pT9HQt78flxlwGPPq+OHsJmFUrEM6eGAfw8Fy0zSAZAO5gQe7FhZzLW4evAS
D6sII4to0l2YOxCI66pOOfw6MgGX/KSfoOUSJY62cvqDmQwQpHfqrjig2co8+lNciYht2VsQ+Vfj
yb3hwz2lqoCBNSJ8E4Jg+ZmN55TIXlE71KJ+W9kFIXnWVq5Be+Y32hNfbdKqE2vf9ZFfCbAim+fP
YIUBYx+jKOFrpnmfi9RBeSR1sX+C5IrXFfI5pkD6Uz5jYXHaQ2lQOlEdvfjGORXfwlFhVcy+G0Kb
ZVojHJ04FQNLNYNebzzNLNlpiYHFv9a4vMMleZ7Wzua+lad0a8do+ZvcVfaJMU73vBokGO59iVng
Rzz0gzKuibrRDUBVRZw/3TJnqTMTbmOfyv3BAIH5NGY94XgD1z+6uZ0x2WBY0usyVrco6k7Cvlzj
rX4n5fG/l/iSA7cjJmcbRPk1V4kU+9MyF4fCleRcWPlEY8pxnyQxgjFWgBYIOQ+wwxbhjbHkZgDO
ghUW0MO+BIRqEZJ3U9PMcV+UIAMc4HoFN/Ct9pTkIOn5rQitUPQBge+SwSLcW02O04vcwh/E/iuo
/B1vxkeJhnXjoJkyszjlRQyteJISSj7u6QNRWDw/chTiuiwSjTv51EmyYT65Be3kAPNHlsEBEDoi
b85y3gV0zD77SikNwIp4MSDZsDS5qQq8cApMiq4SQT7j+uHjYLA/gfrXsiOBrkQDwndQjrL8kvaY
Vpmxx3VriK6WlXLW0JGXGepR3WZD22G3pPuk+rAfhB8BUhTDx+cMAwi7nPazAfs/R7E1LmFDsoIq
fGBUakwLgFm89WfcW2ou3syFmjmgwFD2ocEgbHUzeD6KEoQZ39TOL6719s1CPAns/7PgENIKcpqW
qRdQqge2LKUv7FCe3oJPAI6MArIC+mTASzixUiJwfhKctoeXJlh2NncyBE6nYAwWeQwUXHDQOTAQ
IKhtaH9A5TkzMzKfhjW7c5cXxZbbXX7ZXA489BpVFNwN8D7ieQ/NLvT1PhcurqoSs0kMsarPXPkN
NkRnZMQTUizqDBeq/RV4eH8V4SF3/bFi5udOweyOIaTyiNBmsY/3CdFU3RZ0cmI8jROcFiWMYmLW
TGZxui2XHSHT/ywtQ7D+6D2EW84dqmRzJJMvGTbSm+Wry77xG2dGxXv9LibZFQhWBNMDwQu3P43Q
RrpD0JgKeKlBXbpjEZhyeJagTraP5NSi8p5i8bq8eX3K4NkoQ32njwLqHiV01JXrHwsfcBu+qoLo
HoxOVrffXaj8yk+DK87KNJGDaFzeAnzgycVy8E+vcLvrq5Rv0D+MHprv2TG2Aphjxfp+QsVRqMIk
b0RQd5sPlYxz2xRBHTqN1c0CpUzwBmwIWhYoC1EXeb1Zif0xvFQpMOxgaUdySe3gPazwgxncX+Ke
RVp3+v8NRfOxDjlvOm7hX0Ck2Psc9eshYHnDN415zUbYJMB98mj+g2tF18ynBcsbPVkEDMl+/3hZ
UkUKx4gw3gxiA4f9l2tkDJi9/0TonD4dxFZMRrFcwT8RintliHAhCMgdHRbwl7D18Y0RF0zsu3e+
xEvBECjSjo+OKraAyNhrLXSAyoKq/nzBA66pIqmWZZCOsZx1/uogHc4NW4QMVaq0No+0aCYJvU4R
AtLFzljpjnDz2iv9Bkww0ZhjzQRLDM1f7mDoWgi1L+CeOYPWWpiHj5IEyF8e0gxHm2Wd10P1JPD9
hTQD991IQNCB9KqXXK4HvTD95WOEhYpZa2q8G2mdvst9MRzoUSkhbsKXdx6Rk+nzEQj8hjSQUthT
7mlM8YzwJzzsdOPmQt4Y6jIxHtBKV0tBWvA4i0ie15+J81kNboDBlG+eu4mIuY5rEk8ogz1AsdNO
sgsx3u3bKidm2M5SP1lptorCjBNjrUlrqirSGDnt+XUg4TrUJO28yhC5kGxzPXMXLc341oJRrZLA
q/hjgUbhsVqqPPn9rv4+pE/XIsliydagIJKcNxHYv1ex6jq8pq5PpJbBbznjWV5iCYsHD2O9sL/f
mEwc0PsQ8TpAL7JoKqD3sAGiA/S0yizZYetbZaSadexnt6ZHrU7kWMH+WDg53Pdozmx4WSoYLO7C
XhYnSwe1/rRUFo04Qj8achb0nE9tv2wvtK2yVABbGKaFzCw5X2QFO/XHEq0Wo3h4SrmmqGvmg016
9/MQN6UMx2UEFenSkrNXRDmIuAiWWXEeEx1+5BZr2ga5avkkLp67eBGGp5BXYxjriwdlip6yN6LB
Zbgt2E//OUl86d1qmzogGA7hUOngzooTzCYXYanjPq/ilXnkc62k0sHMwkZDtRdCEWAw9b1U8f2t
8qcfIF8lwjNZ3U1DQ0Gtzsaj0y5rGCCzVgsJa9fGSjYPHczc+a/PhD0pZFq+Wke8VXxpg4wfb4KV
RgybXDl2z+NhCIPZ2BIRHD3Oh2zDMMRcCcEoOUpjvnTYJAGrmfX5OuzF62UnA2zNbk7C3vQsPm++
uCDhmi1hy3ysVf5sjZMkPuOOKEpxJG8lxwn4jtPQ0KvAEokbsVbF1pAcREXKOk5cZjBtNEXQAZVZ
0rMyBDXmLVuO4g8Q6mDZQI8DwN7x7g2e8ohozcS8qiMq518fRlJbUJq+4GOp7g+iBshFxXgRA5qF
pqAivUsfoQlZm0sZoV7qMLnff4AuworTxKLe02gaUuGjjPzHJwEelY0jikVH/ensCeK3LSV2u/Um
T4OtRKiYZIrV5U6z9/GEWYrYzDnpBlc2vb5A1wcwUz2LFA5whNOeUyQb5WUHzRtznXXw6LBftIlr
otdUy4LkSwf5OZ6QKkYFIpg+8LlmTy2mnT4+6xCqRjKNBfl/UOWQITIAXPl6zW+mh+t+lxOJRvjy
wd6YUREjuLhzNj/KuATEY9F6tBBjPF+5Xl+2iRmQTlBMVH1cto3eJ1Tpr18gn3i3TUS0EMj1wfe+
ScEk0R+THZPEaXL2rzxDaeL8yG7sXQagTNkdOb4jTGK15YEhBhT4+kRbxhvb/x9BzaT7ru26Upe5
pZw1Sj+/Tp8tvdmXSGARB61b3yloE6eUuhBEH50N6ypseMjjFFlWZqFUQNiJXHZWpEK1yhDVz5GR
rWYyIh+SxBATTdNZouyZuPK147sK8fvvf+udrUsnx45pjJAwANx/nW0UsKfChGn37QoeNgG0zAPl
BBxV7nvl47m1xI32U9f0BO/DPMwP86iaLhIQEK+kaYUyx38CdEAJa0NfIQBYJFIE1xlVOF7E3h3I
6gRToGOUlVNrTc4PJjFjYATDtGJMxGEo9zQM6xOO5+3PcLxTWuSFj7/KDqlSO+ojqPhRK/Rgmcar
vQcJwh6+fyIiw3nvdzeCxH7+0UliGs1fPacenbRpEudTkGCzNkxehPyZWFNS0Sj0hJvNgxvGYL31
+KpnK1HGSdHlnxyp4bFkCh3VnhrfyEZNaHQOkgDIVlG0yHIGRh4IOC/apYuEiZ+5EETjsQ3UpN+b
Q2p8HLhcXmT6GC7kQfDLOguG7Vu8yVvQLqiy4SsH7c3VqaeUs/DuV3yuNp9v3P9Ac3HIXSilcaCO
4P9wEPg+ykD1qfmtYgtdOSXE3fXhTUwxyHFuZ25tj7Pueueu6/118/EixH+A74UgQarMa1AIE9l2
XjhrlxO8n3tpYA1H8uJ76Oqp+AFC3umfLXQ356V78txDAZCYQ4B1Rk+jrlxXze9t/fBBJSXwQVBc
S9RLPeqb2198S8WnNbZhgYKpkaBS85QXyybzQnGGeW9nVLoC0+16GI8S61taaQ2wPOytprhb18OI
hvM4QuAbiefKWhUdeHg9K7BW2uyPlILfXQy8OTBV+P1UKHnqe+SMa11rDPJVOvlSSoW5Can3xG6v
7gXuUe+TZZ9dzO2CLNAkU81wz7rMgrVmvcsfnLvhrvQdO9FMencnH76KFIsi12XmnVD2+NSmATS3
lxqcC+PQ3/vTy1qg/xVqtJB4J2YWMF5+B1xWoi7Rz9tDh3RcKGN7/T0wrbwQ77UtLxex81QmPvvf
V80fR/1EigLpuCYuGe0Tph0+9ek3psIx6+pHmjGMtKMUgHBs03YuPJj9brx/72/wtX1ykKp0ziKS
gEzzIcReP24aLMyndqccLHq2BbDeY+FFH+08Ul+oW7zvfcIGuJ1GGpHC0lwe+xfQXjrv7Xi5mR6G
qDr0Tn1nzJ7SgdBUI0iuCVeEuXY6uEibnPiDrbtqmcdQY6pzn8K3ym4mg+r1jeTNbvH3bKugemuu
vdqdPJNnNOM5hcqNaIQqMYnV5qL6ClY/Naqb7C8xSVVfWW5Dwt3Wg53pjsOD856VC8gvT7Kh1fJH
xZMg6yLtwohJul4zBp6KiF7r4eiu63RmovlZmNzmgROsB0kDQ5U70k4pU9v39d1J3jiNQMnGQFJ8
IgtVLuX08hLu5ARKfgHcvXSFkWehLJcgCMooSHc6/dBYowM4R60RHXauxbkFkLhqwP1l1HLZabhQ
B5AUZ68QWUEuMIUqhEaeMdy6rOn6jZqQ0+480e8uzipHKregc4QbIv1umFjcJl1fTsBOf+0qVE9x
jxtdHHE15ZWjwa8Ugq0KTSrTYhF6lhCXzkor5RJj6L/IULz9XT9BqwILp0Ia4t91rfLJp9dazoLf
fGBmqMIlZa+rICAq6dxSTn19EYoxikd10hHO/7+vKcY1sPnVibU2Aa0iw4EanrZcPRmbClxqHDsl
niwPXcqv3HcU93+Y1v62eKnr6jui2QM0GtK4+kQRbXhi+mEP5hR73Z5wocvPOnzvQKqhCnQgNcyq
GY9Fczso3Os7LE1TITGtmFx8GEzzOwn1tjrO6OGJ6tSI5EhxcyJ9fc/wpLDgyars3YQE4ajOQXUK
sEh6dmzXGR849pqmuU6H+932zUcKfqYPMKnrDBrNlZVXoLy1oF/KMesQSP+M9XJmkgFjL6yEjlFk
P2IP+4pITCFAPPohaCv7WbyPfoS66rMrzPDyJZ3FE5c+VRx8b7ci8gmwlYYlPMaQ8D66Beky4Uef
9YonOPkELB2ZDUvro6oS0visRjV+APbLuw8PmXNxkGM+OQR8KvdvrAkq22ZiZ8NoXjDzLgnyQOb8
xAD8ec0QcrMHSNhRTiJCxsFXGPrHIz4ZxwjG3V5NjUw9HjRVds+mnZ3CeHEbcyZ+fA0CupVa6kEK
ic7fnif+1cyyjUn4L4IU7IsfUNXQFG4Jtls5L4tlDEPOPKEqgZIHIqeKuxS3Ifmt/Qh4co/dfzm7
Vz54OjiJDN/5HI067JQ8tnnF3V0ySKM+330YIzv5CHRYqfWJ19z3YGSgaIWgbDWLWOM9/ejEUMwV
CDsAhVuHgaCY+rFdd6ieDoW1W9TIyHQ561NK0/ZkHjuyz/LyWGtA4XLsJN0wFVszcGIKAt54enCH
N+SbKptrnjXZ9xqls1YUBmFaWAdDUczQUOsJNG9cG53AkQhSpZMKaLyxXk0qzDvLvSouhCvuonC3
D30Mu/7DTK9sr0bkMt7WpevWIiPy7hCC6xOpNMmstQOTxpDlxDFEd5tIneYwaSqGp6jjk9g7L2aY
yGV33Bau0RHkUsKHffiiOI9IHkvbiDph1LzSijU0TlRGNLDV3pTOb/ozsRzEsJ1H7yZ/mBKgQPaZ
9fXpMcGHB65mqVTP+kGLQod7189bKLWdTZ7gm1JRg10+hsR6rhY8qXIFXkI7qUZKC+DVesG5p+iP
SaPR2HAtJg/6N31PGdQ/6icpiioMqT8Hxzqv17Oa3PXn6RzRv6Jb5ZRGEL2RhTQQjzRHsFolajGl
6y2PIsJqucgSJ87ja65oMR/rtNnzA6wORkyoO1OCP06tGcFB6GWwf8W13GDPicMQOOAZ3vx12uV4
o2YqKtVMsTenQkznfzrdcwsPGN4uPJv+WeJApmTo5ki+EQZTulwxRycWa+u8/pPwmEOMvAM7mf4p
TEe9buN8kVOGqJIPgna/8qV8A0D4kEtNRDr0ggq0jpwzW9q6L+U4OphPqAzqqW9VtouMiT+88ASR
6TqiaHohJgfFebRct06WOJr5cqvkzA/lC3roZEmimicI/fqM0XkDg3TH4P2pOXmg9q+q/cKq9vOt
6XyQQx+zwkhvrecg5b/C9nLHeQoPOk/7r+BFmOe00u3PsEyYRKzLW+LGCxIDJx8MxJH+/oBurM25
WBOvyQkNHXjNEDP5GjRd0L8abmoeZTIMBlaTcZBBeYJ41CedcsCAeC8qADct0Qk6zfwMEoDwxcfH
ENBEX+HxIjLRx9oA5JSXzlma7cJvu10ms5x6ei09hWTB6HGHUibTXc7c8r9iQSN2fwA2XtwIC6OF
4FdWpNoBMVrVJhAIXsbM34K36on/q/PLrfC/mEZ59EgDLuapwAaPQdNvW5RAF6LEQdEpIclitLXm
MyGr/GbeXmA+ZNxFJN6Ibm1iG9iO2rSXzAxQalXx7B4c9sVM4uQ21ZH5pKEwyLcVVZq1yMyABhk6
ZGHqJHn82b3dDlQeMkCw7jUtTsyp4fglKZHjTqZFAGK2B78wzi1spoiBugTzVyvL4BUqjQL5UjqS
mz6a2T9koBvOePd3dmC1srquEaSK0Ywf/yEeB6rxOee7zA19+xkNw+ySFPXLoeDGd9F41Gxfj/cT
dAlpa3JHWVhCwpb6MegPmbnlVUHM/c6hZew2tHeIxnJTRFoVRrAyoa8yBBM5rDgdCAChxTchPnU5
nqPAMuzOHyGmmoEK1QLkL9Feussccn6RLXLrX5GDoCWQxI2T/rdzoSRnXzNEhvjKOWnp0xzk5Zvs
KSFyH1Ra1xh6ZrF/rZQFQaRe+d1ztZZUjm/cQ+LqTQMetJxNY1JouGx5lr+TOTxV531yQEN0Ma3C
UTLBm9VxnVUG60O92cSJvCN0tJyLGCWkXM+UKBDZ7MZx2twpIwhwtDVD3SYYnWIXsm0Damf1cdmk
Y+6WpUgQx/epk3tPkeA1ISjMS5p7eAqhpGflPjHtCe3NTuIAeJKhpgWQ92MBNwCTfSbM3kHff83L
H0oTKR0Q1xm1gR+IwglB022VK3Yjqtkb81bznjQHXKlirRUiOqzqU7WGClCSzF+YL1AgARo47Y2R
dMoOL1V89EwpuDW+iJ4cnTtL3DEwALgw4Xk9xp05SKwl+1IbvWHEUdkNXiIKO+E3UrWe3ajboekR
I3f0ag/A+nMZWfA2D/OuBNwQbZR4PuU9kY/8WmSz44tP71VFLkCwzjtgyAZatQUOfhj3UO1Dp5MX
Cm4mpywWGxxjrOwMgfGySjaMw0M/xJrZdqU5ElWSEGuvmpAYkBbRT0qEJFVKptPYLTGRoh1XomCD
+8BKtT6UrXaj+g+jq+Q047zSBN5ZgeLoYOJJf+u8KSajhqc1OR7VgE2i492yxYNrBjNfgj2sE05G
Cyf3Eu28NlB5whIT82Nd2lFcyavWRPsyLZ/IjkX3WSLoNCuF/fon54Z1jIlVOT2OVxl6wY6j/9i4
eycALxBH9wkCEMX4sFOegMRE9mkeXKWmBUkPgmj6fXmeiL2Wlei6od+m5l49qOLvvG05MLoD5L5W
+VJlSX/M6lJCJX7EU4Gzt7YJcGS8n+hTwYju5wLStWNu3xf0y96kRRQLgb9I8u3I9bJkqsKS0DMY
qpicuCGds/orkjE8D2KTKUNGrP7a0Lwj5SZpfLmKETX11hGYAlkMCR/tv+QkN1TaPrP+OoJAN5fY
aJZooGiyv5/lJF/JrNt1GO9jAfyw80+a4gj0mWB4L0ll6i+ROmUNwftAeb0HSQrTdGcOsS1wjOBa
aJeF0ZAhhQeJ/bZybiDLw6V3cRi454s6xR0VyOgfURqtpZPA17/95V8rdBjdPHBvttaRWsp+WqJo
C5Q1kUB4UNeOMYCOHmYExpHL2MOkbqdVpRULVYNUn5KH6wjsyKzrNFTJAZIWNKI8BlYSaglE4fJr
9XjreJGe8W/bcfimwAAkUFZ9FBRtzjw4U5lCcIHjc26aRQazppkq0aZPLCp7Sazf8UTB4j8idpZf
blYG04T2bnaVY+cIevMLZi+yqmWrvIopNGB1v0JF9kRjsETGjV49/qQikxhHYy85qTqtIsuGWm5k
2YJUw/W+kd/hdPwanz3OYaOG1rpi6Ariwbbvm1H94q+FOGnjU0ZZFwHwanXtCGjkBcnTdonTsFBG
4RxrKCkDW94N5rnMaZyFDQVWgqJ4gjcTHKPkom5L+xWzlqw3gsn0zTUMRhV/obfbufsefjua10SK
XlRenX9PQ6Y1r9yqZAiRPX1Xd4vOXu94srK3AQSKZlnrt3RLPQmkDftlZN8Np4KICWLAUNSjlkac
7BMKQkeNEZSJaqouUApZzibQcsFBkHciDw3x6HsDg3xsmq0fajOtBEjkp0Rl4UT7iyd1HZTqLLkV
D87ko8Bk4DPmFhtxtOBHxklTiF1cixrG2/uF1NfxN9nE3ahKfb5MA/+mo/drS1D6wLW29AcM2cpL
YxtB6gI4YHmmCOLk3eaquNAysOPo8liSQpAUNxSck8UgAUrUxX+jm7eVU4xl1/1w2cbNKwaYmbOa
+l+Q3WDUVDgDjyUdnfW0WE5Y3Q6g5iRw7GARtvhhic81dWpThUiMItEZ/7HD5RrRDP5oYxAEdmll
0SnwSb/FSW36lmAvrShoPjS3ajmXDdUnqMPchCPnb08dnP/jPHm18Lek22n5OH2VeOC/cB/R5d/G
dhKBiWvJoXbkxeWn3xIu7sVO+X3hXFDX2tB0YTkgHmZIw735xhcQPQUUpF/2tdqXv6Wls46vhCyP
LnukXRoqIG0Ru+lb6y/QTS3X00TR7fH8MqJmc/3TDOCnHD8gVschKE/HT7bkwHuHl9lLvbzxq9iA
cSfzr+v0QLTr1jz0KhtaOvkQzly0GSNiq7YGiYZ2mPQoyY8zno7fmKhVeuTRWG96NZgp/M6l1blH
PDQCIxZCdmkF1IWXJJloSd2pq3FT/VZosklHHSvftd3KczZ0BRhoMjAR/vXgKOMQ7zWSFtJZ//ok
CupO7Jvo+bm0EWQOUp+IMZNe03n9YZ5iBQAXKMbdOBbPXgL2iPNfFnycEEJLUHrJePAUsdTy33po
GpnCVOgRhJAJHR+I8EeRRdugc/DU5fCllWEepnyc/qsPQsa4GLJHX74Gt1jQ2OwcXr6/261DEjqv
02Ipnt4f6+J5QP4FMOlmbOKD3hMpDCPTMS+tN3wUaC+XDx2raV3yhp7JT+3v+liJnCqwuXyVM3e3
x+gFdk488TVJhtw7T0P2U3PBPXg9UoC8OKefwNbhF0AMLswwF+gWx8qu2ErUDKMxqbabuXvPiDFB
4T70SkMJHqwrjx8GtmkrR+CV7LW+f6fJWgH2yJSg3hWLq9TqAUPad2CkSJJR4tvF9+nBaS9FbEGl
yzBtrCrPkcCwZMHedwiWE7zo5DCh0HtYQv5izpOpiAg5LFHO5ql6WFv0tuiiSFCLFdXHTJrP12lC
SW+/FoaHqnksZOxhUFUqo/V6jnxEkbdcxP3dzeUF04V2KyVC6usu0PSWUmgfdEGHyHhkl998kH9N
H9ipOjmWC3aAGbdUqJWvMGKuOltr1caK5QVQqaFT2FTK9qI620lnzZvdcrPSSZKK2CcNB5AYOQA4
qBJ49LzoqrGogcreBo0AiXMnIL2Q6c6JMSQI5qxBtsm/iz0KQvX7guqzek8gLH351eBcfdYrIFsV
eD/S9sD1XHyUuczR1cne0c0D0C1J+8r7H4Okm11MiiUvodKA8IHz71S422sdJzspqtIZEv5p7gKu
hWiAUy5RNwUQvucvwDGYt/d9l04wV0QohgjEZf/Fc1OiWKyLlBBVdsYd2YeS8MQ89k8UsqM67ime
7cSiTM+kQRHp6G8gLCDq6tB4AnF8dGGn0pBiKxzD7rVqVUHYnZFCXl87pLwR5y7cG0fToFEOjSPE
WX/4PPXj01T2Itk/CXXQsEMCmAUXo65jRlBGHC4nE+JqphdVrU38almae9hOcQyJr7HAFpbgHyYn
L7hTSHLvbQM9NkRvDWah+iyr7Xjo91h0mj8njCkUBrhXdNeeDjzXK4BHKr/OCFBp5LLWxrV7s2N0
UB3H+X1zzJ3HNDz3ksbQ9sTJk4TA82zhmkOnM2BFK58MyMOxARAo63QVVgpMIDOyZgB5nml7rwlH
KFY22YNCGPMdhGWgOMLN8ktMS6ARUn477LbrLCsnA3gbuzZhqULvXhYShyjjQym4hamUZ6p9ycSP
z3gRiA0+MWOYFuj1o3X8mTJikYka04J97RAE2BRPyFXVzuBF89lJ/yMvRekYMoqRQcFB2zWB/MEQ
mpShp9DAW503TfIoUrzuZToO72/BSyXYDzg3YSrOaEFm3OjiTeIK3/EYob5X5hlq5wrtXRlHftfi
IUNQSB3ovkgXmfNZDWk1nCWsRLYaCMnbBMzEdw2HD4CKFbfV/j5v1QHAoaicNuW4mPcg5eepzKmZ
WkNn1P9Dyxambmq0WlnomlhMnIFE3e0Cc6DOQF4Uc1h64+8pDwfHEV6D4+WY9t1mBrIjZl6JWveU
wthCBhDjptkpBTRM65GEATTrzyoci5WldK5rckQVE9fDb3tpJxtGAE+O37tBlLsMs7ZgSA+L+K5A
A42xRH/N+R/TAEH32QnXBseMKXkIUw8HyrSsQPXpQyF5omhgR4SriM2nNM5nJpk1QkdBQTrJVK2F
2Xm6ngX3Dqa/o/aMziDuIuZAuCwfYRUyLh+ldwhj2c6S003lAYngciniToBPFE16H12WgtsS7Bbr
QTvdpd2Qz5QGHlqwE6A8YoKYc4d8hnfujhSVyTpxgwmXAttB0hjB3XCVBi9xDMVbGCWer3JvMTKO
YUxXMenvuqTfX9d8QJvhxHqVjrZm7pEHWHrPtHFaPXLCUbtxO2URbMk9OpgLqcj1sZcuCOgYJWdP
e6mjwCoN3R6VdGLuMMfTOdLxzWbh6Pyjm6AmzDM/o6FQCG2Hz/Bpx0fQQoG+OT7C5BZfOv3Lkxju
V5bCn2rd4Tb4Vnh5rn29f1DkCMOkgWjbDWtzmpbwoss8XJdYYqRbSaW1vzJ0GHq3s2KK5Ikc9MZm
1FgzacYjtitNMFGnXSzs6OiPgVoPI+y3igWa3VtkJRRwPfyHb3x7sYYjbHMcmJX5VjGkptVvvkTI
QCNQrPLlUoycdSKYWO2e/LMNjKSa0gR0o/YTT3QjS5N3njVYhs9ytJvQkJFKVlfI2xUSi3136uCW
W/nHzchrnHEAwJD0T1dgT441Gs29egQjwdqNymLwN67V+xLnnSryNXJgsdkKdqa8QF906S/erlan
FdzcXQpFO1/gjNC7G901WnbV05QAJHqPotZE0qdKAoqOybqB8uw4OqPO7FcoGRsDPbTvqXg8Foq2
A2LoZS/lPV3ezUJ/wZmUxzqZLaX6lwBXJZljUvMSeEMvggRAA0BwTGkU4CL4nbKY+fDsaiwJjhdz
+IcG3NJgVsclXCsl9L/Tly+rnUGvrjEuLgpJfpS+8PY7CDioc4TtqMPh2Sw3JdmL/EXILnmuAHB+
vuxel4iYGLPB/pSbGnR1rZiqTbDN0ykcaY7P8AoCCw1VtptbaEOWG2C9JGTI9XrdQBxMYDk3+4HY
/dt62iuY/t+W+GfAZ9/MLg2a/oiLFQXY3CFnY2FUnX33HhKtuRscoowadceX7+elowYzIMVRgP3A
q8J6k6VMkm+Cl37yAeRB45jAShC6HmKhq7CnviLJpn99KKX2DtstuEHpK/VmW4r0CzdIW1c34y7Y
99qHiWwl+qjIsQa7zdXXCFKYSszxjws7PMS7K72Ohx5dxgwkbj2A2PWrMK0+UTXehIBL1Brax8mv
V7GTf04v9251gGRbaqiN5Zso4xqgg9jWSl2FtF2jHxTlAiGK2g6hrBSN5cVsKfRa0YsyhDxyQiFq
ZVa4q/qpzwwZHU0eKGbwO1Qu6csrfP/QihuuhWS9HqNhAc9XNAPTN3lecj4Yi3/ZjO45UOZZG8aF
PatItl2EzcX+hFpFW17wvXLVPaadYadSMcDYnG02qAUW8heTfrHQktVvVnXoGSrnUDF16MV+fvdC
Wr/nmIdX6F4QRugkQjhBCE8g8mUOPTtmyqQ3XRrTl1gK8p6V12oZlCBgiVT0YGlRNihgzRgdNmB1
QBFHOxxx9LkF/5LNeD5qm+iKGwGQ2sILw9tdJYqXEq2TlJ6tMXZGKmP2SQ+hF5PUcfPR+9jPcdVK
AXBHqR9z1us1ILXPFDmoQYkingpEKlI+mzORUYxbD4viXjICeK2El+eDZMTpWIn6tFcCUy/e9xtq
FBAVk8hzeW66bH5XNgWhk1+VBJaZVuo4fyAbCRiIpvVdBUCBPUOrghVnp+6OCPe7Bc5VLhnVgSjs
fZ6ac5i7HwMZtDul9k8x1mYhQMUFClpMNmRunKICRST4c0uw8pUJRl+uNsTWRjWrhft30+gdkOvY
W4o03HCQvUxX2pnhsEfAlgZha7wchJbepYQ3ySe1Bt5snc1WzePyun6B8pbN7bNJs5IQG0HdiRth
hROlcD7ixT+n1vTJYSeEAa0BhSF75Jkh063d5JRHsydq4DdXm/bIcNQ3fZ+lF06iELeuSqU8Kd6O
X5IriSe/A79jj9aYNr+zus9o/nKafv0Bx+3/bspCPXwNv/8o9j+ZvcjxBnTdzg0MwwuYWzTCvjPP
Il6UQhk3u49j/EL5xSxuw0NGBrxOYOsNneNzScdYvt3AmYDJvOYmku/8thhXZ+XxjTgmRMgapRAY
CXHQz3y24lVXADIkQsJKks3vQmAhFr7kI6h+omSXqGQBa+mhM8v+WmZPvsJuSoEAOIlAQT6Jho+E
q9zM2kmZew3QT6jlu8/yDnM/cWDU4y9aXG++Tp6zZGAJxvrQHotFor8WXGkkS08A7SWNM1dh3dR3
x+/S4zgn3DTHuSAV5rFXPL1Rgoyqy3ffJBOVzsQ/CHdJsjCU3wNK71iJNVonaf2IIgtUpjakfmTd
SsiChgMFt6NSJvG9YZlvNFdCXfJOwIgRfn+Zw8rSnfAwBUc2RTPoqiD9Be0aDkbQCepMjSO/GRGs
TBaJPfoPt25GnriKai151rJkfM1gll1aVSDt5J78BYCyitM2xSaDtb4TlkZ0hiJydzhRegpUJ2LQ
nXMQbt5kAwPkjBqW4xZEmEou7EK6qBYz8klDYEjrxUoAwbaRBhnL647E5sUq5sb8uq8/8m1Ev+Gx
yscx3tPLom+BFGa9+vqFtEJ7ipsC+CcT0i2t/PDHcMZj3lhiQp8v8lqKQrwxxyzFrz7XbEkIdarl
4eQo4K5H3wUrDXAck4vUNYQukCB30lTpFA7hcF3Hf8iwjxZoEHnYQRLPVlsbVbN6YJt5M5oe1RFu
hrqtVIdKETsQnyWKCp3OfLuNCHpgKbOWMkYOJWLjPnsrSKcDZAFFBASSXMHhgshGpbDHSswl5mB3
I1P9teOWFDJ1diS0UjEJy6QdWnnOMGUEd0WCu8CTCz8fUQRYaIDIfZAQmv2V22dOh4HZsj1h9A++
h5T8ZKIBNET8TRFiwnTZedu77ox51H2ySyNZUhgv0j/QxeBdArCchlPkaTw2g0aDaEJzaD/dJt3O
VDO4mTm76jp3wbyjjsdfoU88wHmNo8TJAFokqo2/R1tsNg7CZBMnE+Cbl+QsgwbYz0haWDIHglBN
WGXaYownmXqZjhA1q8d81RlanyjCTLSUkXb3Gtf6lnalK0m7UYjuS9EYqUnryUMJjvFcEMS22AKE
jgmWDWCPhjHcQyr6oH3zUlXOFu/yAC7C5XzsfH644f2d071E3Q4ApIOnTCpr2B3pe14Phb3IV3cq
BsfJVCY5knYFJ7AEkb9dcACzXm8P44Pohk31di4UXj0u8UsWBTJ4hAafuvxgLLWi3Wf5CCxqOZ8s
6IXxynWgb6noU9510sm1+55KLoMfTkMeUJn0iWEqcSRnq3JqliHOvfcDrF3BW0yP/iKq1wQhlrrF
5G/Mix9x5GG6yHAhCLuGD9129wMqCXBgk7S8Ce/jECsOiNYVWwHARiF1zi6006hkiAvchWUOP51p
EyABAV0TK0nCkFxQQ76qIgrt7aJhqbfEBoQqGzMJenWYM4XsxQNGGaeYrlpeLiGdHblemdKT8ILj
kNp2RUHEQhiUgeMLwzTu4ZIgogG++WV8huQE0bST3lT8NV3mv7/oSoDJwOU7IXwl1YBTPa8WpKUZ
dPDnrdN+Pi/fzeAC7p8rN2TLV/cnfrcPc+4UhGP1ZWRxirr2d/rZ3cbJ0Sv3jsAovK3j/+cEJXM2
0Ba9sAWHJ+qg0Qd+Im87KwuIZ63I20mL3oLn2E6tp1f4B5gN8ncdxoivHRFtFHyCBH2TpO2vgW6U
iYv8C+kHB+Lx1cQ92UlIQgIs2Vh1SM9rqwC8T67eQVnq30rLXNT66CKHessw4sW6BRT7cEUyrcRx
faOtvZEpp+Nnl6cTvtNTtIhiM8dzqNUCj4zbsP14gr71hcq4MFf7EqqW0xjZpIqQVnhwhC2Tvtem
SsX450fVkEAIXj1uAaFyqKFEIbSGhw3IpoLDcw5QrD1YcVUp4kMSEmWHmLoCw9voz2DO44KFZAPu
Fr6an9Ajq8zasQ6RM7L/8Uu7eGra72z1FGyKTSX8B6Phk5r2J73jrB7fnq27/0v1LroWYkN54gEs
7qDA7vT5ATxfOkWAoGP7z9OGZGhXwRqHRtuc2dhUzjFd92EXQ1/dY5BxxgRELwyCzatUcAP1MhOV
z5fjSGhHRLElZXkZcJYuFXzYdDv29CQ2PqHyMMwztxSNzJ6SV6LeGUis9I3CLLdqKPa1/or47lGb
x1MTqfQ7c1ZOW9tRUHIsZEptd69NbfGXuR9e/ddH4F5c/iX7hanhakkgZTsDb8+pdgLtMpmEdORb
EQ0bdF3X+EaJlwN3Gd+NlYtel5ZrP61s1s/DnMKtdWWrb6QEI4Z3nix57QIUayNvyEhByQgh0v+7
lvP7M/6mosFjl6hlEEy30CKfq93yF/yka1raRdM+LshP5es8XmZGTPHHEXLZpumNpluJFbk55haE
Jy9p88TvVqIRBFaFiA8jH8CLW5I9kd4Avqdbr8ydJj/D9sPug+oagXLLNp7iUtuTqcAXPSC6JtGj
EuPzTvUvUY78Sm26MI9UP4/wCk5zqwcfesa9WiazIODs4mhNJZqiJ8Y0TWiaJrCQwWbuY4nHN9X5
6UNo72gTzMzz5gQMt+PV3NyK19vAqwt4w5MeQgd5qqiQVYoUDtqdNFPNTWCXarLZbGABsWuSiTfN
ZTnPzgekfBZJpSPysmkvcKnesWP1eGrlOjZQAWvb3wJKHOGEF5I5zpSofLY3PV4ZOpH8fo0cBA9F
btvjTZtEsleiP591qPc0xPEobw3IJX85v98Tgz1+KhYYaYXVzrNsZDmWlIeeleabSWuDNaZE3mkf
j0SCRXXvSYcJM0qhHlfhm2qzDgVKhvuRo9RG4PlbDX+G1tuQ8UWyBMe5GxFUq0PHvSSKqAsaDD6F
lxm3pGWEqUM5CkbD43yIygOV2DkrDx2dBf3z4Y28Iyoq56edz0Hu1HkG4Oymt2O+WC2Ea38XtYIy
MbyznPED5M0BCmz5I9ajB6PPC0/zWDiSu6aLIm/N7uOBISxDUYZsHQIuAPiuzYVbfCQdbsztLnfH
bluc8sJxlN5etzLdYhWd0VWTbNV+fVPku3BCw64dTxdJmh2x8+VReCJ/StgF9+Peu87lmxvSlWPO
+MNh0Q8ZJ7Jjzd2HNzEepoZa8pT4xtUGgFAWN4Ikh36nrMUb0t7T6KPcxg5a3RJ2hiQyYXmVZqhe
mwGRWbAU1XU9wIKUSLfyyFUAwTf3ddHSij6Lcu2H+FB2T5jT3jAuWOYYPD6ZfIIdmYaiFuRezf9G
YiVgMuHBUFbmT/9Xo0q+cePVx1urQ54OC05RXCkbIGOUevaGBC5l6vhPEiJZ5UoRHfqe0NFxZq7B
TL7j+PBaqM1kVfOen7gO2FfGaVzpqOjpPm1rY64JLnhW1vCEud86c5T04l2boyrpIb/lCcQmuSaO
x9TE5eEJnplm36gF9iaPWnzgCHGGBFdJvZr859xqLV35E6vXaUOehHZyLtjerW2Zv072iACRndTm
aWcdfn1krLutBhbJLEUBIvSQhNUAQm7hBfuAnwpmKevI0gmuJLzKWBLKRml6o9C6MbKNfTo7fh35
Mx62OLwj4Wrku90j3ZdWGpFkXWiHLoiQPRe63lSTE0/ZGkJJ7UmWh02fnbKFIAPEdz6yBc5KjWz4
CgF5bBOX648fp++MrbuLRQbhIIHPmUaPSy0vG2A173z+3Zm6EVqhwnwtZ/0BdW5Ex3BJmbgk06/i
8v/AjhcWekRVvqOGCFYDVNPSMZAptMfbeHHkTTDi0MX6JYpkVJkSaSkLUPgWBdKUhsjP9M5EiRWU
fmzqxQ+/SXIR13bTE3/6D0ilL6AfTchawwyeDJscvWfRoyM9bssP30PP02QMSSfqSCux0Yhfb5h2
EIJKImi8CGfsaC4yx7CSjGvAxae1lYIJDGfJSpPe/cuHWhB5igWLQNM2v477AYq7wepdpDX7poOt
C7Nr4KQquNqblQjFnTMfW4zf3MW/ErOljeI0wFZNVwrnxzAEUwCb6yr0JGnQnevzHVHXFS7t82/u
mq71hmYT3YKfoVfe3jFXB1sbHpWEqSx9jRRw6Hs2YvT6xP6To3HgJjqz+douo8D05SR3FfaXl4ki
hTjAUXZrsSD5qy2DXWBNj3e03JNy3sJPVeq3unbs5M4KudknfFI4GUM3pw03v1riu5F5fV3HQxcj
u7b57479i5D/oDp1xQbgapk/rTOfpqu7DMS/MJ8StunCOqn7xGzr/JzcM8CJBLXunt2bch71uolb
4HJ+dDqMX6NnTE4KwFeKp8HDFbq7OfthQK+kyld9MncXwv7FOBNkf4nzE/O03Qam2vbMVXl2u6y0
KDXBjYZWwng9wJNfglXZtgIB09FAby8e0lXgfOoMwpzdESRsjmPQPKe6qz/mK8qYHH24RLzHNwpR
hQ2puwqQ3olFo9HdevbAS9BkHIpuxrq8OM86tWpo5XkJkVbAWXULD0qCHPlUsCZCyASjG/2Dm4Ub
DVaFMbKGZsWOX7oxGF5jS5Z3KafOBtL7IIygAnXsn8nr/iZ7GTpXKFLxcjAP5icACLAQ0GuZC9Jx
c6sxvwCJx0EuhQzZz8cjYSIlCDSoLc0Txda9QxuK6sZiVkqsxqGAwB4j+Frr//UzFmn8mngWxw9K
QglZ17zi4soBPSUNh69Dx+bLvRdsQzd3K4T7LA4KSHHM2hOm9bxhbqkUKqw/tLuew1+HO4mpaE9Y
MpdpwPsYGikkSLapitEZKL6Q33R0Jd55Bt6CkqZYanx8N3sxIJxVwv0rlqSdJebXQaj3pbH3WBK7
cSH+j4RJ4xZ4mffG5vQTzZ/SVFc0qi/l8SUFpAU8Ej37rtnjUWzPmt2ZTJBl//leyDSD6OAQeEVK
nUq1zLWYczl9z2h2btWOvSXIyrzVrnY5cuyaXfJDnYAvgCSDk+lGr/hHp3LVTMEeq2Cd7sX+rTzg
u3UV24+XaQPd1CLqS/5hfLcRRrNg6+o1Pn36JNRJ30X1JNWDVL+h0p5tFDl3bkBXsnjwRtAU++Ab
xAZpGxuLkpYgbWTfLsw/XXreaTeL+mFtqtfPRfGWor2MYccTgo1I2GXl4DUf7X9qplJYDbgQyNXh
NEPut9hQsaXbAPf88A9EQoo8/tmxGKsWtBfn0BO1/sm5elRqCorWLw0KbX+YgtFK+ZvRHcLxMnBD
BCgw7klcBZ18VR4o6yK0WGfGQ77sXgyx2OjRTFPFV6prh1yWBWpBIOcDOwSK7MNNSsTEksqPKYQ/
shoUwBVvRO/kqf4+HbcxX8scbhRm0SqjOz05CJPQv6ZfZQJlVMuv6k5cDjhdgFEFDSRFV7wUknxE
Wb/P7C4oYXjDvnwTZZp8Y54itdt9prWSozDngLeWda5ZxoLOS7cxuuEZka4GVelcFiefaEuKycx9
GmLeQHTWUj3Vt9IxpAy0gJ76eAZGKggPOCsQSNnlO4VaPr7LlL3c7wzXv1lyOI7sYqPg8+dsqadC
BvM1aKCdQzKMk7WlNDLHdKJZnOPEcWGTV5N3sNdMLTgh6DU3jmTweto2EygLxFiKySPKQGw7k2sP
jyMXVMLKRxj6EdkAcad1T9TMhbZG+B/mk1PkT/cxFJcCm87fs5SYZAl3bzFndsKIxm8w9kJqTLK9
T4NYGT0/o1Dn9m9r5ef3P/AdE6JLskuafIK4+TC4n9YMxRcBM8duzR7GakUl1cs6Iaxt7/8Fm9vL
cmv99D/hoHGaeu3JeDJO1sNpDZ/1Y+Jqar79LSGv76BCcWSv3R5t07Q4hWzkKxyRsZwMAQkpzFsq
sA6HWhJZ4jO0WPaPVWBBw/UBRJqthodxhxxrNMr2+C6MC/wKCXxzMJidyuQLeftChVEOan8TVyPB
Y6quKuwPz7OzIt216Adm7q+d35b1t/+H7OuTx+fs2FQ3TyH5rBLWWuPxwAac5IZb6z4lheFzwRRY
76nI8IJo4UNO0l8V/fSRr8oDNUm4yI8zVGWiL0YHIpdLe6eD2lQYPGGbc+SMeYUsG9zfsq8X/+wD
u3UkIODdCaNTQwnbChF/7bm+L+M3cBsbR032XVqfoBtyR2HQs7V+7ZBH6QPIPZ/fqIXRfhb/QET5
Wr9YvmNXVW1aX7nK6QnATMnqeu1Gw8MpHOkkMkJWd6sHntzr8cnRM46GvsZMJ6v4cZYX+sgPvEiV
vBNqJc55SWG53VW1xxo1QeHpftlpikO0HRt6OUAB8XhTchF8YMoLvBisFVcP7fZfDFBJXwWCvB8s
t12iM7XTiaklmGjobws2l/rCH6Y6qGAahAt4vfT1ZAkp7E6ASCJ1I+9/wk0GprY4igJTq8sYTjg+
of472VJNn9sBRomHQXqKzBcPPv+sCj61LSuftgSJ38AeBFRFdvRTqD1efYd/YJQ1/VWd7ISdM2Yv
ICLGWOOOXG20FuUHZA4ZoRQHxw82QUwUU1n5z36Juse6kIRsbGYblXv7IxNPylEvVZqJXTJOoE57
aYczA3+mv9qVfdlT05sM9KKz8REC5QN2CXEKcLLkYP5GSeI+n7TbIh3JgqI/juy1TKDwsiDjnJI9
/g2Lv0qn7zPvaVbRofCY0IZo/Y3b3JowixVHpUOnJou9OONvE9OQ150HYaQerQeSIvB7dPZV/vkj
I9830CrcpKe5hMJhfm1D6G7wM6wbxBGpzSbCFEzk6N2nX4tU/7CWS2mN1PfHt0/xJsvDswkF6HC1
rgxHm2uwQk5MzJhl0iZ1e3aLikgoBjELXwptNa5PytReiAOAfDYzOwt1FfBxbd7PHGO7voIOUtPs
fLFTysvRtycrpwCauaEr1eSVNAG2q46cIlRum7vW5mBDpFCcthOBpWBT3X80WQeCjg04VI1hYaPv
8pzzhncAEfLSAgRmS9vSfK1vEiLGEviOLOfsvA/gFl5NkeQxFvtBTB5lFTlXyD6nmRoNF+1FQqTg
EXFrRyfLv4maDCQScz7AhVTR7ze8uX/7L+FvWORjb9YPwghfYlsY14lCERyMhYF9DldgWXNNGxjJ
WetpE/WcGP+G81U9/cLXUbYD8/rTAD0J9o65wEzyWvesHodqgezGm9718km3UvdxAc1oMfkD4ree
vP7HMqwrB5Et5+VPy5CP8ILj2WLAy7xzGwTwdV6ZE9fn2/IzlODgGd5wFhV+hD1wxE+mZIkx2NWA
EC0wpicUhfZJsDAHsxZIWRwYXJ/tChjWtlRSlzfTwiOqfNL6zcxSEpeLZVfeL6pHcKuPNK66lFbF
2DYPkADV2wy+XwztL7JMbROsmFaU0Ha1YePYK93bGnczfpTlcijqyh0WzIKWKlBraTRmQrWE8O3w
GYsAQhv9feUSsCFjeZ4izI9Mo61luwMo5P+N3Di9rpF+6J4A7eR3hP2sTpkoZfmHchu2deNccvXh
eeYUz6+whA8lt7hoyBRLMR7LwCH125Xi2rXSX1U5vN0vUO2j80dE1TzfyT/Wg4kXUSi7OxRg9+KV
gkxpmEwrz+KxZEwpF5ht6bq4hRSdZ34/e8Rl69MtDVoyG+Nl+Bpe9tvifzTZpt9mVDyWn52xl0CS
xR4umAUlu8ehV8BTRXnikf+PNzD3kCZO6mTvkchbk2r65OYqUpbWPU+hUsfh6Pq1qu17mJf/GyEA
UHirqkdbgxaabuwoAf2I5ZkztMAJjHF6nTum8fqJJuMjoOH6HP1lpi0C+FsZfHe92dMt8tFpwvpE
YAi1Db0wPFj9YFA7wKVjiFGJCQ+0nqDSp1VhtpH0T3IKdWMm0VRgM5D1mPeqPIiNZzsTaaMUjPYc
A/b+ej6MVEHsT88v0TolumbTIennfmp6cyQUXuCDywYxSqQ5fExeJbdveFP0/xdiDudS+VWbzkcN
J36uMMTYLRJky6F5HXstUp64VOhrdeCOvkpkj/yZRFlI9zM1Nn6PshBT2DMy+vFqsFCJ+WLk5eaw
Z5xZUegRxqeJ7eRPykqB+whmvk4g88hoF3eFwqFbIJ+d7c1sjzqbVnMVEOgclwyB1p5iIoS/ZfIr
qvtZz51tDYQDuta1xnp1GxFZc0Iaphi9V+ssy+CXhfDTJlUa7gci5f2WItM84JihMQi8iHi9LssN
wbXzdT1ApSm0uLK56L5y6QDx8knFt1cO+MZjA/ubc9V3m892lkO+7HqT6met+RKybrwGE31f901Y
/Yk8SGFTXTN6sOyiHx5GepPWwI38TDSredzMxJ74GSUa/qoQkQBhhzjprOlRp1gcWEkqpbWc4vGP
Mb1kiRZmZNwmBjgpn3QHmFnl9Mt7D6i3346tA+LYu/lKAY1T2pEj3X7SmRGhDXOiWA4lebAgh1qf
rsKPmGrDJXyIi4TEHi5LagjjshnbHUdNT0ReRnz7iSfTPujjazt/ZsDI7byQyARLnT8iaGQkkjae
DyRhpjDa5GSvekPLnOBBQAfyF7hZgsvN8o4VwCU5Q4uYt7upLMXZeePKSnHlibBkgxNGX1VsWlda
N6BJDvAm4H9wRzeQYMkYlCc2ho8BwWZJ83ubbeH2p7n8eHDw3TkroYfSrP3+zzfPDshr0A6jVKs8
TMPv4QQyJE7MUu5Y88RmbP5yyiZ/KbvCJYj3yv7AqgQfXo0m5wSI0PyEXHzLjH2CIVXO+ZSvdZcA
q4p2jXXQILbgRiQf3ip/wDSUdrwgAjFq+z3TdRVEYApr/4xhIo3wPxgNy8wpU99tDxaGTRNlVV6K
w/kp5fSwvn1UVAO/ko9h+G0K0Hwqhz6wMxWxqMIxYxdUgWOKLZx/nAq/aky0gIxcURFA/lyVDA1U
32B54NjzCrGRNJIki5irhO5Ts8CYZbAD6oXjf05E0TfeMML37LJtL/45aUNJMhbCrzi2GmY/V3y0
N2Sx/LqVcF+Kz8Xf05Laqt+tpjvLk5xfET7a0C4ZcUMgGShKGJbHB9wjbR0Vb7v4rlBAiWXg4/Av
Fod/2yb596pxdgDSp1bNR6eXSaDuo2mKulHiRm2E2rhrRUAyHdscbHfYESZc3YoILSuQk61JP4UG
9PYLZJ/DZA1TW76/+cvlSrVK2PwHc3cKuvpI0aBqlkqd93UE0tL7b4oHUM7QoTp6uZAl1+1u3TgH
Tgx+mquHasaH0sW3FBEAyzSN40KWRZsPP92nRc8EiEQqK0bX78lMiCcOjy6I/Xz9AC3oT+iioqbq
Zj2Cl0fGgxOuZB/7YqhIrty/QhbsR0FMj9zA9yk1HdryxSOvK1XrLKpvj/RMG1Y3d+AfIVgbtr2t
GfxsgXARQ14U/8sPTFaUdjH1G/NcuiVFRCLVELkEZ11t94hsFR4U5GDHQ5dnKOcRBbFeqk0+45ID
OsB2KB+IReY1BGScoB/1qkdBmSM7jVciOG24M1hvBG9G36TinSd37AeFPzj1bPAMINWVPsSiUmVv
TYZEEk2NIeafmsudohKfgNhg9cNDFAJb4fMxWUOeosBQaONmIeZ0VbY6/Qp297ZHmeC2q9/7pnCN
tHgROria/q10AfuRTr8ad2y1uq/mDOUm1TM7NJyg9ISycf5iJ4VcJWFYwKemUU8Mbq2Un741ZlQe
zvrMSEFshXm45xYNYeliIFLjbc03dG8Az8TAH8ul5EEzrXPIn2rSYnHZOehnFmUIQKTXMVo+VKSK
LbQO0JvzWjZAgwn5mkYq7gNfDmo80X45Th20GLvWOnch8dzXGUYeptne2lh0hexadwFVY1Qd8eDw
ztXqUFFzZlQro+QAi6I1ogJWTLHTGzl+fsjKCHfpgJCLG2gIa9PShEU61ROVtFJcNVJ7fsmlWxv2
N4R6TrusjkjAjdEIDcQBiSsNI93Z0FxoXRORlhDmktjsIMKfGYwxgcs2VPp9mXwXmn9R8M+mXPs3
rFcsbA/rWfArD1BxyYG7EEQEOWsWhSiC5BNPzD9N3UFRFh5/nH6jq2D89OgnqivEnMpiDZT97kSY
BpvRVhocHKd/XBj0R2d9a2nyKakmgeiuOd9RKpXARcR7ZR83oTi4kbPa1z7i7bi3qvjmhPO4LWgw
RE94o9V7WUGNmlxCZkZVFZTSyDX4KTr6jc547YLP6AihgXT4ne/INafjoCUM//RKHXTLY1w3fyU2
Mv5VZHnUP40FvjTAQdEtnosO+pP3FnyjKNuWGhjfdKMWQXw9SHThDBNPsHhUy5SStAzBXUUQLS45
gYza4Dg+CRfpEvf01bg/NBQaRFYAoSzah1TO+pw3zcTLwIXz7PnuVnpPlrV7/U2jPptce3OARmd4
QAv4Uy5CV9Zwsjc5gj3dXw6BdhiWJ8hrEmD6/tHpCynKZHAdRR0gKIgLacQWVLkJOaZ3CrwVdFt4
bJccxn/QIVIoijXDMEb4C4Z6O4AkLgxEdyq1KjoGVIKLHPfuD8bvBilElcEueSyri6HA+OCLr4gX
kBHsmHdT3qdyhCRR42D6VDYBiehvYDvvj9uA5sUCDg9XiwVrHK5B/z2zKKnDfPtyYEbLWNW/Kr6Y
uZ33cxYfsIhjfhTJM9oiCaXFtNDFVO1LCflU51MAxAzPMe5Kq1lC5TridonQqYovC2xIKqzTMNzZ
FzpA+BL/sohzjfyMISNB0gUBrTZ5qc/DSY69OSD3cJvrAT7XX+JgcK0WWEepsuA7zZ1fB3vonUZW
eUEb7U+91LxWVrZf5yqzpeXdCLofgmYS9ks1PWqClQWZI4frQyFHIobYqH2fyZYeGdCkI1t1RNvD
aE8ML+o+pNHmbJR7yPz+aayRQpT0YzxKZLnHbWBvgfmnQxcZZVwAfPeeNEoWoHU90ShSkopU8/J0
ctkkPn5tkiWsJmeBY6j3ofOx08ZqIJo7QIfGG+uNej734jJix7Dix2A8e52xgxhsbo/R2zIXzF+y
3xEByxVNkMWC/wdoJp1YJGeUfeLQgmjPpqRk/L/VJ01mV5Vs1gDJopVAVr859FnE7WIQmCL9tbLi
mOGc/PktGkFTp3M48UXYRYDectVmYLvLwIfytlBRInttFcC09zVwVIIIM0Taa+QwXcLTvhAswYW2
wf+VrbYg/2RD63CW3J4kncz9D6/wsu2NjkLmnlhGubesDIi9LLD8qipDP3TzCTUybuu3vomxn2Ee
ec1tRDTXF2vPs/UG4prhvfFiU21I/nTPdn261V90BVvCqzBHqIhXMcSeT3V6692JSubxcQoNAsC2
MLI7iJ3BLwnDIylkT8OUajWSpP/gAhacaQE0BhrZ3P+1C/8s115mbq8u/LwF1e9qEscA3S/9BhNa
mSHP7QycZliBBtRFcfFXSRCmhFp7vYcGHBymm5QhPnjkajlX2Uv0SEwRvCdUgMepm6Do+PKvBa3b
a3nTzNdzRrMiSsMNBdPK9t0MsGr+zaR6UqLm/uBnD37NND85edUR9yMpLCrbnr1zGSK5Xh5rbgV/
TMvBHdcPs496MfXqhn0wfKDLN4tBBiL9os7EFH0ljbcvBrlX12q3Ugg2KtUdcqsLVmW994s5Ifqz
phy1BRVtp6qDzp7uaIxnWZadaR0pBgR+pliOQGj6dAUBmEmXrXRC+VUGjmDvkQMD6J1N277WTbXO
nSLel2rpyoNg2fu15VehdAJDB0+oMumgt+mdF38Xou5L97Y9E60RsYkBaLmSemYb05ZmYQJxlkzE
7hmw1OjUliD9Nh+SUK3OjPEFqwjLi5XPHbkEEFefXMNpK63iPvHDIrxc747wr+1a+uTQ3FJJYP61
JNfjtY2agQh5fJnG5mmn9hIsQTVQ2c60mck85B/itlcp2V9J8h33dkRblI5LCiLMEL9tO+go9cUq
IaKDGStYOmnj4+NIiP75r9Zab0k/BDHuRRQqi0Hz5fETaoj1paRh4pKRc2EpSQLyhAevIGODMumm
On89xaNC8PHKO24pOOJj39qtvy3s0Ac9sSO0wF73iZaMQ108igsvbKnWdl8uv3gKuXVCbuSJ/h5M
RuXHYNJmaVfCAUymgD5RQ69d4SHEAEli9TlnKXqSR9EY/USrJNCoZsvq7rY1rCBREnONsEMMxHwC
hi5unh501YnAVNXXMN77SMxvP70Y6G81qPAfFHF5i70F/35mFJ0860McMfVoUixyWjZYdtbzrCpp
vDSInrbgPivBRwnu9x5ZyJV71RCvoKkei2S30/ReOCNElPnxaKLSik1hqhSeRr9dOxr6QStc0dET
dD6N0bvQJRLJXwsJY07ZxVECaWiHt04Ev+gSTy6vJvAe9GWYI+BsaTvozXtcD4kqjeh/Vxd84NDS
Y1q+UVIesuebBCwIl0SGy2h5w6Eve8F789Y0Zs1hLSZnzen9iskhtSOsdduZnmnH3JGyUSzOLVq8
SQbip9k4QhO9a/Dx9GGOZNy6+Uvld7RGKVfqrxsagYj7ikgxUW74vk4AY6obGaKHZRaJA44vxqEo
4p4URbqiklpJVFnQiXgyvCSiGOuLUgVbpUJ27MasYY73NewlQKqVycqnoJXjtfZ/RHFgdByE0amt
8X8spnwxdP04clQqI0BinjezEMNc8pS3XHxWs4/bnsZgKDeI2iwoKIbYPRRuV9Qv+FKDroK/3rom
p2sX4amqW+NPrzdYeqw6yfLUYelhckjEw2dOXAz02QimosJrFVZljl1ME1zeJCWf5C5kICWeMCLT
XgJeoJX+f7RJqo9mhWD0WcSd9EEu/IbcBcwNiMrys7Ann+wnBEavcMS6KtV8Ug6ihif4ETGybs2T
abIPCNB74bf5f5vZlArYI3NskGvplnCURZHKAK+Li1oRKiBwwq6OBEl+VemRlQD42Konsx5rpgEC
2Bny8BQvGotw9oNitMmN7R6xFmwCR5NFzRdRlV++gWGprct4YRwtWynofWCFIZ01OF7EmsnFgroX
18/2ZXdXMS1ZWVLcG0KHOo8Lf6d7FvJFWKufcjvfpUafOLYmsrjfCDaCXB4tgSwJ/1NPXwuCpWN+
ZCpf0BDhOV48Ce48JhLlU4enoo2k9WBF2RQiOdopGxMVnNQHx5gWiuAKTJN9nk6y12TpJn3e0OY3
sKI4XpgtfUwmJ46Afy+P4uTwoR2vxb/BIVn+WiY+5TwD+HLRCHA/qouQyHq1AP1tpyYSnaUVSNc5
SG0dvND3lW2cx+kU4jy8EoO8Gyh8jWmyaefQ9LyDvRVWRNrI0HDxWVbhbfJtJOpAaro097IPpOx8
qXlGInEaKwoCc5O1ZWHPksF8NAj/p64SOU6c94eLzd3jYVGRLQbsD1KFPhZPv9uas6VbVbTM/u2b
PzXzTqsvMPd2t9yiM1ryhsth4MHfdNDd41qWToOwli1W7vUZYuhTo8aLljWxJAJp9Asrv3rAEouE
bopM06/UHfhemSWwXAksnCUio7CgS3jg676LZ9TFcqrhTFTec8Qol+4p45NSWov3ddI9OetOSV5x
u2c+whTRL9nCb6JAu91Zkgx5VE3+bqw8vXHlKIeayXrAGAuM50TZX3feUwTyyruGJg+hBkGb6I67
4ezjo8V59Qae0z2ikeMQwX2dCLjD6Ni2XdxyYkUk/3H2zjE7cBJfN7kLxz/ubuH4taRFma5ooUH6
uL+uTQ4BO7a5b6N+YVcLM2Vnoy0d8aRpM/x/2Rr9LO85AbbIFJfP5TH9SrUtqXb+kf8xTWCKzeUj
Uhs+k9SAm345YKK6t+p55Sfnsi/8+yCiMXV9rbfmwAi/u0Mg7ynS95wcgFh3KUpVwtuO0d0X5+gH
f2SjHmlFy5wmog0Kz5Y/TtkwxHnRi9J79vse4Y7ybW382Eo5TTLHbwnnX8/01v/zkJ+Tucc9NgTq
r7iE4tUVg9hsMAntX30JUTQLlNBCkUnJnmrnibJVw1EX5pCXAqwEAfqC/C5yPhVJWCRoMHki/u4i
aNTVUCes0dXLBnE1FqM5xqmVlQkrMblVwBlIexbxqGQCsfKkQFKItLjF08bgm77lMTFTASHkvPRy
J58vxd/hZ2F/9ze+hJjJbxsfGBF3hy2z6sR1jgkS+t8j/aZAHwYgx9/jLG9F3fMI2Ix6MFpjl3Tc
5u8pg7RwHV6CZ6TJHIwO5imscO98HlRDuvQXTR3A2GV3X6iY2GWtgc3mSrxLTKnkc/cv6Wfj16Gc
h4T92gguNsA4LFdcCDamPI+Jgdcfx44QlSmLmaACSIm6raJU1cw0W3RXCAnNqNoVV8BCA15Y2C6H
jUdb1lB4z/EqEhwYPKTsEMi0UthT2lBC8lOAAZOijLf4lsOijn1Ck7hFt7L59Qy9y5kKPoGAjtia
MHyDJmkb0M0v4d+lBWBMdtC1K3/1bQrP0ou1SPkrnyW7LBwyr7qbkZr3fZruHZACETvDYIykFy7B
9YSrAKGO/ex6M008H4tVo553SU1J05L4NxJKqRCxIndFCD9Kg1I53QPwg89Yf5x+nV9Ex/lzL5In
v22szUGwEYNAn1KqG6g2LV87rKHErcayz1cH2QuH9sXU3CkorjgF7jE4cLohVZkWZANNfc3hjMg4
1bdrarOF383oeKzXsoqbrnridFKAxwi2ASkRHwY/yY8P5pI0XxIL3sCGtS6NYlginDM3LUqAvWW9
afzVeLYI1K6j5Pp600C0BPKHT+U97cy5pVwVGYzTpwW8Zaur7idgAmBB1DfGnAu0oFcfODqZyo7o
QSB8mft9bqnsHJHM5GCfxXXOudv/GDWS31He0FS5k8bbghnSlwwVZjpBrPsm3vklGKMlcgIUJkWY
PgAM2sPejUUntb18dLR4IImW4r18XQ8ApkQeEWbl/LSwk4ptKtN3BbExLZQhiMOTrJUN5dsHFduy
dnkBfkexabULaesORVUnhzvhSJq0ETyN/nsMu0pLSg20rCH1VTql9xkbPCpdaO2CEAMB42GIG9RR
AfI6mwBji2iRI0LxvzTua6HdTflerp1Ai2yHGX2Hg3dAhI33Ba68eZVChAjAei5Ya5CDmPmNGXzM
PjThRBzD12KAFFYW/m8BitzGzlkpKrQJ7Cj9plx0xB2Edw94mCZseqt//STCLPW4s2AQlFDj/Ula
ThYka7+b8QmvIQ/HT3kZ1jDfGi2y7ZAtBn/cwNHYoE0F26K2YxVZ3A4kaZ6/fTZVa63BI5w7lkww
LL2R3K1ku6eSfmsTZHEh7qURW+WYHpMS8k21CebSYOYdeVYq7Iex3YLhhZSL1n0XDYUY0Wilyz5/
5RPZAg9yHmK/PekO6VuP7Qgm+xRg1ak+hLczAwq2VluGXlBNAe+tea2qfluMsRAQ5TbBePFpHU89
IutWE0o/2rVxJT7Z+q/R6Pp3R9ctsJdMcgvehXWOwFIL8QxD/OuPOyVs9rEzlTjjofuJiwCKliwe
Td5OlnqK7X4EfTiXn0wj6L9yI5kAa1sXMcePy5nCppHisfwj+v2jbM2HFYSpMT/5aoIl2VPD5X/C
xrcjQnoJJGEq7vidyGwohtRm6R7Z88Xo3G6KWuyaHECFxmCcfOhz7POc7a6FhNPE9tVH5j79H0F0
/zLAT6zFTeZknORyMpExidXviwfbvSwPiITyxcAKFerWL4chq/oGLqU1cPUFA9QZDUnOOgFQANzl
QkY1tCn6LKET+n8y3xsSyQ05NNaOH4zpRn7OeF96/xdxVHZkuaNK1dGrOoAHDuF5WDtqy+GHtU7W
ule6iINKT4musMAg/WQQGEDKhoAA41fuT84RzUX42RJ1LV7KRA1XX0ussCZf7v+xlWJEncEqD1BA
YExNVuJF9or8yvDRxjXmQkz3qDfXc2RkyZNNSNE+6Dl8wWiYYUmBVUXpFItNR+zZaWPI/Fq4KEGC
uNZCOFkEOGRXleLYxFihF+Ab4maPworn47Zw0iJ0MRxaaI+xcj3de0bhBoiQxhF6hfhsDuDCu3z5
7bDAjQIiYs2Yf2FhJSPFoaI5m+T05o0VuxuUL2xAWF1MyJJcuVor2sQdpm9eUBxik6mhg5Maj/wT
K4JccmXsiDXK0m8av9kK/SwapAt8FzOhbQEUUZqPGa6MVETBXEGaziNOh7NqAWb7ZPFl6H+bLd/P
fvCv6+Ijr4jd22iwj5UA0HF2oaEk/useW1MQUMdwpt8xU//UuYmISlWc1eG/BRnAwJYkROQdQUhd
AhWuEmKhw0J1nAF71FFTlMrGNVMbAVvh6K4aHE1HtaL1q9nNORvhi7/TtJeQTFsoG+Vh/GrHUjH5
+2sul+A6whz+vr8NIYVFvcQlfUNb0rzPAg916GE5xlSKiIk+bXL3n3aVhFB/nPPoYN0w98nG9Ub3
b2Kkc6sJnOvXbj4vipvIgBrFasxICbJ7O1eMd5u16R5jfxjE94fwsd3iYhxIIeErLJC9GOYf1yC4
7G6Fr8Z69Z8+L6HTd/G+qZQoHylm9PxLFSrWjdCNTlW9IHOtTS9DdeePB1NoCRxbrWy+BlgfrjV6
CP8No8JnQcpQp9eNXgHiVcarLnjB9nlmjn8LxnXLAPe7NcOoWGC1hhwUdqMfvxKWV1rDeWPCDwrC
8AbU0vBQbsdYUwJflUExGN1dhQuGH3bhuUJ2aW3QgJRAGj0a+7MFh5/qOys0/a/RGdKP6TRbyt30
y9U0QobXAgIjtrAw8kKsHUF5v6lm2fFtDCFAxbz/pZChNRUYK6OdE2NdIjb6WELtxn/Y3Yi+afcL
OTnc/pJyL24/B9tUrUKPlmII4xpDGooEClTOG7DNmekBdrKGz6ucsbJ8YUDW7S1UN431IRgR8XXu
726Q49FVgo4XJ6pBeyq+1HXd5pocKQ0HWJS6hrv4f6ANudC7i4WFnUBdD9LVZK82BFgaY3RgmuAC
WijULxlL64P6Dt9x9knB7TgF288rDHysCox0Uc5V6gut8Tqrrtw4lp/Kb0UE/heFw8LkrO1FBX7x
pbWYvg9WAAehHLXrtFVSxD0x5RG34SzcV4KEzR5Dj1Fk7yqdQdYGDCvf3I9LSaF8Rz0tHW6ntReE
qqe1+1EfkEySkt0rwd8FduvM/xErst2HrwKLxFPmoNV+47b4Ep81Jk6sbwirqvfPDw+t2wyzJnTF
gK4WeGVKYmPPJRXlSNCxLP06suzSr6MKWu4LWhgKQzENCIriEy5rC7PIgaklsLChJMIdFD6DTFDD
Uf3fycqjGPPS8TAPyoI38LUJw1EWE3hPgifqRhJiaD/yjBuOeVXkgRMnaX9d15I9VVkDmgFTfpYi
wABkmtCf+2S/al+1M++5WBo6OiqIbhylMyCi+tXQRSCCQBgDZ3RhwzFCOMJ2OXRT3kILyiLcpBmq
14AnYriTcifHZKkn7wDwq1tl4PJtQHYOsX3JOBf9vK0KcRAPjnQm/ht/OtT/4rGdTMFI3xt12uo+
Ih1CdKPj9qO3NnG58wZdvxV4T2kX6csQxnHEBJqyGIkFkHCsorRBnI5+kS0l7oRFjBdBdr9lSC5o
rqocNOphO87BsryCT6MXEXahV/hfBm4H19qAu4dKM0m/px84VQg1+30+/8Vif5SlclZQUNZwp3gs
333J4CWLyDLBXkF9mzYdDEq4bMUae0HkHmBc10833IYtKNDNZ9G4WL6688kp/lJfKJcRbTyQjqDk
l2k2y4mUaGt4CdjVg2KR/4/j45KkGdI/xgrXTEW0VV8iswnZ26XVyk0eEfEvmOHuhJqChcqf04U5
XgKKU5GZQc37XStddZjBOZUhML4oU741RTviqwpitvlUViSJd8fsvUhRRAPRxWzDMHCFtm8HvA8a
vLEjUMzmZ/xIVH5WO/fNIDNlUxg+y42rPmihQ9U4l3zVsWNbukNUtGz3jtJQi3/MQwezcIhink4L
5kxRdH+Ujmvxjy1MmpmyLm8grdOSMIWWT2DP+iIujlHvN7RrfHeeAuiTZOkEvlHmshJFndbCIoIY
hn7shcvYFTY8uSRTL9Uf/s+TV3xeF0CncgEgZ5oFqfG2VGfDNK9WrYfsz93py8sUpqVqnW0UN+37
P1vZV0UHqZF6A85Em/l8xAIxF5V0MBOYD1eYfg1HST5io7DOMXKr4YdgbFB3R5wxNui4czvkv17m
lzH+HnHd/H+PtGjtrwtBsUjTWNg+v1IYNddoLS9iJUWij3VmgQ9G+eRgNCDmjwAx2Qw45u6fC3iW
TPzE+zxnR1ZuOXg7jjut4dkKhzLYy3cmqzNviMtGDdHCDd8NopZhliZaomuvN4YIf8LQfUdJa2pt
y6NamNR6qtvmwJBYChlC06aRMTFS9CfcBrpu0DAqoVcj0Rv/4qz58DvD5kB0xYtNnVylMjOhyH51
0xZJ0NHFHC5N38QxGyIST5Q6it9oRCikdlhRAKE/lAZ6Mum/Vctomiw2AaInrFg3+W5xdbpM5C2U
7sRjuTp5TGPuQR0WPbBtngzvgTN6z1DF8wCP0oP6l2ppAbkYy/BcWEyNaoSOJIeyXHzd2RbpjumO
2c5X+FEGcCXS0DBjrFDNERDUW8B7VFAbVJRF6Z4sXCzwggYumBwbUTh42DWpAcGuL37ZzOgTweTX
LNO0+HNs/vUWahGYBPtEZJMq3M01utnP4Adrl5DFwIYCNX3X5wtRBjTimsFRoTvVxljmrPkhj8Wi
DXptlSt2DCPDMe83QUVLqdpLF/5RaTlGp3f+Esi/V9KmZ8EtFHwJxYGwjnGE40F46r4YsOosCpQ7
S25WZtkW/dWT/RLT2+D3o7ziH6TSH0PkWsQileKkfW2IlCwgKZIzv81Po5daz2yWpe/fSxItcjTN
8nZFd7N4W2QjNChd/2AfTjbUMtJ9I2c/z9vOxM3Q7icN8kW7SG7mrkm/9OxixDs4zjTqGknyJV8J
yC3j4eCUXHVbRH9YRKw4suo6IPr3oKblJ0c+5WdqlQEubeNOSwSnpb3O8UoQCskS92I7QuAgbf2e
kr0P0bdAIRUm1vUlM/EDOzy28OD1BuwcHIU9fRRtcQnc5wo3zFuHF+8O/yiU5+O6GqQ03P8PC88e
Qe4FT38Im3UmnqNhpQPDG0eugAVgS6dXM8mIO7cEY3iGXQ6fNNJlKnOBrr3Ac0owMUArkR4zVsuS
MKQ+mWZkuSpRmgTC8H6F0+fZPeJzmdqjjg8dzu7D/Ga8RJa+DrktNl56GjFvd0ORsfnnzTZYbFki
14axuxxGhTtqG5OE4SjmuQTVg7ZUsqNijCDTFrN/AXvN9ug+z0XHpStMRcFwSnyc9MxlV/a00dt+
3DSau3gv5cn5zuLp+w38EOSXvDzrQ7XNp7HOrN530mnMCXyJPni2DC84OD+Tx2UESifw46WYljoU
yjkRgr7AxOwX5GBwSPT+aJLmMoJnmEXL2DbXfEDcGijsOKOl38uySYIdwE47oRlT9833b2aOGw8G
JaNwRgFa5pItvIYILYmKzs9Mo+wBFmkutjG1yo4d6t5S3cjOI9GnquvaeSa5MgtWPlneCByoVZT8
SzmopjVDS3new1IOxSFEf16vOtLVOC+BjdxW8wBneLjh0djzExRqUDmgTLEv2Zt/d7W1FZcJ3iDi
RHWZAWuw1qYdR63mhJYi+tzN9tnN8WptqFk09MPhgD4lZV2qa2kznbEFXF4cql0fsCo4SB7PxXmg
zeHMecwxPfKuj91s5cFUIKRGsNAFladNdY6sjM6Fb2Mr7UhVCQf5tdHamDl+oMnpveAiGgnl+uSD
GUOfDPPrPqRaYfzr9K9eTX1QNUD2ke0VSDbMcgn1LHTaoeJ22pgS5AE5n6p79fkTG8fjh0N+hQRh
PnoleJsLVgDvDpn+PiSoioGZ/Zo7dkIGxC7OezK5pEvSTzz3HCab2EAK74bmnCNh7GZEs+9JuvDw
VzDbuqTWkEYB8hRyrNdL7s8vaV4upbuDlG7snxY72693GFlb1IHMDHgGz+eGPlv6bRtNLVPdfi9f
wMBaYunOET7MPq3hQ2FS9sE54aMpdEfaH2jphNOFPjej1ZFa/2t+JZc9dVwkSlMEXdv7qnqlE6tZ
X8R1ZdxMVHJFXXANYcg4xEhS76cl5buxvIEOSRUqrVz5amyRcae/6/JIGbGGee/9tlk1WS4nFwlX
eCWQLHbDiHHl9LuHJGaVrdllQU8W7c3Yfm6JhKgdpznosHfSpAW1HZnVyDv9u7OUfAFu0UWPf9eZ
DaJoQb7Nsinn+kYrciWDwwzTOv/TdfH/MRJol1Iws3IPbLfzh0RZycMyC0nmoE9lfaUhTO0kQO0W
6ez0Tw8v/gyGOxS6C4al3nUHu1C2FE9F7ViWYUAcbTJM+X9kq4EUpW7A/MBWJ8Wj9sROlgvvhzkb
IrcOqLNgyY/RhpYB5oVMoBpFUn5PtsRXGiMd3+gobmaVpIGiLkFt2D26p+JgcA2vNKXmskLoEiLn
dDH7MA55zsY8zVY+MhsyxuHWCvvKVHDmaWElKZC9zA/TkD6Fq/o/6YpbL5GDua09O/a4mFXYPzOp
Uu+ni2jqMBI3WYs++Vrw/TrOEt5ZJ/dZsV+BfCq3qHYQGRsCPvrTQfO+ViEyFtsuGBqUSBJY/zd5
YofSuIk2DzhMl1c1rL482kjGxsQMQQVpe2whzzp8Gpbl9mmv2uWKkFmJ+TWc0i3acoXNq0lCPn6N
MMOpesroMc7h0Wq1c2JBdKdXf7FCCN+rM/DvQCXAqj0E0mxPUDdLMMqJNCgGxyASGxYDxxvwBTho
o/XNtJwTsgS8o1mYdGd+VC7hCwh2TrizAKhtHfPTuGj01gLh2dp/H7q7A13sOUmhGsCMS/FqIxt+
Q3zSYHpTCbYd1Ktz1jYVEvYruH8B/DS9UQYPnrk0Sb7QSSI4IVoTzHygLrDRL1bJ4PFv97NoFl9p
pKW1DaAI2aPGH31a6vTNJU3eT7p14rWRgAA7P7tnCTMhRlPkI7Sj58drgkKYevfgjymsMgryihuD
GyIOzBwFlR8ImfyvPNASI3lcuLyCUw0D1g7CvB0XjOStmTIJ/2RiCq5qGfzqoV5rKmK5CuIiNtyc
N7oC3c8dVsRSjWwly2kFGawIYg8zuBoOXN5R6oZ5+OIIUu7H6d7J05+KHYRgJFV8CmeJgd8naJyH
d05f5cE7bXMF9dCmdYydKD64+WNMvCW0yvd9gYhXShEQ5UNPk8XTTm1+MO5+788UzD5pJzj8eugq
cc8G79aQRjn3IXkGcQFq7Fc4lB+u+/xNhO3SM5i2ETgkivyyVHTZBnmV/XKwXGwvE9mEC6U0V7lh
TtUP2LdFgcAInsQqBeZZGGbgukazHM3np4h6x1rg2lKOIS/Hp6cmGFX2M3Zm05AVDddRgO5Le0vB
eGsO3AdZxleHGFTAiENgY0v/lTBWqxR7vluWROw0ZHaR8ZkD/nHtP+kNYISUz4Dpg+egV22XnpDz
TAhzV9W2ILoSHZMikLjjoUqMFaadoaPk7peh9f/p2btC9erWNmT/SiM/xb5NpGRxDzTfKy//KDuF
KCuO/brvS+4kY08rGYb4K65VEFrBN3d4kFuOrl7kPPFV7Qw62pospKflXrxBDx980ajX0qfrbEcA
naOery3tgxfuKNUKEBuxOMxVUcLGKVd4yq8QT2/+coBTnMFRWewgSqdrcPH+XilfksMCnJcgiPah
KPN2qNqXHGGaygMo7pHnMGKchrXCJSlYWNuPAoUhgm+Qui3sknSfcUKH6b56qsuxhx41pKvO/pQ9
qyhlVBM+Tv2m7xORpoPhCzblXMUm+j+sKM3Pjroh68TBxFiGkW3r66KFudBghjt/0PqFSarT39Np
0xiqE0eIC3iMwoHpUQOAVbnNYyOcFJFVS3z1yWqrgoDR25dsgyU4MXuCesEGNNkr/zysWOMWQcB1
gFOFpAmRS5HfWXuEnRHJLmHpo69mP8zl085llCKErA5WzjsD/EPa9Cf36LF0FtbLOTC8OA1IheCv
j69LQ+KJKkiUzy9G+d6DdIwaQL14CjJDYogbW55vIJt53wtDyi78xc/15Cr6WH3q7MG31/6kUSpl
U9XDWGmrwoWFnafGokGZyMm3PZUaXx1VQ4rzFROdDyfn9lj2AlGWpUAxXuc6j5c3ciH1p/iFBXCu
kfqYN6VZW8KMxKrFQ1r5mG0wfWo3hs8rLEJN85SU6GzJve2vATygsRCOU3SFpz87BMPBTySQz4MP
y8Hx9ZMfofAViSFusWMEKxP17904q2dr9/ZnhT4QquOYWypxeBRM3ebv/tZi3ynZ8Mp3s1EwBZTP
kwbLrOLdDmzs4bpyyIljSZD14xhpM8OFNs7dzbbUmJg9eVm8d+M2g2BB4u/YNAXMfXlqSgPx8Zso
T7DVUQHqhjKWYQdR9R0pbHDqkEVIdfdeSSXa/qz0+2J4LPJ5kp0yajCzbI7Eg4/n8Evt/NimbQy6
OXorqyVSmBGqykbi6jGy3leHFtyjXDX0BU6qJ6OL4gM1Pf49OjdKv9Jo7KG067NNrlLlDkTI11nM
9P9OpHDhkPYynJN7E2CQaNlKUjpGNTCFNbYYRvr6uGtjOxImuewc+KvnsVzgLviUcP/w7Y14P+a5
SgkQUZ0fMe3eTvonDioZZvMBOPFsF6xAYvXaa5pGovBCuOhkpfqQ9cDdB1z8q8hqSmWVcsyjgVkz
Wy86Mif7/4ASkrIEFnkBvsvsgTFDlqHJCy8Bn1pmxumdK3SKXH5ACUipGOM06aiWPXv/cHJqADRz
j8YyPddWqjwsoCbnp4ua34tOvaBF5yeg9XoI0CLGin3m3vdfBhD0yVU3AzUPx8XMI8NOOeYVPXjJ
vDxU/opmsJRbNF+KUs+UhdlO2wmb7yoyG9ZmzWMBftBwowQKutPgVAiv44NeLTEQVPNsdd+sOGtS
koDxtUIEwu8QzUt8PKkjQsBmWRlDBwj9uvTQpRFVwCkPwE63jffGZdgHoZDhZX3AhuNPDsABkpai
/ye0afHyMC0B+/4TbqJRe09ATziNLCutSid8MM9wr0bP8ceyFyh5dx3r4J95MsN9dBpqFyg0NFep
pjq87TLHP8Wmln3ryIg7lghe8/AzpKrs9+1aNsz1lWomkwV51EuN5olXkkXJE8nfuFn+PVYy1p2U
89RLzRorCBjrJVhbkkJPBUSDebj7Eb5hfHU9dTFwgM0QA475xvl12G08L6USFGIE4lLwu8Zza4gr
gtMQjhA+uHLRinFJWEI02cZ5yQ+Ubcug7ZLa+O4LYKQW2l6VV1Q4y1z9ou3OPbeTEseEl4n867vd
gOAa+7VRR/udghO24Mxkv1FZZTf7bxidaUsAgMb/lvSWCIKw9wAb8Cc4cBftSzBeNiRq+po+CNct
flAwNqjKKsMfFCSRQWhEO/Fr3kPj5GPGTvAqtBupceAFHp9urDO0Kcqp2BU4hgfkejmmkdKM6C4t
262JlQIoL+LDSc71vgdp2dXBsoCJ62Qxln2PhsaYRlJCf+/Wm621FqeXtPChVy8nQZYRzhZnQCmI
J9YLu1bUQwWFrH4t/stCx9YfCenXQM2Y9wYzcjqfqJLd10IG4wRIs6sK4vA9cnueEsbXzdHizo3T
vZW1ScmgBZVnXNX7BeeWGtkEfWAWtCRw7I4i6oi+98ASp2bnosuE2jkrNAMxPpeXAaaWAfct78jM
qtc+Wzqrv8N8fBhm7ddlb5XX6QZJTyaWJidjfw/GeeOIzsa+DKVaKrUdPwfaFrvHYTzUoS8f/GSH
nF0E/ato3ZFc7LyYenWRWwN1lUxd/HqaQFkLbKdUU90mqqAjmSM8yh8y7WXG6d41RFDjCk4jhxny
i3zeG7kf2ZVOQHB0m+QtdB36hno7OcmtSluIdv2IdqyThx2OjAjziiS8ZikOPrdxW5gP7YYm0tiv
OZgQm43SW9SbDoIqIeCY2F1mrkQDbt6vM+no7pFQ/bgVON4FEPE86Q2AkV3BVikb/asAep+7v/3Q
VxqPxloGYIW/OmtJh6yh1O9iOyGPGKL+u1mMal7iGWel/C82X19FPO8IjPXeXzpYXAc9urp53tQs
Fg6MBIpzfUQXqPQQVF+O1hsw40dkPF8Zg8ketDtX9XEzHjGLqe6fVsilJGUdr1EY4N/Qo8Zy6CCj
pISheCiCUuNCvKeaOcbFgGt81pupCGtlyjxw9pgC2pkTkK1t2R7s7qP9V/yBE/y8IS3f3jt/G3/r
fB+cRl99De+WEPoVfNVQdRlbT9A4w20ronLrwaMyuJfId6uu5FyE5FcMIHjSAI4i4DVvwcRYV9Ei
2fqxWEAgkMl7IhiqquKdxp9fBmkQxjpWzQQpGkAgXuhm+dzL4qhSCIu1m+vIcI+kJ81OcR+OOk11
xSsAdbAOEUUT9na2BazBThjbdXH0WlnNP8hvK0sEr+gJxzhPsJmFGIRlxF6lT7Q2sij0NrxuF0Dv
ma1HIciLTIR7nfPb+1Tqnv3BtInrW1333fll8n9RMIKwmsEEzxP99vKYtTnfvvbaNTf1B6Wwt23h
0hSNWV8nF5QXdVK/F9+MTobr1zyFA6R2qskeJLgVEwDUSE34Y6/HGU6nar8LIlc79WObuwRe6Nkj
vEHslOZVzmKzq2StOjofFWdBydXD2/QeijL8MUJsOA3Bd1FAQnRIU4Ncx9LeclP+mqT0uEpCvo7F
kBwHOXDWTM2uwSeKQo/cLqTFEZDIqQXoaL6wpwIBbAgWXb5W2G6KGIHNEYBqrRFh+RYN5PWrlQy2
13LLHGIUcHYZyWY79dSW905t1lcM4pd3RaJK6VjpecIm8MOnVm5CM6xvvx1tLa6+bS7oNEZtcbWO
eWPaKOvyanOyiTLazfSNtD9IkJ5Wsy3wzZ1whVwwXYKrgKY6dRMSo/MHVwSMsK95i1DR/1Lbtqq5
qiXrMiPjpXdcdIHsPxsx6zwnJAfL1HfnqKLVtnbiK0BAtuz6thsZVmJHCI/zc/h8oC+6jZWFGPFm
OFRUxEHBZ7Uo2spVOVWGRSjexWCThp/Jr0Cgos3Jf3izZHPb/P1tUwrv6NzDm321ZM4qJ97o1wIH
P/obrO/X43IKExeoN7X5Quk7rc7HzGru4MDrZqp3gU+lu++N3e4vk4tAjf3AsHTMkArIW3KRadT+
PLCk14HCK5zSAJytUnyEDwu+eKsReRHkMwH0KVjDKVm9cv4uZKSE7J7anKdWZlOV94muIULC8gZH
kjyOb3/Es81GBoGUBCPmZMOREylzOEaUIa44g0wooUdX9Moos57lc2tfSfBaBmLfVb56sr2g0Iwk
iXUwmkrednUR3hQ0a2FRUDIEnVW+2yIRmmeewJCKDsI5CiNyInSsM6s/9oHIgyoCSkJ+CFgGh5Ar
mkEw5jkez8b4O4kVEmpq/Xrv1ThEgq2a7OCmI4x9xNF8CYyutSOZsx9Hyj9PbKcenQ6y0nicjBlV
+xp7yv+PLUzHZ2hRJ5hdOr/M96T9ZaTr/1+kk35tf60SZ9SwyDKM+WarUB1TvSADWq37nBhcpylv
T5mBa84ioe+w6+eTAa7k3csZEu5yLqGrW5Z6+VweQay6KFZQTpQgLU195XU4QWZkZNiOEr0HSsgJ
yFKDaAHH5m12aLkSVfIozf1tfiD/afsFoL1tgl3nAz4ANDYeXOljwN4slwjeuYvn086LtRXLKQQP
JiJa/1HedcAwc8dFEe06pZl4EOXPrmMOB4YKsGId1Oy8kGVRtu98FyNtTkKRSDmN0B/eHV1eZ5Jj
FajgaAOE0MfqwSjiwyVQKwHYIl1urkMrz1att4smc8nbfJjfI0VOrYdejiXs3eSW29tnDwSGHgkR
Xl4Tm+pZ8rVOX/aOBDUq/nhDCsDwUgo+94tPd3l5svsckkkqIdjsPVSO8eWAEtO5zeQKblvszlld
CLwzAGkkUQMvsuKJC7w1tm76kQ2ot7jilLwEK3R4MOLjQXZd7KyuHUQ9TKGbAUHuDkA7tjrsSgjd
GgvqcQc4aNq5taLjUXpsjoNT3WU3GdHlktKimSVJtPkqgi53rJX0rxtjtuDmEEmwbED0xc2jc/Ir
9LTPDauAyDlhNt2793Ro2vb4YEbwUlSktOAPMOWv0H9DVzLLPyPBoIvw4yZ8pSau/YKuGKj5zPlC
uIVWmGqLy81NtMVOklTVvuyulAKQckgJnhXodKmHyGRIbCHnHmYbsJA+sXs8CgyAe4J7jfb214kq
XYPUWoU+EiYu7nJyqzhY7yyXPVjbUbl8iAD0JaWLr2UzhdzYDGyHOAEFxLAvs3pH19OG2fujGH5R
fLrNMRroO2P9xTRS+4fSWBuEHb/a6VxJ41dl+K7/yVjQ6YsDMsVA/zLT42gKvf8p8wxd0Qx30kJ0
GFrd0dECWIr4sUOO9nteuCGteiU8t9sUMYP//VTXt1t3WVVad4VnYqHN8zbQ64G7bXNZfEC6GZQQ
FVM5UKB9+ns2wOyBnrJt0XfK7C89WsmPRq1G/UCs1+/qU28Pne+zo/1ILwgbc4xlx8SnQixaTu6o
hT53GAqc/kQLjSpmhGrEtk5WB01uaRd9DdVOOZA8s0pUCDpPC1bYZHGYZdrrLN6GckFmcCokTjuW
ex/riytVQLrQjGGAHAbNN89w8s3W/RIiGGtrzImxPaGO8bjknj/u3M1DMyHgXsQd130nkFCvagyw
RTbIZiQGIeu/si2ld7uYq/RMXnVoBaDsgdj690LvOzt5ddiJvg3qUd1CFsvs8ReO3DoOeuU9dZ5K
cN9MEZXhuOtZOvGKRH3b47xpPZHHKvqjGPtbr78q4/SyNdWtesF73+W+5oXhu+Ugf6V7J5iVLbMY
wXqYWlV0Z27sZpOGZ7lc6oSCmbw2sVHNRrumRVVMGZ12N0tIw18eZoJPdDl+xMHuuxwgaI8fztDB
FMXzH72UkeseU+ENVaQ5vQWVT6QCbCAGRbRUt4fySVVYKfIecy/aRD20hzR8ldPvoD0sujPEhPn9
YsGWTSb6J7jnPvu8hqgG8v4XGapvqI0MJbcKr2p5ExBPrlJgkyRCvNsI6CJ2CsPndRsDA80bFZCT
CHsckZnwb4jwVzhzVK7ZWQtakgRvR2U6P2djyPPnAqT04Nojnld1IYtVJIwIaBTN52R/7DhY3Oa8
/JP4NsN6JVSlQtK8J5eWBfqO6+MMBLKH4oqOiecciK79reIXmwCW+Cko3jfxJOdQcjrTNBp1kRwk
n2objteeoz63upeZ8arzNSPFMGLdm/HQe1/l2tS5nrQQeYzpbtfv3mX46/7jDkwCfZJvHy9t/TxW
Su8vfmu06FGg7KeFCrUgrdeVx298F8QaFa68QoEHjN+dCaRdVML8/OEC+CnvB5oRNjiqEWm+TBKZ
251bzNqm0oQmhYW/AVn7hho2EsfywiV1Wsz1mCGuWNjB7YHU4rc9Vafz0MSWfg3tvKJwz+j6GXgv
o5MfwFfgx9sHUUNxkrDm5DGPcSomb9TF87+7lzxOckpotUMliytJShZIZzOEmgAI8Pwel7PR8mUa
TI5i6FtYk5mzywAFU/8+NlOYzItFK3TR5CzS6D191cU1j/jHZFRjHXuoLQ9Z46s+FKlZs442uoed
I7tlS6NmJkZ5AS9mkEV6atxnB0aTFrGNOA7NFEjBYwbQ+/yYd1AFffw1dpdOwjZqYCtHsjrMGADJ
FDb9xvP9P5WHzfDzomQUulkCSmFIR6DwTG+tlZIzYV5AqtKVLXVH2e9ijkBCRarqVSGO2WDksRM3
uaZ2ZGeCRGtOcrbZ9WN3gPLd7PVyb8nW3GSXtZgQY+zEmJMlsdnBbDzNea1DvlMu7uDbM57ZWd4a
N1yycix+3Q6CVTmQSN3sFfmwwExdo/tRXiYYuL8kXERynMzMTXI+309lXaENHhjPwh5VRytcty8H
p1vCyYT5BqdKufFtO18E1w9vGmZYR2h1w9+I+Q5x9BOQNnBXuXKCnau/axEZyby8XSgwcKyivQ6Z
bx9gpHV2jp03+yvCApRPznVhth4aJhKgXTKCcK+YaG+F1E1D87FwD44C1NCgJLBKRQw7+lwdNu3i
Ec1d5nqjrXOxPJ+krgZR4E6mkxu+d9jttsbCrYeu4NdVwGLguJK9B0PWizBep1amy/4Y/aWk/mN9
VMZ7LHLEJpmyAp35gzPdVH1AlNEcg808S//J+mQx9YRQ5oHd1wG/Hu09aiAK5xfDiqw1p6Grq58H
9ycr5ZS9I1wRj0dWpfbI/QhnKUHOs/ClgQ62NBV5Yn/3m+mziJg27Wnm/LDJzUchGDfX+bVzFJrU
CX6bmJFu6q3zSS1dFOIwsOuo7N2nb6rTvVpkxSjHxXSMIYYPiGlP7vHeA3JOrD+1LiK1v+sFTFiS
fPPXpdvJWsG9n+1wNTqoAH5bvmf9Mv4prYDPFAdw18LJCSaaUZ7pxTPHxzB+ZbreQIUg5+I/W+qf
hZOM740zhBQ/aqThT67vpKHu6vtvhkTNAgGjViYljvBkUmZoZON7i+yilDcXpVLdMzRGNqO73Ux+
6iqWpL3XsyMrqpti6UXIerLxRvVVTyI67WdyF6rywSyG5MR5jS5bHprQhTQ7SEn9GfGHx8/smBx9
GSjPx939ysH2VAd0G0yvGBjM5MA7ECzKrtatWpRbpqFQLG4bIRrrPMtO31WtsRSkcKRRps2AcxEW
ZmK4mGJ7JsB0Lw+h5GLD6vYdr2dOH9t9CFgoQvVYj8aa5to0R2bn8+OuK/C3ldm4DgQiLZGlT9De
AoRfggHk0D54YpDQ1QQrnwj+8H5h1RulygzF0wfkM/oolf/46t79UT4emwb1yyKu4g33OAn1zcLh
eALCwhnhXyFoY9dxxpLSBBH6fEv4wwV+i0OpWFra3PjZLO7JuXGYGE8Ie1NMIK/65qUbEKvJjNUG
qfw3MWbPvRyhVeQxcYvUFtQ0MDWTwsNhAQkdHbctwQVf6fm6gXu8YBWaAoEm/Khiu8mNFeXCDtwR
DDUmRZ4TEtKIoD9MzGs3aSKzBnvZIx+p3j2BI75Czbs8pA38tjUS5Liw0zc61uvTTzc0sqi3DgwG
qWDkO49Jwf/JBrcxnkN1GaGqrXbetgQTuvUBjc6Wn+xk5SrO24zMHm3gHBybYnfIFRcYaYhQzWh5
bHnXxHyHecZl/F8aprzKnVptuXK16iXzX2q2ZV0fvI7lmToA+hBmDR/16cOKLzqmW89hNNNsOB8S
yynez9ygZYHOo2C5FIJ/UPIhdXgTE8DwFIQP6EpPl/g9gAkzZirGxacqP8vbpLyliSb0RVQWdd0f
CHB+K0w2mIwUa6aoRTUbOHJR5dQ7+hclQPKrYXRoO6XOxvM3x7pa1/vmCUIcmi3aiNv9UquXEj0o
Tn/XXQ3uhjO7pVUE78OhC5/F7T7/kWvMBbgy2tYtURR5GJWaUYfl4SPJ8kaV2t4hH43GIs3KnhtI
kzVIIym2F/UmHpTiX6Z7wgR2cSqCjYNQWNNNJYjgxCux/QdFk0xTE/f7HUZKmi8RQekaPH+Y0a89
38m6PS2IeBo3DeOT6EhUR+d6txFzGyPmXdDoYQSKKiSjz25QaUdFEs6MU7nlZoQnjK5hbNcqswWy
JYV9ZRxpPF0WLYVjcp8G3/OyqlOC3cTcKL+tcJQAi0WByg6nVcihr1DpsNqaYdKlP1u8ZKc87YbY
uz5quZ2v+odSfLZzewsJo1J0xqfLQsgoTvuxO0Z2yXiLz+mHDgl6NXOSgjdt9i5pphuN+o+/QH1u
tuEkLxzBx3FTUD/CABZesuVFqQGh695AF4Kk0yJyq41SZBsU3V1nw8EsA08ZmeXkwI7EWyZhfDTC
+js+AVHc/BZuL36ER4p1I0DTF8l81x8d5fYpuQ7x5I8xLpnO+JsOvO9f/qQvELUPbYUwaAxp+38d
A7Mi1/Ihma3Ar8J+t05Bclc5fFo45uw9hCmVzlP6wcl+jzRO48ha7UDVmnpK6Up1ZLx/eNXElQBD
9AU45i0g6RKKYDJ7MnuHIdVrUMd2TkgPGSknQkSS9e3bFNa9Mi9ml8uwfLaBlEKhS0TSHJIifBtY
Viry12Wx3EZ7iVIPjZ3iZ/RmHgnfoNJpD/YsEJNbyKFJTmvYLzcayxMc8MNAkK4E3Kvu9afmAXiZ
bpyYzI7ivvqJNoFO5Kl3kkCSLe2aA+JG7hVgmpBGjgcSmXNPlgAWuhYXosX+aPWQLNn/UI46q7hn
ZrluGohqN0yfCDAPL/sWjzo5f5QZ9zUSdAKlCRZhE0cfUB8x3IZ4Zud28v7TmGBe9RpV82y2WbZe
1xF3KEFObqKoMVoLurhiES2pVUZ8+vpXHgMaQjZU4dJddBCFXwFHT4ExUgnNC4E3q05ciuvudiR0
2Mj+LMmPYTpUBG9+TLSSfDxOdbxCXqkRIuRkSSnSy2FtEBGjjPBz+QLfO1yOzDpX6FdP1GLSjCii
C1Hwgoqb4CAyp6HyyOUyBJI9AxKP4SsqaD/uFhS6irnJK3iQnFS9dtII+Az5i6SaFUaQCajmRJAy
f9JrTJpyiE0wLZHfD+aVqm9LTpgoGPOJKC69LAHgyhA4bnndsJ4qTpPVJWbWMLqDaLVsHQthgcpT
aW01HNJnSkjP9kZS1QDwp0gmYZvbvgA9BAZCy/tmBrHoRr/ljPupD70KjMGjiCC2t8K71Dh/IFHK
0TRQXFQomyg8/l9AeP9sxtUX9FGmo3C6ij8IDqY7i2ubEa5EGHYtktSgYpBUt9PDb4pJ7ORBnlvt
g1Py3MK6yzGuOuC4oBPSXmOb5uJrHsN7wUZ0iP8Sv0AKTpBTaxzOfByzGIcDtnwDgENbqZVX4/x5
9jcxDLrJ5Wej1YImhdpqTXK53B147F12IFN3WTEGlM8+sOlOyk4PV8W8dTU+HXf+X0AncH6SjCQk
w/nzDiGjUPZZ1zRIEEnTP7l2HmTnku0g26pV9TMaBVSY0+sfAAKuGALmfDJiETWRUPpXSfh45BDf
RpCevJLmomebG7fvzV+NcSUFVl1vcjwzPUShRsIkcVGgEsRAJU40K9r52pblrUAolbPIcYZ9odEf
fTR6UYFBhizldSMaojzNQ6KxmYLkyCiFfFlrvse6n+Nea0ma6G7DRlC3pbEyhs+f7tA7RmB7wzAQ
QDF9gTStLoCwxumPjeYwgZZ8fnV6Hqtt/PGmV1WOQXNFnxKPfhbP1nbGOhQ7ILJLF5J5ZCPqRi9/
ISrYJZx/C8ceJ/K0mxe5yYTi7QYzcDmb7rRKlbIgcEkHzPoRsew2oeOw8MOdnB1C9eK1GAQ3+bQi
nqx0WgCUzeMUtMmPUgA7m6JqCRHsjQBJ2jfdsX7eT4SOdbEFQ4bk6RDZ7LbwkZPT8adQQEUV5u3R
IpWQCV2E0NLn3oXKVYU2w8SvuztdT8lsFp72zj8Wc1MTtJZuHzpWt+sCPB4+ailaj3nZoxXJML5q
W6YrdkbG//CGeC5TgZJ6+OjqiU77lzk50b8CTABd4IdvKVwPFVNBp00O5RCbmr8gzSHngXA2toRz
SzGyX0gReWsuF5KGzFnc318p34dZ50wjEkbMed032Sf4c4awJpUPF98tsxqqVkVtSw3NJbBKvjP7
8mue5POGhnbk+hvtamzu1FvhI3uPTGSI+KPbAEztKu5Gfa9wDUQm7tr9gg3w/lnMp3S7f3ooGFB0
3CmAyu8Lt3c1ok7qJE8B1tR7thINl3eZDCUhFVWPLQWlqCIzn+8Rxh0tQcIHlu6FlF8oAq1Uirkt
x8vnwK5G7Dffk2nYPyW1WAhkxRn0vPRJK+vPgUWyie1IMkvlzA291IkFWDz5w3iKRSoOJntR7G1P
Npl0a89/3PeUTKAKGwxX91cczq0WlCuEEJ2mTYuHdtAY7gwHjYbQ+vnGa7HuFshDygb0//ykwGas
Kbo5Mo70jSelwvGE8CHc3OYuC813WUsfEXlcwadsI8BKEvIqyUGCP47jrvnbaPCAj36fLoeD5Eh/
DXaPu+ucm1TGxy0bp9HJmaBSCd5t9YNd3+KPxvXir/wEsKWRaVDMttTmAbKdFfo4rBhpkAtuBfKL
FxaGLjnpw4dj4s/2zf/Uk4eZ8lWXtPirGIixoeAA1EA1tgYgTJsCrIsKTDdt8sZKmmaqiAe1GB1M
bbV/B8nk5HXiHPTTJ/f+4bbypV10K3OsZ5cdahk1zI68CGaFweznigOt7NME6GVEcaGXQlxVaJAx
5D5/SVwzP9LOoqlRFTVH4HXvuzmZ58CKFa1EmVA0xFjRLJ+X08Rtq1P6aQtNKiR16rtDpsG8zkbG
62apZmYxS9J7sa6mmKF2ZlyhgvULFHD5eaSzoh2EhwfRb7bMi/lF6fxVS9UwxuqAxOMNKFcyg19I
lEx5Dkvk3K1Nes/ThnMSTQLUdD+aduftlDyg/ggkRWhG1LsqvuLl/8th/ws7x5LtDN1X/XL2M+YC
IwreXkY3VyA4tyxICo6ahNEQtmee0eV7si79K3hUMCvJJWMZB9ErA4uSrAoEFX9PxmeFLRSg4gM0
/gIEXcNqIKFiVlWCqCXcimUhDkvcpal0Xfe4cFWvfwcOBSPCrlknFCDuW6Wl47VMbjmn4/wtio2n
0Wb3gCKNDtEF5tXBhRAxXJT9UEG7Wav4KSpyGh5bySvWeNK8TSgB6YVPoXB4JAyLbZzXl5lkIzy3
uTGFDXWCl5piA5DKKXNMdrA1aykF3w9LS1sUN6z6K60lDUY0P5Q1xFzgwehQlTVxfg3DYeD1JRwL
gbyrmVVPCR4LshZW3n4qjdiSUMh6kF/DCxArpFLTr+Qo4ls+FPYJKzU4doeWiHWJPsoxPHktzndc
sefFnZJTsQQqRzXA9T39c28nwirKM6HlgCFRwR2B5ApCQAlR6ZBrUB75ikqq28wKDsmwHOSWPMjZ
EfdmIU6VQL48k34YevfuOOSWA9ihchLMsDvf0tIS5U57ODemLZCuh3xVQ2mKmEpMm+Anhyw+FDLs
JH7NiJHrH4bCVdX0JVhCmQ1cmpYmPUI/deXXXPrRS0ESDR4NVtY4fZIeqmBWnIJK7KPTPl58V54D
I0mq4xLYfR1gg89/5eqSi76x7slogZw20CeA4Wq5baSbbV0n128FuqP2SICzKBKuG6dMhNx5c0Tt
LIb0nLUchiPx3kWL5yBVyWvyzHX4WdBdOwovvucxv9eXo9bxX/7Dc3b9/1gr1UEEu0j7PHGiX9RE
JnBjnPEY5x/ZEQdVFNPMl+L1LMat5KQBKRJJg8q7YEiG4EiBTWf2v11+9kbLMKkcq7mqSXRpYK7M
sP36e+v7Ut3/za6Vx4Z/leJOHzyvKdcPrpTs4xx23K/wiOeAS5e8kTLu5yJc2LEIW9ppLSiODwhM
r/odYW9bCjzqUNnPiAKv4z1UkcaoGvz0rJS5Go2LEX6l5ije9WVzjSkJXFBsbYR+cGZm5XQ0EZbA
dFowSJqqUVogGFRgV25vmdyVI3Oom9n8BTD4GXYXWR0YJkrPFSCbt32FZLtwEDASOaImJXlzC3OL
cwdLwWeaYOHynkv1Y4xjaVxjzxUG7y/SJUQPxHUuCGJ+OzWSt1gkGWhPdyUxKGHNj4+Nd6Onzr5z
hpRxy3oRL+oc4JTeIdOVbEFNGmgMp8cKL3B8munOjKgG4bA7/iy6Ay84FJdkOuYTvANDyyd1UQIy
IwqIoWdr98gimdmDeZPb5eiJOha5YQ1dFMN3oLAnAlGd2HC8AvoaLlBJXbCQYNLmn1rbrOF0n6OT
JYUPgRqv7wMJkceVzsAtwEWoeVJEE2MLgDitM2hk1Q0Hbpaf2paB5my4NXhGV78rPkwJfTn7fXWl
8kZCxvmFFRt8DNy+5gdH5fWZDvRco/SV0lsmgoaBdRTh81tQoub6RNSabvHD3R6RMXkSnVYtIlIJ
mVGhLG7w9MLPGGACV/142PV98qQSnvzmv1J1L7BpNXBN0UKVLHhveGEq1hZwd/ztqm1u5oqf8Tkp
q2UwODCOkwzxNjFE+fQPo8CR++eB1QVIGZ3Uh9OELu5zgBWlsunmrADi4W4co3mJXGkIdeejd0KY
ViVb3DaQjuo1jz+buWPVBC62Dx/iuvtOty2yB5kd2+nTUSzqL2E52TVoQRUsbo0Nh64nL+i69Tx9
1ORUAGJSHdd+GoKqL9IgFxYHZfM0HNROGaGUrCbfS6/8FZXLYzWh+TNM2q/65VRZ67KnrgyV021G
9/BoesMNSGFskeFezjk6Hxi/79lruBxodFTzI8IBomymapU/9VzVVYTpcEjE5wRL00z0GhCx+a2A
m2mrtbSQNHv9j1gdXZC6LzT8ur2StGIyTvKQbBKIgVFqJNpI6/zkNOb/cJXTyZiKYGV9SeKX/Atf
rahhowuqA5VpePDfypRvDB9eTCTUkOcUx2PLDh2ZUI8TERAxDNt65q+Sg5HXQ4rODiaW00h2CAZE
eXQnNdzMXTnsO3pXKjbM9H6XYvhYnGvpuxLSqasZwZ+Cqaef+tRQp5234H9EgwW8XGrp0A2UtKzQ
vjH50ScXIZNev92MuqY4jclLKnTp+Txx+khYoyQu2rPWhAR+U5EbIVuGAtctRCiAGUNdmbc89OyL
+DImTu2Rl5hTtXLTA8KAKQ8Um8MWUd0BFJrLuDwQAh/PmPi91fsxFcyn8Riv6BL11FqSCSI8tRTu
jTpaXjHhd2RCJD1sOowt
`protect end_protected
