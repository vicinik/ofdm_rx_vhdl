��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��Euc01֜�eֹ�t�|�(���.�W��:R~m��`��E[8�����<g���v�i�I��{��
����ߟY�Oh�Xv(��M�Ձ�S)-&͵
�N�2'oQ�{�|#\"u��Gՠ���.#�6���k�)�6�Ŧ����W !|=�͛֓}6,�{�2�-����Xl�J�M$����90�㣘��4B �4&�����=�����ǁ?�J�@oZ�&'S�&�[C��j�o~�8�iN�*1@M�ū��hP��>S�n��Cr��V:���fJч��W���%v����:`���$���C�I��զr��6�}���GU��щn���k������ǥA�A�<��)�EW����a��aG`j��޷��ե��o������������c��/�3�x�	�̮�[E��#`��ȱ!�t-���7�vQ�X(�V*��=<���񮃓#E߿����c�y��<	�N;*���D���5�v`+N��U+O��o^�pV�L� ����;�7���=L�V�S������ҝ�V�E�e^\v�f[���";$��n�<�w#G��xA�)�Dй���~�m|`�G�-�(ݣ�!}q��aL�BP��9Z	�=t�WG�L#���$?�mqFg���<z�>	�E���]3੣�*q.�Tr_�%�9s�/"�I���|1�6g�����B-}@� �",�Ӧ��*��%��	Q���>�+6��}��N�.m���7
`� �� ;j��YP-��ZҟVƄ���ë
��1�t��#9o՟z�YbB�݉�qc��h����(r����P�\���X�}�����FF�9�l��c�6��,���gkԓI�cUe �׼)�M!F��H�"��_kc��҇T��J�7�1��T�flb�w}Ҏj='�Tc�髇�֨�������[0�(<���e��"�j�s�~B��i�<�k侫̨܃l��u#\�O���$E�{�鮈�������i~I垜-P&p�k��g�h?�� 2$zKёL��R"i�5T�	��*P$��]=m��ַe9�18`չ��%ǻ]t��{ԝ�	���Z���r�&i�|�	�c�W� �%]��	�?�8#W���9�W�\|�Qzv<WZ�m�����r�!�b��7�'��ы�ӯ�������{�(0���1g)��闒-��\d�@��F��ɶq���U���<qgz�l�R�����J�({���������BuI�-�W���I w� �9�na�#��"�ozF\n�cl4�94nej(��mI�n��(��.s��c� �*�ҏ��_\�k����ekoݟF�4�x�znh�Q_8���#%�p�LZG{�1�0�K�r���m��3������PV��O��Y�
��n��yVs��"���0�m]�	l��~$��u�+�]�ra�Q�Q1�+� �n~5��<,�M���
EҘF�dG��
����|�>�܈�Z�[�6Ј]�XP�њ6�HRU�+�X��K�6:�@����9Oa�FI��G���c���JJ���ZP3tF��*��~i,�#�wbW����o-�+��H*�P�1�����?c6���n��� u��������\)�˜��S���>��2�	�I�syL(:�s�/��� �A嗺v������{3J��b�S��:�o;e�[����O�d�~ J�l�]�=B��B���rB#O�������]�q���'��$%I�b*O���c85m83[d��2�a�d���1]߀N�L�4X���Y�n��}d=���Gr��!b�������h���D���io��E'��^O��/
; I��&(�1}�2r9ڨ陟ǘ�_���y�]�����U���d/����L.�X�6�I��#�3���2ղ�`@���!T��ЧX$�Ibs�����=٢�ʼ��Zc6�ýw�fy�c�D^n���iȪ1�Y��CM��Mj�?C���ʾj���f�����9�Ƞ*�y�D�$5�b�Ѷ8���s��(�.�����3.}e���ʦ�a��Z�3mg�^Ys�).������,�t=?٣�xJ��<������6��%S>\w��SR����_K��Aq�k�܄��Mp��A�~Q��e���a*���F+C��_ 4Bv�}1�Eq�u-���*���3T[���dl�ns���*:�� &D7|N�a�ag�0:���!�K���ڥܶ�͊$4��61��ݷ� ^ &�5wPK�@��ŝO���HC�Ws���~QJfEO�����(I31 ���M(ƈE�ڼ�4�E�3�׳z�B�Y8vâ�����b7�c�2�B����E����,>��vU���g��L����m s��=��A��lb��cΒK��!�^����1���Nyc'p�^�&�xd�9W7/�%��b�8�>�|��ؼc�Įg�g7��u����}��|�0/r¬��9�%M�k
��ϻKh�;gf��Z�$뤊��qx��YQ%��We9Ȯ/*t�����ך{u�B|q�6��d��*x�s��@O�}A�
�C$YK��O"i�W5��Qp5=��Q�$Ol\�A����w�`�y*3�'�C�S W n�.T�0_���|tѐ���J�u�]E*�9K7,&������^�왕��#���,/Gg�Nu�^9Nx�qZNngjI�+�m�"5kti� �ߒ����M���Ў�y�.v���y�>���?�\y�KxHv!�2F��WSA����_p���Ș�r⼎DV�2��1�4o_�ݍ�-'�u�2�u=<����$��pŎ�t4N��+>���9��0om�DI�c��J���3!+�9����ki 2�n�|�E��-�M���Ei�ʡH�G�G�����������X�m���t�,\�e���$�"�G{���j:J��<�|������`���p{S��	?����$-g!�O�����Y�l�ӥ�KA��V�%#���s�kY�C��2�U������S�a�i�Hg���'�H�9�՛X������!r�BY��bG[*[1��͛�[�,8vL��LMf��I?d��[�q�Y8Bw)�^�`_��ĘN��
��ۢ"�{���������h�ر�}Rv5ۀ���^/�v��){� �u	�U�k��UH;Ej*�t���Ue�Bȵ-�U] jU1����.g�S��%�? Je�3��X�F���R�b� �I��o4�V�<R�9/�iq�{�y[�@\�#	�\� 9¦ �'}0�a�f��~��*E�!��YE���Ȁ���|e�
hm��l���Mk>٤^܇1��E��a��k4�h�oS�����t[�d����ᗜ	�yT������3����y����l
��*�k,ɨ�/�mCu4. ����(�YӁ�;�E��סe{>�Ѫ1"(��,sIQ����\�Ǖ�ώ�7��@{�ʅ܎OJ�k� ���z,*��Dn��r��	�����`��V	Ǧf@���g��KJ�,��*����.k���`-BrL�&����w%Ƥ�Y�"EϠd�(8�7'�DR�Ɗ'Xk$��x���'|a�@t_x����@�j&#G�X=�]8_�D�%�������k9XFOΜ^�����9np��5o�W�I"����� �����3"�L�s�.����]{ot�x��fD��wr��jLN�$�[��z{�/b�ު<��ذԕ�9w�e|a�H5�L�>�+!P�V	I�}�QRiU;n��x�"S<7�MOj���5ﶕj�����e�(��H�L��o-b��~64oO�ǆn8^�y3�	�k�����>}�W�Z�~(�pRo�'�&Z�tl9���e0�/���7&���4s�1�_:/Q`e�_�����H���¿�7kO��|��B	K/�;��nP�f��HO*D��Bp=a|�FXS #Q����l{0��ع�{�a�'���hzCw�'�b9]�@����@ ��7�<g�%h�"k�p��AEHk�-
�wJ��7⹋W��<hK��⽼���P�@,���D�`ǟY���	UFe'���x⏞��&�#�l�#ˡz��-=�U�8��f�`d0׭�6|h�W ��Mn)(��[�ˑ�噘<M�O�|6n|�����H��E�5���kG�����^@J��0Ak�f��j��HO�}P$������T����/�|�{�O�|��Rw�KY�܁!�QD7�H��Xh�O���s��g�Y0Z}��]��5ur���8EY_WD&�J�à�/Ej�[��C�*e����]�y<�3A�t�{4��M��d�� Y���Y.o����ާ)2��^�0�:�k���(��FI#�	a�*�='%ڌ$���*��Ѱ�u�4|������������Q?-���3fU�AE�Z���"m$��P�r�S�w�T��ց��ެ�V�*t��#<�`6F�$0�rf������maכib�ku���m�5>Rٱ�����fna�^~R߸]g�T��KA?�SU�[�^� ��x�hX^eo�����<,�^�}Y����O�,iۂ7>�p7�i�p��P�����b=?�+˔�����_=�g��O=i���$�<����[���n����=����+�wϮ�x�|��c����R��2o����~=��^hf9�`����s�ɡ[�������e^v#4��䮥�����H��K8^
��p�w��[�"[~����l8�Y���K�oD�X�M���N��ij��'�&/�k�5Cp�hC��j�������6�;���e n+%	,Դ5(��DN�\�Y9]�Z�U!ʰ^��KcXc���x���a�W�)�d���K�g�P,Ŕ����@fہT�t��2f��P-�y�Ʊ��X\b+�0{�h�hͪ���y�ї��gG�2��n���LA
�V�u�j�	�w"q�_K��L���� Š�7�R]fq�/_)l:D�$X�c����5��]e 8��r}#���g[r��GD!e�:�aO>������)��iyC�t�ǽ��ܮ\�8!�/f^�����҅G
[U�=�E��(N�t��ig|�`�Q=��Iк��� ���=3�H�r�c�3QV�"���ʋ�=�鹆34��Ǹd��5b�2�9ǛaY�`�W��;��v%=�����pZvU�>�kЛ������=JRk��U�~ҝ���3�[�|�E�_��#�� `����CQ�naI2�Y$Ǉ{08�'G ��8g[?CR�Of
&�3'�_������n���@���EZ�y�,��(1]���f���a�z����[��4 T� �Ep�u�񉉾Gĝ��;b记p`ُ�5;� 5��	�Oi��m#��?iG&���^Rq$(H*��P�=@�XG]�
��}�u�Q^�)�!X}7��y�$vH��`��y�Æڳ��YѰs�}�
��}������/�J�_�+�N_�#˪��w�L��A����ZDy=]����~4.�`=�����g����?q�.�h�0Q�,L��w�`��O~eKiAb��x˿	QX&�HI�f[�����gJ���?�Z+�����bA˃�]�I)]l�p���9��t�ɭ5�b�����j��L���_�H�m{A�V����w�)�]�$�0T4�QZ+�ۅv�=�Fͺ�B�������	:b���<���y��9�\,U�nifk��R3��q#@�����b;�ؗ���e�L������5m:O�*�U�li����tv��ѵ@d�7�V$�$Ƃ�!��q�a��ϐ�x�G����Dԝ�����Y��Tʎ��H� \�oh���DF[/5�`&K��X�&{����p���c�FT�:	�,_�dAl�O�y� %�(e5\m P�T����.U���"另mĐF���l�%��-v��2�?qgKt=B��d��R�h�P�gl�)C���E� {�Fdgx�t,�mC��G*O5����Q\:dB@H����_��Mጅ�aΆWM�vI/+����߮g���e��$���5������%���h����9� ��ɑ������k���V�rk�p3	�$Mb�}s�O��+����ey`����&��4oJՉ��~��m��@����Q�RK�m@W<S��R��V�L
�k^��O�T�8�_t1�<7)�ǟ�#@4	CɦI]3�CqEe��Z���'ǿyT��S5z��B��J�-�[.ŭ+2j���B����+7�n�R7���u򃦟�pq�R?Y���mQf��z�y(*�	pU-"�z�?���Ls4����'ߛ��D��4}�Ls9�	��d�}�U�;q��SXE�l`G��k�اrgm��#�R�qg5�s���7��ar�MEQc�G=�r����K�(B.u�������¢�q�`fyj�/�X��ק�aѷ
b�z��Y�nB���j���zGQ�M�o��H��5 jϤ�}�6`���o|Z��xr�LZ��d��T.��i��h���(G��hBt���dW�����Ī�v��jxr�`��A�(7u�GX)��A�z
֗�@#��վv�3�KK�<x�� �� #�2�ݟ�0���³U;��g��[�U"?isIsg��8"#�t��Ȃ~W����`_��{���2��:��F�kA[�07��Ӟ5�s�+K�=�vI0�5N�me�]$��ւ�u?܈ߘ��\n?�K?�Jg���Q��)���V�]n FxA8����՜{q��w2����˜_��,�^�-�]BU�&����ms������6������o�πW�G$3�������e����������h�8Y��h��Uw`
����ۺlsh���2���4�DY�P̵b�.R(֔��=��y�q�Q���Q���$��d�C��=ux�{�i[�v!�S�-A*Re�ѓ�$-�^���M�ߍ�3���Q�=�,~&n|mƦ�O�wZ�t� �^a�z��=�\����WD~�v�����沗,| 7ަ��-��n�D��ߧ��{|@�*	�I$k�l�\���:v�V.�RWm�{��B�♢��������l�c,8�$�i��,ɡ��V�h�i��
�{8~Gue���9W�G�v�B��C�`�Nc�pg4J�&o�����	���+�Ӽ�_�=��u������f"La'�D!�qj�&��V.4����bzw�0�	'Ag���{ws�zh_�~���֢�x�*$�h����k�z�N���˚_�M��tᮮ�\Y��,"$5uIm:R��L���P��rO��O�`���X"��k��8�B���:�D#T��E86����?_�*Fu�	�(�ك	�@c�����&B�,༏n������;'Kg�׳�/��ox�^R5�ӣ+&R�iy,0�jB=��$}�@���������M�c�[��E�f����ܵ, {m+	){;�97n���������t���܆��Bv8$܎i&�FA�TP�㟊�$I:�Ƕa��<���)�5��4�d1�R7�6���j�͔v��{	O���|IǴ����`�[FT�qӥ�K�n����ʸ��8U��짩<5Q�I��[�uF��Ec�-%:�o(�v�?�QQ��c��Ci��XɆA���`��P�����/����l>�tјcי0ƭ�x��PЏ9�fkA���0� �=Q�1�Mqm"/�| �U]Fn��,b��jv��4������42�y���~^��& �r���v`�����n7s�V�W�xS�5��(�Y�f��V���qccq����`�(�:}ԳW4��;L�B��WT䡻��}:�pN��QȠ/��PD= h!�Ţ��W*Q%�E��Yx.� ���m��ܑ�Z�35���񲗷"�Q6�Y��i��0����E���x�y�xě�i��ťsC��=�1"��3|�k��+�,=~Jg��Np������l>�� @H����lsqf�a_�@��Bh����	��J�!H�Qڨ��rK-u�8��gx&�W�F��3�Y��!=��W����ح��{E��[v�~���N5XH*/�ٿN����7�|�
`|��q���9����t�W.]�%���붑,U�(p����z�\'����ht��"��xZ-�e��$댁ڕ<����,Y��4d}"�o'!�g���>��I%{Y��<SY;q�Ē֗ĸ�F|
��m���8�����ҒYGߎ�	g�x�~��˘LL�+g��_�ݯt[��x�	I.p��c�G����c�U�d5�׀6O���Vgڋ����$��-�v���#R��Uf�i!g�{�`��d#&���i�i�:{	�e�:Z)�H�R�x��&xZg4_���ڮ[�6��!=��b���Υߣf�]����s��
�i�0~�R0}�V�q��VB�N��lz� �Ԩ���l�gޮ���%��0aC�lO����s������ʹ�EQ���Mo�>��a��e+	�U�����uv��̟%��xTO�qej���V��R*�����%0:u@d�D=��gꄏ�$�`�J �i���Չ@N� �+�� �������bu�������f�2�%U|���F/i� �!1�M0-���<3���v18W�G���;I���œ�h&ohf�C�L�Q5}O���φ�ɓ^�$��1+I+��:��֧��Z���"���W��$�?w7s���[���@`ͭ�4�߳���(6&b�*��0�yrl3��	�}_��t.v�Nf�t��?�u�%>TH���0�}�+#���B/k�'��`��w��3]���K�՛w7�3T�7�|R��J�k����M�ȶQxzD�����ƒ�R�Q3.�� j$��K�骭
�T�0�B�pϟ����B�Xq�EC��R��IԈ?FhЙp��\ԧX�4��j�!�Y!�0ߗ��_�$B%�� �(��'BS4r��=@Glpu���$���~}\G���{Q\|u=�l�g+sd���Oc��w!R��ʅ�7}��˥��Iˏ��)31��9�(�}b|:���8� ��v�5"�컗�~M��������8V��O��>K�9ܸ
p�r�u������xhd�����!H�0:`�"����� C,��'��~��b����M��w���ጿ�<������������Y;؀Z�d�Pő7��j���
b��a-hX� 	�c�D�gg�ȡ��nl�V�hqM��̓��^q6�]?���esK��	�/>��9v5%�i��`���כ��U��\���i}��"����ש������	�~��`	�Z#��Z}�pͦ�d�/?:G���-���u�W�Ě��eb-R�L�o��.�\j}�
T����pd~Z�o�nZ�l�����6rق{F>I�H	X�4`�,I"�>y����!s?�{2wnl�
�"FyجW;j�j�ȥ�aj��Td�,(�ϛ���'���ܫ���YٮG�P���%H�;�}\=���Y�f���'�X�sto]w�~>�B�F��*�ê��UkS1+j٦���5x��_�������z�D.�IRsO�jw�ipW�67���=�d���� �JC����
[q�b�����֓|��ͻ��x���Vt��y���k(��jŃ9����ܽT��ET�cL������O�xd��%����ԃT� MzhTX&��ݲ2�\z$2�qo������>��l���j!�w�����@�� =�&��$���Ue��6 ;�����X=��Ftxt���{EgE���X�; 4`c�G��N����BUk�^ۊK���{J�!M��
�@M��CS)$�&�y>���S($��j�wx���,��W+\�KNh���2�P(?�闀�r����[W��c��0���[�}�������gQ0{�YV	J�b�r x�"�89ַ,�:�������H�H�i��E�2�d&Q0EO�	-"Gcu@�w�Te�۔g�HD�z%RܣR�T�؆��Z�Z~0�f�`����� ���nk�xa��u'�jִI(?q:��*Zwz�����v��	d�"����,�9�B	ĵh���z�;2<�r=�g�*�y0Z����Bl/d��ٴ_�n(:�1�ŝ�ْf��!Ot�����Jl��*�a�b��Tj��`Ē<�����y��2c�3��A'�i���4���3$�`@� �5����OP�
�a���e8�_4��D�
?����'{8�����>c��dt|I��L+`�Q��s2�dMB���%�p�p�)_�`a �s�$�#gK2J��{H9��������!�*��gӆʘy5�\i�g�!��N�G䫋��9�/-�9��N��
�X:ŰY�5�!ɃL���&A�Ac�Bɝ�����e#Rӳ�������A2-�/��Ŷy���>]Vͱ�G#(�Ii�s��ʱ� ���*ن(�ۊU�Qbp��~E�����1JPԂua_X
�r~���,���z������Of/��P��`���{���E����,?˕ăf���8GL���~B=������;A����=�p�G����.�C�2�\����yr4/���7�j�;�U����(t䑒b�ٶ_������xB�v�6�����K���JN E'��ʥ��b�>�蠛�l��e�R����}�%����z\��+�BaL��5J���)��lU��}��s���G�����"�_>!����
���"ٲ�s)�1�7��8�Nxѯ��7��rՑU���&jz�h#*c�t�x�G0���?v;�������xɺ�ѪE�U���	1�[}�d��C��@M>�f5(�N
H����l�ӎR��`C�����M5vﺫaQ<�1�{�v���w��?��&�	���Ц�\�<�,`PY9E-$� ����}�E�:�D��:�����4$�3�	��,��@�lF�_$�8��̤Q8[!�$��h�}�Cq�b�+��ݴ�?�ɉ�ќ���s?�_W�?�p�B� ��X�"��n�@#�	st!S�J��H��y�WH�P����3p��HgU>�.�@�����B�:+��'��T�s����bFÈ5ӲU�&�)���0�g���1�;�R�A����d��S݃���;�E�1^�2'�&���I��M!r�ړE8�'�����W+��tFF����
e��^H��h���8��A��|a~k-NL2c��IAJ
;���T���d����"y�Q=��D���iE�r7Ґ润�ݖ�?�.��^�8�<xLY.��ł��>9�ȋGm���LK�qB�W5�#�����(����� ��xb��F���:�% ��I��*�լ�}v�Ɯ@�b��$��C�T�Y����(x=M,�ᾧ��8��1��q���q�`A�����u77W"�z�P�s��2�C��Y�}�*�x�}Ɠ		y�h6�U�t�Y�m�>��ã �vz�.It�e	EŶa�=�����p�"�7�d�w�M�O��l�[�PW���\fxcW�>*���}/m�gW�I�������V�*UW��F�|75i���YL���*�;~��0`NV�1���]u���ϋ��>�,^J孕�򅺾~���ԟ�z��`-7i�gy�R��_����,�\��6�eG�.ȩp����=7�B����Ee�'2B�e���I �g�A@�iky|7�pvU��$��7I��1�7�z�lz#?~�/,49?p�$3�x��a�*b4�^ﱔS��D �ޕ3�j���J�5г���Z��ZQaL��A	�&���ߝ,мL���`�4��GE�3��v�n�H&�(o�g�αM<�Rؿ� I+��mo2:��R��Ao��W?�g3@{Z8�zX+������O��%�%�ڮZŐn�gi		��f�9:z\O(`����:@��/8~%�J��N4]Fw)✼��bm����� Z`��o#1 ����'���{A>�L��!�Y��tŐ%��ὰ�Y�MA[J�+�N�nXlrE<He@�r�]�޾j̷��vQ����꯴?ӛ�5�&�is��-oúӰ���ɘ �0rT�gc���]�
���Y��l��U|�|ɡ}��u��\hVv�a\ќ��'#0��;HI�:ө��ˢ�^�����w�"�3J1�����z�I��Xaw���Bvs�$.7@�)D3��O�,&�Bd��#SNej���Oc���\��=���]c�����>U@\ �=�qƁ�B�n[�3��}�E;��[���㲷�
�~a�C P� \r��dF
g�}�?%h�9"{s+t��w�{J	��/[�i��ށ+���"�I�?�%9���]F
/���l��lQ��������C}�?l6!v} ���W2�=�D�d��q�m.@�E1)�u8�c�[+!��`�~��sۈ�%v9���MFCtK
���F#��´�0�����z���.n�v2O�4#Ž��튾�z�<֩�
ҍ�6���f��&YL�0<g7@����(���]z�_�h}����>����@�NjV -�O. ��32����շe??`E^����Fb%Va�g
dK6���9��`Lwy���6���|ݡ]K�K��\3^��V!��Q^�G��;$�Ư��ʁ���Rt�p��FG/���U2M �w��2M�o�V���{5�Rz�?�J�¤���U���7��L�l�?w;l���C�*���l��0((6-G�Z|}�G5Uwr1���L����qV�9�c���#gc%��>>u��
������/����諿+`W����kQz���?�G���H_U�n��KEb�&5��*#;%{�qpc���PY�7U�`}"l�ޯ�~}�D+q�/::>8�RkQ��Y�W��.�3p*��9##~�vG��y��7Li�>�z)��߰�Z�}�^\%�]���3��4y�^�1<(�:2P��V�� ��"p�"�瀶�jPA����Jz	FbE��$*S��t{��:��y�ܢ�f���[!}��G#43������	*t�|���	�IBY�9nJ��D�]�pQ�a���F
.ʘ�r�����=DҔ�ľ���i$U�)�`��T �ai������'�v���a���J��R�.Y	��Q&�I
p�z�Y�N!������5������Zm.BO�����%�B:���]�B��	�t�A��6$ms;�σ�+Z�c��X:}y�w�
Tj��1�u?iKտr�x��$��k���Sh�/��e�`pe �Tn�$�th�Bio
���]�z�sss�ͻ��L���&��[���H�^{ڇ��վ�d��%)L{يX6j� ɇV�0�"��EmM�t��w��x��9<%ǝx
��u©&Ȟh�(�c3�ݡw֚+��+���'��y��ٛDig�a
=h�����O��_�Wm�u!,���&
h��XTfC�����H�����:�U�k+#�u�c1`*�I�#k��@�I�6 ��4�Ŏl�1��1JGu�'��7�1��cbwGJz���5e-�c�Lz%!�Sacᕩ
��|ˋ��}�_��1������X�b�P^<$U����0@��N[�_����z ��&�䀪u%(R�-����Ib&!�Ԡ��_�0�bn-�cQ����f�qG��G"&y2�&��jql�����?||=rN�]�[1q�ޒ��?�u�h�tG�!�}�d�s'�z�lO���4`�����]�c�Vc� �vp*�d�ü�kJ�ڱ��u��C�v�gkt�H1���Eq:٣`y���o�-D�G�����kE�mH�'����7ś!���6�!Ke䟳�"����(T��ɲ�F	�8O=0͜�[E�ʲ�{�G�����+_�OqQ���ސò��g���-ߐ��X2�u�����ټ��N���dv:��� ��������ň�cd0�s|Y�v8nn��6a�"b���}�2p�c��%�-n���%�|�H��ʰ�U7=���x|��?���!�y�q;*wL�d�� F��B����o�1��w�k�����T��3�_��@�c<ZI×I��Q
PHH�ٲ����s@, �1�6�c�L��Z��_��[�m��y�9����`�c���
f`|�~�k���?�mi�������!<#�Tw���&��v��uz|P�8�@f#�n�ԀׂҞp������)ؠEQ��Gݮ�-�,����|������,���s����JG�!R�n͆�40|f2���Y���D��
储�3묠Z4xR�� ��b.!�ԭ�]7�=1ՕHR`>��ݓ1���*o-i�:m]�����%���V?e��ɇ�)>LQ����yJQ�Ć�2-m�f�9B�Kx��O����T"�vH}I�����
��aa\2
�LN��*
B���a�kwo�p�3�sXRtDPxG)7w�Mz���*�s/m�D{e��k�����#u�Zj�+�:��]�PX�I(s^�m
�0�è��&' ��b菲��h�hC����6�6x�!?�Id��l�y�?H-�S��5b"��9R.��⭚�6�"����O�ў!?���v�f�	Y�Ve,�/�zZ1�y9�~��8�i��@@32.�&ʓ+�v�L\�v�1���T^4|:3#
H8�	�^�?��ܔsC�@F�S����&� S�m�p���hP]�b�y�ǚm��.~*�H�<��e��ѧ
���HO��2���ԗ��X&����%���r��r��P���@/n�*�G�%:
�DS@6P���A
�	�5����Rw���E���Y����
zS��}�����Ȣ 2�/8�Z�Jf6(į{v���UǠ����IU������-�yR�w ڗ�XD�m� =���*{+��K9[��5H�">>��1@�&�}�y
���,���'�?!���dF�<���~ ��g:�TQh�E0
���U"���J5-��#&/n9 ����X��̠���:���Y����G0E�bgx� �58��6����17�WW\k��ff��%�q��=_�1�
c�LUgT��1��l���=OY��"'�]���D��������uL��)�٥�)v����^md��ST�F�����ϊ�Yjh��2\�isn�e�S!���Y��#��[��X�����NV[y���S�d!��c#]p�BH��}
(G h�H!��@Y��BlI8�eF�-�p7�<�B��G�|����lS���5�8w#\�e!��𾧯�Q�6h�+�:��=	��S�[/�����c��E}EmD���� >^�\@(���;�Qe�b�o@cs,�k���zd�]��B5X�-]�6h:�;�	�s�/�L@�0l9�YW������6[��LS�+@^��Ey�0�]ҡ�/M��E�@^+�܁�4ꪱ��-�|�J�L?�#�$�*a
�FLy�P��gt̸+y���!֘��Hi��F��ď8[��/NnK��6��ť�8j�N7t�`Y� W*�SO ��W � ��íj� ^6��<`�F�&Uy^_U���\`Z�j
�Ii$�(�Im����^	$����Pj>H��W.���:U��@����7�%��6	&�U�F�6��p����61�H)�����t��pI)�ɅZ���픎*�C,��8`'s��| {1s�~�&ӜG�"3ș {�+��#�,�.�D�K�
 �&l����"�]oE��.��#�yR�/B,_�"O�6pNDS+*n�o�ɂ
��H"�zě3��xC���%J���b.@o#eN�R��C�P��T�s��s��f�'gҳ�%qQۣ��zW݃�8o4�|�ֆ���WOM�"*?U@��� V8���ذ#2���5�{�{`t������GMEx��&Lߝ��Y�5Fg�+#D��>>�xb�6�z�p^sUS�F���5�Z6��<lJ!���m5���Q:��;���ޛ�h^$"�a��|���U<%[��7ȅ��:13,�����J��	��K,v��@�u��dv������`�����n*j���F҅C�GoC#F&U�ܞ���6e�X��+Vg?��_�0�Mn��, ��m3a���Q��M?�ýJ�.���Η�����tN�R��R���� ��l�Y��v�)�>�94��#��E��|Zg��
�e��a 
�bX��ػWde@nհ6�o\�G>%���a�ߋ�Tl�"�������Ki�8�]4AW���mXP�Û[�P�L�ܖ��+D�7Q�}�(�%D�th��t�*��"�ͯ��M�PI-�妲P���1`9;���ѵ�ү���$�
F��9�ϖ�@q|�M=�q=���3�a�$!|�Z)��gp�����ꅺ�,����1�}0��>[�H:���
af�yF!�8{S�ĚK�||����M��_n���Y��蜗��T�I�N\�u� �9�3�����ˋ)Z��{fM��k��$�4;��K��I�湹�T�,+��t��(��[�,A�c�#��9ĞZ]+HeNW3�h2��Z�P��@��B��@�������T�����51Θ�h�mXI-�=��
#���W�^�.�:YC�+b�#�r���l�O
5�	%���b>˾�'ڲ7z��eVe�8�cg��4��_f"U�T|��ꮉ̏0<L%l����]�o�a��4F����O��\��Lx�
�@�05B-@�)�1K��������A�yIT�X 8�<_���a�2�CǤ�6c���3e�%Q���������஍br�.ڑT�:��>�ؕ��g`�޹�^�SN�W6 n�}�+M�P+��lw��P������hV������q@2�а��On�tG�SO�8����J���?I?I���䷔���H1�rc;"ecdL*uM^� 0\~�b!���K%$��lB+�/O�SYz�t�S	���A;��3˳�!%���/�N�O��6��r��"V���W��{	<Z�_��\ϳz�����A����Ze���&Je�u�!�Rag�Ô�/e���<f��W�-���Y؈櫽�x����M�]���U�T=�����ϺDT.N�gﳧAm��=ށ{�r�����`�����Zj�P�*�Rc�l�?aY�Q���1Å��o�)�< �@K23QC�]�A�: = �Ϥ>��,N�G�j�L/��k��["��,$���ǇCw1��K��r9�J5 ��#��:��I]T}IIJ}�C�K"+OWE.a�>Y}��&�|��~��]�Ƭ���p�l\�!L�w������C'E��qW�o�c�Շ�*)R�Y��ϫp�g�o��\�-�� 3ת�.�b^�yk'W������*�=��vv�c�}'T�jU*�>>�0gY��+ �LE�y�V�c_VP�J�W�v\Qw���Ĩ�!v9�&	���S���q�z���K��U��Y��>U��R{GRVg5�Lۜ5�1i��1���b��V��|>��`�W�v�E��9x�Pf�N�N�x� '��=cA��%��.cz���+��2���K��%�Ե��.�`lAIf4��o��3O�"�gr-,��-_���4-X�U���1+��m����"�FA``]��Z�;�NyY�Az����`id�K�:�n����H	����KG���� ��"�k�O��Ixlɪ��54��ALc�e��~G"ǋŭ�q�毪?�{D� \�^^'\��c���S�j��-ġ�&n5����ܘ�:|�2p����Om����s�M%��!џ/����K�;��|����S�m4���h��?m����c(_��ʽ�1�N���0������x���c��^_���χ�9�7׀3P1�4��Jg���{�C����h���^�m��; HLQ���J��]B��h6��j�	=ca�!/�-w��X+��~�V9L��؋fʮ�����þ�\Vٛ<F}g��&��r��ҎZ`�.�[@��Z�h6����?ejBs�9��_�������+�4������_�"82kQ���P��N��A-�@]-8���Њ�я�pĤ��?q̦�ӱe�J��,u�F���|q����$q�¿��Q�V�s�䎯�-h��/f�Z�[��m
B�;��U�oUP��&�l�"�8��z��O��3��<i�9��l��a|]};��4l׻���.�"���7.�t�Op����V4C�4QrvN�0p�AV��k׆�ς�������l��M�c/��¿|c����޸��s�f���#ý���h�@��z���״8�C�7�8��<�8�]i���e��Z�gY�v/51'��0��.�,F�B�|S�F|��G��$��&X�0kX6���G��O8�ѻ�.hf
CW������<HaR������ks|�*���,���r ͆�	4��6����n3!��'�v�,T�t��~�I�#B��lw'��H�'�щ���9�
qx�1�$�b��Q%d�4Ib��at�@\%�����V��Hdg����gV�Z.v,l1M������c������:.�μ}-�ܡ\�7�����z۳��'��5��� �q�r3��]н�hݧ1(��9��W�0>���H�?�#�JA�����P4*��4���V�`���oc.�h3!��e=A/������q&b�Ӱl�󂏱�����X�[�a(c�)��L�^�X5:���;�t#�'�8�{�+��X�*^:=gy�1�P�M�]1 ���V�1��@�!�>�i�^f��k6iϡ���4&Ww��`�cJ{8�j]�+�%grH����8�8BM�Q�����������96�W&݃Ka�
�0ɛ�)
�sϥ����T�S�ª�B�z	�l<a����Y���ksd�H��X'kZQ�ĺʩ�Wpv<��1�ְ	PwY�	׸1_\�$��ݚ�$�2i�ae��Ͱ|���\�
ٮ���K�� �Tq�@_l�=�c���<*�An�����||�hA��냿J*�l-o���@x�ts]��ނ��۟�j���<�Y2��9�s���|�ǉt��T9���s]Ь���m8R7Y�y����a�Jd����oNUx@J�-@+Ƃ���?�NZ��>U�C�~e_�L��;0����^���n'M!��5��K�����q6���`1��YE�.,����m�7H/-z�U�s?n*X�Wxܽ�	�R�g���((�tH���b�#ǣl��6����L:�/_#S��!��qCt��xu�W�e/y#P�>���Ն������1����[���k���q�g�4��uK���u�xe��~��-Ds�q�֛�� �&���W�e�p�yZ�M��X�Bẘ�*�,�-�a6�<˼/����4�5�Z�$�B/������i�<ÒO�n3*M��堥��{��ܩ�b3�;�}��s�R�*
O5^) =>,�RR"�F�Ҭ2�(�+�-i�Rx�wJ�Sۦ6�O���-�z�u*s~$K��.���a����禣��۫_xQd8�Z4-�k���Bx/Y��oO&���lׅ�ʎ��
�#D"+*AUZ���@_P��P�|�O��z@����VJ����@�3�@e��X�}P�ĩ��!`�_;І=j���L�������wUuH�/8m��p���<�z6�s:�8����Z����`FΞTt���2�Y$�;�d� Ts����˘Aef�X��Ql>��}uԯ��vH ���6,s��J^�k�5T޴�rKp�ix�PX~C,|����+���RF�!2�|ą)"Ҫ�7�E���aAu\����	-8w����ǋ��h���Ch�{}@꜠V�޹DjE�y���Z��X�`�.a���K��I��#����Ӽ��s��(���i�HZ�
�zR�tE�*��3�Z�a\�΀��3dT&|�L*�2Y6���+�����B��?�ɰ�Np�m�ϩ��@�Ǉc6��!u~�U��ыI���K����^ɢ�hg�}����M��8x��n��p���n�0v����������d��Rol�����UHGbs���G��1�����ԧ4x�M�9����]�q��rG�@ _?~����!y��X��?���
� S�����P���`@"�[�G���̈kMa�Y�4R�D�s�� /��)�v�p�Y��i���a+4���m�=�#k`,���	��T>@�Wz�P�o�8��KA	��kud6��������@P�~�}��&@?k�j�
9�C���P��ʭ롣���2�v�N%N�X3$K�`FL�m��&=���/��ְ�U���d�A+�"G�Cg��)���bѓ�d�XF��ze2��<�������d����20-ՎW'�&;��^u̚  �I�T@�׹�Jf5�(��7�y�+⒭�R+�C;�Hk������A~������5E��x5f9�>�ۼ~p����CPx���r�|�7���ҹ�$���M}�{��j]� _"�기�19:$��2]S���pE�+�`y>��@�f-�q��}iM75��V�$h�?u#�u{�wuA���P�N֩_M�hp��։����DAh����g��!�P���gb�$3�����l��*7��r1�%�н�s���f3yt�%�O�m��I�R�X���$�� �.�q�Kk4$�7����Gڤ>YQ�x^�K�z~������Z�h�mUl�1�����\2���Q�z'W!�'sG��K�M=d&0�T|�5��.n0�2�m��F{<W<U-�̆	�F��AO����	L�]W,�{�{[���nc�;6?&��G�#rl����8�d3�30d��Æ��f�k]�ej[�����J����/k��Y):Z����/Nj
��}�I�O�T�Pl�"o0�F��XK��
1��LљJ�����*"�ծ8���6��<W׍y��C�97����N�"�}D�]���깟�sH�9Ϗ�(��M!���:]�B��P����}��2L�^�9/HSS�rWO�B����5��U�.t��w	�'K��)i�/|��2��ե��8��o];/7:y�1oDφ�%����P^��w�ʓ`q{�L5��kƤ�n��+(N�׍ʞ���v���uN�Z���ѢV�6V�c�dl�����[����(R�s��T��Mh����]Xш�[�X����N��{E���e"}��W�9r)��'�/H/l�QcO�6!�D���g$��l�p��Z+xv�>u��ƱV�����llR�� Y3�����i6�T�$�h�cq"/��)5+�(a��-t�2�CX�u%�/��ڵ�14�Ͳ]X�I��@�u���#�y���tW��HK�#pb�\����颃̖sJ)ٯh{�̿��v�J�XOnpf�x7��������>�dD��D= �F	�:�`��H�r`�)����=J��ļ����������z�퇳cC"ϲ��fa�fmJ`��:m�G$�Mՠ���w�ö���%#boa�(�^%��L5Oh���6��ͤ5�k�6v�;����`��XY����2`2�^	�˼W�c�� �S�ǲL������~|旜C��S^A]lk $I�au����D"��N�^� ��t�|Rw���,&�;����7�e	�+��a�u�*������>xc��)g��w���G�6��y��h��>�x�7��N�0��3�m� ������c�'-=�_p%�g�uн�&h�lb+=�.���a��E�Iآ7��V�} <�1�Z�Gȳ��B��cJ���(�"��Ԛ���/�Ѝ,r�%�NO���[e��l4��ܔ�� �)|E�oRts�_�gL��eN��e�mw w[��c�s,�l�T�N��0m��IL`��tx����ϿhaNG0ǺQ&��I�Lc�Tr@.2!�~�ۜ��D#���'�]��ʁkv�����ʗ�c��M��̝ޚ�=,��+�k��2��_�:CY� �	2@���n/$�ݡ)�i����p'٭�p8R�K�n�o�I�G���]b�N%,	�e����˰�8�?"�������ga�;���?&>.�5.|�j|��b?d���m�F��6���d��m���5�㰈�R�'՞�ϣc�d[2V�qZ9����:)(ϱ�C	ʕk�����S��|؟�N�I1$�uN(�������)����Ӛ�	͓�Y+���ێf�\*�`�:�Ɍ�H�u4O�Ծ���?���U�m�4�Z���\���Q��1������ ����we���K ,��q���B�6e3�o���CSN6[-������k;j��W�az6��L7X�
1���wR }���� ���tu%����&j>��,)��{�h�f&����84nJ�Dy3Y�%�/$����ڕ�:}�<�rGw�i��J�1�C}+���n�ŷUq��q/�Bf��>+�"�7����6��G+Фu�om�ܵ6g�YG���Z3��/��+K��rR�D�;ة�N�AG��${����6M��"�R���:KVް�Q_��t��
ܖ��؁ң?��Rk*[���4�6�����em��Ǧ��$A�h�Z�����x{\Uj�5�>K���5�w:�n��H؃cq�xD��9.�|n�B�z����-Ύ��󄺁�Yx7I�.�����`���>o	���]���\����b�z�}��u�mgU�\p同.Z��d
�$?Q3񎋯έ1Af���1^?���W~����n����Y�b���w$J ��J"�2=\�{ Ώ��,B��j�5����~�hj��Y���(�q&�1(�\��T/�;?�#�k���-�b{�.xǃ+� %:����6CN5:��C���6uƌV�п�.xQ�PZyB����l %�N�C,���'Q����_ƅQ��3 ��"�LN�}�^�,���s�uu�Ub��a�k�+�>p���_��9��A�~!rVhl��o<��՛�J�lN��5�%U`��D�s�����X߈��4+��hwo�R���>������G�LȮX豀�~�V��;����`��2n~�6;���W wR
��WwA��dP�S��:h$���<a?"ꬶ��?�7�T�J�hLt�������!�2��=�����ˊȊ���� ً��-C���!n-�Qs�|J���>�h0��֞Pr���Tf56'���)�.�q�QM���Yd�H� B:�����w'&5dN��U����8�
aTX�1�g�UZ��B�G<������B�k�������])I�]�hٔ5�
�T�
��/��B��K�Ġ��r�V���V�����Ϋ���V���@_��2v���B7]?,�knbn(z]�x��?�����G�1%cF�;�Fg<�L:�2߫�cw�sn������n��(~��K���Q���Z��o���'���G<A�k��cO.�i�ծKn�8�|kYu�޸T��RJ�Q�L�)�
�����Q�و���c؈e�bM�}Ի?�#�t,�Wŭ��r��r�䧆O��7?��.� (՝�aen�����% �3b�߫S��iK5R
��c�DYΑ X����9�A�/�.u<d��	#��[*"��k��B�
zo���{�i쎈�#9DEk�H�$��*�}O!ʹ�Wa�W�^��+���a��t�S��èT����<�.xd��A����cJ��Ώ��d��P�o����Xy���JŸMz�/�D����{}��,��/�L:9�I,UV�d�AZG����q�m�R�?�c��ܹ��Y ����Z�w��?^�S�ƾ�G̅ZR��S{ٽg����D�w^]���'9���beF2�v�.%e��Q /�^3ϐ9%���;�#�֏E2CM<�
x?��OT�]����ѓ����C��,�N�Z�<�n�A�_�#���N5�=3F�Zmu���y��x˛�r��83%.u�>=|k0����;X��q&5=:��|6����w?�S.��&���Ю\����`�&��L��w�����q����Im\���a3�dI=����>v%�)Tt����g��W��_�]��k����qB������H��h���a�!ʫ)�b�%�^}�U25n�[�5�0��K�D�2�AA��\�`0�ޝ��@���-d)��	���w�%�ݐ2X�
#��<��C�TP�0lU�/��T�����N�O�T8b3Т���{Z4������	�f=��b�[�㞀D]�m��y�db�N�$�Qٿ����&�����;C<��J2 @K�'��3~���9)ʗ%��Md����J\�����K#�Z�l����$�GvSc
�IH� q�fB�>z4o���*N������%�C�z,��W��]�Ju�g�@+U�j+���D�v��$9&pgdy��+��(#�ܡ� �p����!Y�t��� � �?�w���N`�mY�X.o�����ʺ�����	!�BG�;ҧ�3ݜ�<�ܶ8!L�.���0},Hи��u�%���tl���.��ӎ�u�W��e��ã�?��o��<p+I���l��VU��f�����d�
���1=O��Y\�T��\Fb������#.��~92���j}_�g<��I���2���)@3�e;,����_����S�5YM���(�.��t�}`��Ӎ�p k+���� ���peh��r.�������WL"�GqFg��!<$1��e1� �raf��%t�_w��bC�����R
����������Ǚ��1�yL��ˠ��*f�	Bt��`Qj�N�e8`��l�T�^8(�s������`�C7Xܨr�Z$��Y_Дڄ�DI�_0:CT�]�>�����pfr@�jd�ObQ{Քoxi��D]<s�@LT��t���j�������x�ш�|��>Z��ns�i/yꄾ�l-�mJ]d`��u��"g?�<�N��t��z�;�P��S��9�2�=��HL3���;�@�9J��X�R�[/�4�p���%f�'�[���+��}�H�=(P &�F�ןÕE�KzW��v���b8���&��S)�]0t ����+�� ?G��k����D�r�B0��^�� Y��Hp��9��M��7P���A��ɴ�PX�Ğ��`��4\ưG�0-�Ï�Ƹ}U��;I���F���a�J��M� �q�n�[�(�b�3�j�X�l��n1/қO-~b��T�>+k߃TO�(�a�z�w��Qb�Rه��]�(�YE��9����Y�J|kt�_�����5�#�k�՚��:7]�IҤ����ޕ.�̺��&BKA�����!�u��6K�{=��Μ��u�Lf9J���rPG9����xz�_��%�r<y�t.�}�I���?�q.p����,�mE���O�c���� YiE
{ ���8[YΧ�;;�u@�s�`�Y��w�2fn�t�Rr��z���{S�g�z'6nuNX�B(���J��ڦo�G/=����9j�d�뉐��*�>]4 �c�L�)KG�����{�*���?����#:�e�	7�b̒��+eHg-�f��d����aF�=C=y���
N��4	//����L��$IՇDp5.C��W R
�w�2
���+�392�m��OG���$�C��'�.���	 ��x0A���|��ńmc@[���Jb�ß?��xA�Ic-ݛ"�{էK5j���=��5��ۭ���X���K�4����d5-�^�j�J����[��AjF`��Q��R��dD2��i�yڜ������4��_�R�PnG���x���^<UlV���7�`Ӏ(M;�		{�LM� y}'kh�[ސ�)>ܦy�(��jB����!��]G��X��'�K����Z��}�ۑ�S8�K���7a�4�L��l��%��[D�z�*�"��$��{=�������TN�%C,Q�����{�j��������"�,D�yB��1Y��e�[�lfYh�x_����3��y����������x?��b�m447����<�n[�5�|��V�L���{ݸKTȖ"fv�/�?������0^�Tk�0����igZ��t���j�.F9��G^�|KtR����Һ�l��V�1�_��
����{y/��ug�9�Ǚ�.^kbΘȐ����T��sB�K�.%���S54�3�&4�ϓ�8�7���X=���4#
6B7�2l��Ͼ40�p��s�F��Ly	<�Q�(���}W?2իr��*��ɨ��\?1H����iy���cU��:.i�b{K�.z)͎�A����\I��{+��� �51�j�	�,�gbs񪍆�-i1���!�zl��lD.��
��cե��I�nxչ�:��#U��ڬZLT���Y{��l���B�R <���trA�<?J�氂�h%5,n
�?��a�w׀=��I/�U�/�x��=~G���\9�G�p�_��<�0�����c>6��y28X��a���!�}�P�r���V�{HlaT�����8�+F!�dm���"`Ԯ�,���F$0��� ����=��|�
�/� M{��'����en�<�,<6�񱷻�:_^����(��GY��	l:{��Ļa�����no&�����T�"R�����&����)�W��I�0@(x�j�L[�z��XK�HoFY�y����ɟ�d8sHPwRhz:j%�7o��� �������#��Ԧtf��|O8���C ��yVþ�h��.�����\9�
����kH�����d]?bo6����2�x�`���;���`p��03	b��� ���7FI}�3�>��dnXX�V��������tIY|�*He�qy����L�t�:Q���;��'�_<)͘�̘)"P���������eZ7@��vor�~��9�5B�pC�*���Yq�:���l�FR.��.���coe����*+�;-�}DX� �3,��!�p�	����)���1� ����_i�ʍ��������&4��や�1[�hf.M��P����\�����ry����	��Ǭ�~�b���C��Ck�N�� yoV�6u�.�|�&�L�l{+����fY΢~:�4��.��HT5�%'�*���+�Ѻ���W��xI�
�;^`�/�+�uTY�$JZ8�S��~��`j�~�ͭz����T�������h�dr��nY�W=ϳ��QY��(�ӛX�Vlշ�����E3m��i�I�?H#J�7�S���P��M�@bh�oaL�S����hIy�9����jj{,�U�\k�Ӎ:A�]�~2��3��XȖ;p�������BV�6��2Lp2)*`L����P�eWM��պoY�#ǁ���~B�	5�r#�,�+9��4�Wj�C~(�����}"�_̯��b4<΍�p�t�Q�m8~���z��񪦮/����xOX��/e�!Ur=2U7!X;��~ �ƣGo&���Ze��ND���;�^�h�� Si\W��@�Xs���:=fV;9)�|�*!�^��p;#�<�S��+Py��\o�����{y!8n����-m�5������gL:�	E����K����?���_Ec�:|7c�g�¸Nl)(xI�-���:b�sǒ�c�ӢвC�B/�4�A��R�3,�����F!�j+��A^7ĘGf]��_$�p��:�W%�:T[�ԓV�
���X����T�g�k����{E5��k��z=P���Z�@1B;q�F�zl*"��P�ݳI���XTF�8{��3Ū�>����`6�  }����]_��0��/�wH�4���A�H*��e^e��߲�+�|��U��)v^>�%4��Dr%����-e�f"��)Ф�t�\蹠�[Ɖ��K��vz����5�����t)x�"�B��(1�~��&�[���XLO}��+5[�Ӡ��k	��<��<%��i(�e���T:��ᵅfX≚V>�.`��8OH�)=�(�EJ�>Q=l��{�J3(��f��/����[��%�v�I2�� 5n1�o�oQ
����[�E�}�����cH^rԽW�%��m��!`PW����v>�sw�_�I� ��b���{ԋp:>�	��-����R��e
�7|_%1��"z��ժ��޳��o2�D;/u�Y��8"���v�^Q��z���9��^��4�R�>���SWi�=��:��/-�!���+g���w����)��x�$2c"i_� ���\���J�Қ��ǈ�w2qo���Ce�)��U���[P|&�xF���UO��fG��_~�-��J>xFi|�&I�U��<55������
��&�KG:I�̅��u79�j�@��-^����j�6=0�?����ج�����@V4��5z�"�|�F�1�i�'����x�힍�Vw#X���>��� ^$#QG��N|���Rd>]2"�U�5{�k ?�X����� �: l�Vd��;Q���2���K%�a��˃@���
�TW�y�0��-]ڼR����=�/�Z�bC�o��l��O�!���w��ӹg�|_&�Y�IL$���{/��)�W����,������Z�hH��������
R���������j'v��y^��f��Mr�*�k�팵)�5-�,�0��e2Ҹ(��x�h���^ł��oN2F	��9�dQX�����\NH�T�OB��h�i֟<(
Ȍko���j��Ky<�
��z'�Z�&��8��=4�N�(g-�́�'[�,6k�A��������Z�K��\�l5b�k���[��/�r��zN,;�%Po\���BI��4�E�������b� �x�nb���!��D�?���>�T �$���}~ ݽ·	�$%k�.W0��C_��n��g�{�t�j�p.��B��O��@���K9g�b��VJ��c�"���MI�	���F�yx<�r3B��Ū�j1��|])F���X��<r��hB>�	e����k9�w��&�ݷ`dҿ���)U�zXs`>+���>V�.��N�?��s	E>D�ܵa�W �]����Ѿ$m�w ��{;P���G�2��RY��d<5��s�+DX��+��z�r��"�	�1zxkwD�~��x���
;�M�X����T/g��D4���K=�ټ�S���k���M�N'r�s+n�O~[��m�YC>d��xb��Ŧ��*Lp�<N��1P�?s�&�ۦ5���ؒ��c���.��{ UHhjQ����~������J����wCU�S�=���.���OC�O?<Gς�2�{"�*��@1�w�X^�>��WV�LF.� ����p�g��2%2L��myZ^��gt�IlC�u�-����[^���P�u��˼!M�o9&/MI�[���$>�.b�|����e<h%
+���(����}eŶ��o*C���6 ����놅 ,���j�nvY�B]�Zb��+�����&$[U#� �FsCi����V��SJ��]+�T��F~�sa^�~'�o�ۢ{�;�v�^�n>�	����*�ģUϘa
�V:�rpr
vV�:ʩ:��m=����Z�>�+�V���!�apɑ0#V��}\�^���bv0֕��b�o��/�h��J	���+�
ǟL�ۻ<��hlP�W��m���J���������,W�Ҩ�;�dbm�[�ND�l���T�ḧ���jBpI�����"	��[X�p�ۜ+즺kM��/bN�ތʆ9�
��Qŉ�7P�E��e6���k\
�����r)7c�����r�:��:RBOmQ��ڥ������ꨎo9	S�jW@���3���.~	�s��f�X��f�'�~�`��`��l[d��,"����7���8|?�[o���d&>��p�p���5��b�M�#�:�S�Q�8���bq�[5]�aE�"j�|/�W��m�7�����PM�K��Nmv����a��S��¦f�?� �W�^N�K'd��9<|K5���Q�M@�L�5�t֋�~%oG�c�S���4��|�\��f�z���EJ��80�V���IkNxic�~��<�U����/ߦ�S2�!H�>�K�"*>q=vH9��ڙ?m�\�O�\��`�YH��i�����W���q���C;D�(�~Ǳ�d�#`�b�A���!���Tq�ev�bc���Bn�K��v��hy�ǚam3�<�jί��`��T�6�����i�l�{Ls����m��E���*�{����+h�R
�o����S�h�?�:�
8G�j�7�>U��e�����$ይaY����%�*?qߪ�F�%�	�w2�Z��K��8�Zɕ��8��������U�Vq�#RQC �6n;d�e18E(Ҏ>k�Zgxg�i������̽�b6A>����U�B��E>~�#����Uj�,��F��f��U�Ǧx����c��L�~��_��]�"��V��$����b���4�Z��i��c]���pk�sPv�q��e��|�Z�)|O�Z�1��S��%\�'|�&�	�:_�C��N-�K�ԟ>+��艐^1RFq����1d\�-j��JT�������	$7I�
�oN��홤 6�ꉧ~V��YA5x�bI��o�������5� �7� "�)z���V�/*#GQ�!>YK���$P�X���a����i\V� �
|2����^��\;�l�w������?��H(2�"wa�%�u����U�ầ���e���6��nQ�L|"����'+m��K���e���������:��:1����Af<ݮ�,���ݽ�;���/k§Ջ����Bw�0��H�V���Q�Cq��7n"�8pt�~Je��ś'0DL A����i���ҋ!�( ^D��R��~��ů��B�_�CM�����O\`�rn"��u��/)߁�ܵ��gl���x�b8�"��f�����s����L�Cl���5V��~�< {)�7�1BU�����r�S�,��;�Pn�Q�2;M�蝆�F'T��[�V��u &,[��_���
�԰^��K�l���D��u�@j��㓧+v/j&v��;��C<���ܒ�>9���L����K3VtV���J���_��@~��:-�#K̘�r/h�`%��<k�m3�l!�!Đ��pj`r�^�Y��d�3M�=SWأ鮓6��G���g�s�ך�n�)O@�k �޻�8u�hI�ڈ��jQ�Ӯ[@�^`[��<�bW�}�c�٥8�!�$wd��F���iLI���0C�
�	�eA�H�ۙ�I�Bo��02M�L6�`��_��>�T+6���ҵ�:R�Џ���A���*+�y�>j<�����[�E�}?�ìd��>���Xn<P�
��\����1!6�>�<�9�^��r|c�e���~�p�4L�_���5*���u��JX$)�T���erj*�_8g)��vY��@��V ��v�q��1�����r���<���B��d�����'5�����D�������E֙�5��V��
wHL?� &&s��Ч{�F%-����T,5����7��S�W��A��ɬm�U�-�0Uٝ�����k�b��ו�Ȭ����V�<��nRz�z|���Hʦx���0-}���$."�{V�_lJ5+>������s��|$�F�p����Ǒ���F��#u����9S� �[vq���pcf�������x����e%?Np���d?0ޏ2w͞��
ۗ"o��|�TLOv��TrY���w����F�(��k���P4P�U�H?�����b@��v
�뤼��ߥlQɍ��v�7�xXm���lz�?f-�7ݏ�HY�{�ĕ`�e;f!��Z�5K���C����Wl:~�PΪ��.�|D�L'M���}���hlx��x}뷔�3�Mpm�P����Fy��� �l������I��⸅u�FZd�
|(����ah�����5�5�;tu��C���4�(H��i�Q���1��jd��"l�p��y­��3)4�륱�(�J�׵�Ǚ��G3��"�TtN�KP+~�����P�ˌ�.��I��?�]�Ku�G��.v��ȡ���%6��]w o_ ~�f�G� p��?���cc@9�S��9z���W�Є��7�c��!Ԡ���s������%�
�N�}�voWëw�c's3]�{&ԧa��3��gz�ou��1=���y1h� �9+=��n�Ј��z��ͥ��T��7����
 �`��鹝�3#�ۧ+���,h]^ lt���Lj^�C{�"�����Q�Z�9^��;M� ��
m�]_P�M���/��L������x5Y �h:w��-c��[r#JS��jjR�!|�jF�:~t�{��GIi�9淤I*�S�0�u�ARh�u��l���َ�aS���;B��pZ7n�$�����*C�%t��K�ۅbг-u�Mm,����F��y_�� "�t����9��Nh\S��l�(�l*N��iVp�t�t��;�d��a�3,�"��R88�?�J9�S�)b*c��l�~,?}�����iS�v`�\� /G�ҵ"jd�N�հ@G��Ϡ��ƌzp-�?��L���<����֫��F�]wP����ŷ����g�"�X�m��]�+9@ȅ�m�[ꆺH��k��r���b��S��*|�l"�2���ɠ��C�,�6\{螗d�� ��LZư*ƽ{[+�� ��<vT=�#4P�D�`"q��\L;*�Xe�J;����B��L�-E��l_��_�+�Ok��b�(��N��3�GS�u���������pK�L�9�?%�2�|�}�2
k���j"Z�o�I�撨�S۠2Fů�VG0���Y_�w�n���5�=uk��)���9�,�*���<� o<h�4�/Qw��[�v��m=nR�����az�lK�� ki��R�e�b5��}��������6����F�H�RU�;�ô)��
^|1P�N{
�GȜ
�#&1Hܤ�	����J:)�<�����Ei+��%�JkS��<�J`vv�9��k��v=ҘƳNJ^�=M;�0�1g�b�;�5]�����v�eRHG�@��j��[����F�NN@�r��7FPߡ@��:$��.�HL���H���)5��4ᠶ��)��)�^�}�����&q����BG�^R�[��;�Rg�L�Ј�����Jd\�����+�'x�_sH�r�;fF�$�\/�����;�r�i��_!5 ��vqA��u*�@��� ��[	����pB��r���p�������=�6��`��U��׶ �[J>���Nt�G~��")蓾��f����g���]���Z*3�b�ω,qƣ!��d&<��1�d��~R<��1��r��'t���ه.��f�Wil�4TD罰e��S��.Ε�<�.�&���������'5Q��\��L_m|�-ɴ�Z� ������VB���ƀ�l�>��`��A�Jڸ���å���[+�2U4��$̹!ɋW��F�"qi�*?\��Ht�"?�X~�p�:��ْሂ�2��
���5��y�a�T�+� �h�������7c�/����G"�2.��l��.l\n��)��ʲJ&z���͈����ϔ(�^'��bq�p�\���d(�fm�~Dy��6���������s~"lf��2ۊh=�����I�e���V\R �����{u�F�g������A�� �yO�a|u;��7<Y�]Or��y�{2��k���Y��lxh}/���:�޿o�k�!� ݩ��y�Ԯ�d�Q�G��y,���!������ۋ��-�m�{�Y�c���e���P&�\���3��u�Z@VnS��=��O�B$�������E>�y�>�ޛ��e�����7�3x�Š=O� �<�}@���9�ɉ|���g�P�JG�=Vh�o*��ǟ1��6���t|!M����F�6vS8���7��~�=}��5a��p�ؖ�N���������X�f�*��v��H葻�lT;^CN���_GPm�LEN�QƼ�����e�׆>ڂ{@^���`���3��g~
@,�>a�'h8���H��)���`+2(����]����~Koz3��k_�6�c=]m�����J��,��0���n���==�ix� ���x^��q$(�\m���oݵ�� t�����8A���o$ �]���}��!�J		�an}&]�̮T�����;Rp�|�!=l��;���1��*~�����j���ܾ�a�.���N��0h�3�`�Ԯ06��"�Wߔ�sF���:��˷s�qT&1L��E��#��̖�Iv-���<��G�Y U�*��h<��գ�Y��C ��a���j�.��GQjgw]W��	Et�!Q�B?V��W�:Hx;�h���w�U��?����'_��g�ߺ���ݥn�{�8q�h���Q�R&�x@�Ə��������;���t��cq����N���&cI�H ǻ�0O��d�3kو���\s:׎��U�BZ%|����Z����^�-��}��@i��?�r�P�����g�k&��~r@O)se����p:C�
R�Q�R�]R�7���e����ݽ��>��aB��wC�n[;�ER��� �'}~�q�x7��M�,sM����awO96t��A�'��� �r�b�@��<D�\�iD�v|���E�
eW&G�d9�Iƛ�ؠLP�����E��kl/�هAP�1	�x�iQ�G�amP?NsJ�}�z����G�K�S�'��tSǮ +��1��W+u�m����\���DT�5<�����!U'�u�kg*l�֦pfچ�H.�����W�Y1m�*U?�K!��B+�.�XĵVZX�i�8X�+3����}�����ĭ�l
��{���\�B)r�p�7�����"*�)�H[�*�,�lH�Y|J��ӎ e4=�d7P�-�����O������1�P˲�;#i8wK����؛GQ�/��EFW�e�"%��x7�"��-,�T�3�x�@��%��7ur� fW�Bn���Mf�	bV1��q*�7(�6�&-�52�L�����j�8�N3k-�ǚ�t�2�rH.r僼I�l���>/��Q\�ۖ�(�*��-�y�^��^d	�va��"Wa;Q۲�eX�2΁y�ԕ:�&}-_�Xk�
���496�!��u����69�k�]R��1ko��`!�ل��,A���4eF�~�c5����_���X7H��A���7Ц�#^v�hm���`�M	>��p��%.�ږ��ׁS?�8���G��`3*�iWKt�fRd��B�9	҆Uҳ�)U@�D��FW�y*bF�����[Z8��rWm]Q���n�z:�.�t�JN�?�lQb[+1��(�R��Q��zʴ�?=���?�vi����$�I^F�U�YE&�;wNj짢w1Ei�+�f�����md֨�㨸��a�f2�V*JԈ�㿏�#�x�o����9zO���ˊn�UEJ���_�Ŕ��&���T�/6��n�?�;K&���\�F��}Mj���eE�/9�Dq��~��2P�GU�Կ�4�[�k.=ܬ����.G{�^r�%M�����SL��g��FNq	J�ܘ�!G@4Lg���6D ��lUD7Ե��5�@ן4S+���Ԍ����%�8"g��A����dm���8P�� ��/��<^1�� `��㳭�[2�*6\w�ƌ���i�B*��^�kWr�%�:y`Z�cf+�,v��D�C0Dr��яL�U��9��f���NpO-�e&l�u$� ��R'��Իn`H�,��Gq�I�pQ��*�_/'�i���{��@��@-2����uW�Uw�?���e�u���k��o�=�U�Eqe�]���*�����o�wʝh�&x#�R6���Q@���0��{w-���~`qM��T��鍉��f��i�������TG@�]'=���@ݛM�YP/0@k�kP��d˗;�-�y������`�Ӱ
�8G���n#~��'��y����p)a��1,4���>qH�g	>,�DK5����m����M��A3��e���?0��7�7���z"�S!J:<࡯�[��Yۻvӹ�Uu�2�Ox�F� �0�-����(x0[�^��om�����)�i���2�d�"�w8QB�)�d]_����+ Mo�0E�ǔ���#tRaOn��m"!;]s޾�Ud
 Ֆ�k��� �'�K��'m���7�@l��L�q�j�"��|��׳j���erܙ�������=�'�M�f��$U��E��Xٿ�
�f>z�|Ӑ߷�!v��`�*��bk�dO.<79�{�%?DbL����+8�����;�.t�.�.#�y��:��'s g�o[�8�������k�T��W� ��@�ؔ��]��ʝ"}��@Î�1�T�qEB>So����ё#�:�)D�N��j>%�Ӡ�N�+�T�~���H.b��ں�v��cW����]�p��p|���R
23��Sr��`��8�S9|̍��.ԓ�<������l8`ǧOgG��H�e����M�(�u:�������d4�7t�u%T:�p7�)q�_�wy�"�,2�8r�*'����[d�B���"�v�[���:�ʐ�)���R�A��׶a!q#�)�KGd}.��\���z\S��0�����H����SB�,/��W՝J�� �lk)>*�C�㕟��4%����=���AХ���j���bxŮ$r�PE�q3��@^>�nG�<�v"��ʭ�@
��g{���ĵjW�3��{@���*/�y����_./xq̢��i�FU#:�w�{j�qWf��sʛBL�6��^5+w\�:��`��=�u�`Hd�����������DO��?d:����Jr)��^R�^&����.�Ox�gXyã\�ƹ8�}�u	-D�@�l��Ƚ����6-p�\ixхk"Ω��:Y9rC5]>���E �Wh��!DY[q�2�+�d�U��+a9�V\p?��cV���/�gF���A`���5�h��uOؽ؊�ή��/�}^�yN��:G�95v~��t�Yqg��u�f+�HQEf%2��ql���h0�27}��q���\K!jI7s
�]ݡ�iN^��ҧ�d��?�O��.�%����"��8������� 1�`���M�[�Yx�����~s�QD�3���<s�o�q�\�����3T�P���iXE�d�#��a���V�@8���@��{		778ޟ�	>R�L�]���"v��P�4�I�5v��aOX��$@�-z?B𝲣�m����WU�!��6��rj�g?�k,1��`ƅ5���f?g����^xm�2{)�꧷Ǟ�p�.��N�7�G#oU�{�s֊�/���Ă&� Pa�{۷�k?3�uE��WXF�MH��g mމ[����ie��'�oj�&�7ff��Bo�:4T��@Z�s���&�{����^�q�����P�/P++�ȭ^�z�i3[��΅�y�;�0I��7�q�Ȑ�Y5Vf�f�z�ӄ�ò���'%��j�7u�j+B%"��:M���/�H�Th|$n%���K)R�Y��QQ��S�s�؎.0w�ݬ�dl��0J��ca�Z:ԕ��f���^kI��jt`�8b0&؜��)��]��y
']��MghcF%�`�:�F�jx�O��y�����s�6{�u���t���5��AQzb`a�h�isi��E�u\!k8ah�V�"p�_#
U�h���ڃBWGy
��Vf��uц����&'�}������%��#�X�+4�%� (�b:�� I�Jz�y�OD�~�a��t-�i�Xtj�j+�F�Ǥb�KJgM��:�Of��Թ�۩9�&��Ǖ�e���VHn��NC����]��F`(�����9%����hD�Ԓӂ��G�>��&?Q�3����7yw�N�d�P9�����
�$J�,闗������ ܆�z2bh�<'��~{K�^�\����Kҡ��L���C�>�k���	��sA�ԿhᠺL��hɳ�MW���$%�Y�Z�2��u�t���S���뿝��o���Y�l���0�i��TD�Zy%2� 8|w]jo���)��l�kp+]�>��%����I��2<0ϝ�=ǧ}aT�K�5���C�MT�W�fop����а�6!�`���͛���HEH$�R=.�U�^��:�'nv��J�#�.
�j��WƵ l�ω��,�	�/��5��V��)��r'q$ì/$�?;s�-/�b�ou_<Hf6��[��d|ί��u$�����gh��+~�,��;MUg4Ev΄�
������8a�]�_yk�X��V
��֔�I.t������?�|nu�ܕ2²��p�}1�b��4����&P�C��zR{���4X24�07G8�>���G�	��+a ��O,�8U�vc��T;�(�tj+W�	��e���jO�P��0���@9��C�J���x��i+D =��**�竀�w.��$�%B�G�P��H�����>�Ys�aQ�(�9Ч�iQ�P|�H�|��㜒��+&�+�.��𔖑�r��^~NhadI���q�0�ͪ�ӓ�f�+9�����5�.��p#�Ap@�'���,(MWT�#����{K�V�I����yF��rg��蠍7хvM}�:�DC��E�<�6ǳ=J��b5r�x����{��0է4�0I�q'F9�ٷe#��쾚��yJm�S�؛�� >���ϲK�l����4�9t�զM�N�s���i>F5�wk�+�t���d�c���T|���{�ӂ�7�Mh����-g�\ ݤͩ,G`��覆�o��o��:��E��;y���ڐ(���o�|�t�������*�Rf����_�ҐCe��W�O�r2�q�ϳ]�[bY�Y� �P
^S���j�"�+����{y�jO"�P��j�-��Tz�q��O�a,g�GG���� ��D������3�}$��d�Y��ZG�F�s+|���p�<,��##��/4���LE9���P�q"$)�+����fA�ݎ�׸��K3���K_3�m�WhH���Mv1�IL�~N����S^�+��ur��p?�*��B�Ca�R�`/���SrC���t��J�;i����UӸ�\�7a���'�1> xiO޿�@�5� ΔA]2�����Ǩ���ÀXl�prKt1!��(����9���?���/�:����%�	�y�93a�{�	@8�F�*���R7sc$��ѥ����x�e2dxe���׊�1K��Z(	��}���0�����I���F���D�w��^�:�P��x�+� )E�H *�7R��P�����C鏫b��?����їd�9���A=����g����&�+^��~�E��P�21Y�<ye�A�݃*3��0��}��"3��h������\)�s����aE���4c�9�ƾ:�	�+V��~��Rԕ� p����@�\�v����g,N�̵)m�V�I���
y�9�A/���`�62���̴�c�	�P�\��j��\�Ÿ��Z�sW@+��0z����V��Z�"������,�����>f��)Ï�R��4��p�����a|����-l�,K��踉�)y�0ۜ[�.�*����jZ���:��˒M!BV�Td�p���^K�h�%�Q�G��Z�����M��P���K� l�@��*��3;�Jנ��ݬ+�ّh0zWj3	`3�~����,��<L-�UHW�sW��!J�3��@^\w�`�(3~eͯP�;��'7���ײ6�����Pj�;���͕��?�d�*�M�c�T��C����CS�,��}J)=�!����S?��dF�5��Ń�W~+�n<IPϘ�[�I��-���n뭢w�N�ť���iUG<�dJolBƏ M���Jf��f�I���A%
h�~3��]p�57��[��;�ҏpr��j}�Fj���c�M�Hl[6�U9YTඉU�U7yKr靠��	�Pߢ��wx���0rk�yR�3Ȫ@S��Gڹ$`>(,����/ _&�mN�Y���,��zɳ����_�IC�����j��xש�Kt1
�60w��^&])����R�k�S1<�����ݑ=�-��`�i"|<�*� �znKJ^/�����t��h�Ӏc�J1�7�ܝˌM�CI��B,�_	_�:[ĉK?�ܘ
|0+�9V. ���{���p�Mbnr������57����Q!DVk�>fA���w����a��MۍZ�z�}4�r\������$��P?�]H� �E��G/�� =�1<1�;�����L�>�M�	 TJ��U��* ����C!�X�[A�=�C9S\��E���Ɠl��?��u�����DI��o�礌�,����)J��+�m��I����4/=���3�,�8�-�+�#s�|(��.K?��_�-�l�%z��Q�g�4g��=hed��t}��VC��dҬ��6�߫v�i~`^�r���FRnV�={�_�G�	7�y�n�^��<oe�����x!g�5A�A%�x�ZrD�k+��˕�(�� W��l�J̨�V��\lVJ1�-)9��a[����| ����jHP߁����[U�z���<{A�)3���OE%�ʨ����Ծ�n�[q��L� bxs$^�m6^���ʊ|�7����!�zWm����9�a��6f�!
�'�#a�{�}|�\J'{�7d�Cl'	�d
�E�%�!3����:\���
���z��7%��|��P���8����E�B>�����A�$ZW����{G�ҿ�w��u��dB��?}/���
�m�:ѡ�vuMA���ĉ��(i.���t�E�l�i7����3�*J׈S�[ޝ���"J�~Ť�P�g� ��eB4�#����TK��õ��(HbS�N�����S
�|���aq"����KV��S�5yFZ�ĭ@y�tɺ�TZ��{�nQ�c�)����pq m_$JR�S�����N'`�6�_��+�&F��B$a�a��O�F�
�%ή���YK�yڂ��ٌ���%��4R$���IS���6x�S�6��Lib��o��pş�s��y�D�x%�U�ԓ("7���i	�#���Ҟ�	�yn{4�f]�0��6�r��y%��T�{�+�����5��ŢVY�b����d�eE{�	����F^��
I��Yie��v6�1�3��8��q6c$����s��́=rx%�i��Qe���=2)L�Epbw��#�2ڻ#�eHʴ�ޡl�Io���G��#�t�(�T|�Se~5]"e�$z4V'�ז�{�X���pզ���&�����Z ��
�{�`������T� ����8�ii�����X�1�*cԱ�CO���� ������"6h��2weӲ�M����5s�{��� C�]�4�"Q�փx!��V��}K5Q�?�E�zM1���v�q��DG��v���;�H�������~�-��dM�==���'YQ�O߄�\���� ����ΛJk#a�MB���q�6�c�*kh��C����j;�dX�|��^vw���E}I|0o�?�݅%?_��0�����8T��c���t�q�������_�a/x{n)����)��
_=~��m4�{TgW_oyiɋ�%�Xw�*P��k�ZY��kճ�.bsR	�E���XtGPHQI���c|m�q�=��fn�|D5^h[z:*%#W����ᇮ��Ҥ�Xr� �7�T=)2��:Щr�/��,}��{cb
���@:?��z��%a� ����g�d49|��s�c��0b�ӏ~�g�g`k�<I4���D[�Ȩ�
8��y,{V�7:��Ğ�]����̫sբ���][�&��/��Σ�v�dŸq�4�$���A\k���o'��}���.��A7�7����ʟ��:>���tn��Bʋ��&^jj�� �C�[��MS0�o�}|�n��Ԧk��~�����f���EO��~�`�{�����Q���M�p�%)T.-�x�Rc(��Q��:�� 1����Ӌ�w�&�\\Č����^o@6Ǖ���U�]N��ܯ&�!���i�N1�d�K�yT鯧6��:]Vj����ߠlN=	��ӽܧ6r���2I}1C�©{w"<ݢ��M+?�$�>���5iimU����7� �H��A��-ű�&����g���_M�l�w׆E;�C��n9����w����X�K���z��0�KGŖD僁^s�Z�1; ʋ�-�j��=���1N�T�V���-�8��$v��G᩻	Y�s��[tl'�����+":E����R���X�f
¦�y+�_Y%��y�#�>���X�0\ s���L)��HEe�u~.�ܥ��F�Sꪾ<��@�S5�{����`��U sX�|�6�)���^��.Y�����D,�q�vԩI9&�=�*�:�e����e������c�D�v�m�0��}RB��q$��SUg���1}��fk2���ۯ��y����V��Nkܷ�(���p�=<]A������3�j9���c��饩:ʊD\A���탏*ԮY����#Ƕ:�+�EG�Q�]�N2��D�_p�[R�6�"��(�vQ{i�Y,_!V��6c?>tk��WD�o�zh&�S�?��N��E(�{2
o��wa�Y\���C��y��&�"������E����9�goy�}�>��-֢f�s�w'�$�r�����Lg�a�	�k=T%��f��zz���[�����~	�Cc��)/d']���T�h��f��U�m�Yɮ#�1V�����cW���Cdt�&W�M�Z�����L�,@����)	>�$�+֬Q�;�-I�n�ô Ad�jxR>�1�	��V�(�6�\t�ٻ[��x�G�GK忢��&P+��h?'��OmV8�fqm����߅�~��
��Z��sSr%��YE/A*nO\ET��=	]��6;5)p5���;ֈ��awbV����?gr3�!$9!�EQ�P�"��^2EZ&1/��o�z@��0�{ç|ʾ���,��A�Ύ�_�eѹt�d�J3g���^jw3���n���ɰ�J3z�on^�>awV�9�4>[�(o3�`O�d�=��Vɀ`bp	�� p\'	��f	?���'~��Gn��- Mr����F�|�n ���������fIr�[�~�1U�nl�o���i%��ҩ�b+���.��[�������6<n�_=�}-�
pƷ��IEqzӝ��KW�
,4��{���s6�桎We�t^�+8�{���Ϊ���?8��;�N UzJ��*�﹄vy��s�R��9?�X$j��2��1�rL�ѧD�k�s�����tօt\��e~"8��4�%���'F�A�ؙ �,"��C�)od�~Q�z�u�����iAx0���|�YN�!o�dD6ͬbr��L�����n�A�a=�R
<�
��<���V�!����ȑ�����Y�h��ֻLa\�c�j1��K�v!���%����(u� zܻ�R��$����nR�������f��F ����u�1Aah����y�:��pWt��o���,���,��Y��,��
����������3��a�;��ӗ��p��؁�z�7K�rE�3��xn�/�dn�$u�XG�?5n�ӟ��u��Td<eP�}� ��g���3d��E�ѫrj�g��#P\g
���;+U�F��ߩ�iT��J�w���v3�>Iɻ���m-��!r�Ä�8��#_�q�t��D�t`a8�"'Ĉ��N>��#gK�#��}��f�2�_��8D2�z��>ŧ�HO��8����Di͗�Jtg|m�@�|&�B�o����vO}PC��6��>��)�-�~n�i�G�����h�|�g��k:��� ��d	koC��t;�q� J�LK�����/}�o��Ud��I�~ɚp�v�ցr��0�]Cݛ��FAm���P8���ݢ�ɨ��`���)�B�E,�J�_m�$����+ӝ���fi5��BN�N8��֛,mG����$k�E�i�!T+G���[�vj�8٩W ���-֚05'��N��l�4a��(W�]=��x>����m��� �&̃�^���|��0��5(�����r�n�q=)��$5��d��'k�BU����ؾ>|)�%\�o�o�n�n?@�Q��B!I9��^�%������Q�ymst�F��美d�g9���
Pf�؟p#m���2�1Ddl0�h��zv1\y
gz�s�ؿRXi�aB�5�8p���{���K�4�\���!�]-�=�d;
�,�ŀp����P��5��}��-�֎�����'`�˃5D��)�JDi�MNA�Y�-r&>��dP��6P�}OF�!���>E����
4)�o�
�@ል7�=����Sa%	o�f�]�
�A��ǛCJ1��R$�kW��z�A��(v�<o�-x�p���'>ǌ��� ���<û�&#��9�������Zr�%����z�.l^�\��N���F6�t+�p�&�	y�
�l�E�ڃ�����۪1-͚
8:z���geGN|��0JL��B�����^f�1(���u�l�<��������{���@�u���K�ۂ�P�R
��b[D`���ߦr^��i�h�"2���4g�>&��iU�=p+��"� *2�2�:��ru���G�^���nl��q'={��&���b�#2���d/��;�4�.+E�p�b�<Np�a�������G��� ��d��Q�U�#<�O�cJ��6h$]z���V ���x�CU�t�0cg����~	�sd�q�֗Sf�8��9Q���Qr`��԰�&�3m����w�����@�S�چi��Y��^�����b����k�m����x����T��YP|JC�����(�N,����d�T	A[��	�߽��
+0�'�X�����_�����$��~�0�W�{�U�׀��˷}~[`�x���IBw�v5y�3q�'��G�	�U%g�7�z2���� �Jٵ>�4���g��-j�@�b#�U�n�����G�!ח�sY� S���D��"��3Nj�]� ZD1�v���`c�+���DM�]@{�^�.a��~�8	{�t_�!��H&2�L�d��Rd�l���_�A���}�����b��w�"H�r�Xe{�[b5���X��ђ�I>�z1ȼ/����``�J�f.����'��q�ZSP?#�c��t�AҶ�Ȁ��Z�n�u�c��2J,'$������F��Ul1���~� ��������Z�c@sVL��jF��� �0iYpS?�B�������Y��Ā�z�X"�M=��=S�����lj>{M��K1a��Ukv"�� ���x[F���xI�7S(p��Q�A@�������5j��'��v���~�+�9x�;'լo8� �����<	�-0��{=��XO�ԝ�G���x蘙�7,��^�`�z�j����,�����aj4 ����P.Λ8{�_KL�z���bɆl�Ze׾Z����WPܲs�#O{CڴgwG�w��MB(8�'�#-G�ƗH{�����0F���1͉��/�g�]��w5�YFha˻oѓcܕ"��m�}c�Jj�C�D�q.77C��dIf*���f��,�v�� M�>9�+�+x"�b�b��$54ӢN?A`*�n[��m�����`(�0nK{��cV�3��q0�/R���M�-�a�+��gx��C3$������h�n���U�p ��k���M�8� �P_����{d2������C�]�����)+��<r�Y^��s��rg���Y��r��,�w!�Ɠb�m�ٍ���8z?���\�K�1������8�E�_�h��/�o�ߨ�~�7x�l"j3���>Y9i$�ߵن��Mhol#Hݟ�9�;�nt|���'l:��r+���
�UEC�R�<u�SљӋfv;�+au
���v_t��xs�a�6��� ,{�å����AQMf���E�0U"e)N�=t� !�r��w�8�¦v�L��_D/�ti~�V�d�	�H�=�d��u�H�݅M����֑~7��J�2R� ���~D_�Np���OnM��^i�U[a\�z���~"<����|ʘy�u�O�Ma�>��Qi3��:��X�>�t"���#W���u�g@cX�a��ط��N1�������ۆ��No�!A9�k��vb��� �p���[ �fv�F.hWU�m}��ŗ� �=�)�J!�l���bkfk��x��B�Tv�(���Cw��~}��1k"��)7�4�"sƻ�Y`H��2tJ����� =ʙ\9U�N�}��� �ÿ�'Ѩ1�����av����%�I/*_&_$�풟SM5s������ޮ��=\����M�;c;Ijw��E���������竁�Q��%���=�nZz爬ywtPw����1�;
�b�9Z���[m� ��1�Hر�p ��ZgU�C�B u�G�ue�D���~`�����S�K��_B���{}�Q�A��t|Q633F�)�@٦��ZA�NJh?�����JvW��4S�ǔ���,���Nc|�����k�q`��snJ�	NwX{I�m�Ѡ�x����$)�qˀ(<�]!�T������:��8ذMK[���K�����������Ĕt�N�D�N�s�`�x|k�2�P���7�M#�a���=���F����<��&q��#�H�歇)�6=�`��=�ӯ��Rl�XyWȚ���h����$��=37+��@����&�N{��ĝ��׫琗�`�Յ�g8��_��Z!9�c���s�i�}%iҢ勼~c��Ƅ@��� -U1���!t�l�;�t�
�*b�O���A����0�ݧ?�,qZ���^�N?%�&����O3�/�6۠�3+X�4~ב~��R=	��G�z�O�
�t�݆O38<���_�y	5ŧ���Q-��;�&d��M��8z�q�.s�v$��"��m��Z�=��+�f)0��Ou�ѱN1�p޷� Z�C�4�	H���dWS�g�P�9���������*!a�����C��M����,�V�s�E7+�#\��W6�v���o� 2&�00��z�s��m6Y�VFod�>B0�e[͏�����_Jѥ�`��;o��\/�/2nDڣE9F�.�!���^K�WѼ����唫��{�Fp�J��:>m�8R��PL/��z����u�Q�1��\aU}{���Nh�ڼ�\�e��q7қus�`k_E��G���&�^�l��Ô�/��76%�C��q��e����>'����$`[8R]ǽ����M�Ex�e�����`��Òc�Ғ���VAeY*5� �M����d�l��� Hheb��n��K��)�Ք��v�Fh�ւ�2�=����R�]��R"��~P��v��%wvm��8��SV��u�Nݣ�s!��`ܲ@��3�{u䩞,/컞�������*�*��Z�5,�����k޽���5�r�)w_k�����^ӟ*��D�[`%��n3�������7A�6���C�|��c�^W?:ģ�E�)`
եf�Z!��\����F�+�����z֗��BzS=0h'-i%0�jD��Tc�Xf�l�n�\m{���_fhn=��t�������*����'�i4�:�W�����~���_��8�Q]}gà��o<F�F^�e���^�WnHџ�3��)��z0)#'C�T*.�J|�4�����4�̭�i$X�D��UM��*�[=�pC��S���T�'���"=IIB.$��j� �o��ݢ���h˛o'̕��� 4n kRV�D�!j^l;�4=w�V"�s�ŵ��)��wh�5So�1c�̱P�Ms�?�lv��� our�B��b�1F��J�\fn�[��LX���K����9^w9V�L�>�(�WE��4��x��'<]R��o$j�D��=L���M��W��M�
�)�!kSnݐx-�$d�ϝ�X��0���dc8�F�jPuz�T���%/F�ǯ�°�a�h��cAڑ���3�c�+3�ٓ���21H�=�Š�4D?�^���p"�fZ�F[W��hK������+�����dy'�6�3��:Mb^��2���`4�y����;�Ⱥ�kۏ����#/u�C�SP�B1S����Ɛ_3nv�L��k�ū�=�I�e�Ԩ�!��9w��m,���2O$l����=U�Z֍�ڞ=2��|g-��N�uʪ��&<f����H���X�]���L�iybR_xZQ����A�6z<��d���U3�7�78�
|6�uĞ��ɩlSUh�t���}~�e8R� �� �
S�o��>K��:�v�n"=4�+��pb4���]5A����+���i��\�Qd��`p�@I��ҟ�"l�{d���%��=��`����o��ކ�S�ƜC�.R<I
� ���iX��A��",�d���Cע�׃el��j�\�*sun������N�N{�̋�.�Y��R���}}����P��[=&Mg	fo����H�f��S�����h{<9�4~�*�iV*|�Hѹ��P��o����KOa���"��G�!mAt���d�,��1���/�$b��`�
�8�Dn�Y�a�S�{��"�0 �ˍo�P��Y�v�v�-��c��rn�s��Q{�pא����u���iq(�������T�U��F�3�N"���vX����؍�98��G���f�"79>�L�T�X�U��4�]z|�ˆ�H�w�y�������T��,�o��GOQ�P�,)Xl��=�J��1��u�m�R�� �k�=*S$CD�M�[�'���M�"`��
 �Ke���."|�h��R��f{�}gvW���,�`�zL|��f�̷�O��=���5Q�4��Q�9�)E�B)n1�TҠ�r��9�Q�7������`�"r���5%��$����ݿ#�	'&�Y� 6Y׉�o�m���z����F��Ѽ�.tʽ�e��q8M(���ˁ���%3�{m�u*q�wZw����Ȣ$[()��Q�SN����&ET���q�#R�Q��=�e�N�s|�F,%E�SJ��G^Z�L�Em,&�⧻�!���`�t���ԆM&z <Q�����-�����H}��l����:��@Q�xS������RV�J�W͂芲=]����~iA?�T[�h���)�L:2�>;�L����`?�����ю��U�j!F�i�b:+�{Y<��ugp9:K�M�z�*2�o��u�(xSP�x`|�"���	&i����U	}P�cro�HfXeh�<j����0;"]�Վq9�{a~@T~��N"��u�c�զ�i�\�n�h�����3��{����hq�viC�-�m���y�X�㥕Y:���K}B���)T�F�4��
4�'����XX�=D�nŭ�W�m��o�;;H"e�o�]�L)ã��2U�Ĭl)��O0V6%f�Fـ��	k�^����*X΄nzwcw��}��s{==�!1|��g�yɛ�Y�H��Q�ݍ��v�'Æ"�&"�])��'nm���I<<��<�Uަ�����4b�o�ϛ5��I��a<©���6�㪀���Y��ն�[Z�i�s����I��u�k�]�|d��J�f�9�6b�=s�	�AJ��]��b̨�4��)��0�r��v7!t���f�x�@�߱}���6�_�<g�͟���U2����ϓſ5P�	R!����[�ukw|@��ٳ#�u6�:j��q�M�;�I��R�5(�3�rqc�""?ېЊ8o4�bV�W۳I�VW����jM�,�Z��l,��:{+��2*\�����+Ͻ�b!���y2�ӽ&"�5���c���3���*�ǚ��֚}�?7>ޮ�.�+�x�Co_�q\�1�_��t�Y;�^&~� 6X��V=��K4C;��y���/���f�:b�0;��s�P3P�(w9�`y<i�j4�	��v���y�U�����8
/eN�Xֺؚd��B�`AS4�ND���&�0�����FU_��x̆����i4i:}1�Ο���7_��h4O+�UXu���7����@�Up�YS�a���-׀)�{"1�����ˏ�D�VB�:�f�-@0��1�'�.�8	�҆��"�qu������HkmpA�X|��VXK�0����l0�3����5K����ip��vi�A�o늳N�tE%�i��V9�Dw:j��2�J~Ďע�en� �*<Ҝ���	�p�1�&�st�����͟d��S�7܇򼾊We�<y���Df�5yj爍�z2&se�J�U�4q7y��Q[S��w�w>�,Y.2�d�p����:��OR�'f]}3��1��yO�{lPq'����^+k�&��u o��Ť	�"[}sG!�ʄ���v������(S����w����Ț���f�����v��<R�қ�b�*��\p��ײ�GAQ4��:�9�DR��r���8���b)�!X3�0?$�!
�����.��Q�dd��2�]�9?C�T���~8���e/vq��u�Њ��p�/X���.�\=.p/HI":�/u/���7���W-<+��+���m8O�d��L�1ż���7bBЂ��� �wo !C#Z�<���Դ>}j�r ߙ�Eu����ŵz�������1�U&p�.Qk����VX��r������P��{hy�1n$k�D�����@�����H���T���El.�5ݘ��ܕyЮO�#�!�t�u�&7�+=��F��Q���٧[��
�bqY,�G6��a�� ��go��&/+ � �"�W(bK,	= M��I\��}I��-�d��gt�!�Z��q�t�3e�D�Δ����enZ�� H�Xi �(�6Ih�0��{�Uo����JTmv"�v�"J�1�s�3�ʒ�����ж�φ�5����z�&����8l0�T�֯B@WiN��[�y2��48�$�C��6+@H�����%���~qu'�Xk�%
t3n��������@0��u3<��Y{ Bt��'O�dN		'X����RݒWT��O�_��DX� 6��?����`�| ��kZs�ᯀr�{��rt�d� :Χ�No)"�g~:J�F G���Y�����;&�	cSС����_�t�0�#�c�r��T	{�xG,;g7�����$�lȓ�93z����m4�deD�#�����AȤê�����/�!/�\�Da5���M!�_�+��G�*wT,�i/|z����V^)�d����*�T�g�01ݶp��tK��G޻4r��ɕOV��1�o��]�x�<ꁍӑ�����;S��Px�Hr�*̓2da��B���ݺ"ك��*�]]U� �)���>	8l���Q?�A#~�Q�{�9� x��#H|=�*ч�hS*�u�Bn�3j���@"	NI�G�5ζs�s+b"��ӆ������㖊�!�C�)�f�s��)�x�_[G�j.�*���s���y�H޽s�������3��Lq���rFT ��O��@�j��1lx�&��Ζ���n�#R|#��d�$�/�5��'�����:��ذJ�-i���LL���{q��+����$�"<c	m��������R]8'&A,T�2��@m/̙�aT_��e��K��kgueK���vRM�=����K[��#
ƥ�}��w�m��?��]6`c�.�=|��>#�d�*5%�,*0&���A�A¿2Y$;m��dE;t�A�O^"�E��H-Jp��4�v���C@t�?s��%07�? �"'K��)ayM��x�2���fWh	�����V\�wT�3�p�����1�ͬ���(�Oh��(��.I��_��;�0���.<Ȣ�T����\� 'L��&Q*ӦM�)�GRUpM�y1����)����
�t�TN@�}���>�lj�������1R)橄�c�"�6'Dfx�9E�f���AZ$�R'@���Shk�g�n�Al�k^�����n�[��>�r��P�ӧ�������~ro-����!֠'��v�5��#??H=>O�O#�}�����OR3#�_Ԝ܎��{��oi�|lJ�dVh�rZ�����z������Ͳ#V�E�+�WG�w��e~�F5�g��n�3� ��'�`�ʲ%O�g
��(����hO��
��=�3��OB/h�U䔰t����4�>�e�}	�@�.D�l��������X$A>mD��q/����a��1ZABLI�h�,���c�[��(Yٕc�4�Ί�z���BT��
E)
ϕ'�f����4OQ��n��Lf%L �����r쥿-��{�e��P�.��L<0��"��$�n� &�9�dz���B�.Y��ȱ�S��'s��$0 �ߦ��%�#��Z����t�8<vn���}��i�����DM�$�)��n_����H�
"H@�DҒm�FCպ�����4�@�B:aL��{���h$S��ر�\�z�u�B�%f���V����:��e����]r�@X�ZN�z��
}��Y�����4s:bю��Кa߾�K���]]㷿�7H�lT�]2��"�S��f�Rp�6-���x)ܝHJ9>����ǡ�M�M��JT��:p�X$�~����;�Y�+zhL6�Xa�vP����Vǉ>!�i��&����:��I
@��ڌxC2P;�ޅ�6别EE�)='�����ǆ��/�����r�����
�L�E�2�����µ-�F<�$E���,o�C\A�����$��ܦmZ���' ?
�s��L�R��v3���(�����|�\�h�~v�M�p�>Ϧb ��/��P��vƙ90R�p^~�儼R L�YX��!/K���տ����eѲ�n�$o�*`WҞ���W-qy�x�m�W�$G��-DB}�c�t]�m'�`�s*V���V&#�5�����x��"�j$�5��4В�P����@q�|����ŀQ4|W�pϩ�IM�8�qE�{������0gŉ^Lc/�)����߉U�,��/$j���D�+hf-&�|�:��(��^0Ha3�O�'��=��;m�]���O	1 '��\8��^��.Ŭ���z7���qd���3�C^������[T��0&�|��k8����(��J��V��H��2&i��C�j��E���:�U�v�o3��XsdA��j��8�`�?��݇�U` ˁlh3�*�2K4��3����]��*W��������E����R�cZ`��oM"��)A B��}�l���uzk���q�b�]�d�/���̸/+c�Q�H[�	>�X����6�.Ґ�I�����C�9�^^��&���O��N!�Ep}�{��O�Hb�Vz��"_[��>a$�v�i��AV���-1%��^`SMm��巑sW��؊3���H4]iN��w��D�Mut`@�;-��������{�T��絁��_D���3p�8��=4�Ԇ���9��Z������$Ճ+��a��`N��I��tx/@s��q!�� ���L���pC�Q�K��_��A�����n��[kSUN��I�a��[���q�&�C�He��8�dg HlG�����ɧAX k�C4r��b���`@�=v͙Q�#TkM<s��,X!GĜWYZ�@r�~��C$L��K�#}I�;C���J�� ���7%���Tb!+�EA�(����+)#��ɖ=���U���D8�PIoj'�\���4�l��7}:�*C%��4��ͱj[憳��׼M��.q���s2���hdǛ{[è�9����D���0g�S�~WQE;-P��+�J���P�DhSR9@cz�l }�hZ׺�- �Ǘ��_�qp1���'oU�j����s�E{+���'�0K̋��[w����}ŗ�B�puZWvCn��J4�=��~���l�?L�7-���ӛ�bc���9TI��_i�4�R0��>��zc̐U�o��JO��͝e���୵Й�)�� �cH�V���Ė=�B�ǣ%���1�(cI�4�?���>��$�Ҿp�.)������Eq���_�G�Jv����rR��6�a�kn�2��m��n��[�u$�����Z���	F��k"r��{��P�m�.�D�֏iN:=-w�ߞ���B�NJ���r��)�bM�:T��(�'���FΫ Ið�?�Eb���bͯ�Д	7��{T�-�ޤ��GG��4y�.@C-��/�q���'�u�f"��l�1��ED�ң_����t���z
T�L��N�J�'͜c�pR&��)m�z�7�ܥ��c>f����7�bZ�+jk�ᙦ+��{z�$���9�<n(�b�\�J�L���NQ�vi�i��o�l��E���������2�h��ܢ<���K�%JPW��p��� ��{�{it�f�O�^NK�T���i4[���\(J�g��̈́Boj�"��̂Ұ�����%�)t�����[���_mG�7�]̮���zR~]�u�&�Í�)�#�4�W�)�R%�w7F�O�z�tY؝�]t}W\q\/Ӗ�+��60�.�W�%)��5�#ϫUr�aZuk���ٍ���i�2�J��h� 7�Օv]�뭋7�&I#Q0!�'l�Q�O��D|�lVt����'���η��V��z%ݻ\���A����2��5Df� g�T�Ĵ�|�Әv�k�¹�����t�28���7
��F�p�R*��k.�Ɵ�r�l��?m�%�WS{�� �G�|F�N��������MTDnٹ���,Z}�;�&�;�W���J�Sf7�j��IO�iw;W�l�9(�����@�������9�O��Y���q1�F}����%��L����>e	9��6TS��S��	�kŽ��� mʸ������
)@��\�A��_3�K�hK���ׄ��B=��t��io�kzu�Y��$O�tRl�ģ����c%(�iyD=��s�#�u%��w��0��g4���e���D|��p+<�ۻ�Qk-�\
	�u�`��� v�X&"kپ�L�q~��DR���<��q�歒�M	LiZ��������*&W�_h^���&�$�~����x�M(�����f�lw^��]4�*�ތx0e����Y�;�'3������1"s2�����9�������$C�����o	�K�ה�T���%�1��!Ad��*�^Lx��1��W�j�ǌF%���ܥ�ޏ�~.�$𼡈]���"i�Z��X��#��,�ԝk�s��Yn�S���I��\�v-�{Hf����ޥ���ݽ�1��@fq4�}#�*lY(@o5��w�
E8�t}O�tMk�E8lr���V�|X!�N�7����:ӷ������s���MS��v���?�/!��4���p��$��Eb8��n�������=�R��qy���CI�#�]�=<����ݬ��.
�����S�p��*~K3<�i�Q[�bt����ƃL����V��5�(�K%U��08�����Щa�� x8�f㾾?d���'<l	�@b���:g?�盠҄�� iJ�a㸀x l4�P�_o.
S���c��@O�er��1�H��rF-��E�e�Ӷ ios����<yՍ�W@�<EVQ��pF�}gG�;�f= J���f�4?�(3�^� l�z �5h���K-f����A���z�O�y�E��֥7
�T����ذEmЉ4�*4I�f�İˉ#;�"�0qJ�"!�b�����X�<@������$��˿���� /�0/w�	T�����������L�U�������D��"u��]�D-���Aq��Q76^P�����68�|��!/�1�0@�9�/��ֶ�㺬����f�
 P{b�?�����=�ځN��u���.�0���=W�j����D���n�k0��i�w�Dm�m-,��#l����%^Aѝ��#IC�b��I���1.ӳ=NSo�W ��P\��COP�������@���-k�x�Dc��\J���-B��(�7��e���V��G#�*�hVT��>`�#<��e����|����Z��D[��0�s5�#�:�b�,˶3��ߡ��qt�Ɍ،as�y�s�;|>R�I8P�����~��������*���/8��˶�?���j�*�(�%�8�`�hܘ���0��':Ae+��o�gh������H��%�T��)��{T�u���K��.���N���n��JYAq��:{�d�#k����b�rQZ�����]@�b�u&�z�Z|�`��??��c�S�c�0 A$�+lԤ��FkOKKC1X�n�-x|���p:.���X'�(r��# �.?��n7P0c&�Z��}*Ȝt���1G��le�������)�҂��i���2:|�oTD8�$舭1�W}�9 ��5-I��뫺�Hf���T� p�:��G-�t�� 4CE����j��7s(Ec��I�@� J'�>��<=H���F�yNM��vg�yo)=7�=FPa��G���g߼�{���Ks��9p#2�� ���D���K��E?5q�����F�E���B�1�����dӠ8��d��5��q&s�;sp���+��K�`"`��;�B�3�N �z��a���f�/�fQJX��;P,�K���ó0�.��c�3M���b#�����4�T"iWT`���ɧ��Д��r�l)y.q7�&�{�Z�<���:C[��tr����&3EB�<3���F�z�J��%��99NԊ��خ��"�u�L��zdEX���D岾���hm�9�uD�K������<(���t��&iL��[�7�{���:9;�:S	ȿI10��Lкp(�*f�p�b;�]VG�k;�ǢE	g�C��.m;9� Lz%��a,� �n`Z��/�Y1�^c݉�R8Ͱ��`G���&QI�-G�r�
���udqb�R�Pz_d/�lp�c�~S� ݇�w�M����ǉ�^!���\h3��1��D��C�]u^s�R �0}p�b#��?�Ԏ�1Lb'`pf!Gc]RZ�+?�^΋u�W@�Q[A���"eA�HJ��Եl��dCr�&�(������Xܰe�5Qb\��]��O�	7u�9�ȭ�5=O��u'
b*Ns:��*�GN9�b���J�-F�N���ؠ_��g,��wx�c� ���k�J碠�=,�oǐ���vH(.�hm֬?�-���޺�p�f�3�c ���E�H��T�T��xQ�:�"�[, �3@㐠W����BA`� �����'c��	=��9h��}��&��3�(@O�ls�}pp"RCs��'H�X�����T��*��$�܅�o����!�m�¡�%��ũQ�5��~�6���:�w�(�D�޴��Җ�f������H Ŷ_[�Q�;ԫ��������6{9,�&�i2m[
��|��b�Q��!�f��X��I��>�>�.��l����_��\��g�8
�Җ�
��C��g�~��z��4&3^�Tu6B�9�����Y�@4)\)��v"	{�;FT��e�/��`6A	T��Pϕ0���O�ua+�m��1q�guSeG�jt���HU�к�V�x�����;�K��L�_6�:[�0��x9��/zͱVwf���O�-���7xJ�Ϋ4�6�[T��|aE�U`�ܝ!�ɳ��&���`�ق岓l�-��4Hg����� �k�Ǌ2�����
T<eu6�G�v�����WBeRh��N?�ˆ Z^�Aˮ� g$r2x��-n������W-[Su�N��c�V�w�ʊ֒";ѵZ��ދx��l��"���� �[׀��ݫI`]4j���=��`Q����.�țX=ow:;�r�m���H�K�h����b0t���ng�fl�7Wo~�S@j�,�o���IlkܼϺ��Pt4�5ȧ]�$"�x�b��Ltϧ�JW|�Z��T�nD��*�+#$o�����ŗ�`m�j9��;�F�ɂ��d�݌���J��Q��M̑4�������C-�#�K�g�����d�o����/�H�8�õmH�(K��|�Ʒ�����_w� I�(D}2W�L�4O6��i���T����w�G�&IU�$\Д��j!Ì}c�sGk��k��s��Qi�<�����j��BmW��*�j�c���-4�Ͻ�k�7��5~�0m�BS�崟0�p'��HT^����2�A���{�g�R2f���˰���`@Q4�WN$���ha�4���0�&G{����nj�kG/$�Gg�����_��}8�TNd�����<�K��*���j��5�y����=�:�r������������w�؝����k*/�u�Qʃ�|�a.�r4�EPz���)�j?�3r�P�|��#^����&�/p�h*���6a���%q�W�*5^ϐ"#�E[���%G��|!�3�PM
���zD�}_(����c���h8<
�]:�J��S����-ȸ+9�+1���8�guO�"�"aC-Q�C=��^F4��Jx�qQ�"h��I��J �v�C��9�E���^���ȪL��Q:���^�*���9�N�<9[�4]�0�F�}�(������)0Bѻ���k�:(��&s�p<�Z�hz�N���,��f��k����_���~���N�u�l�?�e�J)�A����n�4�b4�i-а ��	���u�8�@bIc���B��1{Ʊ?2��|<گ'I���_����l������P �ïSfpꋎ��Q��#�8�JJ}Ax[Df�j���3��
o��z��_�$C��C�E����\}Ǧ]�"���L2�p�D���y{.+Ȕ�2jxk�d:���Qr��Q}<c
�g��<��s
1^/��+'[�Y<
EZq#J�9�����<����%qع&�
���<�鸞=Iє$��*v�;o�y��E'�UV�z�F	���U�e�X����H	�"�
���ǉYe@[���6�@ o�fC���o�s@��/��ڏp�BbW�4?�ح׎�QP;�A�%�yZ�E�x��l��`���9�f� dI����9��WE����Y&�y�^6�o�&c2��yĺ�PRyq�x���r`�826�}v������hY���,�H)�:W��3�x�C�f���0�Q+�U2��&����š�yV��{�z��\���R�j@L�c-q�??FZ���ӴKp(^ J�>ƃN����N��8ߘ0�J:�4�)�	?�+��0���=�,1��'.Y�;�4�����R��p*��Ww��VCW�H3�7�q���`*lk���/r�ݽ�J|ۀ�,Ҫ�:��{c0+E�7��1 ߜ$�?V�,i*|�M<]�?ʹ`&��7mHe���
�FH	
7�<lI�A���{ŷtAi4�A�=-	5M�j�>�2��v(R���Z�9%Fu�*�SL#ꈼ�p!�Bt��cϯ�g�9�#i~67,�`���Z.��&j%˿��=Z
%w�b��D/����zo�z���j�~Y��0�]��e��l�k	f��O���ߋy~�*.u��&�&?
pR.XbJ9I����yj�8�^�^ˇ���j֗��~$J`�����W�r-f����Z�~l ���$/:V2�'�S��23�*���؏�ҫhaTo�pe���z��+�aMn���������I��p^�It��+�rmax���#+\Wrx��N>������[�K�W��L�=�!jIǲ��ófdv�/'���'a��D�S�:p��Y�t����8��rT�K3�l>�fv�%��1�m�	����T�����\A�<��(Y���=��T&�b�$<���Ա��?�������Vf#ښ�g�&1T	Q/RxC5R��?�f�������Z�L��%<�k�1W��R�MZ>�1��fgUGЃ%P�bZ�6���J/2��\Y�0ri���x���k�S��]�
�q���_r�u����\�	#���ϕ��E�81�{65�!^�O��!�yڿ����1��N'�ê��mU��փ�?���'��U�s��)��o��� �(����J�Fc���'����M�pnp�/�-D<i�fz8��Ȩ�k4���T�����1>z���*����^��M"̂u����!}F��^"SM�۩3C�����5��&���^��+�氜�y�p�|���g.��D>UZJ�����L8+��#p���|h0�D����dr���j?nR"E�4(��s1C]��t>��sVȤ��_s,�R3:q$�=��
�����t�Xp���$H `��b�Է�v��4D��*Z���v��Q��:�$�����3>���� ��(O�7�}`��Vfs��A�*�ُ��Պˮ�w����}
��ຫ�!���B&i���h�pI�"~��Y���^��_��U��%
4� ;G�([aB���_i��'�]L�����Ś��S���7I�Y���(kL����ʎ	uP�Q/�
^|�)ԁ���7�"ۼ3�6y�\�t��Q �Mr��a�b펍�v��D~K��ϕ��1.��z�&!v��R��2w�;Au�M[w@���]Fl��c������!�]+V��H���e��:[��F2@|��	I��ǈ��d`	$�T�ܻ��_>����ű_��;�t3�����y2�=kҳ*���j!y��9]����ڊ������ُ|�	�Q�2���yn�F�����U�'g�ӻ���,�U��8{�����b2�euL��܏EL�#�e�Nr�u��eW�g�`~�	98��5�?��3tr�v�yQ�
�3 ���cu`������l��9mW��Y��j�rإy�Vp:�����8֫�O�l?�PE֜єK�d�%�	�}�	�,�y���}TC�tz�.ȥ����Ok�����?�9�������'>��Q�7�0g�z�ƲXX��M���{��-���54Q1z9��dI�\h��_�d��&2M>'Bj�of���3��Joq\�ʓ6�h����؎z2A��n� �6޿�t�|<���]1��B�|8�t�\���^��CHy����3�{}�Zd�Ee"nC$��Q*����P�KMn��2�n��nӀ~�@`VA�ze�n�`���@��A��p�؃�OOXϑ��0Ź0(S0ꇵŭO<�j�f~C���C�m�"\H��ru��Ő��qb6�ԋ��d9�<������E>����I�$��6-��I/�w?����pM�E��@ Yib��Y�q��\
}��u%�Y�R�Ҟ$��2���t�ψW�P�~�����|�y]u� 廜 �U ��+O*��R�^#�z�)W�U�s�=B�g3�#��1j�����>����Ѷ�$(�������^UYl`��<��(0��t����cC�{���B�*�y�7�t��H����h�����q��d%n�����'���޾q���av@�6h�EmbA�/_&�0J���;b��yg�e� ����UXs�Ź��k]d _�dn�|@���?w�1DȦ���� �(�BHJ�ǯ1�4�۝9��=��[���]������F�w$�x�:w�m�ʩ�x|�g�`+�A��/P�7���jCzn�$�8֥+��ǽQߒ�s#��g~4a���$�Q^{a�ZhZ�b�N����;1�E�p��_$&V���G���p�l�(�����?��,���sVC�x����D^�Qb��_9h�\юi��K��O��Js�ao�&O��X8&��ܺUg,��ȯ�:�4Z�����}+�nI����~�{��������彼2�>�g9������외_ O8�P_��SV��8@.=�@���I�h��'$��:��Dg/�����J�x��OMf�,��iX�6#i�v�����8��9�^a�퍽I��Ҙ7����9|������2�3���KnYV�k�
b=��;�`]���lXkڿ� ���"�p�v>L��R���S�r�D~Z���(��;�o������A&O�LH��TCd�UJ\w���7�����o�#�X_<(�r��.���?��g���[�����`9&�����x3�`8J�[�v[@W���������(�G�6T�nn.!��=<:��8�8K�����3Em�@�u���E&p%*D&u3A�;�q��ބ�FС&���:_�
v����yC�w�	@���e	�G��h<A���o���VG)-���x���wNsW��C� SOžjז���WV���򸳥=����D�X�Y{�O�7@��cȡL�c�)Vb�P����!��Ib �������$:=�tk��g�̿K��W���	5��[Q���Qr�@�βX�vBg�[A�:3�J�Sn}T
���w���Z��'������P��)�ބ�	��a�&CWfaL�O�XA$m���L��O��r�A�����n�ȿ�	I2X���Kƒk�R�Xuz� [3t��#�t�Q{��,�W{4��ِ��PS�	j�g����>õ��nB�p��8���9�>P�C/�b�H�QU��n�ͭ/ѫ��?��M(��e�u��(%�̝W�R_B���r�&Yy�(�0qn��
_��/�u��R�g���䫾YNbu��I�u��Dik ��(X�"[�Q��BB���(�>�wl}����.�ŧ��z� �DY.�s5C,z�����Pfn,�$�6�\m�V)2<l)�߱aRc�ݱ��Q��m>n��u��w%�е���6�t����v#��#�m��
��2��{Ɂ���Ѡ�Q�?�,?�lΨX�G��(�q6�\��h�0Sq�o�W�T�8�h-g{ē��w�s�������1n��/��Qnތ�:os�,;~�S��o���*�dj]
��v��\��H�9�	�^���E���L9osK��Г:��p�rNr�F���>�-Fs�4��0���N��-Sڋ�p619P
��h����B� ��#ն�����k4�4$��y����d-*Br���G�A]0��_0��l��}�S��1ȝ���A����d$�F�5i�!�J�>���D��
zE�EL��p�˺4"�����G2���!�7�X���a�#)1;�M���k�d�;��=Xi0uD.i��>�dE�vܠ�����6���v��úHG!�у� ���+�˦�����[r�C~�����sX��o*䜾X�Rh�����[uv?X�"t��JN�X0�B����2��t.N�m>���fW�B�B��+<㦸��3s���,�JY�YBEJX�!�o�w9�K̽��Io�\o���������6i���>���`�+��m�E�����0��}�i�mO[V{�5�}�S��O���ї�-��7�K�(�|��j�d�<	�P�e^ޠ��zC+�y5��� �;��%C��נ�м�ħA��5z�š6����Pd�G1v>8�iӃ�p��|rj�ƅ>��Q��üՋޚo#��� ֔e�)���j*S�+��T	/ߤ)F��S��5�F�����'�'�H��ϑt�vc���e~.�w��*��8ʶ�ѿ/�/Wͳ��((�+lf߹xнj%���1g%�F�i�����߸T!�Gr �C*��L�k(�.��V�B��/A�%KpM�I4��`���	5�"]�^u�����������`����_+�e���p2��R�T(R!I�K�o[\�H���p��(wE,��h�=��j���k�[���*���#7f�`�Km�R3]��^��X*ܬ�-l�:W"l��q��^��;a���Z:V�gḣ��C��S_:r�F��� W��!��3�W����%ښ&D�*p�¼���&a��{�����Ȥ��--�- ��⧨����t���f�ֳq2P#PC��f�����،!�&��CM�4��NM�;\FV�$v�	l�|����Q]M�k~N��.3�1�,���jmAE�?�g�-&g�S��ko�����?��,��ρ$5�w��ڌ�1�������?L��������o���h����	0qZvb�i�n��_��Є���C���x�~o��!uՀ��̉!�K���Ů��j���Ň��Bw:~���d-��ڥ�㊋��14�,�o��1ð+���3���>_*�<j�O鼇�&k�/r��% .��Py���Eoo����������Q�u��w�?VCj����>O�b|q�[޾��PvGJ���IP��C�p ;ٓ����5&�
_H-x�|���٪�&V
��q�"3���r���UmNu�Qk�G�C���}�3�u�	FљP*�Y������cǀ��{�<������A۾��d�p��	����x��kG��DV1n"�!��R���N�����|���f�S����/�u�:>pC��[K���3S�7�G\��K*N�,_��љU&�/�"�&eo.|�:O LB^���t�������=V�g!���'b��j2��r��*ǵ>f}� �tB9��΋���p� �2s����_�`$J�8�S*�\�&[�$Xҭ���I&N{XC1+��g ��r��������&|�"d�*>�a��D�C��nf��= o�I�R��Cr7��>Q�����<6j��g�Q�<�A�R^_�$��|�,��{��� ^M�%��W@ l���%*�k�9a�Ą΋�M�O{D��c2�;��E^�i��c_�b��*(�m�\p��Sl2V���~�y9�m����8��(�n)�O�fZLq�7���	|�-7��� ��y�imnr�\$a��E���wUڎ)_�HZ�3�C܌I� OfGMI���Mθ�L�%��`C!���)y�ge9��F��q��� M9��;ͨbz��F���?뀖K��$ ͆����t�����ׂO痼l���א3@^�VΆE�|���d����"��w;s]گ@�����t����";�b-&����O� �Fx��Z+r��Ib��OΏAʝf�[�\��5J.�:ħB�mT`��;HT�ej���5�-�O�����gi?�F㐠���(�:����	5��a#��\��o���8ֺeV��پ9��o�~��d�n(�vZ5_��0m���6Q�i��۞�^b��:�0J����G��� )5����J?ͻ���V٪��A���E�Ts�>�߉9�����H2�Į>*'�ѿjC2u%�;
t�r��3��n��\7����U�D� �84�ZTe_g�tW6����x���]��C�ݗM�Elp���:s��ZC�K�$S�.A�qc ��1m-��wjU}���@��U�l�J��&���k���c��\�?X*��6#�bHl%����T%;��:����kڼG��ch�﹭C]�Hz������a��0�°{*7�i/k럑��Ĉ�űg���+�Ä�5�֖f<K3�.ff�qGf(?��U&���}�=^�� ���d���A*w.=�d�KN|��E%�������	�V:���_�B[zkT �<�]���71��m��[G�eS���uZ��_q�ǚC���b|+�+���~�pe����9���)5�Ǚ~�3�Q�Qi�l���C3����>�d����_��esY�N$̎ QŹ#���WAA�g�藘_s[(�b����}8X�Z�"��˰X��gO��o����X�O�|��~�͢� C��7J0��C������f)�gk&�q�8?+�o�bP5�����g�M!J�q#�=H�/���5��]��(��vՔ��r����7M��H`of�\���ZqeW����S��i]`�#c�z4숊��ԹA��qHz��I�kԍ��5�×�u��N��n�~�Ũ�:4g*ϊS�-���Z&�q^1��Ʃ��8|�qbxb
6��縚ṃ� �(��8{�h��.3h�;��O"q+��{��:H
E}/	cv[>	�_n���=�G���O}��\�Y�S���mǫc�M"�V��J�n)@J$lq��S{S��Td�kJ�U��]�Y���xK8��V�ʗ��tv�Ӵ��؜��x�)���g8��� ���%Ov�_<+����́.3l!�v��,� %'�'y=�M��t �qN����/�2Т1��Z�	�=��};r�r'w��$y����j�Ӄ0O��'66v�N4���Q��
�d���I��tjy��XPJ�� ��\��D���-e���k*l�Y�������v��xmrl�Ą�!+�f"��a���f3z��]��L��Q~�$g�3,�/��W�'Ez�@������ʵ����4�2�Q�l-%����As�U�	���QF�"|	Һ�!.R���K12��)L��D����j%NTF���_F��Z��3���mIo9��$P��0�����������x)�(ڳ >��w����9��/S�R1�'��L�I,X�4{-�>t��컻*M�R]�#�f'�an���$L���}�C�����Ɲ_5!'��e��B��O͆��+u���5��W�]�pr~�6�����e���~��$4���	�q-�8�ib��v!c7��#'G����5�!a4�UI^E Tf����a��PȞ�6��V�ˉ/�����"����OF.�ޫA�;�I�K���j�A�6���g6���rT>˸X�b���o��0�}t�,�Ɏ�>��<�����l&�O(���'�$<6*/�r>Ͷ�^��s����]�8f1�N�D�0�n���iv�4��3��3����)"5宽t�O-��֢�5��T0��2��dWzy�6T*kܘl��T�P��o2�����{��]�u�_��`���� �T�9�=��դ�RIHv��UT �ΗrQI>-��N����ae���ˤ���O�V�˹^��K3��b������YB�+��,hx�k\�L2,w7��I>`"��,�S�[m��3e}��1�_�X{+̠�߿��=ᢉo8������,r*�"˞5���B����ehUp �cp�9F#�9� 4_u�<��SA��:{��͕$���
���k��G��6S���l��Pr�����0��k�PvF]�P4t�t�;8˿�1�FRӍ���87��X���3�jcW2U�d4r�=O�!�wGcQ��0	Z!R��[ûx���r��9)�؞$�<3P�F��ĕF_P�[C-=�_����A� �����c!�!N��2�a�9'N*�`�cZ�V�VMqt��>�5ZZ�#���νڠ����y|��~�"�\O6�����Hr��m�ϐ7(�J�߷��f�Hwb���bI��+����>�H�ʺ��� G�^+ȹ	��Rl���=�쁗������,Qm_k�Cm*'C�9�)�I#�K�`�����������o��Q��DRGҀ�Kx �I�P c����V"�r�E�c��?�t��ՠ�ϐMf�蓦T1�V̇��L���%���8J����e@c8qo�W�)��� Է�$G�ȱ�>Ư�glw��Y���Wd>Tp����w!�b���n沵%��Z���1�P��CG�<(8�5_����F�3ehv(�2�z^&��� ��ab���]��hl{/Z�����TZ���}�-Í�O;������g�'�h�C���(u��ѯ�����=ʕ4�Vfu�Qc$�sQ`��e��\%@�7�l�+���|�k"B��M��:X�~>MS5��n_Z+���7O�k�mV9�?ԉ�w$A�[��	�U�߀g�-�~�P>XM�- жāf��)� n�K�f�o�-σ��xmz������uKm����@��K�C��;[ŭ<��bvӖ=��*�og6��C�4f��5U������^�ٓ}��s���K���^�gY�I�%ޮ�Z6�xA��_��K��s&�H�¤ v��2k	B�}'s��I@k[�"�H�~���:Q�v���L�ń��w*^I����g���]FԈ�[�j��};Ty��ۧ����ǂ)cB����A�1�)���akˋe\�Û�#��ܳ�� �]RD�4j�#��!I�y{
!c��գ����
n6�[���'=��Cd��v7
0���l:�R|��km����\[Ppu�UP�q�;.��|{"�JQ~w�
$/å6s�S�$�ȋѶ� Ox���M����Va� ������^�lk3���l��2"��܉�q�uU8Y��9�FTy�0J�a��_12�h~�@H+�nr���z�������Xْ#V_�}7&Gx��A�\�ť���x��9(�c^�X���Y�<�(#��(�����b�����n�?���[`JX`Fw�M� �������b�0Z��{o��-��?��t��%j�D1�l�����Oi�gu'�UOVBD�"P��I"�W�Ԃ5��Fϻb�f1Ӝ�W�wwcv��g��;�y�[��Gxx�Y�IL�	W�nhY�A[ㆧy៧��{���׻�f}c{����<y�����*�[t ��.Ռ%v���>ϝ��U'�˲0�EӲg�8w�ZZ�U�����Zg+_�`�u��Λ��g��<����f��<��|@���xm�oL#3�Z�D�Ս ��
�f�B9�;�@DǷj�IQ��D$�]�]ހ��y$�b�h��X�ƙ��7���`����]9���C������ܝW${U������(�<']�%��k�b/Eϼ���-c��}�M���1�V(I��8ft\Ib�Љ=`�a[�ECS<����H�1c�F�.\ı����W�+�>`6�N�)Y�,��Qc� ��:�î�����9;�g��	vM���M��fn��l��_r��E9&��YxA�1�*�Օ�I�����M-�>ŋ���4MM�!�#Zq�@5s.t����{�K���)�D*���������f��ᖾJ��92�Wq�&�X�F�{	������K��9�������Nꋼ'��x��&vvh�z/�O����t@
�H��L���x���k�8\����m%&���g��"	��e�UM�E���u�sK�L��
�M�̖�CKl6���P����M��;#V2U��P�Aaͽ��2�XI�TK��R@yS�$��Ya��nB��V&\oK��$P�Y�	Ԛ�)iV�['����3I�SQZ�IH�#���2���L��1�cH�B.��m�A9�ǃ��u.�J�cC��S�d �up���Q;̫��ݝ��`q�l�`����?1��%�d�6�E���ҁ�T���[G�i��!�O�ѝz�����]���,��̃Q�B!�+�OJ9`�ׄ�R��N�[)�Kơ��O͡e�*s9n�% 
l�S�j֡�M�4��h�q8uq�]�f9�p���4'衭�-*��,j��7�G���ԫ7֜!p- Q,nIL�?J���s��&cǴ��[��F�*�n뛕��3	��������t�����q@lx�	���*$P	U�!�h�� ,k.���<�e���b�{���(]>�RH%@����a|��|H� S;�`z����b�����i��j@��#�l�)ܛ\.\�0="b���`�m�ɐ3eck�{�|�Ë���<+�0���F��T���}Q�i�ri�j��磓���Ek�Ci�[��2�#u�J�*Q���M�k.�K}Ľ�/�xo!`���@�C����<"d����Lj��_#�ݙ�vQNy�}�۴$Pr|}Σ�����ҟ@���jde��!�B�+2T����y?G�̓9�;G���^bv, =��Fk#.��?[C�?��iE���_|\����Շ��A��z�O9�=j��dz 
dC���V"�rBx�)	�6�%�G1�^`��,�V��X|����d%XYB)8t���1��A1�g���K)������P_���?�!~���(�%)�"�*�Y^������ _ȍ]��V�i��:�֧}E�����=���W:��
BN�#��.22���!:cw�k܎�O��'��|���o�W�<�e|~� �����#:������)���C~Ic�[p�ںHq�������Qb�.J,�5���"�bʴ�<�-?��mU/�K�LCzp���}��[��2�:�W��g.����vс��%��VFT0!RǶ�_�w1���Ō�2W�AT��wY�B/F�W�M䋷+���ѰJ��*�����͂r��G�a��rQeK4��iy��
��q�U5qI���b�<\�sA�k���O�JN��F80���|s$�PX��kR��~GnT4�fM���@۴��>�7 >����O��U=LM�&q*���(e@v &W�hZb��A�c� Y�8�b��G���� Ry�c��%Y��r-�n���Q�&��]M����9S!�t��Odc�V�Ċ�ap!Q0��xQ��ӆl�� q��Z��>���q��OW�&R!�s��29-��~b�q��"�L��!��}a�V��S���a|��m�ڰk1N]ϼ��>g9�={�s[^+�
{nV�1t+�+Z�LP(��6���]��ݿM?�r3,С�:��ٛ	fk�E�l϶Hl�iSo�0�n�����F-��]��lBIdߖ�f�1��	&�ۮ}RY,��SA`G���r|�wU'�}aS,bY��hr��z��rzv��,+��T ���DJ�D��t��W&t�d}�e��Ɨp��5�(���;.�����X2/�RI?cr&׮��e}f����Ba�U��=YcT��vބ8�z��8��� �&X!Z���2�׿�w.h���!Vk����xU\4���3����b
�)���ko�7X3+ڞ{�OR���tu93M�t�i�=������y�ɶPpp�H�ʞ�{�Կ7��������e;J���G	�ES�嫢U���0�Д��~_���p7FC}���
���H��q[��a�����-:����D;(V��?]���\A-������er!FG��9.D�Q"ɲ���TFY����)a��s�c%���7�*��z���P�@肯A��[�{~�)�X`,�R\b�z�g8�xpM�GVޱ���yp��[w-���=
Xq�&�\��٘��<�	w���W6�M���3,*ﴥuH=�����,��ץ!ٺc�~��<��4O�;���3�[���jw38"id���M�(G5z�v����:\�
��������@�^*P9��A��d ��

Y���1�����t�e��kN�c����)b�e�����aQs�[��`�b8Ԣ��u�}��_Gۓ(�񟴿��4t�_���K�8h4e����]jR�A���g�?�b�������%l.>���	����;s�*�s��Uk��:Ũ�1�Z�@���x�Ж���eH/`+��s�mQr�ٳq�}���Ը��kx>ۈ�a�^�����ַ��5-����z�
9��$��RBG�5�I_^��$�V���}�<�J]ʘ�����Ol"쇏�/�캣o���'�;�߷  61�A>����~��j��Xv��B�X�@t���.?#�yդ�	uĨ�!�b���'3�{�^�aC�7�N�(�s�+��*�O��G��DWA�|T�J+����ӉC�O�e���J%�\}p��'g��d����>�ӷwN�àU���ės��{���u�T�/[��+^s �L�8�Z�@>S0K��:rF�M���i󃚺�8Ç�%.�-\�K��ň��P9t:<� J�-�E�ɴCe��񢊦�~�M�6Ғ�{��
�[5��l��1J�XCB���xx�����+)��I���v`t�i=^���;�T��3�)H�v\k��ˈ�y���"9E�ʇ��j�AE�����eT]h8�����Ԏ���6�Mi�WZF'�h�"�+��@h����D>�5�]c�4j��Ƽ@7 F	w��`�l/��"�&߽��^@�Tس��P��{Ԕ4E�?7r���gr#>c����Bh�˔���?h��.J�UK�I)i��L{���b�B��%xw � �6���	+�I�^�Q3Ω[�	�!�J�T�����>�	t�@qK���g���e����1��ދGlb?�\ t�q>Eq 5/YK��.��-�7�
J!6y1�c�z��(�g����H��`v�����ɽ`�#���$��O��k���������=CSY2��w�H8v�3y����Ӂ�_duT�{55���\,��V$'��&َaC�sCz׊�$ރ��6A~�<L��$x�MD ��Vl.7-�H���������i����Ml.��֧]��p�[dm�M���h�O��VSr#�>���K��M^��Q� ���w[� Gu� ~��_��6�d��ە�!�M������[&uf��u��;I�3����^m:�w��l׀�˼r�=�
����uE��t�r�Y]�X�k3pV$=��J�2��0����aB[:I��_D����r�6����
�A��9AU�P�"�~�L�<��[zӂ>]	�۔r��E��(�Ϝ�Y:����S�.�_�pӈg"�E!}��#�I
ڒ��g�]�ش��l�ʧ;��f�'����su��5����ȵ;{�E�}�_�xD"RU����5��A�on�h<S/�~��f���H�Zj��&����7'xӞ?B����� ��\�ba^�@]&/j\6P$�*���wc��q�~^��,�A��?�� �*��cL3v���g�G����09�$h~ۨ	�nMϖS�Ȭ��P�@�%G��p6z�$����js>�݊y�sSb�TN/D�3���W�)���׿�ԇ�H���I�>�r�|"���a��՚�=��i����CIYU����9�x���@��d�Kt��f��=	qYմR'�_���!�1D^���������2�8�<[N<E�/Z�Q>S�"�I�z���-�c5�(+I��W+�(7:O	�hD9IX���	bY��k3�:�Z����N#c�^��0��a��%a5�X@٩jIy�p/�u�k��6��}��j��Zz�@�:�6�P�Q��8�r{�)���p��ʪ����u� �r�O"��.i��B�v�;�����:x�+T�r)b�M�A;�����S14if��r5�c�	&��a`���$���ۡ�O��qJ!�S6�Ԑ�R"�K�I-�����}G�P���c��X�ӈg_a�K�舰���Z��s��;��>&�A�d�O=^_�(B�}���]Z�4��Ͽ�N��'|S\o�%)g`rC��9�
�:]�ȹCs)��7/I�N$��o�ԑ����Π��SL��cù5�ǅy��!ڂ���S��>.�
~���� �%!砥'-�� @Α��w��6B�E���aQʱ=�&ms�S0�� ���������>$��F1Q�r2Z�}/�Z�ލzY6V�#>�I@�XY7�_��C�̤@F�)��|P����B�$;�By��!ndj8�*������=�ˎΓUi�u70R>����N���*(خ e^D��*�PG���,A/�I����+��\-���]�O��ΙDU�}���~��<�������a.w<�N�0 =�媥@���)�;N������)BymQ�\	b�?>��*�Vn|��S.[� ��$E�C!yaHy�0�|V]R�,�x���r������s��UTu��+��Xٓ@�+��X��B���'\�ȓi-)�ö}������Tf�щչX#A6��g�}QQ-�����rEA6�j���^��lh���6 �{��.n�8�y-�� IT&1.}���:����9����4�ot팒��
ݜ)��t�N����l�X	�8糋jP!�j �|����S��~fd�YŶت��aIk���O���%�C�kE?�����׌I�`��M?v#�o ��sТ�o�F���6�}���ie%&���R���0�}��X���jϻ�7�]�sz�h��;
�̼�e��b*f�%ar�@����'�5L��[H���:#7�^F���߲ý�I��x��@�ZV=����f��
T���C����՚�u�p�D��h�g���$���X��*@��2+�V���A��ť��m�N�D���Ѩ��ܽZ��+�ړ�|L�sx��4�xm�]�r�@\6`F17]C�M+�����K��d�x�Ƌ:j��U��+g�(�}�V��z>����@<��3?���C>����Y$��4��&vFuw��ꆎ��\�f��"Zz�W����wJl��A��������a>��I�?x-�2m4��#O.?f��f�8�X��=O����� }�
��B����-��% -H��Y�6(��i�G��I���~�B!�m�ިH��in�((��=�
'�]�nJDE��/���Gc؜��a�Z������m��a�\�1!�])zE��rU�����!q��<C:8�*���eG�Uv�$�i�2���'����@��_�E��u���Ƒ3E�/�M@���?p�5Ч����_��U\[��<��uxnlwKM1�)����%�c�W�x�_�6֪�4X�]\�W
\�P{؞;b�2mn�]֖-��Lӊ6�T��W���2f��~�T�pT�le��.��H��C�sq��gX�Չ�g�DX5Mgj@l��w��z�p/�Q6Zz����#�c���N3�^�t��x%��C���l�Z�TO,~v
�㰄����vg���V#�� �#'�J����,We��?�{�:�S�{�zM�A�_�"�C9�?�l�/����u|ׇ�@%�"�L-���ż�Bd�D���w5g+�s�d��3����C��=T).u����E��ЗfM+C��$ib{͠�#@����
m)'���{e�1-g�u�}�nC���id|e�tܗ������H��YN���G��%���`�����o5�Y��2��r��5Ԣ]��'L�������&��v�m�)��W��kwm�8-
3v��31����ޟm=�h6��Q{a:y��x�ͱI��G��r�����	����c����6E�fD��*U1���9�n<����s��JI�d ̋s���Q�NM���u-�f��0@2m�"I2�+>2�_W�3b9i<��'[htGnA���X�0��A��շ��.�Ř��0$%(���Y�i�L��ƌ0��	��u����"��Wp1Ǽ���@*
�A`�%��މ�l���m/'��;�֜9Y�Y���W� ���K�<XE0�6	zH��U�Y��Ps�&�a��7��9�,��Sݪ�:����I��!O]�nN��� �R�2+���
V��WU��z:q?1av�~���@[�Q�y��Z"�N>F=�Ǚ�ٓ�z�\U�p����N'�[���w��UG$�f.������*�k�]�m���N�/�]����f����^�I���I������F�@�7J��D���Mb�X�z�~���Űo���tL���l��ԋz� ^�̄c�����qC���G�H5n�S��á������� ��CC���S֊�!��#?��Cmnm���Į��,SG��C\����t�w�Y�b����\��z0aj�����=_Q\ #7v:���2��MG9!bio�i�Ǿ�YR�L[���<�X	��<$�jY�G���*=}�3{ ��;9�bA�[�n��r�`ި��	EuU��M����'e�-5	�bGZAk��?'��d�n����81�;k	�W�ȍi��ャq���¨A��i����A�������z�Q&�$gdq`{�)��g*�U�(Gcx]B^���ya��u~�U�z�Ӻ���f� �1�c�R>ʴ���.\7��26<��^�|�G����3�ZzI�m;S�L��7b���;���/��0����*8e������r��/����Ջ�����i���bk氻Q��;�eKd�ww3��>��f�����������Lz��s��V��3jO/{���9�u~T��{`
�a)ȼM��Opum��� G���k��.�ͪ�.u�I��VrJ��e��෣���n%W��7CE|�eLm�ʭ��4��t~��kvoI��� �Ǯ5��E�-�� On���F�Dp'�D�z`w/��QP;)�䲰�¿j+���;ˊP�kΝn	_nmP;s,�r�%���~)y�a?�a�g�ږ*���
O��O���x3�/ȓQK��&��od�_���^O�6'��h��a�QB�a�8�����PE����[Y�C�I�W����#�`�=~8?��U��;�h��0�:iR!^�\��l�0���ѹu�%�B͕�=����nK�C�l:��
u��ɸsOuL.1a]�*�dt�f�l�c���a,�ÿ��Ry�BA闅(4���C��B/ሑ��#��5G�q-;������T��?�lf�;B\SSmcC�ݓ�}�t��n��T����{a2o���6�n��n9}�,��-�&$2GXo����լ��X���y�E������C���p���W����p4���J�~�3HU�R֯g�eo/�B�@.tO�F<��z�4�?�Iv޼��dR�Ox���Xhk�f��߇�q��]z2�	����h����n�X�5��G�4~����
aV9�J?K�XCZ�JR�w2&Z�9��ӠSl��˨̻n����%��/�
/���Mm�ޢ�v�a���O�w ]�XT�9/�e�H�'敼Q�MX4D����W[��0��	E���[1KSK��3�m?�T"���:�[�ǨD����ZF�"�'l���T�*��h�K�}�f�.<vc�H�,A�q�.
�R/(4̺���ԁs��ר2g9./npW����k����g��&;�<rV��Ҍﭼ��bz����v��&���K�ʓ�� qF}��h�JD��=ĉ��pԕ�n�߫��S�®� ?B*�'♼Z$��*ڤ^W�J8�Е4Y�'mkO��B�,�����a����q��1�
�^��8As�Γ^���*?b4�(���u�/��^'t�Y"o'���Α�D���M���~M5��������t�}m �+�H���7$n����Ĕ�b��ĤP���
�E�����-��B���-*�	� ����M�i%
ӻS��4	��lRt�E�0��~�( �p�@N�	ڌ'p-������3^y������J3�l���f���;��R�P��� QS��_��$ B�PX50�NSE"�%�k^�9עe��82�����Jẍ�`z5F����g%������ �TY�"�a��(�6-�#�^�5���a�?��ȷF�.P�
�8��kM-�v0���d�����[��u��~�JaT�#Z�S���.�q>
V��j<-��&���Ǵ:Fxg�bT&�ꦵ�œ*G4G����0�%S`tz��ts�L��X1O7���x������g�V)���"Q^b�`�y$�J�(Ӂ(�ޟ��Y'�*KW�{\2�����|Mﶉ�����W�Eӂ���ڀD���y���3����-KЩ���}�`�GԈ�}w�ȼ�����};a.� �7�!�.��!�!2�	"p�c�~9N��'[7蚏�f;@�iH�%9B�o<� }���q�y��FN�	-���;���[�q�'ȏ�b�+&;�D��e���r�zO b֗!�>��
6��$�]-�7�b,�`�j����G^﫡��Aޤk�~{@e��Sˉs4%M�d��)9�ïv{��`�vRV�1}�������gi��h��H�ŀ����M,M2�}:��2�X;:� |G�$9�E��)��x�Γ��������Y�nֻ�N�o��O��U�T��3�L.�c7�'R�xQ�"FЗW�O�=ń��l�9�ܭ��no6��>��k�]uۥ��8�k��%���"�fbl����@���@Sٞ�b8�jPՓ({��]Cر���ǯ'%�A�q
�x;�>בSX$��g��Y�vx����Vh�5�?�sx}�d�'��?��@C����R,���i����>��pN��貂�G̃��(4r��jg�{�<@-f��2�{�>�<��0y�_.���ky����yY�p�'c0�ۄ���L��9eDH�Q�]�Ҍ_~��l+�^`/A'%pW��id�f�R�n܂�d��S�)��ψJ��ߵy.��WɅV�L�=�M���D�=� ���
.�^��:&������2w����6۽!�*��8�p[�+�s�-2�ɜ,� ���ǀ~��;#���: ���L�m4�e�}{�k���u��m�-�U��@��Y��ľj�:������� �跿��Y�R}�q�%^��JS���ȴ.vU��p���%��~#��S��R�4�1ou����uQxT���/bMW��,�LƑ���}�)�����F��n�[��i�"�Q��׭�g�����D�8�;�
��K��:��3I�a��w<he�\N��p�38���r��15MH��?k�V�V�zR,=�MbY46Թ3�C��=�]��]�>�`8�rU�_2�������GV��b�&�'�w�!-�>��@��l0�d���^;_`�k�fm���.�@Aѱ߻���O�ƚz�S�$��6W*���~����4.�D}�#�s�9�XgJ��h{��,��z�=�5C��w �����9����`�S�p���J=��^O[���5	J�A&���v��yW�.[u�F��. �yR��Gk�@2l�3������6P�5�M�4���=�����1��`<�Mbck��]���%G�;Ʊ�\p���3fTq6J��惠��[���H:��>>�,�, 2����g�iQ�I"��t<�c�����C�>��� [���$�j�|Z��%w>�C�Ah`>�*��N�F^k딍��ԡ� ˕ �����L�Y�P�nK	�&{�'�v�X}�}l�}�C(�������`%�_!��k�v:wن�����N,��� �WL6p/�(�9XR[��L�ye�vh�F_�����P;Ȥ+����o9#�����3<��XǕ�7Q��� G�ID��F��@�Jtw�����6��-4<�ﱹ��������T�K]��t�w@ �9�h�:���[s|)Sb�����'זX7���{�T�ԧꐓ
�TS�A�4韱#S�-����ϦS�}e��!�p�|��SF�nY,`����H�G��C���kZ���o�T�@9'YX��˗�Ҿ�Aƿ�v���IL�/)�W��P6>0S�9�y�ښw�!9O`
��$���l�J�G��#�K��{���+���&q�D��.@o|��П�.�w�@o���a.W\���ѩf;v�M	�b��I�f��l��ؿ�n��(��/�Z�:E ���1��o	���L35��Q�	�T������!}RuQ-%�����).�����j ��\��W)�
�Ћs(���E��a�Q������V�%�,�(�L�э��;�I��޻>=�����0���12��<�L��Q�h���9�zc��<��;p;� ^�&=G�p��	
�Q�fd�#��`M�@�G{\ـvcѿ���cJ�n�ﬡϴ�Y0͊�u���=m��i~``~�g@%Ք��s���o��-��Z��3����®�x�ǩ �{���)Q�<&Q�71�Έ���*�$}ܘ��.[�+ޠ�ݖ�Ƚ�m����a�tY�:u��JkrS��[z �n���{�
�Mw�F���ި>b�������o��Pc��B�C�<��,?�:�.��4M�.�N�$�o�6�2���-ص
�舥��I-����,��%O�a�۫�ME�A���x�V���3h'/��ţ��F���H�G���Ze�>�*y���`�SaY�jHa+��0?�.�t�X�7�	nШ�n4z��<^Yo$�7�{�c����Y��$���W�a����A�5%ɭE���&d��s�^���
�x�X��)\1t pi8w���|���F��WF�y��H���
Kz���oЊ�Յ>�n&��~�J�řɬ`q�s�;q�J��T�%�pגn�X��d h8p��w�T�-��okNNǹ(>= �N	im�9Z�#|e�oZW��L�j�ѳbmI�����`x��n�����k���1�;�2��Z�N��GL ���S@� q�>�8�F�'ҏ�׫�*��i�ʚ*c'�UǌONH�U�����9�%Hj�hM�q;��x���ubYW��s?�
�Ş_�Cr���I6��j�hU͇��a��Y�u6����oLei�ch�z_>/|,o���;!� �{�I ������,K��wƢ�N�2��ކ񞻢�����~7R����zWs�[y�%���8�b*�b�0��d�g���q�x�v}�uUIf$�פx�Z�������!Y9M>T��	C��Yν_�t=xY�V�����Q5��y)4�������v��{�`���'"x][W|�}F5�^���M��%.�<�Ґ�\T4|>�F�����rR�W�j�?�)�Ȏ$���#�=������i�Q�#��G�vs�Y���vT���I=b�1M� ��?� ����+��gC�����{(�5	8�KD�CKt?LD�]�dv�=@=��]����y,<[3\cQ6�Vx3�[""a5G|��S�βڝ'�i�$y���`$8��;
]���<���	�K�b��Iw��$�V�B�ѕ�%���k����8���3�Em(0%�?e�:θ#R/��f�X!HG�bIi��H$2��3�:DΜz�����O��ܹzaV��%��>v�J,XB���P0�R��ҫc��br�ot#_�F�fk��l��K`����B���^�0�t�~�����s�>���5=�O�Z�'�뚲(�43�{s������J�j{���xo�.:[�dPy�)���4�݄+vtm*����g��8x|F#�s�/`"����~��{�GQ�w�^(v����"hE�cuN�����Q�O��$]��,�����'z�4��ӌ��V�D+1��צ�O��C�����0Iٞ���5_֪>�o�/rP��ˮh!Ss�\�Ml����Pw�s�be(9��6M��T�f�A|.����Xo����� J@ZO���-�x����pP�;'3Uw?�����W�hkT\U�!���kn
�f�wz	���	���"��ϒC<8�{|#E7<�8�~�J$gE<��Zc{��qom��#d� ��Kj��AHԛK�
�����9�@Yj����'��'c�.�E9�l3TF_B|�)�^ĝ����3�a�@���{�3:��po�d��*����+��Ŋ���K�Vz3��S�m���!�S&S̖�"�γ1�g�k'�rc�����UԼ�cŖ��G�,	a��Z{ۙ���#��~x��И�a�2Ff+M�k��Oơ����]]���O�����{+Q?K��YG���p�ns�uG�X��
A��O��x�t�>e�唑W����rEő���S�A��V�r}3^��3[T�l�M>5�W.��@�!���˔�����1��ˊd�����A��@V(�g��c��=��+����u3�pE�h/d��@>Pu����F;}�>�NHD h@Y�@d�s��=�.�-Z5ݷ����2V�1gF�� ��&����=ђ�%Η�0n\��P�[J��`M�/�_���B�af�(�aU��A��L�.,��y�[��J �CWQ�A��<$�
��c�A ����ӍN�l�7�v�&��m�B���e^%*�mU���z�1��[�j�ڒ�F���B��l5;�I�ջ�~E��&��Ѱdd���@{L}!Ʊ�������Y17J��οP�z\��{*�*o:ď�of�B �����F���ݝV�*.`�&�Q����R�o5��JޗK��_|�3����,诤zo5}�t����;�΀��9a�<�@��߭S��g���0�z��n��7"�V�P��)���
�ݼn�t4�n�`�?�L����!���7d]A���q�k��gkό!XJz��W�γF1����[��m�i�����f�"z�ޜ��ˠ�F W�<8�z������˯�Үs&����?=��DL��:˼Aq9��Q@��*d�k'Qy�lRt�|T�[Q�Z�l� ��F׸-(�p�o�B���������N�t�y��`�LMb(�!�c�?�Y��)J����昉�4yntk5Ao�4f��=Qv��}O�Y�/�d叡
%Ȼʭ�)����?����V?�p��}N���ܔ��R4��y��]��GE�1�$\��a������<5�	��C},O��N���<�V)���p�P�xN��ϖ;�?�%�RK|6��2��<L�*�k��GdDF�;��l[�ܪ�$m��(�*>^)�� 1"��eꠥy����d;�]r:'X�p_ST��p���)Ty\8+n��6ɸq:V����ش1�Z�.{/�K� 7��I�^�O^�k��/��ߍ���7�΅)%~��SH��qf�,�m���L�{��e����B �7�g�t�S���zʉ@8��|���f1w ��7T]S���dT�	��8��iﶬ;B���>�R|�� jR��o��0�i����hՍ���yƋ|4�dR������M�s�+4i����I0�q��}rT��y&
9vG[�>Ӵ������J�+���ڥ#uc'��Pڪ����t�/��� ��| ��g:���Q�O�"nLz!a�M��{\�#�UR &���3�aǮHtS�W��ޏL+�N����&<����f��M��T8�Z�)���Lz�-'SjN_R2�(�G�d�P���P5�A���t���e�c-Ǹ�D��UQ�k�EF0��ܜ5 ���%�rM�Pw\( 3�K�+�K&��&�n�;:5@$3M�4�,���AJ�۪���	:͵�	k4�\�����R�a� ��t(D�ļ]&�@꾦ߋL��l�:�OXk����+ET��uSBObɬZJ4s��{��huή�Ȩ�j����;��hfz�s�O�GB6�]F�!�o})jEk�n�����혨�kDa�{f[�?��s?��Pc�����E�<h������J�FI�qI\�1��zN�A�
�HC��ݭᄇ�T���җޯ��e�PԶa���=�"#�J�8���;	F��9�٤巯�RֽR��Lr3�k|����!ut�j4	|�r�#��̾�5����!Z�|h��D` O�2���������ܚ��o~ su��E�m=6�7���)�EG���4@����dټ}?go�K��[hkÑ9��3��bqx9�,�x�7$��GUws�W&��ږɯ!Gdͳx׿;�ܯ�a�`t��PJ�n+����4/���W@���KM�����D.ZhcT!K�h������>��������Tt8�]�X������1��m�MơoG�`�g��蔆[*����� $9�Yɐ�b[��Z�{�>UO��>�_�W����8qP�F��tZP'R��A����������m���	q^��>�q���-
����	���|&��+�|�(�����؄wU�&n� ��v5��\f�M,Q�lg�i)�<�.V���!�z�SU,bМ�����T�ԓA9��t���)?����ZJ�i4��I����l��W|��91,⁙��ll��Z��^�i��\X/p�����L��|`�}��_صe�&��V˺�N�'�f�[��pbZ2@��+a�pXJ�:tY��Q�@� 1x}���lt�>�3�"�T��f��aep"-��p9�q%�s/_<x~��he8�h�ى�C�5�u��Kv4\ɣy;��ЧlJ��z6lj�s��{��a�^7���Y�X'�gyDYC[��C�s_����
�-[���:���8���`XQ�EQ֊k��΁���*�ԩCq4͞V.��,�	�|R�|�R��1�RU��Zt8jM���Xh2ٶ,FV�Nmr.,-�a�'}Zb9�ʖ˾fbM
�dP�t/�s.OOU#�e`Ȯ��6���Z<f+=A�>���ƥ-��*�e�/n�h��ĖE� lF�)w���^��O˹�J7`���~�Ld�X���}��>�K�?!H�0���ĿF����Q<`0�`W���L����%}-��t��t���l9=�AԿ��63��K%yf!�*�?�����Q���]�]v����6 K�Ⱥ�M��OH}��LJZu��aP��Z���g��h:������������pglZͭu/�FW�;d��k1N0�c�����cn�ן��
K���9�5��E&mH�i�G��t�J���������C_MN=�j�^F��X]�Հ��m�?�f��W����ۉ�z8O�_���b7�d�[�L,�0w�1���`���[˟�춠80����F��۔j�x ��}�b�^��Z@���L�Z��Ȣ��lt�r��[��۳�P�E��	��:<���'X��J5ƭ���G��u)92o�troM~������֦�Oy�G������"m	�cF�]�
ժȈ�,���^3QS�~1��Y�q��&��WW��|�܎��e�i�o�f0`�����+���QB��D�W�SW�� ��|�WG�Mq�:)���S���@�S;��/%ZF�S�3�!�$��PPz���5Md,����J��Y.���b�:�a�[�
��ߴʃ{��_�e;-G�k	��y=���x����,�;t*G ^�E��noײ5�
)ؘ�5����6��΀fB���U�T���ߝ(���ړ����8��\�Ļ(1��t|��g��?�rk�i�T�DJHa�7%�)��_�{��ڨ.�VF|�Õ�{1�1��7f�?�f������AUC~�b��Vvڤ/Gb�/4�}"؅����<d5]��]��pbg����-�]&16���^�T&_75)xoP�j���+An
���q��֖@��t�����`|�q�l���%��;i�[͋�� �e(�[�e0Ǥ?Z<xOҼ8�1��&k���^��G