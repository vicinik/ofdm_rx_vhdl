��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��8&����[,���$� Jkj�P8"�~ꋐ���fi�O��sebZi	���'���f��UlH��:s�P����h�Ǿ�3�ra~��f!9���wJ�zX
8��.H	^U�.ȨN�"H2��<�+1��zA���Y�\o'=Z�:�7��S�%_x@�m<���I�Y��@yA������'>��jcsr��� �����*Ce����(h#�����$=6q�
�o���.f�p���`��R�3Xj8Aq�a��(�|Ō\�����K�S9d�������s_z-fWO�W�%�K�Y�CI;�8���jj�6up8� ���{�8���7�s2gX��g���,@$�����Q�̳�]����nN��]�ϟ��:��G�s�z �9�!_�Me/2�C�{`9�7{�?�I8� ��Ç�Y+�\���|E�n��Za������7��d���= �_η0ȼ���*dX��(y}��~կ�y)ЅeP�n���Ҡ�P<��H�<*%��kmҬ��Q����s�"�E�C�F���G��E���Ϙ1�)x-ǹ���r[�E�%^/dt�j;�&�|�f�e#�~ ���2r�+'�B9�	�3������c�[;�F!,I�z��P[�rO~�y1^E��k//�/i�,��;6ѥNChT48�%��ק�;v��؎� ^2+qn���p�I�#�hN�MFm�{��=n�=�I�_���r��C� �x�d��a^�*�_��(����Z{#9��򭌑��q�n�w1>����,��b`������l�ΤCߖyp8��"�f� ������D)[�`%儩`G��v�PҲa����7D]��^�����Z��I(,\�C�g�J�Ʉ��SE�?7��� �nhSY\�����N=&1\�y͹)�!���z�����A�ٴ;-y����\�I����f�4Z�*�>����>vl"5����o>�q�Ot��j4.�D�d��-���{:�gՠ�J��Q/���I"2{7�SJ��3����4�>�R�B|i��{LX��0�V���/�?S̡�_�"�y�@6�%�@�e԰K]�p��Iq��>*��Y���#�q�4 ����`��ҟP��󂱘H%G�]�$�@q9�������Go������zG��?�Å� 7hLj�y��L���S��6*�����#
��D�?rk��]ƌã���+����L��H���$<=t)�o\fo<���/ro�Ӹ���
G|[vP�'M_�b�/4R�V˲ߠ��G�Թ����mxXO���a��`֣�V"�;�TR�9r���̩�R,��fBFgj��Kr��Qe"x���K�����?��˯�
`��>X�S��Ҫr���`Ċ���B�~.^�T3�N2�ĆA�kh��ܡ	�6^5�p+���_�`�uyx(�'�w>L�y��0(r/�x��5o)t�h}Ǣ��	%��w~q0��)e/J�{��=oդ�Fx��-��#cA��]}�����m?~��l,�����^��a}�$;̍���@�E���p	��d��?مQf ���B Zu[1�=������*�;E���I���W��D�c�@��ò��nZ!�5RG�ꁏ\?�*���� ��*����z��H�ϊ�[�.`�$Tσ!�y=e&Y@j�7G��)ɮB��%XI�)$�ݒOʁ#���ͫr� M{����W�]�����q�חJ�e��X�/�c��t̙��
�����N:�/ u�F�I �C͕���Fl�}��$1��s�h}/�Ma��9�����6,
����2Dad�d�}���`�sK6f*S�� �}+k�KZ�;�=O��[D��p2�`��I0���|�[ډ�P�����xV����~G�T�sQk�=��H����b�ky0���q���t�yv��[d�Mk<�r�rA;�C=��^@M�.��0�̛�%C;��8����m�|�B����"]ŏ�^�<�c���c����B~��7�sKT�6�g	]�oӆ-�P�T�t��c���pC1�Z����Y	K�Ӣ�~�nQ��Ͳ-W�T������*�9�d�qJ���U,J�{�^(��"I�vm�����������T�I`Ҵ�m�� ^�:-��±a��eP�p�'8���c
x��C��~��`И���fo�����?i;��ڕ�U���u�C--ҚJ��?˛e&�1� ���v�F���g4-��N���	������go�W��^M�3,��D�x)�qf?���|83�s,S�b���+�y��R�,[�u�`�j! ��#�r7�2�{6t���Dbh���I����T�+R\C�E��W����z�(I�6�D6C����QY���38�d٥h)P|�]&�K�d:1�k�M���\�NG��LZ��p���@*q�`�����}�X��IT^�[8b���\L�Yߛ��sc���{A�6�\���8v�����p6bצ��V��Ϙ��a���@ޔ�>�i��U��,�7+-��:��=N�>_w�\=���g"��3��^I�@�I(�ad*{o ��L��\�7 �4j�Ik�{�>�*�Y���^۾��ϋ�1%5��H:�T��*;T۬�3������]yN4�\����7]*���פ�dv ���.8yI����h�޵���f9\W��U���Jyж8���|�@��1�d�N�J��q]�ח� �m@���N�Oagx�|B�� �\Y~���e�a��ɾW�O�/BבN+�����-��W2���Z�Y��:ȲX� �2�<B�`c�=s�����i�y���HE�Le�Ȓ�%�;�@�%�V��y$���3rjGK�j��W���m�4B�.OoF�����0�_Y�̟�i�'��f��	��;�A�`��;�.�Ǳe�p/�[�^���+��NB�}���I��Ev�k�!����~��G�)](�V�7��&���E(Ȯ�,�8kd��a�Yk��ؘ{V�����\i���<�2mN��aa���R��sue���yE�81����EL����)�RZ��8�ͅ�-yk�/�r��������n<���=1�-�f���{� ��7M�52i`P��C�1C�^Pب7ָѓ}ޣ����<S�s�S�.3����Xϯ4���W:�	Q�������>�o�p�,�}5T���= �.�K�?'�`�,m�jSZx(���̗Af���6:*��g?��ԿZ���!C�%	�7��A�4"Ww�}Qpg-���/����%��۽��ʗx����.���w��:�S7,����:[ח���ֶQJ*a��C_F���Sk�j��%�pr_�3MH�J=:Y�
ٌV�YR��4��!ia/�c���q��y��lƊB��w9,Q�VN�St	k��$񠕲�kmΠ>��V/>m���r3p�쬈�u���C�1#�4������jk��xŎ���cb��h�᫡�dȻ���<���p��)ѵ��Ȼ��F�٣�;�׷��LaQ�'�k�=����6��L�i{=��n�gvx�s�X���++��:�fa3K�X� ���|���xm��Ù�b������W�(��]�>�cXY:>�"#ђ����-Y�qִ���d�a�Vz(���(�;c�jtz��[�6ߙ\�M��+�����}�|pm�N��QS���N��g��s��Y�_I����	<�dX��В��y�ɛ#�/|����jT,�'}ivw_���K�U\ݹE��<nK.<^�N��Շ/o1-�����E��b�����*>��KZ�5���1,p�=ŗ�0��_�<�+�-'N`y��/����+JI��X+�GZ��c��@-��T���dф��^��$�ֵ����E��A�$����g�����&(�w�Ʊ��]�I����l��[�����a��Aj�*���|�=㴪w4�I;%ݮ��`��	-�J�
cc�ݬU����31!z�AB���L7�����Ϝ�^��Xi�k���d�%\�x	�Dv�O�, ٴ�]�Sx���j�W(z��}0w,9 \"��_0��Z{�A'���=��\��-W�L�a��Ŀ�[ $dQa' 	�ʜ�t�%�q���.�R�<�\�U�?ż �2RB��|�T𱌏��ԃ���i~���w3��~�#%��U�����Y�ؑ��i�?����P3ݫ����A�����p�‖tO�*�{L��29�� ���-��"R�����nӎ
Ƹ�RM�+���d��5f��ј���jS�[��AW!��J�Z��hZ���Srh��b�oQ�=( y7����!�1���.j)4$��,ǺE)��y��@�x��o�4��O�@���(�b� }���;��I����7<�1��:��)�CsGU�E%�̭���	28.!ZIU�!�pm'��sv�r'��щZ��'r���8-�lzf�N�����=~L����aeI�T��jB7 ���H�}M���a����_Xa�K��MB���5���]�nsJ��V�F��bax��������"`��e:�L�f��q>#Ru���7g��J`�ek�A�,O�L�n��s�eSz�O��Κ���ֺ�ّ�)[w��0rG���!Fu��24ƞO?�1�3T�$��1U��Z�Ynt�Y���a�$��*�%�v�{��(nn�I��J�^=q/��_�#<��
�m�������Z"��::�
�]��\������p��1Y�9��*��J�h� ?n�@xw���	��k?<��n�Tύ-�mf��h̍Gan��rύդ�==`�u���z%|5s���*��t��&���u��bYr��O����."xO��~v�*�_� ��K�V�|S���g�7q$���CQ�6���w
-���Z�&s��e��QA]@A4R�bWʅ�L���,E�8�ia-��,z�<�R�g%SS$���tʎ�)��`��KKE����~�k�*?�>����x�l,����l�O=����nђ�|�X�nH8�)�a���PN8�{�O��������]�0Eȁ�����i��_��u�� o~�g����Yr��5�G�⏩��s[R! ��^7�'��q?,&�B`��AZe-���A���p���*Y���V5�'`Qy"d߷��F�O��= l�ܞu�|����-o'��CW���8�b��+L�:�����q5���������d�
�O����C��L=���ؐn���Ӧ!�2�$����F�����m��fP�E��Y����<��p��O�E���xY� m:$��? �h+h�BD�>9��'h�T�,��G؞�91��� ��~�E*��Q ����TB���
��Ċ���;!�5J��0�rҺ�2��m��/(v��^O��aK���i"S�&&�0Q�,�d������t\�G�$��.ʁ��m���C��V��*���/�'(��/�;%������R�4�4��9��2C�ȋy�,��`���j�0MVR�w%+L+xic}�ӓ�b"V%0@�lzV��g�ϧ[S�K�[�ڏ���v`�@j�R?GBo�ȡw Q(d��[ٜ'�=+�)��P�˗A��0�����Sb+��w���"x� o
�J��v`�+,���X�w{U&��v\˻��S�V*�UY�Ps�>x���akYiM��V����!o���z���$��m�<LUeK`(�y=�n���ǆl5w�2���Q7,�:e��Wb����!P�c>�!!��*O�����/9�:=3H<��0G�=u�U�1v�.�#0��i@���_z9Y��k�_�!Df����e� s�s�Hm�� S��V0�T�k\8�hڪ���@־���n��?�t��P��5y͡2�b�פ��*�*�d�]���6�´�Uߜ�+�	�>J��/�$Gu�\B��eI���_y�v�'�D���w.�.P�~cg�2 ��7`g.���K+9COn�uE�����%Sf�!A)������`I`�������Q�H�Mu�q�����Ԗc�Ɇ��}�ԉ��4q�`x���_T�?�Za+�=�q��Mhy�=)s0����a�Y���w�i���_�:�,��B��gMf��#5�x�2�,J�٥���G��}�1YLd�����?!tgMÇvV��MaH����&�ȔGb:�9w7ȯ�����!ݬ�8n�ږ��+�!�����Դw�C����ƿ��
� Z�
 &�m����0������X�8@-fUx�$t�ql^4�
P]+R�@���S��D�E
JӀTY|0'A%N�kH����̽s[G�e��[YB�|��ѳh�G4�V���'�#zf[��:�f���ԯ`j2+Ht���#�#Q(ªlo)���`��]IV�M�D�9��*� ���ƞ��`4_Ļ���@��>�~�p�/����E�\�b�q.��R���>ߊ�R�+����	{,���`���h	�Ιs�تN�����T�3@a��*�2h)�YK���w��Y|��A�y��0�E%/,�[I��jiB�<��{��[�rkX���ӿ�Q6�y�)j�y�\,�F�8,�Lk>�����a��p�����p��sQ�d
aŤ<��EiP��d ��p80)SDP��ApOLHhؤ���04�����q��T�^��¬�<A����T����@eC�ZwK��ŉ���PN�{hr��n�_H�k�6��Z;O�4��O���O6��K\8{�4��3e툿!�N��jg�衑���c����M�9��fx��U�ʍ���>�S_
G��W!�%����P$�
���vB:Շ��X\�YY����������](W�M��ɓX�s�	.~>�V�����*���Ԡ�/\Bϗ���_q�Ry��y�VP���*�MN�^	�:����wL��� ��Jé9��㒭8p|$� ����L����ߚ�B&Śx�����&��������h�C�*Q)Y�����fsG﫬��NRE��Ax���[�n�*-���i�w6�� �qH�ϳ�W
�D�QK�Tћ1��$��{&��6z��p4]{ٚO(�!Qdߧ��g�v��C��������]׃�?�tc$jZ���6��{ǒ��x�b�4Y�2�2�L�+ 8�a�b3��j�3��EVZ�5�h�6q���o�
�zɂCD	����VH��W+� @�j�sʄArPt��5���,�s���������`ᯪ$��0��6���>��h�*���Q0� \��Y�4����g8�c@��I����^m��H(�(g �v��%��~��ۘ�Q����f2�n�X�U�zv:1,w��D���w���1�w���TM�)cQ�j	'��ӥ�R��%lE	W��c�<�nl{���O{vSb���������_%@��N��΅k�����e+H�5ɰ�+O�%����\�QF��l���#���~���k.9���2˚������,ַ3��g�#�{�`7�����,>��j�d�,�f��ou�6�"Ɲ��PD_3�6@��g4���UQ�f�����H�����MH˵lb[�r7��4���k3&�(�T��L"���f���L��F0~f�mwI����Eb�׵���c\'M߆9T��9�������Û�6>�Ay���x���&v7;((���H2ޑ�z����lU��`��~=�q��3B}C�a�Gʄ0�S*퐆^$F�
K�l\���TJH�[K�M:����	����cWk��ir_J����:q�8��<�M�~���?��O��2��;X2qo��w�'�� %��&UbJ�	
Nzf�g��~<Cщ�iG��5gW��mH4�ҫZFZ��-}��J !���4�s�,��fP�ԑ���(X�;��^��Є����U�!e�z�L�d+�@B�#�����~�6���f5Dk���ӱ�`w�z�(}�>��qP�2�-K���R�]�2W
�E`�0��P�>�4�I�<�@/0�&�
ɤ�z���Ik֌���|���K%�U؆cA���rb�9{���MJ{u��xq;�ڬl!쳁z����P���լ��L��9�4�;m��7*̗��6�Y��*�~q`�s7���e��v�*��W��ۿ,!M�^���F�3旃��\�Y�r/����|�� �=�o���n�4kɏ��U�R����]�n�@L	���jG�=�F04��~f�'���È!r[���V�>�Z~ �5Ig�ϺÊK�[��!Dנ4�?��i��י��G"��\��V��6r�@ْ��n�qc�� ���j'��"�1�Q'l��C��AF�`5�^c�T�7Ӂ��~��Cn���N36��6�R�_��$YS�+�ƞU~����sV-��1�b�"Ц�!������{� /p��(Ԁ����O1�&;�j��yG�l 8�_�h���cSs*�{��D�=������>	��̵8�� L,��;�w��
���Ұ�1
˖[��l�x��Ml
l��4�8tg�o£|\%ӭ��[<�{��&�dvvJ�����F}Ͻ�7�Jų۴��R̶ nZ���	���7ӺK���!֭"�Q���rd�k�z���R�5��	���VC�~�!�{�Mڷ�~�����2��I�v���MօS�d���������<����~�*�gR�r=�xe��� ��#�j%bL���֣ۇ�c��eX�,����9���Ƿ��G*�i���� �����$7{��!R�=��U��$��2��p��s��)\WV;c�ւ2������M������&�A`��ŀ8�6�9rk�:s[J{K�A0��?/���m@��?_rv�W��� �
W��b����pNI��mKW���϶�:�&�H��������v"5�=U�����#F8���}�Y���,@U?$0yB�,���� �1VVՄ��
���sQ�/�닙�/r_|��x��l+��!SN�a<L���l�j�rL����&��D[dI��x!�xIlw�C��N��bv�#xD�JI��lCkI�أRn��-��7�i��5��[&,����T�]��ğl�E��0ys	�������X��j;�Xz�]��$*��H?}�~:َ�|¡�qc&�{�F����F]��r�Ǆ����'	荓��J�F��}Ņѽ/��4��U���}�rK�VzI�,$1���l]+|�k��޼6-�-���������v����Z)��4��I>@�ݩ�Nѐ;�O�������Ȳ@��&����I/%�>�D�.x�`�F�m9�aY�=:<�a���ʸr�Qq��$�,8t�ʹ��
��=��S���Գux.^1�l���]0h����&Z�]p��E�|���{�6ԦSBI&W�uyQ��t!d�js*E�@u�����>ߐ R�8Yh� ��c���o
��uL�ژ$3F�#��B��(�n�C
MnIX�Ⱥ�u��A�&,RCA�[���rC����|L]e�N%��c�:��	V�y��s���`%wZС��C�,i'�7����k�Z�6�Ʊ����]�*%�o/A%�*c]��>i����8Z/&�+�&�&5��W����KQ���(_Cl=��n���l�����EYa�.
����ǣ׏��xZGd�
��3�3��ec��ϽC�b�I1�C�<Tz�[�8���鹢�w}��JY�Gi��񐞝�wx���Ac���s�	�LP��;Cp&�V\�]U���n�=��/|��hy}[y�N�yV�,�m@j�@�ֳ�v��A��~����F�]�A�O���Θ�ʚ���x�� �P�D<�pS.Gvk�(r��H�������Q����l� )����A�b��"C�	�Г6(��=Ǉ��ul�K�m��G�xץ9svݎ�^F�Y~����{�N��Q���j�}h��S�x@�`6��o�Q�3;��Knk(_Q�7���)�����bG븾#]dsӤH�Vx1;UO,��C@,հ��Q���dzA���6@�}�+?߭�Y>���Ϋ���kyw1c9k��1(���%v��#o ����gh�^��Y�pbvk��>��I46�\��,C���r��D�sw�(������y@Ǿ���S����1�O��Ħ\�l��ń��5_����x��T�R���fF����r��Z�ю�6�Lǡ�@i������IC7he���k�ھ!�}�V2Y�X˜)K{J�$nP�(r^0)���y9��^ᡢ����6��i���`y]،��r\���ۇB�I��Jŝ"���7�o��	p?=��]�`�
!�"�yp9�4L���$9���5���Q���!瓄Fn��=7�)��eZ�m�/�q^��F��Hd�}1�AMc(d��ow�P;Y �h���g�����\��sr���H����O���_�,h;�H�MF:5z�P��{��Dԡ��'�S��3�ϒ|rh����ma����YN�zv���<]��a^qS�@C ��Q�4�px�N-��|R��_�
O/�QT��d��Y�yKg>7/��q�K?���m.�d�/�h�$�D����Jǻ=$j�앯��p_�<�(�-�u��&��;-�Õ�KH`�,ӞX�>��C�|�/ �koDʣo|�VH"Wd�"���'����.���|�U��y�AΪ����5v�E�S�ǈ���3��|f���<���P!;v\�s�˃�1��`���C�$9;8ɮ�hG�Ó?�׫h��/��xN]�6��nCU���y�v�H����a�v62Q!��xt;����\�j�~�iV�E����x��F��
�%�dՃ�&�a���R�Ǒt�\��E��[wB�:�>=��l�x��8�~e��p ��Z-U��F£ŅC(^S�$U����:]���vk���G�q0��c��ُ	)i�&�Do!��%/O����p<�����I!V�+�����aU/��z�f�t|N���@����S��	�[g��+��|h@><�8�,�*�hLf�6���Ԡi�$E+YR���%r�JL�ob6-4L��֩\����G��M���}��f���s ޅw�y4	{���f�&Lul��V�_+� ����6y�l>w�� kDW�xZ�YK��:��u��`W�wE/|UNPy3zH�U��Ԥ7�[�SZp���.$\��5i�[-��(�d�G��e��sei>ѱ~U��'�*k��� �5����4c�� &��;Z�>�s���P]p�S�0��^E:�]�I��,T4x�)�D��	�,��w�B�.�~������X �֩}5�_��ʠ���V�����Ҫ�em�I��0	����k�#�x�=0R��:��eSn
���𴜝�����m�ݝ��}�����1�f��L.�"&{5��);�$oFJE;��������%b�������睵��d�jd��/㈍�0N�6We���G0�39��XH���p���5�y�N���N
���;�B���󯕾�yH0�?(	C6�P����
"�]��׫�t��c�܁�n~��;�Ծ�!,M�� `pr��_$�d}��ײ'�,� �`�;�����C%�G��ά��}���L�w�gp,�<1@`z$�v���!e���� p���Ar��o"��AuNm9��9Õ;�� S/�7���W��r������t�^�꽮/t�v���A��(��=�=�ѻ��������d����=Dr��۴[.	,C���}H����� y�����G).m�Z��B+Ɍ��$��S���g�`�Ǟ���o�/x��l����)jO���*h/d]�S:~�#���ڍm��s.A���X��vַ�Ђ�
��9�A��0
�Fa�R�R5/\��2@;�[����!H���|u����v8x��6a�]�I��Ձ\�#'�4��.�ω�e�򆻖�#��i9���;�%�Z�s?
��f�{F/�6�3t}3�2c�:���@��O���1.A;΃C���\��C����C�JפG�� K%�w�nF��`t+���/�GpiO��^�	)*��SvҤc���d���MQ���֚z�/N��~�ީ�n�l{����5-�+��cGR��UbҴ���C;�l���8"���Pa�NAߜ�,Ӕf�m���-�{j-�-��	ћV_g��Coi"U�8�"�!aj6*f���?*b8�-���Qi���|��W9&#,y���B�%$d��1��Z���A��(���,F}X��{�M��!���M&
�[��G%盂�膴m�E�R������5Q'�;W��r��0]"�[z�Lm��B~��;G3P�_�J"f{�S��'Y�����'קּ����a,�"9����9b�5mK���*���9 u!#%�E�s��,6z>��A��n�rN<{#�
P���#��H�-����F{0��4 ������B�PI�{PVi��v��n�����&������D���>^�j1 #��0I��/.��d�'���-
ʟ.�%�hԪ:uƅ\x�E;h?��PV��{��ݝ�=ʲ8��T������ͦI_�O�<�T�+��M�lRf�c����ڼ��/�mCvs��2�LaK_}�Ù�#��Q@�&꜅���G�x;���;�F����y9qt'�^�E�NH�����F$6Ld��fJYg�����>��z��
�5G�N<��Q���i����,1�.�p�+��$�:���2j�R�q/����*M]y?c)�@CC
�o?�~�]�W�v��4}1�_��)�']�)> ���Tj�b6��8�b��ir��uV-ii1>�M^�Hy�h�u�wEk�o������<��2����t%����'�Ə���d40#�Hc�E^m6�PC�ݽߘZfg��_��T�Ϳi/����^�4i/o�|ɚ�y��S�B�a�� 'w+�5|�#W,�1y���K��KG&���u����rl�;�K�۬��%���?c y��d���{7�!�ňLށGiq.��_*��b�gU��������b������T�W`�sF;��kTd�իu�+P
�ʌp^�Q7{*��"7��.J|qH��<�x���
�秖e�T��y2R�Ie:U:�hI�k����i"b$��{~����1�y� r�
�eu>t��`��j�R��F�4R�dQQ�\�����sa���#�hn&1�̳_��mȲ�5�{]��l�)2�D�P�ڙ���R�L�tYY�o�<���I��d�� ���2kh��L���D@���H�l!5@S�.�+���������%�
�C]�u�n�)�?��,��?ĈdC�y}�������>d�%]>�z �����޻�}���s0D��	�M����Y�{�v�2zI��N�̞�-�m���.��.Q*��ԗk{�}�.�l$A�f�p�A�)P�w�g�7F:�����a��-��w��D��m�ҮU��6A�9T�G�$���R��YDu!˓QT�E/l1X���G=|�Ԅ̸��4��w�R���d.�I�RÉ���HI��j�O�d�br�����/�cU��x�N�_���.7�)�c~T�F��j�EB|};wb�}~�ɧ�.��y�_Q�j_�\u�u"������es<�v@��� ���=��t9SHG� ��[���.�a�̜���TV����˰�(�����y�d�NA�*-
3�:�.b��X�TS.1�yB6U��qf��R�8H��W�ѹYk�L^�K�ȋA�Ս��E�ms����Z s췫j�����S���#;�C>�VԽccn|���ݷ���Ud�(��k3t@��H���6�}���,"��#�،��t�Λ���*��^��d4�/K��:�m�~��.�L�\���cS .�u�J�C[j�|�o���?�f��(��Լ�����A�H�L�o�0�]��o ���]r!����v�!_e�����8\�5��Ug���z��ۓ�*]�9�,(�M(�6fG�S^��q��z���"�_��"�j5l9A��̕&[�e�O��ū�SӲ�.��:aI�D����V�{�	_�b�$�k����T�ɳ�~#t��azXk'ϟG�El��[����|�U��"�8#y�P�/X��i�LT_���|,�*G��a�Ι� <�`��N�sէ��`�C( Uy��
��dI�1^E����7�^����Û�*S�X�]�l�L��h2����I��/�C�=�BP熟�y��o�w��NeOJ�T2�A$,^�M}��+�c��������3׍�p���Rг���28Ũ뫤k�R���7�_g: U�������8��;8d��� ��Q���{�{�����}S�겙��/��Y���M���xq����k�Z�E�'� X�6���'c<�Q��E���Y�W�N)�:B9P<�#����F�8�.�a�a�/�_�_$�j��E:7��[�n A�Xh���Ҧ��t8=�ޱb!��|�K>��8 oZ�a;9l3�LLP�o�W��7B3��L��>��6�2)����~���+i�Vp�SA?ڙ:K���'�����_=9yP4_C��^}ȝ�K��A�ǁqF`�0����Tq�2����}u�;�ƚ�e�0h��v��$��~���Y~g�uk��q��Π��C����C`���9'4��O�9Ƕ�~�8DW�����'��Sf�0G��r�Y[A�*Ex�	G��k�%��K��'� �Cw�D�#͛,���z�aM�����_I؄�E�U���1Cȃ7*���C>.����bV=a���@gn�N�s(���;����.,�7dv���d[�YET���*ݖ��Eq��A�������;�r���;^D+5�/0K��4v9��ٺ䯉�G���3DO�����b@�Q���2�gE��ܳ�~X�����J��*����Tmi4F�y��gY��b+ݗژ��U�_�<$���}�1��QG`�`�R���[��PM��ԉu���`�5�����c������rO�F7�2/m���f��Z
�P�s8��j��]H�cA��Z�pK/��Ŧ�Dĸd��6!-W@13GЬ"@�=tN����z�0bўm�D��d���G�{�Y �@��ʒH"�v/�gµ��K�-��!��W*�(��p��B������ɝŞ�
�[��p�lN�/���,=����Z5A�+��>��d�Q�"HspN�W�_s��R��1)����-%P�.�~�\&)�G�����������ǋ��=n��lP=�E���lU~�Y_y��T+��1j)9�L����}V<al��9���S#���s$j��;�3<7��T�0^���F�y�ӕ�4(�Ҭ߁��BU����'P���"�M��A����f�$K��[5��ڮ�#���Q�7����zX��.����ԋ�1��U��@}q�. �>ٰ���s��P�g���~7���Cf3�oS���nO��(��h����n�A�YBʌ������{vQ:`��D� ���7Ӛ��|���/�c��У��H�,��ἠ��������C�v@�U���(B����������[ rwsh������I����!�$�Lא-�:��Byoəj�v�H��c��"�;��
��RB=�en�q��|^5K��J��@b����hX�Q�7f$��S�Q�=��"�Vo =K=���L�i��gpd�'��H@�v³����@�F���Ȱ�-{��Ue�|��UK���PB�Jz�t2צ�E*B�jީ���1)N���Jԃ��;#���"ٳ�O���?�c���na|�eE��.}n�U�&�[DE�@:��ks_�gF�G�C�}��s���A�#Y1�	q<ӗ�)�2>�_8YZ �2��*�<�����R��_����4])jG�����d���ק7���ex���f:�S�5f��R���y��S��R�/F-���!:jf�B&�=���-���.2�W\�	���ۇ�}��g-����DDr<�u�W���y�ص#$dX<�΅��2��9���C,���{ Z1v��-���DF�2c�-�8����0������$𗭸��1\l���f�B��VF�����r��D[#���y�¼��?�bgx�������س� ���q��*�u�����#_+8���󏾝5>>X�����*�^@�%#����g�8c0TL$�A�zQ�s=+��t.����Qጟ�_�G{����HK����ϻY��v�@yT?��e������s;��(�w��
<tU+��t	�����2JU�Bl�:�}B�Eh��+F����[7l&J�8�Jh���rٝL~r�΁��!��i�֨Zݴ�|��6��r6-��a /�@J��"V=o7N�0��㢪��o��p �]Q�i���ҋY����.� ��W"�M���y��rsr-�l�{�XcK[�C�_�w�2#"{J��O������=�y(κ�l�����K6�̞�,����@]F#�w+4FFF�x��Z�O�������Ws�gx�t|�d��g���W4�� '�q�h��y��W&��ښ��2���ɓo�R�0��n��"a�"�����V��݌�W�����xdc�����%"�v�==��$�X_�42K�|��6M�MRa6=��w��w��J��t�ʬ?�}0��� (
AX�͢$2w^����!�dx���U�J�f�)]���r���!]��Ad87��#��qTx{MOw�A5Qq���>�yu$]�^��<���r�AZρ���\@�vg����lM%R	+��~[�vO�h�gE��!�I���K�LbM�a߻>����MY
;!��$:�(���H=,B>����������d����J&R*$���zl���S��N���l�7lB���s(r�
M���g��j�"��ܚ����˿�E�Ը&"��T�N4��I����W?4�=qL��_�\�8�f��NY�4�"�L�4#
�y��u!c���|*�#}o-��U������e��EJ��}V@��5����q���9��I#~rm_��X���f!���a���jxm2\h�� �à%|�ZJۍ1;�9��S����=�g�N�w}�ӽ�Ο��D��zf{=4a�zE�;\2��00q����Ik�Ǚ�_m��H����a�a��?U�|,�� ���a���xQV͜<��כӪ{��GL?O+��&L�S#�3�e��$�^��Ab~���2�+DA˸���(��O=��'j~�%B	&��Z���5? ������IM����2�Yr��Z��4��jN5���N��8�u��|B0��B���ZD��?��t�:�Z�=�a��mީn.�0�IϚG����Q�%��]�V|?`o��Q�J��� �]m��u�?<��g�
�����u�p�+C��9͡��J��jR;��$��j?�0�����bz#GZ��BO����cuP%��G��.c(j�Zz�%	׮�%��B��ހ�e��
�)���G�#L�����TJ���^D��7ulc9�e��!�a�t#��_"��S�:��CO�Y��[�#����4��������M�������8�*��i������㛇��k�P�5�~�����\�J�W�X�֌� ���P�B}r]B�|���RK��#��c�J%fx��^���x�g������=сimf|�I�=�>����&W���;�Ue���!%7Q�ڪD�(h�ki!o��"|ef�I��?�X͹�4m�_&hZ�NC�T�a����d�m8�\��e��r�Y0�#
�Ŝ$3���3p�v�J�K�ϫ~^2\�tAȸ�=��[�`H�O��������ʪG�_����O���I��.Q��̥'�1�q7��$�G8T���>j�n!#��ސɳ�N��P�	�7�h�~Fà��7=��n�C21��E�Ý[������Z���u�4Z�+��hK���a���N�C���8�_~ �����4�#h�(W��f��k���&QP���lN�A�tJ��Y#��;7�d�d�4)L
��X�{*���V1.%�� �-��%���|��+��d��$���a�j��4 ���$�c喫�B
p �<���e�m!.��	����(Q܈EQtX�&ǈC�NUL������l__	p/mxܯп��:��+g�������$�J(Ջ�B%ˁ3l ���C"+��L��K�hBB�֧�!��/4x��3�	��Gq�OP��]{|��z@���d�qwHfѸ��Y����b�Ip����E����[�y��"��S-�3�����XT?wɆ�ehRr����R�� >�LD��<�r֟���������=JL�Q�X����):�%�t.E8�Ťs�rh���I�Y�������o�x�S���[s
��Z�lo61!���`?4*jA3 +�<�"������c��zM���Q��c���N-f`}� B�qY����HyV{B̝���/V��5������B���U^K	̎�Q���T������An�o��ET����m
���"!�����+�I1�����	�a�W̳��ksJ��ߋX������ަ���g����U��7�O�N�P�u�/Q���k)�҂�%vu�1��	(��,p{U6�4? ����N�s��j4�-��y���e�Yݽ���k愲��g�{�h��I����kmo�����֕s�✄,z�%�� q�]��2zw��VѪ��Y���K�۶�UO�{��E�g�:�|`��q")h�r�?�j��!=� �"2VǴL����I4˳Ri!.�P\#e�kY�~_�ro�ބ�]>k<^��T;Ar9��˞E��Z�o*ǎ5_.U�w��|���K"�����@�o/�Q����̙��<����ib�&W�E���Г
!�8��x�ʄ�Kw����y���$�$�y)@r������j������g�0�R
	��7n
��s�ݜ@�zن5��e��EsrɆ�֌~t�2��Q�1��]����ԗ�2_����7��c��sD��G�1�x&�}��Mi�b��tƭ��� E�R�~/6�E���F��*
@�ck���Y)1��k�`��ejW�����̜G|*k]�":-a��m��9�{l���ɖ��b>T��3�T}>�&�>d��)P� �z�D��J	�hP�D	��H�����H����z�O��-S t��D�`�c�W~^s�"�	n]UP4��+�O����/�V��D>
��uV/���u��?�G@,a�� .'�e�n�޾��t���+�ŷ�95�d��������^�/�S�J����@�sQ�����t5���F^b*����O(��s�L�#m-��c�c�����Ӽ�,�Q���p�zÒ�?#�'=�pi͂�W��2h*4�&yr2���U q@2��	ݿ|��]�`�ڠ����$��S*�n"�DZ�@�V^WB0i�a�M�\.��l%`+�i������/���f+�-��nh����m���P*��#AW��(I�����v����ԃ�m����c:3m�I���6k+0�4Xt�ְ�f�>��Q�Б/D~�j��=ҵ8C���h�ۈ�<6'��^c�p��Q�o)�/a$X�L���MfG�`*��i��|Lsp�G����gE���@����ˤ�IC=�l�E�*��_��X��	0��jK�T:��/�^� h���A�Ӈ�싍B�г������u���牾ޟ?KSWא1 	���z^6�a�S��z~Gt�1�4&�H�5R���<|J�	w��Fjꏉ0(ّ�!��z�q��Z����`jsNɭ�!>L�އ*D+l�uW��J��l�F]��~��vΎ{�댏n{�$h�G�[����|}�5���#�0�S���;ĪŇ� o�Qt�tL�D7���gA��
O/G�ܒ��_�4�A�d+UW�:r�i"1ܨ���R%F��z�
f��rn�����#Gj��H(M�V0��9,o��[I��\a�N�2+�m�u�E���]-(C6meE�I��}b%�[T�Һf}�9�U�c
�҂x����w� �$�5������%F�`;Թ�m[�U�C�p>6��	��ލ�:��|���m�|���8C]�Ǽ���f�^W�6�V�Ƌ�H�����V*�%+f(��-�wV�y2����2��"�TJ��ӕx�lV]ߖ���RfD6�5i߯7��ζ�Y!ڏ�YVCA�N��(؎�3��m��K@s̈́�����]j�������+Rv�m4ё�F�*;���5aE����=�Z�0�T�a7�El�򡆎LȪA��.��;���x����QMמ���6Ԙy��[����@�l��2��B ������M6.ii�%�m��ͨ�n_�;����W4��� ѕ����;�I>�R�i��� ��32XV�\4��#k��E� ֌�
�84�5�d�TǬ�}Bt�*�y���K�&����z��_�g��.| Q|��8���3Q�Y�]�u���n�hkСH�?Zt��/1�CƜ����9�d�cG�1\Lb��B�C'YI��S�aǈTa��9�B/!�,¼�S�H'�I`�Vf��l�JZnn��\i��q��x>$I����Z�݉��m��-���}�J[" �w��ڵ��1H�8��[��	��=���?sj7����j�2/&ħ���	&�S�M��b���3��'a��bL���ξ|�iTR�s�����f?�L=�Cl��pmߺ^�TyB��?Z�o�I�9����h�Ѯ>VA���I��~��m���ЅPw���� o��jZ>�_أ��Gr��*XL�KE�~F��)�n�9x��J���X���4���Ji����� ����_��Z�,������뚨(���]驉�n�Ǿ�P;���p�F�q�_I}w�<,ۋb�f1�K��LA���.����jVb10�q�o���X0w��r�u�4�dT���d�ɖ��zn�t'<�K (��]���~��=��rB*������į���Tq���9jeJ�B%�/����a���IEJ�=t�����\��!Q��N�#��-�m��I�η�,�����Asq�J�A�D��R�n*�L�)���V�Mxz��T�0���L���+��������ل6g�v>yp�z��T1��a�t}-�8xV�~�U\/����W~(@��2�]��U4�N�/�1�1�Y����5��hn�(Oyd<h����E�����ڱ�+ʐ%�}��DJj� ����-��d��cB��%��Z$�8Q�%�F�y ��cU�r�0�s"�޵Z�?�o�F���z�C��^���3�zltJ�r�a%�������CIk��p���T���V�Ԅ��z��N����'�9�5�#y^�g>o��8�t̰L�.`����\�g0qk�v���0�B^�$`�8OKe�k��e|+�Lx6�B�٫��qπ���~Y�s�2	2h	��ג��ΝN���O�sa(�AA� �L�Pj[Oz
�ű��d���OYڹ���Yf�wU�x��^�y� {r��ڳ|:_��Փ��}��}�ލsFA�|Q vEi������q���0�#0�Dܭ���¬Ɔ�]0������a@x+'�>��g�aE����>��瑳\#���U���~���j�%��mo�rq�?l��z��kS��*Lw��2o3ڀ�LlM����r�^���PVp4Z�LylxߧÐ�]�-#�$'˱Tm�v��-nU�κ��]���PoȮ���И8Ѡ��]W�XI.�t ,nH�-��\4��M�@�������㰴F��|[<��$
U��x�z�ᕣ��Z�S6z��^�/r��G���F.@ �X���DSI�4f4����59�r��L�N|���uA;��a?Q{�����Zv�6�����Ί��P	���z �\����E~t�i������+)���Y��:4�F�����c������*קK�E +� �>Z��2�0H��w��&�+�6�S���#̫�"��`*�nO�P�o�8%�'g��3.�����	���9�;���l��+T1�P4<!��'��9f2���N����&�һj�-&�y�BI����E�_��g/�m�_��L�����`G՗��{W�L�$�q�?L/���яlᱯx�X���s�xj��% Jy�i��M�|��k��Pl_�(
��]Ί�9hN;z��Ֆ|�譃�\F @t�Z�ܻ�	�s�W�iO��!�_�I�}�F���s�������JB����a�搅q�k4:T���`��|1,ay�#>�
�z<�h�!�����+=/������>7�d�_P�$�t5d�?�nc5��ζ�f����f�)pY[��jG�6���\1���!�Q����s�&���S8q��m���@�7'����X�p��[DZ�vB��*�+Je�v ��8�6�jv�a'ǀ�8�_U�Rr��i��Fy�����0��MB�<lU`aa)p�Pf�q�EH�Ȁ�� ��k�E��N���.`��]r��j��<t�V~X߲�ro�ݑ��ݑ6&������aFJ{� ��aˊ��2������m�U��kP���s����ᇪ�|��f�m2��1� ��Uh�)0�J���S���n�x�������xh�G���ν��c���p�Vu�[	L8Jh���V�N��B�ؗ-+��*f{4M�-ڗHoc85&��G�\'Pޢ��y�H���	�g�����SV�+#,��qI!F���w�(�	rB���̴/��Rئ�KZv[j�"�_7�fzA�Z�
U�:�/j���"�0�\:�VJ2���U���d�g!��մ�[XK��4��!���x޴cf6-ԧ���")����/;Ol�H�HcERyL����ˊ�R�bT�� /�ޛm��H'{��G��?{� ����Wg��ȇ��յ���w�F��Z�E�~�����~GٓX�ӯ�@����X��$��[�D�UA|�ռ�Ĕ.�$�P*����W�&��Xr�E˜�f{�B(=
l��D�j�K�	��J�i]J伛@F*�X�+��Q��F�;�4��E1K�f���+��B���ɩ#,��OO�[�`2���4t3���$X��_T�C�o���p� V�E�Zͩ'���G(�����z�U�XW�*�뀟ǅ����U����VW+	��k���ڥҬ�o�bP5�b� ɝ��8����ч��w�׏�\~C����i�(N#��c���Xe�VA��^yV$��6O��X�V�,_/�R�*�/��RC�N?"%�G;�"N�=gz|{	��x��n��c��_��S� ��4�f�¤cЙ�md^���l<ܫ���T�Y���L� ��kk�4��<��2mnVw+���/���:��!�JɃ~̣��W�$Mr�B.�{F�����!�n%n+s�ǖ�G�NsN�j��>H(GPx�������I���oi\lg��eN�dΣ�)|�i�8�5Z{��j#x�	��_���T�&�̨�GK�$!�%��Ze��gd)�J�^��i��?�e��'�$o�r�'W�ib���!��,a����s��u )=�j]Rf��.%�rB���T���	�3�tf<�"�Y�� �5&��t��'�H�� Df�w��M�r�#��
��e�\,�1�2�!Y����l��f^�P"����7۞C�RmOm�~)���%l
)|�c�8�'�l�}G #����{�v:s濗�N������|�L��=	y�#�¢�2ҼQ0��s
�O�,s��e��Jգ:�7q�BlV����/��֌��X�a�~�{��z��H$.�^�_���Kj���X��N�e��H;�y�t�>����;eҨ�g+�����o�_r#b��.7�j.�ĉ^)��:(�к�������=�����.]@<[��;��oӻ�Lt�5���4��EB<�e��?{��_��!�x�6����0a-��M�ܺ��~sn������y���. /Ր��a���{��`#\׭�O�ˈH�"�Xb-1!LW�ѝڦ�Ima��i���e6+��°b�`����<�~q¿�d��2� ���{�7��#�z��&Z�uck����G5Z� �Q�P+��V��/�6%p�mؠ^�γ*%Ļ� C�m����X�	G7	����I��_8e�T�14���M�5�  �������$��tR�����j��(�����������m���!�7ß׶u3��H����
g&Mr҂��V�{�B�s& � ���P^b�}Nt�H��ŉk��9��e����w�ņ���n�:@a�8����ɩ��k7t���wր�!|Z �҄�*2���OHʰ�f9��G]�u�Bz�>���l�M�qgb�K�����L��O��nE���.�J��$���J	�b( �泻V���w,���XKl0ɻ���I�5�U��Rw�~qm��_4C~1�/�䜷�\���z�0��vg�;/4��,�VW1�<�Xq��vU�VGիc�?RB(�������'�[�PQ%#5�1�W��aoض>��5�h4����u���/���L���ŀe�����'^
�
'�)��-�)���Rk4�2	td���O�p���iW%W;�NU�$Nڧ%`��D閾%2}���  S���7X:'eR��_�y*�PRP�x�s��G?	*�;�{�2gMyp.��(��_��R��d�F������T�^�
n���y�2�wl�:ڪvnM��]i��I�-�G�P��`|��n c%��Ѯ�o��7vڗW�J�0V�pB�/A��5�.�[׍��q!֡���4�w�قG��l��#b
�r�>��A0�������}H31�����V�h�Jꃕ�����v�`';�ǭ��������֮-w�)3��ɦi���g�Ѻ�(
𼞷+wh��%�VXI����W���WB��O^�_��Y�A��nVK�a|�1����t��H�;��$�"�?��U�*�U�U��"2����@f|٦h�1��(Ӛv4I�G�DG]������Ԡ��v`��. (Q�b3͕$���{J��Ir�ꎁ�b��ua��r:���o1~Ik:�h�,­��Ys�ѻ$�}߯Y�q�-v�NTz�����>�x`YYqw8(�9^�eX��T;�s�Z@34�S*�L�L���������Ρ/!�#ㅄ��f�k���T��l���6��> �����Uxe2��W�V�m6�W�-���t����U�3B?�f�z����Шu!�[��rxG%���f�y!��ۦP��[/J."a9T1f��'z+v�����/����lu*d?� G[��:�G�O��$x^��e�ZA~�,�'W� ĵ���MZ��&�[�U���t��ʲ�-�\�Pd$���O9C��Y�����<W�	+���ueIm�z��uۘS�&�h��	���y�F7E���nJV�<��n��4�����\b��������섹�y�t��aɚZ��zn��\��`LuÌM�S�P����d�Ɋ���������;���ߥ����_��J�-%�fY}qeH���1ŋ���s�������X��lE%k�{��	Q���߻+���t����ܻ�JZ��T�)�'��:X|K�A��,�P#e��i<��g�d:L���C -���j5b/ ��)H�;�%%P�b�?#WFæ���?�($��g�M�������g�H���Q�̬�ߧ��#�!�����U��b�-\0S�7�u��N*o7P8=�@r�@�S����w30D;_�TÑ[��F���'��o�l̛��ϩ�x�CQ#��d^p��s�"��s��;���۲L����;�j�H��d^�l)C�%å�U��l���X�DO���fCC񠈭
T�u��._�ش���6}��~��j0�U_i`ҶU�R)}��Q��ER�ݩ�ƙ]��m��Y�l�*mXi>�O�^� 6p�8'���_D&:���"ol{!$/��5q(�KF%���8����6���t��v]�'�:���f�����-%690]dͲr-�y8��=It~J��t����7�u
�JD-��`k4B����3
���ݠuGf��CN��y;��k�ɔ� ���Hh�B�N���Պ[������=;��p���ع�����T� �.����9�*�{�}R��u�8�"b�8:�f̵��b�U����G}�Ȭa|@�F@�ݑ�b�w˸�ku�f�J�Cmb�è��܂��v��Y���]�q�q��攽�{��N�Q���ˑ%�z��`�R��="���{����W��ag�����wZ=�]��hą�kc2�Bt'���Kud��hz1��³L����S)��Ԁ�^W~�!TM
�W����Nk�0�o�����$�j���(g��Űj>���:�e��c�ʶ��V��91�"E�0�c��G� �*~S7��+����)�	nZ��W`�nϸ���g�v�|�t�.u���+Q� ��ۆ��ϱ~�qa�9y�j8Y(u�dt���q��/�i�;��bBn`�j"`M�>���e>�׊Dd�����[V"*7S�py�[qE]k�{N�_�o�M�m*T��N��aF*6J��+:�{��ZB�_{bnhޔ�z`��$�R�A�E&�+�u6d �c"�x��uȳ����Le�]d�},l��J��C+�c ��e��x~#?����au���Λ��1�;��9���4,�������ԟ���;��<Fd6ÁQ�.�*5��#M&��_��9�z����(	~U9\vx�	�ѣ������pC�M1Q��U��S٤������x	������ &�k��a1��c�W��[���g�nnm�a�X�1jϏ��b�AP1A�F���L��pf��@�C�C{��x�9��zEJ�V�?n�E6��ԑ��[�W)�ˡ�oq�?��{�v�e��1	`���������Ll��k��cl&=�j+o8:mg�k�4=�W�Q#L�7�f��[p#�I�U��ݢ�DӨ�,��YK	;��D�)�t�����?9΁��KTa�U?��,�Ǉ�?� p�ɑy��#�'*湂�h����n��1h� iz