-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1o+b7UloFYH9N2OlBEPI1mwTOXel5LLJJFX+l2M9hNWusxuBE/h9uGGAIr/cecVvsdGPu1MlqFIn
rU9KPiz2CjkYD/gIiccrEZUIZRot6cDcl2qT4kOEu/g2pN05LVtbbDU0sghXynHxMt8Xv+2Kvabb
LDPDcUv3VEKfpOYt9ExO8WEMHK8EWjBkNO6zpW+oR07A5AwGXY41w0Mp5JkYTHUc07wywEV/B/fr
57JaPiI4aEIygBXbVbF5aKQSOxDEeu7ZddSuYgbimKGjZH4qvAk0ZEigk85Gj6QWYrbAGIRHBL0M
aUbep/DxXPibIa0O3vIq6pudhKVqDcfCjEF1XA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6784)
`protect data_block
E5b7QhiB/6RQnrw4bAmigPuUR5Kq9JuHD3B3/53foz7jVZ7imtWo+8yNHfWLXTqjk/LpQ4VVqr5e
8W8zAbeqbZcPc1tVDvGvtCeMv02t7sfTdvSIsJPAU8uBUVaYENoqpY82fYa9PpwllGWPncv9BJoh
Gc8Zt1sFqA5Kx5rJbtAD/moiCTWhu8MA1IA27Hw3cTGVO0GTMIPfskPmwJM9rfUyrZAa4Yfprcb2
OZDv8ObvfV+cLWmyf4YwptqXX63STFuZUEdt3p/WFYsl9THEPTHB1jP94WNiGCmSSGOxw7EWrMNm
fYjCKs7Mt1e5/2zVNB8RYBNWu8/xJMkWqAztq+sz/iGjGU9tnHVHSfVK6wgOLWuzqqMfYE+PzWuK
GJsCWIx5f6l/rQ972JU6A7Ifs8Flg++PJ2M2EOM8mwlRbmPUOljqBw45JLi3kiwoIji7eqerxWUm
cFL4nhk5VDre408eEfMR2iVYwei9oxtOTviadj/xTODmefx1YmY6EjsGyAHWLyK/ihubNuLwn+c8
XhKhNYtOpJyare7tMps+6D9lxrvAwXCSpnV4nS6D7BkQlQHmHYrNBZOWVyj9RMb85SzwvDA5ShDK
bTaz3aL26NKw/09xBpeEp3yZJyblcdaWfwh4PTSA/lKawXe0wBa85Tj17v/ZzjxcpStqusnQL+14
fHhMGy7l5TqHl/FZpMUFcP9BQvuQ1AtYCYhBehWTxgwpfmQsIV5avH14KTzKlpMyhtxMzx+HrGCl
nBgY6Xsc++G1jPLa4roTKIsndfTpQE3nLgKwSKyYs96XQaB5E6MgpPEUoA2fQSFXjbzCoHVDRTT4
IjIFjBxK6XbcR+zTY+IPOoa3tgPoXiJdFYRSXeBoUBSpheSPhcRjnQuBco4m5eLlYNdIc+GSw9MW
4G/VbwpCSHPhtPGxKc+yTZW/DiCMBR/3qCEwFQ3uCxjOJA3b80R5UmE0AKRgHYEXMCxHauF/aTpm
epXDPrfYCqJAXWoSH6PPLbz69mI39gFAZE3T2Wjb4wJtS5Yveot8+p8J1eVtCX6txz2H3aSkz5sz
uV9fw1q4WGHP/tQVGLThh1gLg+9VAM2pulwE/3Ciwx6RZESrObQo+E17H4i2UO1d4+RDvUBXBVH9
9MmsBgCZs4n+p4XuViTEjY8Qt7KVoqK9qVXMuZYIP1Sh5LLCc/7+05vF8k7DCbntWuWHtwo+ZXiu
9xqklOeJ1tw429dCExTFIFzZ5RxurF+FGuemqB6IfELp2WCgIWBDpGTrH+WNkZFolnP+2HUMy2u/
3ZdL1xWQWb6FNeA27xSkR/q8oTQZZtEuPszYQaQYhsbfIW0h9BwBOxQEK3pC3BSXmut3Vdu1fFdZ
Zo1KhO5ZxfrdOryrxLdXEmuQcn7nf5+uwaN6LQaQ3UEPcVMNK9RU0FeRFqPa8O3RzzbG1j59PtVP
GCMKQXP6hWsMDLIK8ToILQVS1lTzzpYSf5c0nX7tQkB0EpARROzx8s2YNiYkg+K03TqH7IWQB6hZ
5aoyoC+YIYbe2YP6u4qUt+0zZ1kuPBjaYHndfdV3JQkj/ttHGYfeVypwIntlaKQZdGGUeXJhclaI
G+u5Uj0Q2CUp19+K6JMCpynyT/U+E6KMj0z8efkm9toObn5JSWwb8iec0PyhtHRmzdrFNFqXDuLn
NyG9L4BbNf9zMiRug4vbiYnP/0FlyrNbYV03KAgoLfRjgFyyNb/V3/RXwimY238+el4nulO9xK3v
u1zOoopXbj+4/2PKeZNZvJd5dXYMg/f3Rqt9JFhG8iTDi+T0gGYr1xKxmcT1Xbe7HnrcT4xwf+t6
nNpDH8H/0PakpkEiZNCnWw+oolt2Ap24asvPvioRpaILAuy7NhkBoyWawHbrwG9s/uMVpMCDv4nP
Qd/oH+t+7MNPhFxD771JtIHFA1VB5Ym+ZoTnrUVCc0Ivp/Pv2KrzRzeAEC4LAVcGu39MJWdfqxr/
6Ipbeyvt63LAEx9b/ht8dotCtQ2GIXlPtLFZ0apl3FZ8e5GAbLRKHEfqbNj6foThItSMwhUKhNxx
4ViyvrNHCjORh5HARqnUy0EiQv/2VBggSnphjPVIFBSwaNwCryNufH24wJm/owHJ29H7x4v0+zUH
4vRWQlMx2VQQm6urNMIFVm0AD2Zjwh2A/vsgY6am7ESk7SkUlpL6ChpAG5egiXCp+6U9NmAbx4qu
IgSXw65LCQvBsOA96T2nhMvYqUEcVdKHfCdIwic/4Te2MrMWuxBdiPHEhuxGoiQHqlqAu0tArN+f
k0bnINqdW2XqmFnPb51/jQxDJmXtLQnLSkxepU3V3ptlFVUSIWs4T8WFxT3Bm/yoDWC77KZyshqb
8NnzZe+hxqD77fTp6Ed0NcqcvLzbWChIj6F6mQZRS7PeYfIcRu800mN6PYlTHnjT/OJ4ASJgNmrC
xh8Wq7x/gYaaDC+go9qqr6ZsESLAbza4vUwy2mlG45DkaItKyfQ7DqHpHCTWKOkTGNVCGfYztc6e
rR1++X7yB6xl9FE4cT+cJlTOTM5CeaHwCOSNllNc0GdFoXlhTH3Z26gdPDF9wh19iXnWGw86/7Fc
6BNCugBd5dzmbJGdoC9ozIJkjA4SsLbEh+UKuVKtwPBvdDX0ZlMYpXkVwtlOpnlaIjIRuMzT25lB
7cwjemTYGXFdwO+QSYAE7KkKrKb5bAffYKybuuXVS/FyDj/jANX3injSsThou/eG+vXlaUBAyI7e
iGRo9apVR/snFJybq9oVpKQhugXvGt1QwhSF/zf0ng9nntx0Hk611pxq9n6Wtt0kgHQh2SN/Pvy7
qy+wdAoUh8q/RuIAkYdJ820fTiwJUUJph+MofMRhcO7eIr1EtkES6zGuhcwnfnrcVXVl+zJBe0X4
eMyZuSJq2UHewKbw1RHcl00Yuq+Zox3ENNoZaU0ngEzLp+TZ4CxyF93HouUPAV2MVko3iV1Padg9
IRxLCYFkF8IoOpNSRNgbUJZ0jmWHID+H/oihC2+GBKpNElQdYIEHgtlDz2HQd8obux61fgFbr7Ba
Kt4IAYuDLO71r2PYYgJAkoNWWScy2CLUOhcjLvr2ovz9i23//reh3XjPbQtJWjVJWuuNbX/FTjIQ
5aeaohepbvcJQWPvD0gsUPrggQVJEC/le9+mQjsy+l8vA6GZxGK+RJ1xoHJfn39QUR6fqVsiEqYL
dKxM97sIOhI24buV7AmZcnOqq6+CVs9V3DgHTQdfHgDKzAoBeE/s/7/PL/xtUEGtcj4yGuRxEy7k
ydwPdWXdFyP1H8Jz2BTLOtNsbXOjs5p4rmTcZ7TK5njauwum691CdGGK+2/nd8lTJCKJ/kEXg9HC
FTmUf6+t7AH42XXyel4kcHJ3OZA1Iae/kxccskU6gTobUvP+vp/EEU43I799FiEAvZXXG83t93vd
OfbNryk99V+botUGA+vIc+f2yEFsh+LtrWS4pC2K2DZ3r5gLIqWNvOdBd2dBn/ikEXsWKBrtsa/S
K4K4LJ08TJfhZmIYgl1haIpuGrUZpfg0Ap7s+cmwb6Z0NlWxyhVii+AbM6couUmq699TsJEjPftx
V80JownmvFEEbZpA7z5mpzi3brnL1iEQlA+By1UJssYFY1Td8kfYe1w0MZf6rcbVqsrr4L41TnJ3
Iij7w//hZarU62q9wOChOP6E2e8/xx3LpPJiwUxfD958Hjfe3Q33aNQM6hX71iIcCCqQkmy2d1vV
DBQqC6bETY0pq7G4skP/6LOYaU6ROPdrbrcBgzLrDem6cdYXOdd9pQaJCnBl09Z1XuRmhyONl1ub
myhHzLH3J/bfLqgAQ4PjuzeKRRY1SsXfKX5mFuIq4jUqNZG9fHO1/TigWm0dRHxiz4HgOiu3W5hy
HQ+dMrn/OLIUm9mtF5/cRasvqoLJ8s2MTMscydlfcipOqiSiVqNAij+uSppjuOJP2pLFCcQwBwiU
V4N4w4rAg9LCiZ9dbAgl46U3GJ58idLfj5XLWFhdBk/eSTtTqnwTcBZn0G7yXAHF5vFN7nl5x/AZ
PxGaay1U7XX65nkcz4dgHp3rYd2dnv90H0UKLLv6GVsdCE/Kb+qkqiNbTmETLGiwbCILqrXcZDKF
yhicDpqwIJY5YH3QXO7xrbP9Ev5zGPYrlUfk8/IEGEQPEE4gsVRq4UeLE172n24XTpfI2cZpSohW
haKUIwlXruZ4UnZ7EjpM0s++blH6rjuM6FXgC/i6RWaP6HgIer98Yj2bPWg958Yfgc5RpP6uC9cw
qL5nOdFR/v6LtL8sob+WSKUo60zqI/Z//kumgcOfEvR1W2YPCq99AVsfJObYozM+sjtZEY4yD12F
5yjPmQ3sYt2ezLftcSPYgNUuiOHBuAZkUR7skoNnkhooVbkdcyIcVdC1eNax8b7sROgeXZIaZt6f
hJYa0jRCu6I//Ij6HD6iJRA64OPqGRbHgN2TXyV2bs5gRk4OJfIwaiYbiUOlW1T5Zpe+ubK08If9
Pz7Snf1P0jd6qV5DVHBCPN90OUW2/YShFyPwJEsDP8LeSV75LI6B28pTqoOs6HOyt0X5fhj5XBNq
LLXKkUZBGzMpnPUyKSEUNGHxOGhEgZQtewaoFEMPzgo4KXbO/fWz2LO0B9BoTqi3JHJc/LgthDyr
buBMi3OxFDaKARJ5R2Eug3SwBjtDqkAPbjB4XeTmPsRcIhP7Wd06O6SVvfIx8YTZecnSv5uLEKPt
+tns1uMN6rCfy6MEvRxyUhlFdEP3aD5KW/RAXtJHiviz8LBNTEBSnUtGW22xZmGVPSiLYetcJYdu
43FkouAe9jrSS+KNIb2FWW4B7vRIb5HYKmVtBISnlad1mU2T8G50EtIEYK7QH/jS6GHMCbl7jGvn
vaPJ67rLd7gLj8IdJ0n9TmZkhwkcb/kaXxAsxJI4ySVW3+rITWJEFg4V4wuh+DYJhYs4xtfl5PBL
SJsbXU2pH/rjx3wvccxsIESqLiOwOl2HRYprgTP3CQJRctud9VDX72VBS1jyMITNmXjdShHBmNwQ
ax2CFwtTqNUAyhiO+y9u2Bg1SD27Iq+QDCSaA79SGfQGBtMsmgQQruSVuR12q0sJ5t03DaO41V2A
OTd3w8zM9r9rdALAcZOkgAixRS0fOVJWJRVP4xcE1YiysRroF+ZhV3NIZzogZ2O6dpoFUGgyxdR5
OV2IQgIpSoneWAZeVT5FX+9nmxqWbtIBAFfv4RogPeTa8X1LGY1hR1+GrT0CxDO2XWpA0Y4cWv9O
lDSwaunXQEuVnpBZKXxGEf2Geo+aHcR+4er2onEhZBNKsg9U13Gt+MDWFx0vdRMjbUCdxZldvymh
uN7VGfu08YzOY1wmQXVrtdNy5CIBATHsmkRUuctiilcbNSnitOzFVzKmyYqaM4Nom/kClXM43vm+
sXVk13RVPK04zhB5uHNbA5BAj/BY+BQrzVRiAOh2iSDKOkgOtfsOCOFnQ0n02PwznoTlrGpMCckY
Qve9FtU+YkWt4bg2GCzgTwU3ZYZTh2l0P2wAKU8eqfAYQhWat1XmOYhFYUeQjl+1fINJp+7lKkLV
BcUWgRlHi9O2bdVT3Wmi43cAUo53ZBhhToBIpQ1YGU1nz9CpJ/EeOOsBwz901+quEUVZnyLp0UCB
HOL6fV+EUrQpLHYDIv4IyXOD0do1v6rL6DBJLw460vnph3QENb14Gh0i1XluCPN6rILEkgtFE+di
fpSBnxslX3R/L404UXYvpCKTo/1BiNfQn9LzWqreAjwcz+RdFw9RJ4T+/RpwxJxefL5dfSw4pto5
oVP8aOnrx0x2M/0qmZyNlQChtSDqM2jX/EebT2Y3KjhPFtuwqpbWPmRwBMnN1OEk3TqCr8aKqP+z
KP3sxHZaqfMHseyMT5FK521RsgfrjsJXVP10AAxVmWR/bu7aI+0fmL2oOuzYKUANoplunz42pWnn
CUOGsukFTVmhpQPJXaE3YkG8ocvEKAkvuEeIyDHyjOpw1wkyBq01K/HDPQOEiqIJxaij8TmM+8i+
N5peX9aN3C3LnQOExhr6Cs2OBygekPOoPjkGXC5H6+1JA2JCNfcYA9cNFSTbVZKmC6utLsXkzLq6
hRjcCua+7TaJciCQI6jwyNWroX1e84AMVQTnRBkQKgIkvwk59T+AordQ0GikQ479nS5PvUp6qqD3
mEvPeT8YxXq2UCbiIw/GrQEueHKXM5ecIzaxUQ8ngbIZGdCMXadcY8y8q+ppwGG3EL9+T+Ozn0av
XLZS8pnw1gpE7iz5wWAgucpqSpOvbcdgeHzZTzjFLWYeq1Fd0A3C+qooGdI57Sra1fIzahO39dDn
Xt3qaLROcH4bPN6GvIpJIs86ItU+xy7fiCn5oTtQLjgc2hAsJA8tyIodmI4k+M9tLYe+0DuQRf6P
dACbU41zVxQGPMSy2q0VcF1NtGY4fwBSv7OP8JEbBsC5EUercZUfWSsySxpsYz9oqTyhlEH2yfKU
MaT3muYMVlUEYPqTlEqz79+DtbmcwUVmgZgjm7OFgDKMkZusjhmnBlMGGvAOdJwdZf+qQhYuSZH6
y6bp4YcWlVjgI361uOSC/6X2jyHrgQ4K/wg8kxcuGtNtqjZrIHzsfwHhQsEaivYD8V92RqXEupgN
iy2i2z+vpgda1j6KU6D6YyLEjG0ITpBJWK6zIV8aPCktMaG4COBTFusAWPD0e55nHxkIULQzyNu7
qE3+tLexlfkQUjTBOvdPzdHN2F9q3TzyX2tVayslHKbOk2C7+BMe7B3EG1PJ79V+LKLbCOma0ar9
LueulHTpgrbZp1ynrToA7SxQnVVBzFQjZt3U0aKD07a/0Pfph3J46A3t29juYkjAWKK/sgeq5JeY
D7G26fR8I+7yirLDJNpYTJNqMJJqswA3ul5B5UArgeAWRP2NI8J7ebVgxBOww4ziA4O6dEnSEl+F
aNjF78kCApPjSGVeQNUrdkzSLojC2huodgeoFYP1jSEE3YhS74J29Y2agOFYKQvAd+ABjUlL4U15
7f60YWMOQdDR9B3JY/qxEemNtoHylnGdfxyPzu32Q4bR8Bh3N7MM4/CorHLe+daLwNseDhQyXfxJ
K6Er30NjgDjWlfZm6Z3pa9FoBzVLQoocT7lxVSkuc8av1afIx6vdH3TrLuMGIPC8r1NikWCABV8U
KVGb483ilPUgkkb2vuryigJpzlGQEU8jr5U2zrq1loi7VrRAcNRyuuidvF08irUkXE54Vy4xEOFL
eYFb3sjPdF6z67Y1oc8S3ObD7HdaqYTQYFznyKbNhtVN58edndbANhIg0LkcUbA6txdYsVvwK9lC
1msspqRVbzmPYJsDhsnpIeIOZegFBqASqHzutWO2D02HmnP8/cGH6FAjgT3eCPD5t95jejRIZF4L
B5Pzx3l7Vj9oBZWsEj7T83Q2p70Rb7xSUUCoZ9bvO7tLgfzH6KUyU2uXEvboiUQpW7zyTC6P6HNU
YLlOUtt1ooa4LDp0WEqXhSkrpgSI7hWz5C0CpKKL/DIZ7VUMdBTuMU3LhgAFFibZoRBgZPZC9zQg
lIHq/XFT/H/muOFepb/CECw1A/NQAvjd23CSMfZ106uqXoYyj/QlegUQtCXi72m0K2GmNSp2Krw1
kulVslFIRQ4KjWDocrPFGmuxh2Ol0iS8YYJeo2OjrTEhcb75DYiG06v8R2jLVNUzths9R/flyEOx
lxO/S2f186/rGC9PqX/Iqxq7qU3kl3K+A+lALoy9ebqIE6bY8N6YhUfNioW1Au94aOyp/GefsY49
9xDNYMc+r+Y9/+tLw6YIiO2fGXxaD6Tv0AZxPwxyRqYk591EzY5qPw+snHjChwS4Xodvaufz2en3
nz7yY0zTY/KWnsfDdGYUB1WrIY/Mx7hxY8b724ffmFdctgeDNWhTStSLeGfd63wecw7eUR80Tgv5
cxrJJjNh0IYonMAxcTHbmiQksVy1V0l8dIY5a9bMY73/mTBo8B2ks/wSjD/kh3LTvU9R/d40quDk
uEKjwEuFdG2VzjGpPpJ+N9VgBaCevRnzbyatDKhjgYxSn0pT1bTXenIUxM69IADkAowRpZcuqjd+
9Xr6t9PH5/8VuFEdOa7BPLJ2DlMcbUDvQjU5VYrylqnTUfpiPlbbTvPU/0vJrjccTEb0Qi1d2P9d
HTbYwe8hMHHQcggPe/foKGxjbY742Up73JRnGPV912MST2D8jJfThzt7waUC2+9MoleragyPek67
IUHQQuYj1qzRo6xBkgCFz3lgfSnMtwID2DhVIXxuDWQNP3UG0+8boNFUl5q029s70SLlrzASWaN+
ZADSoLXUu5y/u1sFYaDmoU8TlsXUJTl1EvSrrf/N4h5mgwQIxeFe+jECDXNUl1gHHh/5GBWI8wUl
a2leTvv4Emr9r6cITxuqCC85jqikZ3EnvX+Hze5xm4QQeisPtjSs3VEsGn9R8e4c2JjWadvvRLYh
9GtE5/aBB/GseOA/TaL7TuvbAPtTF9xHkG4WbZcj0OqEbwU2g7HlqWuJ/lMHvDmOqE7/k3fwKJK4
KNGubVwRDkiHRZl7NktIShW+IrCt0Yl8iDZcmXFIhXaZOwoRY4jteK25Q7+FpRjr9nHxdNzAxS75
LpwGbHsdME0DyUiAFZ/e7yblodNH5AEzz9UInbIPoRsefrnlfzjjskAmFM6n3vjFGyQMyoCY3UmJ
b/vZIBBHO+sDHBJ2G+pDsJAkIOY2rDybHoi+93qY/OVE4lOEe/s/+7QTaMUNqPC5dutwHH3jSVwC
SQGv1B1qyRjHzjVDkUuxDkCIasZ5uQnPDbD3KFJYgDKuVd/i0VyglvRU88tdreon4TqRs1NP0qBb
3RyR88zA88AocBSU8jTBF9a/2gRdvs7JkE9eeRssQP+tMp4438UJAJEhmfBdmh4YXVqkfGUOnAza
VNfInzSbBOJypzz0xZu9uDH1cWAs/I3XK9dtJpqOpWt4jqvV+HDDVea3h0trbroXmSsvplh4lP+4
3TdGdOGMTjfFIX90wuDHj1XxoYkLd3NXcXKWyPOsD+RuIK2H/zTRVLGVWARnkLkBEBk5T63hHWN3
jQ==
`protect end_protected
