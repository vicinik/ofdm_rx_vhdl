��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��8&����i7����I���ƣ��G��غ�]�=�
��i����kM�^���Ձr��~t���$ ��揢�W"�2QReK��>^5>~�#m�ªUF�����>���w�a_�0��Q��YQLܱ�ɛ]���E��ZC�lo<���!Ú�����g:M�ԯq��J�Kֲ�C�C��-���.�Z&����Y��"~��*�K�1o��阔#V����:�$�K�Hh>����~�{[���6����S��J�/_`�����G։9��#���rT��#n�2M�n�G� b�?CB���*�<_L����9��X���^�9���̂q��J�������Js�
L�	������^'c?y��?=��N��y:e~�Г"H����{?���AB��cN�5��~�]M�16�:���<)�K��ˤ��ȥ��yr�L��|s���?y����/��8-\3�ۓb�L�ɗ{���̛3��?.2�{J`d�����vj�4~�v�B�nP�z����n��4̳�]�� q�H�����V�R��3I�Q�����ͨ�}�(���|
��A!�n�j��q��y9`�������[~�oV4���vi��]j�	������Zp����O�:Y�G'�����f��m��T�˱��:�dm�C9��s����u��Q�r�豜j���c�O	��_S@�	�YȒ�ٕ������;��h�5�]}�U�*r���,�4
k�� ۘ��I�r�3���[�
d>��?�x���ǉ��Ѩ�pت�~L�z�N�#,7�@Y�;{���Ǒ]#Ңh�����3׍��H�����N����&V#٢�Zd:�w����=�}s�(\h��7`�9�Λ���7(��^�S�&A��r�q��k�9=e�[Q��##�����FJ�7��Cӝ1�1�}?���2±�Q�zP�,+~���	9-�&�|&��Ji@x�۵%.����Ȋ&�_jMQ���7�?�����ə5$�� 9�� �)N�)"�����v6MDo�,�@�̘���,��k���&�-v�\I� '��k�7�(�;^�]�do>�$�F!#�m���휬"VRݎM&�C��6�P���gZ��<�ߌ��b� ���n��<ޛ���(RcC�����G�d%C����. ��?N��_Z,�3wMhQ����[t���2B�t�D�OO�"e2�%���(j��R}�E� N�,GH��I�~�9S��*�;o���ST�kŃm��|�A�V��nO}+dlӄ#&&ʾ(�~(i\Y1y*��{���o��m��>1>�0���~�.
g�{X�Ш��&��BB�)�ST@(��dQ��$�^��k&��Y@P�q}&nQ����ǑR�Xy��>���}]��&��X���!m	��>�f�[�34D�7&&o��'P+���Kt�U^�K�oU��1zR1�Ն\w4���Lgc&ϫ�;w%p�H7ؙ�E`�$�*���bl�����w�n .����7�$̈�f���ޔ}y�ǹÖ�﫳�d���L+��Q����8�$�k),3H"���8X
s�v����m��GWAtT��E��|2��w�
��2;):��5�Z-q��:���*��B�y�Ӳ3:�^����o!6�AV��S+Pq^���0���yN�f<��؏�f]����YO�hZO���Z��Y�:ec,|f�����ͪ����s�0��P��l���
i�^�x����C�̩��h�R��BW��P����y��3*BJ��~�n�m�B�C1��w%rt.���5�ǧ�<;�kx5s߮�LE�H�3�1.� 	.$���a�����ҕDTF�36瀨�(	"��ƌ:���͕}��1r �'���nWY��eB�q/��6��|TŗD��+��
�Q1�I��T������$�z���jw����V�wagSH*ʦÇ�c�9��;��&�V��,�Q��2"�i����E��(����?��İ!K�h}�/�<o2��G��:bG���b}o�Ƞ
�/���"[��H����:_�����5�]Q^�?��*f�m����Za��s��E���?D�^��7�S��V��_QC{dr�/	f,�-[���x��)v��6�x�����hN�J���h�'��|�^$qs�1��������p;&�͖��$u�^�%�yG�� �'=Z	A�u�o���������bˀ�u�$̫j��HL����֧!��^`�i�а����feΌ:�!�5J!`v�QX����8?T�Ď��=*%�]/�"nv�M��Ø8{�&��R�Ѣ�q�O��j��-n�����}��d}�
��g>¯��%ߔ�q��=���o�S�������e����)�2i��t�|�|a哢]���  �0Pe!挀��F���$r�9�7��F|Q�ȋ��9I$�	Bs����6��V?H[^��P�;Qj�+͌;��u&�$�b�(�����'�Fj�PY;��
�p��)�<��E�/@(0�1���0�-��L��d���n��&~�9��c�~u+�Y�`�0���`D����P�J�.�-Ʋ��7v�JJ���9�Gcd$Lt1/U��2|�YRJv"��"��'��#���ȿv��< n��?�Ҁ��o|���K�^0ժ��l���q�l�+-%�6�R��/�-��6B %�Ŗ�dg�?�o���E;�/�i����"�*YϺ$�N'�SN[=�Ƥ��jረ9n��CIV�����Y�Q�����E�/���k�<����j| �(SS~���Nu�W��\�f�t�Yx!� C�	��P�E�w��D"���:�?�^�2�rB-/�J�T�p��8Ξ;Ĉ���l�E���9e����o���WͲg�
��<�ۏ��p��^��&R�z�ٮK��ub\HȾ�'�ѣy̤��l1�9v;`��0� ���㬘ܑ��uG�J�� 8�U�Θk��^��8�`�d�.Y%��
jeTB4�&(i�kc5�\�9O�Y��4`B]5�A����L�`����<�\R���2�R�MML�mD���1-���)�e�( S�ę$H"S�j�i�V�aLэ�N"�6v��֭1��\�s����6��B��K�G��Hr�	� � ̝Z�$b�-'�an�e]���2s��Okp&����A$�z�+��d$�t
f�jGI}�"�P����:ru�S[�W}�I��մ�z4�^���Y�+�K��~�x�T)yk�k��\�>b��]c� )�43�D{Q�i��d>S��* �N�{�_5ᴠb�Y�c\��CP!m��
���PTWx���H�����v��񊀻�j�:�q0����Y�D��)��/`��AÿS�d��W)��PU�8���)_ #H��q���sH>5͢�,]�}E{l�p�:���C�q�>*4�`\@v��;�1��TG�ѕ��4~)2>��5K�筶����&q��Hl�E�'�PO��Y�%�� �<�0߭Ĭ�[Dp�b���a%�iX��R��+��=1{.!�B�n�3�w�[�D$�F�jT���8+�����ݜ-/�_q�x[{���i�9*$T�4�m��Kk���iS����<ư�M)����SA���y�
�_��1G����|�n:�(���>����Zy��!�	_&����#��;Dhg����S�7ih�ɩ�K�ѵ��(`�#}��+�H:�WG����K��x�
b愐�.�9���©KC�)�H�U<��ZPEV~vi��Z���*����b0�}������L*��GW#��T�0������as$�3���b�����T�I�wV�:�~�u��[A��i�R���x��3T)4v�뒂
�}�*c!t��GJ�k'����4��1@�H��v�ڋ	-%��U�&��u�t�ı+����9<��+�4A�u�A>W���!����"�o�������ܡ]d�J����ϙ�8}�?x0~	3D&�?1��U�h�	Q�I��S_�'�J���G&ڽD�n]�����C҆'\�R���e�O�� ^!��"6�[=��j�`9�b����4��?n�m�kp���р�wVZ�R#�|��J�v�RXko'38m��V���>c֙'t��tIn�f���c�v>��,su~��C�X"D��J�����(�9=���VՎJk� ��Dz��ԄO�F�$�#M�+*��Bƛ�;�7�'�Jm4��s�����(���8D"Kî�	�bL%���Ť�.�̈���إVR۩��)zF2��3z�AXJ4?�<MPY�"N��9Av��f���Bb�C�rC��Z{�@��^+Y3k)��z fjË���)4ֈ��s��v�Mҩ's���WO=1L�y�C���A�8Q�}�9=��a��=2�3�^�ۮ��3��ly7[��}0`V�ֈ�^�̿�v��@<^Hǩ~�h5�;>�|����n��P�����ц���BP���e���f��;�h��ޘ7G/ۣ�t/J^�?%x�=��F�"C9>��&=��,G�����!�<���ڜ7�6UR�9�,،�O�Rg�Is,��9�7������|��̋�f�ѨJ�[reҡ��,���G۝,�0�����y�wk�?GJ���Y�aV�'�*d	�����Փns� ]�_����3�v��[
��O�ytk�C�IT	��l�6A'�fх?������������*�<}�r��� <��E��q�0 �+������Meˬ�TN�Deq��v�������@��]p��[H:�t��l⏇*y�q?�M�0	nmGkZl�#�In�Q��0}��"��RCp�]�F��/�9�v�m!�����IpL����;�ޟy��"X�����1�f1�
�S23ojj��X)���25	|K��P]�h�<���!n�ƃ�dڹoJ�����:���yH��F7��i�g7$���3�K��h�x����cɑU�#>�=ߨ:WM�H�հq��'�M�1��q��%�\�A��B���W�u=.主�9�[�~�c���fnhD��E6��v_I�g�ˢ��U�¦�"�Z	�3�X� ��7���8��fўv9�6L0��I�)4y�f������.fy;c�^�)-Q�߀���ӥ�=���.	+z�Q�B���D������MϬN��''�$7����od��}}쒿���V���I�랟~��ڶ=�z��pV<e��J%�QX�����a�<!�U��x�f���L�V�jg=�S�lLG�4�r{���F?6�:}P�ge���fw��T�UXz��9[�ǚ];6B����[��^m��&W���|(w����T��&G���z\���і���ƴ��Ѹ��U_�/ ꬍ����Ⱦ0��x�x6��n�|�� ġ:w��=�\D�:>�x�.|@�B�r��p�겸lG����j����
��ו���(������Jj:V��P��|C&.����[Fcܟ4�z]��d�YҖo
�θz8~�2�%�ra0
\��7~,�
��)%(���^����7��pn�C'ƞ	�7�)��e�Wn���	yd�
-��.G�(����bH=׬,4�X;���*TW}A��7� K�j��l�ܐŗ��e�o"���2H�6�R�X��ؽV8�����:�� � 3&����\(���G~x�m��h��zd+"4���H/;ۉ��a�허�7����{lN=5���IM�>��o��.�v�^����T5{�������p?u��PO!�@��K�����,[f��1pȉe��䍢8躱 �l�����s���s&�ɵ6M��>��u_�IP���Կ��C�\9�y���P)d�z�{�	b�x+A�YC��$$)��ң*�Y3"B�Q��v!�͏�������$�1�K�I�iz=���b_=r8I��W�����zi>Jo��h�.|DݰM/W,�Yn�&�*�}�����w��Cr��V��D�/�5a�7� 4�(��
�}+Q2���=>�&�B�6_�I��%]�-4�BʣC-�2��O�v�{}���LTN:MR��\��	dV�=�N7��m��f�N�ϗsoYh	;%r&P��p:��S����k�|7m����ƌ M;˳%�*�
�U�ļ��a������O�<��G�a���D�ڛ��h۪jRDM�e�����ab<Ku�����캞���{=�(�̀�"!z��!�^[L�	`�e�2�w���(I������z�19�,_(t�y��+�a]!�t��u�77ن�ڀ��4Lی��䵯e����6�gwX�_�?��j�j�sbL��m�n��{� =�}U�P�I��芅�
:A_5@���]��5k�O�u?D��Neb��bb�e�a'Mg�S+C�`�q��p����:�0~{�3�/��4���R��v�+�C�W,~������6�Pn�4����ϧ���!J �RFf�ÛCk��+^�:_:Q �Ĺ4!3��BO�:E�,����4hZj����6-[�K,��<6k��r�!ꉙ���oL	��=��Kf�̦y�˙�2-2�Hě��ꉵ��}���ޒb.X�s�� ��5NSJX��4�M	����<��Qx�+����ʮ��c<���q#��	ǃ �4P���pj�a5���3+q�wL15���9&C��TN	_i��(1��(�p0��U���i�>����a�{���M�<�+�,��Cg��oG�����f_�:,�՚P��LK\�촲��9�e(2�.��I�8��1�����b(�`��xezzQ�;u50�k/�D�� r���<�_���2 �s�O�7��.�I��_�Q����<	ѕMW��g�xً�դڐ�p����jnI}�0��/w�c�?d�@M�}Aꢴٔ"۾AUC
�?��=�hT� r�F��L"���qt*o]�=�x>P�S��ޱ�� �͎�ѱ<4��	�EKi̷S��uO.𗌙 ���H@l��woZx����bt��$�d�2fz*�>K��4����q"c˓�]�M��3p��p�F(��z&��>jN���Z>�M7���@���w�ً�ܳъ�q�c��1D�^it�l��%�u�u�H��@g2T����T��"�U�^��v���=�~��P��U�S�,�$���ٕL���&��m��aL��p\�H���[�ѓ��f�e��p����ّ�ŵ�����a������RH�2��d�&ؕ7if���K�����"�XO���pxe��4���#�j�]��`�у��d*�XO��㥊�����|�ܿ'����+��H�2ς�,�]�Hu�w�7^�����~�I�q�O�DÕ�.GX���YP
 �Wa������oGo��t]����J����J��:W���fGY���t�d� sHW�gv*�����5lA����q�~9���:!(�9�0�z��C�l��9'i5ȷ\xR�]H%�������y��ȄY�GW����ߗ��}K�o&T�j��V�з�����6��) ��˲X�u�̚J;�@��pB�K���A?h�3�{��%�
ZTB�{�4��n>�9Ŋh�5p30i�l��q2�~�!�Ti@Ns�.  �i[^��ͷ�R��'���o:�`~�VU<5}����=��S�.�B��lFJ�g8�s�j�To�(t9���|���]��l18�o�>n|��7�P��P)�aq�{�6.ȶ�����6�UO�n��%���Ȏ0�Wk�$.��Z����nVIHDx��UR�;���]�B ���9��|����"ԙ�J;P�犊�×�J��4�/��~�m]y*u�`7����(
@��