-- FftWrapper-a.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

architecture rtl of FftWrapper is
	

		-- Components FFT


		component fft is
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			reset_n      : in  std_logic                     := 'X';             -- reset_n
			sink_valid   : in  std_logic                     := 'X';             -- valid
			sink_ready   : out std_logic;                                        -- ready
			sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			sink_sop     : in  std_logic                     := 'X';             -- startofpacket
			sink_eop     : in  std_logic                     := 'X';             -- endofpacket
			inverse      : in  std_logic                     := 'X';             -- data
			sink_imag    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			sink_real    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			source_valid : out std_logic;                                        -- valid
			source_ready : in  std_logic                     := 'X';             -- ready
			source_error : out std_logic_vector(1 downto 0);                     -- error
			source_sop   : out std_logic;                                        -- startofpacket
			source_eop   : out std_logic;                                        -- endofpacket
			source_exp   : out std_logic_vector(5 downto 0);                     -- data
			source_imag  : out std_logic_vector(11 downto 0);                    -- data
			source_real  : out std_logic_vector(11 downto 0)                     -- data
		);
		end component fft;

		
		--SIGNALS



begin


		FFT : component fft
		port map (
			clk          => sys_clk_i,
			reset_n      => sys_rstn_i,
			sink_valid   => 
			sink_ready   =>
			sink_error   =>
			sink_sop     =>
			sink_eop     =>
			inverse      =>
			sink_imag    =>
			sink_real    =>
			source_valid =>
			source_ready =>
			source_error =>
			source_sop   =>
			source_eop   =>
			source_exp   =>
			source_imag  =>
			source_real  =>
		);




end architecture rtl; -- of FftWrapper
