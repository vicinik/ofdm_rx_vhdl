-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xdsVKWRU/Wx/LfTALR5FtQdZKytgwFMz2d+OKCvdsg3IPxjUZyjwH32URzM74eCAuu8/6kwaMbXJ
oSPpm7gGYFKGxh9lzVm9GxbS8tocrrHPfhV5MTR1luryY/Ho1JeMCBO3mskjzY1Kq1nLkFhTZz+V
pGW44NEUryrxCNRULnTJf9w++eTgfDpTWgiWJagnH4rARtS/4DxrwsyOK6a6rvhWXBPU8C3sXZLX
rVn9caoFYsfFmJKFcFSd+/bdcEy4mz1RFUd36YM/WhPkK+IABd+UENrrdy7uHZZtNjHZ2fOBsu5s
Am2Qg4u45gUQmpz9aqPQaOq/y0PhaYrCU7qPtQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6208)
`protect data_block
+FnJfQpxGtD6g49eAOAdC2OmgHFzE1MNPiKlEUo8RLhUs2Dp2pGD35idn5sKKmBj7M1io/6YbRQE
Y5nov+qCxhwWp5IlUzXg+inneyO9T41WpgqzO2seOEYXZBnNBHnuMCHQbhymQV9nO4jI/cXGrUrl
W5/jGfBjH8pLNGtc9VxeBwVFvRwInXiE9SoEYOiViEn8pZV28ckOQLOQ8zl2VCIG7W+SXLvtiqiB
TBTI4Iz1HPeobC4Eh4dnLZPkWZECpVQLHKDzSw5b+fW+0BSqbnXeZjNSQ41+wdV1V43L0lUULIJ7
/hcSeaDj/wPVopQ37AdRICPf1w4CvzZk9wlU5ylm+xitJBz9nlwo7LPpm8DJaiCzSBNG18wH54TB
W9K8BHfKDJSJUMLvlYSFBBei1CBhQviLyKtxpB2bF7tPYFvp/Xec6iP7K82RhqnjjItFwHvzTn6L
2VrRmgeE5/8O4J0lTT6m0DUlEJuPr1Gfnkvs4vmoLonHma/l/A/9t/d93xw9zx1ppqbg9qJ9x7R9
KZJ7W7x+ApdDHVd772j4N4GWbGMF2VFVS6c7s+ManA2+LQ0XuOwdb1z6C3rvXwrUMhiw49OaDDi+
aozdy6f9TgXgsKvWGthd/tAWaclirGB5y4POBFDkZ2sNm2dh9BMsyapxn42mIEjVfKIERta7jEJU
gIUDp2ZjzKn05XNPw6FiqsZSGNitY8IryKE7HfeFcQW77nu/p7e0AFMjTdgi0wyWW/GH5IxC8gpZ
du2grTZJkVmwBugCxlL5SumhJxkUGbVPsQuA2H7Rp+28sp3vywsXBOWlf5qcf+Jc7ktGanmtwqiF
ooLd20ZevFgLw0DDKCX2+MvGa26aFFSEzCfxHyrZ265LK9JZnbBRbqE1m7uBEcbR97GVxUXcmy3A
E4Mkj+fT/xMIeMCWznzzUTbkTQyf0Fp2eoU1c6NA3Gzh/7M2CtcwgnfPaBHtDxPUjksmHPoo59Ag
HDiD1jmJNp2i1how1FLIx0aUQwPaIRpB0fu5Xtci3Xo41R/V/tFbYEdQQem1ZjS7KffcShWtH7WR
rN4pKVkvDZiym62UbtQyZe9g3QH/+axHIAS1dZNqRvu6v8or9Lkh97pyZjIcGdRJsQDwYHwC0+NE
gBGyRy/kD5SEr0vEsnq00/C/9g98R8vkDR8DKX2kSph0iHXD2NhNThZ7jqPmjd0yPPgAcgLm85ap
g4OQvpPzKnLzgMp0I+6gDdsrOVabfsR0mBwWwvLSQ1dqkUvcbhR9TBNEBi833UbhoyIa+iJ0QvOj
YMPekFKUPClQcFnrJSchfi2K3CD/4jU1Khd99InaEi7ywQrnAdDv+0u/DdOv7eq2iYNDgqn2xFV9
a8DE3W6kHtiDTQgFNzJwcgJrklNGFit1FYMBKdJxpVkVQrwd9UX0+goBRgcDURQSyW2G6ABer0gC
LJCKxlyY+XhV8Knl2bERn01lcn0gVscKHr7XCsz+a6055MJ7trM9Z8TzP/XGEhpKuz/3eBtFWKQ4
gVMhv2DF5kjlg9RAvGsB+eubNoOOrAbJcOqCh35Tuyt9fwUIw0M831mJiA6j6n3g8LCWw+eUNnhm
4a5rrm1HHb1aakQsfG+rLZNR5Mq2kDpU7f6USZlNMx98vXUVuCdLY4jLUORDdgOSM3/ZqjYlli+e
Z+0BhMrrbgl3eo8oO6UywflYMKZhzUNnDKC600jCADfClhf/dRA71Rm3VLY7I0m6OXpGsQ4AD6ZY
0FmUycSM9AEIa3yfBKdqSzxbKSgj49py1GlH3HqwiP1m/foyoBad2JEa3qVBNpMnvRtwfjV5ecT4
8B/DKUTL6xeIJJO1+6KrGDCpNiW1AQ+ebJg0w9+rNXtzgcrZBW2oNtyvgqCNljKFgZ8/iC2F9UYD
qkYYVTlJHnDHONpZiztjTVk9pZcJNpBLhW+xH8z+JCXnTXnJlVrgTa2XWK/dn0P1GaMaLfn3sjil
mZSVJ/TojE7aLYDvchWr9ogqvw5RK9NeQcYY2jHZOzisLgcfQ8DzyAHntIu/xI6qzLoM8BOZnxFF
LB2HiM5BpCe4KndG5Tfuf7UhLrkV+11rZk59xPQu9NHUNo/WTwuahVufDpUFtuRq4YctW2ikwLPY
KFsF4KT1b4hqYTa2gi0OZ15Cd7hQO407I0LJqrNYktfLCox1ao86FjitI41/R6/4KTtsa02aNIcr
pz3KiYpPWPg8kiolCdDW5fRQGVmZJW2OUJabovbnu4axGtMxV8LAHKvraMETt1Tmi3UlkV2Wp7l1
EFZ1O/xgqMyZ+w334e7OwX3d8kESyEKFis/JEL1YrmnvUUMq8ZjPIsZalo5UBh67zV6t38bC2K0o
7SiDzqdGhTnAb9olYEplaCI8suF2vo+Ayroq1umr9K/wN+sVigEAfOM+CBam3aK02l4Nn/+07pIg
q87AhAxbBLaVpafheOPulREgGXm6cEuLWiqjNot39ml4W7HVfg9BOWrwfkinik/Ky+3bDubro+yJ
NOfNYxv3FiQjT8J3V2OH4AcITcrHrjUrms6tgu5Os0yd7SZgHGW1Hhmna2AKAgLZQS1O8MnY5LvB
n7HiqtgDEze/LhWiDP8lk0031ZICKe0gQSUXjjyxw7uxLVf36WlvzhQcXxwWBVihgNtosITFh+UN
FG/86Krx7H0yqaDNPskhPho987ZSGtoJ5xp2NPWDkL8DFXHchPmKxgAo0/WJt/Hhw0HgWludQsNX
jrQcL0AoJkWL2s9dJwoYpK1k6Ii4Ss2T1bjfwJ8IXokrKGAiEGUnAOeXdZzFIPhNnQ094OCaANvR
zXj7r6vOhiJeV/9y9TyU/46yp9Hl/LsFr3DpnY/mf+0IdO4wFrhnsQCLyINwjYsQkWE1y+5dCEI+
s4Vo1sjeprM8NmZOlJq6+ISecVU+S4iomSJajZoFrRWe4WNJwRFRIrak2hnH86yqJQZg2a8sBHNl
LKNkTAbNpA0KkYJXvFsWY7v4XjlnKcvLWrqObBFIVF70QIfD413ntdp6Mx1YbfrLC06yNNt1WbOj
avB6ygvAJgnOty3Wva2CQ0X3WE6t8ghEgoBdQKgNGbLvhUPq5sHdMZF5lfGojN+SgnXFy4MFlj96
he/+OsKqdcpvfgyR++rr3fGbV4fWtYO1Hno5OOKqALDKBPpxQpJ6yzsxZzZ0+e/VA6yxvPdii/K+
eANA5L0moL/VXYnHclfWGkGtpqlQEp4sGPKM19RzmxdYYwTN1Unk5OgaraQbxP7xFnlgHL4YJDuz
0eORsXJA4X1O4HqyyQA6h/rXx9mMckMY+YBdkdnnPiXeHucxhoRUuy8kFCWWIaSjksZhhRmYwcb2
4Dq6c+7t2DZTFOI9Q8UOsJii9OQtxiNDktck2qIHZbByJkMINVL4Oh7YbRqgVfGMyygOdGiMfEBX
RgwKTZNr2yxS5K/xIy4l/e+dOg35s5bQ3gpZxA0RS+Km/J2+FzxoC2F0zTmHWgyZZb61pXv6jZIZ
4lm5quHa0AjQnFbpEclLrv1T8a8paQg4wElI7ZhOrHk0xRiz8mMqUIx/P+VwhAWUCMYJSQJRe4Yf
zKaAvc98hUs87fH8gbpGV0k5BLOlO3yn2YV5GigzTZ5+TFZ6ZS02HXgANhUC19XTGjPgDrx4gSSf
rYmySHWuTa77dqm+E7ZdyUXEvt77ekX6xckZQRX6aE34GKK30eXH4LqMdy1jM8hTaCgs3uAkknEB
nxq+Q0No57nJPqhw9BnnFoIx59DiJmSKyrdTASPqCpLBSkXOa705HO9BaOivJ+bFOtian7vgPw2I
2oTfLFQYQwSZMP5cmpG4B/DkZHPNIlfk1dfy4DEtMuAcLA/QyAJBoXbgQrkNYXxN6RUR82QDDh/f
2ElYe/YBCzYUqLc4vP2ud/gwZdJ1t6Vr7vN74WqQ14mBwpLU4oJ7ZGRsd4s75G707M/UhfRaKNwW
QBZ58xshxFTlYtr6EyzHlijfwaESneon7U22dd4PYzFU2kfSrP8YnmLmyUXQAKcNflNt6sCUgOaT
6aJD864Tof18Rtb4HVnODhuFZcz8YdaKhJ+tWDbo4R/QgKxSc/e0Qrtz7D7+CbegPzs9VpmyNfcy
5Smhg39e+573+fzyMopQJLyj5j01K+vszK11ru7xq1a6llPgRfRGo+OlTDOC8xCbQ6geaOlAYzT8
ZJAwoVGbTuoZJ/jDBFh3yIK6zeDrMcVxDvvPzHS2YBXLnNOzjMkUrsHtKuY2TBPxgi1mcV9ufuYw
PzRp3hdBtkWTlKzOLRtA21VmXug7P1EsRI4HmZxoGUK9MaiTnIns4dIabO7d/p/IYSyhr8OEmcd+
8+xcxff6XVfFMukbgFndqMr+BkzcuVSNp4v10yB+k7Adb/lY9G4IJbr+o+Q3KXe1CUAOyZ0NIkfu
onWK/ATP/vbqXQXje+dPAWaDxMqZExsKEkIKLG8tCyeM+3B96vy6eE+yamHLTDiWgN3WZwtOe6Tb
hUSqj0+ajmyukjjA2WdbwesJ/aqETewd2QQ8NcpA4OyQjWDtF93Sn1eFr/0BYx7XWSodocceRokx
ez4SOWhlN4fiLcqQusKZLKldb8Ug3oYbzEyrixFeRO2OJ4eEUsHNWRaDyz8RRdc8EiRN6UVTnkna
b/uz22+s8OOJsijXO6VgU2UGFsw1wUQooRO0C+ND1YQuwj6BpQt9xpLhs78weTe/O/hEH5A+EsV9
f2K9qgGIL/UB0RJIP3VP8gAJcWftCf6e1ACjeN5EjMSHvmBkUKcLibgZPMwFEKD90Zv38tObWvtX
L8IW84Y8yTbbV0dUaYvdVLFZi1N67GkISLwEoVOfVnXEwZNTniIdB3nCgAum1enH1jIaFoxJpPyJ
vRc/uWUaijlb9LIdCG04Xq/TOdDcFdeShZ0dtKHh7ccBIK4s/iM6yp+5k9uLkvYT1lR3MbT+l/tA
sWxr1EmqAxVFZsaK8Yu0OAjk7T28oNvptEx1f9QzWFsYS3WHJV7Fimj5CKjKIdaTgyEb/Cj8Jzoz
wkckZSlo1sYTWKkJT1pjH1ojpWtQwsSEkD7e8QBYJ8tqmF/k5YT5tRylXcdMYH7FsUAt6tp/1A7F
jvki4V3lZO3hZId0cAEecEYj87YHXSO7TRiYnjCSYckISx7ThsWxWolcWO4Q3FVNtNHlJpBEYbkL
X0STj1MO8VdVkIxJWrIPvtA3Zny/v/qWMvyvulTdoDQPTVm9Ir2ccEx6dhx5sDKOl89jvtMrzUDy
vOAzJjGXAZ9oYEqUJPQwA23WXeeGbp98pptnDp7xfChiiAfQtwx953FGC0v/nFZ02bVWVlsI+k7v
1Am6zbesh4blOJBJ5GnZd8N+FUobhS2QxIGkkcFQqG81ehAPggmXzk/DWJ15+vNnnjOvYHxYMCXq
DUw1DSP3pBN/ZQ+4ZTn9l04tySSR63ZsqRZzngnbqn94mV2c0xoqlNxKP/PyVm9Q+74vpndFHXaG
WARnKe4b5sntCiJNzJTAFC38RmPQQhuYjoGUMFDZmtdKzKRULPsruoCYQqJTNNaFHKqGODjmjua4
dBPJAVQDFW4HIDR8vprvYxBwoGWbaKjP0XcD0afUnqgAjakyeiRUxSEjSg3YwJ5kzM1XXccFMo21
3jItv8HURYDUm+VjWTIr2hJpJhJhNU41wRyahfz5Wil6KrnkihAChZkWa8sVf/L+ZhAkY+ncaDHA
8aEuTyLxIcwv8HxEgCloffeQAOXO7CU8vl8gZkrEHEdtRfYrKQAf7nwpfB2WJxb4I0mfcDjIb3hX
1+RSP8faWiFsYOcw7uCwC0jdhTeGgTtX1XBslbVBVIziySzlE4K7ZuL1Tgr7d31M3wvJXv0gwO7J
jBvKcJuEg3C5E/68Fxm+UANschsRSD9n7jaT4HO2MPmQi2r+3NUHdwagHGZWs2ma/9z6yskkgmRu
o3UZwTGbnwVT3QATXo3t2Dg0V2iNdNvWOauIcueBtg+pKL1FzBmm9gs5+5PhLFqAMup/O8RVVVp2
VtIOc6C/2IgO7uvb8EtV2/WsOz8cIA9ekBJJgsX4h1FMnh7QsqBqHKLe1cTz285HEak669tpg7No
a0+TpP6Yy7MvpDF6O7BF6JrL0wXlGk2gSvhhYDJTPQ19Im8cAg91hUN8wRVnCYgFhXQgl6qOqqZj
s6eTIrczSVoyJUPtV5i4/0QJTvC318+WyEFx1828SocgWiKE2+PJc6VdzCvOsqRKieBjFGeK1JUx
uSVXT6ZHFS2YhXjeqF3D7FoWKXbH953T1dYMhPXupQdtBGZ7aRsRQhf9rAcQ4+3PJtNdx5/XWz2z
eRPCz9xXh+rjfhFRcDY9P0GOgr+ej5GT+anBKD/EWrBQec9tPgaAPIbBg388wnljv5UGzQiA+JOs
rM2BFHp/vnSJ5P0ZdVd/BG2XQqi0gWz3FnR44hTGTUbiI4TthoeODt5cyUgdD1VgIMrl0X3bU/5p
ob1PpCC0CFmoRXPDEGwMBEhzu2egd/boanSK14n/2W81qeF5uxkbNi9a2ymz9trLGbfBvleR2DXA
9EwINhNsn3modZKmdHbvbxgW3M1OASpWMmIr+zloyBBf6VdpUpkSCSBDB1SfuLNkk0T3Y2yWxxIy
KVD4NBEhSBZPYMOKFHQhUlyElMG6cMuYIV7wOPkVi5LwBLm0NF1EfT3X2/SGFPfkVwY3RF6Rhfyc
9rfIz0mDLLzTteQpkesIB13jvhbN0WEhlHrItUzCi8EwWkWKOnMjMQocftTN652eUHsUV3gMTv7O
1H7iq/McSCPe51LxHG3aV4+W6kLVLJWwsGdgB8bnW0q76aq9PCDIo6tu7iLmJ3/G+V3NdKTm6BLu
qQKowwe5E3xcGlfVj3xxJ7cAgBPGCSqbH6L/v8s4rlwWI9AvnqWjCRu57ilRYCeNcDKspjQYTVbl
CilWLyNb/L4FF0EVL7HqP+wZqbVn44Jt8Ul8wYqiOuoS5AlvOhJ4DumKtSP1ZCg5JJuSdgVEEfle
rueRNlZX55WW9wJAXR1ILO+IfvG9fj9oC1WcFddJEtwZ8rOQ7QIMf5UbWQ3uYhCnIpmFI+tvsU2J
aQKyDtIyhrfqmXPRaLAaX93rduOKtfUyoSwE34aelYt9YT2gdr4Dtl5H3gLKWJF47OIvVofi7H9V
v4KisCAldOfaaMNOd5swJlSqwHBrVTMRcPXKQGKefNDWFAH9gjO8M0vNpKAoIn7Qj4vR9HvdEIjl
xOxXdiP0zxUVhb97GJ985I9d4Xx1HUCw7nF0CiyxhHDdhVXsF5qAakhgFfoIqmeDSa67GL6ogbp5
573r7CQXdTPNC/p3yT69lFt11lbQkRNFggJf2ukMmRkt/xlONDfi4yXyMDdasgzqw11ufKS2gnDI
q2yQCZrxTQzVr4/Rv/8IvIguAwLlKAuiJxb1wb29TDgIXnoUHNjO17Z1xtkg3cMJ2n5cWnscrwvX
Ov51FWnVaIzFNSSkmvGQzafD0VEBKDknm62BXr08NhAmQRaVzRVGg0XA71huH5aajFgwpDBXgmyq
f0UKjv10H9OmfufQztUcdvVMlcKtflDyIeL5THKpeqVN8P5WtPKj2L2oYM9ovX1kBMtp51m5ZCIH
qpZAYwuh2QQxTxjR2XeMuZiOSXP2+9U4xH8MGu01lcwOX4SOIBDfXRB5akkUMY+okiUK1G11SipA
Fka3DajcM84sVWLz91QqHL6AtkwRZpFiOJPY1qFsrHiDb5sRDZVAGRfiWvDCUMzdID/CJQxoyupr
Rvw5GKe6k6UAl9bXOc+c/wJgY/HP8AHGkiGM2xdJ4+DclOxoz0TPIlQmiZ+t9bJac9aMYVsa4FJ6
ZFW2cmTle6pfdA5UKWNE/iVSmAPfKasf4QtJedoDrvEjjyHGB6fB36mg9jN0PTScVCxpiZIs1heB
1CJe3RqHWCpQQPuUeSEdEeEtHm3zzdWNRmeQnaaG1XA+LH7vSGDqfY+gDNBXy65IRGoDEcuuuHSB
MAITzgXZVD/ktY7hvdLS/6gfBuzj776AZJygJgMKYZMzprCCNEdTbPNjxKIM1MlXUgLhw9V9hrfP
NyN8QlZpXz40B5XBF485X1vZmAx91tqAcCLQqm71oi9ojhGC9a0OuSWLi7PsgRsglhfV0r+R2231
732k+aGGIiB2oJ7zRSXuxPYlWaSYbc5fWTdNWBkmRC8jX7YnwxIyQE5oXWlYok7xVZKzFPYlsV5U
LTQ+r+JL56kGMs6XR1N3852iro/yLnWSCR8T1G0HwSxHtX7rmtk32Nn6AW1Gwo2zKQCFWQ==
`protect end_protected
