��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒������O� KFe�gAn'�i�v���k@D�	�q����%����#�����z>�zl�"��:���B�'�fC$0�����D�`��qTܜɎ�X#v�t`��B�y��.wr��<G�|�L��nQ �&�wG#7�h���[��]Q�ó�Z�m�䚡�)�z��0��� N"�`t ���YL��4���4x�Fä�c�Y���t�T�~ ����;�(�;tL�3��~K/F|���G�.6t,��<%F�c�6�`Y����+P�T��f��~B�[��IO�~��ʐR+/8�H��-�s�,�Z��"#rY�6^t����k�*zU��5s�ؿ�����{�����R}MdQ%�F<�� �N��h�jʝ�k@w�'ځ]e� ����̥V�C	���1���GVQg>�lK�.o{e���	���
���Yz���S��<���$z��^[�IMF(/����WI�aX��.x@�ؖ�"λ�^�������ZVt�vD��)���2ke�r�:p�SG������@6k���G������q��@Oi.���i��\�;������^MO:�
��+1e�"�֠^C��ù��+׻��JE��7�6z��ͩ��t&z��y�� Q��7�(��7Wh�R(�7z�cpF�� @O�n	P���?d�͂�
��I�ޤ�*�
��2>3�3ɴ���&&`w�u�OԪ�CF��`��E�@M���	���s�jw�HH;�l,�*����yE �/�o6�Fho�[�P�6�z�s���8��%)�"�� C�p<j#���3��S$���n��ʪ��@��E#� �,z��=���!sI��S�Z���r
�2�;z���c��1�.��5�|�������X��R��]��{Q2�c�qK���K�-]2�V��h�!xf�o��!�h��u��$�EZ���X�읭AX��g�A��;4��Z�o��"��Q9^0�8Seӂ����Mc���,�KB��Aԇw�t7+W���(;?U���2�[��P`9R'^˄|�4�s֞��h}��X��Y��+.��N�k\o~'OwG\�&�'{�3D���U�ԃ����d1�Z"�Q�)P�-?v��G'b_�S�x������5xN	m5PXT�� �"������3
}E���8�aM���n�3���PU�|�!!�1b9��#�ah�)ǡC��_���=�* ��+��ٌ�l��[������*�R�
k�����	�_�~F�(�ҿ����E�jo�+<�k�f�p`C��U7t|^ǈ��DJ��`�	KIXB�eG$�M�Ǚrw���ğ�a�H7;�)��j'��;�jJ"h]�I�����I����c�C���`���s���	���,GiG��TE����%��^��)wsZq(�3;BE+0��I*K�LEƛX^�:K1դ�'�-~�Rm�ޑ�M ���a.����/��kV��%�8ަ�=�{��$_�H� c(\I.] �TE����t�3���9��k��^x1z�1��'xS[HJ^�z=��*��g�7��%��������4}�l\�?���W��X>� �E|һ��$��>hs';^㠚xF�/+�k>J�b�%Zf2��r�#`�}p1ǭG�W��0�Q3��E�����8��5PHv�¼Y޿��i*���ᙷ������0�����3\�8��ތ~ \aޕ;%�cs�a��6����G��V�,�|m	|��?T���֖�OP�I��EG�ڟ3�T=w��]�볈�שd�쎸�:��>������q�o�iq�Q����� Y��g%�N]���AĒ�q�%�+�Q��*ϵՂE�����H֋�(\w��Ђe��K��&�HUc�y ���w�߾�
��[&K��4],��L@���Q�9�z|���P���vje��q��	�g�aYi�_����-2#Y]��F�\���(�~�����h�e"/᳡�S�)�,�!�:�F�2�}��*�)�U���eޮ�p�C�u�� S���һ�y�0�~��W�c���U�^�fɥ<&.�@��+DN�t���ӯ�9�Tqr�%mV�	�M���-��q��Ɣ�`��)R{rܑ��~">�#ax&��2?�u��j����1���} ����i랳\;� �da��C���fvL׶���2�牙W�;�[2���W�d>{���>�̈�\·YI�vC&
0����/(��1yaly	�%1�D*�x�8�&���mJI�~�,`��V��:h>i�,ͺ~��ݝ,�b�W"7Ko<,)�Se#q�����-��L(�^&��晁C xy�e�rRD��0�n4e��M����ѫK�F��������{��MV�^�l�S�X�D�1Mj���A*R3�,]/&~v��>�������L}3��(�H�h���C"�� Y���fluD�k��(����r@��"�S���=�T�kR�TmJ��a�Ӱ.��v�sh���da�[2\�G�:d�g��p��l���*+�c�fԲ��Ӆ��R$�ŴZ��U���ǈH������*5�v;��Ϻm��qC��`�'�&�FK� k�M�ԅJ�� B8��Y�������[�������>����n���0H�O��6WVB�/ɣ �9r2����>+ŉ�? ����V����2�Dg���&cB���*�"��-q��ڦ&e�2�kBb���8_�X��
/��7������"R���е����߷���m���Z!j�5]�m+Y���X�́pf>	�Y;AZ�!&j6U����`,��<DQ�E�t}��"�Y��l_m�Q�|�A�	+�A�M�}��5�\��Eֹ���yjķ���ci������<�Y�`z�����-o"����|��!�]8%sG�ӏ�x?9�o��Y�2�3|�tnnu��ʕ�YI�v�9�1�C��̲�U�c�+��h�vm��zGVLc��6�c��؞�i�o�\Vv��)Z�s�������g̨x{g��#�Uf$F�=��dm|V�ׇ@|�&m.[L��k��F�Ԍ����<�O�[i*�/��a��_�t�ٌ-EVzI{���Jc³_0�L�[�� ���4��G�S|C�BI��1��l!g%���pQT+�geWF�i�/~�l�����
���VN]	�*�:!��O���R����G�Q|-N2�����k�.ow��?I�Td�R/���H����8�H�︚�k����9eH[ m0&�C^j�(���<�u��j��Y��8Ƕ�L[_��}�:�����7;�7%�V����r���qj�� 6�|`������;��""'�wy�4T	�t�^�!�5��@�R8g��.�R�ȫA&$����G�����M:����[�0M�ި���S��I0鶭tZ?�����s�׆�^?��a@]��s0�Ꝅ�u�s�1y��r'CV��B�S'5�>d�,��R����$[�0�#�A��S+A���˨��m���fIx9$�w���hFtc��ݞ��[�ɀ�c�ޡJ㾝 ����0NS�.{]��U��B)�tKbBS�q��t��K��k���,=�z�Z�+"i�E�'p�`49�*.��鉠�)�i��C� ��л|�j��|�������K�9�
'��Ѯ��t5���y\�Iǰ�]��l-�9Q=X+T�Q�lîpj�Y�E��ZPA����,���:��f���{�9�!�-�,m	�Bc��L���YbiH���<dڒ�k�g[��� ���!��)7��Lr�(�*��1w�
炙�v��b��hծEw<b�E\�]�nnf��GuCZ�u;-(5���r|ϒ�Ρ�6��a
B<u�AKᒟO֞�m��Q��F �cf+M�J
��k�@%qđ"+6wr��'�#��8O��U�zk�Ι��Z2�zLm�V��/�����h]��,�g��/�6�aA�.�o�6�.�gW<C<���k������C0�&?D���k���^A���`�7$/�'*<�Ax<��}�N�5jr�O!l��/���Z�W�sQ���ma�4�b���n�l���YI7�l��3�ix��RՂ�g�/�&��ܣ�19[�Kqg��ow��p����"�8?�07H',�r���扫`K#y�[=��̲����&�T�"��UMc�Y�[)ћ�l��3(QҖmj����&�L'��_%]����;2~��������o�;��-�4~E�{Ap��3;��+��Z�{ƘL)t�q�D&���F��p�o��&/;�<��ւ��ljV�e-$p�=���E׵-���yJ> ���M�m�2���� T��jK�IkQ��3,|h�ǀ�ؑ���H���o��ɫR�����o��~��6w�_X���� ��:o%9�E8����W��NjG�̺�<A3�ѽ3�����-�l�VUfex���O �C�����|)S�Ph�"��6� ''�t��hF�(Q6�����������S����]��!W*���[p��_�لS�����0%1��}�A�}͵E=����f���Uf�i����AB�"�U�.�Y61��r�?w����De�4X��o���x��T�s��l�82Jm6�l�p�{��-�#��Ye,m��f8ܒF��(��P��	��
"�C���S��';Oi�p�e�P:W`(�46���_3�c/��~�=��.��Sk�z��Vj�����&*:�g�F�
@�jCL%E����z �~�ˌw���)%_xL���[���nQ]Qn�C��~.�"v@�T�S�Q��	�EM0�,�,;����h������cҐ�����ҴW;�Nm=U#��@�'�*��aHÌNŤf��=��S�V5�>:-HB_?Y��%�=��o��&��.��U����k��1�?�uC�NY7��<��.e`>��Q;|�5��Hdwn�Y�6����S�����c�dd��ܗ	�����ӄ�s�%C�ۘ�K7g��ɝN�B�&(^`�9(Y�J��6��A�ml|� �-��B�$�tCR����[@�PF)�藫��!�P���מ1���ѵ����`��0̗�e,u�3Z���뽫�mӂ`퉐��Dc(��OOd_�7�'��n���z��r��ȧ@�ֹL��dG�m�1{6�_��%���Hb6���ń��� �ns�*G\1܂9��7z�>E!2:�,��-�X*c�C҉��1]�.���_;3�]�! X.Y����K��vG	��X����y�2 ���'+�����cIX�ޠ��Y饏�6�Iɒ�x�)[��7F߳��jL"�sQY��H��-�L{e�u��sC��;��H9��G͏U�:R޵z(�Z#�Z=�n8xa��V�QwSFt	�j��y�y��mL
t=���������4��H:P��핷��1��?�h^{�^/��2�%*ܺ}��U�
ʑ�gfn�8�Q˦'�����x�b`�3�E6CQ��� ���br�W.U ��>��U�hԚY���M�k$�A'a��s��sq��``b�[r���������	Zf2����L����*_�<�f��g�R�u����6���/��Y�m��B���<O���DS���Ѕm�o ����k���*���uz�<^W�$�}�#`1N�� ��?����	�d�{2�w�7� ��W�w�e���B?>k�9wD/��/��9�Y,b|�Sq*����!!��Hl���:���T;a�{j�+�0�nI�R��.
|n?�Z�VR���ZS�����]�a��}d�bNՑ�v���Z������ֲ��y�� �����/~��1����./�/��A�;�j��v�Z���%����㵼L��Z����ӑ��K�E���-�|�t-f����ވ�s!t������SD0��,LeV��Q,QX�5xD��*heS�D��bQ[l��g��Gm[��l�mo�QN$�%���!�8ȡ� �W���A�����`��FU3��F���bqf;IPO�ٝ���$�8 �;��0L�U��Og���S�@IN�(���$=\�q��#�B:���P��&�U1i�a����ic��i��΅�U���X�"�L��b`*r&1�+Vd� ��BV@q0D��^?��kQ
�`U���K%�3b6��Q�(��2��%Ӱ��
E��:�ɿ�X��2G�>k<snmON:����J��~���K(~�r��ƺY�~Yn��^6���cr�a�Kʴ�U �l7SS�����`C4��]�_^;�mВ�ܱ��GD�~�2J �B]*�|��AV/
�����T�"�ˤ�xgޒaT���iXZ�%��QtԘ��Ut+�S�S5{�Ͱ"&m{n�e��N0��|/�(��Vd��l1K���G2,:���e���歠�&���0����N��7�B��u�JQ��&�R��@��~g��9�os#��kf�p��k����o��L�ڑ��v�[
��s�q�S�r�}ϩ�G��O�����Mc�u���t���B��k�H΢���a�K�]!?�������x� ��Zִ�^^NVN_ڀ�m�&~i�z'DhXō���
Qu�￢���f6o��%ŀ/�_�o2wbZ����nҺ͚\�%?�"����q���6>�p��jm�o���=��Q&�g�q�q��I�a�#���r޹��ӻ��A���b�u��ǳ�cd����>Y�<!��j��mj��+7SdPT��	5�c�j$����0펊��+�|#u������B<܊oĉ�X@���ѣ�v�����nj�扳��&��XޭsbN�}s6��,P�$	�*��{��?��.ƨN�Z�xvx�}���Wd�����QlK� e�f�!GGړ�ݾ	��>�-��g��Q�j`m�>v9�)}�CO��x���6'Xw�ߨىF���v�����U�c�����s�����v��(�� �)X��ƪ��`
q�P��[d.�QtŔ\ ���J2��Q=��y%v4�ƛ|b	G����T�	��.�����׆�W����0�-���KYA.K��Y4���ӑb*�u�D<����5��A�xi͡�	9�a�z?��_�2�F^l������%^�W�Ў�rX���
dy�UOq4�v?�H�:f�q�"k�y:��!���� w��}��0<�N#�����r���oO O��}�&xOBI~~W\������0���<}i�?$@�E���F�Yv�%��x+������L��J�@�g��]A;tA9������e�{�tz@Eg�7���R�r�ǧ�?� )Q�҅*F���@��rZ�B�wNQS�;�݇�o��#AQu�vv���K <�!�{�@r���C���	|Ŕ:K�� �J������J���*�k��$	���I{���'�������P��(c�9:"��P]sz�]���-_��mB����^#GxG�y�sG#ƒ&�~�?�84ke�r�ͩ?�P[��/���,{-��V�Z��cJ�G����� �m.�uኊ5G޴e�ɸ��ʶ�d���E�z�k��?�p(�\�>LP�52�Ѡ1{���b����pN_�S���S�t|��N����b�Bl�h�vw��D8�-�N;��S���'F�C���.F����D�4����b�g}�bP,`&M��6t�S��ٿ�%�{�F�B\��[E���a���v���gey�"�l�j�1^�3	���ϫ�v<7L 6�{�-�٫�Q(����е�8���'lś��/_S��8��#eF�����0����3j8-R�l���Ŋ�|� b#��H|Ƹv�&�y�6���]�x��F�X#�:D�I��i�{���8�R��Rxj3ौ���ȃ��R°`A7|�HЙi�D]��r��&��Z}i������IZ�׋v�qҐNVB��gl������G!��xZ�|1QK&j��̗,�IҦb$zdxp����gأ�G�+>��"��sX���~ҌR"��M�K���>"�e�0İ'a�=i�l�`8#x�١�*k���h���8^NΨ�pDwD�O����k��I5@����*����BQ�S�E�:9��ʻп���;'�X"v��������Պ���e"��������%dC�i	ׅ����m�q��o�bˁP�'�V�AR��F|z�B�~#\�x"���ܜ�n�4c�Su3:R�r#�).�,V��~C%HE��W<%�ҝ�ɗ�^k��X��Oyfk|J�B������	�+��J?��+Ȱs�$J����'���uP@32Ү��H&ط��f�|W_	 ���ڠp�A�Y�r�A������a�\��.�������Bwֺ\w$�"k�Q�&3+�N���Jҽ��4[zU��(��ѥʘ����i�0���;��&n2����YO�_$^�^�� +�8}��qp�1ƟwWP{���c���W�.��^���� ;)��4���a.���PC�[Ɵ*m����� ۫���;	���9��Uzb7�5Kb���h?=��:zl�l�4��d�g�eRj�J7��$�"��g��u�P -,����\�:�L`�����&��zFȄ����b�X��y�^:�r��8��D�����mJ�Ey����ں/��+����_�r���{;�jm�:&�}�Kd O�f�V���Z!d��>�����	P���Mɰ3F
���W�Oi�\�Vz�O�6:�Ba�r������oT&�\�M�����/�u:D6Ĥc%f�o�y�qҷ0���A;�"�����륺#�|�ҩ�'eUq�[��il#hr�����ܧ������0��.`��şf|7�)��������|��B�<�ORh;��Ek����z\-	?D��+`���Q�q�����F�q��������{�P�e�N�-�`��X�s���B݉�8egn��>\����x���_$Ի�9�q=t$�����yt��]F�b���⊠��P�ۿ���O���n��R���]��I8��C�d�0{�CFN������G���� tͥm���&aR/Q~�j[[�R$+��ǎ%�������v���Dɋn�E���T�Rw�}a"��h}c[�hu�h����88��/��N����O���N�,��hE�G�C6Z��븟�1��'��jt��~����t�3����מ{���VL�u�Y��_�T�d��X�$5.�����u�A��u��I�b�8����Q8����U��n�:�3R��(9?4�����Q��~dC-��0��ƩT��$�vܵ�r��=?y|��'�f��\����9���\#*��l�����5��od�$ӝ_�bʬ�{�rҢ��t�B/�@'��AR�ī��`+�ᗠ�9�|~m2���||��g6�F�݋]L1E�Q�x�g���F���H�a���IjD�\3�u -e�?۴-�¢�\|Ëj֕�a���A�8%�U�����|:e�#��O���?$�Պ�U���E)�����*~HLW����L�r_�c��1�5�7������m8�d����Z��ݤ��$�I����AVzֵ���Kz��w*��^.~(��/x�����g��u� 4ա[0�o�V�7�Ⱦڐ��?�����!�����O
���w�1bA��:4q�RPnY�)pD*Pڕ���0�?��EmC7�I<9���p�#�W

> �ҫ��9�a���~���P�p�X�>%�3J
�H��� +�[�6 g�"9#�F�M�����bnٶf���ƚ����"�D_�R�$�o��-k;�ƞM��<��0�<u>�.���S�oL=̊qo�i����ߏR�դ�0����ޠ~����-#HBz� _7{�pa|}�fm�[��<K�7/8�+�擳���
���%� -�k��M�uuՕ[�7rn��K�K��3
_�ir�=P|����`����v}��%HǬ�B|���U�f�?(&���K,Ō81�)5���� ����SV�w� X�a�A�Cq��wzK�7�%c��5����W�����$cj���Dzl�q_K(0�9w�/j�����I�`�#�j���	��(1�B4W���g�y��op+kʮL��H��* �6dɟnb�]}g}��H+c)c�t%��4�k�o�!�ljޕ��Y�w�eh(�����S��v���%l\�8�q䶨z����gE[N�:cϮ|W2S5|*�L��؇p�iӂ���9�j ��
�6�KH�?���A�i ��#��__
ȣ�JT#�zF_�(C��/���I��0aP�(Ob�P�j@�{6�1a H��L�q�$j���
7ء��L�3�l����#��p[ժ�%1��L�ʴ�W�c���+:�&��|r/�2K������9�w�}N���W�"6�h2"�t�*>PM���KMM&`�,���'�ވ��������k���Db����^[K�'�΁� 3��r��Cf�j�&�DVw���?A�[���(�㎸۝�P���9�;8��a��1�(k�IP�u-F6�<�d��pz����Agk��������k-Bn%�p��l9+�=��!�_ț��ӑ�{�w�(�F6�3��Ѽ��)�eO��!��ɈW��r�{qL�WO���f
Ùb���Wq)��(|}���[�h�9�zAt� �ޛ�=����&[��ݯ�e���'3�_�\QxF�悊U, �=���VIƾ��(�=<�
�*2�bC �a�6���-�WK�/����K&9���3}�#�������$˰���ޓ01�H)#���`5�h��"�n��r�l�Yɯr��R�99�÷y*̪N����i��|�35֑�.��&�#�~Q����S��x	SD'H��3�a�q�c:��Xɷ8bCo�6���ݏ�6�>;��$~�=�'�.)���d��8����w"����Lg�M�\�(H�P5� Q ȯS-W��>�w�&*a���A|[�o��k���2P�,q���|o���d;��b��q�I�.���B�ȹ��wp#)�@mm|<
��~G`��G9vF��1&���c���ԯ��:���<Ě���Y�8eqmFh��>��j۷��܀zO��4J�x"���E�99� �-�d���45o�I� t@y��9�Q.��,@�$q���-�-���uY���X/>�_�%v-��3�=�'Y�c'��~�W �u�����|)��Tr�K�n}��฽������Rz<��	=��긃���7 h�Z~M��/>iuй�ܟ�='���q�3\7[�����!���V0jZ��"�y�)&��,4��(�2�\g	AV��8��x��10���x�1�����`�n��N|��
���Y��Z���VWeQ���Xw@i��	�^ٖMvŰ��U��"�H��O`���\R�kO��~"y�s��D� v�6�D�MIys�p�ϧ�8崾����;��k�_��A�0`u�r�ĽE���E�@MY�-M��Z�t.��K�ߚL��ϭ|iQI������p��v�&��Vm:.d��*Z{D�p)��s64/B�<�+�N����hnϴ\��i8��#�����`:�.2j?6�̢=0\�ox�����yC�xl��2R3��f�ĭ}+�I����gfY��VQV�6AI_��:�jd��F�LU���x�Q�>3�&@O*¢�����v���`��Y�_|h��o*���"��[�E_�&1RI�pYR�M̿EHR����딍�V��m�t������l�xm��\](�Q��X�x���u�ݨ�uT�x��[�/H���\�%`�k��}��hT�6ʯ��*�[�\9�:�4`�^v�`0ӭ��>��������]�]EU���	�1��Z[�ꓥ�� ��p59��fw	+���&��iܭX�b�L��ݧ��k���+۲ɃJI���w3ȦqH��[	�w�����iKWr�ɤ�ˑ��d��D8�~��pCo�P$
��#�9�	�fH��
c��~�ҹ0��:��Q�]�1rb�V���k;Y�y2��hF+��%�d�^����Bq�A*��gGO���2�N��p�GҒi�8z����4C��o��7�`�m��3�^��=/c�����ԧ���Z7��x�����������cm��X�s���G ��0�K�'���9��A\���|S�)�8V{�AB�/������T�ݍ�C ǎ9'b�a�7��zj�s���.}iJ	�_Z$��B[�[i�?�~`�����_�[��[�D/PE�t�f�D);�a���Be��i��|2ر�S���|i	��:�Z�����[��9�آ���$�Z�t�G��g6[���S�$xj���7Ӗ�h]�b�XQ��,B!�����	!	8 r�M�!��@��I5'K���|�Cʩ�,�n�̗�:���5�.��l�X)?����9s�p�,�����I�b�:�����ҟd;��lt�f��]~T�H�d�qi�w��t��UN�O|w�y9�J66uSy>B��?���*]RKg���b����H��C����Y�z5Bׁ���F{��'ྋ�N+=��6f�e��	�|R�:��،W��_��5�L�<��e��|,���Z��d����t18:�ǧ�y��A�'��h��*�M���d"�}�˖�y&Z8�ڀ7����*TIN�TJ�}�7�����O�\s�t��*�5�sl{X��u���hD4��R�'2���^0F�<�H��v6�_x��b���� wA�Ek�!F��Ed���. 1�ۑ�l]J]��j�.S��l���w��̗z�o�z�E����1��7���x*�`��M��U�y5����L��ծ���F��q����}k�s�+��jB0>�̡\®�lx�&P���J��!=��v�ҝ��|�-�(�m�7���L[4��#�^(�kR�ǃo�i�إ�3�n�B�����B��Р��F,�Z2��ݩB��R�z.T�=4 ��]��ͮGձ����ᙝ�ms�������N��%P�c��t��L���/}�x>�����]���|d���r����Q����7ڔ$"n��ƣf\��]Kվl�!�4
���3sl|�Yh��_���	~լ.E��-�+ޔe�S6�������w�:��ZzGZr��K���鐼��tᚲ;vP/��X\V�����5�{���Ȅ�Isj\ă��~�s��~�kfqͼ�L�*Xa��iy�A�w����XjE0\:f�J�!#b;pN"}nI��]�DXg��$d��K��E	�os�-������F�M��6q��%gqB��=m��{gw57�+�Ҿ}�T�_�9"�h&4���ۖ���y�/d�E�7j�X2s6�=�� u��	����w� `~���3GS�f�kj��:��U_����@�p��bz!�b��/dsB�-����8����|��}��� ���,/�a]X�E�Q�W*��^?пyG�c�����d��H�]-1Q�F5���� t0�i�����i;��$����39��#��.����A�+䟉I�? �b>�o��!�	k������h���4[�#� :�����m�}�N ��Iym�����t��9�<��u��s������2'�����8�>�J��͗_<�d���U8I<�w��z�� ���K�����''p�����zܾ.������������|��y��py�ӝ�����sN�!�	pҔ��;�vɂe`)�+�
v�Wa+�/����ʹ8�L£)����0����K��3�]I^�d&�Fb�o(@p�����V�� �<t5��r��Mv��$��A��PG����6q3S��W��Z�Wq���k5���r2��0��=�o��qu�����<i��[)�
�똫&���R�f/��G���WX�b��y�t��$��ސ�P�(��d;@�y)�����nH3����R�t8� ��,���*�7C���d?D��Q;��X�5�!��z����d��9�V�MH�n�6.'���o����Hn��m���_�vy��)�㤣�IIRo�����!�y�r�*����֦Mg�����w?��;��u+Dl�9�V�;#�X���(ӟ�AU����2�H�_���zßu�ʀi���-�&nan���9�K)�ý@� ����Ȑ=�J�)ө���-z��~�1��2���%Vq�}�R��-��J�N�*�0GA���\I���MR��)��o�U�nu�]��l�����R��������q9�cE Z@��ȷT})��`	8�3,P����g��Z�j�`W}�^Dԉ@#��6u`�ʲt	��>�T�_��n�ȯ��u9>�>�W��ɀKEQVֶ��73��?�2��_XE�4��C�c`"��S�ƅ�������Uo�P��L+�U]�����I���.��ܟv9g���QJ���O��x�2����7�G�+5}'��+ʹ4�J
���X�>�� �n�=�h���kDsK^��ǂra���ƕ�,|+�˩�![�-u�r�-2�m��T):�g�HHXR6X�g+K�V=%ۋt���8�N-z"�8�'Gz�F|G:3%,,����D�k%�A_�P�?"�~t�EG����p[�G)���x3�S�(�XC]饣�u���S���3�V���)�>\P߂Y��
I�e��7by�����F���� �D����$ 5����Zؐ��g������R�!	k]*���I2�"���ҥ%��3�Z�������oO��q��`�]�<r=��4�(�7�>��`�	?qq�ׂ�=�������c��}Ҟ�㪥F���<��3��h#�7C��b ������1�T�Uv��;Ѣ'|2��hӤGN�i���/�7�{��Cd(G��{|�
�E���0����>��d$b)ᖚS�Q�l�X��ZG��҄^݃�SMH�����%�ʖ\��yŒ���kN5����-�KXbX��J*Aq����/F�pao��5U-�2T�jҊ[��?ޠ�Xj�犠�JsSY�L��5�gK��J\k��;4dd���fzg��P�������l����A�;�ǲ���� Q =ϻ	��f7�������F�M<ie��v-']�L�=��"��4���%3�����*�S-�7�"@���X$x`P����%N�jɤ�XۑP�g��J�>NhDd��TF�'��C�T���(��-B�p�:�wǀ�'��IZ���	
DT�|��*Z������ꝖO�&�>5[�G�h�vl���G����m��&��Qw�lI��%�����m�,D�*&���;�$�Jb[�*�Û��L6����{2	6B��UHĵ�R��'!�W!�u���ZG�-u,�W�|<%'ys/E�2��Pul�G������V'����q�dn�~��^y�/o��Ō3Sb����6S�h�����W�sS��997��u�`J����ΠH����)\�~��V�_AF�����s�ȵ	���n;d�P��6ƽ��<��Rk�_��?�*B,�V�bD����-�(�	�:��iC{P1�!�!m�L�>�(͜�y�p<���c��S9_H����{(���&�ޑ�o���{Ƹ��Oy(� �`ֽ�
���ns�F�#�ne��$�kPs�;a���L.�p���}u�a�P��W7ד�޻��з�O7���Co\��W����̀��!sPG�ؾK��N��?c�V���-��C�C"�*d�x_yЖC��5?���F��fG�	������R��&�m�����o,�v˙d3����D�AҤ�N#o.7��Q�{�C�݋O�!�%F�:0K 6���V�@��"����ټԊ��YM�Z_�T�ra��VA��7W�x�d�bO�<3 ĒƐK�0�\*�6 FӍ�mZp�U��B�B��{2�1@6}L]}�P��������d�l���@Q���]�̑�0�����_���dz�6I����4j�cn$ ��O�c����t&�9T}�r���Ĺ���I'���P1i]:q�^�-PJ��a������ߎ�
 ��QLr,㸒�M���n� ��+� �S��0b�fK��P��Yӂ��6�W����jE�!5����]D�ř��o6c.�}�UM�o#�q�<���2��y`���9�
W��m��Uz}��"�vc��s��tA*�B�z�Ai��㸌��;��e�D`��n��	�|"�"ј<؂t���X���%$�t��Wo�c�4F�0�ݮ��@���5���b6�SY��w�3	{��?��v�$�E{�#p��Y�A1�<>1Qr ���,��pD�(8L�:L��!���1S"���7|�Kܧ��$)�������C�1u�>��v��^L�Y������=D����O}��뫞GL���m�p$"�v;�Q4�W:�Zu_� �k��q5�J��A;�5s9۳RF�.���.D��m��'c,zs:�Y�vL�����w�qJx�����$th<�ş{D`z��������D�chs{�vf7�Ѫ$��[�UV�	Ю��;4�@�"9�:��C�Y���j�D�y�=�� �mB6eU�%�d`��Vi0���C�ʈf�f�1�LAϧG����k�(%�R�z��/�zͮ�\���`[�Y��|Kw�@�Z�%*���6�L`R�Q!�����/��(M����@����?���t���9�i�~�(R��x����{ڋz�t��ª�{p=����w`ǧ&���He� {�UK4�HNX�D�]cڵ��[���ޔ�y�M�#l�%s���ac~����b�U�3s} ��f=i��1F�ss���	m �/�N��.L��y@5�F������$W(HŊ����#i�?��i�c���b��{��)�P����҄.�����h@9��J��v	��e�'�����6\��8��N�Ec�	S+�5#ժL(>����x����~Y�"��/�Ҩ/Ф�����+�(m����+�-�B|�4�_7�q{�� �>�Ē���1�z�L��+�a��[�+X���aO-������%΄�'�s4�u���w���	���0�
�VeV��|�s��wʙ|�Ӥ���ө��iX��ƞSTJ��;Qɿ� .s@�3����ŤT-+!�s>^)	x�?���\��W�!���g�/�
*��������]�4�c>9�C�9aX�Z�Z�e�tǭ:��,��0-H�H�%Bk�!�ۻ�o�uMVD���b��ވfc4#�g���~�"���
�N���~Q����EoU:׋�Lnԏ��ˣ D9�R�I5��&�;�J����Ii��݂�g�u,�����Fk>r� m��[`%��K��m�/�i1K��|�5�h#I��v���տB����9�Ӄ얱�hf;�T�T����@`�r,d��x�o�Z���;L��n��T�(�vz��Aw5� StzH��آ�Ս��z�*u�B��x4�6��%2�%/!>9l�A���h�r�_<�D~|'�/Oz�_�\,�#GǙ��t8����І!`�DS���(�!�Y��*�w�������cˀ�8{iU�W�D��M"��m�'ۆ]��p`��0��!i.�Fr�����x�]�ݡ���A$����:���/}��2u�s����*,[NW},�H��4co?`+���-���^T[��|�1y�!:���5�89��N��Ì��>��~P�|�^����=n��`�&2�G��H[�����R���7J'n.v�ʦ+�����d���`����(	X�0���>�m��ٌI�֡�C@ϊT���؞ o#��N��,�fh�r�N����ih�XDl��+�x' ��� iy\�!�o�h�iQǅk˦<��^���&� j�&1Ié�6�h�_�OM����_4Z��������d��:+Sa�%I�%$�\�[��ykC����f�>�N[���t�J\岷�rp�v?9QZi�A�k���$�p��G�8����r�����+��9N�[��`x��Iq��<��gkf�3.s���9G�Ӂ�&�����@P�]C�*�Xk������n�E�1l?��k��(��[��n��q5䞝���(��B����}���\����te>�b#�Eu�D�,�-Q,�ƶ�X�(2^ؤ8�k#�ٔ MQ�7'�J{
�B�1oA�u8NW�ln���ry�#�7�����y��6(�t�3��yi�*�:�L�ݥ+�dY~�B��6�G�q��� i�_���E%��^
��r D؆���ګtK�5Vfhn
#=�W�����"㶸��ʘ�7^A�"*!
d�dv�r������<�079elFUN ��	��l��J������#.�ܵUi��ɣ�n��O�xi�v�
"An��r��������)A���K�
NDB��$��?�����4J�?.�o~F
%��K��nj��>z�����YK�3S�A9�&������´�g�58պI�=�9I�ؚoh8�)�>��6������c���^^��Er�^�yDK����ů�����3We���lD[�ko����#��� �s��`��Ȳ>V�ezrS����V4��H��#Zrկ����5�	�����?9��pw<d��OR��s�)A���=Qa�t΀nX�P\���n��Q{K����Sibp�r�B�ع�WmG������~�BH�	��j����|N@��Uظ]¤-?%���Ḥ6Ȃ����R�'��:R�۔���#$i�6�V��,�W�(�0��\� #[MA��V
0)͇�����4��a��&z�6�&�.v�u���ކ��y%E����ר��ϳ�#d%^x�k�M�v�:���!��8�S��5�
�q�����x=WA��|E?��(>Įj��B���vZX��}��pDe������ɻ�]�+�<�Uzm誖�q�' �6��F��݆�¶�Q�+5jp
���8���#J�1�O
�'^w��g������X)ׅQ�~�4xޛ6+�Y.t�W�q�A���\��Wu�m#�J���*j�*fk�QՊd��x�RX�W4�Er7^n�f�;`W�>4�W�7����ZW��M�ɽ�~<��6��z�����LߟCޙn6b#��?»��>��-���Jeɺ1�EKw^���neb�i��\ɽnK�4Fͧ�rqt7�=�$ӥ�u����7$a�%8��τr(p��\]3}N��>+���2��ٶ�K7�,������7���_��`�<jt	*/��K������N%��B�a����;vZ�@/5᳖�{hZs��u����x;��$xsJ ���h�[	��o\H��c6����EW�ܽ}H�Z�x@yM�s�v�&A��ږ��kr�֓u	}e�Eg@�p� S�.�Ӂ���~J_��K�W%Y%�Qs��o�Z�hf�k=b񁶐���MbȻ���Q�N5-g��R�F���@������W�;ƍ;�]^�k�jX.|��&���K�?qg�"�*t&<���O0FC_l�FJ�ȼ�������J���J���'��Ԟ��X��������^[���V-h'���H�3R�k�q&[P�l��,'�9Ow��Ke�i%e�� W��9�RN����뻕��h�f�Ro{�������b���dV�����k��=:�;?GqN��z��u(�k�Y���"�5�0a�=�M�bI����)�o��%��h�'�G$��ƪ��FX\�!��70�zDq�ㇾ�Q��dd5@�6�W���$y�P�|{�GRao��'l��
m��ܵ�^S~�)�#�Qan3�߻��]�|%,1۟��<����d�}�)�A�����3�.�3
��ȏ`o2)���@��g>*o�e�lq��9��L�ǜ��N�+�l�����): �Y����K��`"��Y��i�P!�R�J$�|!/�89%����U��rp�"A!V5����F��*�m���${��a���kE�5�@}����Odt)�߷���8��"���'go�J�3��?˸dv��Ǟ�(�Q��W���=v���Ԃ��b�j`���a��C2q�����хp�!.��t�C��\ �o 'B0�΢��9��/�
r4%�i}Y�+�G�\0@z�,���-'As��ې.J��ظ����j̳x_*����͑1�M��t��/�P�g�! ��C �-b�Io�]�����?0�y꼳q~�{��q�K�B5���>_��߼�f�l�C��Q����@�g�����b|M
�5m`�T��R��x� }�my�F��,+i��2��q��I<W��(�V�U��x��]�m�>��π�mǐ������uIɚ����j�f�6IRT�X�DZ�)��=�ʦ%� �M�$��?wk���%-Ml�@�"K(,�����/��W��zf�c��L�<Q�$4## UԱ���چ���u�I0���0�"��
R�s�!�1p���K8��ʑ��G����B,0��np蒧���z�F� �6�8�;pi�gNq)aL����;�� [1-<� �&��m������*|l����ߓ��L:w�)V'�,����K���o�K~Asۤ�Z�D��=�M^p�>�)�f�'�vދ�Z��<R��b"�tiS3�8VΪ�%��#����]���*+P�.�Y�`:q]n�G�3g_�ѯ�8���<IZ��^�x�fE�D� x�M}�?R�/f/�� ���0Pç4,�*����X4��װO��k�,��1��݃B&%PR;��ތ����3_�bi�?�
��w�<��Q�%���
f��P��R���
�m����6�������ކ)>$?[4�|;��\���=fa�?.�W3��6V��^����ц@��@��s5�	�����Y��dl���[���<����ZN��k��2X���-��5;A�R��Ci���]YM�22��-��r9BV�����]�X�R���]��"J��K�Yd&Q�H=��r�\���1�����V��z�Q_/�5�[��T�.t~9�a�J�����Z+ߒ�M`Cc�C������րg�A�M�E�С�3ݯ��0γB��'�9��5��F*9IQ��@����I��x=�����8K]3�",מ�8�@���G�=�I�)�1�Cp��V��G�ߝk1J�?����_,�1�œV�M�i�������ВA"KU��&i�X�4�_�����8�2xc�������'��׉��$@m�:��H��f��MHxU�>e����`��t��jw��0�=A��KI��p�4d��s���E��j�G�,^��e���""d��ʉz���{ԟj�?<w&0��ay�9r��h˿b��3-�kޗE��A"E��O�`� �	{>qyYC�l#ZJ��bL����󳏢��mV[�/O�N�p�,�*נ�D�x���x����J���L��Chyo������y��~֭5L:qTx���J~0��E����r�~���*�P��!ò�~X����o1�C�ǘ�}���זH�F5���fU���"�@ާ
���m�UQ$�D`vvv=8�kA/_�����M$��&R���h�k3W��?�
��Cl�Xl���u�x�1� ��Q��:pgP_C��9n7�l��g�Sx��/
;@�R�\
�-p$ĶL|�tA*�A��g�"3������ ����	0-�fLĶ���@�V��k�EUfq<�خ�G��Z��m�D��-��$3X.d�R�L=T��.R%�#�?1n������>�^"w� ��9w����O]�hI���e��c\�P�7��^�޶.g�8G!�'��O�>��S�����[;0ʹZqy|�xt��Ђ�ss	s���S�x�Z���d�������G�ڟnq�4UdaU��ƠI��I�1]���x0�y]�K�]Z+��Q���il�^�O|8�ҼɑI�g��:ض�bfFi���}�
�)\3��x�z��[�8'k*��Bl�Ԛ�cX��uA�w��'ة�I��>~�PG$6*���D�7��wt����F�Ͷ0&9�I�5��2�3���3e-Kw�|3hm��Hhp��Hi��$�q�U�@�p�?'�ͤ��v��5��*�6�I9�k��6Ȑ��̛Ci���̐�bhP�r�썚^.Cdf���v����3nzE�c��,J��� �4��K���5�G�F�e ���i�&n��1ɼYDL�`�Z�mH�Z���!M�ˬwm�3�d���MF����i�B�j�4�#���:����Wu�D��\�� \=�W���<�+�qD�w���x�Gc	�~r�LG%�1���P�E,k_m�1- ��T�#�ܧ�����Uˮ�E�J�pF<�����}T�݋�V��ԭfY�/����PA�c�p�a����n4���B�_��:Ծ51�����߻l�v�ۋ4����4|m;�M��30�}`�۩u$r��H%�o'}D�܋����5Z�M�F#��+Z�[�s�lϫg�{�����Z%�1Y`j�.|��X,M�Ø<2X@=��˶K����F�x�d�ܬ�N��-(N/����͖�2��W��3�S6�z��	�1ܢ.-�b1��sO��r�YvW"fG,N`�L9Mz��� <1�z1�4�J��a�S�$��"���W�n�������ݱ%#��y���C�U��J3�Tu��찵<5�#g������Xl�q@D�,��I�\�>F.�%��J�l�@�+��5f
�K�bk���Z��֭J�*�e�w��i�5�C�ǔs�U�����_�h@��L�i�v�ɹ�>Mta�z��+��Ye�z�r��_?����O���1�B�,w���c�@���`ucx쩺1k��F��k�߭U�03��:��"㥋�uG�ܷ�9�ɍa'~Ց�FH����g*=8������!��]��8@W*0�P+h9r�`a$"b}_�_��F���.��6�McW�3�P�;~����M�weV�A��]S�4�3�`[�#rA�ukf�s�K�ƜWkU�RD��U��K�+"o�>y8�1ʮ����{�����!��94�J������z�[0~�p��g"W�F�C�X.m��UP�3A�u�U�4���[�h��,ʙ��[WK/��,Tg'�n��;07��$&ޮe_p�9�<�~G�Ng�o�����H(���J1��b�$� Ps�.t*�&⾸:��t���ᙐ�B�a����_����BJRt4�	KH�_au�x|���.�}���ǟK[L�Xz��\�y��!�����-b�K#mW��`��0�K�o�f\�!�@�lk���y��A��l��5bUa��q.ێ�<��y���e�<�~-M�;���dd�8��؋���4Ȼ��)��"O|�}aa4_ᆧ���6<Y�)�Z�w�&��1V�@���.)��N8
N�)y�����܍"��,�N"Y�n^�.����W	U9NMO�M�+JU�N�����D�p�+3�c>[����-C!��Y5�m���ބ�d�����h�x�2��ꊱE�Y"u�mN�Vڶl���w�����Q�[Hs�[�T ���_$��Ա���� ��)�[�bv�z�	t�H��߱]�i��3Fm۪r� ��K�R��k�O$�O���q^Sm��_�h5�8�%����zGM����G� ��;o3H�Eں��t�?>w*`��v[��U���/�)���:r��_�����G'��\��V�D�����?w��W-���W/ΎD��2�(��,$`x�>0�Q�$�是��u͑X6aB����Un5�/�)ׄ�F��yc@�t�O�㜆t|�9X��z~<o۬ouh #f��]������wy���͊�s��������pV�.��FK�z�x���=]�{Fa��%�,*����G�wN���穏}�g�E�;�O��]�e�Z}WmpҔ����.)���l���w��!ׁ�;X��е��d�i�d?���������tm���ų)>���K�מ��gl�D� 3�d��&�l��T}�T@�U�g-�yY>ww�ȸ�k.�_J<ë	�9d��z<i����v���%�K�>la�i���R?46FW&���}�V6%��1�b�~���W%W��v�%[L�}�|���9^?p;qq:���e�!�� ��l��p�A�p-�q{t|�~�˩>�Rà�R���l��kn��rd�4�F����W����^�d�R�ܿpa�O
��m�%�w?:������=3����Z~'1��#���ꌬ�Qe�.����q�˃G�O�u80�������:T�Ȅ�U@@l��.�q�m��/K'�ڑ��%�c��K���h}o��	j4l�m��k�~Ee����f`�����[o�����0Y[4,Z���i�L�r�	ՙmZp���[�PqX����-xjFZ��iPO�XPv��6�iNɃ�J侮*yݛȉ�r�=xvא4c�I#�� i�ݜCL;��]�,5Z��5&� �[ޖ�^�t�Pφ6H��v��d"UN�BG�A��!����ÌG�����Ȱ��� �RS���ͷ&�JR��L[kG�[�a�:�^������U���?n��w�#{x�Vj���,$�O3�i>�{�J�$�ǳ)�$���dK�ϒ&�鸵�^};\��1�Iշ��t�gy�Β]����?�AV��}��� Y�9h|z�z:���'�B���z6B͍:p��	< �-ud�S�j��@���u��?v�(Z���+�lA�c���
Lt8�5nU�AD�Ҭ�������&� �.�Ћõ�s�|s�H����ө���]��\:'�4�)�1!A��T[��Ze���<p��QB܅ӎ�?��&�M�}$H����������|"BL�C.
���dNu����ep��>%��v�OP� ��4��m���EU5�A�)Թ뺾j_�NE�t�f6�^2�/y�3���>%�N;��������foº~�o�4{��zP p�ռY�ԏxv�c�Ё�?�L��Z��锦�H8;aN��SZ�ˢ��x7�d���,I̱��m���i[�F�(����#���K$��{��!���L�(=���*!�z���f۶���ȃ����:�n���S��5��?����V\+E��߽�N��M�1~��E�׼���Ԗ-{/����n�A�k�+�8<j�/��-2/�r��*=��$�y����8j[+X��7�n�9��n�?�u�=��T��ۋeDR����6V D�s���X��O"~u���4�bbn�7XP(\/[�k���N_�L{��r�2��B��S��,�J=@{�g��6v�wX,$��v��a���dT�폒�v����?��y��Ig2Z-�ĳC��˟��ε���x�߹���9��jR�S$���d��:�n���'��\vt�ۀ���YRj�y�!h�]���8�O�bL�#�V/"6#�9L����*>!�w��fj��sĴ<����
 �����R�!}����i�%��[��)��ɵw)v����ى����gd�c���4������՗jLd��!��(��m,�����i����͑3T�:��
D>�p��Yr%�m�3�i3>
���$��o�6.�4�����BR�9t7�C�G1~��A]���uS|1M��ɶx鯹rE���;I=�~�1/�I o��R��I�����e)�	�Γ���Ӵ�xm������r�/���ΦR��A<�>��h!��p��>byPh/�^���hAS:Jץ���g���#�Ԃ�q��?1�0������ULGLwj�  ��%�������B���N��;f�
����P�����P������T���RU�:ݳ�ðeU\N��]!��������k/�'?��\�x���ؑ�����'5'l��:d�6g3N-tG�R .�"t�k�i�4�yڻ_֫��W�م�������v#<Uw�1&_��f�h��g��	�/E�Fg��|�e׉�	���6l���}��kN� 5�g��0#���{�a0[���"�1@+ �$H�hۅ�)�OI��|.B���ˈ��w8�|���j��j����u}�+�m"}f���D����-hN��fg�3<��F��`�����i����Y�n�Ʒ�%88���y�@�u�x������*��Km�I���.��_]<�?���QŚ�������e�9�M�����A���W,���H	Y�������WM�d/E���(�d�O��xI�8IZ��=��)/��l9�X��{�B��eX~+I�g�+��:0"Q��ޣAvwz ���3bi���z���T��T�"W��5�(�^9�]C�i��H����,5ppPoN�� `H�8��0��Г�����8+	a�;
����E�$��n�����X�Ş^i�6vU� ��UQoT��������z�Q���OtI�O¨Ul�gߛ�FTA+9a�+�Y�@7<����[�,�ԩ3�.?r��8�7.F����8�.�3hZ4�1/u3Y#&{��%%�*��v	:��wx�%ʑ����^�So���i�� D>W�x�x�Z 
T���z��w�
W��4Z��$�ĺT^^ �*ǞCx?Pb=���M��Cݝ��9T�� $xD�t�'�zJ�2M{�jn| t�F��p ^QneY��|q�58�,���doO�%)��f�m2�T؃�.>��Aۏ纪GO��e��׉�h��c����۹����[kb��%�V��؄8I�\���X][ �j���R
B�nJ'6Lݫz<A�����+{�r���j�����J�^K�X�<*��k�	j��Q#Π���/����C���:+���S-I�Q;b$E~�>g�M��I������c�<�M��D�\qW�s�f�� ����U~8�UJH� V�5����ø��Ϋ-$W^�lU?���H���u�E?���mR�x��o��+��&�m�����km�7!1j��)x<t���f��V���^t����O�ז`����.�6��5�����92�{�A���NAH�4�Z�c�V�G���MWK:�Y�L?]R�dhޠR�o��wG8ֿ�cs�9�ߟ��ăk�r�B��
��+M���z���^C�H&<���L��:�p,~F�h}�ެ�(�:D�H|^���8��/9������7�I/v!t<LmE5�3��E��F��ڿNN�w��� � $�lFQ֎�){<X�nźZ$%�ܕn��)��:�m�J�ⳋ�ś� oVkF��=%�j�(��dd^�=a�_L{�ԙ�a���F����3}65=؀�$#6��"�i1��z���tн��F~ƴO�8T�p�e圡��v�[�9l�����)>���� �M{T2F�p7'��^C�t�M���fc:Ӣ]�:��-ŷ����Jk��4P������k��/���T#�4��j��
�Rk��>�7'����;��C�Ge��,�j;���c*�_��Cĉl������J��H��1X���E:IP���w�#dcF����0�A~��3!�M�,s�4�V�����V�D��.lص�HO�q�.�oL��%�.C���`�w:UӘ,$*�JO>V��f׫���w���k��Y����	�Q ��V���aD�}&�쁕t'Oe%p]95���(D��$3=�E�,�!�r�>0Z Do�""��KHTp���;UIP!���A������v��l܊��]���4̀S�����csM�C���� �tf�vF]Ith�5xM��T��ÿ�ح\����wsш1/N�!<+�����As�F���A�OH/� ]��X�<wU`$��m��@�w�dM��Ԇ�ҎZkS���q)#�����I�^��\a,�$3v�d� &�H�p��~�y7ȳ�9�Ct��Fr���Z|����kd
z��\a�9r�,���ޑN���2#9�~5�/ɧ�����AB�4E1�VB}(6�k!��̣|MjX�+(�D�f� Vu�!�\cLu�-c����鲡���Zc��c��;��͑�@�3x^�"p�T����؜�R8\k��qaU�<��W?��V���"��~3)ǧwAa/�O�ގG�H�b�t5�O�����X�.����z#7�]֖�}��T,0��a"�P���Bm,�������q�Ļ�O_
w�t�0ŎgH�j��<*�iă��t�1��)���z�NKyځ�'2^��b�a+��T#�A�2���N�{ c��5����+��'aEc� y!qO(*8�C>�X�M���L��t�4��������?9l�<Son����h0p"FC�H��?�:��5�t��܀��=�����`V�G3���pq�sN4%�S��d`O��_nԊ\�Wh0�H���o��D��;�% �y�벃>����o����`�~��+��SW�ȫ:-\�rv�M�'��]�c-���;!æ0lؿ�*��@2���s��ʪ�Mum	�jm�?��Q�݋za��S����V'+���,�����T�.�W��_f��7��gp?�<���;�+� �{U�f�NB]�ȿ��hn�v
	ܓ���� mSZ7��4�)���h��oS�" 	Ɇjr5/r�6<}$�jh��kƛ鏺ެ�ҕkls,��>i��������"�[��2C�5w��ɀ3���>>I����Ȅ����B���ػ���]�ꯃ��l7X�xvO��E���~�F`-J��.�Dr�$�1����DXJ0ǵ#���ş������,[��O��r�tǁ~�3�"j]âKs�Ǒ��	+��h��~q/���D��.�	~Z��g
�~�'f�䰼y��WO����!a#s*�	�Y��5�����̀�D����3���s��R�4��z=5�I��K+�K����ힴ{3"�dP����=��p�4͍������a:�
�4@x�= ���	gv� )K\�����e�]-7b���*���',�{�&hOW��C5"k^Dp�:�2��@Ϝ�cv><BG�:h��?i�#뫜Dꮠ�8ą�
В6��j8:0���|���\�
X���w�ģjG{���!rx��g����b���Hf�������ĥ��l�F݈ �ҫ+�iE�;Lα�6���O���-!2�f1������g.�m룯K�H��������?&�l�w��c�+�\�2/>r)�9`��.^���G�u� �6��%�6'��GM���m-d9]��>�ߺh�l�����^ID��˗o�8�=0��Q*9}���o�1�?��b�k���ug��k\��9*�R�\Y��Ub�����~H�=u���[�-;�?�/H���X�{����*���O�>m��S�����Z��@xrX�2|�`���Smӄ�:���8ш*9�܁'���][��nK�UN7I��l��m6V�-�V��.��\^�:�\4A���p�e+��lmV���0@	�o�2f[���m��	����+��\�pm�U�ђ�>=�n殬~̷g�笤��cP[�Y	���P��b��B�޳_����#<�&òg���H��%��uk~�}ʠw��x�lեX����-2�V��Z���#�8���ȝ�V���jh����2��3D�<8�\�5+��JL�uL�Z��Jv�.������(������\!+�d�`��R3w1-�Ł�,�N�Y�-��j.����|aj�����}
���-��N�F���g���M����q���&�oCf����NV����W}�/e�<�,�՝�b��,�H`Xγ���8գ�"��l�Wx,��u����OpL�r0S#����[�H�<`^���D��+�F�.D���90b27��5P���ss��5�Fb�t{7���@y����p=�v����p��f�3=�@Eb��I<l���������uܢ�c	�;�}hG��h,L�&h�jkP�u�`�s��D���;�6öX��J��}�����k�gQ�Q�q�k��O@�Kݳ�߶����w��G]�~A&6ɀZX�35|.�e$8���Rj�Q��Wi�^>�i�h�=E�Dk�Y3�*--���M!��F*֑M����c��e��d)0�#�� ����6��/��\̆�Eu��^\�v�r�������`#j0-!�P3�3�W!KJ�
�� �}�8'af#�[�CO Is�m�h�hL_~{�O)���� ���7ȱ� ��B|\s��51ם�k]��#�c�Ҡ!�S`i5B(��5��&�3�f]�[��!��j���U���{�"�;eҸ��9cjݤ���n8=v�_�K�86�*.Y�4��
�q8*�h��������k(�P�@hZ�UD~�IQt*�E%"�][��[��>w��0�m(��/j��da,���J$�	=�����&z��)��Vl�)7�3�H��l�aطh
E�
��R)�d0��H��y
��e�r|>��2A��2U�(6Lz)���*�ɫ�[� �e�U�h6�!�φ7J�=>e>�,�qU9%6��4�m�#��ܖn�Z�F�1?�ritI�yK�TK��Gj�8��st�)cZ(o7���(t �	��4%�x.1��4E�$�g4�k�<��ۭ�O���r�	�d�ܸ?������"���2����׾���D��������WM�a�U���t�?���a�
@�j�ȝ��\3�y�Ŋ�����l�Ǽ�/�F��Zi\�t`G��z��P�;@��_L�)l��΁d3y�7��>��^��BN��Z� �O��\R��H��AL��_q����&g��3~+u⧸P`�L޹페�,�'�I�g5<�Z"��g�_M�iEd}�Dbђ�9�σ��ۗ@�!�;J������
�<�I�'���#��3|/+C��#���쓢��X+�Σ̑�]_,"��c>!}��r����T�P_'�l��!�m�p��e��?x���OIX�1���4����|e�|����7�3�P�i���#ˏ#�v�Z�.#�f:w�ikx7ig@�_�f֦�)c��d��De��ޑi59n�Nâ��`�`�ĉu���C9?`i�y�
�w���Md�1�2��C����Us���V��"��~-z�8R�	���tՑ�yb�M��-ܝ�!a*�7ՀJ�����o��i*���C0��"��)|���,J�&x:#�b�fs�;�D7o�䗮�ZK8�*mH����9�k����UB�Y�ڀ�z�t�E)��6����P�j~%|��i�9��@l ���e�EüT���%b�Sч�������h�����:+��:�y�d�t�A������$�BY���[z>��b����!�ɘܪ������V��n2�Ŧ�OHSQ"s�D�)R�>U�^�E|>z���8Ê�!l3� `35?�	P��H�i�B~8o)�H�J�	�+�����}�܄�4��	k	033���#ƉpD L���g�;�,�����B�q�kp��1<�mIq���B���$�5v1�t�񹮔�^ǱjC�ΊLf#	spYWm~�o�I�X,�Ҷ ��*���E J��-�ԋ�d�v���~��2x�Xb��se�rmH�(��H�1vofǿ�n5�ܵ�tG����)�Z'������v�z��R�J�^���o �����/��)��K��H��K�E�<w� g���7 ��_'|:,tuo�ݫ/~dL�z�re��P��K�Dp&�>�\�4(G�8�+>�:�K8K������*ur��Q�m�$�(*'���T�.�&�24��%��̪L}�w��bTؠ�Zw����	7nR����}������=���5�y�x�P���qv�S�`e*:�s	��暅�0=�#Q�nZC�F{t�ɋW(�e�l��D�'8ω�]a���I.m
N�~H����>�����(IR5�n��#�XAҥ�Ի�F�+����2	,եJNrJ֢�rY~�;�-��'k�v>j߷�c{l�MT��x�ҥ�:)�~���,�{�q�L9)zݞ�k��7��[�_GDe� (��B��,	�����nv���n���/�=r�t-zr�z{���UB��#j��iSm<�F�2�����v8$bh��܅����8����-�\���q!�x�+%�Wk��)?k���
툐�Te�aXќ��Sx�ɲA��IABzA�2��#X}T�JkI	-�aܑ��R�T��]K��*<82<z� �+B���1�1 �|���א�,Ni	��3�?��T�ʶT�0}�d_:퀻]D��Ц��7�����,@��70k�Z������I����B�<;p4d*����Y�)�C��r�����)�g�eT�YR�2U��������[��Jp��}-�9�n��\���kx��q-����������l^�ѕc�����z�mvAȐY1Di���I9j�mV���W�|�G�e���!�������f��A�;n9�+�u�x�M�5�?p����^�%�q0���㦎(������.�p[!�#���x�c[�3��h$$���m����yzxF=1b^'��d��Ŭ�ޠ��Ah��ë�U�\���c���S���$<�b,�l����N����Z�DE��ݖ�3��! ��T(#����	��U�`�,K���O!Ů@��pot��O�PyB���.$r��j��>����i�̩��ea\�L`1��7��+���J(+wg�a�e]\R��w�e.-)�����Ȧ�>�����f����\��pȸ��V�@<���C����@ rCf(�qͶD�_�@<�ɴrW�������l���&f)=|ӹI���XM	�V��P�:0=7P˂�U���N��"喨�%� �n�#jv%����88�2�V��n��qL\�58�^�l��6�-f{�|�#$���:uş��c������/&��uO�>]%JEE��B�t��Z�?�ϴ��OK&狱�������.�]+/Ō��p�s��sI��L�D��}�n��EOӇJ�c6�#l���3~�_|e47�4�ukyh��|�nȆ�$�(����o�h�����p�����{g�ώ�}�*B��J[��]xNGI�w��u�����eW)�Y,����Xp��Q}�A[��	��*���h�K0�vTZ��#^9���Bf�,B�>�����=���S`ڑ��S�Qƍ���Ec��3,{�Y�^R�ne�_���1���`��NW_�MH�����@�a�`�=���f,�vƟ�9z���6#U�g�_+}��|,�e��t������Ƅ�4NT�ЁEh����@����t8�����!;;b�HH~dq�j�҉�y�MU�p/�w�����)���ؔ*��Fx:��7����;�`M)̗뺔<Y��P|�$$]�\��i����0޿-s�����!�D��]C�����czWl5�p�>hp=��D��=R���KEs6�PiWH�w�ûk���A���s���S`���]@l�`�}n7��9�xB
Z�1����/�u�ͺ�U�G)҃a���8�����$3�X$�;��)x[����	2���വO Y���7�����j��ҭ}M��w�.��қpI���%��k>>��ۀ�6D��>^V�g�h�%m凣f7�;����� M�U�y�)Vy��3<�-��su�*b����U�m>]�A�WD���ih�^��8 uI���F�W7T׫�j�(��L�g�{�6��P1[�i�� ]2�A�X�h�up؏�	���T\� �?l�e�S(��+�'k?��K��|���`���m{��"��?j�*�8��9�r)vd� �*�#� �w�4��rR7�e�G������m�5T�|eϼ�Z"����l'��%H�p���7��X��FK�#67v��\��A�pN�@h�7�L A1�.{�4x��\2fa#�߇LR��-_
X��0��h��r�r�ţ9��-}��$+C�%���YXFnX��NR��9I�c����_�R�$�	��a��z��4��$"rLS�(� �j�1f{;k�����	��Ԛ�A]����p�t��d�}�_�~�xdvgn{+/��iT\�rU8�y�kq &3#����=�&#�y�����塚PK
c� ����J�i�Hiܛ�fy*0
F�_���*1��Q&Ɠ��V'�mޮ�ٴu�~��e(�Y	T������j{I6��`�79���/�
�CE�������<��=���4<bK�������4_���3d���D�	�23���Gj�ǁ$���w�-�#�,]�����U��ʹ�� N~C{L��A[�������MZf '�;���-�@�͐�3Dbܨ�I᮳u�v֘P�Wp