��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��Ȭ�SWC
����ѶKP������e��' )_��2�.�I��Z����)��)+����Oq�	�X�$o�
�z�Z�G;"��B{��A�A�5�Xq�Ωm�Z�4zbv^ӭ�Kj�dy���V\HG�P�uP������[��]������%�Aiw�����)Y�;���iY�g[����m,�	����0������wʐ�Vf��C�<<�uE5���8�t
i�婰�'�j�>�۸���4�A�DY V@D�`��\k�ؙ6�Z}�f�%5tǶb��I��r"$���MΙ	���\6���>��*0��k$~Ѻ��)��I�Qp]��/�.�z�_0(B^��-D��E�<x��" ��k�YJ��%�$8Q��4�R�x>@n�\���g�ft.��7dνK���QO`�Lp�P��9֏���jm�\s^��&v�p_���6a���*�K�s��ȑ%X�z��>J�c| L�E}�TC���Dpv�e�"�Y�����ڔ���ц�������}ܷ �N���8 � cէ
{��5��Zs$��I�K���jF�ui�L�f������pb����Ʉ�������6�H'1HP���Xwȥ[����>��8㩢�}�T!���*�K�^2�n��u�:Ƴ/ñ=g�{R�$��c<���=�iB�Kk�z��7J�v�6���D�\�Z��_��Q����f�z%�v��Ă7�!���=�0nk�r��6K�ܟ�Z&�17s�}j6TXa5�%�'B9ɿ
K*�������]n�}�E���Tf�V�s��c�QK1
���h�$��u����D�h�;S���9�f�2ԓ�l��h��@��K}�	:��}��
W�e�#�N��6lKEI�L��Gt{tYMZ�Hq�\��@v���I�VQ��	`f�����a���FT$��ldٕ	�,ls2�jeZ�iڗrW�g=9�}�{�O�P�P�i����گW�9��߸�r�w�NqƑ��5�aY�t�Ɇ���b�a/'��P�Kq�m` ���E�(�ULjS�/%�|\�<LN�n�
�H�3�#mh,D�Cw�|�ۭ��_K"v-��O��E9k~��d��@O����4�1)+��Yө/��)O8'珚�4Yx��]�O�L)��6���{? xM�~Lʛ[JG�D���>���唯�����$m���M=�:�T�b�8��D(0�l�8`�f
�W6=R��^�.ۿ��p���tX�Vc�`�Jo#d� �ρ��]�� rz�0q|���X��5��H��g�ǽҊOR�'��Ƅo��?'mj/$�@��ª����`ޔ�n��a��:;r���-~�\���/586X���7>��y��n��Ԑ� �+u�nf�r��Y&;%��A���͒(�Q��f�F/$5�侎v{�/QQQ>nB='1I� `p$�u�U~-F�GX�W��۾���+*��sB�Ɔj�`�sB�3X��aK����jQ���tz��Ge�h�>�]l�O�wXu�i��4b3��F��F�> �T�w$V��hf&�.K-�/�O��s��CH�J@Q�}P�3��B�S����l��Y󅜟 O,�,�m���0T�I���RÕ��>8h	(��UD ��,�q0�%�������b6�'6�\��#cly��Joh�T�1��҄K3c*���sˬ�/�\��b#;x6�����X��`���Âj�>e��8~�ٔ!<I�����/e��c��G�m���Z�ǒkN;��I���r��e/4�y33T�J����R`��Zyx�E:y��J��j�a5�P�Ɔ�^����I�?@�`�%�$�~��b��[3��j�I0N%Y��^��T�*j&��c	�~���PF.w~�������\��{���F�q�TMr�9���hx�"b��vʸu˥k��
���Ʊ'hA��(X�q��!�m/�Ur��^�J*}ۭƴ8h {	��k쪇TsQ+С��E���� �P��/C�Z��eg��%J��҅���1�[�rQj��鿱</�Z���������u�o����y�4@���5L|��̨����G�d�D.��f����k�F�\�$�ɠ���2�}�c�_4�.�A�/�0ŻU����0\�&[mmuo�g	H*�0��Q)���E��%c�����R!̨���d�v ��V������������r��=�d/�Xw���Z�K�(�s=��3��G �vh'�^[8�̱���4T Tw�m-�Vۻ�Q��g�g�,��	.�/M0G����/ ��a޽���_��~P��!�D�0c�aқ�Y���d�S����9D67�8Lf����a�|@S�a�� 2:f��J�Jhn���@	V��)�kݨ4�?�G�Ʈ(ϼ?mĂ��bgR��塯���>U��r��AX=��+\���q��ow���cr�p�R����X��*4��a��t�A�l�����4t�� z�t��EE�K!�9N(�%����F�Ne�-���M5��OR�
?�ͻ��E�r�+���( ��j�ԫL�|��p{Jn�.R���[�EA��a���"���aǀ�aɨw^�
4�{�Z�	�.{X^|s�t��r���踐q%��Bv�k�+VS�Џ�B��T��{��\��� d�#�����_�����7��v�z�PH]��DI\M,>��J�h���=�x�����4�=Yg9���	O���l/���L�e�£MeG�#����\���ć@��4MzbB�-I� &�!^�u�9�-O��?�5�CArgkG�z}��0�5��K�ZY��/g����35Ԩ�x)�GQ'M蒵�K]� "�_�\%���H)ї� ��o_d򦫄� ����S���c�Bg��f�>o"$���fz7��U��&��d#r�_�Q�o1���_O���k�^q=U1S�H��o�w�S+�� 9��pJއ�܋�f����!<�!@����~��tx�� ��_� ����4��r<�k��J��m�ͩ���Q#�c#���I7�ۨ�x�:�種lԖhcQ����x\O��^��A�9a����P�4y7��o�4^n��|� ��J�^A{K���2ת��e/I��D,�q�+�x3�h�<�p���-a�Vh���]�3N�@gU��i82��^��E:������	�ˁ۶לX��k[��}4�s�A�L�/o���w���ol��s��������@�2j|3x
#��zujq�d+8҇����m(G��.n71 $57ޱ�){�H�\8T:��2q1��"��ܨ�C�Nm���.ӗ�u5�������#L�+���o�b@��6<j`��:;�>���Т�[����.&C�Ft�S ��P�Ϡ�_�d�)g�K���b�;@���G�����h��p:���z`G�s����֭Ɯ���J�F�@�9u$���B7�l��Ua�E�\��W�yKn̍�qF���t�q��f1}���|مµk��E��B�;Pb�-�A��>}#=����.Peku\B��'���Zh��Ow�5��Gu��b>��tnɸ�ꮪȄ���&Xൈ����L��5�^ET��/������u>�NnLO����Јӏ[a��q�O;2˅��-|l�6�q`r�sƎ6����7�>nn;��yA����o�=���"?=�H�@��C��p�L��Kؔ?)��>�Ѷ�$g�p�R@	���<��vCY����L��3�%\D>R_RE�EG���1�i�������o׬�������-eKX�8Z[�̾Ɍ��OԬ�*�Z�^��Y[u��Pz�a���̒����&�u�%��;ʐ"G�����&6=��V:9�NX%�]��2�$��)J��T�rb��2�4�362��QC��!����P�^���k�4�Zd&gܥ����+��HI���ET�۠f�[Q��|{f��M��:����}{�^d���0�|i�nX^��a�Q��]�k VWM*6�I�-{Q�?F�ꎏ{�0���[k�Q��*��7��{Zє��]�K��xJ:��)/�������ذq?c�'[ .�p���;�A��CL�5P�w=FQc�n��e�EBlj%p�R3�4o1|��㼝o�>�P��:��Qy��ؤLow1��d�p���f����伩I�b�!Æ]	\��C�ŀ2�VEq-�xLM�;��د�ED�`N����~�c�H�,�`�e�~pmͣX�_;�'����?�X\�P�fd_9^����+�K��ȃ���&p�!h�	BJ�%�>h	9�ZԮ.���|�SW�/a����j8=C�ͥ��%��U���p�8�Sy�m2�lc<S5|� -q{]��%�`�?\��V]�+�8�5�\⯵�U�!`���v���<����ݑe�.�k������#
�B�:����L�y@tVJ���� ޵�s�����X��C�X�C+( �-I�"Z��cc�O��R�U���^�'T�0��~	��d}];�1Y��BJ`��U<�CS�S�s{���c��X���!$i;%�dXkR��'�oJ���[�3=��szg���j-V�㴾AuT�w��~KP�tެ�b��W���g]��F�2M�f�R�����PW��c�W[g�:8�1(�r�o��L̮���u���_��j�3�B ����&q|�Mt5��SQj� oX�� ���"�О�1X�-dAl2�lhKJ���wz��a>�����;�8�$���g�;$�Ӏͬ_��>Gx��0�6V*��m�o\k=���|���էg5���'Ǧ2th��T�r(B<訨J@� W��\u��SG��l5��0H� ������4�\�#:t5���@U1m�Czi6�0`��u�g��߰Й��5�u_g���[J��ַ#=Z���`yD�����
tf��<�'�-��1`E�o0���d'��kS�מe<�t�L��V˓�E	~�����a�e-G�®Q�#iW�8f6�l���L1�G�r�V�D���A�k�U��a��Jl)r�QX�\w��w�F��=
u=�ƃ��y��qV��s'�w�dȘ=��(ލ�"w�Y���+�ɯ�4(��@���>Q�pʦA�&�*�2�T������G�2a�6ͣ1����/�bM��p���+S��kt�Ơ4�Zg���Z�����~2���!�T��E�X�� �e�]y���?�OvC�ܾG��5�d��b�*3Uy�RR����-a��I�o�΃R�iha�~$�(T�xDBy(�&��v�l��L_.�oo�E����>�qwF�s�kKX��w8LS�j �1���~��~fu�Z���e�Д?�]��ߛ�0��ZCL�;�*�0\��s�����2���M#�p� �?��sq3A��	Fl� >Z¿h�6�{�(
�2�/z��3#��d	�rPn�y�P2a�)ÜZ��%q��/qeNO����c,����*lT��a�S���"�_��2�G����"�>?�{L�?ΕM;��6�ܡ{�@u����c�j#�)�f��A�M%4��t=R��^E�#g�/M/��O^��QM�N:}����g#Z��m3��r��\���f�_&!��Vj6s�s�����'�X�(`�x+;���ǿC-d��E�޴�|1C����e�HZйQ̲�+�"���s��U����Z����Q�9�dK�fY�l;6h�ۓ�O���m����嶘5.ؔ4�Ĭ��빾T�7{���UY#��^&�ia�	�;��ڇ�P��P
r�fP�=������.'�&�^�?��Zy����^�6�EG�����י��^��D��<ճ	����̵Y&K�ɓLV@H�Z3��*L$̈�tIxk��o�����*�	����ҁh�?8k��jQu?"F�� ��A'2�Bj��v�vy6������M`Q�~n�/t�6LkQ�*,�@{fT
Ǳ��l��ID�ŲC_�;䦋v���B��s�#�h��2</5&���/�٧u�)Z���q
��^C��r�~�$mS�P2�b�KJh�F�O�?�Bw_enR��V�\R��*b���t�;�;��~Ш�Ú�!�=�u��_�+��j`�%�%P_�~l�T�5=.��&4����}�ީ�9��!���^�#.��7�ݭ��y?�?�G��:�51�ˣ��*b�J�ң���]�s�s��HV
��!�T@Y�w�B�����/�Ia~y1��	9�w�	9�6�t�V�8F�&�ܫ���1����&y�M���f8eq��om����p�y��w�V�lT�v��YЙ�&x)@��$���0���x���g��n��w��v��C��l��}lB��<�P��L�m#��}z���!�3۴?�x>�r>�ZHҟXj�R��w�y	���
�8{OT��ۦ1�ۂ�pf;�]��f�aĂ��X��7�'�Ʒ�i&��S�p��8�nR�j`�'��(6�b�L�~{���(�iU�~����&��A�u�U�~��l��=b���Qj2b��j�b�d�Y��'�'ȩ3����!7�ja;m����%	I�TF��+X=+����R�<�T�����L�uI��DX-"׷�̀���o�@�����	�3:M�3[��C;
45k��S��{������1�u�9r�%����֫�;�(��V8Kg�6��(�Or�n��oG&`��)9��E$�'����:�a>\��ae.b1��_�ԫ�쭗z!t��|R�y�u��!�d��2��=�N�W��%�*��ްKw��9B����b\�=�䗑y��wU����h�����o�E�u֊�i������Q�F"ngS�Ý񄎇�ằ	O�]p{�r���]�u:إ�F]~lE��|EHwW��,	%�X������/;6k���
=FA�{�M�q�$�qe�>�.+���
/�����N������u���7)%��Yp��v�!'I~���F��L<�茜�uaB��i6�6[Zk��:f���̧j��p�߮ݩ�$����}V��Ѯ��7��Bۅ��'x�Z�ٜx7�ҍ��{kj�FW,��*�c��Մ�n~���r���\�`��
�vg�5��X��}�}��Y�?�kk�%��<:�!﨩W ���Ր��)|f3�ZeD��y�>�#&�����y���.��H|�]jFH�2՚u�qթ��gV�r�c����-��}�
}D�vO�������{c]��"����{w�4�L�t����+���ș��bd?/�K���B7�g�k��/��lBoENa��w�A��e_9cۇy紧h�����u7W,���%�N<Z�J��Ld���g Ŧ��'�*�ǺD��6��F4�i���u�ER �L]2���4�Kes� �Zl��g��}6ݜ1Hk5�?�Fӱ�wP*�R�^�/5U[9��\,~�=9�D]��U�Ty�o�l��J&�f��>���R�����XB*�iȝ�-kR�4B�h)�������3>u�4|�FI�g�R>1)�4⭁�uz��P��' ��0BԨ�����iFu�vii�7%`�1����&#�Ӫ�H��*��+Si��p|D��w���J��Vs�O�&l��l9ͳ^�~�_��"H6`��F�T{(ts|�sD�R����yM��A�d`G=��ב��Ȥc5�űg�,t54���@��<q�6��Gp��U=�'��hNw��<ӓ0,��&5�ah@Ҷ)�́Ӫi.CI�k�8T~֤2���z}ډ����RX	�>*�G%N�,|bB|���=L����@.��-��M�ν�F�b�â'��nchv�I����pl�J��YQ����p�?V��A�5��Y/�-�7��.�6��������8T�=r���|��]�dl�n�����UÒ�;�Ȅ9��F|�� ��*�]ch��aR0�	�4�67��f��d�M�}Q��k�J��|G��x����2[�Qb���Tݥ��|�>��=�`��g�p�qP�ex~P�M/k�"-��{���|�y�*6��7l᡽�9����?�ԓ�w�ˬ���k�l�v.��Pӿ���82ݫRP��s�	��t��A��2�v�]ȸ�-�Xg��L���f>�(�IQ�P�C���lf~d�/H�,}B��|ˆ�{ܒ�?�B�(FC�����!r"Y��4���`Dݯǉ95�:y�ʵ��y�[��~r���of��������b�F!���"E���];cs}L�'�6h�1�>��>�ζ3ZisHoM�e�J����[��ҡ�n��.��[Ce�T	(��Ƿ1�~���C����C�������```��>��������9��TCq�" �=n`�X!�폮�k�g��1�(`u�.o�泖H�>
�~q���V��ڿ�ӯ`����J�V�:,��Ɩ/'�`�S�r��5�˞���<tXLJKJ�i,�U��!Le	�y������kqV
(\_M�^F��SV~̋zgǶ����2���Xw��u�����&.S�Ɖ�3fT��O�C���1�OT��&�: Y�x��Vo�ǌ}1��zSf��a$K
<�⑵��Y�ʍ���X
Ɔ���37���&~���xZHJ����ׯte<���PĜu�;�-�fYRo��>�E.���C��bȮ�~��P��9s+�� �)�P2��$Ŕ%���~؂��Iϰ���jFQ�*�e5o;5��|`�A|�~��3��Z ��߯T��x}$�/9��]3Y���Ϭ�����A�kZ��b�\�K�tsxs���]���3J�ʥ@���<��B�[sL&��Mb���jPB���7�@x�\c��ީѬ������0%��ӓn��>Z	��6���s���E�����џ�K�w�Ɗ�k�Kd������ٱ��J�mP@d��agz�����sV��6���<�#�B�1d1,9��̌�|	n�ӆ�f������񋈟���:V��l�9m_��2^&�q߂ ��	Vic���օ�ز"�Q]U��^S�>�ZKI��yİ(��H���gx;,1o���7P��m�H$ʘ��T&4�5'�ZJM3��)��)��}�d~2�C"�|l/7D�zʺH+���8p�4��ĩp�Ш�nK���N ߕ�'�����c�������G�9 ��-2ɇu�-���LI���(8�eC�ij#ضx�kK��*�䗁�1�ظ��'����0�����C�"+N�^p�����q�vD\Ng��F��)� �\��p$��j*�߿��`��F�#T�%��E��\�)Y.t�t�_������Y�o�T�e�M,O�}��.���qYǔ�[����&Fby_��=5���h�s�q�-��_&�xGʭF�R�3��ڛ���� 9���::D�rH����$��+y���_�A=QK�����"��g����R��gS�.҈��w�����r��� j��H�@�Fm�[7(To��r���P�D�a�m�O�q�#Z��L��v/��\ˀJ��e�T�������	� G��(r�M ��ᓕ3QJo���:yH�5��a�;������m���T�
x�y2l �W�D��鱛�|��|3�]�9��	_m�!���L�h��,���}���1�6z.��<�Hu���#~ �;�w���8� ������l�c�^�ⴄڊ���Qۼ�i��:��nq�Q<^+n�4���Ħ:6�T��Iќ)�ϥ��v��T 7&�\ST֔۝��������������P��� g��z{h���j�����[Z���OCw:���DC�h�)��p[~����;�f�ԡ�֜�0�� ��y�DXܑ�'~�n���1Τ��ϙl�j4�>���3���`aH�4e;���S�ꟺ�/f���u����U�P	x_&(�ϩ%��������]���3'��>0����PL�Q�J�yh�&S����h�MuN��w��b�rn�5h�����b��h�G�;+Qʂ?1��1[^�mOt��%��6�f��b�]D�["��O"`�NG�%Ǩ���0����`�^mU�/U$! ,�9t�
���F���f��]C�Bt�����6kT������r2�7+�3�=��r�������l¸*�.-����"&�i�]��N�9:+#q���G���7�5�s�w9 3��G7�
������A�z���	��CoD���G�ʤq�Y2�6O%Ir�L=,��K�3�?�Ȉ���l �{�(�	�6����}�lh���v��!^���S8r��`�$-@�R'ޞ~u"͎ňm��%<�)֌�b�Μ�'d��b��g*>R���H X^����6�u��=0}W��H��ުO�526^p�3e�'��f8%p�=W�3$�����>u�o[��Ʒ��F]�e�����s�SZX(��c����sh�R����c�n([[��=1/������{�#M�=W#gQ�#��cﲊ�<��{b3N��$�����p�!��.�`i�wr��Te�6 tq��7Z��wf4��"�>~ZK�n���ת�����&��s�/���o�����ጬP��*+�5f2�-�Ml���ij*h�'�Zgw��������Y��WL�t�@|��s(�P�#o��3�4��)�Jl�`��t�a�I��c�� ��f�B��8ZT��J6���VX3t|�`b	�JK7C�p�CD�l����,�uO/lj
�LVA��ݵ���V1���+����	n�|�0�C�3*�7�҉[��*qU��/
W�mCS0]8�!��=[�m��D���srD�Q|C,� Nh��9k+
"�8�&M�D�~�DAw�k���M3����(��N�o���M����*������*�@�s�~�2�6�,E��<u~b��bGc�#�LJv����U�!�XR@���x����R�$ퟅ��Q4��h��g�ڄ�(�WD$��M���q��/��D��V���eb�R�̯��b�Ue|4+�Լ>p���1����A)O o<[�u���i�}n�)�äͱ|��t��(�qC6(\|w1�B��M�6���O���	+�U(%�E��������SBEsO^,JY蓩X��}XpX[B��6*3�	K?��l4����'�cr��bK
▪�2�Mfh3�	� ơ�~�)rg������jyM�j����@�ϻ��┣2��!��L#l��菰�d~�{F]��ǩ^EQ�$-x��Bk$uZ�tj]s�ɪ�M��C|��X��S$���ʪ"����4�Q{�����O-�B�G,����*�w-�f�6f�?�Q�j�"dͱ6�/ܾ�$�X+��N؅��}?�v���*��r6�xK��KX�A�u��`������ԀB�b<�O�FIIU֗�T�-���a��A7�?g���\1+]b�(�:��wLt��$������V��RO�B�����Hb�eW|EǥIaG
�Zep���zх]�փ�:x���VV�}1�m�`@�����'�4�*d87C�[��M0X�ʙ��c ���b�A�t�y�	��l�侷��a�jΒ{vV`��dl�z�K$ZW��N��_����K��%�ɩW��:�_&�&~C�}Y'�@��m��b���nU�Ձ��Fg:�� `M��i�����}�3���`k.0���2�]�!Q��?���%�4�����ځN��?On@���,��PH��}��R(�IЗ��7����e��2l�Q��#i-N_��H�b�Q�h]�T���k���1&r"�[a���`ݴ-5��ِ]
צ�p�x�ӟQ;�3�<�I3�d�t�2`1�VF�aL�%�X�3�ۤ�S��]���u3��(b-��Q��2��^�u��q������q�'��i쿖����[�AA)���p73��`�T�gE�1�Qg��B �]��o	*�Q�,v�G�&]�A�M�"�|ǉV��%�[����Q��`/i`9�v�=�_B��ʍ���I�7��m���#��]ץ��n�Hp��%���ї�+�ъ.VĶ�B�h��\��ɒ?Ͳ���w�_��B(�������z�G2n��My��	�dD_����}ϴv�6A���O�b�muʒ�~)
��P�1uF���[���h�Ty��s�y�x����:6o��?[�ur�}���K�x��5o�g0Ͼ	Ճ�Gƅ�n�h��U�D�P���F����i�"��$�������Ҏ�H4��[����Is�r�k>�Qd�!�d�l:�o���<�<_��)U�o��r�����Jk4Xraci�?a��l���{g��Ԝo��U9���n���u8ؐ!��.纱 ��a��@S�xaJW{`�x�vnCm]���5+��d�+�Y#&P\4�˶�Ъl������Wm5f�����= -�F��I��1�*^R�C2^��� �aރ�r�n�������o��+��Ý�1Y(O���WF)ޅ��]	�����L�+���7�U�?�VKbzc�:��u=�����cR���䜻����F�B�d�� ڃ���2k�TT<{LE��:��t3R�&j],tqs꘼ժ%���3onH\��帽i�OwP�	��ŎV�N"�)�˕|��Ժ��M���s�����ށ�_���~`�J r�\��..���b�I��6����7	U�d���V�x8��������*�� )�7p�Y��
ڭ�h�˨�?�>gj�,Kcg���1����O�D`��PaI���3�kT��Pu�+fw��\\G���@7�LY�.�-T#*e�P�$�RS�DN��T�^[օ���^��ѰWqG����,Uas5Eq���+Hm�e�>bj����F~��yZ�>D� ~��G��^��bh�b�-��h��]��s�Mه17��	�+�������n�"��T��%�4��$�]�!hG5t�l֘f�`ƍY�V�J�h�'�u��yL���x��c�k��F��e>3')�A�WFH��a�A���}�Եj�q�����C�Ns���)AN<�4��ߐt�2!�w�W^�Բ���kP�4�k(�B(���cϜnŸA�a��`����1N�l� #0�tS~���=f�b�_��see�C>L�j��|�jx^����\�u�:��K|F]���V6�ʧ��H��E���sUjbz	���W��e�n��,C��H6`՟T��@^S�Yϛ��殲�|���dhFD����ָ�W����)�����е�c�o��{ř`���4�����&!�����S7���0��iJ�<�@=���X�p�&���[�O �->�Q�`L�Rֹ�W<�{��3h�1x�	eV�;�8yo���c ����|$x��Go�KfWݰܴ��������(x�K��ق%�F�JV��*�,�q���ro�[��-T���?��z�V�;�E�t�`�
I�l�K��#�*z�'�+�V|��uyẽW�ѴD��u�xЛŵV�3�>ƭ��-/���9>�|2"�G)�A��!�v�/F?�թi��\ep�qEU��qx>@���0"=Ytn�>��n�_�Xoگ_ƺx᫧��%z̈}��{�$髭���e�������8Қ܂��1�Ƌ���)[F59��k��9bb�u�`�◫�6�+:4���A�b�>*��Q�Ӹ������C�S�ns�be�öXݼ�/dv�,'�C�G�kx���Y���q+Ӫ���k?G��e��;�1H���t�����q�$Pēֵj㝢�\���ifzТ5C(�x�"J�ي�\�p�\$�,�B��X��'ز��������im�/-(q�Xs���ؔA-F���v�t;޾�tvuhb�����[� ���.U�ү�괂5��s#҄���M�59MB�r�ki�aR[W���:��6*���p	U2���n��xjI�J�Q��Z�����9�D?��o�u���=��Ps�����6�1.�|8W���N�}h�Y'>��~���
t� �_��/7I��X�+h.(ո�p��t��"��%CL��O�}��Dbr�k�:���ı��oȺ����`��J�C��k�ú���~���ځ����r�pN�?P�f���q/�a�J�GK#����h��3�,y�R��Z�AE�[n7�����y����56s ����Z9-G��-�<�z5R�����y+���*�U��I�v�ՍyK��BY*#��z�=��~���� z8n�� R�e�cg4:�_r��wj
� ��j�aA,�	�p&g��niF����Jl�)@�	R��3�m��j����_b�&	r0�x�+.t	��\��虎/�@u_B#�{��ވ�@���%Û�m�����
�9�����uI�yYN��!O"Kk1S.���� �-s=��I�8X�-K���Y��MTq�\��'�^������J����xj��@�(h!��E2������!nJ�m�����vZ׃�\sFɩ&I-	=~>bOf�����tWA#�0��%�D@�Uv�'v��5,pcf/�W�./'$eu����/�D��
�U���of���%f+m�w݌'�B/	�.��p%Ja.���~-�=+|���%OZ�j���h�+F\���'���8���h3��#��)E5H`2��!����-���4bf�qV��$�<b,j�vDj��#��,�7)I��r�#�R���ÁȤ��cM�����T��i���<���ˠ�^f�v��9 ��~�e�{a������+���f��k��j�A���Q��1�_��tZ�0cK�:W.f��C&S���3hV9��H�?��! �.�$�p[����^�˯Z%�+84�� Ed�XF|I��G���5��G��k#(����#�.� eLO�Ce�z&�(��0�'9��!.�/U놈��"}�/��A�%Adm�d7�N�D��}��,�xo��
=7H(�d���xʅZ�3$���J�Ny���ƐJ1���ϣ�j�o�)�ɯ�\jc��̘`;�H\���g�����ܶoV����v�3�:�J��3��*2sS?a�UFU�g�Wąg���U���cp�=�/{�P$�~KU������~��N��3��\W�w2�3���bu��u�&$-S��c޶G�m����Sh!4��N[����h�\w�K�?�:�����qS�&��R�?��;.��K�WZ$�-`&
sNM������4�uK�}�l�`�Fc�ӌ4Z���Lg�i�m�0�M�O�@;��&�k���%$N1���f��a܈�v1�5�BF�r�y��躨u��`�Y�K�f��3:�*k�=�*A5�&��Ut�%���=3	���J�>JVW H~д�IGuS��⻴���A,�7���Z������	��q�Z��Y�/��IW�"t�3u>Un�͊�蘄��-���>+~�i�q����DM݇a`�m	����u��Wo��NBV�f1W 1�Ȟ_5U�SGj��z[�bk����,�@F�3��{���C!w�G��H����o�����F&�j�q�!kTY��w�����c{�O��I�z�3=t��(D��%g'��WI5�1�V;��3��t�{8���+�����ҋ�K蔩`2�>��֍��_�.ʽ/x�9Pe�$r)T�������l"���(���R	^}�v�X�����Tb�G��r��j��� �ի~ɅL���6�R?�X��]NV����3�[���g9����j�������d��������C�m�Gc
$<�W��mF\��?�d�6���0�:��[�R��f*�Ɲ�$e*@9@��E,�iU���Yba���9�%+}�J��	���Gkʍ#W���R��h��ax*�	ʙg������&��島xq��_˦�T���d�f�q������nb/y��!ȥ>��
�L���_<����!��۸����+g���lr�. �����f��*QQ�����U��p���<��iD�9m��qY����<5>����YSQ���#U>���t������ ً��I���1{�x�V�"N�H/3<h���ԲU����o+��8~���N��b���%^�N�,���15�|�L�)qn�� �L�c�6EaŐ.�>�&N���z�&u�&�-�۪����:�N����ЉE�2x�)u)N��0�����~4���i�dS�ӈ供%�Z|iXV�.G$�|Rl�u��,>�+�K�Zp5�2.e�bE.�r���k���Y>����sM�V��$ \�b����?!���[��"�Sg?j4����Q]��vIs��Gj�C�BO;Q�j��HE����^�-{K�S�;�$��P���`Ȣ�7b}*�I1���FUY[6MJ���#��u	�&$A_aDpJ�q��3pZF��3^�s>m�G�p�C��a��U6p��5�</�rk��%��y�uq^,�*��#�M<
{�I��g��>4�O�W�.�&^V�Q;�EwYE�!
,�+u�e_�j�K<da9 �[�u�9gmIR�����E�������]ڨK
 7Q��eN�t���=
?1���'��Lv�M�J�<Kp,X6�xq�����yL��qO����sw�$�ݠ���\���^?�~@(��"����/a������dkd��P`���R�A
S���xfh�.N��8ˏ�&�k��{�p���;�?�ٛ�CKV��cDY~&��X�6x.�]������q~B%J�}�y�%ڍ�`0n��'Y���E?�X��ҕo�Lj��B���>�D�̱;�]�k@f��ߧ�5����$<4,���g�`�KHk��Tf���+�-47Y��H�gq.�L�&���@�:EQ	ܜQ��=B�MF5�F�
R��4%�7Daj���t���R�&8V��_	�'����u�q{B����_��r�!��p0�M>�� ț�ٿ���F��b0��JΧ�{���eO��֪7H~t˔�H6��[��;�[z��R?�Y�.���A�$рI g��ڍ�w�K�Z��\/d��n�W"��m:"c<n*`��%��[��w�*� 
��
	��?_>����Y�']��H�7����iRa8���{t�y?�Ct�)�'h��V����u��6��� j��v����)��������@�J?���F���� 	B��Y:�,?�e�x��A���¢
$`�g���{�PI/#�a���(SH} � �|,S�C�9r`j�^�X���5~�H�*���p���]e{vd2�̮["���y�E���`J�BC�:+K6�@
u
���K���{K�Q5#�f�`���^~T&�i0��:��vꈚ�Χf�����m�(���xη1;')cD�=�rФFݩٯ�%�p�|Q�d�M�K×x�h�O�b���� ��/��6Ƣ���V
�<�����9��iQWQ��Zq����=oJ�Ne��?@�p
�m��v^�'i��
�����-X��!GO~��c�(^J����B�`l��9Z�5�'��ٿCL3�,f8o�?��W��$�g���>��cUIXw Wp-�Z7'(w��$9��H���ĬZ'@:��u=�,�wM���k������昹�k�!F��S����|�|yn�j�43��&�K����bIW���c�w�s������f7���޴|Op�@�w�0�F7Q�ZTҐ���U�.#104W��P�R7��.I�7ܣ����#�/L���,륾�0CT����P��j}���^�]6ت�mEN�nTe��J�nV2���#a�P��@k�-�'|����w�t�[U�M�\�L16��9�Vb��(o��- ��Q�����j}G��
֒4�F� �UW��[ZD+G�$�[�i�9xl���v����	��$��rB%4��֥w��4&'�:V�)�/����.\JN�����M�xvk8��7L!���?�|��7͑���K��=�,�o���{)���n���x�W��G�_X� �����Q.xq�d�����N"�ֵC��8��gr��B��_Ӹi��7�����p�mX@P������h�P��/�/FI?���O��k�g���~�����)�f���f�W70�Gr�WT�<2����b�����R�qofG~����ۈ�)_��P��F�V�L�m,�D� OLw/���Ib�s�&
��=���q�r��T/�_�O@�ᖉ�����"G:�)���O�	�s&8�xŃ�%��%����4�w�IﻑY>�7�{f������l��	��L�p��ۉ�w]�jw�O�(��:�>o�r�Ec�ԏ3g�<m�Y2��#b*nr��	MkK��g����jMn}���J��w�rF���R��\ˌ3T%SP-�B���ְx��D Ѡy���3�0�`���6�4��C����;' +g�T��Tԍ1;�p�G6�e�#N��Ju��{��"��i�=	1����ذ@b�*��oxƥӷ�v�r*i:R+Ĭو�V����
űK��)�Q��
�	q�-{�h�-��Du?m[,`��0f�����V]6͖�p�|�J�}��L���C��^�#Njs��q���V����*-���Uh�Q ����KOr��L�m�W�\�]g��CP�w�+!3���e��P�0)�,�5()o������RN<�ݻ�D.T�C�\�&��z[|Vp�j�������Ai��i8���+Ea641����ݟ~�G5������ڕk���Wh�{����/�����������罍2��YP��)����� /�g$ךҎ�q�tǏ��3���_Ţ�Zl��8K��:���t�>&V��}�1���
߷+`_HY7�Q�,:=]0R� +/����(F�c�ǔ�� o�e��T��so�iG�oX��+P��d0݈a�씉��9A_�x-5�z*P�՟K����D�q���G �x��%�E�i�],�ib9aD�����ЖM�