-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
flPORkp04bcy/ShyTI3nqw3I7ZKhEqyAANL0hdQdFwRtMPdImEb0jkpaXIGw3AshG4Yt02Ea8CjI
Mpcx22Ekyy4yKbI+yIL7/4bhDwEP5gyuIwEINhbMqmwwpcw3zqaKNPfRhlKRZIlEMxoWSE/hkGVy
F500gWRIJ3rulfecxe5BixGCSSOrSdeC0iQReUfUYZQNChSMQlC885VLEamWNodU4qzqmCTZ7Zsx
aGjsaZ5tq/ddVvjDZ8v37njm5M2fGVR0NdEyCI/QFwJDfms+vZRN9EcoRgNkisjimCw/IJUcy+eC
1q90CdQDdV8qtgZeA56a0Kht6BruK69nv5viPA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
fkzL6wLjHYMtl2Pe2YggO6TDTQp5x4PZXIVc98gPO7t452nfcoEXVZ/cpgFOURVs2XzTXgQdKOpF
9kaj80P23V0g40RPRqRickdUB2nwmPv1ZTroPtKhJAJjoEYDOeSRD38VZuoe1OrWqJ9gMVoL1RQ5
J9GvedtOqi23gAzWvhEY/gGEuUm5DhXaLeLiD5rpdFBt0FI7ZEH37Den2/zoKzv9BGtiB57MPsA0
tJxbJiZuFnJwnf5E26FVlWC5+QBc4d6MQcDPDoZHLarum/sQsb4N2UvnNNLnej8+6/qHQ26Ntbpc
GdsYXOTaFQUulOrKq6cCJCTYIVjX0gQkSgMpqvLMuflSbiymcpkJg7XQREO/ULxF8U4sVV7hSORK
4E2Rq34Amd0pBTLQpffr4bIIlVlpbFx37KzGLz1+gBLRuje9B2KSJFZR+u4SiTL6r/76h9RkD6xU
JDhpb6W4jl+rKNF+300dirPZxGMfrM2qAPzxJlmiFaSFsEfR7ODG9bD6PZw9N0p/lbFPEZArxTpS
FoxO1nWXkvtfRorISIeZGTWxNjamkb3BSU5kTu2Hg+RPelTW46+YscyI2Ht0+nsrvgJQ6bs+UICG
6Xm8cIX37WAoG3Yb4OF2s+F994WPpDyh0zMWjV7rpqPoAthvX49g/2/KshpG5BYOSnWOuEpXI9Gf
NJGO5a2Gq/AIx/oMfX5RAOas3TGSWGS0skC5WjtKGnKkOQkHgLCTM+46xvC6lMQvgVgdm4hNrdWG
f6YAV7TyF+BX9I1Ygjp/3qGHdwtFzt9x+lj1ZFo6xWdcfdWCvlvGvqdNyL1KkYMYdnhzOMKjQUT2
qKbfZGo/WGmcGI4bEoky4V3j1w329GuFoZUY1ZZviDJ1/nkP9GndD+MP5cAERAUWRJjUpOXQfDTA
w49xVtcF3bQfeqqNcZ9ed/eN0mdwVYKTX2j0gFuWc7sEM/8Pw1NRE+ELXkoZH00RLsnWa4Via+nh
fLcAvbbeyYuNCA5vAeTLKxU3zGFwULIrwnbR0I1Wu7TUnib29GNkZYevrNXlwfjjvVI0Kf3SoMi/
t3Wz8+ha2mZwQkjPsunZE9UFNwCqKU7/ezXYmaYtuXpMJsSjqdTRVgVmglj9k6QEElYRkyG166JQ
k/MiJCN9CsbdKKN3bdtks84oVSoRSnlHx92B+LFLYireRKVS4r4h1s/0F+lSnMudPjLHaT/k0Veh
DDQ++JVJlhoN6ILL4Fp1HtT0Y5+5vZyTtGUN1SZs6cuV251lUHxrMXKb58+ovw6Q+LS3Jb3mB/Wh
ZkQXm7FWBRKVnDUPkUqmts4ul3GwKhUHO8EYkcwUOondF0lqKaQih5suDd31NUPK3w1b28M0+RPj
km/bh7fTIOg/YeQYsGIj5RLWu4rmLYyIOWdomr5pPMDpcw3S5JLuArwQCkMYuEb0phdjYciYUdWz
B5LKj5d21vQEOH1B6hAliWgVMqOnS5DXbscU1Viyefo4DFXYai1sNtI5nHzFfb6e14QkIeGd3oyT
e+kHW1vj75taQmNqBhqsdncqpbqmVduqai/VW2Pr2/Fkw5nVVW/c1bkEt0EOlgCDsvxM+RbX/OzT
rlFt92MAa9NcmFKS9AGbVU1TY39AxQZaz4N/bvxGqS01eHTORL8GTIfBfvKMTiIwCBZBtcz/ri8+
+AaxtaufC9vbp7PQkejVfR/MOuIj9iZ7wPvZYJXQwNJXPaeFZVix95AXuGLqEpLnh4ah46H1ePpf
Ahdj5aFz0dY5MrIei0Oqwr1FKOvQXpLmVl99GIFr8facFBrz6x+6ZVyhnkO1O7bg3enKKir53NpP
0cKjg8Sox/rOQAH/zVCqR2Amzt4IxK9Nyl8L66OtB90Ebh6A0BLCqjVldMmd0xnHKdM70xBG89pi
8wNKyhCuwIrHiAkkKp5lq/t+O7bl0Yu4NAz/rTgW4KhM/upZ3PG0S0UKUPtwhnrheRO0hoduMJZU
5eFc48P9tkQYtbdERzLiEqu2L+rP+5It+f61bIeWPGGL5/0sNXhD6gROYSIO0jWhkEf67Co6k/WX
EUO38dNmxvcLpxnRQDZ8BIRGAz3bbT76AD05F15TugTJsqXYrgKl6aXX4W2dRZJQItOPFtHxfaeQ
kjillSi6MgkkFmunLI1Hl6vXrX7sbrBzmtnwDLXx2291Q3KGWTg73pr1gRvAg21j0PZZLIG4inP4
AEe62ZcmavgNiMVV+CRqGk+nAqSaewgVA5xRXksQGisLYaqas5xfws4CD9dgkYOaAx887woOL1fc
wvM0fGAju7g6/voKcaNFtk8oF7EReB7DIdkWXgic/tyrRVwQEDxJVfLntfrK63kVlsNH0rdRgAY8
x9stMWwG0zAfK2eF4NeNPfNKxI0YetYn+lpXfqmiW1q21P9SZajq/i6tfeMgie4XuxJxN3dpHyEE
36F/bZijwLWHcyICvlT1uowJGiHK3bO7cW/niP7XFiJqhYyV3z6VU2ZY/wpl/Xk+RJKB7a2pisnQ
DSFZzfLc/4uD4OPwoopPbrJdQeuOiv2xPFqdOeE4ao6CeWifMS5Q2BF29/v9PWWd+P33hLwzkyyR
PEwL91i+xqqfuSnsAexHq+Pr2zC7cREDp9CMaY9pL1y+sTOps0IwYz7NqBXCK+r6Nln1VDpzwPxd
ymOH4Fd5MVCAoGV45gxbFA/Kp6wMo+sX+Rp3Td5S8SIQnXoZwozIg2d+WomEbBIIrEix7CGAlxaO
lH3NBvlFthyf1lOcYuiQEKMoAMXB5zy7GhQ7GJpefNkjxoI8Z165J7qBT+iUAWfgtd/4DMXYRswo
u/EvMz8OjXtT/pr69VPrMvLuli56Pyc7bvlhyAKCQeGj6FUrlGVDUCMVpTUej37sGDMkz1tjkVBn
MR1PToABes3dirCrnypRp5s/kyqtWCwuqTgxwIYXSebo0ut0epHNpgLB18WqmElPMRUAQa6A67IY
J53e3rdrII+PlKG/vowMJitFB8eHwj/eyeYKh4whXXeGFFx1dTedtKGF39SjJ10JGFX4LwPEUeRA
uHXQMw19PCud6jByGGoaIwzXa7D4mkPUkoLgO3bE1wq+j5w1fRFa2PEiqLKXOb3cAXdptw+caflT
Mlj0Ky84d/F/YerSHAj/TvtxHsk0plqbMsyKmkqLoDc9EIzkZhec+rajkK2G7qr7RlFRMsw/jMKf
ZmBaRx49OLUhM3Av2LoHVNpwvfVY+iZOX8N0DVAQAew6SYXcRVXa8ne+//763f93ydqKHjrimJGk
8/ALh87RiHAjBnr/Es3fN3Gewkxm3A+eJzpQK7NlG6xhvsMq4Gjtu+CDog9xltLSqTJoVJkVwcwo
7L3iq54JISrHhkzOxnzgXTGQF6rcNEgKGEuAR1j5b3LGgNczkWxoUIXh55g0w+t5/p+VK9xtVUeT
r6L/Iq55uIcpNIDIqMUJPFbNn0A7bpNVW0lRkzrSdTxr1z5NuqrFzII3d3RkwHAF7rlbQ3Lnv+Bh
cle1z8pxTO5N2S4LsfdAiQjDZiy75XLGG+V9otXv7pVuNvym5TtJbSvbgecuKpe5oU9SXCmbxaP8
QZvepM6Q79Me1sCuADl/5xsbhX2+UA3KakBzKDDG83r5a9Rw4IzJVmWxfZGimWPskrWJYARa4hEi
s/BRoJitjSOw8AK16y0Mj7gsAl9ZhM6gxjMO2cC5VBetYWOfx+FFJbZ4u5P4Lx7uPKJ/3sgSrEea
r6KqOXNMpB+O+RgZUyQeva+F3Bzl27FNIqNl7UzRkHbPX5rv1EjGwrXfhfQvRFeEyMXGhrbU0zpS
FpkeoX95qlrQtx/7w/Ew7b0edsmFdD9lmA7jhlHsdri+wbGkDRkzHk039t/q6HSekx6fYMbTsKBH
GM88EggMNvXfBDfwlM63Nr55a2F5r8fSQZF3LLGDzd4J7wS/VUfUK8E/i2Aw4zT4JjxLP8Mc+9Z8
LflK+xPSWqLwJv5YXDQwduyvTTKJr9SNfiZAmG90Ehl+FKuGrQbslCFR4tQyA1qdnlA5yv3ksOPd
6ajU01A0naCpDfNX26JuTmglYQjArvzBYCYPQWyL5es4YgWxYwU81yvi1Qi+JbI0yj/Ohq/TYIoY
zTn9ZxNMejXghzZVX8c4c+wwTrXZV0Yzybvcye1PnVbgnw4ZJt4KHuhCg948/z80+7HHW8zad/ms
FGLCHNuBVPEbVsFbEoGQasDE/f1CJYEON/8y6XH92mrxmWTRCSTni2JPCUsgu+MUQBtAyrjUMrT2
r7/Rr0ymxzrp52cC/5a3tO1X1uG7ETcqq9qLPewKTMqVUJ5UcO/a7AiZfcn7MOREr0PCr7ZM3J4l
oVOmvUUcRpUZG0dQoTbgeDeY73dSNENCJ+jDp5Er/wAij9xsm/goZYkWWaM+aVKUadPxKEQ/Wcg6
IKMj8iasqvaXWMiUT4ieKq3Yu0siLi7a+VkA1pANjL1VaxFh6Moq+xUyJ63foAJZdB0CGQp43THH
ApcCrzz5bpn0jnC55zwihe2iufnwGR0MhCAYQkkORsmbv3YMNIvaRPfbz6Cr0D+vLH7u576G4gSL
Pm144QJM2wKworm055Tdb45Je2kWX/0u/9GFvVgLdxzEb1koXIDJe+I4cNsjXqchXuR0hLtVCF+/
a7QTqkv2HzHsMKr8IAOmN32r7ebcUwnUYerdTJeCLhpgNFbCqm0In6AYxLPdFI32t6L455f85EDJ
vvpHK0NGjceR5Y4uW9KZvFVLk7abfpMr4VogTefEQfwrRemXNJrgZ4h8GHmFxmCwstaWvJ8lynS2
QMdCCNRmw2smKQjoFxJb+58DsaxgK7kHbf4WOYtK9vXbew0OBRNKTdlW0/G+KtIM4a40Gy56m+mO
qmk3AZndgZKb/lHgu7/W+fECx0tNIovPqPSOZICeg5uzXDbeAZMXVDnSy61RVTWttk7fawEfVCRF
VzbosFNitgGFbb/rlponjk0Bcw/6sOxEKMPqx8KYvGH1alwOH21pjMnxEC76fI/IOX9RDKDOp4pK
OUWrjQO3AESug8U6CHpqgDmodgXXOAWuZ5L/qLYNNzedZ2vOQBcADVnBtPsAl319rpfq/T+cjLma
0ivnBVwTSzzJuc8dj1vFIdfFezXJGBwtq+TiJsphPJY3hgTMikDn16b5lKaS9D7obDi6Q6G1v3V2
yjK1J27qshc1+b6PY0lLJVM2TM6xcS9nidD5YntrGWKZ9BdRBsqczWxPa+gOZJopZaH5NnMFUFqC
5qe7hnYyxbZOLSRIN19OWTqUlcPJ9ZwGPoyesw83j9lO4cOcEHjGjQkzdUvKRg3L6FqEiTZCBbFE
X2TQJ/B7ZjTe8aNAFABAYOZfuPFV7n8WUpomVXu9xDOi+c5BYl2g44IygnwjObomSdt9gNPactv3
tnK+ZwN9ewYepqNZFWMjSseB+cJe4fGie7CYcpW4IBbtZxKStsSWy4CzVRSPKTQUtSrifw7cJ05/
mRshOHdfDF4XpnYkdmRE5xHCS9GqxvatJcsypRxYESJWsTotsD2ugRT2vqrQQ4gFcHJWJ7oSD4Sm
T099IddqDTDvbB47heFQnPhtASLtVmvcm/ngz/PY6dglGmD80dU7I97DB7Qi7dBnWN4pxpB3eOE7
z9Gju5Ju2yl0H2/ZRFBwv28aQLSyZanTPu/dZwgu+PpZoSxOHyl3BvLGX9CdOoBsTn1V6IVrBf7h
aRfXQ/E2t6CgO0hINZg0nT3C50oIN6wZTV5c4GlndlzMOBhnk3cFaymoChvktS7zGQClg0nfq1m7
qvvsPNKhB/s5QxqbAXa2tFSn8dBnIoMdbGeamGoBNPjBQnPcjwjQWPiZWE6kse5Ai+y8Val1fR6b
5CplZMDw7Dnk3ZlpvSIikeyPP8C5d/d+6X+Gc3Xo+4FfcrwDPY/IJu1XIRwlJ1i9/BPl3UZb44ya
n/z9Qx5qh2w6TePyxtxSfhBlEYwgUeSbOmo1lNzPzHxmobvEX26f4hQk77L98Ul1SP+O2GilRtHY
OwfOvAdsnDH3h/DdcbHj0IzCMwCQS+B8OHCodlcD+3+DIZRBbr2BiI4Uhgy2haKeOusFZG4cspsW
1N2Z6rSh5tcvmSPFfu9PZhNmcdM7BirRfi5CVTQdp8pl6QzzBR0R9pCMMnUsR1Vm32FUUd/h2Lkn
G1Sn5vsfrE14WkN0XKA3YeZ1EawiQLhIJuhPPWWPUh16UFKNpNrkmd42JwcrfigEzvyqKw3Ay7+m
/jeEUrhIbQFfUI+qOpUZ5grutA2KjY9ta38q3Hgj33FtCVUdEurkOt7M+WVx7LGE7mGsavliy2HL
dNokTgdzNKNvX/diTUa+pQm89m0t5wL932XZyoeX/w0Kn4+F5gow31Y6FZscZW3zO3YMn9YCYwlB
usSNSCi8nKSpRwiELUvPZbfh6thWM/x91OI5EZWDEtEXBXGVW2Yz2ulAKHi8AAtyTzoLMYm9ha3s
9eiTTe1+6GcAXY/fifv5kUb4/6s3XGZyNMU5qFO32X/iWX+70Vh4T6EDOf53jJnISjjDSAYD16fZ
821k03NvAu0osW96xA3jvNaLNJ5Sj2saSom2fyMovpXaSNe+fBhJI0pOovwV5tXpvdNQmn5mKkD7
7Q2aYMd0EtOBmCpt/FSld6gPsVtJj2F5gBlSpGILYFLufFqhDLII77rQPAeV+AC0X2Zi/12Bx2Ba
tkfg4AZwOFDB8NMTvuGM+ODMItIGOjYHp9uOVNnLp5yg01l6rYTMd2KhVe59cVwsVkUpDkC2tbfY
OMyjXnyZoZdlyLTZUCXrmmbQpzBrWZv28verjrfEzJQ40iZgj1N3wh6W+XNZWxUJmwr2P7Ru8kfK
u4VpBlpiEHVROzaLdrPN04NEYAo+7qqf1CGrrL2FPbE+VhcVolw5fxcpvq/RoAAOXc9dKVJopG2W
z/CgTsH6tmUW0AQ6VMbT3XwQCa3PMHW369mjHOWFpRwOs85VRfblyt3Ly6SSwlRBmLKnotD3Q+tp
1Bt8I6ApSxvY71TM0d9zSKZM6RSySD3x5zxToOUGT8jMy2A0/sP920AwT7QTda9FSZHDaK+N7BKX
snboqKHcy9Yfk7OMtT9E2rX4FS64xFX8zjWTzphB6DCU393hRUr9YUgY+KuFHpQ5hwRUr3xeW6c/
+0q7ykI0zhL6HqQTfuMPimtyRszX6bDybshtj/hqtwI0UxSU1Vxx5BkKhQULkwZGw4LW0bFkaKsm
11n1WxTqE4+C3L4uMcQJUrTFwMDlwRVV4cuabAj8OekZ55ELpoi+B9bFKbHEAuvXAcgQ4/u/jxLE
vq8qT6RpIxDp5Rp8svrFfOn/VtmJbfv9HZ+Kya7YsGBVA8d8s7FYBtrfkJBVbaJNp3lXxo7sa9zV
zWsUefNeeq/REKOuxuTLQ7zecAB4NEl9M9m2NSPo+qhAe7VdZ8AXWSU5MCcE7LzPhI6MV8nfr+zp
59lYhaPTd0tDCOcKxllG0rZZuk+4wutKh47Okzn1s7pgWsTulC/oHZhwalZYDx+VXm2V1gv/nXUK
yQCyy4378liTFtj/qTXVSJKE7F/yCQTYMZ2loxVf+to4fid1sI+eMKyhHdc9l+YrbpjqTu8iYCH/
Wa9hln9WICUD6u6x1+vQf4+EaiXZHmoxtwa0I/QDrzNRxrdKMv1HYszrRyw7fpsc7LndQKWD4+Bn
FHDTqBmUaKL3avpYB7NhNVoVE9WmpFjBHA4r9YirRs73kDKSb6Hhg0FFEhgnmoswoE7qBihL2nhz
sT09kIvRZt/cU8xHGdXsrRtuZSsBlePRZVskD3KoQjsXfOKybRlZ+ILPqk9d6aoKwW8E+hMDdc6U
xuglPdng5elNHOR6ZT8mY2IGCneTnQituU89gDDkCA+UA9zbcDusAHnDFUrVYGNiLxDt5LGwn3WM
oPMS6cqsnotE27RrXO+GPyT8u2/BA6cA+ECHQhOyEeIZgE4d6lrWqd32oK2x+9wh4/rKaIGRqoZ9
B9fLOlaGe/MXneL88t7gzGew9xhZCYaFvlWih65J2nnQg6Ynn2iL61qPocRS5SXGhUJodAPuWagF
gQp0ER1GefIRy6Pk2aBlvXUJbD72d9c8xWP9X/3+6gjoY9xlM3NxP8ff6vG1jiOSZKISETej0gzH
qkckUjJCMSYfMI0jIO9/k5bE8rZ2GeEEXZmQ1TGC2zj7sycMHRL/RfzW0wyct/GEGCmF6/S6TC8G
cnnP98gHcxHqtyjSXGHLk39bIEAJLTKKUNjANyLTFSQa6ps6VuNOtQtUr5KEZH4rAy5jI9S0NKQM
ZDtfYObaK5NaQo0yX28o292T71cpKKUnJSquSc6gkNwTCHfqfSJbnOIKTJMA5ChaAxa96MGls67b
F8QmXe41Blm68LU9g0UyIvJiCNtWDthEaFStDAf9TyDJ4QUsWks3aTFFduLI3jIQH6fo4+49CZSx
kY4v4YS4dISMnNJzYsX07oa8LC5Z+yD0bET1jhoApWmM8EgZPE/XMkaNBKEPSbPufEWt9yI3f5+f
2BLmiul5anvS5nmlKhHPWuneLBvI5PS1Kpr4nzNVh293uNwhTXXIUPvgBsCNlL8lhrWhZhtpCsbS
Vy9noo7WTrPBzY2+D965uXzUFrgCbBYAmGHmyNUHZNuct01bwqzVb2XhhKJCAXi/kHzbDiH10TKy
yCyaGJf+l/Cig70kjnhgGrlf/yjGtUvZhBaRQJmUPkaJii6yeOf+KiTe4tpapZB7CX22657bHdE3
lHg+UIXuFf5kSyoEIEOrj35nPwbH3VIF2Xyt2Lvo41yee8O8jR4WrVhuo+0FCW2cnQERkrxa22ko
h21LbJYYIgCN4SedQtSL1C5DdnEsWlfBiB3miqDCLYWId2bFDYOYdtgafSqz+5W0DW6N2hBbsumN
87xnlyP9qWtVFZqUgQdnjHlVwUfgxyq4j5GmLr7Xufg9INzCyr+OxU7bsRSGdwxdePRsiOjWTSJ+
9qVBpjOuEw+KSqpRSmSlecfaohLw3bHxz73z43zGLhjN7V9nvOcJocW5SgThEW+QfpbxJpjTnWdn
0bIhio0nSdrAq6wQ7lY8lY65uIEBygMxFr8j83e/UbMc2NEiuQ2gMCZGctS8FRjSi0SDNu4h3ytF
IZpzmqMLdqysKlzZ4tv4uCspP4GXBWKtfwCgybPOxBg2AtgYpEafwUlMKEypMnrVmiPOLCLyp7TY
6FIiHAgwORuEFg8JEillQYOFEOK2ruAAskSXEbzv69fuoLtgc/XWJT5zQuJLf7Eds0xlsjywwGzY
DPF4nGPlhzrVVUPt5UaI3o5K4MDi9paqlWlZaepXzOUKqlvuL3sQLLZKq0kpYobW/pSjKVbL4kSx
aP9ADDvJWNIwdlkcOQCsnPBGiqROR39agAbst0WDAo3sxU1uEzKRWc69d8i6FAAF+jfXJm6V6+6N
umcCRys1thsifgDlMHjE7sKAPzGlyAYYKsV5r3vBnUYeH5zC6uswQPQ/Ibr2SAu189YFcIeFWjOz
vEbQM46Taz1sn1pgPdU7bGLSTO0oO4PXRLo1u+bs9jCRfjP38JwUNWt3zFkGRvZNKnLLnhbDjOEW
wgHSlpvh7AvDkaGoTDrTT+98YeWMyW86jVWH7eKIiEKz3yvUKbwhQlg+l4NkXtiM0g/8O//g1o6+
USG2qH8ngHP/s57bIodZXZxiQtbmboKjDHEFeykUHItTqaVJZqrXEySRPGvvkRFBmy2oPd01qvGw
1y4T3W78Kx5JdyLiR/3wtZ0gaYZPre67LUqGEHava9p5S4eLTBmcaUyuCNSJX2tRpy274zk9z5WC
Dywn18J8r8dcKRQe7IeGdZTDatBi7fH8enQ8bznvX0aPC7thDDFhUgtKKk4nOpMyG5pDGp74pLVN
M5WY7QSr8ut7Usen2pHz3sNzzSU0kl3m49mEjI2efFOnEdlBcIbAJywoYRjWOJuiu3TccmUNf7wb
I8sw3ECs0pE3RjMMlkGLry+llilHyhMdnm+mPfILjmBsEg3HBfMS1ra6xTB57aWUiOAkS17tP/oG
jJukws2CsbXPImU8mY5e/f5ZGW1+FS6YgGZTA9YzmBSgSnhSVJ0x15LXaVCD679YDLRytrC5LNrm
ylJOfFbVoogMNtqvIwWsbr5hHpuJe2XwZrAchVq1/Yh0MUxelBd8vCaut8+3AOZeP17rveULlVkK
qHqJ8bRoD/7lDRJrpbrCeiP+VgtzHwyA/WiROIDDHoFFsnvBWkYiA7vBL7TOpI5YkFI+J3ys+lqp
PR93508qcvfeisc+5XoLrJgsjSIPPMdE109MtjfMuSimfnY1KPmz0HtTp/KKrq99rqckuN1w8yR8
axwyasi5ieBsuqVoOtzngSGN6xga/gt+Jbu8uCG7javTKlGwlppeKVdSB7+u9Xe5mnR9XhkI7GQ2
4BGR/lrHgiprau7vNsa95MZQlyjlisRNOKIHqbuhZj9OwU0a1YnDQ07Pwgaz3CWOO7WWM6zT2tFV
keBzgdOSDfZd0Tw63EhUwjVnVh4uKnUjzuJ6pfeWByxVo4wTwgp/jU2m0L1DjuVRR+t8jcCwe3pP
b7/tCSCgmZvDQIW9W0n6wFTkSAJx4qe4hGHiy3i8coXqIzgPwUxy6LYEVKEjGnF/PyFfZUkqjBLK
gmomLZdgMKU2TYfwtCLjWDBVAAi7tovjrtNH3Zl93Pe4x//AgAlWhQ+adXgKW34tRchSmUtf9jkk
zqOdmz8rCOoHI0JQCaoIYLKIRVwqM/7h5lHsv44Kz4H9usmMnUs8AqdcopTqSibYafwqFLNLNd/l
WOTJ3wYAW8PQJ/InOzddRhYk7KXh9LaqFUYFnHuqC8Q0ELx5vtyxARO7blXDQMYb8yoEO1d+sL/e
brIIdt4k9bWVtD8Z1GgJa8n2giod1BzYFudBIrCz7dabkbV+z/q3dvQINC41zuSV9IjViCbaAl6v
`protect end_protected
