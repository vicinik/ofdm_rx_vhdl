��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�G'?��,���ɎĖ������T���CiC$�
�k�9O��g8���	����A�s���Zs���AL�ҏ��J���}i�د���HB$�%�H�O�)�WȟZ�D/�-�^4"��Z98v�o�,��#y1Oq��bq����+D,�=����Z�⾮A.k����>�����tЊ�U�a����Ci���]�"��+����c=9I� ����ȞP��q�#v����V���mvV��Ty���:FE�e��S�]�$���z����ـ{kb��#��I�PP��D�Ӿ��V���W����2��!�;��-ю��0��P���G�wq*���7�s����H�rM��"I���p�v_\�����5�$q)1�)���[� `"�,�L6��ǒ{��/-)�T�v��� 2n�����<@�?��E V�>7�ζb���s%G�4u1�QKh�C����X�ΰ$8G��7P)Z�����K }��q�Ro���6��������៹y�39�Z|�v���)$� ��e�O�^+F}�5������{�����t�C����qcU=���ے���z}�d�Ji[�6�G&+���-?OC�5g[�?�.|��ᯋ���JmEug�1�#�o�e��`,L�������L�z��\�C�!�=�
Ȓ12�'|Mv�x+Ys$J��R��F�)�z���-$�Ts5��~�`!���^F�]K#�5��N�t�g[c��n�ŷM\ģ [A�t((�8O�o�����P]V�ž����(^B�ؒ.\�N��5���6��銵���Փ�u߬��O��DZ^W�|�~)��cFw���R�Z�!%�n�uB�nķX�\�}�������-��y����1fϨH�]��Xz}��
t�R�{���[�`����Е��Hj����I�p�$�����2'���|�����Cǽr�ϫh� 6�����o����Nc@uY�=כ��1�E�j��j�)����!:U��|���4��Zr]��eFdLl�ÿ5t*�}s��%y�0O�M{#��v`�؛{s3Bn���T��<{,����JS9��v�rO.A���ߧ˸wu�R_�_�de�z!*:�/{��B�0�n��2���@	�f�T�D�M�ϼ6��ʡR������G�أ�t����/�1#[|�3�n�x�;1��F�P|�m ���T ���d��2% �9uj�Qaz����^��$�W����3݆d��y��\�/��"���C���}�㼟��OE1��M<�D�����J&{�5�
L�Rgw��{����ooI��|$�����@"gO��%�,Nx5��Β$�պ�)V�Z4�&]鉖M]��۠7�	+Rd���Z�a3��9.c]�
F���+�9�>c��j������7e�g��C-}�q/Z��	�b�7l#��-�����Ś	���
��)
�V<��յ��&�|�wm��[_�e��s�R՝�������0�BL����s+>6=��C���^�w\�s`�X?ӵK
4on�=ŌX���a�g�WN�i=(m6��(��׆Z�3�#�9v-��u�f;�V�Ç9��Z���s�χ��MAu�bЦ����٥���Դ�h�X<�1i�S�l�`[�ś�����ު�}V�4�ħ����"]�3�1 ]S�����w)����2u���X>�-#�XL��j:l"(����1���c�q�숇k�٧��8@�?�[	 ��1�\3ƪ�'�A�#�F$��il=-��LƄ��پE�9	|"h/Y��+J
��ͬ?�e�t2�T2
����T�VZTP��Uloo��o(Z�
L֬�q���/)��'f
���0�$�%��c��Z�ї��lt��i�ͧ�,�e�2�\��I�Mr����Cfu-f�%�[P���%90�F���ž9�b� 
���>�R�g�E��9���}�X��G#�Mʑ	G���7�p�m���$��aM'b���gH��!KM���������$��G�m�*K9��\^���{��������:8G�93

�1�r�w�Oh�(���9 �M�Y�yJн@��A)�l����Q�i)n�=������RSh���_��$�;��t�ŕ蟧
�$�:�ゎ��pC�x̄h�oݐ��C�e��RXD�RbDՈɭ�B&\C'��P�z��}bX|Us�B�j>���������	�?^ᵓ��FZ��;8$G�"���۝����+H'�we�;�t\1B���n	H��s!�K��u�cu����s(y�	��DV��ď��7��d�侎�jM3�A)�_lY�y#S(c�ı�1�HA���$��+����j������ɓ��&y;2���瞤��6,f���n+�>�B6V��=�p��a���s�3��4�˰f�:|beg;��f"'��S Iܳ�=�1EB4��OAa�"	�2e�C4��m<(�?jg����+쾘���Y@E�� �V"�XX�1�황N�귫��=�zR��� ��f%��5�}?���4Ut2!k��6r�ꘗ?��@����n�UA�D��'R�nP�����1�e�,n0eL�t�92��nR��P�5��C "����T9,.����r!�&��a�c��#
��������Y��fj�t|��K���u5��Г���e���ui��G�?+�.3V�� /z��fey�]'�I��Q1�����N�}n�ཟ�g)�0mkُQ�5A��d�=z�H�wd�I�H�e����ՃS�G+�����L�?�
ÃW���RD:oT��O#1���K8��a��>%U0㪟Ȧ�/�Mf.��Kć;���b��E&ֈQu��Y_�\͗ok�㔘Ӊ��T�>��VlfYGD�Z�_M^!�SZ�9iveD�Mc�L�rO�����:z�gO���.��k"7������el��J���ճ��NF��;ǿ۰]��+(�
�"��k5�uԧ�X\�M�Ǳ;�lmB_�n�
����l�]dZ���\��*?�er�X߫y�?���oeK���F=�'����Ί׃�*o[)�+�2�����<;v�%����#��('Զ�Ue۰0,e��� x~9�un}˛T�����t��}����>�H�E`��I1�4�@MjDV�����q%/�4J�����-��L���2��1���4,�����&z�r�g��&�Ҋ1��=D�����l�[�q]�?�o_״cE��Ae{U��	hO��(�j����
РI�b㵄'�"��Kֽ�$�
"m�d����st�lu�X��Y��)�$�LRM�Ԑ����'�w*awȩ���*��C,%B��>�&~��G����r��#Wc�l���h���;�!��'w<�����l��7�7���+W�*�mu��EǐNg�e�y6�j���Rb�l%�5�Uj�~wfOYO�Fsߑ�Y�YE�Pm�@�e�Ƕ��V�ceN��G;C`���Pp��!���u.{�v/��b��W���2�����x�^��gIA��U�گ��7n�u��O���+13�ǧ0��u��^��`Ub&�}zC4���΍�Ή^2��{;�jP��N��R-}�p�̕?�r�m)F�zM�:�L<{5�P����5F)�Q�W*;?݋
�޶�]�(�t!�pA}�!��o*چ�߁�%�S]d(2�#��8׃�8���V�6�W���"����.?ޔ *�y���W�lk��������Z?�yN��rp�jl{ͬW�˔��sh�Ș�A���M1��3���C{�J#O�I5ZM9*��۠�C�Z6��LsI�`�Y>A��m�*s"pR(��5$�v0��{ ���M|����U|!_�_e4,���+���Е�{ʝ��풡f����I�������zB6��M3pK-�*�b���Ց��ݷ��n�����?D2g��a�pbb�����G�`���\����7G�|�X5�;�Y�=r?��{p�~91��EyG�b4�	QVƩ�)Kw��sВ�e�Y�ClA��`�����L}yu+�6�]��p�A{>î���E!�iɺ��������ʠ%�Xq��ʨ�c�f��*<�&M"�v��g|�u�?��i���j��awK�XM̈2oӛ�&�z���3�Mz� ZJ��������B%� \���.i���닻�dWyqs��q9��g�,)�B���pth��3N��P�x��]��[��~N��I_X��:�P$���5s��H��!�����+�$�sF�#�'o�ܗ�R�(��դ���g�P�������?=;�f6��S�T��I)�^_"wțD�X�ŝM�Uޅup-� G5�g)K�?^�I+(�-���8�><�bC#�������@�n]\��D��RQ�>�v�/H���Fkj�e�ك$)x^9�VWv�U�˭���ߥOI�W��MD���Ӟ>���'��*W{�~���j ut$0ћi[��ډ%�g7^����b�9�F���[ ���}�k��l�Q�*��
�De��^�DRi`�<��aՙ��vz�_/cw���LK�C��@�1⼭nu��v���v��D��L�iDt˒{(�����K܁��8!Μ*6+7�7+5���(�3�a�Ϧ'e�