-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RC1bx+VpyodQFRNj3nhUd90vUd5/qYZpXzulx2RXJZTXHk2ZUz9QjU6DgthgpUmDDeo4AZe5Nsh4
awW84I8669wNLQxVzXxsqQaCNNsMW74jm3SR2e6mk0rcmQGcbKBrjCAwuxUshxkP9khjOcpx2S8r
OgjDscPAXaSuW1mCzRiW7cPtHsn0aQtdQxds4EHFs8HVSqOACe6emsHDs3V2nA5Z9vDz2mmBQaup
50qeLvbBWKZpOStDf4T1TN+GV81RC5yDyOLY9/XMAsWi25AvDmDKENndsva6ThQHA4vfpj1V5JNB
wNpf1QkgoGGQBt6/FATTybKxJ4EnJlXhf6LLvQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
ihZ/1dN0ZYfDAecg0XZ8bnNYNjOC8xeKPXgVe3WwD9F+kaTa/rzwQFWvar/3DJL3rF/00LPI5vMl
+Q0q3DMN4UHKd8S3tiWY2cFrhCa1LRAd1gYRQN0aZ8OldxTvOblud5afA0fryrEgt+KbkNPQPlve
G2dxz4O9LiSN5sgcuZhY9whF3s9C23kZ7uC0GN1UHOxMsBWkqrPCNc8cFbukMMXmY1XWGK83hYP9
RE1uRwVQMNV02kYodcs9m9ucjNpxMbliXsODmbHvJjb0H3tLVtPdqFphHDI70CfzZO94CUj/rogp
F7gRY2aJ3AVdo5/Ryx9q4fXY2Cwj5E40so8d1HpFCPGeXvWuhBM/hPSw5pzgfjG4gKph0YZyXCkx
xKmbBcLqLcqTaYATifsULM5ChmEwgy2RQN9w9QVEQntEol59P0NHx2ZAqmuFv8No2eb413PiF5fr
+LuE46oR+y87TXxBJOOyoqfJsTXkeytcfPqodoKHiDhculuegXBs8TluLUbJYrnUvI31tfrIXHEQ
FPU4zrA8mCS91KlJcXgJTePKu+UTkvSmGv4tAzQxriSKAxEAVy/eD9SzFYAM/giWjUXNsoxANIpg
i5YN/JGZN4yu8hR/dgjq7ovF6P4MK3KY5dXtjJ8xJSlkTVPO65GNv2Dvswiel1qDUsb59oT1pU4G
FQQJH1NUJByzaA1mjPktC1AlTZklhA+P0TTjKsXG25Vedi2U1QXAEeBdr8bL80Ru2mc4z5TrGdVG
mXdN2+Tb6RkZj3A+HfLJ3aaLJUM64i1CSj+a61RmC2WTF0scQVT4jO2ONdkOElHMqFAU2uNerx8w
l7DG6I0cl0MprpMWnX5+2AirJg1TMhIvyBrbRwtGOBp683UsnjokGy3V/8dSgUdZyt04CnaNxpQX
Aouxry5Dt83V6Ozq1+cSkd1FHVlhHOiSENHnR2jqMps2HhJgENgQakJHbYcia/wyYeHMRWWFo4tm
vdN+7V3LT/Vlh79T6TSN9rFYRHLDc7ukpvcP9P4dweALnWRKi80IylildN11XMa5o5pcmgMudicZ
yvnB1jfzy0DfsVK62MB/+PWWvgxoJSWehE6szT/F2qK2wC6VxEHs9AOyz9P3HkwXvkcCcZWD6O7Q
f0BhUPG9xW70/Q46stW+gtUuayFiZBi2LR0x8sFRk7J0qE2Kan91rFBayqwox2os20QPQ2fvihwh
OgCyxBOEq/OhhsQqqEr8oWrE3p1Ac3e12uKE+Tt60T/OFcD4M4gAJHdAvrfNNta+OHrCX15zUkb2
ddCMjPZ/juCAEENn4Z24uB3PjrSE9u3G2pfq1lyZB8JoMIHGPMnb4mGk89BpP5hRb4dCHnz0fzGb
Ro8eU6cqFYoHu+smvUbq7ZFoFvhHMgeRnwcj8CQ5f/kx8xybHTI3aFq/oq0PF2+g0S+K2HGsBVMP
fYAGZQo7Nq/QAlsYJULiAPFqbqYOB62m1DTdscwoW/sBJw2D7lofbxGhygZuMCyUEPGQ0ZOGIHV4
6nMOdTZYpZdtDwbZnMtma16T5XOR8UA7NA2XbnQAx1lhELZ0yAn4a6WUCIDpWH4Bk2U/DfXsHmlk
S5eJe+H3QQQPc5vmRJEwDRmVWqKkvUSiAupGnnQieelA9/5tksHSvr4edUlLZnp078e92NXB+Wt+
XwtEoUyrYthn6xitQCjX776M8ytvfM+0CaO4SJaT+8RZTkoZPqbmwCynOGdYUxx2NpVlyU3y3VC7
Gr0WXJogRChvGFArR6QJywVCvIaQYGovssYXvr90+gFjj6PgLzCEdAZQSmlQjgMlnCpLr69PniCw
b+HdOp8ECOUqwE06cw54uo6areSD/OQiawAvm37PMrx+RaiMh7+b35Qo6tteGOpJT4YCdmKu2xNt
fWBSDn3fN6rwyd/HgqcBGSiUu7RQTXWqZaXYG9lxXyRB87UzrZ1qCrBtPZpGLFFKNDDaw9vCGAuj
g7CdH6Gl0TwfL70tQv4FWQUCa5eyKBUzbwmtxPYU7dKlozgHexV0bVqLDxcTU5s+XD5nbQ9s8EPB
hhiZQ5KezEzf/pxNZX6841eDl3pXRIDs5bAm/JwiyJ0KDCqn6uivB2xCsjKkoHkupEM7qeeeTScS
JAqwDA37sNpPqLh2tFYnuUa2q+KrjwKHSuAt5qgPd4zzmpbnZarqc77ZGkBmoXKT88dFjt29KFfB
kb+gsjhws1eS/9xMs3UzTzB7653mhjA1IdVdFQSxNZysQYC9vlZ50H0/x4HnJ+seeRCPTTx/z8En
MUPknj3Cibz1TE8f15HBy5+xMRL+L5ORM45oZnTpKhs2rrG4SnujDhfeuyHcmWItgLPKtA0vzs1v
qhUvrqAJ9sr/FgMSji001i7nExDFmf/iuu9ONsu768wRlQluiIcbRij69RN1t+al1hyWrFmT9crr
MO23mo2n2zXMq9S2nFO0p2SPYwYMXeDF6LQVO+/5FjXi7ectL84R8cGzo7U9QxA9bRzhZe8xxPVn
wNzLTHByuwR5tvy5zKyMbcOoceb8oDt6o78GUPWY3qeSek8bepZP3qmigJozL8ojbEE7ncNCq9/5
3TQBj5b9xWaDvgLbugUK5G8j1yzc1YV+9NBP5uoOV0xgsqv2Rrg6Edt3qef/WF83JgsDPoVfBsGE
yNTGK+hqWnYgJ6TfZdu0osLYsy902N2bbHa+AlmRfD2RA23kVhAeEvGMz3XX+u6rNeudr8kO4r+K
bsaCJGb02qE55OA9CS53PVjMvZWqIEUL3iXh2oi63ZK2fQWHSoyJ4RQnBJucZcy0UchlI+zkgcS8
lc1M+xbb5SpTExTyX6jQF29pO+QEUPokp6CoPX7GUI+u04Q0Vrt0eHrHpFIpRK7X9AMO1Yq7b0M7
81xhoO/4dvGwe/nHZJKpoqv19jDgosup4Cpsfg8uabp7Hv/6FlS8qDo8zbeE1HPKT8Qf9sTI+Ca6
HVlb84aaDhzcsraa2zBaCrFs1TYZWwLel0n0yjW+Mvi+2fixyUwn+4KPk+8+Qb34PPjOVY5WOGwL
JVLmCa88fdMVLPiQBKiksbt0Tcttten7xH1IA5rUGWzSsu+pdcJK6lkMiab7b8JKO5URIgkjMMQl
5vJtd7wbePnyQ/9VTD6reBLjC8Fjs+lsABjRhGCc6XiL5YXr8P/JcFOvnlqW+CKPQY1nRd5HwA+v
a5UmNUVA1SQ+gZk77B8W3LwzswaOln2QROjVe1bdYCcswm73vyV/3nbKAFwUxI/KBCom9zTa0WXp
m6SfXbjlUsTtWnTMRF+90MwC62shiYa1brinT5OvyuGVZXzQm7s/HENAQgLqm9AS79AQJsfswVnU
VRbjonoaYIjFlhT0AwYBD+C1oH4yofsro87PfxEwI/R+pFPhz1+L7dnfgBRRabtHyc5uH9hNY9KT
VyBcKDDaXTv4UWykd+9zn+gxAVTQ2EjWxYFaQwSIjaFUOgjlNCsdwg1EPfhF1V9vJkqhKJkg++9j
fVRmbD+l2rmZkhDkFDs/rqwIVOlvgckykX4Cjt1tHnSkGZXe2op8V+DwUmVPBsBThJoZnmRFXIku
KjyIb9eAgQKTfS/faNo87QN6S+CecITx97GmrDwbETfpI8WMXyGH/yv1xAjaXNx4G35i9GJIkty/
SIgbLyMgw34x0MX65Nr151TOHQaMIi/YaVxiB+cQrT5XROnSwJNZPMMbemXWEJVbhIXGA7Hz5OYh
YcOAGhIyMijgmXf45AY7YscnVZ73TR5tM1Dk5xE3h3EWd/oJFUkEyyHwg8d0l1JXnS8avKifgUot
bSVShhVHD3lCl1Zqakablub0s/QSLDqP7nGWWGWJbnUR+S2ScVJ7lmgnxijsz/IuqZSXTn/fntGO
vb9UjgxtJ5xtlthY9O1QlbplpfIxWHdJjEykfaOLT7zYi7AOaeo++TIGN1tUY3TAZeOK0rRxrpLv
RDLPX0m5qGKRPe13uf3aqhGdDsUFMr4J1MoRgLaRgD2CXVUA8U2HJ1ee0c8gzoKGoQwBCH9Uq4EU
xqtEzuBxfTgJ4ZBdjDnVCCJUciOnWJUwIRiCVFmqUMKaqQg5WxNFfLT4pKXV94xKa7ums5GKXrWa
xDB6Ru+Zr+ASBa13IkK3Lmm7lyNzL5mSVQzm+ua6ocDeAk0tHmLRQBryLh39s/e9vp2WRcnPkxEF
Z1DgMig/cTUZbrRPuIBBYkMUKDmEIwxVDvW9ay43QCJncQlskGYy6mzSO8UB4p0RYKCZJ8a2KMKq
cvjBVZ9+tbWm5q6/YLiy1gkwwSYz93KVR3zInVGk853KnICIYRspr6el7kScoKLzuE+ilZMvuy8s
UIXg69konD+c3sb6ae5K+pRM55PKy/35g5xVTLHXiUInGzNYdDmLhM8JyfVSd0nH+0lus6nCGUn+
xY4HlqsxVuOuACUjKiO4A4AC3Vw2tQBctf9a39Wq5JXK4woSH93k1XUonxN/wEJuMKCFCeZ7oUMY
A1iUntrtXFScYBN4BxHl17J6IgQm0XEpMOA3k4w6MVlaUCKH9qS8RoVkZlmiFl8JIBsND6xOsBTM
39i4Y1lg2zmclCGQejWnYQLwFV7XIjcqGyKl54DEw0eYjXcNAMNYdlfdtkh8jDZFz2pMNkbHx1pJ
x7RHKpqWfAFg3FWreRksg6CIdim1v7SjIud6u65TDVu1MWQN6Z74uSQhB5gokV95HpgF4xZalDN6
DtEBU7xkCRBtZXotRJVgucKTCW4pe/bnrF1Yop+WXPB4ESc83QqjuwOpXbvGjyea2b86GV/nz7MB
JElaWfp6XGs2rmS8Utj+2XtWAE61ufYor6MCS0zV9UmvFzNsUWygyr+24DuZ/jipBjIPbHtTaHTt
GkZaKNalpLAoFbAzQ2g68iFO8nzx76R5RdwyPUbc78U9zhfmsyXK4tkwhgZL/E9YUnKVxgV2rA+6
3QobH7WX8Wk9Jqc6A4N3K++6NzZhBO31tQmhI+Al0O5fbZWS1glWFe+2tBqAostCObvEB5AqxMqe
g9pjkkRnykUu2hq8MkXJXoMYHjQ2s5L0bnPxiDapSfTDAiwegXGg4mKZIKuugRn/k3JLtGE/EbV5
SCBMOhEDtefgtnHp1UgFiTt4eIoIp7LM/IrD40zqm8DtQETKMlhhFHFSnCNeHHJ9qALIrebGoQGU
s/Ukbo23hj8X9LvL05UY8N9gexazVpjr7XXYVljNDEMlV5/xjmzgqo91Q/1u2sqIkhNeU6XmtPnC
eyxoxMAkYH1e1eBEDgOX2RLjWepSYPQQANbe1VGZ51v9vahNmKG4uXB5anPabos/nj5TeQ4nhlij
b5BodWECcR3Rs0W2BHw2WIoRHrH+E+mJEqSJdszuI2R5WZMIIc3j0sabsuQbayb+HlESG+mtGWiw
bCK/TyWsf5qz0MWhrtKfujXz/sZ6J+Y8SHlSMQxkhxxYLegSCsLberE1rc1uHHOE0czlt6MjrqGB
amCFFPF9t2j3YUD3GQpWOXxIo8mnHM1pAfAr6S3t7Bk21c+pImWt7De76t2bvSA3F/o9UqEiutYL
9wqj4UIWVPBF9ErEfsJUjXk4POZ4ithSD3BfCZURQ3OQw7GNhTQT76ILlf38hQ/W04D77faM7uDZ
pMkHPFf7bjHsXXRcrFuRUMWsFrPE0qo9u8mSUO6RtUhjSc9RjyRLvsACShHxtyWWjQXOacT4mDGh
Vps8brQNxe/FJXknRg9OsTzRyYSAib1rq2eAogEBZlhoM8fGQS6iHPdQeFT77xmFsQWB2Q/59H8A
FVzNyuhq4MEMHubebrPzvtB2whjgVWd4tqgA0NWcqXZpz7gVWGwtZbwbhWmegjXu/FjVa+pl2NVe
XkI6gfHk50gkCRZ5RqkwFt/8ZyICuPrH/aW9uyKdlB5IsLZVwYalBnCT1bN9lABCANfDHZ4jQXGv
BjVp9hrWfTkXKSoXJjNJHZZMZd4PWx3dRz5I7lYEBuTwYp9BhfFeEaylQlLKeY+ar4UadqRM+ed1
odMhEtXeGH7yhsFwAkGQR5+KZ6p9c5HqwY+v+AYEjPrNWbMUDD99RTQ/VNY7Q+85Igy0ytPwvkoO
PCSCKevj5vW6HfTZr9BbZLcb2HqmP66emWxmK7kFKSeVD3LCX6XZ+QCiBklaXJkMbuD+9EGXVKCc
P3rFVO/KZuLFOVDbcZyoVlE7HeEBcHC8v5Dq+oN7AE7ioRL4+a9MeLaVlllSh870Sy/wj/LitTPm
bamo551PmgOo69639sjd5xWxykA9sYfPzFQK3w8a5RQpgYlIhPHTGeNCF1PE3r8VTmfdQo9qmxvi
T1JHy5RrlKxmx2cz96oQzlM3KOnfxg0pKFtz2MYvHps9AL7idlGG5+pN4J5fxDZXaPW0foKCDFpD
4xZr+MvP0p0IPT4JSCgbzutWoD1VnmMCnAJXlDJ15cHsWdxhPN6dRvo6FIyuJQDuO1ja4ZA8YfhX
cz+/fX2yheTx3wrHE5E4SGfR5jCetZBzaC6AF1IOpy9wQf6+8yqK+v4Ve5WnMoCkYwrpz8HPqMsr
pulKeXMN27XMemEeDUcDbN030x2rLV3AuLHRZpCGTspGPmiNeXePRyD7nqSqpOmaIaJxgNOomJp+
v9DqTjt36cRsljrTy1IdGnXMlgDA4RIrH/9FZUI7Nkd+tJeGeNukKBHBT/Ja1kVPhM06HWtfMCvj
IMttM7cl71yDgjyFswRzfqNXdlzwfxx7M/eNKL5D6RHPXdCxWwT8ll4redDmjvfa1Jy7PlZAY62j
SwGoTk+oOzolZdv2KXe82MQsZdqiw9QgfxwU9PbBlB0aRqLISu0ChP3ZtTYPFu2wQ8NRIKNGgXvI
TfAJcySFWad2hRUr8zSwXI5whScsoR44eJX7jfPl1DRhMULnPf+aUrJS3CESY2Uf3+G/vl9etNuo
HQDPWFnUATXQc1IWAeEQb3K1aR6DFizqKJbve77Acy1SSLP7C0xsCjxUt9Smn6svMYcW6X8GCt3e
68Duspwt3qrsoVqDCINKfUPIbr43cxgwOfZtG11F2cMhG6GWwK8f+SwXTntAC7DT8kfvGJeYMLzN
g9CyKyJCmgvhLNmoWUVY12pB1gKtMbXFGxTalAhQ2mSKtgWs1KTdHhf+1lVYj83xJ6dcFT5JnngC
HpH7ZqzxtfoNyVzdD1e+j+tt8hO241Xamr5q4JspyD8A+KoUozF97fLOM/cgmegCEENCcDoHoTQP
LS3WUnJxbWROLSGu0J6W20CGjutUjVW7fLsuLQxlTVByOaUBRQL5A2WUkO9miqNx07nw+aru7TIo
z6FBBOi6EqtJAVDv4PIaJ04v+4+zykzEquFZmZVXlOz1i1p0XLM2UegC6OUyLpYqsM+mViT6KzbP
DljtKCAvwT7MdbFR7JXo4TRn4tTwToaxd3hO9AGYtIRlpLCYsC714LbRPY+v0k0MKIluXIE1F0i/
Vqai3B+YPcJ9LOI0nESxsN2rYlN+zzg87xom73o7EjzxyMJT/Hmb5nKI21jJz8WNhogp7NbrWIJ8
EAXybxoileCgOdkPjnX2XcicgItzZcMv9Upv873utYIGTzztS57cTDVb8PWyfJokP/iDvnJZqxBt
TJtvGVXVW1O3dShrcV4rRXfqICqkqGeMs3NVzriV0br2bgxnofMlxAcojIx4fAXay3VPWIHCLAGi
rW2KHig0UV4uTthPlgQ8nCXI15nps1qMs1jMYHmIVN5ps6AafPr88roUhaLdmEG/is9tkwdpgjRb
KHOQSC5s2Q7fbP56mcqZLEIuXYfaRJTTx4tHHgn8Ta/3PUD5Nx2kYujAo4vA0b6aO68FbnFUrLyE
eDZh6JpcE2wBatKURUOWDGIUXPg1LmRSzhmnniL/TVvDyx4XLSQfdiXEGb5xw2+nBQdODh9Lyjh0
g8xPHDPwWeQcNID0w3xXFy7qWMru0jlh3kbkYkv7tKe69Hl8QIV/O0S+k4pjo1fpoghJKHW3urSP
053aFsWteNw4NcmJ8HtjkjONRm2AraygXhFdcVVP6aOAOEZvH4TaR/YWorueq1zhUxCyZIHRXVon
HMtyMYEsbt2baBrzlDUKvgDJUDhTvmH5jn/7C8pn0X1hibSO914G79gP23yS/5u+rH5zNWnzOYhx
iP4fGhUsaHAUy7wmvHI87R00DCIdM8Wl2K7zhRVECgpW5dRNt6QCrdKgEIy2AcaxFEWVDciPasbI
1JrCcIqj27TYm3QpOxLANLq+7y/cZIyj3YJnvOrMDXwc/1Ezg8TjFZNT7LzNeeJ0L16LGciCZt9k
LK69xVGxjwoQMUQ6Yh/pNNOKQXNlQI1WUtjtP1DgbGeLbDAaNs6nthnov8f4Cjeu5ePWWC6SJmsZ
Dh4IvDs+QK0ljtc1z+wXhYRwIcQp3NyVfzUIAJt23I0E/uzm9AEJEErDEc506Gykji9i/eSXUKft
ChePucMmhOgqoyx9LQ77EsVBWsLTBVpaq/v77xs3J18/nfFMGFryOvCOHv7kQaQWHvulwPo3C7Jr
45vKS6Udo054DkWfp/RZY0QR2q13F+MW7NqiSqtl0EKss0nlISq0TGfYpulN53n7pKuBaKQUmzyf
l7elk8DVRtOLmW0MqhBxLBJpYSVn3Adf9AdZf7Nz4x+/BAs2fYycEQOmTBzKurQ7bP2dRpY27fZW
wcVj4WJyMPzHBpVzroRl7MuGG4lAJ74vheN7sDuUNAUfFoTkGy390D4UPXK+fujpDPfh5M4FW82p
cF773a22BjLAif2dO34MTHt8Jk7aqO+DY7LiJb6uJeu1VAXOeWJT8q7lKoM2k2Fnx1jkev5V6Fv7
Rj0LV69h5qTs5cW0yAh8uoOBFK5bZXunk8mZwcrLvAoMcJD9VtT5j6k3s92c1WXtnRgDmQJBElGF
jgurV/4Qtlu/Aq25vOyRmYplUnEMFqg6tZ0PV/LwL2xWki6h+KooQ/5fI2SkPvMsrQe7gXASfBAg
FfYUOlh2YU01YJuVG4udxYst+nlLlR471uBP6mG2SNRpbWe2p1xj9otwoas4uURorqvqckqQBt6I
mSM/nmy2D1EdVjaxCT0ErBTxusTB53x3UTt4dcqfFgrOEqX+3JfFASpVTs+qZhsjXZNepr5IG/Xu
b1PzDoKg3zo5SieThMqHYiJ8XMoL0KquOyH0QX3LpE5nKJJ+UR1vYVNoVVmmRPIrS4UEs83yCK4g
DN7LNLufCETgbDok4x8IXhAjQiFxhxya/BICtaFHyIrAPHf1DC+pK3iGO/KE8Mb4J4DzlI2ubdPg
puZjc46weBs8MPwLecMKXVOe7hMOxtOgDOnQPeZWuWm8qHAeJQoNAo0C2WJQIer91ph0L82M2dZN
9yubJhQItEdl4UWwy+4wqKmh3M3yPkILIDI5lVWQhSs5DLjiH1uHZvrRSx0JiojTtCs3VCs5rPbH
qA1xXLAIdi0z2WFTU1BS1to4JVimGdOocWB5aBPP0dFe3Wu7tXRRlNGJDcbEO4wLnqTPM1EuLbbL
SYgNpX/F78DXEsDNS8hupmkXsa+Kz/LcHJEZuD3K1n+VYHcjLXR+ITRh/vnPPxb+XHERlK+IqrlB
C5cj9yRH0ZSX6MKsM3ylF2O+duLcB0cV8nPr/JW0+p6IYCDRCXcYNJna1nRcksd02E0fHCpiidLa
55EBhP+n7JZPaqfIcySuBlHjRKl3zhEgxoXpowCCbns6tRT8O0JJfD+b+RD6UhJZDcSN7GnYrec5
4JSW2PBrrcLqG2FgR3rYbB0WXeojUxI4H8nDaj4lb9dT3qkNizwtiCr7bQXmwFmDlcikOzZzXYqc
+YxWY5f/96No1JEI8s1iZPQe1Bz+hpbZ+Av+wffElm9bSzt58d2n1FoCXjcQwy+cN0oeADtHGwJq
erF77Pdz4FCdOoF+BbKKn3K+v38/x7MjuSqrzC2Xz3Y8OgXP8TiYrnVLMMMa7ykKCWkdeW/FwP05
HSY9gkSoWvecM5RyZ/7olZhFbWk7tc5xM/RpmanNn/lht2+YCjt5hk+clGZs4UvUJ7apsaBpaugW
d6Om+/7kdPW/aYTVE43gSpEBHf8yVKJuBTo/cDdz826AnU5FMvfsXuNvigg3M5TUALWJA+ObrNHA
LGigmIkSWGseIETIvPfDshOYj9JdnT8myBex7JhPBbNxohCneYuTA+bL/QlcNbiId0kPLLbkDKrt
qmSlTPqllTXwHB1orq7Q4+Z+XIvzUYin+PNDn5gqNitKuzCFGEkN0zGwJWp5Yj/WFEfLZ7ILOj0a
qtUlQ4ub57P1R2AqUGq46ohu6iToSFRRcHlFtjhxXrf3wg3YO46TcHYjIE4y174POW4i4kDQVTUO
Xd19K1sH30WoT3yPfp1pvacPd/wW8uJ4NygAV6MyEG0KWT8B6xerOJpbmAWFOFw9WYIHFVqtnNLs
yTin3Kn54Eqo6rdZULIrWyaNd55IhcFC5ZhXBkmYbj0+PYiNrfOwn08gDVMe8Y9DRTZO9ztl2IEn
GR2EYa6v0xmJ0sfw/6c4ybyWPGQuduqEMmqulcYdASFhGYUF0K86y2KNMN+QlMq/n3h7AKMLdNrK
QIdXS33IM1OrgnIky5dwMpdNqXk3wGnLqdyzGfcTtJmWAOFOR2oe2zVPo8hYtm8r2LeT5FPFTf00
D97oNX/I5iOa4NmWLS8Fdn3tN0KHU9uXRAp44Pnjz152rbSrH/RbcqMzeyrBFyKDrPaxyaRWyagq
1I7A3DscuWclPNz29rYkJtklZAbc1oKHPdY7gL54JKJe5dFhNMCR9KxEpg0ia9mGGZXorhNQwCHc
30jw1Oda1u2OtK8bUX8cmlFVkdFNY7P5xlWveZFushn55uZq0rqSxlKHpgqZt1lIlvzX2k5BvrFl
CtS8cemblQaJc+j4UWxyxrurIEnssGWQcKRiGNUAfpTEZmnuTxLkXBKKxaFoz/ET9QucVyZhX1xx
58oqFOj/AYV80Q/tlRk093ecrrUKE5yBAHonjgIbMojj1dAq1AbI/lsaR75qj+rk8h5ndkW6zDRw
MDW1/fHm+ZiXoZsQvdS1NeRHvEkg+iorbr6C0m/LJZojMmsiGr7UgBCrCIPHFl6+XUkc4UwOYaPV
jJt88ZwnCfbk+bAQdid802mRFWrYIQBKmS1vabVG4jQksHn4HL9ChgDmay1scL3oqYB8TIdc/pMW
pe/17YvznKfHLM33jGrZTaRZB2DpaG0WUasMfb5Pn0tPATBCW3c6WifQoRCt6UVgKbC9l8qmhGBj
xZ2mhO0xC92TFPtZnCe3p09QbE1e7f0RDSHmmGMhVKxHP+3C+78rYFs8LIF7miVRRWpco8yLapxw
QApVTCnb/Ycv75NdJXVGX5XTW+YqA8QTeJGAL1d7BSOvBNa7y/kp8ogtxOdqjUfBZdRGNzXBzx+V
Nz4kENFMXnjmAgJOYyKcIraHIaEIJrP/bPGuOOhsFakZMji3vybuWqidNUcNc3Xw5FwD2+yhjEnx
uCX26dYh9kya3itQKTVXUzRg6lWrrwZT49I6/hf/B0y1D7cJnVIAM7liv6ZtutVrbPu0Yrwsb4WX
o/EXkWOFoNBQRnSbsP0sMCuXoLFy0YKYEkXhPCjTFfiXFVfYjGqfkARrgaJdfvMha4vbZpd4AXbx
y+YNdwU/UlTWCO78dcpJWldRqRQFLAKGjwJ5Q9U/znttejpItWZIDqwSz3KdAHxQAZze4f+e138x
Rxj5JVyUU4Vs9wVadz+EDyu1koKzd4J0q9yboXRTibMLaU5sS/XYgj4ZDmMYW2HW7q/Q7SNlBsxL
xSuJiCq4I2mDsnzMvTxbWJyUca5wjKfGU2vMioX74jUAwCHkA9HXQvWNKrAceySHDKq6Lo5NzpXC
R/m8b1/MMrO3f0xP/YCrx/E4GRpXzgOBDqH+D0+8NOf52mbXhQKKRYj7r/G7eDWXwkUwJo9qgdzQ
6CsSKbXRvainpvly8o6yvjSh2T0aFpAwiz+8Y7eK1VMsZXaZnet5QRsFQrFs9tBb2cDpRf2f8AFR
06FueOuG15Yv/X6oLVTo9FlZ+gTzkIiXYoEUAci1aUxCuhB30rxcVlXefNMV2ePxMb7X9OUeCSiZ
lwWZkEudTDSwZIxtYA39Ot+Xl4kjeo0s1A6OXOkaMIJyo2EuOSkryBmZ4VIO9pixDPf4VVOlFy6h
vaMMlmEw+m71MuzzuuxQxWL0THO0QNw9p2S2uAeqB6DJ6MwgY3Y/zKJx4n2bXBtKtadmVVNlmBgn
pQktmvTAuWgodi0nl7I+wKse/LaNY4P9eU1oDMs6kKr1zZkHuUlkyEKnteKKynUaVra9tLe9zE/5
0N8dI+g7AxjkODaDZcKi6wnODqnu4UvIg7xu1qGWjLrfFgg7oMEiVX5Bxncs15BKHJiw3HY271IY
1aUe5Kzr2JVlxneBao8rDiiA9OGPqVjyoeyz6EyX76J3iGibRgfgTPTSW0z//OBRp5doUpAefy+C
cjwyPOsUFPi9+/8it7SbMtrua1a4ey7aXIag/fehQvZCdlFORoPggPNoX6jUwbqNW/ZU5oz4Ckxe
WhLW5mf4ijQVnG74Zjd1TURDsq0DRX49s5bU2SaISxguH/6Toxsk2jnTwzevyZwBGgEpUB0Qs3Ho
/vxYXjxVUh8GgKlSP87w6nk/4+ww5Ep8BFaAMkfFTkw8NNFc5WSOWPuIlIQWsVFM1WCnBtICJdsR
fVbheYVUQjhKepSv3gFmS6gftqWnCX+BKPEkEWOWZzdZErxP1p4AVEUaiAUhzdWuDoKpM0tO46fH
clwC200cA+W4acLck1c5gPp8XytfMRBrxXthEsrIgJG2KToA1FmMc/MgdmjOaTks/+Hx3mJVTgC6
1BgC+coWh16XhuKaW/zI3MC/uJZjRlcxeVnPTIXyMc8DDMQtKm04x7YAJ+NFCXnMJVELg0JFKDv/
kjiG9b+bEdFOfAZPk6nrERsug4WGvpaz6p/yepqa6s1TUS0dGqah6bEN+m6FuZO9uEyzp2SFiRkz
ZeyOdGDDdpxTymjTgCGvlyNaljiPpLB8iGRv/dJ3mNVB6B9ax/2pvPslfQgAe7uATS2jjG9rfme+
XediksIV/a43oG3C/XL+1HeT23o2ejIU5/700isu4WTKZp7uf+M3/p1bhGja2nKJ5brZ6qzQYHHN
bGm+lwtgxTX2DkdMfEfrlx4fZV4xVvtb6NsbRqWnff1zLolW+FezT9pmwFbn5j3URTFd1/aFhPoP
SSdd0t3PSoG/7VDBb7/w2P9OWDKnFLq5pc3v2mNSIW+5CbwURxSnAYqTDlOuy98yflnNGxa2ic3H
TDNX74ca8iuEKHyP9VtY+5kwpQHfftwqnPkfKIvWh7y87DHMgC22JBXkeac2C3F4BjJ7vEcp8XDg
U9gXPgjQPsLCQ3oYXDigaDvT1Wh6HFytxf/3bXQc2D/XanGVxC+L44nBOtNHYCh6an/Tx0JCTPOh
sI6PLykRqY6/IHgWK6tbBtSOKajpWenEbhW27/7oaDXvU2Blxsp/aDr03Ta2pbo4ts5g9Y7r4qoa
vewLGc5916ZBZ9e698XEIPpX3oX+rfjfW8whPK1fLzvVWDaA02WsswCB2XTLt1lJLpLbSQZxqBKT
bWRRur1pT7unkfiL4nLsCwhHIV4wp18inbKdPxOYwpy3GPQ3CzCz2/HiZQlsVk6oO1/eiC0=
`protect end_protected
