��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�CM�3Dm�+�r�)y^��A�Y����ޏ��B�h��=M��SO��,���3��z0�}�ٰ�d��J� ��� O���#M�[�ԾA�u�
�>�+I�h�V/Ҵ���y�]�r��^�:��Y�V҄L�6�}��/�@��su���f����g�^�/�jԺ��������n���_O"R�����ײ6���QiJVs�/u�����X�UO(kpt�~fp`ɑR�/��i=�����:��Y�d�����ĸY8��&;k�E�z&H����y�m��C�>�;@~��g�����`���X(5fIp2�=�
o�݌ڟ)�(cZ?4׻�vPG����T w=�2$�e����8߀db�TR5��C�v�H�a��J|.g>z7�(�cDY�DxV�ঘ�.��a�X��Y���{�v�0�֬2V�2k,(U�b^w�����650�s+�{\f�x�ޞ�!�����q[�#��i)=U��X,��^���l�A��R��f���h�F���ͻ��[MJ>��E?̑���f�����^AD�X�Vn� ���U�xig��ZR/�L�u��+��-�@�p#�>�d�\�7b��4�q��n�?��ԼW�WPĖ�ȃz�c�
���������->;˳q�׬bѵ��<�=���?����ƚ!т��Y�:�	���u{g�前ٯ3�������g��ovRk ל�	���Ygd��m���	���d�pOz,m�^�d��w}�h@�'�^�7�]Ӱ���"�U4�����]�_�+̚3n�F9�9��gk"E}/�7����Z�4!�juY�ΘL�Z��$@渼��!ri�g�w���xܹL=I�B7�%��+Y�N�l�6�v�W�DO�̨�N���<��Y��D:�p;[�$�7�{}�3:QP��*�y�̷�=�1崹�1�\[�9����lD%�q6F������7���VU�n�H�F�G��*��#���VG���M��!s�E_c��J� �1�d����2%S��������v��_E>+n�gⓑM�m���r����fQ�ư;}Zܩw����m0��<W=NtT�k�q��C �(��e�H����݁ךW�Ӂqq���и�9�,�t������_����;(�'lvB�1��.��R��L:�@lb�NK �E�̎bt��I
�ڈ�oǿR�
ڇ�
\z2�ɴ��Z�S�á��W��!z�-B��v#>\���>�V���5>t�Rİ��<?��Uw��5&��P�E�7���cJuJ�|���F�j�P�5,Rn���W�>w~7]����N&�n�T1Z��.�_����l I/$N��LT�2"���X��ސ��,�Z5ϰ%'����K@�#	y�|�Q8;�a*`/�oԹOy������1�}@�)�+�mU7 ;����G���Bv�M��nNh	��0��̉�5�yW,������ �l�a&���v�y{[���zBXM*��Ӭ�B�r�������t�E��2\��(�Aώ�8<OŐ�K�O*�i������Dv���N}�(,$�}cY��q�
�=�7�
��fkE;���Pg��*Hf��,g2�N���,FZ�o�?x�^�!.:O����D���g|,��)�3d)���Ld�C=LHq4����e�(`�y�[���S����5�Qhiw�%����	��5�p��:�����m�9�T�/!��me ���@�����2��82��©�Ϝ�_��7/G���M���
��E�<o��7"$�a}�����-�����{o���y��{���~ԜMP�$ ��9+����V�.+�cw�uϵ*{o�˚!�/G���p>�=e��h.�)�V��"� �&�o���BF��k/�|��P=����pN1� �T	�cC�y�ZR'�o�pk�u.{̋ʹ�<FAʵ]�+���%�@���>�{���E�'K�H ��r�q��uy�����y5'������=dؾt&�v5�ơK��s���Ր f����W=eh������s��
�R����}j}8ʙ���MF=�/�ގ Çy3}`���'W<�eCv�/��f���������/��VF!w��n�pR�EM�:��:��H,"4���*ɵ|��� r�8�76��u���@L)e��.i.�~0N�V����iU�d��R͵N~(��^�8]I6w�;�.⛕U?u71�8� ^�J��
���<�r����5��E���J-�i��*E�������o�4Z��*�i�gp���H�jioU9`��.H�v�{<�L��@�\�=L�4��m�c�Z��j��m_���*r�'��z�-�D�>����u�R'�H��.ЃD�̾�M��1q1�������@�$�QZn�f����9���'��.��2o���-�V�'��o����/��FE�3����/i�JJ2gf:!�AFn/��8�c�{�& %�d|�]Ɗ�n�� p\O���v/#�vɗ��2��rD<�� ��~�53��3M٭�Ǫo���H���2UȏU� 7�mS�ʘ4m�N�Ys��9�5K�3�U�lU�h�����^MA(δ�/�Z����^)�� ��6Z�>YbM��k��r"./{�e	���e��O�$��ǯT.��F���/࠿�g��p`(��v���C��K�h9[2ǌ-q7��2���'�]���oi_��
�
%���� �>����5�����ũ'#�5�e�|����v�Mu�[���x��'R�����h��q��v�qC����':�Q�)%۝$���R�R?�����wk<dG� ��aL�P�͉Ƥְ8��6�i&o�E�wjc��ݤ��J�&3"�4Tj��!ˀ�f_Nj��>F�B+3i���;K��̢DA3��\1K���e�30��^-�UF�	?f��*��Hk6&�'M�s|id�8Y�}:U�(%��+�D��q��)?;�|`|��g�H?(�����$s��Ճ(TMʣ�f�i��`M��SWmss���y�[ �Bn��o ՘<��P}�V��b���;�>;9��q`�#�ס��B-	�<�`��a�9��K)�7px�Ҕ�[���c����ȑ���T誨yk�m�	q�x?0B�H��㤌O��<$oX�L89���	�*�{��ʤ+\E�� ��ݫ �Hp?�+2����)�_ac���o�A��0n���x�hs ɳ����N9��)`��i���MoN�V�:��x����8����d�ң#��~i��|�@cw0z�P[�cI��U�w��>#s:7łY�T���E�,)�Q@S�M�`Y��/�hm� +π�T7]��R��3���|�U�K�Tێ^�m�~��\�ϼ�v<���>��kJ�{� �m��^C�^C��Y��EY\z4�\.9���M�āӦ�b��B�(���:�r�r7Q~�^�.��_Nt����B��e(����c� k�ya���INoE�Bt�����j��������c���r�j�8dZ�Y����dI ��UpD�V��K�^� }A��8�$`�j�Fq��ςà��Tfޗ�X�����K�7�9��u�b���̃���QD(���E�ǫ>�R��������(۷��]��{�x��+(�Ac�!{�P�\L ���ks���B�����I��`���g75�`�<��Q�L^*9��_�^&�ϫ/�ѝ����.޸"� "h�9��/�K;ώ��U��TH�!ji?��� A��Ð�:Q�ޱ1鲧�_,+?�T��/a/�[	���@�"���T2R���l�"\�8+|��3�v���o�lQ���,T���Gh��Z��(@�|��l���fꎒm�����ʳNh����z�%s`��6�A�"�F�������w�]p��8�j�_�	ܞ\��Cҫ�Ak���}��[�R����Uv}xE�i�����>��ҫ�8up�Z��qI��l�����P&�x��}��9f���_�'���	�
hj�+ܖ�X_\"�=��;�������#/�� pE���8]�?Kp�����L�d����o*����/ɬ&X!:A��7��} ��Ƌq�P��_ͣ�Wx&�֕+�<�/~��+Niɼ���
qM�f[�a�^�,�HŻ��9K�C,r&��kؽ�g����apI������,(�7F�	�"�S�Y�Y���+z�:w�Ck�pg�2������o�:��!!I�C�ye�Tr�}ۜ�y�@v)z^.�I^v�&Ԉf?����]L�$K�+S��8N��`�a�nM� ���;�v�kjTT�y�f�+���8b�oj��$��6C+1�}�3����c;�6#k	��2��[޽;Aj�uXCs��gU;3c1�OOڴc���m+-�����QD�� �x�x#�|���Ů�@?����vaj/?���h���U�� )���Ո 9E�A�6]��r>�H��&�#9
�0��[=E"kv�#�,ռ�Pu�B�E	by	 �)vQ[}ȝ^��r��vj C(O3�>�1�c[����U�#���Ndr8�=�(�@��T��wP��p�>�����Z]���V[�����x~͌���X�0�u�y��)��f�rmsi5Դǐ>�4����.�vj�B&U�R`f-�����A���1J7�Ϭk�pck��f�_��壀dr�3/�^����t���Bc�	��#\r���w����\��r��:� �[�o�� Xmf :2ƨ��c2%����T.*{0g|%\�E�^��p�V��Dd� �e����ú�P�x����c����a��1��l-�De�-5�/�ǝ����D%�ʋ*���\�zh�۬�����o�߲��]}nE�ڿB{��,�����U�$���k���HS)�w��,/�̱E�ʫ!>c�S���0�^!��4ޫ_��`r���#9x&t��^�eNM�pz�]N�� ���(2�5�����q��dGY�̂}s�g:�����r D�F�'w��+�����$Gw��*k\,nBT&w�(H���"'��|�b1�"��l��9�G:Y�sC�:,�GI׬C8�'�B��XL���\W�a�ua`���ߘ�-5No��X�.����AL_C����E5�?2J���)E'u}�+S�<
�|�Q�4���}_&R�~�0�%"]А��r����}GxC�ĩ#�����7-�����jGex�H9q|������U��%W|�6������m 8_ �B�<��ń�;(s���;N�����58�
ˊ'l@`#�[`?��mM\Y����[z��}C����-���Iʊ�E��L4�0��k�S���˹*Y�@q��飶�������{c3���6���H���U����Ru@����	�3R��Jdd$a�>��D�v�'rf	)�$��~��Mbٕ��	�V|{�F�~���c���H�hæW��b�[8>dQ������Y}�V��"�~����V��"��� k~ˤj��F�7Y��`�0gHm����:�ʿ��h�=OA�fH6�/H�44j�r4��f�
�������8
V�^$���*��4©K��*wf�Ɵ��(i�T~�jݐA���E��ĀL�P��b�ݶŭ�O���i킃�|������� �$���ᯨIF��r@2`�6�/�aB:v�k�;�<[N}_���2�Rn�����1}��BGU� ����s*��6|a�'-.vm)*�:Ѐ��j�<��#-e��fU�lq���ɒ��3������,����\Q��E���7#���h7Fb�(J���E���~4