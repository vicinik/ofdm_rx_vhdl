��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�e:�G��PV��wOe�X}�+�1Nܘ����8�h��Ɂ�J�X������ɾ�~i���U`��(h0<������ެ1r*����svZL�S��u:}^��;ra`a��� C@�FW��R֐c�sGRV!�)@�1!B�������� �9??n3FLIq��ݢ��FK!�5�6B6��\η0o�������@��z	�A��@g|�D�Ja7gӽ/_Cn\�K2 -��Ǎ�޺����kx�Eߑ��a�%�>!;̀ёg����	�[�YF�z���! ��3:��X���:|��RF֔�  �?R������a�?����k;�z��BO:��~|�ё�Q�Ǘ���j�td��忩?�'.�à{g2M�D�χV�E�i>c��d��*�n_����a����:ҹ���� �QTف�.j��P�"�i�
׃���˻���7����2:4��s���*��� ���:�A`����)������uA4f�n|��x���E\�d�=MЧ�Z�ɝ�9t���5]��gԘ�Pe�ӯ	_�K��SOʙ��F������Op����n���V�E�Ynb<X�<�*q��~�)����S�#A~�Wkpߤ�.�-���G�Y|�ٽrF�b� OAw�;CEj� K�'�T�pO�|đ�=I�(��P
L��w�r�.�Ħʖ��t�B�_�x�!2)&15�ȏ�%ٖt�e�����Y�_i����c�e��*��+S�v�Q���"��z(�
������Q�uv�m��)�s�v���dn�3�����4���&�,Cw�����#v����rT�"<�����"������fÕ,*���h��y�9�xZ�b3��W�u��S�)�\M�,��_z��<�9��@�\���݂��-Gx��j��L�@u/ܭP���,�5�粓F�<��1P���E̚n�w�4����[���Һ�˂�*8�D���51[�v�Z {%� w��}�[t_�@�<M���z��x5�1ܒ��E]<�(����tP��Fˊ��N��Pg(�O�E�z1��O@\��=\��z?���~Y��� �D�.�q_t�R��em���<a�����Y�P��c�v�ɱ��\Bv�W#�q�ĉd��
���N1gBeP���� �����(��b�p��3����xfкq`�p����
���	���Xn���W�s��#�q��GΥ�܂�u���s�8���At�p��\��nmp5�P�1� |Q�m�p�jh����^��[�pp�w��a��c�"Q]9ٖі��3:��D�Ĺ��{r[J�/�Ch[f+W��͡�}�Lק�,,��g@ī���{>.�)��lkv�m;IjXq;�uoQo�>��jmO�W4&@����Crq��;0e-��+�����G��;�����(�5J���\hRPP#�7lc;b��R;�Uư<�(�	VՍӋBx����ߌ�� p?��wY�b�tC�S ����ǝ�ȑ���N~�&�O%kSCl���(H��l���68�\L�-���' �if�A?��'֢1G{�ـ�]%��.*��C���P�U,�+���o�ޮ����a3�"^@k�tR��Ӿ�D�|�F:��0V}�Eq�b�)�����4&P�?9:��J��&$���V���>�6�0���QV�A'l���`���Ů?6P�T��&лk�l�s���E� �%�Sy�/lK��vNݍD?�����C�g�8N�%Ny��Xߨ�0��@û ���c�6!|a�-`}AAm-K�0��L�#ڗ�����ՈlD#DgI�&��Ef�C��m�s
f�!��n�֭�s����ű��"o���M-G+����-2�V�@K������CS��q�ɿ��z����;>C��Ǔa4j�.� OOA��n/���!��t���Y�X����r=ǫ:���'1H5j5J6�|%��ȄY�w���o�d�C�X�ibE ���;�rېF���Y��y`�0�E48�����xz�}%n�x��� �D��8�w�8r$��:�Rn5
�� �.��/�E�T[��;"��c3�)睵g
h��P��rj9����Fru�%ګ|;7Ҝ�������#NR����dX��,�	�����	FB�'��f㓳�7�1�yN:����qrJ����P볶9��?CƢ�����!
�x�I�����̍��OnH�`����PЊDl�F>�tT���x�ʼ��Fߌž	�7\����'�V���V���Bl���(P��GsIt��sQ.�����&EC���4R�jω���b��o���p��t9�1�o+��㥒���_�gÿ�BF�CO̄���v�� �Q`�	YnX^b�E{%�":����QT�Q�D�^���o������8�u��?-W��G����0�Q͔����Q�[p��$8{��=O����s��V��$��ɍ>&�o���^1i��\���=p՛�~?��cˇ,M/HN�FZ�2fak���#��#�Oo�+��B ��<���\>�2;����f5`��A��Y��9}o�k6�=�mqY����ܕЈ4F��f�4�Y%��2��}��F��zOQ��D�z��e���m�%�8�Q,H�G|�1"�7�fv��M��	e�h���(x�vY�K�i�kpT�I}͟������'L.��LN�KNdt�Uw<�pԜ���E|�i����ʼ��y3q��{����<�b���0���P���ߖ��Ex�B�0�`+����ɥ$��+ڨ�|��-�Q�B�c[���f��d������'��ygƂ�.�8��f_qF���Q4Ǆ�^go�h�B\����Wr�䴞)���m"�����L�H����`
��Y��4&�����į�Q�pS(�w�R�6Z�!(�,�qC���{�d\����������g7�W��q�\M-Z5�æIX����݌OP̎��p��[�#^���ȫG2VY&���As��IO�0�V}*Q�,v��3}H�}�Qzf��1��o5YG�g���r�1��ep=̞����7��\Xt���ey������e]�c �����<�;�_k��-�15��'Vgvq�;`I�:���dF�������0�TA��0�q�J�&�%ZY���3�/�*_L_�!��'C��h@Sa�_;Ha:�
h�O��1F�����v�Tu@s
G���8���J�ԧՕ%���Ȅ�HE��(������R�Vub�szi���
=�v�����ײ#��Y�Y���t�%��i�oίoEܧ�{�-�W�R�#�u]��j�3M(��ȁ�CϿ�|GPt:$W/T�j{!fE�+~��Up�/ja&g�Ey:�|����/|�,�6T�t�Y�c K&�o�!��u�L:��` �@����L��F$l��$�y�^f��N�Q�w�'�w�цy�k]�M�$��L]����ڔW���2���Fϸ!��za>����}�p{(������wE��,95���P�X�ë���߂�p]CF�N*CdTY$��{|/u ��T�]،�;�U� �u�t��3�S8��4CP�}��pY������a�ׅ���0�so��+����:.wS!R���c_�A�PP|Y~M��GW;��eU���>�$�P����R������<v��Dx�Ѫ��K�4��I�ŵ����hۨ�W����¾oO	TA�8K�rs>q\	�D|=п��݊�5&���6��R{����#�׈��U�ɤ^kS��!��"J:IPѷ�����H���ا�qy�5�e� �P(�˟Y<`f�o�E�O
��K�b�}�)�ň�˸w�B#�D���n"��p���`1�E���%�L�&]�C?�Ƙ)�����;�o��%Nv;l�������w�to8^��[t��ԻbE>�1�#����.w;!E���1 w�%+鈵+��?�	�B��z��.A��-��R7�����"DQ��T���98?���6ō+�2�,��l �Ƌ�Ԭ�pI��9X�՗�h(h,/���S�l��
���Q�lDv'���TD&o�������V�Ps�#G�U��Re��Si�H�ShC�Ew\��@���`;@H�)��%��Γ,�AO#�Ҕ'"Պ��^*��/|�8�}������ !>��4��Ӫ��c�y��^�_�	��f ������~A�v�d���
��Y�[�	����7�C~cL����ֻ�"6�����\�������������Һ@�Z�LÔ�{}�ﮓe����j
.ڗ�לO�a���k����]
��S�e��n��KR��(Ӭ#I?�-��g	�\�� �8̳C��UVb� X����P����w�)�H f��-�y�x΃��f�#�g��j������5��һ�k�D�k ނ�l���0B�j���� �V�H������6�yTs7߿�_�����$^l���m��:�w$�9pD\�p�J�2��s��.�̹�� i���>��d:.�>�"��ۆ���Ȏ2=�0 7ߓ�`m���B��'Ŵb�-�lp�O׆:����5���l�XWŏ�$��d�4,x�0�2��}pt��-W�~�3z��!t�.x��O+�.5�_7����������z�x`��ڐ��pT���0�5d��J�[��40|�v�n'���	WYPM˷��c����Z,�U뽍(lrs&��/�e)�y��H�|Ѧ ���t�k5)�
P��J%Үt�k����=�)u�;{�/3%�y�����cS����0- �`F�n�	=�0V4W%C�;������
@��¬�3p�����>�_��ĺ��U	�{��,B�3�r�ǚ#6�A�6����](��nԺ�r
�,��v�4�' l4#	~��ҧ}o��X�ua�Æ�;D��#�ݱ0v�$�H�f�Q��q��:p�a��tÓ;��э��y�|���=�Bú���������šB
mH_����֧) ��.lA��y̜\��YA���Y�;<����p��Hǯ�m����8\�Z�*������.�T���3 ���<̚W}�RN��t��X�0��F/��>��~���KF�5��h�9�=d��*�P7請d|���%Q�2I�{q�u~�~k����1��Z��x��߽��D#&��Bw�����wn�2c7����q�^C<��
��Ĝ�Z"���1���y�0;�P�%��\%:W����b�s:Z���A�]'�n�y@�l�Y�;����cYOnx6�ml�7�v]UĽ�l:��Oܿ�����d_i�Uw� ���P����*O� �!�8&�`>�e8�4׎E����X�f���UV���x�d�%�[B�^籸��Px�"C��n�X��S⬰+�[�#�y�x<����.L��Y����)��d|�vI���aNud���|� ��	L��,��OWOB��Z�7*DM�i��E3(��S��6�%�SF��[f�iGQl��i��s����<�'���wv�BK~������;�g>����g�_�%�>��R��#%�)m��*;���;e��'kf����9���� �	R!��e��.�vtR«���G|Xj�3������9�z$��0���>�iv{d��T�*��Je���%��Z�2����׫5�� ��k$���q8A���|�؍��T)c�a�o�N�/�����m���uS+����~i�^e�����Q3�s�|��������7Q�W��I��4٠kd�H�N���v_<!V+�t�&��p���7���jL��B���I=̧v,V-vE������9�*����:)06�9!?��a$g��k�����VB�8};?re_\�;�g��>r��adʏ���F/�?3Þv�w�'#��ev�f3�F����Bo�ո�o���ꀰf�N�\��{w��E����i7JHݘvs';��q�`v{r�]ڑ�P�s������4줎�8��N`&���"��ۘe�JaG�o�(��uo���'dp���4���uKf��[�eC�^y�/�ׯ0�i�B��t��X��l壙*�/,����M���5)KZ�C~��,�9u�"ۛ�oKYt/H�p����)t�>Vtٯ�N�)ʙ�8�RY��4�BS�|B9�JdK2�(�^���~-�m���/���׏�cX^.)��F@�jɮ�29����6f�?���侌��f�"ض�Ӧ���o�9�Xh��a��˅������0=3lM�m9L�k�/^j}�heT��?����r0�x���#�{g��(>����s����AS�å�ƵZ;pW��������FX�]�����v|�~$�P��&�e����Y��F��7cf�:R�X��4@˴��=m������G�j�i�S�_��0����]V�.��4iߨ*��*��6~�5��Fɓ��/6w�L�k��t��"<����Xk33e�Ǝ�P�׊�4Io�xًNxz�=�+_�S�ke
	v*T���5�� NG7dL��m��{)�5w
�E<3��(�Pʔ��-��j��9�9nD�6n��ؘ�J�)���ܗ�V<���H Z�7?��\�.�-V<�U ��B��Ot���kl�ڽI�,�}D���u,sݶ�t)R+�V���%o���/D��
�c��q����Z(�*#��X=pG�L�k;\z�'�6W�HԐ>�7(�/~$S%B݃���j�q�v�)B,/_<����Fǔ�w�EWd�k�
�i-��]o��?�4|�!q�bw2�t F��.g�X~�z�@8���.��A���4u+Z��ݼ[wC�w*I�_��>��z���֖��J˷�v���n|���N<=V��\&<�)i�G�G2�;oCI�^a�d"z�9x�C������ �`��M`Ĥ��?���_��u�i�մ�Qd�(����Kn#E��NU�a�7�����K4�-�b�FvM��%'����NQ�[�h#8���w������o�yM��H{�PN�����_�r!�!� �Ԯm���>qE~[\�:�&��8�u��.�.�N��U}�/����x*"M:쓻u��l��Te���Ξ!T漼YuE������X�L$$b5~+6HF=G��O��s�`_�O<���b�!�oM-{	�v��Px�����t��gVRu��>k���Ƹ�h�<A��2�-�e~�Q��2�|��|4����{	�;�o�1�XvL���N�.�-��̓=w��hO���/ė����K��Q�d{�>L��.���M���N4w�L��ߏ{�P�Z��S��l��"���t[Y9x�0�p�6L2�x���;yűP��c2gj��-�\�p��a�T|�o�B�H�
��as>r�W�wT7]:<����haf�Sm���/�i�A��}�D��
Dao��n��؏}���G٘��iv�V��.�;��LHQ�>RY����mP+$H�K@�{M�N�=����~E�ȥ1̏�x�\�B���?������d�ܢQf!��Ik^���0F�~W���q�� ��AEqD
��r����2��)!��9Äh�R�_��(��u���m�����)p���8UMe�s?Ju��,���#���C��zE���p��uKI!�>@KOܗ�C�RcP}3I�SSs�-s#_Ч�: v� � �#��{Fec� ��w;#�t<^Q�Ѥ:p��w���2��/ ���@И
 #�PF'0NRc�"9=ԝ��+����,��Β��͠��8i�4֕��d0��k�����Z�({QeT?]�J'�L��z��M
��Fb�1���9@���K��r=;�d�}�R�o�܄/����e��k�����h� �!/��IB�i6���}Ę�T��vǃ�������3�7EW��$�<�k|�����"����<�>�ȣ�4-���h���\�#�F���4�E5��М��Xж���h4�;w�hByB8��v�B	P�<�s��7>�j�����6ڌ�PK�2x��\�����_��M>4Ô��'��V�M!Zͻ�]!^�r�5�xZ�)����z}b\�ѯ�S!Ӳ��_�"�W���sSq��c6Ό�SS$U�:���t�K\�m���;W[31���8�.Jy�7�ߩQQF��lVB�:�B��S,�W���`	��ݙ�"�XWꯘ�Q�l����x�/�Ը��EZj���#V}VHa����0&>�<���E�l��nQ�]��ƭ'�<~���Q���J��Z�2�{m7�{b[��,�ƹ��#rҬ�dzt�sߖѹ�/�Rg*�����3u�NL���W���_2��$��8�d/�)�� :3S�'����Z l�e1����$��5缫�z��-��g|�	�(���R톯�Ɂ��T�[H[�����̌H��,��\9E���e��}p�:r̄�@�Ѝ7��M������u��Z�1�<�����'���H��%g
귇�:�d>Wp�Ċ��*���F��Y��[d"�X����931�">����ظ�2��P�=���p!;=�f������_������$�A�����FlO�I�61�{�������'!U���뿥�}]*%���P$�H(�5��a�/,p�:k��j�G<���W	b��{w<l�S�Y�܇Au92�ydƾ�"��ML�J^	�8��Y˺sx������q�D��{K!�o�k�s�", ���ɂ�U�t�|�g%)?h=9n�Zq���씳y���v�_.27�j�gq��� ݳ���^�tc�xrA��9F�Yr�v��,�D�%���n�Y.$/ͩMZ��*��v�bטx{�u�����ˡ��4AH���^6�ࡓO�|��x\C<D$B�Pd��X./�n�K��`�w�����0��\�cI3�1ۛ�̪o�_h\$��7:���l@�9�QoBv6����v������f�;���Âb"�eI��J����]��������7�()�;����9jq�OM_�|��;OV�#����l#��g5�/����  h-r=��y���m��u��YZY�&�X#��?����jȽ���:������^8�T�{�����<��+�</�I>�bsG���X������>.�M[:��P�A�6�_��Wt�m6�c���W��9(	:�>xȡf�~�/�����dW�T;��'���v�=EV�g�&��	�b�@n7�Km�K�+�F�P}t�r��+X5�l��)�qs]"�C�{]����W�܊�n����޿��gݞ�ǣ�v��D�ʚ�6���vd4�뎎Oy6���yC�a���ւ�����Q�gi�8n�_R�(\�)��%
l�����3B��J-���g
������?��r���,}��Ɔ]o���2�WV�S6�����E�n��uy�?,�-�0�5߉~c��1b*gp�J��\<U��s�WF/�L���w|�����N����lR�Sχ���%U����օ`U�ǔ�>���EV|[2��/)�A@����-�;edل$�|D�vє�VH[%T2��0(y�Vt�hU���X��
�S�����o{�H귘����:*�ԚĹ+�"�Cި�	<ʘkoR��*d!�k�P\\���#��~zY;��UDY�� �N�σb����17.����W��e Z��D���)p~�s7-��`Njpٸ&��A5"(AWلB��[8fK���ྑL����2{�$z[S04ٮf�R��4&V:�e�F�Ղ
��'�IO�'��1Ua�"��5�W1�����qO�a���(�2��zeՄV)X�d�|��Ƭ��f~�9��e�a��w��fk����p���^+�I���!sIe4����;��ҳͧGИ; ��"\�(GXJ�0�HuN�Z�Qv's� ��z�`3������bY�ˀ;�C֙������Y�菵�az%�x�O��(�NI��*�ujne7��3�24�x8�"���@
.~by^8K�yJ�	�g+R���4���#,����O���e%�my��PF�vS�o���L��8Uu~�x����M��><;Z��2P �#7����!&��j����(W%���h���~DY�V��]�$��v��X(_������q� �o���V�e>�ni2�W��4�oY��8-�4Uy���K5���d� !��4��������K>�1�����QH4ӿj�k
���cy
�����C7�tԴ����}7
�f�M�Fg>K�iGZG���U
�4Px��D�
��M���{O������(�@T����EݘY�e~~�~��AK� r^P@��\}�yE<� �X��c�*���WU�c>	���m��̞ɩ�����������Dz�H� ��X��h���u�rM���j'���NN�I;biL���p7��jˑ�+@�Bp�ΎN��'�:ap%k���4�������Z��5�P��=��>�?�G���bPǏK4ȷN�. 6^)�i�bv��r *�3�������Y�ɕBA�3G<+W�m�g1xb`�q��!�N�}����1D��Y�8�� [��oWE?�F�+<ρ�{�+8�ў�.���ɡ�K�f�`OmY+���hea�P�W��h�w�Gbl'��J��}_�.^8B�Dޱ�\Ab��j����
�3�YrF��g�bL���J�6-�<-dUï����ё�)' ����5������fp����jy���c���"�r�y�ϛ�ɟ�1�W�������C�̻1��j�������0O	��>;1j������j��H��gH���!W�R!�v(��=Z����7w��nXu6z��<ޚ8�e=�˻�@��XK']M�J8���b%푶y��X����NԚ���SN:�ɧ~�R@��WF�?r��Qۉ=$�	�����F-Y�<�o��~{+��l~Lb*;�+G��xϔ��k��/��j�k�"|�I�����J_��0��T���(^�	��>����hw�j��P��tݡy�+�~"P�(�VЭ���s�|�y�(����͡�Jj���˶��@ �ީ�Z���$�4�Ι �9�G�H"$��[�%�E�kӕ֋3?R���,��t����]�h�P/xO�\~	��|s�
~�-��;��u�����]o��� �%���>��b�.���=9[>�?�qG�T��3k����h
�f�uo1��͑��DC-~�	;B	��_Oy>ㅳ��!����<�j�;�}$����R�Bq�v���m�X�r��-���2uG"hê�f�����x���4ZBr�뭢j5����5�U�.��;Ц�.�Ŗ-j^��_��93B�}V;R�|y�E��|�vf�p�yzaKG�9�����c�o�O�
�D�]�br�E�h�}aY��	��������[��T?~YG��AE�WgY�����/�4���P6@�
��#�tD���ԋ��- �$ ����dX3к���/��,�%��'�4 QZ~|�A9cZ�������1.d��<��2��� Q^�u�GL�Y#^�MW��שc�=�� !�>: *�jo�}�zez+4a��z�$����Pf�E��!N��6}u���{�o�L���mM!�|��gg���s�����-��I��hw��M	�����\5%�z|��ס#{�i����y�и��x��7�E�� ����.	�L��������<xO}G#���7m�)0PWVg�-7�A�yf�.(��!�%U5"�D���?\�DN�#T��b�w<��m�j�osMp��;H���Ӓ�eOr���M����Z��K>�޽A�w�o{���%
��y8�!�&G�+{Z�ŕ�� ��@S5'�C��o�9�W��^��X�Hy��D�\�7\��S��n�;��Y���1r�LIZI�)���rŷ�,|0O���e{H,�Y���D0��X��T鯃�r�8*��4�tش`�* ͻ�N�Јb����йCͲ�.�}�zʖ?���>�)�!-
Ջ.m�I;�Ćqi�m�	Ɫ��t�:�̬�d������&����8-LQH������:sg���b�Ӳ��q�;}2��OQ��yv��ʑ���ϝm��_�I-4s��7�K���9ݓK�pX�y�8�J�夋�/���=]�4$���Z��9�� n�1����.��e��Ԡ0�������~��<l+2��Qd�1$uO�~6H�i�?_��n	�j@��a�q��pMA�`��v��'���	U#b:�
O1Ѻ�Z�_k�ۉ"����'�n�7�^Roy���p�`O���艸�##�
t:��y"vj��s���Rt<�Gq�B�Do��cCM�6Ha�΅�R]z*9���@����AD
�<x�����V�����I!�4�U#�����-��A�aHc������o��k�K�� )L��h�1��b��oȀ:��"��Cx"8A����@���P��f����d7P�\�����
|�����V�Y7�`�j
m��x�u0�����_nx<6+�I�}4Tá���h"ay��pX+`�ms�s��yKvD��,���g�ƺB�O�n�CZ��v^��p�+�Ѹ�'�1�WHA���P�E��W�Q;K�Wd��C�6�6�I���?_��+���uLV�Yaus� 42>�;���We�?�-
Q�<gR����֩�u�L�"�oѻi��xy���y��g��Dt��v�/�m0f�M43ጷ(��2��	���e28�C���<�7mt���u	��Fj��g���x�
aɇogM�z����S���:*e;�f�Z2,�ƄW�sȡ�Ê6a��%�R�-��� D_5�T��'+���<�rT����y��[�J������WƤ?+
�-/ ӹلF<e����|����
���7*�/����I�t�Y�ݕ��{�@�,���&4���[���Q+��ˏ!�c�=��m�F�,s൧�D�����Ѯ&�A���ec/c-�e6~!��@�7 ϋ"dˤG�K�%��G���R"��b��S���eS��So���/��U�'��j9����8�d����֪̫a���tQ��u�!���:͟X{��t�5C~�4�m$]#�^e3��E��s�yO3��4u�O�sʽ;Te�Q�i���q������[(Dm-tfD�
:|�u���3���)o�M��Q�==���kl}F#�v��?��ğ��	QO�ԇ�Y�O�`9�e��J5'�{D���.b5��2�e��L�ݨ��:غ��w�6�M,�Co�ʨ�g��{ué }� ������v)�OZ���xD3B�y.6zQ��>x�R�8�:��F��SY섭�A�g���{/���w�Tn�N���}6
0R��@�ztD�uK�ɀe?U-2x!m6`E�14�D}�ǫX�F�=߾Z�6\-;��9��2��"E,\�������+�E���	.}&����h7l����{<=(�^LL��<RF$L�BWn�	�p3�#y�}0?K�j	�c�����Pl�Riڡ��Ӎ�̀�1w���9_nS@e��bؒ`�I1�	@���h���gc2;�tr>$�~��He��x]��Tywr$�v����4���qρ��s7��?o;�1h��1^瓗3���$X/�Y�[��gH�.��@�\~��y��*�(��O�Ŕ��:]§ɥ�֡�G/&�\G��E ���A�ps��y*�m�s���?�&à]}0k�@>��`Ns�or#pA`�v"�L���(�)��^����8�� >��	�T`bIp�xtA��{0�|�wj=����b�$@Bm״�����ʺ��"��H�\���+mU&W�-m���Ĕ3���א�j#���tȩ�d���4q_�A�ƙzq �^���xx�0xX���zW����Iӈ��Q%�������.�Kgf�ğ�B��{bND���^oK��,��4�VO`���Gi�����Lj{ �nC��Ǎ�ô杸�����wˏ3e;W��:��ЋS	�
�$�εK��� �畷��D�NA�	�`\!��L�,�r/0;]�~A�[�G6�aT��b�욯������N>q���DE�쫄�D�`4�����T�hs�H���Z���*�ݫ}�f[���v��q�K$ҮF�L��ҫ
�׼*�s;��CX�NU��7��T���Q�'z�[6){�l�LY��$f���I�)\����O��첂�]:�c5ʎt|�˳�ve�)'�'��j�Y�b,C��GgE��{v'Kź#偱��3���c�w �t�F}ݹ� �6�h��氾h�{7���L���qƋ��������;"��c�m4˷`u2pS�	�i932^�$[(��53�؜U0���ZX���د�8p�N�
�?d��9�>y��b��ra	��`��`S��1�gPvɮJ8�T">����x�Ҷ>�~�U����Y���	���mzU�!@Ru���~���O(r6�BF�d4�.vB��O�yU���Z�0~x��Ѧ7U;�+�]�b'$���Q������7�������!�}3N�T��Q �s$Mj�cܰQn�G���6�i�By��i`�r
�k&ԓn@^�!O�N͍�*�[��S�ʕ���D��=S����W#��Q�r+z��Q�(X�����u$�B�%v��O��j�ޛ�;����A�!S2�ӊ#8DTYŘ�rr�]+��l�'��D$.��Cgd�+��(&��M��~�����C'9�0�h\�G��J����g3T�>F�M��6o��wt�X@i�i;D\Eu̧�J՛��xm�a������Y�sß�<��9����l����9�*(C_�;��bz,Q$������"�;�?�S3�J�|�\;�O�3	Ǐ�J�&���b��ރL�J+�[H����ؠ����Q�L��8��,1J�� !Ngo!2�9�y�<������䰘�%]����=��BI�j�� LեJZhV6�N����T��Sj�`ۆ9Ґ����[�&%�ƀ4#�B\�a\��D�N-ȥ�1=�Ѥ(��03s�]��Տ*��w} �d5#���b#{$m?������=�źl;k�J�|;6��y����uu�Q���!�D�,��H_l�+�Y<�'ez\�j�����������Y��E0�q�ٸ�b��2-~���^5��y�m�)���?�����nI�:a>�D�!�[&*(�U�+�Qz;��d��(��-��J���ϸ)�=H3�� �x��H���Y�a �	A�Zx��]>��:�Y�#�f�ʚb�5�:�� �)!x<=rr�U���8������ .h����@8��T�Ol����k�cV�a��3Z��28K	M� �Qyh�w�z���%p���'x��M������eM������@�x�KiE���W���Mv"��Z56�� ��"�Mu�9�V�)��#��%���:@-rsZJF��_�T�,����m�-g�<a��|��y��\�{p�wrHL�e��U�k����DZ��;殉L\j.����!l�ގ6Z^�{�v��6�	HZ��.Ѯ�*���x��G��	�8?�\c�I ��MǙjP*�4}OBֱ� ���cfI<J2����Pp�~2y�ڦ~K���Z�t�x�PQ�#�?+3[���Nؗ Jw���<Ȩ�P��
҈:wp�ȟ�m�z�1i�nĕ�VB��!,x�����!��g2��[$6�p��\p�шdK��c�Nx���"ľ�LL,�1@�&;O�.�k.��ޘ�:[��_ˠ�,{Z6�j[}YR�d${���m�
b"�hT���W������[�T��3W]Ck�(�vϜ�yh�ۼ�c��w)���6zC�6J�n�vGg��z�)k�;OӪň�/O^����0u���Cu�8�«iI���<vהgn���3��GJ[�5n����=��s�_&�
8�=U�:�p|�7b�gHA�z~Dl�KQ�%�=鹐�S&�7�t�R�o��:Y0��Q{u�mm )_@I��u T���b�{3�X�0|�K3�BX�3�"Z'�vU��ԍ7
�����C�,���QF��uk1�`KK'�Cw6.QCmIpI�ɆyEz��Wm��bIG:�p!UI|=k��D1����"Ɨ2�A/L+^�7ɧ6�:����J��a^�U����}S 'I���y<&��8^�ϣM��@�s"�"p����Ra��?�%M*�>� A�S���G��T�%�;FjV�ǨU�W�m�o��{�6��#�m��ػ ;��>@����=<{$����;>!���<	�w�[�o �s����hP��ߘ� �,k�{9TE���R>I�_�\�p_�^�������R�]�u{1���7ט5�I�k�#�^]T���ڹ
�ni��*P��:|�� M�l���Z�n���suh!b2�@�B��≗׹�����B�{sh�M��q�C9�>Zd���T���������~�u��}��ޡ���- �#U��p�:��^��W�*i���v���.z�����1�����
C����� �7���3�2*�<�i{c:\�~�ߢKd�1G�]��'f�}�b;݉dQ� uwQ�ґIX�P!��KzX��YZ���ɩ�[貙G�=�A�x4".1�F��C�^V�d.LI�R�P�|-gge%#=ڄ���,��F���8�q�z�߫��	�ڝ��6H�1wP��)W\2������R٭����>������������s�TR�L-�3�2�Ւ8��=�Cgo��sa��%1��D�Q{:�+Ժi�i�3)��/\��d �9�8��G������i�7N��;P�������m}ۀ���'�̝�X)4��x|���+ĕ��{}���a���;}{
a��M�x���r&k����nMQ��,U�B.(�F�#�?i�v����r���%!���\Ė���Z���b� �%�~�O}Eܙ���+G?�A�IJ4��C�ۅLjh^�W��IvHi����.*����������+M�ˆ8� )����n]u�l�XC};\���`��+���*T���|��k.��=QP'1��3�ˏ�h4�x��rU���h���z�'�-�)�@a�6dP�u������$s �u3H �o҄��z��-���(ا��H%5��SK�^���u��Rw�7
o��JX@6�z�_��7K��V���o?O�	$T!<���
 �tk�<�-������!�7r0�O�@\(�	���c��,��t�v!� bq�	���!-���H!�t��܉슉��#�k�0�M[�Nf�-�\���_i�dG\�'�H8��c��_J�S�.&^�� �e�c1�o��>m[���2b>W<��mzIcxbT��+�rp @�G�K��Ѕ|8z&!�V�pXC�]��?�X� ��3�	���<;��E4���+�9h8�݉�A[{e���k��a1�&Gg-��+��������������G��er��W0����&}��i}�N"<�P�I�~fG;�,�*Fm)E4vG�_��ne�4�K��Rbal�w�(��p�c&�
pX��@alH��"�ܮ[3��� c�,<0;�5O� 4x���.�#�2�`u8[�>I�d�$k���T	g c޴5Ku��#)6�ƗoX�S=�;��[��w�֢��R�H������QN��g���8+���R��1�G��-[rQ!����}�.°�G,��m�H���\�]\ybo�VK�hd��)�uO��_�;�����
7˯�	s_��tol�g��F�毺v��.�4���gi:C��l��{E`.��� ���P.�Sڌ��}"[��jv^�3?c�>��r!fG�y�&zln� O�/O<��5F�j�T��ݪg۰�*C��������&90o@�3��M2�y����bIcʞ������f�Z��_$�38�6�¼��&fc��ѧ@C���B�@f�`��]�Ycqd=�	X>*n�&?ԭ?�<AR�x�O7S�����B��7*f����b/&�gz���ǄĆ�D�B]�ud����w��F m��z�,YO��2������]6?4����n�����OGi�șr��Q��$��焑�t����k�GJ�!�ծ��3P@	x�!�"o
F��-D(�E��xkn��6��p���X�N\K�QUWS�?�����,�Qo��2��h�M\1�I@�H�[8�8a�L%�i
�kKe����� �g�#����ʎ�z,L�B�H��49C�:|�d=�����'5^�o�I����4�-}��Y֭>_U�xB!�����
=��
q8�S9�&���Ľ����w�ɻ� B�x�8�M^بՔ#W9�(B>B�i�c�w4f���0&��eP6[��8�F
�z�5�!�-�Q�Wϓ��+�,����,����3b"%�^^駘&�O���*eFg���� K��)~50ߤ@EER�⿻�'N`P¤Y��yzX��4f�`2���%�� ��D.q5��i�HQ&�z,da�)���'[�v{<7����AM&�`�)��F��dՂ<N@��V�½���Xߵ�m8�踲�-��vo��T�� K��}I�����0��](Q
Ex wߍG��:��2��B?C�ņ�p������q���y�ś�K#X�j��������yÐ�����RT���(Id�AȦ���+���}��)[��;�Tҽ� DσH�@�Ϛ����Y�^(�<��'3�*�M��S}+EE�U\��X�F%���#r���܌O7�Fc$���9
ofY�?��j�(�3�ض习��9�������h����nׯ]'3�x�HL�
�O�0y�r���YVZ.e�[�?�k]�X�o$gˁQV:^uc��&.� �� ��Y�EpF#A�U�m��.��T��=nV��؛�Q��WI��c��u^�w�d�i\?�r��[@�?�ؐ��U>$�	E�e�G�kq�{N���͋�ӁF:�`�5�����@�f��4."�ط�ƙhX�Ǖ6d�Q��cU���Nn1 ��_�:Q�T{n��Q�|��be~KL $8���H�+�o��_l++�m^1(���$7Oi��ncB��[�XP/�Mz r �
o�� 	h����o���w���)�	S_`��,;�hB����Pb�b��>�#�|����]�<e+ēg�E+Q�\���r�/�y�)�̊+�|(6`����ݿ\[���/���Ȱ�VA��wi�aj���ǿp�`~��4�ب����	#���(��X�/��<d~����%Qt��J�����yY�e��뗷��?��cs*��!�(|�(�iL��a���/F��$�S��Q�
/M!$j�Y8��u��|930���\�y�,ق|_.��Jq'Xt�x�&rd�����`��f������k����D�o~=ȴ��%��(,��u���aH��g�����̱��Gq���ǂo%�$�[�r�"��\�H�2a�YOw��S���Q��i0V%�KvCPMݧ&M,ú�EFSk3�H(��L����'y`=FMMu�h1���2��}nZ�`��$�X��Gݓ�}��)3jϷj�ѣ~^RW�:�h��
��G�~�>�8�m)a^Q��,_#ΉN��nX?��ƅ�8x���`RKS�+�0�% �G�TkIA.�F*l�cĐ�)i}��r YԪf�B�&f����7������R�*L���Ѐ1�.�ʆ���C�i�<����fo��ɪw+`lg�ZQ�Oi�M�Ʈ�2Oy<_zT��y���􉍬66��oB�gG�� .T/����K,ղGr6x��g��G��-~GP�T`-LҕKy�_l���	iN�x`�b�_�~��5��M~a��ځ��~���^y�є��
����ӏ=��<py_k=-��_yg3M����ٸ��u���bd�6qS#���&��6���f��1��c_Eh�}Vo�r� ��o/�)7�[sZ�?�*�z8r�1TC{k��V23E����G��ɢ���<�7��yX$8�Љ�.�I�X]�ϔ��`T��g�"��nH_��S���G����VO6��^��êWˏ�k�Y��_���]þ��!�DP�L�Aǆ�����q�New�u^��c7�*TI8j�	�s�qLz�f}�c� By����/���x�2N�$mf�+w}�܄s~��x��֕؍�D6�G+_�q�og8�j^
�.T��������a\p� �m�c��`y<z^�\�+��V#�%dA�؄�_��?7J�͙�A@DĔr�r��=9Fr)��yع=��]52J�u�}�S�	��q��ߝD�
�,��9
1�fO�XV�Ex���i�Ӣ���q1L��'�� ��T�|��K�D�F�B����k�G8�~e�L�9O��u(�j|����_L����b��	�$�7���zz�j %t2Jk>�=��w�m�����ŏ�>褑��O�&Rs� �zZIc�)T����.�Ԩ3��8���z���˝v�!�0����^�QF^OV%�u�wv�@&�37D��{�����;T0�������ȡ߯㘪av���o��\S�|Hzn��6���=� �RyKs)�.t���嘈�B�;�|��Ȏ�Q�'�|�+@v�/κp�)\K�P:��h�!B%y������4e%�c싇.۳WE|�������B��<
ȅ�p˙:��t���&`���|Y�r[V�8���:< Ko�7��F�G�kF#�m����4��E���-���(P�����(hVp�(��F�l^P��.�Ad.��q���� QT���aqZ��T����Y��*%s�;b����5'�=[�^6n���wJ;	�f7�A���B����;�.��8n��+�2�
2mۆ�ӯ�����zH��/z��
X�u��3�4�r;A3[8�f��m!�c����խ�	�۷�YV�ysQ����Ob`�O~�l�6�}F������֭�..5�'��',���X�>'pI��8<��w�~�!�S��Ƣ턔=
�V�)�|�[��/��*w�3�I�T�'CPۥ�e�d���w���8�����).'���itEI$���u-�P��P�L�
�G�cd�"��z�ko �d��:Y��%6GM�d����"��t"����@:�Th�K�q�7W ��m�s=���
�$+�`m+4��$&YԘ�ٌ��lG����N{S�=qF���\D�CNun���c���Pa�s�>��;�na,�ؽ�������-ׅF?�uP�V��җ�K ���y��@�[鷸ͯd!���<Y��'c�/F*/z��%�e|!p�x?�0j��������?g�^��T�Y?1������ߩƑT6N�{�� >Ok`K:��jlm����]�[�ա}���[���α �T�|6����9c}'�~M�hhZ���� ��&�E	��ec]�F��5��7�� ʻ3��6����s4j3#���C�?��G���l����W��i��̃�g��5�S>5jY^/[l�i<�<	��M� �U�v�`��J�'�P�۴s��߅�5(g�{3�s�i����P���sO	 �kQE��u�+���s�ß�R�'<:���o]�x�,k3�EĎݨz W��k������z�F�Om	LpI�E4Vm���p3����t�Z��a����0t��D����N��t���˸�������}Y����N��Y_s��1�g�(�!y<���3��A���1��Gn��Hъ���^�٦�oC�=dK��q#Q�#��ܐ�����2�Z�}�s���W첨�َ�	�b-��o���\�1�P�ǍwAZ�����-�O���re�J�s3R�'!2}�)��0U�o9Z�FȦM�|�Z��*EG���s"⸂�[0/��C��SK��8�H�bXp�C�
`����c�������̼����/r�Û�nf����/����R�*�tp�l��	d#�(w�h{y�/����:�&=ͬ!u&���*0i��;��� .^;o<g{o��G�����9�A����EwR���%�Q��N��I�ĺV��BK��ܵLb������}�j�~��q.���1R�����ϸ;����
�L,H�����A��xu[$��qFB3 ���6B/�Ob1TƵ��0�.��f�^���F�S;��5qَ����{�pez�-�׋�[AI<�d�z`֑\-����{��l�A��U[^m����:F�B�s�l�����Zq� 'p�aLv��L=h���NY?.Z���8t�q�+��7�D��w���V����p��n�7������鴰x��{�U�
	���Vd�Eo�J����v�P���x���Z���N�#o���1��O9��G���1z}/����M��� R��D�l�dG~3���g�N���@�@���?��M,0�z����{K��,�����<��]����h孋WA[-��v�N�uH��^�<�Q���~isX�A��v{��\�fA�$��9�0˳��@��;�L�-�@rF�n)~E�ċ�<��#�pDO�*�{�$��ޕmryt;z�:��\��q�0a�})ɤ�K[�f�����B��@�V7W]Dj�B��~�W��d�ٮ���ݕ��W�������w��^�3�a:����uw]���l�t?L�\C�!���ͻN�Nh.�3������)�wgF�-Ⱥ�:���p���n��n�f����0��^aoh�3)k�@v��_TQ��%aj�j�Z��-���vC��?�XEju�� �����@%�7g�����!��H�z�Ϝcyf��Sb�%s��7k-r�*y��gm��>�sw��p����@�m���Q!��I��� ey0N@��m���m����d�A���y�ˠ�3]r���L��p��#�`ֺ�T�%(�N�qzw�
�1��`��jq0�%��j��w~C����<m��d����^�Q,uϦC����� �1��C�[��ՙ��pWR�_̽���j��V�u`�70q-OQ;'�O�I%�/������`&%Tk��%z��Nu��gD�۸hp�����r}6����@L�͡��
E�ax|9q��'k�OUGt ��#Y��xI�4R����G=��o/��ڤӒR�$#p�O$>OLQ��,���=���#p�d�&-p7�]����N���늅60O)?�O_����v�R���'~�X}!PD��7��^z��YZv���s�se6Q���S��B�D$�j�-rc�e�4E_X�L�;҈^��'��mq!gSL�����ͯ)�dtI��G ��`�N�K���|r��%^�GM�VQ�ŹNl�����Q�v��ƴ�b���\���ñ3��$�,c��_���L?߻P]�z��Z
�ݤ>�SLn���_v�6�B���h X�H�{��R�/�LU}{Y�
1��	�I�%3�@U�LL+���5Z���g��D��䁓��v
-3z+���r��ٲ����Z'DQ�6�{&m��	�BZWY!��s����n�_qި��J<E�&{���1��tK�����R;<�"m����t����E���܁��JF[�3v��JwYC1"���I8-�
��R�t��4�Eͱ8ˁ;\LC6����S���hU���%>QZfe�ڌ3��3�P��
3j	#Q��YR�pK$���}�[.�k0r7k�җ�{�k��6�͇z��k���'��N3F�"���D,��0G��}^I.�i�4.��h��Vb�wW&Y�1o"����AB�;�L+{<�yވC���*���~�b<��� �$ܱ8�[�:�8�Q&ش��C�1�Ӥ��6��z1�@J�+������(G��yG	�\��4������׸�p٥G��t�V7�� [�?Wo'�"͒j��{���'ez��t��n�������-c�Cޚ~ 7NAk�X��`�=�/u��?��X�牴�I>1�E�(-��.Vh��a5���qCJ�x �Ut���eji���8T;�V*��*�� ��8���WP|����Zp�mbZ�מ6�g��e�Y`+"��¿�S�)g��8u�����9�3�R%G�u�3Z���׫�w(uj?�����K�4��?u��m!9�zQ�������?\�=~J�_���\��G���7M$���
��|兆�Ѕ+ 10�狼w�����YƘ)�m���T�V�5������
�z�	�`��u��]:�#wi%�O�&~�^L:�<ݕ�)�r۰��
�8v�+����b�qW����K*9�P���N�˼#;\�dRk��{�D���4�&h.��]�I}r����-z�/\t�e#�	�:�c����f���_�vN�BB���0g\j��S��D)��$g���<�̲�7c}�x�c��,W\A6�|�:l�e�^�������*�Tdo+vj��y���\T��AU[[»l��U9�ɝqp���J{]1�V�S��t_i�z��ˎ'�2`�Tp�S٪�ï+�2:J���