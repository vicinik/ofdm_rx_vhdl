��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒���8���#��\yo8��^W���S�@���kg���Y�źA�����"�v�F�"\
P���DL�7(6͞KCDg�rJ�߁�x��zl�;�xi(��9�r��	��¥�q먮���e�t8�A�~�z�L�v������۫� �+n�+��B����V�'��U��QB����:?�
��q{�֭�c��*���ˌS�h<�ה�M򅿮��vm���)3ǉ%�ǝ�[O���(��yB��UY��5USs>�E��U�B
^�(gR�
�]����(��������2T��������Mա�m1�yp��q(���l%zr5eTY�!��������];O+�׹��Ȟ̛� k�a�o����P��\��î79b�9�P��ttI!oz=hִ�8v�F�9�s����U'�Z+��V���,u<I׽@K�T��܋�ɛ�z��ݴ��&�[��MBi�E��6�N���A�N!	����������X�
���� v��?���;;xZZ&d4Z] ��d4�)�E{.���VPޒ���r�.��$N�CzO�*�)4��1�;�{�8�)7I��<U<�A�>D�Z�4��X��K29���/������\��5�����p �n�;�wZX�Q�H����r���y.ђ�/N��|�>� "�j�t��3(,�?��O�������<��P���Mu�s�\�,�,9p�������Nn��8=�>����t'F��r�z�����E�(�|�:�T>�@��-��鶫�'�Tˁ�j�3��d��$����7�}%-�#�Sڐ��ILȺ�s��4��h��K$��MS��T���[�v=j�l�u������i�9�A��{�<'O7��Ս��`��{ k�|�� �i�{���M)��W������x8��rB�3
�p����N]Yq*��T��v1`TWyo��{T�$Rd���&W�;��ܸ���g�(�!��da [6l�QPHՇ�:�߀D
6;��i �!*�[��?�jb�?Z-��dq����xj�O��P��
g�Q��B���J�p�gE<B�*��P��r��� y�đօ�N���'F�$>~�YX%�����7u*-�Xk}̉����PE4]g=k̃���C���0]]��!�<�g����������1n�o�0*[�_3lwj-�0/_SCt��?O͘�/k�|>Y:h��^P	�Q��6 o1esYV2��<�2C.��%�Hl�d��w�Wh B|w[����C�y�J��]Z��,�����F� G�B�`����d��u�%C��1&�������)���/_qϷ��]��T	6�aG�/���!�c�C��	���5w�5u	��<��u�Q�HbB���6�'���%
|��+G�'\KV�j�˩\@����C�f�m{X�E����
.��@��oP�%kCRZ�e������򾺭��~�� M�A4�(�����XXͤ1�yX}�;�Mp�[_!�9�_{��]��je�^g���4I�����DDe#p��퓗�!@�u�Џ��N$�F�8��Y�
����xמ��2t��c�Rd7�`S1Џ@�� �Y�2vȜ�iY2yB��	i�ɺ��<i�ޥ^c��˪��p@�+'C�|yԹ~�^� =6�ʊBR��c��O�,����n	ɝ�F�
��c��/��H&�a�Uj�M'��Xt$�����-��_����T�	���ͅ��Cq��֦|�FG�l��t�*G2�D�c����px�B�2aK��t�	�3�W����{�	r�2
9f���I��V�w]⓮?���fB����ڜ�) �f�q21 ������ÔS������lzY�Q �wb��P���=�K�Md)(��c�;��#�f���������9";	G8�d�0��s�A��좛��)D,�^�|T�h���i=�"��B�Eݩx"̍���!a��Pv� ~<'2B�D�r�z=O��<��N����o�Q�B��o��54��Sr���۵�S/_:xŮJ�����J
��i�~���7�o�!��(&��+8>�T�\�]Y�Vչs��_"��H� aZ�� �{ͩ�8r��B#�#w/G 69�S����4�dF�E��5"�ê)�٦�I���/s�Z�%��>k���e��8\?>�h-�%�*i[�
�|~m.E�E��H���am��ZS�!z�H�Z:�A������5���{q���5�
�Q!�2&������m��c�:�7ec�ɸ)eݷLW'���GL�2�*_�t�!�M&$fO`��;i;��E���W���Vwց�L-�I:ސ���js��Yf����g�܋�o�@3ڿ~�%	9ZY	wL2�w70,a�b�G�d] ��D-�>��a��&�dƸ�K��yU���#ҩE���t�~SYo�~G����_����_��C��-F�,�R&��=�̤��S����Q�"��$ry[�ܬ�2�:kNJ���s~v,����$�z��ݜ�f}�X���`�-.=X�f��>SA�}Ey��p�J|Z�����`�Ph�,�O"NO�(�5<pW����!�-�%�x��(���E�z��)X:1���&}jgxr@��"��9��b���ӻS�}�˿��c���S,������>\L�n��M�k2 �+�1���_1d�r��љ'w��Ǧ�|��Kn�{��r �fL}1���jܯ�z�w����l���i�rR�-�
����g��V�%p������G��a~$<>�"������:P�Nڄ��KQF%���yЎ����	a�w�/��^��ySl�*�����ia�����K��t\{TD�]4A�"��oˀT:>�)���m��NtR��P��l����S�38A��9���ѡ�c��R�sҦ�D���u�vX�\W?rlv��v�g��=MB�:�a���ိŰ�=���κA��~��)c(���r�^��"�\`Be���^x?��k��*1v�[��0�,-_��g���d��<�!
�e]�1�������qc�Q^���[݇Iu%*9g��5H����>