��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��f�)C�� �P	�wǫ��dK��z�����
X�Q)��W�a���sgy����[	ky��F6�Ut���Y©���f��؞4�_�F��J: Ut|����f�y�J��a�}{�}{���Lc<��Mg'�0���#����2۷����a��is�!v�0E����R���	���oc/�6�XiƆDQ�'���=�>ی�����V��y"v�bF/�B��.��}\
F���� Y��� �2�سo���M	���n�z��mqC�(��i�6�`�I����#4O2�}����|�8���)�ie��vo�P޼�硱pbǶR�������iPB_� j�Ў����-Q5�	� ���4"I���x��d������(������b"�T�v��&��M$;x��<K;cDF�TN̫�.Ę�������ݝV��Q���Q����z�B[�n��5��*4���eU3H���~��4W���%��-� xR<���[�gBɽ�ѱ/9R�- l4P��Q2=�l���S�?,�b��"�v[7D��@�fsOU�%׼�-��c�����|��2�jȚ��[Fd���&~��R4&[<U�0�;r^�嵣���)�wρD�#k�1�fE
��@�LD���F�?- D��A�w-w0�'�*e%m"���q�M֒^ʊɔ�f�F�T��
����2�s	�Um����q��#gN�� �@����\f�ھ������G2#�gU$�5�5xeK1bk߿f��;��~��̠,�Y)z뫚�:I��C�o�s�;3IlU�S����@�4��%b1�j��s��M�Pk�b3��.�v�����ƴ�㽬$�pTux���HϮ�y���ϐf]�awa��G.7Q-2���Jt �c��g��/��p}A��G��}H��Z�e,J�	��û�l�K2{�/ �Χ$�m�c��`��'�VF_�r��#�9ɋg-�vU���[�At%�G����u�W
��>5����G�Ţ��$�6R��Y���el[N������>%��΁
U��ұ5��k���{�E"6�&��"�QOI������v�.QX��LL��p�ug����:�,�4�����6$��p3!n�d����\	�s���f�B��Ǳ�fn����-f�oz�;{��Q��~D��T���,.8a~�Ъ�"&�z=�M��_`~�xIʨjԅ����aoF�M��bœ;�dVjU�
�	b���Ԡ�H���p|S���;@�W(9L��X��5�Ѳ0&�.��3ܠH_�9lT{E��|C�u��v�3f�-50
�7�k�:%`��m�
� z�VA��A��	�ʫ-��ٍ��}sMC(�����۽(Ų��`X���h[2~���X��_���]el�v]�9JS�Gx���]|�a�Wkl�8�U����RL-�?QN������+�b� �(084�^]a�!�>��X2=Q<m�5iD������
�����fTjO��PKf�9�/A��C��V�����`�Z1n\^S����I�l�5>X`�s(�
�J�:��͍i��*W�2YjM���n�4�9ױq�����x���ߍ�|夞x�D��o"�by�W�uB����[*�OߊrY��_��Ѭ�M}��+x����-:����?��QFr&H-��l��Wd���DD[�j-�uP��u�R��{��M�;�xDy�!��qp�LBY3q�{��Qi/�����rNz�c�O�":���ఞ�G+�),P!��<!��������s �r�R;m���~���Ě���8��J��G\�m�c����\�%x��y� �&a>��	{Qz�L*���in+�X\��X���<d{ڝBfRt���h1��Ǵ^������b9����b�vŖ��Ajϩ6|�nʐ����o��@��a�~���t�r�TP ��&���ڽ��;gEҁ�x�D�Y�J,�.�I��ifub=����H����_��p���t���p�Ӱ�$��GSU����t�Q;�d�4�Nu�/V�gͰkt�y��%��m�Ll�[�.�+S%O{(��WK %�@K<�Z���f���I=�`�����N��q��'T����$cW��z�F1�s8�*M	&OZ%h~�yp�9l��!~��rC 99]�L*=em��p%L��}!q����$]ocT�w ��[^�"�z\6�~��m��qp��S��'q�w\I��J.�;ۂ���Gi%V��Bg)O�������@qE/�j���J�C�lҳvK�2�r��[�Hɘ������c��M���:�X��cX�P�n���u�%s��%�]*�{o;f���P4��.l�L^��	b�&ι�>�LfDȾ�st��9+Z��/X��@�-N���I=utn_�\="'�ό�kw`��A~����ջ�TV��<���B\�9:���]��-zEЊ�9�B�O2����z�2��?	<�<&ߏ�8`o��w��O�����X�E��<�� ����	P�UZ���6��t��I�|\w	<��^���yЌ�=p�J�:-�����
�z���HN�8lg��yYR(�����B����݅@�ѩdd�ԑ�@�:�:'����M����$f�i�}Ζb�l<��.izu�
��V�3�ڪ���H�%ja�)�BF�L���%6(�K�rʨz'.�b<Z�Q����2���K�jM
:�N�I�﬙��0b`��@�f��1��{/���4R�S A��[wҷ�������8�e�*>������wnrɘ�Us�0�O�}x+� �={8d�R����&Ni�����j�"2m�y��e$�����v�g�*ش��['�$ ��άl���յ>��Ixf�=؂a9��̭����a��-{+��'t s��r�9���
�?��0*�֬Z��<��̎?�wA���2�����Ͱ]��m�F�e�t�p�<���Dj�f����������|�~�A��L�<\�_��R��~�UEfN�U��[P���7��Yf6��@��> ��o�Oy=p���y�en�!����E�]���'E��]4��C,7���Y5�VCe����7[F5c�S!�݊���)�hc�'�Ӱ+ȑn�?���e��V�a�^&��A8�|�׽�z�v������m�$^��c���`�Po}���0FU�mZ͉"��2���W�+���؇����H8�Xuh`����\J�Z���Դ�c��N[��zޝ��d�S�n�Ԣ�?e@��.�j�5Ē�/�X�@.�h��ar�}>08��|�9��"pH�`��8IT�yl��x�d��&�[��FR���Ƌ���&IZ�R�[z��9~Uݍ�#�tvy�
�l(����Q�=gmn5{R^�%s�U&ܴ��I���}FC�A�׽��o���n����e��U��Ue�2�m_�4��;�
z�����QQ�/�Xxݍf/F,�g������j���t��񮕷��a7a����@��S=t,��XE-����)� f���WX������}�P���[��Zhk�
��aĊ?�%|!8�Ӣ�hq��kbJ�=�v>@k��ɖ
j����,�qq[�T9?������iU���V����� ��5$��������.M�����v�󼗝��O�l�Se�FZɁ��)�s6(ਞ�EOu-��`�E<�l���<�@r"�i4X��i�an��nR�O���[V�2�M��=i��	��C��@�n �y�Y��'���&.�Q/��O��RB@<���`qi�� T�0Gv�g@+��S�_	Q�T'w;$�x�:YF�ҫ�[�cY����s�9҇�3Y�N�����gs,=�3�cO���M9�	���pW���h�,e�9h��4xF�����e�I�q�ݶ0y�K<t@)���/̔�\/f�n��ʵU�+�ٕ�wH�N[��)�����m���57!k���V��V�ĶxT&�:Ҡ"��,���VR��v��3��'/M��P��\g�9�t?4�����#�{��&��K/�q���P���}_�FJ��A�٘-����`���j{)���|	�	�j Bm��kdjB�a�[�ָV(����?���FU"�
�3����(�ɱ�l#	-��Ȓ�D� �6j�B	n�W�rF���t���%�'�� �����3\�s���3�;���[��q��s�V�Yr��6_@�o�A�B*��%f�d�E�%�ӅX��&/�[�P��$*j	��C����Q<s����1��@�{�P_�6	� +ًE<�0:b~.�zځ?ǙuϦ���Y]�z���ݼrǂ������K��.��G�&�CB���z����8���~u��|v�am�_wG��A���c�) ��,'n������+���J���.�&wǷ^¾��Z �6&S���!��
A� ����G���v`�SS�*ݓl��:!!����?���ǮG=D�ɵzc�VGCˎ�[JxG&�@�wQ���1�១�8��"�.B��u����/;���m:��\I��h� �$��]�?Sb��ovb���f�ŕ�M%w�~[�/��UU���DJ'���5��&�fhC���k��{�zqW��j��e"D�^� Q��d��j�=M�$֤�	�O��/os��P���?��K��v(�g@��dkd�A �*(������-3�2F��'�5#��k
V��6��!R�`�>�T�;�s<ˁ��5��d'Jkm�SR�8 �#3J�+�
��q�?)�@(��k��~#�-����E�*B̓C2�Rq����s
@��8���DS��K�a��X����L������\U4X�f]@ݫ��ϊ���>��ŉ��o<G ZN.���6�N�129W�jS�IJ�<k$`��ݩ:��z;,6B�b?��b����M�a�G��c��L�\����P1�b�%Ǽ��P��8� ��5C�������M�5ڄ7bf��BB�{Y�7�s�j݈L��g2#*���e�����gk0��sBB�P)�d�sY<�	�{?7<�t^;�)��3�qK���D{0?.���kB�U��xhM��)����s��Ќ6�7lq^`�����8�e!ȵ����/��������������� �t��PF}��s�'��xy��قBc��R���_��Wc]n�C;�$�$��VQ#M~��M� �2a��1T`����2�+�n�%��s[���fm��~���j{m�J{��G��uM�7��ǋ����(�S�zXKs��0���+|�22
?��V���L'�c�2�r|r��5:�q�?��;-�Ox���gA���I��Y�3���#��D�nC
U�m?�e��U� �Ϡ�����|��sm�m\`���N���N�q� Sh⧝�S'7n�]e9 3���������E�� ��(�����n+��Z�/;p��xܜ$�����Y_��͝�߈�XLHb����M%5� KXm�j���A��)�|�Fd��X�=������`�~6�S#_��ßU�!���zBp�d�Y�M>^���|��h�7g�Ծk��S��YE�-�(�*5�Ϯ3W@�^��Yc��	�����$K捻�c̳��9k۸u��Q�0��H����64-SS��};\���串�>�[��xo�#�Z����{4�Cm��%���-�4�
}S te1�q$�OG*x݈�G{�EN��X�"�G���r�y�1��| ё΅#�{�iL��n�@l[K��Fu��t^FTL�:wK�/�W�
]�4&�F��+�kp-��kf4��ڂ�	=����o�x�
=���Ŀ�ܕ�F��8���A��Fb�^�z���,�ב���Ф�W����p�u�:��i�MJ,A�*�$W���Oa{~�lSc����@e	Ea�,�	a��G�u�I	�����D�ġ�		q3c��0��낣o�pd�%���l.Q�}<��˼�/SA$�J �]��֧�Mуo����M��/�r�Z�zXFkPPW'���T�.�Х�c�����dk-��b���
�4	G�\��ԯ��2K�3��(��.�O��i^aj4��`���R+`%�wMYhv"Qi������%�������-Ă��v���7���#~K0?ދ��7ŏ�x��{���ϥΧ7r�til�?R��[ӯp_ <%>�qN6A=LD�_;gJ��p\��P�*�@�h_�U�]z�V�ޞ��Ǒ���z}T�Z�&�P�������5�ǰ�{O1\�s���Wt���.�$�'��D�O�p���Ї�a�1%B�d�g����j�8W��c\A˼�$�q�WR�ܳ���{���Z��]�M&�oI�\m{�K��,�[X�^Z���eQ���1���wz�62�Yq��>"��Vq�k��^��U��S��ޔ|v�3eV�pC�u4r�5 �6P�_i~�n=ī�/��Q��S�
 0�*����x��Ѯ^"wRǣ���@�ud~�I��J���*�SM�N��A���I����#�Eh���g2�2c��Ju�o�*�KZ��
��&�~%���t��6������NkÛ*?�Af�~��!ߘ��˓:9>������HR.�wF���7
��p��W0��#�1�T��l�CÙ+§-��,��9��aށ�	�U&�s	N�P�L����`���Am*g]����˨��
lR��?���b�J�.K,��
;��z��FRKk���ә��AE�}D��B�d�#X�����Ai�bLґQ�.tg�3�2M>d1�Oqϟ��(��Α��j�+�%JQ�7Z���LU��|C �J��/��r�/H�.?z���[}�z�E�J�@A��u��'D��)�V1�Ɍ��iw���hNYB�y�:��H�� 3xAB�5�p���q��aT�W�kK;�BT����4m8�*��1x���������h4Q4y+D׬��*}��p�٭?��63��q��w�1D���~��-`�Y�����7>�{��a�e�����(�E�6�[EE�;���ϐpǐe��F{�u��10���(8�� �1������ܖF'���F��`�u��7��_�4 JX����J�R��X�G�l�P�}dZ����@"k���I*�5h�
�YW�GՐ�}���a�+���|��ac���uD��te�5$>j�������Ã;�<��(D�A�j��DPr06p����k�6�c�7�	T*�ϲ�&�(J���z�iv^W�E�P��#r�@����gW�XW��/�ܖ�*N@���W�z��D
��f�
e]��LF��V>LC �i��`W�{-Z���j��B�p�4LZ��9Q�w�m!���O�;�4?�n�?JH���IE{x04o"
��_��7q�H.	�2�rs8�i��g�߳BT�9M�'�4"�ps�d,�8�PV�S��lak�}�uU��U�q�� ��Y�E�t3!����f�a;}�荌���&o�D@'흪�3�e��A�;ޜ���g8x)+�7�_RU���>�gE�\{uzP���@�qu�Fu�nb�J����My;���������C��kú�����}V���=�.�OC�Nqwq�����/����3��pT�f~�2a �O��5)��~P*�D'�74S�n�P멏�uiQ��G d
}���?����#2^�F������j�zޠ�9r��]�����5�\y������s�AgoY*k�Bz�gx�_�M�ulF"�F�^S;����^il�vj����O�<�٭O^�tD�?\���0h�0�F
!���KF1��0˺h5�J��_���x���],z�9�x>Q����c��-ฆyb9Z�X�SW�����N�R�8�
�ݫ�Ƙ��y���x�J�����M���c��
��ř�o����F͇E �ѾY�u��`�ٛ��9��-��?>P��:0Nu�X��2��s-�B��D<q�f�*j]�����k�3&>kñ;k�m}��}����?�\l��:����^$z�Lo,9-s���v��AS.����oL2�}�D�l�Ь뗽�9�;K� ��r�O�_����쾥�ַT���E��!y���	��4}���h���&�}����|�ZlmY��h��A[	J�����t��"熹!e��9�-����=2C���QܣT�_ئ0��lp�b�ԥ�գ�c=^�hPEJ�e�>�9Bb�j�:�阪��Ж��,��H����q(&���"�%��[膘�֪������aV��5��bT|��B�M�ln���RL��2 c�T�N2-LUx�E�����u�NMz�CO���_� ��[;��*%�[2��*;�U�f��RrtNA�{�}�sw��k�}|2�-4jDcB�9:̰r,�+��N�� �ؿ<���ɸ���o��\��O��Go�k�oǼ.�$� b�9>s��(�.��yR��!.WW�A˕/D��[[�)��r=m������cK�X�rW��4
�4�#�>�8۽7��D�o��@w�$�F�W���w��%����B5���[��Q���H���oI�'�/ngeZ*VQ:�������zU8�+�x�����D:S�t�ٯ��l*�(�;kɔ�㦮�!'�
O+�u����.�Ы�aJ��"�|�ʟf��јԞ�i�gy}u\E�ZL��G�����6�7~��eZH�3�������ʌ|�}ݛ�jf��x�R��b��+(������A�&�jn�ФR�j�w���zޱ^*������N�65[5/��@�)Z6&��Ԍ'Xe�xn�����N	v��9J�2f�c��1UA�y�l�@ð�@���P8A���L�%G:���q�h>Ծ�AZr��6#{'����}
X�����.	|�P^,�~�]��Y�a�am�ި9�Ū�����6�I��-�]H�31��̹�\<�9���SV����׷&!�>�>) � ��Ӟ%T��v�)���]q!�^m�_{4o�:)�!��]�K��{�����2��
CR�A�sZBc�\�R����KK�1��ْ��^xG��wϹ6�ќӝ4���"
����NjO2���Ȱ{y|�X�E�l�����.�PfVQ.s�	:�M�$S�7@$�2�,[�hи�Y�T�r�>Զ���N��~s �c�v���]nуPC%�[�P���-3h��v�x���V�T��o�cwz%?M|d< h%�ƞ�^z.R�ӹ�a5�>Mw}r���U%�B�v0�DR�bm�;S	]����W�rX��ݓ��>"���2���Ge�p8hS����=�LBO�L7��G��\9Cdr�
��Zj|�g�K��wO�����n���9�";'3Q�8!����KTrJuH�/�/����C���r@�-fL�k�' ��
wd�9�9��=N��I
���	��BS�i��p�pe�z����[�L>���l͐��T?�,�3�����{a�����ќ��9�h�/����k1��c�~����Û�T�F��
I!�Z,�̸m�u0A#�v+$Q���Z�ju�+a�r�C�>�}^�i�E'�Ӈd<f)3�e��>q-z�k��������Q�#?�g��0&�n�s�iӠ��Q�/&�:@�#���&E!�`�-P	:�dd8-�Ů6�
@��#`9�f�I������If�h����xOjF�`��D�_�l"A����k?������Q��r��?T34Ei2зlh��l�ϭ�'O����,
@��ݻ=�/�Hf�	��ʕh9����i8?����y/�Q���Z�}�מ������`~�(p�bU����z;₣��Űԓy�n\_\��/q����f!��l�X.]�H<�T)tk�vK����틹���p ���L`aL~��!GaB)>%��xs�ǒ06(~W�����8�rU�Z�Bj���ة���e4���jM5��lӣ	4,��-�t��w����NG�3��QYe��ߘ5��w�Q��V"�x�6�"��-v���b�_;�s{��
�^k��{�1�/��x��ŜL{g�kS�x��=�D�)���`�`���K+��T�,E#��f�$^�U�>�.�����9�1z�o(�:�#����1��FCD���� 5���� z�+���)�^�x���W(a���l�-�s�j:�olUg����rZ���)�a��*� E)��nG�{'�!vF|�׽)�zT�/�)P�ae�4T�B7u7��ߝ��r����)Gl�֙�m���뚭�^�0��l�B�ss����პ.�/�tb �����óN�W�̄���`1MHP����ܫ|r�˥�y��S+�@��n;,B}��	[�w��S��3V�h����1�e�
�Y��i��f�o��( 2�Q7��f��<b����L���������3�\��}��k��ϼ�-�On�^ӀŅ�}����P5��>lG���t��.LV�{��[������i����Ufo��ϱ���:v��D�fRE�����ELۥ��4�K �Y�/�Gb��/?� ����1
�����x9���}�]!���k��\|����nG/΂���i�,�3nЀM���+��S���|�"]r
�{o�}d�U	M�9rtѿ���5Td~A��4����7�]����������	j�%� 1-����a�A�R�H�X�`�� �P/C��d�y����⯵{�~��q�\�	�,Y��O��w�M��fT��2��.������4R��k����N<S�`��>�{cT�<ь�L�J���1���Β�M�i��AHZ�* �O�v__���d�A]ڪ�*��p `hKO����Us/1�[mD�� t[��{�%8�ZM-O6�Wv���cE�l#�G8V�{���X{�B(�A�2��