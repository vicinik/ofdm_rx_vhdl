-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YD1nSxjzbwdozrO1/v9vbje8NkNCcsA4/ddo0gKrWeEdx44YacQZmFYRayALKAnP//EAQVQO22/G
g/952hMrFyWtO/sGWESOHPW295crCmJRYG8jJlh2lsi3fpOG0g/KqvyCHUqPhhZA+uc1+2UjYzgO
CIuJZVdDNPHiVj3HlHg/CwC7/N+p5Mh+bMaUoSN56T37pIxhYndlsCGbnNFOH8QAJQHsIiYmZzxu
TmHcLMSaGo3WJkT4Yva2LUdWa8gBLI/33OPfZi9BNOEob6NE22Q1DhOkCLv8PVBmYkqFMWyMHa48
5sDIveGXYCKCB8grNs0YwOdJBaX6xGj0xqRgwg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37584)
`protect data_block
1oShSmfraj2yItYe9eZ4tL7XxPHwqilsGujbXUObS4+PsiTra+zRH1ERvOMbAC4hYRO/ow9uHezo
zK13Gd+h50FUm2ghQnJr1sG1YCn7FIiJGsUVFHtaq8dP6/JhRTB1h9tNO5+rgIuvcS+Hn8pYx9wH
4WPhVmngPCSIbvQG6u155pppzlDx3GLDBnC+7DPjYG5FyY5bMi+/nqw5qriecDOhrlVt3FQGpCMm
X4DYAz+dn6s+aqRaZ6NkR8KuBZ4cCxCVkzu9AwPlMhi6u3+AoBHGuYLFcukTPEjnLAxPF8NYMSFY
mq/5NNzaqRaJ2pW9Odwb5bzjQrHDAVKd12h0djPX8bRw5ujXXutcJMrktQNWgxY5Un4E8DmB2XOT
4nPljYAfKM39xEQzMsA6yMTp2Ttzylx2VM5ioWphEKH1xlVefG6wrPlPbd95e2ju72nh6sVoUiZZ
aNQPfS+HJpjfAeP0GCIWOT1tfNH2jAB2fKtm1DYdlZYTlxi5O/OKVkovBMRDn9tvauMtQgQyuShl
GCFQkMM+hM22Jd+g17AypQNNwo4c0AvOqoTaI6IvM1NHGAnwTOoCADvHi2xRCShrYeBv00IIUz1+
+d4d0UHQaHklijWq3SgeYECwSEZYoDmbhqZj3blAdDaQy9clGVD0cmw+/qfJbWIzUYXG/0lOB+Td
vYRnTAqdS3mxcd8OYVSgMVFizrFhxxxWmyBj1/MUaHJaeEsUw4wJn0sLJmpM1eQW9mxznP28lQAC
VMLxVqhaMNLlGP05TK2KxMmv4pqE2AqN4AbfURz///XRjg+Vw0i9lj02ebpxAuD5DnulTvqp2zVY
LCBenLI9EHpousGRypzAfFRw2H7I0+htIuUsaLkL8zOGNCg68BSb1sNSwWf4kHeE9lRCpyTRGn1J
MJwtL2xUVuAeCbMfhUPlCrHu9GrQknyjWRVvdMR+y3EjbVm+J0YqtLy0bj00fOHLa3h7FvRT2E3q
pdTKgi5zfJ5wPJLHy+NKLenUuZ0UyVwdOCGa4s+NXuAf5ulRgec7yyIAzYeBGgm6OAFfeBAeER4s
phEcub6H0LnARsq7komq4lLDVChJ5pZpKr/eMqZW3ubpNe/lcTHSwKtXXFdKDs0cy2cED/HRQbGH
qPxlcIjDprOY5/4N/gwHhJyDiT33FtJO0fsRHIYs7iJgoi/9Ft1GALMWcvLqWNn4rWvFQRLEC2p/
ewONsy/GemzDdXzDDZH0f/hp4TvrLCjC9O58HKrT7XLyhnSlQqFXXNCJa+abVcRCFLwqVzuOk2XV
TfTFh1SBZxWn6yux3vkHAOkX4VBOYxxYI7uv9rnJseeoeQVm9ITuLwbCnTmSBq8i0LYUi7/6YxTW
C3OVpi5XtwvdwLhvAoJF/+gK6WibC6jcM0oe7lODLsDogmfh6ChZW8wUH7E/RFqbkXJS3O+XaNQq
bKcMY0GAqEfRziXxd0zpNo7NVf66lLnwveXZQ98pkmK4jeL1RvtkXUpIyGOPMq/JlxghK0jmycVZ
jLY4uKhZOIsW+XXRga0AzYDOdTKM6hypLvDgWcWIpxjekoNzQG+vJnE1vyBAOYGo+9PFm4iZJq/1
2THCtPTGx5UcM+crYtrqWowSOAyYhNDR/SMjAJIRdG+fGc3E09Z/0yNRTnVIX/SpW6bp1/ZyimgG
64n3f3xtNqwFdAAS8SJwlQx8K5DqtwWmsjHq1UiCXjImz8/HRzusVBlImKS/n9HMlwQ1iL11XU/k
BcSQ+okNHJSy1JcU6tc4DSNIskXSoeKStvy+i6wFnZGEFWDcApQ0GFHomJUkNh6PQW1JDhVYYD9w
FZM41jGtF2YsYPWu6JwgL9pFuhLfJra6MgjBFgsjquKgKSS8YOFQzHjoskN763PhsF7nzVn+hFz0
OhNk7PqMbfzzBzX0xoXnIiauylO+SmXwuzdLIoqmh0hqujtoX4NWeoYMjQBAhDdUBikJhzvP3k7V
5pAoIT66YZimwBxks6ryHHRtmb8vugs5UT4P4HplJjm4bFDF/y8g0dhqCPRClytgFz163vb7QuxP
scLEnZrCAimP6XuvuxRupu+D9rEBSiTXa4LdbfAQbLJNKSSbO8RBfv2nFXKYiOoNIc6+U1RFrNz2
OYvxCmVufa/ZVxGU9lCenOkPtz5DUTn5Lk8921sYokveL/j5TfiRdhJK5Pe7TvYfo54IwoWaW6HG
vbHABXD7xZuv3MGxPnQ7fWI+dTWHMMng59ec4OUxT+rQMYtn3lthLH6q22UJxNP8FL5GDCeMJs4H
O5G2pcxJ8KR0Az/yTJVP/rKGZEWgUonPhk2eSpJfXjbts/5xEVklfR9rRMW/8nCICk67WhTWg8TH
BnnYyvBLj8BKiE9dIw7pZbMjGkl2i/1GVNTvQvjz5EaVTxN3ruynC8LLqEZEsvd3o1XIuvo4sTno
YZecEh2QCCxNMPrN4ql+yxhxfmtMy+ijafxY5NPzwrti53Vbscrf6Gl/h7VktCLy+498gCahf1rg
IegpYIEvKBimjZkTKhfsg4y1Yzw4EIO6C5anYJzdwH5soen2n1ylkqRgXox1CV4MFnS20Dz5YwbU
xwWiBw1Aoq0m6Tlx9w4Wbge4RK+UEMkg6dSPuGF4Qrnbkesvo4/TxkyOo8DA/smQ91nzhqQ5MxNH
DU2qAKPfx3TkC1oTc178S22C4An73rLd1vtZK+Qs7kkRbSqJy5cDMnsLbAVFaut9lVU2ZM3wjS3r
V/eslvRzKZFloJnBemspCFdeUrkjm94KJqHzJIyRc7iYx/dnp/1gYKu3chazdF2B9WWkaMTATS3n
Jq2UlnYjQGA8m+yocvCbWuuA5M44MKiH+SSbuo/0qQ0syq98BUQeEog659yLiKnH8r/4h979xUeh
sWrCu1NJDkO8FgWJNSdqnURlByIjSHn3MHIm9WF680pj41kf0p9ll2TLs/TEfZ/sZT12d2FA5Vto
9Ku9PH4jLA5i1mHfE/Pi44kJVtlxPp5xzkfsLSIsIQgLj+CVnkYNrn9Lpmu9m/cVf40M7spH0NIj
c7rjGA8vfGva4lQy6KdOco2gHf2HY3grcUtuZynl7Zmu7Jv4a653xIb3fh3oDIIWxhOzTnWKK5cr
3eYAG8uU4plL7OHgfG3n5viHm+SbLf6Rwq86wew9meFXOc6DSgyS0YfCyxs4Ryy1jkxWTkmVt/Ls
g/H6NQSmSBUdLojOg0Y32KpwVy6N72v9Ryv7MtGozQR+l97rLgpMatFR8B0X82MWte47e6ycTmUx
hL7bBCYBmZMgrMvsTYLq8PT1BfFNbkvbHoEh1aw9VnI24Szrovx8k5tpWUGcmddlHtRFifgOOKPS
Q5VHp4vo15tcnK6mF5AxFBb22pQlVfrbfC14qYlD3Lb8ZQ4eWxeyJFfPzkHrkTddpOXQ+LaZRr0e
gcTGdlVjpr8nzi5CY3qrCsH4cA3yN6Q6z3Pn2FzJ40js+I/F/M3l7TQWIChhwUDZAtQoDXhciJTn
0Wh56ujaeFBzKcA2uag10PwEvk9ghGPKcENuYh6P+BzQA0gxC49rrio9dvFTWi30Ua7l0cx8wTt6
sjwRr4VazLB6WDAMpx5yLzEnqnbq38CY752rxDXU8NaYUFVsQ4ce3TTheVc616Cd/zYAHXtOk3ab
jUErk0icHxYjI/F2eIUjlUDUjXNRGKtbi9f3KbdKIZUogxlJbHE4674VCMX3RHT1kSxb62LWU/By
wC2BEIiDffTVlWSQ2VK7cbaUCgyLCxBPhn+xu4d5hH6+Iwu0BGQM87TzLdsCOqxWqsIInprwqxRL
y3bk5iXvm4sSnicvZB/A9ovIivxPNLlhWe1IqwoInSEPWC3mB1mw4ESSC4xRKFOgwx76qZfKlpXW
IQEDZzCyN2Yj6Qus8xlG5aoONnvU15TqFIntS1qeacvyjAyvX+n3n93aTk2igfGyaisucvIGr+hg
+2KXhxVyY4uy3ATGjEQVZBTFzRTikRY7BzdxVVEQnO+S+aqqWE5mISh3IRcXxokaSDgtZBnCKcvv
jsjBFgBq4y+YjemgQM2CWVaucZw+Bo+sNv96orT4P2FXEHWqJ2EY4dPymcyTdSiHK+eGmMRDW5lg
hnPafM16sCt0tYPZEY6KcIiG5HCi9SbqgxqPLKYRZwAkGggZdkNjzJ0KqThNOskAXLRaMXA/ICkv
BzH871zKsIieE5wv+tx9c31Z+gFGlO5dU20DQaZ2eosYEKzY4GPB+c/qvOYr4sLToW+lndnh7Qck
2e7tGaJBsnfQMN2wW9k91chmtfvhFgIo29mexM8cLFON+eqKZ9f/hCv9OluhDODLrZz41SytAL9l
N4/5aTC0EjRk6AJRbLj4N5f1mm2nKDRzi3gF0FmpI5BBTAk6kItbdpfeSC4lqkh8exrj8NDK5AK4
AtMiLHnXFdlfcftTKDLfcpex4mZGmKyu8RSdr2+d83Ek5aroZ2L4GbLTrf/nhwie6U1RtlDgKhjk
j2Eg3wrlLZIdBrDNnBF1B5vyLUhrBaR6A/kGpSCGFhZ7+px4EoIBWswOYXFOFRzSes9Ju1jq/i0V
eWdJGU3vL6Obt8qt+6AOw3Uc1OE5TyomUGUy4jTwSqWZksmukjXvE2xUMdTMxaPjz60A9zpoieKb
jYS1xy6dpNAvwQCa2P63EITNDd0kuWOEQ8SfeB9qyOsHWGIv5twXx2DT+6z38otBH8VjJo4P+dEl
6vGCIWFnXVywC5uAiGojGccjbZwrVOBOfVNqbe3TqJQtPDy92yNaxsbZvrB+8MAqnt8s81GzkSgp
q/vyZgNRsQaqAJvNKL19kZQCmfa5HjCbp6HQJlvW3X1lqdWW4uS6A4PBuu2iZni6MM7ESnU33dpu
TAK/0y8as6/fEiMhuNFXmsSBciGmp/D7tVa7KHMdaH63khHiAAV9vxph1CghtQBFcj+mLPEtWHfd
KH4J5tQUzmnEqzb2FoVUBbBd2y23+VNcFmAfh/vesSDebkU+RsU80eUFeoWC2HeT5Jz+y2Zz0yeI
vgKhx+uxoK/8TY9xiTHL6wjODZVPgvO6RgWzO1EjKvTEyFOi6OHzmU50giSoK2Jat9DE5xJ9lGcz
E3wFOh2GDsmeHMy963z4EQmXxw8H2cPrjG9UFaBDDD6QyOv0Hs0lcwkkDgClko0rHd0RC6g4CdOC
xBzwU4haehbPm1LCKmWzI1T8kq0BRQ/WkYx3J5o9NhQShgoWGNMdFt2L8wGJ8Zpp5KeKAS0sk/cs
VM8xAXyT0rEuNwkH6zUOyqpuxl7kdcAYT/x/hGki5IKGbOZpBdyL9zEdEsrG3lQm7RpM63B6ntTy
UgkG/4F9GLl528kszC+AIagElB82LKDexGHQ4yZ5jqVNNIkO+QkdksbjxNRaIB+iHwLSYaGrFQRw
HqYfoh/isrNTfkDOyJaNBIXwF134kfNGb/rTdU1R0jSltp44e5bDGBPlTyMTpxxzfiSOBDszG7dB
Ih3H8ZJPsd5EkTjaGm626dW6MXclEpHdJoge2Slnqx1ak7ZqSdcdldhzUdX43YrtuOQoe+/MD8yy
ohYCs1Ws5VR0gOdJQYSOQVeLSY8aX31RNi1qGeOfFL2inzTWc8Jp7/8d630CCmwztNDK7W0HtVyC
mrVirPII6Klt2KVnZF/AMpRHbCm9E69wR+uZqdhpAp+++WHKJ18cPLUqrfPwqKwMNa73Ta1y5AEJ
YwLAJfAg4QYTuNGCl7umAaNSVinevruqTc+XwtYqb830THHaV3I37qlPL/oT+65UuRq2PQ1h26yj
q/aO7WDj4HCnDzKuIz0sa/BtJCbeYaHhvY3OIsnbT5nAVmc4dAoGRjSojxVzhoo/VjmNGkXx3Lyo
C1xFEuuQlP7CP4kL2URX6gV6KuJwej3rfMI74sYwvYbK04ewzfCvfK/s2SretezL/WCSF2x2l7fe
L+ClUEiO7/CFAbU0clxBUyJai0V8m5tviEbdXw+c92nZnq3tCP4CUX7QaUCEGzVed8cMRLwfM0Ft
1aq5metDBtroKxy1wN0WfkO1JBLhoXZbc51nJSYKhL6EdA/Bz3h/rZOikHqYWj9hOKWQfU4HbcSV
3fWG1WUZVwzos3R/tjRadpf0VBMmIDGEombj4kH/Hc4XlBr/iksDWFLj8ZUecORNwZQlgaQngj2+
nrJ4xrWVADfCiWFPqU24hRFNcV/E2qx94ORLNSX7Qnz7lQC0wlq9SQkJ93inWQrsD3U7d5xY5Qit
19AojcqFjJ3zLjYiXCz+z9cmm1sb8PHY+zRZ4FX5zT3S2itVkdjHkiuIn2+jSMI4UE7p1BFyX/lQ
OG3LUeORUjF0++e2mIIDWowXVskt5Q/l/FCHsJH2s4Dc3d+YeOroHVPwIr4HXoBIA+CDwQGaFRn5
FOQDcEyxK7tH7n1v1zAE7IGBj3Gffjh4LRhmJ6qfnIi0J8ZtAB7UceQl8GNP1ZJhBLzwvkXEovFC
8+GvL/2dQMgy9mo5N3o3JtrgR7Pqqu1A7p87PZjck6h9wzYn9WxJmPWV8eBrP3xQGGm8hg1Egaiz
BJFYQUw99EAKzc5kL+PWYw0DGnEof/uB3me71TrUscZ/a7AqIOMQtuz1a/EXl/nvkQrZhFH/Nfp4
QzkWVAas5kJcznVFeg2XyNUvD44l+9l+9CLpnWAmcsZbakpaX2AbiQcq8n6/Yry+q8M2tASn7OF3
KT36WOD5S1X6sXhGPg27mA1v31dLWDsqg6l+g3PeLiLkd4XI4zOZx43sjRzQbcCtSUR/h3hLA27G
Cc5v4rMg/KYZh/vJG0T9epqpPCnSt9DJfuU4jAVkVHgz8B9kBRCyW1EQI/Bk/VYNS6uD0GPO+aw4
Wv/zEahmQ+pzg1kUeEbyhiRJ6NUtVpPQp5yySwr0I+DRP6JISXeThenXgtx/Ctyq/C0gKtzx1ohX
GrDmaCBAA/SX3n7jO0GsmGQwYv3tRWNvXZJvbCLLwj+uP8yx24a4kV/f25OFLiIRydUPVaE3scpv
nRaTQNhhqYopJRZtDefspnWXN380sGFL2E8nRd8qJhWhTlF+Vse0xJmbwio+rA5sPXzoAZEpiy7Y
qm++eMzTI6ubooA+0A0dsG0yZ1PFcfiU0w5IolaEjDy3JtxBe9adG4WIzvVyb3VelyQldwdfeF4t
wbAk8CNf5iN3y6cPQZEAElnRSqfpYWIGLlG5DEGdNeD4T62HEtvCcYWrWaWJTC9PQSIVB7iz+Ysn
gD4q8+u17+FTsBc/gR3BldMasnN/zCGX6S3TAdHiDkEFVjXNAkho8FwKttBfrfSK32eBLGDpeGcQ
3DW7gaZduKMi0aDpYUcfV0Ac4fKJE08dlGxK8CV+g3XdFIdvZLaAxcbi/y5G2WYBOANbPIj3wDaZ
6M74yn2cJD/RUTblJb+eY5c6IpjJYJidIdM8XCFt6m9Slfiy4H+98OQchiTGwSvIkX45tYEiQCrM
dO3BQgHtJYc+ZnwcLsoaT5gONAjfKMoF4y/a2OOfTkESCdl2/AuU53o3uHbY3bmsyzCWEC2ZRvpL
DG7N46F29bei3hO+C9OfRjrZLp9ZZAc08LQJ9Il7Oi1S+Jk+N/uy1G6+NhIKl+zYsh8eRsq3JX8l
cDdrfwgdA0PFPGcI7z965JIhVckFdj9fxz/Cg26QLjCzLfYJ6+KkncHiiU3rg+eWfBMnzN0bAWun
TUoW7UmU0kAQnSRJ74qX1rWnrJpIQEHDWE93RB32jDBsnnYl71d+gpIGlCggofLYE1IMSxSV9exS
r4IZb7Hpp5z1UO250ALiUwym7fui4YJ6wdgj/6rTb1YWm1coZ4iBy8m2e1xMUPLoOu7nvrSbdDLe
f31dKC7Xhk07AxYYQLMJvoCU+DQ52q3kkDjolSrcbU7Cz1AAvKIkmUDmoB6rDXDgsCfaDEOjMMD8
SyOpfPFiMAO41/B9RJxBMgDeE9LRD1z03DC8FaT3ItEWbxKOxr9ZBIaNJSyxwFM9D3EnMI6ln2WI
cpmzBSdv7KGseSBbr5E4u8NIztvYbiAUj/78Op6dRX+9+jR/ZorDtQ/zGCX7Z6bPJ9U2HHiKWljg
GXG0XosKhdNO9zOxtE9TUa+slBDx/8IAA325NS4+govGULcZcTjolodD1SDX1EF/+pT8zsHDP9OU
WFZU97k1909hHGwsalMDabNu2KYlb0AxEW4c2DdZSENHMms6LDV5yGnC5S7KK1gIUi6UeKH8b6e4
njHGtfHn3FFM14FsvquRNmzZbaU/c3wznZjhPqlgV6TsqyqUfbLRWpMwwV98T63BzYfmPfdTkkV1
ANmUDv/Y7cfhSyFpbQmmYUG6Aj8OzbkAbpIrnBdQ9w3A5Cn9I+hW5pVhuD+s7A8EutesbhQDpsdL
VrBLGmIwF6EklqwGykvxcnBhnPLQ08kL+JIe9SzOcql4o0oKYobpHaza1OLqG8JIe7k55/+txZI2
F+avJgpww8XbZSyUIA2icMKStHNPJkppPdVHCF8K8izH67fszTmqod++xcWkrX6BpTauSjRjAe2e
PSfLvSq2zM1W7iz/+ZKyVEcKii5s4vHtlCmxCvubhuzsBxwuu4o321Q1J5SaPay9g0cw0MrR7ReT
8shhIYm6DeW8nvZmcUotc2kSbya7G80GrNuXhl9HujQxvftg5vrIqdW7F2ELHTBcEPr/sDBQbG1X
vj+k6ynDiczSh+/uu9YYzxK+q+HTJ3TYXRqhL+jR6YvA5AdIWSPRINtZAFHWF/vv9v930eKp17kJ
BiejoFuf6bL8JnPXtyUBq4nmJNcKyacLtlMRhs5P54pu8514gRacE7Rq6xXU7V1TcemzdP2lHBMa
ABWEYIy0APsHuAyuNmSrIp8FZ2sQMl9uHIVxFs9a16gJN0LREP/dG2eh4Tk7KnTrjxaui86OKNaJ
FqZHy85Hq3vrG855BySulxBnitNRGItNh6397nXtyjWuR0yo5BL4IiilDohBGomXBSSJqbATwD1+
Zc9YYQHWYTQ0Rdd2QupkeSm+tkLhoaf3N+r9OAlEZdNYR4rieR3nOyW7XWwe3eYako/3OhrgGArw
j8it0g93gIVp7IoppI3RvSwMXA6CtulssjoHTeiI76mVS+FS+3oxK+H39C8bgGVKJhtGJees8ldp
qBg36yxzT8o1nuZlmdGb/rqZ5tsB30z3mtLCzq0GoX6fOH9SAGFr9mvpiM8sy96y3L5nQq8BNnIA
L/NCrR57vLf12NCNXQAx/h1xENeRxIJZz1wBaS0YGotOajn4/J9RAH/G9Dr/7lqT+sRj1zMmE+vX
K2+pHrdAhD2QIppFRr/8fQ4wiPDl/x0/qG/yicBs8PgC4zYHkOta9QXVXfDnB+rjyt8H8Yhb8QAH
JCAHx50wD896EoCaSgQf0Pe/2EBfSTx/tQ8MWpX3trs4g83oozDrP8pT470YRhVBcaSXPJoE7D/W
48SVPj5EnIeA2Ypn+1ZdxP1DeO8F2oT1DaJ2lQTrqerWtcd5vm3FjniQllkmCucLSEC3Knzg4iJX
W3oFgE87n8OCrP5yCFgKV25ltT57gfBTaMHChlfA0aI69xdtu2YS/NX3QEZFIPiDj9oLAZ7MGguj
N2SwsfQ/KXRoXZJJasG9bWiXeUaLu+rzOhI1hjaKrYDU/sAuMKPzUevvRoznxZhdLR2x3t1xty2x
Ct2zCgxzxJ8sE8kW0FuPDDYkjbKromHl5iVjU1i0mMVGa4Ld7AHvq/xt1NVqRegyTny2/RXbqsM1
0VjxvubStEt5eIDDrvRJDTtIEdCQc3g0cCtudq35ZgRax7NXs8ywOV+b3xDG1qQMTjz5iGWVayZU
eGfeOBkcu/s2exG7Fq8/gUkH5Re8X9Z5e4CvRtcA4FeJU20IFbHs3pPnUSek5awWFgKBwHEg/56d
Lz5byp5JBrMBFW/oq2igGqZGHURXScgrmRSA9bX2XHfjZZJJLCZtex60fBSCCbLn/Hoi9WuNqqGE
MiYDjUmvt/LEjxpBTFfxWQR5/wB/1mjRq+Pqvuscfrii3+HT9gAYJrKF9FFv9R9IdQSbtIotuR+d
6Es2TTXsJz7TW+QuL077ow8RVQNmQOhUHheTH5mNJcc2DjpQnIAmD4pEHvshDrsmf+OLirwrWTWr
s6Uc2MlQf9DhSXTvNXH/u+P45AtiUb9EWma/IkKZ9NNcVrHpC2VuVX9QNE3c98xY2sfYAcbxvYVq
MIalU14M6mQtFw/36cs+ssKHffHmFD9Z30ZpV05WtdYU5AtAFtuvtajFdcWAoInGWfz+89s7IAbz
uqU9DnMgnZkpuVtHpsCTs1gt8I+cW03ZeX3UJyJ6tgi0FBiFecnJULDJayiXPlQpyU9VvKcWtzQW
d/bWyGIviP63F9sTcuGTZ0LK05ul4mk++gnW8WwgY2jx70yh2WRRNESz4J+Knhcjn53Mn8CNyYhl
q2X1AnkpQ2YOvgMSgXQmGbiNiOMDJEpIp4aNXEuQWDdd7vKBM7mqoDasImOSXwJoP+f9RJOKU4gc
Ce53KxmpaIk5VC+TL3VcTbbjxZbJ7aMDLxuvvHOwjsm4oI12Jf3iiJ/aTlaJb3MO06hOWaG2qPWm
5NGysOXqQvVfHIwUwrB1lq1hz6kSZrb/+H8x7L99kEOQtCvh/MgB85g9pPc3pflaiEKjXgaL3lya
wCjmWrucMPaxsDvfuI9PfGPq9WUPN3PULyz/H0+2rt+/x/mYx03NwXxpGP7Y8TK/p6D6C6efyF+d
tbuSowwm3YY56iO45cnOrWDyb9JZSm7n3y2Kfb041mkfX4SOTd9QJ2+75PeTFPcyo0RLbPPwVU16
nhu/f81TjHhWYHLKjk+m6hLrG3FLvetPXwWFjTBajucynM3ROKQf2Zn2+swb2q5/D1pY7HdYlMqB
zr8ISvS6M12nAzo/NHecpj7DHKCao3v1TjZIQBxZHOUKXupQCiityutG4EzDH7CcSQbhu2xpIbL/
Rm1CjgPf2xTWsUdSSnm9ykg2O3nOqbIW/HWNWZ08pOQVCGbTo9gRQxRsstjyFGBtUOv9eaPsw+9n
0tRv8iFLJYvkc/j12dm7nrmdeb6hJK8xk6wOep72uegqGjhb3mcsm3UhObyc0xVSmzZtpcu/q1YD
56kYYgEggUn3OZ8JnVJga5g5Ft/7Ldw1tb5kDgfxcHdm/0TaJb02lyHvrzOk1/vJlYUFh1nkJKS9
CrH6Yh1CgFT7CJTN4QR6a8tprZNRxYS5EsgJOdn5TsIXGr1ei3wljJBVXwcgRp4i+dnyqQhEj/IQ
HIdxsv3Q+LatettT1xiCnCwPzcCZ+WOdcfVGcty/NH5EqVwE8ov3lIEJQtJi0/Www1M9ff5bSQKp
xisNAIqzZ48SpkFPkshBlmS1Oxua66/r8ZL1YLiAJ1UtbVwoAlcpU9syGUPmHtzIB/6NOavLdc2x
i86bvIPhSRd/4lVVBla3XxGs9QlI+h0wESAZ9QiN16CHQ32dDI/hHdgYi59910mOg+AbZrGktvjx
VRFu1TQVT3cV3MSPCnVESH1SS9Df9ckWaGKXStHP9yjIe3eRERbdX++B54HXN+BXL0og3jnKCEiX
1CcxEdCkjw/kFOybRPNFcNwMCNWfC1ciLMPf9L9IJfx4/dVb2zSN4sOuA6L6Uub/juQCJvaFyD/f
3nJKviZzvSpz8/h16eAbLqUWDEfrCA/uA0Yl81eksTlVleHDHiHZgKtxUD9Gb31dzeyWJ0R5hGYZ
dwW66jDCitr9eGvL4Np3Wn4z6G4mgt7Cubdno/n2c6mmkfABGSInLAr3qtIQcTils/YZYzF7WG80
/4fWtEEV1REVlkAeVVJl5t/402hCvuZdFRpHn/kJyjEFeTukcp+9m2y8cz4uesfGeoz9YA2SxO/m
amwcde0ZWvabWDIvdhoUVhOT71tLaCzhujMBCAXvxwFoH7y0MBqTqyqdMiepOJdI3610FiyKvKCu
/+H40RQmGB+SpQS6NUVqNzeCS8wKdSQNGSo7k3QG9/DtQ8KVK0VwJzqM+wNhIw7G7a9x2zIRVa+e
X3tK9OWADUxa/c+PipgBS0brjtsza66v6W42QlYiD8j9urCeTM7TDowhBgUaClkU/wOjt6YHP17Y
a/sTdEh9kzP6AZHZp+DKfMrFmJiDJ983kXwLDpv1GPe4Qt4meEapQVftK/8FuDcq1bmn6Mghomth
VivBLczZEjrhAbFvxdK/Zxkv1yQmsmpXnSB/EtU1iaeW3cuqBoSzr5tKhzGsmhNwbICcq8AsT6fy
3hZCszZ/fi7qXrRtTZmUny0cBhNLsVWPwOurmaXb7l+EBY2gQObdwRZvy75i0PdP7Kn9QqooLpA9
JpCx/EsPu6QiW07miWft85YLP2kozMFIHtIGD45TlI0kRbT4QEK93XeGHlBDHctlPNMA+W0OhNdX
p8M3eWeDWt3Rpj9wFIdiQqIQ/rvNX7/jO820S8fLiS4wQ8uIrgpmYgtvhM7DbkbpJ/T3Xokppast
K+NkqY6haoxTA16AI9bSrsmBjaHae7EVdotUpJn7kF1kcy0h6xcWUvPVLtc8Ruv3+4O/HaSJ5gPf
E2G8tBPrieEQe06XIakBBdCCKFh4EGf564n2jd03yaafiuncIaq6hzqocDdcFgL8FCuYaDF9yggO
fgbezBcwrZoHFeAJOV9Mh26l7JYfumXwKMQluo9QtmvR+RTgiR1pi8Yvf86UwCuqCPNspQ2RIsr5
1dHkW1tcwuallTaFyEIWYJgZWDsRh2kt3sxOtoPSwkrD27wSHCc3tZi/9dHnNUWaX/r7Cc3xukBp
IMN04qxk29hPSeSSFCxYnQA/8LHfr+pd8Aw+S5y6V7CqCnlNWmmm4gnzb/KYHDsDiuZHAhqOWHn/
L+n3OdWAucbnEwQrGEfVbK+30gPXh8bDKx0Y6J46MwZd+zZzMlNbbKcMHNTeWJbYNdU7JSt2oKB2
rwccHVWp8kvbrkO03e3DigfYj4M2ezEwUiE3JYZVWv4sJqSb4fbgMi4yk3pHjaot+kWtWHr8Q6aD
J+GHycBLVMXR07p5YgLpOYBDU9zz5JmPNxUSLX1YlAs46xb3NKaPMbjp1hPTC1A4kWYVqz3H8HLo
1H1d9W0Hvc/mYNevNC8R5y6pofjz1SbUHKZDaMNGkBsHR3tFDumvbqQKYBZvQOOx/1nKQHDcCh2c
OBL8wwbsfNbhbXNYA9bxv96e/eWvDbN4N/j6BoN5JxBfFkkCgB3p27aWQ59RW8SfXXSIAulGS6CW
DKl1n6sgUJxKEG7VF6U3XmXzviId1xUN88cxiYz78PnJSDobqor0sV4110ktxelWjRIzLO3mCG2Y
l+n0Qe2prV88XobswmcZWjqxzvks5yve3zA458Ksqw963pZIbPcfrof30f2z0HTmJjnIcBr3CTZG
RdZXvCUZdvGm2UtV/gDBO2L8f+RV6nM9H9gky3jMueLolkqYwrNfWpYoChgAyrVp5O4OLN7sfz9d
YI8IUJ6gHBqvWefd/m5qdwAVE4qfuTnSjogV+2U3+MAnyj5MPSXPF4ppDMJ2tGoMxXkecISM1fVP
KRYYlp9nYHqz6cC+mpAkaglpn7frpep2FO0fY1OwcMfgogeBGJIrHM4kYCswpwH10ZIrIDtvhPqB
bmK/bv/fPcCpP01T81MLCYa+KTlUj9gXzbgxyzODIn3GtmqH3eQnGJ1p0MxkO7iBjqaNt8/W+MV/
kZYMVWjdZwi7mDOusNLn3PaxHN1LXLx+gKyMAwFxdZoDeh5KrpR3HZLtWpDrruw+cS5PMl265m4o
Z/bRFeB9ez5vIAmeT8+HuIrbEDZ2FsO0sh99IoZhxhp5gYjWDskoOkjqQKF1CM6FfaOdju9eM4/6
SJJC0kob46YUC7C8tjIuNDj7ply/vIbmYr3NvXG0V7QWMsRyOyH4/Ow/MU6GPN1YHOyP6oI0rbgM
hUsqgVH9mqJJAGuH29u95umxAvMbB/Kc7XqTzngiZyv5kUTeNu8YaBapIZDmOPfeLeK7Un7E5Sgk
76J1CPrekdcMyYoz5JML0q7CIL2EoJZUPLEmAtNDW26m+n2dny9hhGb8EoZZP/6IsfpmGIPbqvxq
iwRNfHR9TINj1RJlFu2V5GkUkqjBfkfD9aahuRMvkaVhdnbn6aeF+roawGE8j87ePo9x2ALT8TjN
MfPgRAM85wCuTTv5JqAhI9P5EWOOfIdmD21F97D0ex8tiAD/PZah+Pvkjlicg3yAu1hSUmiZ5QEP
b/0bq7aQB7MkutRxWXNnsEyJlI9oAeIhPKkkAlGFhZVpbfRcFhfTqZ/Lc6oqp+GiODE+ZijmWc1q
zQHA6cE0hYQlvIv4eyJWkcjvYxP2Pc2VehoNwKrXWYsW7nJiP8+Rd56vIb3kTyzCm/FvbGmn4jfd
f6rSEdK20RT4bGGTk26ymkq2lO8r42WI8j3VuJXoQ7EwY8v6Y10LyLj3DDgHFNmYQvXrkaFcCuUr
YE/C+Z0EN1lxzwJc642ygLxzD1ybcbq6Cepviw9hlzYpkqJgG9zlCiqMqbe2aatpBzSAPQRe0xyg
aB61O/GI++vTa4YoZjjoI0SaE64qj+E8UI8gjg66s7PSbq1glsViZG8eZ5Xh+tH6LOuGy95nbu1N
l9SlLIbdtXiSDQ7Wih0I2ZVOqgYjEs0w7z9iGJkjjZhKu5w495MpbIzdzAEdtlZKTMz6Rckwdv8B
fiuTwCCiU6xKnELku7kMaDGKys3CRbgabxEUxJkOJO4JuTvGFpO4Yh3dgjTcchewEEZ3I8yqQ9g1
hdi7otZR/MOO7K9+5q24yzR7NHgRCOGfDdH2YlgIT0diAl2qYu4n7/AjtXfPtydZprf2sfWVoLpx
6xaIi73M3WUVwOq0p+doAVbHGEnD8Ti2WxuU4/QIXg5Kxw+bde9jp/hs2OvgFDOIalAU4CdA2511
MbQqDA8luBtMTcZN1TFr+U/MaZzrbgBprhljx+CUNwMIighWHnxGoaNbZbnVJ60xEUe+YUVVPnbD
X7ZCU3JuyqFra1Q47YyJxAp+2yBzsXwdc361qJzIrDi/rLbyYfTWbFuEurjt7/HUPS0SiagtS7+D
M+0nlhkxvap+IMWlgio21AzsXC5RBBOrRn6jEk+/pbm86JLuZNhpzjPn4QelcVKyBU1Xa2GE9Evq
+5WxH8G1rRzX4WD77KMEbmW2pbgrGQxUOv56Ljl1ubAHCidApfH8DgKqFcNjeSXVsXzAQvv/6Pun
VJegaSFG0P6JXKQefOxlO4e8vGfqkIp4jGJ5nVqkZamVGn80A7gzo6grixffb9ZD7oZnaT/PhPT+
/Hb79RbVMfS8sbfr5m5rUbXMmkOIi2grQX9wgQXIWuA/atQXkkYvdCgEga+28CWBGi1RQREOsxmC
PwXQrNruxX4p3at6CZdU42ys/eiefhq9G1IR/1Z4P2JaLDkvuQe8+j8mwlG5eGFhIXnX8X6GVtdS
j/8R8t01bO9yb1BGgAGIE/T6Ja5PIKN2pfPfiM/pVFPBd6ZOILy+GN7Ojda5yetzwwaNPk+ip6XT
hxuhJKvkeZH+vO26eevuuqm8lh0h4yAZFo3dh5sl46Z4IYE2CiNxuU9R27FevxrNV52tALyyoozV
V6vn4MXj2/5/w90CxdhZuoLb8STFBR0/h8DwIvRuhEAPx/ir6KDqDcsghxDscGUvGFG9NpL1gnKm
5qG4uV+B71NRQmiQd8chhzEniXFDkI//IOfbt3DGNoRp4Qko/Fa2T7SkSflJUVAs1GCUxJ1NjmPW
si3NNAiBnLAcT+n1+JOVrD6mIRIVAugfKuoBJIkubFd+YeyKHhaPTWIr3AaHHMJBoBsHpJMvcMbi
cofwise9tlEbp3gM8FJc0h0tuDDmudmJ7LZLRE68Y0qlVqrOcxuTLJFa5n0xj7MobbH/UurCgXEp
o8mC5EHsI6W/Y7NVcwB4asMLB5PQav7s1+07klkGP3GJJCvVvbvis2wEzxTGEekg8sy6Uz9IG0H1
kNNM3qgBtne3GGp8mSwZvR3RcreAz7BXt2BaJx3aLRcTU/Z/KEr8dxWfcs5SVuEk4ph7BPXEXnhD
0+CYsr/ToRCfVDte3dkfQMBLYM+FWGeCSS9L8aSyWHyY2YIW/wnOJsqk/FoHf4rsVGhH1rFKCTm2
BFgCojhERmd0rutWL1IGyoLn9B73EagVuXrF006ETmMgaTbT2WTGP/P/B8Nl833WVbXsRZ4XJT5p
Xd/8gyH1RHob4aMca+AAfRE/csLoF01tUHabDw+TR4ngoW1y0kRLFtQhircd5Bqayk11tzQk0j71
7uVkIhsHA61Vcmr+g5hriHDLxC+zJ5nSAFs/YubyJp2Cw2/VZwb56xYBtcKGNywx62QkwNpTnnja
48wjgeK9Im5uRReIF6Qg8fb/nrv7O001QKNp6eHKrm45jMUVxhGwmowV1cG84nbqPZsJ9bMdruNX
3tV3giExWVwfiJaDGqwlc4XXOB8OvKc1YnDNltFmf8DOaBV4ulTDbbPmWwumftM0zUq8kY2YZhLW
MmjYodwM+wbXS1wZWniKFnHvX538OvLyhNUkfaPKNhLp19meBvKrUFrA6HfjcBe7b8RzIG42OEzo
mueYDKGdnED6sFvqUC/5ghnRUykg/KXbipvlP2PIlem5AYxwlc3k6flqcPpx084VeAzZ6IFH85E7
X9fSpoBA+WpqWhdlJdquMYgGJMidIGmkhpb9RYBAJ2FiN+XVBkGHnKJvhMQlu2zL1yd+HHN3Ow/h
L9S7LAQbtmWfLU7WAOuFqFvI3/PQnPSI4YS0n40t5qaqo/TUaLYZOkBuJyFdgShz65pWpkCrH+He
K4IkeIJALiivHaMHM/q24uP8HWdd10Q2M7wTjOHKJphPbQyemtEEIw/NYcwtAuGkdi7d5VZ+UgvH
ambE0MT7FVRV6MnD2Y6yRXlDQXgjIa8gBjWpQa5LRyRgRPDX0pEaUNLQzFDhXZBLwsXsLco4hmnr
GyxxNiu0CNeScXi5svlvi1gYtJdgprt7UqGRbim5gReVfGqOZWLRNIC14tCb5GM5rwwhpY6hoc00
K1/UjdjdGjxG7skc3QzIzGi0QtgW+EW3bSiUpcjaLWWAn8Is2ZNnMYuzfFtm+Twd8p/H4AhnF/gU
k2SVSpA6s8EcImyj38SVCZ+cKNjWPo0ADB0/7FABbU7inGkt6Vu5R9Kv+1p8EAtPBjxDOgrbSSBl
6WoSRvHsvVpcL6jivGEMpzWmAv2BeZSIXDWl0RzCqdiQK2XOTEjZ9k36M4mt6pz/dT7iJKaRS/++
RJBxUDrYbPnoTUnrS+TSq/sToSTsdMZlfYO2Mo7JvalhAnPaj6BhgplUa7r7nCk1JiZHbPS/tcu5
9/elYhILyMG6zpiQ+StjAdDcBs9AThjfgR8UbPlzL69Vy/6b4UA9e3+cJQNvQ2oMuT8R7EQZyQtw
Os8RfUC8zFvJAgQ+ysEBU0JMXC0DtsV8x3WY145Mv3GGQ2KU/vHfcJnIXghaw9YbCC7SXFPhdQ1y
gfmqjKJ4M759PCXe7i5c3ExJPXN170l6C5vL7h6kSLla+XbopjySUTroAhQrAXZeJuV6S2uWU4Y5
BbkgjctU1ztlomjMk8uf67kLCoFY1F/gV906V28k00ZP+Z77qF2oyLFl91XJZ+fqqJmLwh10VkFN
YHSzcCNmjV0yrjTJaFTH/9n69ltKmtnNYIpRPgqWdFgM5H2mAQ6XmN7AnoEpCSBL8c9MBETklGyG
Ti66MGMKVWfGe3CgkY6dF0VvjpKVRosgvtdNRbnWBgJbnDD003dOor/hGfE6fj89I1PXQd5CJ3aH
hYMQhWRgxOd6JFax2FEe7GeEpA19g8EzKEEFwWVzn7Z1WL45Zv+UQ9mMwhQM0paQkjKm+mh17Hie
qpSdsDWontkq+DB+SWd89b5JKATnerA4WxwEShIg8UKleN9uteBlCaiQhK+MDLn/BaCASXwDSgcs
ychW1NlUpF+lqjnDHR/OxZ1OQcgQoozq1BB9ko9HgLMoCfgiEfGo9DO5tm4Ja2pyhyMXfeZz7lV2
RXufB6uJA8d+myUivskc5c+gYgjCwTRSn72wN8d0CjwVpA2X5Um29kN0Xh6a7HpYUqcoPAI1y9vu
4wo1bZtlFsveQPcjBTk15J5dnWhkPAt8OkH8aTKyUw9qvPeWY6B60woPDAqcBoQN/EYaV6cuGRNL
YS9QJ/OF992IzcFMsUM1mBkk8blIyMiM5zC+kMSBI9OMlyCGwlbdZDa0DOqjQhAuoaOKVNXEG+Fy
zVXP5rmtCDWwcE0MmPqU1PIPyJw/AqXpPsmDM28r3vBYPQSiBvRxfRBuxUfiKjOo3SxxXHKTWDql
DLzBonVBdD5HvahbyTIGK01hYd8NAaaYiiNBtBjzpV8MINQs0cuTYkCSIoO/3cI9UOao0xmcGGNr
pDmr93KAu8/5Xu5XaWBc/oNkAVX381fyFOOKn5To2yF4VenVmPmp6QFg/hehVV7ZpGyzwZqxBiE2
GSJkHo+iIRWXIeAIxg2p/RQ842TtxlDxWOFynOO+RS8HCkTXhWWp22KYt/cE9UYVY87J19gUZSZv
/A3qUPUuKxUQ1IdxdXoxSP8/mGdAQooDGPhit6OMKE+7C8vkDMiJ9uW+T9BmK+OeZu520GodWRvM
03P56+B9XecvkPM87LYY6n9s2RXTTvtSFCDoWlMYWscopoBRdq7ZocudAN1Z9c403brv/+2/Fy2c
0U0rwFXrmfVQBqh71xcQX9VjCgcgiHCgKxXwdNfy7te2GROdcor6h+fKFdheEJJp0ISCwM/oCIfc
x7B7AiC5gmGE7nPc0wF4V45cZm6GVNOodhSUb+xA9cbMmqrjaKi1SVBHGSzrjcBoHa4t4BxAqJzv
8aR1dISSjEX8Rwg6mEtsBlk/V1n0d8WhLI95wyrftundkkL4BdqE1JO1LZwVKmIrss3+ZtrpR+VA
Qngef/SGGzh77DPZRxYUDx6DTJWX/EkkscnJweD5GrYbPmPpgZpPbLnNNcXcJzjRPtDGNS/DRXT3
Vr/USqqapNjH1gRiRa6/NfuWEAaDfU34n3FTtV2J+JW8Izz/f5qSub8HRo2BbuKtgxyKmKHByS0B
I0pvgMTg0AYDySE+fctF1uIXF6vIsz0iGWt6JUv6XjCehsNJxOhGZLm2WfGn3AkbIRc97K1iDmHK
UFGD9I5uE6Y4+NJ55JOvwoAeXesbZnVDwbNrUNwDJV9qs3FBdbtoUEDDlsN1y7EwK7z4qZroaqcQ
0REdy/wEZz4ehQtI69AqPHtq8SMQB41dUPsNTlGI+a+ePUXM19SJfoGb+wB2iSsFFw1tQrqfHocu
N0KJvbGCAP3J7ug+oZvag5P404DuQ7Vw31NKlKLDoVtX0GgjUcBIPJZ5tHPKt3gdPjjwDsZCyHXw
N5i0HJDDAQIJVf4EoYdIYShOc8gbkzi9T2W/iaCo7V94Pnfkjl5NZxJPYmwYemy4v0DVhfX7fPoK
aSqLUwIUHHZ39iq537gPXaSSNO/aqZeUQ7N7rPvn5GRQjqTxew6lRYWuuQ98t3zObmdTfyDhnW/k
2/2mhMWgktha7jGvqfaGi4FVQpvepJk/alqldblo3h+LJUBlXunev+GLCsVKj46V9Ragw48RIalC
nIyE79Bo41tE+ZTmKBzynAzTvRwtQYwm1hXt+4I78Mlo4vMSOLKVeMazehseKPptldiWoKCrZyyz
p557ntj2m/5rYotA9OTFJkYYa2bOJohHF6jK5F9ejhJ+VNaFlp2zIPdZtEGWCuSQgxzCNYWyAu/5
PMNW+JEa90e+3FG9knoaYXL0SwpwBkbnO0KgzFZu4ZyYoMordaPo4w34vwcbQsFhlIkhYympK/1n
hs/Ic2uiytitw17M2OAzFORtttp/dSYhw7/2mBnGFwfqf+KCWETu0RAKBt8V4CV+T1+z8iz4/eFo
uxqOr/3yoQjGgxGeHUcFiTzL8E4i05cbtYizqiWkryQoURvsX95qgQdPKOZrZUdLeCTepMxOUqcZ
CWocHG8YAZ2h4Q6rnEQO9YmJwm0mSxWthktn2dZFWPBQ4D8GlNiPYQlhaSSBFmHE6AMfla/Rr5u8
C6tJlOw1E9oWxKZBIemCYECT4Nze7RnEaOsMW4LvkfZCP4b+uxLyuIqP2NJ6QfHCAu2+xTMsVIRC
0Z+aKz3IkcxrHGr4QZclfb01RSJafDNelQe3f/a4CzVtFGh0zrHxlyYbt4Vb7BlB2gMW1iQfNdvO
pn/9GobxBFuHz6yxH8qtp+BJgRsMTbKcwJnwn+BcY6yQNcnhpbTUiRjP1Uph25/9LY6bK3Yuxnxd
r5LyBfFxTQp5QzQOPoO3pTthSt6bWvVWkan0hkZtinRJcFZ15bh30LKsmT7Un0q9DsFix6OrQEq5
a7SPLow14k49FLy1qyRkQwx9qiUL0V1rVHiYX7GDV1+dqQ5Ngywb5AdXuDmaWhNG9Rv7Pt2FVgwr
TboZ0HZsuYnUP/7jYUJ6C7dE6lhcHmEPzh/0FJFc0kgl7zY2Uqa0mfXdCTBj1oIkLFJGnYqX2aKI
f4BXn7aV2bjjqKqhzHfcxQ4bpeTXgxS7xk9j7T+7D7V1p9Zx10oT7tqhhY6uWdZSothoVsQOgYnn
l4BcnVC8lHlTFpckqD4QmbjLpE+T/1h0WHOMiNpgDPQLTNx4+GssWDo99NQyK2bewUv+Qfeu5PUt
ohEtbuk650rJfSYAwes3DKiLelJ76CMjduDHYXGM4GNPR/ncYBXAR0CNK8YGpLoWN8gchLkyjvYp
DyMD4/znzxfluiF5HQAdowtsKIDtqwCWjLoY1il4Z5KIKfScA6y3r07qQon5EqBh8OnbwZpy9DQv
SisA3atoEbJbgUGMxfBalKcZGLR83Qni1f62rzmiL9E7GKoXilSueE3R9dh7tu18/sUxw2Zrma32
pJsK+mcNyLx+FAENuVcEr14yk+O6L+QUYs+be9r+fHvR5RbLTILyB8BS2dQpQaTxM6UxWir0wKGe
dwphsmFWZCsrl3879W8Rcwm7UzGtARY54KwC8zDm+n94hhGSAz4JR/Te4OM7jVCeyHrXLOa7JjQr
g/z86tZokiIqDTniIhgIcl+BGCYnayzo/12DfcUEzdkAcioUtlJ1eCqnNGDuw81+McSkI75y6ZXh
1tq85DfsS0loHUKFqnzLnFFZ91p/zWVk21/4sc06QMifD58k4futszMDsFaroTJFg+9RA+oukbQn
qjKD071C9nZJlEbHCzimzI/52Xl0+DjWaUAEss/PA/42rNa1OqWS45wkz56x/B2BU1R6R479W8dC
lsOXLNfClbqLbarPSdyEm6YFapJWkCFCUmmz7nuQK+34l8+WTOhKO5gaxUpEL4edCsX1ESN+c4AH
w4URmaNXgcBLXyigbuiKsKBwUye/4HUJ0MkZtm1h+dyk5Wt8GXVZ+slQV4u9d2myKzckZkr6Lu/S
YP6nyleRWrfvwr+zjZn1+HKLLxSp0xAVrxtMQYAtfuRecfrMo4qdvsotI/8U/ICO5xjpGDSFa4wk
+o6T15SkINzHnTJWIuw1XaYmjectwZ6Vfme4GfdEu8Oe/BSQZtP4GhRr+J8Bl7DedKea9XofJUY5
1p0eBmAWI6AUGm4QoW5umI9JWeQKqWBfX7AWIhJraetN4SSGVjJisgx+myuPTIZMMZg3QQRDNtH+
Wv8Hgdzb91KMPmIk//NUwxnPgJGMPHv9eKQ1orPx2VBHXlRWBJwKYiuOOWdUE+pMwe3i1ck9DJRi
Ll95RDuw2zvZshPKUk0XH/n7R/mQ1yoaUEGlXV8VwPSGvMAkcKqwCKlvp/2lJkFGuTZs8LKuywmk
AbcrFOui/jlvjIprjj+TQMQOm4JQ4Yqz68qXSUFS3DbtOFbRnKkOUSp494Cy1Vtk+KSOZRWQGjmL
CGe6FUvufub7dveM6it6nS7E9RcT11SRnC7cNpLxRpDlrRqKWldyeeBzE/feaAe6Mo9PKPdoNQVx
hSp0F19kw/6/XYM3mXqlAQPY0X8dxt22bfd52Ce6Eag2CJMcNGXjYfE2rsiSSu9V85qX9zivrVos
F3VwLS+qEv7rThN0MR5d2BT0cUkKnzqcMc2+g54nPJ56jvn+S9jqVsTgX6H7qv9a8Ne6o1XSrRW/
EY6jLW5pqHYqhek9vY4MQn73ezCLxy759GAKh3tFlXTz7l+Ph4JmzXBN0trkgljYgDSgSO6FBlJd
IBdMMKsQI9vxcODHwFvvAhn7fhjywBGoONjUURKxLggqbUvfDCMwb3djdzGTYzPYRCZMD9CGTLX8
NXbAy2p/dQvalwQ1u+PhasOD15m7uz3JVTuPT4hHtXfZtVgacY9q0FqQn5sL+306eN64QH+I8x14
/tfMy4+t7rUeWHzohtjl7/ZsWsk3G2FbZA7Si+A6A6o1GGVzLPpCjtM1c7NsS6tLggfr2DSbAlVF
ew1i9FWhzHN5dmQR4GBNkRwhaEs7LEGshqjRX4ZeGzKw0scUBf1a9lw5jTV4UyCvTLyRQyYkNsc2
r2znb1WlI6OWvk8f1JIG+w+EQ9HUQlApsFC4DJkULDMvyk+0pN11ptqma9HpAQ5tdMjr37wYVuEg
Uhz0ayLBC2findLXRWGFnpNNEp54VlNI+1waOe9wZfRjZhWOmnfozICH+NcDDy2je+6QWQ1IVd+u
pf24Pwu3EOd/8PKL5lz3kegtMAzg2DriXi2ROO5CtQROkmdA2zoaYcWREx9THXgPHddahbwYxkV1
V7TkdqGLAjp3aSr8yqbTDsKl06QYAp2gyctxlsBGfOv0rEvTKGFkPxYuf9ftxYMdDwaGWozdUR8Q
xKyKdlMje5EdZBasCoppA2Rovyt/sQhOVtv8X6L+cxIFEBb6W8kaZfNsIFhhltxiIalhzwaUmqm6
OuAUhf/z8MSX8TZ2aQBuoBdPwHl/X3ZCBsdEOZIREeQrMcHYFh6iiCmEh4OL2D30gHVd5L5tUqIr
Jd++3oQfkR9gkw08xnKfwEmlXLaf7PN4c9TAxNzQVemi2npJcm+uw25n8Io/XdJ/PjWYH0im7AAm
hqsT5ile1kYYCxv76wZX3imYb/Ybyd8j71H0P3o4xsTsx3SsrZtesTIAyA25GbzTEFDKfxnrk3CK
Bg5b4Vadmku6NdvaeDyr8rcBSQzbVO7Q/PGheq3wDSSfE4VRS33Oc/0aiuDCkYfp6CyOVm0ux1mt
QQR42ZFMO+IKW0xFOHksRhQRKr+BmkIBjzvxRNYOTXL4m5MuMCAZz0ZHWDcjHRGQO+QNuh8lgEnb
5O4lGwvZMXJLG5fUu7qThyxdvKwuYq0B0PPEy6Hl66a0dosZMdZgnRpR1kA1CCnt0rmCE9sNrUyW
q+OrlniRHaG9Z7LRAZKL28BzDfbDa/AoWFbKerUqAHVQGdgtsh/SMk2KlF40E+t4VXJWvSAptMRq
+vG9xkeIaSUgOqK5dsuH1jiSxJ94wOSWyc7S+wh8lHMSJlFy71n31d6PkGhmMGeJeC6h5ONQrL8G
AyScZPewEa2r0Jg0Xyab/mPekPH2cUYqo2cyk/xMv1SR4zpWnmSAI68lYmqnyNXyqYZip98XnTPF
ENb7ajU1xeWG1oSfrmor24XwKKejt+roozkNvDlRrapfVM7FGfDtSbDXkPDLEhiD0uHQKw6dlZwS
JEIKkJxGKovynYbfsd+ID0/48mvYD1heiTBuFlGEoqVnYiI2Pt6p1zc+JlnrgR0+oyoxJ4yQ2Se+
OYpH6vVMhYhkYwwajQqgr082TNvJOKG9TLyXMu9IRcAYFcinsc5JNq8VkXX2SSiz+CEcCYdSHgdf
PN1GFG9LbcyUll8exLiKQ/LkuCowcdje9FXuJ4FD66Kq7Elq8KvAoxFJ6865ZXXlkx1dWISuQarS
JYY2MVKkC03+70GOU49zACZrrysWPflok5rdr7xQOlYRK0V5UMgEJRgFqNR2xaGuRyrOcjkuIMV9
5NGRDjk4eP9Ul1Am8lOu66P8Zhti/8pLPRmx1S6i6va3cLJz0KT5txwVoMZEcLNHbKXtb6SNDr/x
dFgg3YXiYPzsE3Xhu1e+Y90/dOQDFC93kS4XA7v9s3c2S9COLYMMwgcPyA56+cHvcNZ8MFnGF0oe
YCjhFVeFlh13GqNnRWqLHUOeqVEiyCWBmMZHr7cTuzGftSvfjZD5fwN/sFSzMeiB1smWGVq0N7xX
1JaYuQtwQw9C9J8dORzw8J2IR1Y6TBk3vmWroMro8l+JFuoR5VIi5f5DKLG1L3LxAmhA6SMCmdcC
Rhd661ug5WpubqukMLTQotiWezkq6tWjXxGtLoTUNeXpJxxe1LT4XLHdsbBkHDtnrIn4c6sA4t9s
HJt0gxL3/Q3zUkDTOYgcliy5Ipi0lHQcV2O8LtF8bu8pBS4ITjU7aHIVz5nSQum4PTvGbmACafhx
bAkNb+CuNcFtPXV2JWckAKTXPItEzA+I40i2g/m3b+kta21zaGacPUcfRz4MCF3XXrD6EZo2ExNl
s1peE1Z0uwssdRrLiexVbDrDCg1Jrv9j0aWFhcyTqs27hBS3yZjNn8OnOp2tFR9huLD8dkSUfG+h
ZXVDKzjXnVfaeYbSYCEn7MCcYCcXlf4f0aulSLWtktH5uRTSW/sTxWTLsEUfFQ2mxBuh6T6YVcdE
/YuRTPM7EyOjGY+8ZNXD4c5+Cn2SKz68Vre7KBSE1C1V4QE5RWN32uCYXycnpAqnJWYOd2YMVW3t
MZk/juugTKJPNh8NWle2dvsAU7AA85aLQRbkkKSEGo44bp1L0biAu4F9rSJFp+aBP82TYSDLSxEC
ChcRuji3LVEEYQYjAMlIOMws8UirQiNrBCTDVee0iuMf7/62EkwFLENnkkuey9kU0IipkNMglk2k
OPKh8kv3Ow6iDdfRIP7Uj7sF613dks2G0+8cIapVDBvmXc6IcVmG+L9NbBQQxO9oyvPoGduNyGxL
oGIgwEr0VUeZEYMMY8aUhtgh4HGeYOkkHhBl44QNAtN0CjHX39qWXf9CPHHn2UNFNiOo5ZwKNkAa
6EtZrZ+4pwgdZaiyfUWJbSAubiMmC6vlwdzVIFlWI6t1Cam0VQlItkiindruZpFLtO7+ofm4HB4W
xMHFgGIwHP+vioGR5HKVB6R82feHTMwgFYTxgjRlIQN8tNV0T6WGNv1Nsr5UxOzHNkP30pMCvj+R
aZAAdVWgDnMd8EopLFup79O9705gjH3B6HO06V0aF4aFM9/qWT0CrWdrTITz46gx9ntW8pcQ0/ik
NeeDFPOCBEie0nofQ0cVRbsZ+ZcHTjnLrDsh0RdgdApnKmNvrwcOS3a/ypzPd3gbpouhdVEbc5zH
mb+fsgExs/fnSWBQWSkYy4h3w261F33rYpxJzc/+2p/BA2xQi63rIBI2WDRJZtvUOe5Tf/9o+kmC
lkPbRxFsCr64VD+qWr+HeQKqhAqGNurH2OE2NkuN45nACRenaRzKs0N+AVI5ijSv31nQtzh2CBoG
7LSo+276bw3TPmOoVkkhmotT7pg5sJdlWQ+U3KlWWFbUEd8Qc0SKFH0eHlj3PcgUUce1J+3t0Jg7
1ex+9j6HFB3CFOy/Fw/0KyHO5VJ7LrNGIIsBpjJeF+IpUy9IoVDKmiW+ZhnoEga0/R3bHYer3V+i
nAyjXkMDdiTDm0lKoLtPuUQe5rzr2z+lfsEqIdaIT5ZEJkF/sFXdolwFvC8pz2cwdPXYMwNMX+Ae
vLLfI12/9rHMDSJkzgsOILusDETHwYtJS2nf6nTNAgPW4iqBSxhHNrI6khCpWQ41qVDPYAr94AvR
Rj2XPONzvMJABXDX/BBors5OHIHNfZjJdDsz1EvXkeUSOZ8C1ZYUDUbXnlGLdLbNK/EcLHqOXnnC
wRRw7E7GQAPt30OSnDGZewx2Uj3jQsRGceD95XLjJzJXL4vERDVdoxlur3bfdthINsOdA3dY24zx
RcY3Jj8FWYYLZ837aRW14GSANORguOpAw7Bc3RGZssd/B6KIlLMB5KRQfwzLjdwYbkIMWVVyptW6
Gtq28/kweuwktQt92449DRdZid+jx1ZnFzw5yT+I9PN6bhYwQMjM48PJkSJjSQrjs+eOODYBDMaq
h16LdwhnQvbDgR9j6hV7Vdj9NHqR0lXkeKVwDvob17gP5hyo+z94AmRpYFUSxPKtV9OstC/UXzl8
aJrJfzSWcSEOXrqQKDGshod14L86+Tt7wc9fqEw5Cc4UpvSQzKau3zIjbwsXZE8GcdRNOAdWgIdb
K/h13nhL2vHvCHJGoP21KE58KuflCCfFd5q+UCsQ5D8aXQnSp0PCT4jV/QFkhPvuExNzWB3DKHO2
MoSkHiw+Fy8VD2QD1i+OgT9OlNzrgMmJdB4+whoDGkI9bdlI0he9I1/tBZ9PAeJs/lvTnpiDu0a6
20BbLvlRVFF5W994vB6jVu8vstxifUaklRppZPkbBCSe2pU08FBjdNNpqXDjykz+CsX7zVosI3gz
Y+GN72w+gxb0KTp4+qZVT8jLA4yo5iona3Blcg542zJxdJBtq/8uHF9JB9ZLVzTcLulR5Yygoala
3YDW+ZkTfYfU8LZYLGZGq/aoKto4hBqreOpUozu4dMY6TN88io3X8MISOIoza9QBLfcdHJWxAAGU
U9S3FVMAebQRgChdcnwiinMSJy2TWueYEQqOpWFR6qHd+xWgJZ39YtAvEpnQOr/tInUYcBvsk0KC
KAatWyzCQ4PnZss/FruQ/XFWV5G7dErMYIcG3VyiEKZHUkeVuzTzD6Y/79ZmOhp1+JcpNqntvlJe
mPTxXOr7UFSNb0+CC1BsDINiAzutHMiICqj6Zka3IkFV5jWvDR7G5437qQdLMmpwq3G492YOukdC
Od0fnEXa5Blu5ixurZy18IwwdeKbTSve+9bnPzjRFe+F8OMMqkcho7OFFCBFdHpUTBUmuhxjlsDE
v7UuXce+TvsdAApNlKf2OWhK29dT6MaUkwOH2dscyuVVIVIfXUsiOohFXUTVOfgH5PIbDkjMsa46
SIRbFO4nxy9kEKMxR6MmmkTKhQ1lgcE6RT+upm79RsVjyCcs7Yz4kH4QELHr9RpBk7UZO1TG1pHf
i37pomKQ27nKnQ2208TIcxuwWFGKryWL2G5mN+18LcT5YU6xdridMjWRpCcHxn2VVh5bZhlbW8NK
j2zT4IFjBlxTyTWX4iXWljF7JOfC3NCYH6nTURtc7LECqxXS9FrOLidzEiQDx+8hISBzdeB/RmY5
9EN9u5IR2eiO5EYhCOw+Dtr4H7/EymSTdQ2gYQQ0qxxWQZ0z0uaej/U1r6cT5zciPWbcStHVUlGo
YviFkc4tO35eeDoBs72y59GrjfjokxtPpil5wN7bkNjmBGeNhYJym48g4hSLoYYRoqoPiSPa6uIl
lMZhtC/VSvPDJtmkSn0RH1qU06XGSNVSURJ62gSe48B8NPrgq9q0WEnV3qJZD27tO2x7Xei3JE6e
bSKvTstpSTiBYd4T6ooWLnqFrSMO9e/XlnsMO5vjCmvcdJMkrwyzqKxkFbdho1kCPj/NBx4VK9Hi
Chw08Wp1FuzBH/6s8uTBnnrlImjZ1ak2TvqYLZETA+1GNfAEFN4UuxnrXrf7myNxS7g9toN7t+fm
bNP4v+QvpKNLN9u1kyfNjqwN1i7BWISFH/+X4C2xAVtqYyU9/6JUfAUE7lQ6Gb9vg6A2KCz0rpON
GIzDuANCC/fvbng0/WlgzEW8yqN/2QdLEk7mKkXo64GtPo9hXKaSdcWfhTcNxctq7uetAPfE8ny5
nNfO/aRQ/FXXnfhCKqDJ9OelSnWIUciScs6DUcTEgWfTQDCSBGQ/QzTBg5mjZIqcfErWUxHO81hl
KLmFqzUlj8C5p9v4vJk8ziCaE71ibH1XbBTW94Xf6Y+VOTxPMxwSEzqvzxb7PEJhIN+PcyXEc+qO
2QQwkiBDj2i3tCwKzmJ/qLOC/3UfSj3cVrMUDHAgT4Mdi7H8Lpj+tHCl0XRh3nkpQNy6GCbG5Qf9
5eOQpXqWXjOIHVU163lcoUT7K0I2Pds0ct+QaTrS6lHzAms/GBBocIBSJIXU0qnXku8aE9xu3vUL
2sO04dw8OyHga2QoQG5+skr/66uBgO1i3EVpbdO1ftvKhbbJC4XXUMcBEdPA+s+ANf8FGzefSBVz
d4sSKdtRfSqBz4wj9C9fcqQHXoQz59BNDX+fiUJxrGXUx6ADiI7h0FqDOj7UlDCWjUiPKUgPo9xD
GgzCo1RXYZlQsymNlK3JrP8Egw6V90VZsyPq5uyfgfuM5ZUr+LMvYuITC758hMhLngzSDcAe+5kr
hBjdAQHA8XwyEd/NYl6ZzU6PjnxpDFmltsMTthOxkK0+H7wNUrVefhDtqJX1FId8bQWjbLaXzWwf
zJSXqYSbnn/65c6erC50ka1mQygxeMRKWyGrObgO4CuV4DJr/kmxvJ0DMRS+jBBDwe2IaSpCNWYx
/KNsCy9p8LNBHZtALyDHOs5EE+pjfI5ZoLLF6F2nP8kqfBhOtmSCZY1olv5A5gPuroBHnpY/UAKo
QtKj8JmINENiMomNlBlJMZzyExaOMUTV4nN1xK1qY8+JL00HkodIHmvGKI1v2xfvpLWYpVEiPE0a
8wwZ9VutCGepszaBYn0zKcS+RmLxT3fd4ljODs9M7ZcemPHXVUiKqG9dXzmtpipQjaT6Givv3Xa1
RZ5O8oYeZfPC2OByvDA+G5RXIIizlwl37/jOlVN/107E30/Qil4Ankx77jGW9Ms/73+CDiuxy4rA
LjIy2rLZPUPz9Q2Rp/rUMHPEzEDkXHB2M+fg6aG1LujxZ0PrWLG5E2h6t8OEl+3afYIdAsGiYUHs
+U+h5C+fqFiRYs2iV7vkClWOfyghfI3CAaIT26kZimIdDG3TzEhVwPKWkGYoJPliXZ3UfAaFcaYm
RtedWWJkf5D+7MQZHSQr4PZxcMGE6Hf7fQfxYom7+Z5B1EHKRBgVw2cOHhQE7qSrYw+sJexAdsC0
MpQawyf4j9qYbQMDxZXmYgyCLLCv+Aut4mIvSt3d14r55KBpuyMdE/kLNveRIScbKL9lKH48OwQG
JhaC9RtOMlbvWEw6GDlXmSqu9Jj8rv0FclWkejoSQwROmSsYyYxyBJgFz3uACAFnGvnq0wakGhLd
1GzsDFvpAx6q4ldU0DEhj23jPgTNxZcCA+4Qbz3slU35oeL77QbWociWxlyK2SUSWeyRJvW2OJ/h
yw331V31I31K/p/Em2W8Ctbq5HUl5CjDCwlvL7KQKAWZv1uTVYtp8lh3dT7Wl18Ro8IhC28+QCCH
m1QeHOPPiaVsEU1mZRwSt2i/ycpjNLOw7o2anbIrA1R1DNJ5m4LxU3eLTDdp6Kn8MDHgjVsMORQH
j9M2e3GZXSjtTQ3J4NvR04VoWwoU/ETWu1du3jxAKKxIaJp8QNMsp4+iX33M9XDYtQlr7maoiI4I
tvmZH6HRSZF/TNRk9d0fYPvYMbRrOfPevnaY5Xbzi7tdnVhSqXHbYvmMumnmOcafNybXJg0CVNTQ
4eM+HE1iRxqadufQa90V6LVTsk/e1KceXFXzyNk2bQ6xQONvJRwG3eXjAOXt8wncRbyuqUPalehm
vEep0upMgGLLoHG6VDZon5aPdoTmKgC+RQNTNixKpfIe2XKJLAdCK+H/1kGiDlV8EKyKm1uHx5jt
dNKJ0pJgUiSytkYtHOwyybYXb65iJ8dsVpwoOgsGB/DstoZli49Mu9wyRS4nwiSIqiUv8W9J+iKT
VfGqvCizEHo4evVHkW/soeRPscA2ocjk9qBauM92HENI7C9krUa/WThCUHZR6ayOd9IJxqkSC95l
d0Nrb9eMae2+HEOK51ZDupOU944nLqTOP8R7QJA4nrBzKfYDu0erXr5YY/KYrTFABWy2btB/V2eR
suGyoQY/WUxsCMrY8oIoHGZ1kQRnhtx2Kt3wAYCMFI0YcyvGfwFpybtfNCx+pxNpi1LWodHwm6ym
fOE2u2DdDxdnUfrL1v+UnIqJOi/Hlw0Il+Gti4F40MFZwEcmkU6ie3DYC5DWfqCY5bjV75rFTij4
vHoHLH5NVVdaAQ2QR/sJocUPHxrG7IuqmJR1TrXw3rMP4Bmd8fO/+NUN467QXvL+oczKSlSBnPB8
bXUV97e0bBKBfdCQrJtGiiERZcwCMmXJosSplQL7A3EoTOfjT1EIHcW1DUdjszL26yC9kA6QSuYr
ZdGNhUz+BR0v26KPrJyhTEuWPEbYyeU7RE5p2gVUvlnoEZN1m2iB6UQs5xp1RmhZ2a4WOj90OBNm
PzTUyaAMixHqyUGuJpa868NCY5P2t8/XYTakj7AgGVTKJ1G7DQ4JtFWh1LNMIBGjzKya4Oo0nmv4
ggEmHuWrbVQ08b1ThFwsXpvtpB6hggHrSUZ4cZSYiEB7kHZ/KbAlSHCZv0t2TVV8wP1WCT1Jrtqa
TK+Wj/KPMNcO0LH3FtQHNy+6O0ZZ9eD4z4utk1sECvvbjdU+RqA4ADFJzh5YKM4YmWiqZsdiE285
xJJu/lIhQLvzxpHIAsY4kUw0wo4XUNpmMq3Jh220sA8BuzR/k50/gr6y/9Je3xA6KXJEaGDL67Vs
YIVIKvdIxvvC1Y9dBdAbUk89N0YYS0Jd27s+0OyYvypvUOOwkj8p3eU0RcmDCcmDyVkEgXZ/LqhO
n0bgUMQ6t1Yrg9zD/VOAoaVToskEyFf5cJcT6km0VYLuidB7kYFr8dsjaGwORkPxiKY3mUsFDwYM
P1Boyadcrpjt1IyunLfSKKxS8y2e+Zo0ruYKUJ2IuCM8g/9jDTdF51rVLHR2RYSjb8XgZXxgZNXU
M9Udh2lWkEZcBmLN+56VekV7YzhRyDfSrkc9nhJUeocAV3rUUz36NKihGVlyE6jTzHLm4+TEpOIa
6wN82Wj+6JAyamxEO+0g2VkObMChdmtCxIKyYILq0D41Ovw8/5o3lStlCcq1DnRtDV+xG7gvWjQ5
FwjA+pv+ngAaDDGqSvhSSMP2At8DEtF1Y/FnBFENZQyKnruQFOGc06azIt+5FFMXTfR4DcZq7s0j
mRhXwCxtcDbaDbmutIF2Dv2XXO90sypIsptD3s1ayql/v6gBl6mHd2KmtIMN9kcQg5EURPkFQG5p
Vbc0qoLJTB72tBnBdbU/ksRHhCwb1zbzYC20A5oSXyZonz7BLYG1mDFEJSyTMwhpE4AD0uTEDqs6
QszTMSYQAvH68o/UePCW144nZh33HUuAG3ObFghJspfgc+zA81OHuACxa4Q7OP+499ynmFFXBJir
7WNaewzntVky+AHnEE6HVmD3roJV1fd2EWN3gXg/0jSxC/7sD/qwDHtDI4nqae7A/pkpEPs3/94G
PE3GJ+2musIrP3cmBOwXO0jS1jGrepHFSg3//ha9HxT2FH+ziwX3jwYuvZiK1WZwrJenNAidcmxF
54DmQXwvUrr5Hi4XfBeKNhW/ILBDLuwXxZWi07nZ7YfaUTtK5JngQUS6Kmf9TuzvovPa8P4NULIr
cdrYYg7mDnL3cOe3c8RRTjCCRpFpzrVFVurOi8D9WvslWiTy61mDEwDob2k712tWQzjyJ+A9vYZ1
s5qPVBgA2ZBzUf+HENtUxZuH+ky2TZ4q/evx+DvVASAoQyEfWvtv+Kpg2bQh5Dua+N+tcf9UhpQt
WScoG94MtCspBugcmJLm6dfUMA+kOvE/W2SWIFvPEV0V8FC19xkuVKmezQbxcKriF/TmjpHdrDDI
egdEk0tD9BHZKvlL6WBmNSn2jUKpYL9sH0VgMujLIb4cLbTmPGcX6nBEf3KCS+MTKTHBZ0bNaMM7
gvxEaZakw+cXY/59RX+RvUWKFO2O2/EH4txaF26yraeo3WRsngttlejOzdyLxN1NZIxTrIKnafmr
yRjuuO33M/ols28sNnduuPzhj4WLnY1Kl7F31WCbN/0Q+kuizr3+lMBDU/u4nO84CpdBZhDtU+mJ
Q1kiGaOuA3cxdCQ5lKkkFqwgR8Z21M84RyApMWF74sSNuObUVTyXhbxJ2liM7d0elq5lBOi40wZ7
cPUL3kfvaBhbr8BYx3MUoQDCuJAGJZZNeBjzmnpPqMxSyUtR67Tl7gdLtDmYH6x/XTPu81oxTQHh
vXTmwJnwvDYu2AMU6kvqEzRMNbzYpmZ6KpGb5CNCyXGwSnDppx2V8rn4ThdneCMqW0d5GbGOzqaO
/Lg7WZw9bBBe/a0K7BurOSORtHMsHoaF3GNUQrPYebBhyUeT1WsaeSskD/zPkslrkfZtNvxm0wAq
SV4Do5ImrX++DPHUgBsTGFi09epH4no2VHbjnzlcDNGCQI/b5H6k1cUm4Ja1JA2UbJMSdylIaa9H
FU8/vnOadfNiOs9LzNPfpBmFPfy34KDK7YIrb8K9Meg8hgjSKp4fbS5X7xJFfMQlm51t3p6i4hOb
2r5GLwotSS711iGBlrBAdYkOpd6Zv1rn+d1/AN/rSoL9OXXpBYlEpsk9bYmS+eP9d3aTn7fbF9sh
XYtAdIbz6XoE/eRA7uzhZlJnAZCtgj2V8v8bV7xXRz4cJYUHlDePmLCGfighUlspe06wc0izlJwX
s8drw3PIEosbrGTMHJEQXKPd36eBkpNnpdoK4ZVa1CoP5TAagu3btaH0ZVtxqf1C+KwzStcrGtte
aRimY654WmTYvd54HRbkIQrnVLX/5xNcfkMkVbSOJ9Gk88ExvpKpFao+RZOHC8IQHMt4loHF9H4z
a5HZRwW5qPmsvWQtfSDskgsda2qGTuYRl0ibe3yLPVgNvQ4ruY6L1VG4uNDJx/6Wy1vJhurSiumb
FIkd9fIZXL5spoj7c/dOtCjfQj3nA7qri+rP0ILHvwaQypgGTLhXuX5fh2rpez/cTgODWfrTcHCe
+aoNhfcpqPwu0v7b3w0xyz8ZYmxvw6dwX6dFTPEvwf5s6JpgmLCcleteaO3Wzah5eBYkRwl8pDw6
h3FOOwFdkkuUB7DJgW2fZdKfMRYdvTkQrCuPHHxlQ/QflsZzS07wC+8KHNvYa7ePUMZ2qI0dQb0I
oYF36s0kyi32ARG9m2HFNrBl5xdv90kidZcKU/JYpXocpriWLj/S6yjMiq+MEkwN6zYjByuCndxt
Zg5jx7OUSgpNm8jC9N8SaAtkF8w/uZY8mxpPDvnuT2BF7hwkO7QdLo7A9BCnts4bfNMfLbW6BXO8
p4M3ABH/1cAECaqLcQgKr8TnZQs+TiFVwQJESDUr4eP9ToACyxPFcaJeOQ9vzTelMA/VrY8MyfvR
x3v4MiJSEj2oPSZS9x6Ls1CgiWeY0XDLooUv5AEmUPav8Xv2FZ2jWRxrqgjnE64u2Vx8sjZC1Rj5
e9jiL8ki/ovP8PoAbU8+eRcWiEgbNfX2xEVzWx5+1qm+OpW199HOwBMEfCtgdaZYjcPb4+IuB5Qc
MIo7ZDlLA4pHhlU6uGAP+rTdi7EFr444TZXxXvkkVspu5kz4QgrswnJNQLQBjMEWV7u2RaeOeo8Y
58JtpYxdOvCEZUQuswt+BOQeD9hJY/irnxL7+AVJAidN4C6AYnIdnjyaXpZcCx6pprGr7pZRBTuW
nfyX364AoOT9HHRc2gk4v+TDA9+gNIKN3Htnr4MYjkYcWj3iV7NajcFCmpbtzx8rPba9smzYcsaj
D9kxNeO8r/h6/f7IlpK9LtjqMApDQVW/0+V+yPrm5y/U0ERpizqneGmUIMGfbuaX8xGpvauFROWA
ZBost0x+g7sv8KjIktVUfDK09N+j212ukESiGO2guONN9hNlHESoBaWaolftBHGqKI0ZIhN2u6py
jDRrt+TXHwtPkKW4PMi8aR/zPhVVx0W0S9vnq+kqPsANw0Iomls55TJpiNV1/Pzz+QGYkwVx4iKq
9OjG+4gQ8TZlmn+XYzYE9nMlCOK0B8881B3d497UlYQdbIytFIOLueVJcvsSUrvJlqFrEuJgac76
zuetIUcaeBJNibOZlS4UGjMKojt76dhjNSdFJSQR+SW5leC/jAOpuHzZ2xC+4lGljLQnHjaT82xZ
ycmPbr4ZibdRi9Qs4fNu6wIi06eRG1zbq9Tn/gxfevi2xhPENYb6a4PrCtJJ46qrIosBWiF8hvlC
R/kv04uxv39V7Gti0tKpJ/uDsai7r7XPeeBGif/xLTKhZE4ARbt5jNZrnhuikPgvnGFJDwR2bRpT
PT/LCe3xfJOXhJ/sUXUM9CepRxe+nOcXpG77RX/Lrc2gZRMmEfln4BNOdH9KHu18cW6+bBqUJJE/
LrZsPQehUkE7lVs1xIfXVYVxWuyHAffW7YDRAjL5Obtlolj0TznLJTYvBRMs6KUR+I+YHzJjshZP
OrPVfQ00BxqNLBOAGc52VYTjC87qKx42N4DIGTBIy/ezbFAYOlE1KeqVDJM9xmkphaRWIQVc1b1m
5EUe8D9eW9wQ/ZuEIZzxrgLU5MhQT4AfR37ExF/fcJOo7jDRvxgfV91y8t93l6fapd0zPmcGQxE0
fgK6nsNiBpXaR3A5FoCJ6vUkIlqU3ZvLPPDZrcPxKpdB0p2LEd/CYVRhRHxCaeqm3tXdWhd6T2YT
2AtWsv/kEsQGb11exZzWqWKy78T56gD9ChIqh2raK6ZAgvC7cGEbeUkkx5i6R097IybotSp1xVv+
KGmLX3xqjniaUel3ONSROqjfsE5ZHG9Agioq2WI4xceI/QQB7+qXaoNJ8yl6z7sLDkn/ddz3zT4z
SUiVygtEhrCIAsF+pjAfEdgbEIyGHum3GcFv0jxsslAL6I9rHajKWxqlpJVyYWNrmfxxlJhmwN7E
ooEhE7wUQ6uKHWe2cGEMkF5cLrZpea+Jqggp1Asibr5NWJuqNd4luKg7F5/HyYDPl30jAjaoWYwk
EJexSln0/Hysbfh4PglBdUdsTHDwPEexIbJD3beukNVPhud549DJT7maJD+Fm6oUGqeG0H6YVW89
JdTBEYyYuU78AAQ9tkAyC/CUJaMFK33MO2uGj7ejySK8x9Wd7M3e4ANj+oBxrO49kMGLjWqO/Yhs
UXkacsBl0o0sK01frnFm6A9QwgTwH1dHYigXEagX+MXD1abBzjxICD7HfXeCwj8BWGM8YAAhYa9A
SbYnPbJZMtPn4jJm6ZuDoVndU9LXpnMEOa9wae1bDa5/nbMOQwEvwY58g54lnzb6+2k20SLMvbrL
fRUa9hHTCvsZI0UscHW+/sFc4AHA1o7KRhSrzPRc+6R5YhhIdQUHqc3dzYXdg7H/G3GZBFSa40jO
D1eMW2H5SsVXAyHVwLgrVsQwp8MOdPnoqR5PFTk4RsRS6uQfQCtlGkQ9mM03PZtUv3jBDc1H3EgE
PndAqEjuMuVBIxL4dqt1jF1Rb/IOO8CGiJ7aNktaO3QujecQwdWBGiOpujssB0lUQZNJDSpAGB88
rb+qPalZv65nm57kXrU3KIgow86HWt2APxu1fXtiTHjK2l74UVBjd/zm05V2N+w+lzf6klX8bW5W
nqL/uCJJOGmqhgMil8HHsIdH5T0edSsbCqfxCNKLL7HVftYoI6nJ1tojeBaY3OekpARgXHKpOhsi
Xyf4L9h6rIgPrghaGE9PgvC6vO8lYQOstqtyI5w1UyhSYaTWUWFhVrzhJBfv75T5kk5KaGcwY2u9
ddydk/G3/rYrhz7RiaiV+CS/OJPNELkPTbNFIZwUwqPgVAZLb+KLkoPaEeqzunziw2xost7AXHFX
cHKzSBBWpV0TWxjSKP3M2IxNV75V0nshgPyKPNqxQ7/dmZW4n2tX+hkVV0PVDCx+GkD7tfRmmgPy
Tr6727XcXG+UF/OiR24/hWCQeyJxHw3T8MRAmGJ0jjmM/Kq+fKdsftysUFEW8R9yt6lJlAeWPBjV
ji/0ZmVkqeGYna+BgNrKdavSFJyCFmAln9hvQIRVCcZIyBQvgFxAKGpTYx1q9blDs2joSiDUiz1/
HkiOMfZ0rCUF9N+k5sTvW6TNDGAlnAsgjwOM4SZSg7W4+ae1edvXTzH6amPZQfUjUSsvFaf8JrP5
1A4yg56FWZ4c4eTZD99bZ0W4BpVrsne7wUXfJ8H5tK3j+046RcGNYPZHzkmNakkA7SA3J++pbFci
ECqbl6LSSdmLsrihosx/aWzzt0Q0Gw7pOpLXb1+SjZWYNiAF4g75vebiwEPLeJHjhUI4kr4plIvQ
Sx0mRrOxMsakCQWDhe0xwxUxf0r0J/YI4kHNift6wjICQXVEdCdfLekBK5i+q1kjgQ/n4yKKmImN
QKlDS6XanMw9TD171F4LEQyx54lGewxZ2Je3Sy3+PvRhtNh6b9YXINJFMU9zdxz+DninJVTuHGup
uxYSzuZoKrlkjGJr4gvKz24rXJ0LDR0DG8WUSO93S+77Cj91yNQzzdabiz/8VQk5xAeAhG5Wf4tw
l9MJQvlcEjwMla5ZI8sOpk0p0novhKHzxsiVwqe2DUypPsG4NzMnMHz6vDNV6iyOUkHDH4y/bLNZ
I1zDHNEpS8Q8jFOL7ezozBVdH7JuICip4CgLfOTY8/RSgFBX/2fzGHh86xyFk1K1yGXGB2oubRIo
Ki8bPFWzPbOqo4y1n3x1JgNCnyX5e81hLDVlkJ8i/uQ14cd7BPRMzmlCuam/ormPw6KQfQopWnNn
Isuf2s6iqzw2a98lxWyra2TC805V0H2pUfHlqDSm9mUmvG9rLvsMQVtDpLTajgG5Xm2teu/4NmKC
EATdy4gu/vYF0HVeDYfplfHj/tzxzazJDIM7CB1TZU2fyKLXSmQ4i975kJQPTdemoJBoXLwNqHQt
YMmK4+yaxszrGZrVy5tkWYz0BosuiXP1AX8zeGgIfLPJq6ZSVsruwqV8wxRDAWcfTF2ZfQCn4S/s
69h2R64jHwQz1a80TR3yOgw9PtMb/LhRMxpqgr05wcshl5H1zydd2xADxJBGDdZWFSYHPvRdaEhW
UTpw5+amM6a7e8JYBaffpiNRylNz8jYcXVjgbmnjI2ADb/eP2WRAwgGNzTkAUdt1e5odLLV5oX5N
1l3uaqMI/g2BD0Cu19R9wj29KmfFHBG8LcqWqOcIeMx6XW4cY64u+ceIa4XkPobs06xEgHi2rKC4
ekgq0N8PEzmYb+naI07eNMDWXPYjVV+PzVEQDAxjRNccdoxrJfbEeyNKCljDDL1FF1oi5oRgtKr6
oo2wXXaeXODa6AnH8ypWio1ZTwoBZACIYPaA/7dhnlm01FSbmtUmRUK3bXcstXWJXil5Z5uW8Qng
xfsVR3ocMgvHlDyoEO2sHcUNeOQlHaBrXxX51VBzRD0gF5FaRCR7UO7SaS0ixGIDKv7hhyNUUQdo
BYZC+qqaefS9MWcB9JoCFQlZ7ZercnNGRmsY00iHyHtwFaDBJq3S5/u1Xpy3/e3v/Sl7ba9RFzIs
KisceQm2DgG7Y06A1hKG6S+VI7JWHJAQNza7iplzWeqcneBF74pbyNj9gbS0fUvn8K8yyhOhuhuf
cy6UxYY8M9U9FzbyD0Zy1TXspxsxBPiO1e9/lbDpN52FYyLtUelnDPVM+jyuHud5rY1yr0TI2Crv
IreQ6uffzKjqlw7Sclkd3ynZhWZkOO2LMgb/GkQal82aaRWeQMWyOWAW1Ry1pYi+mK3lUwVPB59U
ybc5xydnNt1HpdcBCVq7PEdWTz09aeKSRjQbPC8Xv6TlpDTl95JoSAyCRKcL/knnzdE2kPKDZuFT
1+07FIs8EffcnFuN7QBKYyzC97Sf7cWSOzNYBWE1xHbOjlxwNlEysdWkCS3v0X0kAgQh+dZZFTsY
R1sO0FMgoaxm+UcdSzHIMJMPYHfVOSU12lhGc7nnZJ2DMyEU8UotFH4mvLr0HT9Pakbqq0V8ZJSK
noR5uaj0eoYMdi/7YxBMMPW9mI8aPLZagsF4QcCvcp1z8TtQ6FmQfNfG8+IFGa7kekmsTA7mt8xB
BQRkgTBCeuwCpiZ/a75A0bCMjIOvlHoLiuRO45nPSsdQ5z3O0S81fJW/cvL7DKxZcJFomIViscXz
VLVUYGhXROLQNIOuyy3owWwVZIGD2rqNRadlUFYrY6CVUVJ6FhOdLKxfVE+TXd91bxuuPciTSqNC
nbTKuDF0fojKhqEj3xT/rQyaX0UuVv2tYJc5S7YwgMs92uiuornUdVYGZld5mY1HJWPuFZ5jJvOa
QFAoe+/G7zY/SsoJ6KtTJ8r64z8pHShxFQIGuxe5pYvN3J6WZBBjDX0HNrpPdZr7KMdJd563T7+3
09wK2ZoJjzYh/jwtwqc6SIPPr1uV1bKDs5FE5r0qjggoa2OKNxESoYRy/XqSNPRdWMlwoad4scLg
/AE+O3uV+LlhXlfueoiXaLb0guv06uM79kTkgkh9G/WSorzQdu3nJwGiKZJZm+aq7X7R8vfQuozv
b8cUxrBW9lmLJT3Hh1NR5X6c3Rv+1vzHTKUjZDzm8I5j6mFSVftiZLmyBup6cDnFBgeEQhpR0N2y
tijUluKU07/JQnrf0hvU9wrn/olGrE3kkIBSdUIz8iZSIowD8E0PX6naOxl2bYlgbpF9fdfT+xHz
JMRUXTbHW1DS0/Rvf6itC3W9eWEFBWN0OcrwRDRpBzWX8SGavNAMBTw61NeID5LAw2kJZVUe2gAH
jGscvj1ERCGJMKJiqtcW41l1h7jhufj7WzMjSfA9fa6t0hcz/BCNdDhJNc5vp0scmjvpg5+BXXl6
79MJiXChPCV5UD7Xj6CTGjcWJMychea4vNNqc4E8j4YVhmQmIgg22uyj2LJ18YOi9gtaD8fm3YeZ
idz9K+sjTRH3S/YUqlkrty/QivZCcGWkNNgx8EUuEmwn3nfVRgr7Y8mTUORriYojwQ0yJv6X6z/e
rlZfeWfbCZK/k6D9ajPK+IlauWqjF09rUrkbVSy3fC5AZ5bzDsTfHwe8J0KuPK6hFLv7bNALy4FB
C8sRMMITkaILE2SJcR+otqAI6jgfTqhkuHH8UcTB140cHKxkVou58N0F5H7hRgyYVzQ/3Q7FLpLF
fLD+FZJEB203FCyowo6xns9LTiv6JE/lqp6hMjDGMWzyi3YaM2ZXM1TgN3xKRZ3z1sM+f7tPNYTp
oUKcGf2hxaikWtPNtaAbjK9Zgi/ty+5r2S+5cm6z4DC/AZ+WmX8U7Z2OS+qD8im6pldGl+QkfAn6
QZR8XcmLneFbPSD1GrtvNJH2RLrmImkTwfKguQB2MnhoF1XIeD05y78C8DZC5uh3/ZpJZz8lG9OO
SUWNUZCuj0VSHhBjT71Bc9V8blKqq1q0kbL1zBq2sq6CMeqz2UMBn1xM+jvie+2jVULnOFfLpjcU
2AilGRed1aoXyfqV9+st1sqtkOI5IOxR0EIX6pYfXX8VCc8d4TozTZBNyVpCtWM3yl064HCddUGQ
XlEeJPy5uaN0IX9SIhx7/UNo0BMKEPz9Ts/9Pnxm7MRgZls5TISrrPSybAuYQ6elF/pGa8VoHa4o
QCdLm8QNQghN4yQla4TiWrnlaxjnDfnZDz1SUN7SC7oEL6hGhmIKB5OG+gNM5sjdwAM/PlOFHTYs
O6hoONDk4GY+whC751PqbRa9jzjmqUpBYNCFcT4MUktPTkRIb1M5mkfanWkv8Ul0eemBcD/rjyyR
TjlXZ6wPfpKOYTYcUuHsrIxBkKEqmAP2IfLVCEERtkABmlBG8G8Hzdl6z8RWNWbhyav+BdTTKHP6
KV8NHB690h1tgvCxAoB1aghqCS0niiNPc4fO/eH2iUYxeWbcWOLUVt3+3Qv+3AaajbWqymEDuMg3
WObF7gFR3p4YMawm/7iQ3OVpl6a7qhEgZYAJSZpqVxKGP3uLUf9e67kMmKQfdleNKdh65h1K17Cm
iNu7yuvgrH1UfRRmtXtZJoZnUPVRiQ/jBLzXBWff7LARxCxZB/qjiLLV/IXAP14hOtJf1O6VIWgR
qqi7KIBGt4XXUkjVEu0OYpRluTkvK2pNHU5wkPL5tdoG+3EkvKWx9on/3ARVCQWXHP3FJLO1y+ZW
5d7TEaLg3DmGF9tOg/NrZG2Euc0DgMhsKypugJBI1rmXZFtmKuxpHxu6u6bGmqSvG0+VU65IItP6
e3mkPoWr1aDvKCJfzvlqx4mt5qGZw6051TjThyem7Yz3gfOBy6t679HD6ERSgRbK4tI+f3rBLi6T
K6vrTXlXLZhFfqHzdpEp9N/r9C1YTdTCd0ZsktngULus3l+BVwVikMCH2KzKH6z6SyYEBgxZ4hZW
XsN51mpGWSi13OIkxaDCt34HHDLLV87bgtvmCETsucM7qB11pjA3/+9JReXotP73oFxyrUqKQxgO
L5AvWEYL5PKu521Ls/sbbvkMes2Oy5f6qMOSm6s9Rw/T6G6zbSbFbOrZ2Kfmh28JsQeQLVC060T9
/yOaoB9J84stYzzB1D0pp272uyHhyecMdwb9L2oGgINLz2ct1shHIEUhYu+iCFCM7r6GNgq69CBb
46sZgGLBbIk3dZE+8+INBgCXEf2CyiGFXmhbQXO+5Bcgnx+T/v8Ryuq0hkTrN0QJyYfKNhmSlh/z
NJBayhrsSpQV65aEx/9DlpHoEIaXQnqjT5lWtBkU2S253tUdoRPt08Stlz8KBNZ2Y+PwBguAwvUl
f+5LHRZSPr/O2q9iOuWQa8d/Dzhag6+Shcu9bmhRh7tyhzteGjlaiG1V0csm0fnXRSZpGcd3vZje
qlCxqhaWYePIc/l28oImSX/qH4mwCReb+AruM3nqGvHGVAMXFvOXxAgd9yI9ZAywsjZr46KHURTX
8R98oLW7Azeo7mifmhSczsTr/5N76A94Tfyf73uNrxFvk9y93AN3/iIuVky/w0lXYczsNNcgGxbF
f+PfLyaWNf4lB6WRKLKyHmN7nRsW7m7GMXKSOotqhlmvUrV2qLqJeZehAuHsWlN62GId2mSoQJBJ
G5qsETMzTezbjsklRzrLpfZul4Z6/JrOG5nnrz9RculaxEdBktGWCgLdVzJphy9Qyp0p7vYPl3WW
l94QgF38hpEmBLqAXxxV+YgHqKApnyD6J3IuCZXnnvrP7hKhBxbrr2PiukZZOLcOVJckSX1IEjJn
B9l/1SP/zrlQ2z2PReiFOCY7Omsxdku+TPUmLbLoobK+TJLmbFmBntbm2WYh3W5jtAYt40umwoNL
RbC50bnquraXEHgm50TLZIhP6ZO4PycRFwg1VyqM1eSfZBQ0TIJ/jdJKIlsimJRX7Lh2qv66li3Y
6I7lrgEFSvWKMuw8YVLdMoMOh+6T8QUAsksLk1pSunmmdLTSALzZcSum4dBkRuMgK4k9Io3/t9jA
m7bG36JKM/dK9dr2uwtt0N7vrpBJfkdlDDsDr+HemYc62Nr3P2Ew+S/pGI1J3oQdF++0ZOkBr4fq
ywoL9EM6ibFL0Q8lQRonb2bT3GU9XYos/gHgohzUFY3UneyIr/mJZgedM7fDQQDhcfTGHtjSGhvU
28H/yJiYMtLMPTn/lCOAHUd2Bobzn8XMCh0Ne72fAf4sFidXAU6+Jyfz5rdKyM4b+HVcZGq2hS+a
nvHt3jg2ZKO571TZtE0peUGzlmHep/izm7kmOEIcFHP8RtZHVWMVoeFIY5FbSfD1P7RlNjuclWwY
5K4PR+TrvTzEznvkKCoYdKGz5LZnoTowHgG350byfmBFRu82HsRtMdyPe6owHwSGCq4JwpHcESww
8irRAr/s9sqGr2p4TuJuCMK8Y2iAnk7WeE3heBvMOk9k+gghUmwSDmvECw6S6IMe9C1ozPqxdzhH
R+yItbmxrpbwle8XzTYEQU0vtdIkkGZ06y5XGH86XJbOl45JBPpF0cmX0tY+1NiH8O7HpInYZV7O
xJ8fmg+jjxsbvjj5unWeP3nWU3ODts4QPLd0FpWm5UWq0sBO9J1ASY2jereDRwbFripUFzeZqT6W
WyCoLkdAwgPI6mejO1B3rz7ShGvVQJgDE8l50veiWzjK5f6mWx12cmoRiB8jdDmJqiI2l+2LqUlT
pQQ00HCf87QxpjXPo6FsodSgmE9GYRC06qEvHr58hy/8Pnccj9Twf8wQ+1X7wAn4UtxjYp6/J8Jv
x24UxzDjFceJHMhYYO9Dc279b5wE5VyheJYWt2SbsI7SdITweKueLE2/ZeiqBiyBAxf+ldmfyXk5
wM+tOId9GRnW6JrUHdqDBXb8ZFpL4bzDPr9U3M797q6VQ0mR01WmG7709km9F2G7QJtH/FO3dFiG
BwEE3uRCtk6RhmpMoVtYp2zCfHu6/2EvqGz0LHwcffPEDTCnnC2sPkEol+ysekypI4L7ICsRRnB5
Em3rqmsNSeiENxK37mcOmAQ/QjeljPkemvDk7cfm2lUgGY8Q59T3kNhY21Vwkp7spqBwNIHUh7wN
xf5pbBvNTVr0yzcpmA1PYN/buNwiVJaASTg3CeSa7aSzEyjPIs3oiik9uOoDMnHAT/iI7clC7u2A
FM05zCfu2kM/ANeP2AbAC4rEL3ulxNAGhqeIec8fLRDOiL7ZNUgEk8H7AZBzVt3Ic4woIWn37OyR
bnz9byBjeixbZgYOXlT6JF9nTt+YFf2htaomvlPnagyyWv7EnwU2MIPmTw4zMSIwWqw9pbvkrpCF
IAB+UkMbpcCQ4qbJiieLm1tAboSNzYp6XXkNf/bGmIOGHoZ8GfPOeOg0+kVV8hrLwclwDKeLPe/C
TgIU5PkeydfHdWfngjb7Di5iq09Zh1Org8M7fu9I27I92gkjmIYlc39fQXcXxrvNOvhXtp3/Fq0U
BIyao678xd9dtKE2MeXB1FmQzwXDW/ulvSM76+SYTHs1MZZL00ApUtPbfiFH7SZ5b3sOzcevPt7W
P/AFRm+SeYgPinYU44Tw1vEUWmf3I1TsWd/1QKCIrkwNEb1al+PmIuHvIHq1UEt+pa+Cw8w9UPyn
czCqhA2XSASMIGBmvxytRdvx+sFWa66sEzkVunh6Qs5sv4p6IfJXHh2W7MFFTFKqAoCiyt5s39t+
WMcSNThMeR2NdCq2CaNwNKedTWvADBRlocifeDfwNY/CcPLB/gRix9srpennq9AsiQqMFTuWaCL2
JFHBK1SAKQKXZD9dK9qyGOxN2hbWOU8dENIFUHoJOMvySFVBae4yemsjvNiqovxttTUzzqNuQQ/S
YWGs+sjnCjta4t9irevDM2ZBFPzIc3iAp+Fd+TgQop9j9HzAmAKqzws2xP0hXoz5mBscNhXprEvD
AjJfK9YqbHB6tG5+0pXz5snuN6eNHLOn3YUKTJKkfgzx69u7miwyzZxFF66sWE1DO4yHmvvGlwlM
fmy22zexW6Qt8lrFMt2BnOyrd/uU5lL9gZLLpIp4csF94BM0TTEtPzaY3gFekNrhTjAUo/1TzO4L
ZaBZ2sLCSIpsq7FsNeDp6OofUg2HXQNUi+UmmGWEJVuKKPAs+Y39dtcCHuKrLRb0Vm5uFJ83e/Jm
ldZRaxvtHqQfWDHt2xSNVNitrN45KDFz/G3N8aNKM2spSz+OL0R1R2aIMAW8bm3M779xjM0uIqWX
HpGBizfu7Rm07lZsRBOdzCQg5iMzCzTsrVOU74VLA0zwoq1ZlxWXBT+JIpiP2qdIePfAgTo1w3/d
mA8oyfirabSEiF0aWvm3x2bWVF6LEbw2vQp/2qALnTRZsfSGkrKWyTTcNfTzQv+XgT5FkTHOzdYZ
Dp/ZYO2cSBgopxPahcjzo60pniieIBapSAJ8fuVEjGvL4MMMO9ssyKK4kAzmUYG7o7TsXDu9A0f5
N4FfCPG+SRd2gUOZuW8XtnWoByGZdngCPQjc2SPylRMru7FCezjqZyQzEgrcZhSSZHl3VDI30VlP
1zMeeItysjHZWgtKFmnhIMtx1No01EXK2OUMjC87danKjBgQqts7YmsrklXXBv6OdAq2ecIZ27Xn
QWk/RupufcJFqnlzTW7HbqFNSPWGCuu6+s/rJv81n/SVKRVmFBLYkVMIgmZgd4hWgGPbtRjzG7ux
y9LEN1oAgdt22FdSRqe3gQqVM4CcbtO2D5kf+SyIDHhocl/gxIg0HbRHWMLLOgl2UcdQYQsNkip1
O+p0MxvFXLGt2W7MCbyeIio9JlzkcH6NYCzYK+VfNQDf8U6xQcu+JWfeh0EQi0BOcHuRLl/Eqaha
8R0MKsRhYC5iOqvBqJ6AsI9mEOdSI4a8do7n4QwsdXG+poBwqPOzrkgxoVmCGAfrZyA4QFf/ux+s
AET1qMg9qTxqRwU2mACBAI5xhKZvVxBs2+3tdhWxGbbmgwBDRoeju+arxVzDuObj9Y9Pb+x2ObXL
AS69qLEy2TocSHod17DrUZmyxZR/WB9DeJ2LESdL+NRxbclE8QFru2OSxM6zLgwbTu1ZU8FJJ2qI
4GiWxtoZdM1af8VDDw66tChcuO12kMhXCLsNgH/YjoJSyswrJDj4IjCTdPX5ZfQ6cbbYcW74ZAJ6
gNn5328TQ5ksO/wLB0i+C0stA0T5xf9T2ew4C7rncHxLZilIgDGmmwUBOu5xW8w5CaNhRGm+31bc
Gz8hX0XwYtwEfKv/nfkzw0MN1jLbCuS2xINsAO2w3iHiAuAcM0crkOn+eeL00NCknVJiv4xynlqW
RE03iIRiowU5qDNTDqa1PhNt2JwnZXeqMPHkC46z4ryjG6RpbkUKUBd4fPbD1+BJ53og0YVodWjv
TNZGAO/pzxSfixO6MCesMpsAixLdsGCdY46thk39L2Bj15Qt3gGfKPGfXo3ds9UeBD36lohB39we
ArirX9fzBxNdKcbVgjYVJLRzNGOFv76s/oKQvf2QsyZxLajZAeIeP0XUGmx6ED+SrcdlYjuRLCFC
xpJwe1f5gtiCimi5rIhEYzmG1ExsQA/TMkmNr+qK12EMcSEIDwdp7q5z6gfG+sH+i3D29JgwK8pY
ZxncESTpcYQAl7gSQM+6KQpP3dkwxMWZ4G6jI7zEl5SPFiaaXDp86WKIhRwxE7xFsIudw7S1a7s9
QzWV8t4dk/wmz9VKLkpQw/WGPbOuVJq44UHO1bQ7B5usm94e0lt9nf8/ChAP5XTsWCyuCmbE7gwG
9tCVULIOY0q6/jyjaEX8tZb943RS7up83cLLrMCAdp/CdIJeuXcKu1u/Swnd6nCXakJVoSWGXHYp
0i2ZRgfjPFMjn9yFHcRCrMZcDOeNnyF7G7XtX1g8H1WYWWMUA3XuwClh0PESO6dl/QtUqvTXHFav
QIRNyuDuySC6DYMbF3T1ymiyNic4wiMUb2PCvSl0sX/UAEkTCCDcEmjwiLfAR8KRZ6acrnxwGw+g
yWy/z57Z9wvALbKv5/J5sl4GbokJI4jnUK/+e4mTIcPdxDTSGNcQGhUWkKDQ1BtiyN1VRbCYah09
yobTCZY4xn2+S2RN2xqnMK6FwE8WM6JSWUEsGxJ+bGdE0xsw0Ko0+X2hX1FukezWi4W/pLRXVHCk
AaQo0E7qhgjkWAyAlphsB2GGDbDQispUcLJSgLHnajSqUmlzCtLzcHfq09qe+46eeBhOcpv9E+KF
rGznUJgAusv/EeEioNhDuCLLv2QdTfBXVI5kv9w3QG0mORvsl4AritxTVUyGMw/N1naUE5f7VzYg
8bZBIiuRi+hSl/lNzPeOKC1+0eeGCuxyTvd2a1OfnkiEq82KwuDYvXQ/lvnCLAE1+z9KAB3NKepQ
/hm/HgXTpyRTTudfyStw8pY0yqteSWM2LSj9tWiN+DNbrYhvGhZkh01LuJcm2dUvU4qQbZedBYRS
pFIprR0SxJn0kKd7UhrQ/YLoD5XBLOGbvKfdPaNjUfOraOaKri6Evta6zOpPAJY2CYxVY4KFmOhN
wxPSJJ4yxC6Zhk2TuucEtoJXRHAObniPu38NmYJsuE82Xd4cVyDk2uFhIKVfnwxKOH3qwkdz2tTQ
wUZfc4UYDzVsWPc4w7w6he0Z6JJE2FjhNq8rWPocll33S+/lSABbOSGqB5UecZ3TwZjBE0D9x1dL
QIezpP/RTMAisU+1h4XFEKf70FS2E1h+icZwQD280g79KgwjSK8W4c9G8+rhA5fiRZvHVs3bS9yk
dDtgfm4fyHvWl6tk+xMhVXcNiCPD+38LbzSNMWvz6YtvLDd6QwIf0uJ+reMh8XzD/jhqPX9UlZD6
jd3jMgKDj77gE7c3j+XiW8Y21HS0+/9atYE6UKOJo8vfzKtkjS/BFqWv4OzhuYolhyn4TW6mwN2s
UkUNZHaKGrDE22hqbLW4dqnoBmnnfJZ7gJ4pYeWEc9qGVhm87gRVcXWA1cBQK2NUGNWvnAL/mAhW
7F59Y8w8SFCI1OUp7xLNMWQjFCawmL2U/On/+RH+TXNI/VFrmKcBWIW3CRw/N+BjK200oFtDAHeb
O5/amsSZBQ9AsBJk3xi0DQML+ilQQgkgYzCEFW5WZa+sU2r4cR4PLBKP6pmiquZPBkoXIidbNW5w
ncDEUaluGZfUl/PI+MwouZD0hQqAoe0PTSiqaMqDqPsvkRNJuZTOj+aldj2w3Yp8t5IwzxbasfTj
8L7J01DGM5pmFUJj/wPoNkSYRhXev+XO54Nch3yWhzitqSyaBWvASy8eVqqu5UqBypC6oGWL0qzk
Q9bdeWzBfwCiECz7PXPMt8CMwhgqcN6kuH/vRUj2O8zMVkQ3z6cu1/OuZ3yHGYnvRaFTHLszBc8G
oyUuy/D+B7cU5DRGULC1WzX6VmhYVvO/OS0quc4T46fh6HucQkqEQilz5YCCCsnYgyHUrSZEnigN
kyQ9Lphc7R60XBCoYyCWxp1413L7e7UN7CCI1Tcijqx+J8CWrpPIYbsjqtif0NO2BpADyV3CJPaB
lrQD9AmTTzOPN6e0K69WlQC2CxBNqd+tnYYGFeIne4olO4FkwtRoP38LMbAjSS7CSr4QYcXUxvff
od0GNMGlgRypTUfderu/DAb1ZN+q4OjWeQVEKfx53wUpbWUr8V0T+qBiUYefRxa1fIju6wuarW5O
8sgDH2rlMkYnAfutTdD8TvAb/uWWSmBbcfGhTuvD3ps2sLZK9Zohx0rFeW8XMVTKi0VB7cizeNW5
x7BAdOJUBeb3eZ9fKEjRaRSmVWSuNR1STia2DIyd0RJCPonz7+vBMbx/hkOkATes+MZtimaDBZ3U
2QwWLiOelEhJe3d4pU9R13GqcRUF1qwBb+nP2UOwg6jTtrNkT7fHLv7yrNusE0Tp557vNO3JmAIL
49CiOmDlyvJC3pE98oaa3GhSOXFd87XLxkiejQpnKAbIVGuY9vfqjxRTN4vRnf4WQ5I+OWNgHofi
p0AfeZuTAct+nzA77Ae0e0OgpbY3gNRxdUYVlBTCYg8WbmvyXBo4BcjVQVpFS8DHFhJY1onOEPOJ
uFC/I1XAZpGiv2/gYc+hYIqhdV1aFWhmQOnCmqa40lh5ZCFDBCY29qiQaOI8F5kx5glRM7WK/4n5
rt7sjHaJdAOqYk9ouvJyHQyvwrbRRlZFTV7TNhUjoYtrrGZ0RB4pOlcQmOXTKQW+/0AE03NedhMQ
VT7JBNWEh9fg7Ue99WCYpkvAGaRjkCoHSwrBmYvZgnEl7cLTCAFSgMy97rhalTzN62PoAxcbRcqo
AIjFoz3tmMcMLm0QoLYSsTnZsxMn9P+P983HQNK7rIAxMbmss6UeYiBvYD0WJxh5AcHHiMg2Lks1
eIYanAysYcZpt+Mb/t4rlMSQiFq/JGWLYUOI5uVaOMcnxNE7BBsWMK60qsosykxP7V04SyXLmCnZ
QFxo4p+T77vaCzHBKsx/oxla6jVW300u6RUgVTBcVOiIo2HT8aiH1k5jk10wm/O8zZDI1LRMu4Lp
wT886jCAgvIw+U5dJepL/8LCK3GGRfvtsMT9XdPoqrFIPdp7nZFI/gx/vopeBtIivrkmfPtbQNC5
dZuSZ+QlfY3+ryklmCKCTJ294jOp5vKcEC1Ir9hOAUBZXNSCB+86AOToW2uKeeQXyoX6m8mG/zsY
YVYTgr4ontwRIrvEQZQvnDMx+bKaRTps7d4GzJdORHWcnWxNaLiC043xSjfe71D+p+LH4wv3Gouh
XWggqGpA0+sIn8dPYormKeAyCA+gziKpD8u/LYi7MwLvA8CG+XaRK5aSNxRAf10s37EzXX5KnT1T
Dd/ABOLDU4gUj24heQby0tfOg3E7Ed6d+5obBEOYtxSul1NWQirecn7bZIlSsDJOEkz6JU+e7bM8
T++J8SU3UenNIlXpj5ox1bPDviPN0dP6aW1x1/2uDEBJRNPU7dQxFKPKo6R6HUUbHcE2jXRwC9PG
HgDTgTeZC8G7DeTWWqyoYq43+iHNlUDaI6bTe8cKX8H5ucPK6zg30jmkVtglGG0s23QjLWoXmaXi
S3aE9NGRDWXvuj+dn+fk/YYFNFAur/sNAsQVKQz7J39dUBmgxGmIIhHjcXJ73kBwfn3OQoweQ/OH
iA8HukjQ+YA889Qax9I+5XI7DUurcJuzUnMd5OC1gOs634nnj6+5+5m7V8C9siEejjBnFYDGY/9E
/Xb748l+HyNOvWGH5aLOVH5fRf73LcgVuBiFCJ/4PaCCvMh953wlL14s7/YdXL5s94LxQ5UPTHL8
mReYNNiBmLrMaExb6Q5gWm70JFQexkfc5Uuq8tHopEH6sc4DjcXPxrp7JSI+5UoH9t8E09TwnBCo
/JwOUUD6lgZHjLEc8ZgZXzYaphOxxD/sxeUFMSEPYZyHR0d5NiWqfjzOSpN34xCG4p9GK3GiO8dA
rvo0Y2aEvxmhvjAnele8xFrdqAxdTI40Ci4CvFXWG3PGbzsC5F94G+N4lMgGCCnJQLoiPLMZ8MZw
a2kKAJoVhQWY1GfaqXvzixYb4YascCAFpAZgFRBrQCCSnvNJqDwe9n+fE7UREWFpPM4PuUu82JGg
09jhvfqA6Fp5XeSn9QG3/Ikgc9L0Lk2mFm08esWrFVxTpDANvNlPLRuMKUZFxJYEbU8VOqUj/Jxh
7J7n+R9jXbxnZ/3suHN5yuGYrBKRyMuXKZZm7BHN9fh8ZUgaNaDRAkHS5QXNyaCqYKjXZkiSlVyf
ovghbdfdkk7FS08EH/osrn8honl5NhEmOq2cemrOlVwr+4Yc1H6ftRmh8JvbStcSLqqjx1liBL55
A3XeidZZKvmymoHZEPDLWh1FqegawkWFg2WKk40EKdTtGfq4RxRkmz5NyEEt9DwPFzGR74AFCjTD
mRV83+2COjFfNZP1r/1Yf1sGO/NhUF+eZk3P6RIQK18V2xy1kTOYki8AlSYrxhVazjk2t+0XReV1
If0pOiUE9bxe0edYYHwZrH81MW3c/ICYZqr+zKJXVvKDT+n3aBPTY/t2cKWeq3dRRzIVeSc8+f85
NAJZm/O8wBiMQNoWYVqjfnD9cZoK7sLjat4W8DPbLzzn2UwX5tyT8VZ3eO8FXA3mDKNEL8xT6JkS
0q5zCeiFZ5HfK/IIutR91wVUp3Nf/0iqhWdUVxN3mrYqEIXY7/Sxvh+ofQDO49j0PTgyd/Loo1T7
MgIvofXNpufYxhDFVV2bJBzWEUkOpB0DoPQakuvcvbT3oAauToBO67PZO3ndp03YwnsX2LSvdvc4
Fl7qU5x9jVq94ruxrP9rFzCw8mlhIA+yyzFTUsEf9Hkt7TGyTLhvP372lAiendP7ffFz1GxBmkQr
JFpENiL7RSCYVlG3og8WF4M54AMGiA5iMviG+relVK5WZAon3FejO5E5YzKnuw70RV8hn4o6oGNa
UrB23iZbpNWkr2QEVL4D/GAOv+HSjC00TaFILgkIc05ZB/OAkQwSE4y1afuBdMwb2yvNUmCPu/0v
HcxqazouyWL7USGxuQquPPTXUUFj8SUjvbkMZebT1SgIL8vgLuStPm6O1YJLcRT8p2t1mFRk6VgF
23MeUQcdjdJFQ/DhH2N5rhVywqCzb2ArhbdSKPHLnu2we60P/qbvKPwQdHp5QqHR3Whd6Cvb+1RR
oQeKaPiH7GyujjBGLwtx64dexYL+QVWSnOQj/69qZRU5YfVDljWe8xOT/XDLqvV1elD19RDcFgZW
VtJx6NGX7MlMxSHV0VhsHZuInqe3coZKhL56Mcf8k4jH/2JYuWLvCsQFFq9XVG9RvtGs4st97QRB
24ToZG1SS3Cb9ys9nbJKmR8eYDkyvX0ZE2h7w5UznKXDmTAIs04vSaELQRe2YQ9iZNg18kJD7cYn
/3GGuBWgxa1OLydKJGA5HwZFFkGqN9DfnyHNdZiJVq5GvIMZFSwS/e2rAsQDzQSVEtUtqK27h0hB
Fe5KTP3N/CZxWrysbzBznag9UyML
`protect end_protected
