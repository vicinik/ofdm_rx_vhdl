-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
18W7fE5852lCNAyxyVbcPw/eLhLPKOrtLbehlw2e4mTzv/LGYgyrAwXrcjME3oqeqqvxOpEV+ogg
ELX42EVt3GnlsFG+AnFIN+o/ZFbwg6CCudPQ+7m7V+eOYmiUm0mKU5KJHBOXsajOS1sqwAsbOF7b
EdqSL+Dn7pgPUkhcIzyVae3GfBJdPQ+6hneTUzENjDfu9r2So0qz/0mv40ZJIYVvzonnH2ScXYua
VsJgTxwog6/3HIztUHsEpfIW/Nuke1k7tKP6IJEGpgGbffeP/UbRfSGEK00DCrVvBrh8M8G9NF/l
KbqIN9x3OiuUFJ2yAqqymNmKeosR+3gpVJqM4w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25136)
`protect data_block
ZFEYQ5k0VzpMx0QVKo+9tG0vWv23MF1oLPQipgcMyHCvHgb6arzpeNyWKZu8bGGlTzQfz+7fd0wR
oa084zVZInRHrtEJtIBksoQwwQbTZPieVwmlRlo35lYZl2fOX3HWjQnLJvfRbxW9NQCtNgGo3wzw
pD5xSoJYqo7nYeXrjTO80QYxKdoaYhk0FaOA2AVzdqyJOd3ICAQjkYcszqsurhSYwz815OEN0cI4
Rc9SvRBoUpIdvyuheQ3ryY1XUmG0y9pefzs8AWzse2jLAAeRLu3/ukBf98zKoFQ3LypMUkNKq0l7
iHh1M8DhaiO9uZP7uFY8KvdefqhcHqHBfBsLCFbsHcsvxO2lMxyCtHBG9UJcH+91VSAF8FJZMLaR
GmntGVfuL9tJ7S+NQAX63ZjJ1mA6WmX1mT2bKM6Ds2czPVYgic36c8xaMKY7BzUuHDTythbKyXMP
xKnRP5+T73IvTvXGpcqZOXr5nUaJF4ZVPI7zR0wHxnEboObvUqP8WLxbTdeGAjFvMHCy1GpUASIq
bG51qvU/CWSXKh2D84BGnq5bdDrbEbyqUH1ZYe/8z7Oef3ierEe5vkSHcinwxWx5/6ML8uSandJX
JwTTrRl1V2A86tEhcyMgM5BjHhCeA9EHSEplUSnAW5wgdJV85RxXY09into+wIjouOp8gXx9Q07o
TwQ9QTluGals4uUmqigJkFmuFxTVT7t0HEmafRVEcZgwoUSu2/jWfuKf/iRkdkEFR5aKrg1peqrU
orVlBl4jkx5HxaVY3IwCNizkHiL05GCpgbVvKhvacvQwdj1b3x4LB89cy48v1tq1WSoK39rPd6Vr
/VpaMAWjQnYpDeFFqBKpI6s1wurXCEC9R1hl9hIIZuYK4D/YXQL8hfcUT2rDvROpTkf1n0/jQuAQ
AbryG9YtcHodUVcZnCOS520ObbCz5EwNvYpMR6I0alaNA5C0JmRmndAp659+lIfgbKO5V4iUqmMA
7S+5g7Lb/RRgedu4BjQGrYwzR/nuohgOn7UhjbfMJqc/QSpI4xpyXpZPJhfBWX1ePXuv3Aeapf2F
KtZC1z+YT0X4O6eYGaozW3QLa9nNPaji4cONvUFEqM1zyMYEg68czmLTREUXjHok/XpKpF+/NzRZ
1/FBC0EfUpE4H3cwG5yO+LQ7YrJH7bfJrJ0vKTKC8BA38FFhxy0rtKZC6hsWTIkRUOOPHh9tqqAY
OjQhTkuiNELoDBG2qUfKbZNCEsR6dhkVWk8+3dIYrz9CYZHqzty3cjqlVezCyh7NAzuW3vwkRoHm
Lnc2Uvfdp3BwN/7vRHflrAX+XctdOm+V74wT/ve2FUjpYrQj3dgD6HSh63H+v/oEoyBITmaNlaUM
hjPDk3/GTS670c50fq7TYbMYXA/zD5lJTkEo7jt87E0Ayg8s/+/YOiX95pk+lnxGGkqPHjNLNjYj
pVlqpnJexRT9rTopaLX2Ff4Jx1zPjy4mWpGJjIlUIb4iFLTKXI+OqzePFcsXUTCw96P0IeHDrmyT
zKlAvkKh89Ocr3HdT50yyb2Mfc3BFLf6IaXOMsGqVcURq9uDhjlY3v0zR/IqEaio0EzwvLRST4to
Kfo3eF3Cmah0QMXBG4Dieq4OoLDZlHsITT75vJlUI7xizm6jy78s+o0niF69aJEb76TZiniyUaA9
lZKYdh/SD+Do/Ph2dgIVWc9mDjj23UMM8SdXNCjjALvEBjlDGTP+sCFu72U99A14t/ntcsjmkFy6
OaThu/WfpyvZ5bJ6M4/ljW/BbMrHatra0oDlWwQK45m26uYzO4+N6K3RekO30DNzNq97m/kkLsM2
cPoDj5fGISauTEHzCCxPKmCa8rI/N0PrSVOIoaQA0AG7/0Nke/JYl3y6muTZ5y7SjyVp6iiQ2dvm
yNhLz/Pp1+bCwDPpDQZbTCHfBT1CvAe6XGgYZWCDJhBQCsL3Jctt4uhdPIgvQmdJ/nCxOH8QfhkT
hmMoFUFWV+4+aUBZ9HdbWKPDMRUzhEy6typ74tzq0pIJU78lz9242dtYbrLcHEPBWYpTc+PmxZR3
4RkWKTr3Fm6aM2HCoq1LeIOI6FNQ1bHA01v/Qb7OHLrPhtwrYx06ifmAbj3+GCoNq+dFEiu5R7+6
ghHSH3QzFtZ8Bzx8qyYOYDSqZIEE5ergNQosNt6OSiVrO3eZmJpQAYusHWkOOwRPWYT49eqWawU9
oR2rWRMrvNJcvRerdIwvQE90OEdTvCFPeM5DE/K4JFEQtAkhXwiupOSqZts7kG4/fRV4sjJJjzwL
213FgX4zi1gi0sGmjeLUZsPRkActS1IXCVTeL0HRPfW7ZDEero7vZr0VW0WYjO6hwZrjGjpX0T32
KNnia6j5tu1wiFru0gX7LC37rfdWwYlRclDBNkQxdshK1eHJcnrKJEN3/2JBhHp6LWcR7JYIV3kJ
uqMe1lsryxl2liXm0Klx42ODOUWIzY6G7/HEAydgvnqVPXME/54mQiUrdfPDc+xIMmycypVX8hAB
CsXO7XBwDieVZgNgab5xUUSD9C+ANh5Vn7NgH7dZ8U9u3deJG+CImRns8+/xYaU6ZJoa69tUnb38
txw+AAGzb7caCi5fT/cHJdWPnroe2E+UOhV5ZUrl2Dskoc4fsPkAFBCN9TBHsAFu1g0e+7ZTtZKC
uCPibUyJqT8UASpFSIDN58ofg6uodbFg7rHZyqN3gm31vzHVpTKn09UAWK1MlrW63iox9yrnyvI3
sL+mVaqOJr99SQszeU7WGCpAahEfwFHooOQVYTZAwHp2GRB7DoBt6gfOuwco5qG21IV8hFRn4yYS
T/G4qcTqyGiOXsYOFyMU5/hPc90mTbCdS2MIhxjLl+xqDBsGY+IjlBzQcRRzln+f7UEaAObSFzNb
uIvwDIiOFEzNZor58+d0aZpwg1qTfUw5C24UFDIufmzEVC2sEJpJoL853bkqYYQQmsmPCeG4LvFh
IPRkWqeC6zx0+QeolKrWUHYDbewjVgmQRI/sOmC5ym+BF2/x6+1TFf/obeD4wEaEbPwA8BPNN4VE
ZfL5pn0/xo4WF2K5YeS1vCpZLB4VlAABbLHkZ/QG96yoyjs4i3wcNv2Y8RUplfI+ASScgSiDxXDV
VOJJZASLKWFJoNHqq3erioQyW2gliyx+/knHjCMKiNa9056026rHSpRET0YVuI0r/67L+26c4glQ
1LhIrN2LW9KbZ32PfTYASNXq4l+aYoo1rjfgthoSn8Tr+azErYidED29sFRM/bx/zVlLqOdgD2mG
t720Bi8Ks2t9syxn+F9WuD9v1GtMM736H0ifSaK5ZzDBKRajy3fGTldkUVMrXtoMfz8WCoGXkqK6
3VgxnmebhIkZw0Iv3i1y5M33RwXQaBIWYMCwoAn2epfurkJ3PYLkVn5oxxVymtmNulu48XPoiFLF
ciMieejwKgVKQa4O6e8+uqdRWQGsr+C5bJIgclij/VYJwX8Ur3SyqecZxtAqOLT3aQ6HT1PIhuQf
0juLVb/yhqgNE3CbSkVZfluC7GGnc5aeP2k37Fsqr4fet5bnfGk8rSkjLSuHSxP/3yeyUH7iaCJz
aJxTopuxWWxPRdK+4r5XbhvOOF/slBxRk1Rnu2IZnZQjKc78WLs8b9Y6QtEsuI8jnzGO/J/UZ0L1
5ZvPBQ8QdDPVpDw70inWitvgiLDy0IWK1dG6F41u9NY3SWZeu8TWaf4CQ4nZjmVDeQOMOpxo3+9+
3ovZdmInCNvired0kKbMtL8WyFKZGEFIVykNfj/aeueevx2zt0pFC6HvwaE37mOr7rvOUitvn9Q9
BFQBpyDSt6EbL2ebKA9l31IpbNhGGBb0Pu7NztrPe5ZzVkOrHDQBnU5EpaoioF272wqhl7W01HtS
Uc5HQ9hiRY36C8GT403BxdfUyepaY8XKB62QSkWXDjCVJJ8YWWpf749GeElf1TVPBPgoWc4OXTWp
qE6qWDww7vv5PfhdcOpdiM6G9a2doBSAW/x4SWES66QgXIL+aMFFCSkxStnpfoxyTmLZ/jXzc2jH
toycr2Syd7e4+aJMA9GTgfkfMx0JHkLFgCmPD7DmPCDtZ1Q/5QGwyVlYP5an2rYPZFzExsTX35uJ
wM4ahQd08QccZqdS83VFtvkEWoe7Oef/IX4q0mEP3x7jMEFYR088q9eM1Vl4NqQZ02/bPmH7ELVo
03+wqCpw0h6onqqpr+5fxrCPa4GksOd2Yf9H7aMRg8sZN2ENoCrcqltcex971q7Q6She6n8R7VDZ
OjHEA3kt6LQXuLQ/QcCrejwMNk09uQjOZVMuYs7swUKQN271ifA0gQSKhjgUUPp1hIQY9q6iMWTf
wJ01XA0aALbcoCO/RJlqZonXgOd1wsEL9iJlN6WhmXh6tO4A0SbeH0dUaGdyHGkJSEuM9V84y9+i
Aj+xFwaAR8laPyXuq5wxYGYz1YNlIO5xwEpeuqecBs7fp/05Dx710/A/wsYxBqHTKR3GywffuF6K
FJ+QMvEMupby6SefKrM2ioI/K3BW25kkDBQ6U5OpoX4EuqkEHEA5ToZtXb3AnSnM15DTUCVZIBBw
MBMrf+MOzxPMTMfHHeQ9FnUOdiKqMn36z5ikOxIBq2UfwYIqV35YfKBqabPqQg2/WPTniF5WhjuE
r3kbHkifsfoRxn8HOGJOfPVE0YgdaF+Ms1SVRP2Rz8p3eD92WgST8oGHc8OLKW9JtWNlNgyY1avZ
XgukMxS40LvlxAsRbMLnQN0MDgfGdXXuNTcz2aTyrotB2XN1gqVnmLk01k0re7SIS2I5+xb0pQ8W
aIOT0cEPMI4N2rv2Qu3WUzks2PCQqfW8DqwjlX619/aEMZ4k6jSgwXddOLNaBkDafKr1MPEBI+W6
mj9c3o2UsgpZX/Lpa178CU9b6EUHrT/OXMKCOlMAX7UGBfs9b1BzRDiRvWbDoaR9Noawzt3ddVLw
E95Sc1BB58dbmcmYtpJLuTXTXxSAD8CDZULRRHul5Qf44A8CicUteSMYhPClglG4UQbdZpO9g5PR
5DUPI7koYig1NDVOoN/r/Z3bwxKeiSCN4L2xbkTMrAKKiB+1oW3pMk+mJfL48GyC0b5JTNBHaeEw
NVLZLdDI8KXi6J7TqoK0XqAyiESxaZK4+lbKoNabssObNqk9z0wa3E50B1bsT3nlLOnyFgWOFAiz
3gyG+SgBt5M5TBsJAGl4l+9pvyJNV27Yz8hZh9K64zljzV7Z8XBouAKOM1PKt6MEXrIgsmxUSCiO
cVbsivGCh9Zv74xNrSm0gP7wDLsXuQVE+9g3cnL5D8nRfew9+B3D9/Agoebma7Kj78z8qtSObXIi
GkoiVWb9/ZQcZChX0OzY6VihW8iTz6oXcY4+pIvk4E6/l+uCFGVWVWg47Fm1v8urMSNcbpYIiUfB
zv5LSIRFTPkHtWZSr4bLP3tp7qOO8zxp/G/oYL80LJb3GOIph6S+JFJ1FhbaD/vMmg2Rrxapdx8U
h+gbLFk1GSf3nSks4k9+ksigaWIA9C25B+9N0rn1W+dAUiE0BjRsqozKlKMw8Xj7naoN43+qCY3p
u+aKWlMDUyv1NRDP3c3oF84lbeo4h2g0AgmIQWWNH9EvXLeNJl/hoIgWIToktBNF208mBIqoUhUE
pKqb/k2l2Zshho3uBp2KoQKlQM0gh633G67vOqL9JQdlMicraIBR2Q/BQ0sKpitgWtJXL+eqraRU
tZ4Ze/j3bboFh8DwcSh3FjDK5LepB42bQN2+ZoJGTURsPvzPOAAo51w5ZTRG2TGqo4r5uLEcK6MB
qK/e0FrzS0wpAvRuQrncWFYi91fslEd5YOeCUHwAgsriCQnKAun/j5Zv7zMjtfN44npHYbBvJ3ze
7fYWvH+DLuunoQbA5Bfz/vTgth6Dr+99HjpVTnjC+n4f/OhSDqB+9ISnddMTcxEsC3vWCdQL0jBM
O4537AYusOAMNgIarwYdbVOS65/Wh4LbWq8PuvLK48/Z4jJYYndSt1qz8dsfrU82zEENzN53quCx
bJQnVhxEYqk5+YOBslm+h7+c5+MctUIm8oI9W5xg9zfeqUHmL8+XAgqLiLc7kIxcNxQQtQW9dipF
e4iJk8WxpYwOEJS2kcU/S05YN09vFxaEDvEEHOVmneFpjr+CJECA57cx1+JuE/HfoDjTerSm4g7L
aQPxBN0Kj5tue31IZRuAw5oEQOmKRxgWDXAZAy02NHUj47m+9OYhMfmZ7eh6jIeI25HoqrWlxTuD
DABlUQzH74vSj+JGaXHehvGsU+WHoH0WI4o7WckeE4v3p1MuU0ITUZKr/pJKh50nV2DETnyzrtZS
O39ccXOTw6uAtili6MHdmm68cKkcgFa9NlA6ljRdDKDa8p33+bi2Q8ZQLuMZx6jHiXQkIqHU6EzW
Bpe8MjFPV5PUKNxZbYw9v0iLwzzKVstKBQQvyOjmSVLPnjyKqk7g4JYa6PFUbunWo3hFwfZsUU0p
UH8M/nLeG1DYWJc5mbwFn53TMh6w7dmp4CH3r3SU4oKRZvUGOVli8/km++0KuzdDUaGZwmzj5Doh
cYCCfOLwBSOSZ/DDM075bBp9q15iaEKQ/SeaBegXUXAzWnlh5tU2LgsUoD1u5SCBxRESLfnvQFZR
xMyasRCpaZIG6LwwHD7xSHk34Ury7uPU393cCqB3vVIUWtHWJd/xNhANmdH3BKfnzVs1evoRnuUl
VBpDzUV5vhOCCLrMbZfx9QJpflQH7LVUlPXxjIZjpR8hyDpJ/bM35K5SO6MDl4EYFYcDtHI8LkhS
Wr3/l7xycacGuMA+gGxswaqJyClQY/n37BeDlnfRRSJRBl2WY6+LedmtWQdPhX1lNdt6aaZ/KKGw
shfKPwKVLDsuOmSR++aIY56ayb2Bo0zH/9EGJejXE/j5Gkvkl06aZy99LNu5c9Nc0OvM6pkkKT+I
uEC6fEEt5sjHhxSS5VOhnoNF3SAB8IAFjPVsrklNhUP2W7zhZD+IdbH8QPP5A0oj4CFOSbwR4dEY
JZp3MxG34yYU40PHLIwFjRRA/wVCpakVerQlnKs1yW+lQzMXaA589C4leQ8Nwm9OU3tqChHt3ic8
3v8Hm/gLMi1Yz4z/v+ojeGZT40kk61X3iWsNRKhIUunZbuf/XQFehgVZmYaTDJoiONDwymfccJgS
fFKK4Xr+UKRyQvxicB9n4rdH/H4rH3qr7UTPj3nwpb53ldi5FIE7YpsJ1TC0z8vJwrOO9TRucojx
4GMQzArZvHu0PwGC+9dyiAW/+sTs2lTlIUcwNsD4iIGY/svi9MRtngNA5HnsFoZxl+XIcQtCowF0
JMvuGM41NLX5TtuoqBCC3Rq5BEicvfQrs0bs66ilWl+y34ItEaTBgaHwgY2hJFulBE6oGnx4HwB1
+APBJAZBpUUxt/KU7eMSQL6THsrOvyp2jBz4TnKNO7J6/e9Iw+DfnBTYJxe8m2S0uA8pgzcqlHGx
kw79bprxVIKyoPicpK3LtiHMpoF8JQ9cx8tmAmgfWOGPU7oOd2NptonGhKRxlPDmxUBlzr60diUh
vcwUEnFfLqEtFmR0s/GWFGgMfBn/yB25uu4yJHO5n8YhwWHkq19B8ozsK8SoM5elsZgsZX955LMK
gVur5inI/P+sgwfAw27r9m57suXUjfrY8d/s0VwYhL3y2v2GSMZGs4ZGhTnpIJmWq4ZPLUfO48sU
X360huBgisCYl/nTCsblexqQ5wGXpJYSZaSSDPLDyummtuYRA8+tPieefTRTkWvZnt/iMVQCVMIZ
eIzAv0coZtiWCW+oHdjcmOgsWw3kuDOG4/WHc6TKBI7P8YphRDnTwBM5lIxjxXwsgDgA7h473Bfg
7HEzrrbQMMYK58ilGrwONSX7ipLltQlsrH4Od2CCVxKb0IZPKPgv7G4dSizHy81p5gn/4vXyBSkM
tbF4bTzvaH04pue2cuVl1T37apmeXDKzcLWLMO8WzEdmD2eGpRrx1mdCA/ws2hhITU3SMpmz5vzu
g7v6oSkfTqlaBb9sRw3JWrIrzdl3cub1qQPQQYY3n64mcMDMEpTqORBEX3J8j9Jqidyqh8gZQNYf
jWDYQOByyamoomEm90Kn7qVLMiwowPqjFUcX8kj7o2vO9RsNKdSsjmvzWin9XjtIqqq6swfGkJzG
GxMhYKdJj1csh2D0B6f2yTI4J+qNG8pz4DUYhPemy782u/KsV6SkgHoBcuIq1NWS+2zEhK1Xlu3s
AL13wLzxxoXPzSAVT8EHwhsaf5pdWYEdTTxL/0uHDOgIyAsYJ3j5PkeT27yc9PgAVWiXFvEiM+gb
tK5O/m3yG/3Mc2ntHvfadhgbmHXI5Bo3kRLHqvaJVsAapOEukiDmxmsXvfy4rekC8WI/YsCp95s/
kpgjtDhzEuujbF9J04pNBHtxGwAeV0Xgv+XfVCSJYKmoXsIy78PrSBjduX4zLBTYPZ6GmHBX6QG/
LAIibBuhTKOjliaEFaIr/dSmpIwW5LF3srgYGLm8V0j/ODbvb81QubCaBX910hJRrfYlLilUz6qe
K395MApqs7Ntzls8GOY1449G0fFEbFwu5BTALpU3fo44sIg7VSB2BvDoeDv26e8ndKiiZox4wG+H
Uo3Ln0gRoNBTjxudkBvJJx3mr7oo5SopMez7cpemGbHWCQtoFh5y4VpC+jU5E3tpGFMw4MG0JvxU
HMd5M4sE5KPjDCMJhcX/fRafUGScOHWL7gdmlOEI5xKq/HfaNHJeRvRfS5d0NKbp2MCGL+1WxpYG
NRA6S0AnQFIuBJ9Yw4p8UE7aFepbgnwUcIk9Yv15LD2d1xWI0nV67HibhPFLZyQML6AMj8rl2/Ho
kul6k1UG6rbFmnvim4H6E/vt7Vvrpvl3wkGI9WxcID+p4aB9DhjTxyes+e/ajW4xsR0CCdHxUToX
lb/bPvevG3ZCMd2fhXgN1EUZwz0p5P4sJ/wDDCN80Pvt28/hOxGoPyNIHO/6+DiHJvuxYLKvqcBH
1GISpWoQ7nirjJ51MeI13lSWBo+ZP4xv1XZRy6CLbcBad821XFRFWbYQgG4NX8vAlTg5u3PoslTI
FIB3cgoT0NJUiLoNLsxvJ/fVyRPY5/sv2gEx77otQr9bTJYncDWtxzq80SY/xnivBaluGEdaueeO
AzpWM8Bmm0D5yPeeZ6R4v4hxor+0VUfrCa0jDW1edfVCHR+SEco/sUKE95nuQHwW2+wYEvaKJ4Nd
+jZoabDV8gfPlaafLSWec2Fo77fHxwjKZBCqteQFhn/J8ZMrbqyjACBho3RE9BkZIHPRjVKoXIJE
gD0qR5yRzNIZDDCdNo+PVoHGeoXSv9EV6LXb/4DbtAhqLKPuxDNlYvOyTVNc4V25agXcjNjvJuIE
0DDYtcUSkUWuiNDQlWgRI/w7mP7NLJ9+DVIVZvgAFAzr8XfQpy7FX1e/N7IRz+RKUEWoHqg+djsq
uV3NtKzycv6jYqF9iKId7B8nyWoO3yW2L04I4AOLhZ6DNmjIdnx2NLIxPyVLvzN8SZpHNvdFYJoq
6i0PR0VoR0mbUZjpCunPW5NKArlcPiX8qef00h0co4+wFWSWzLPBo/QiMfc6L/Fbwc1baP3cxZEQ
u0InXBtc7JHrvcjA19iFSVJwdriR0IZusU9eJ0P7niiPZJ63UkAS7kLvDKqdUZnwSh5CDMMEwDQ4
v6xzuNUZ+Pl7XLuxirExktbzAm09LfClnnq7bvU67GBzWenLmeDhKC6CuX7OgXVW3riZKamxUmku
Lp88/L5av+CrR7D/9RxPnq6mRG1yzJFNsmVj6OtOkTNZUksZs0xTfMwJlngduwCcOWzuA5+YJFiB
th0PE41mLr3K2tcWy4UQEOeFN6+nSAWnuEITghZi2046Qi8jlwnWNL/yiuekvf2cgeIw+e06Prqd
pVDPTVCVVj2RJ8i2nq9gfx4vwChzX2qCKoxlBA+Zm9/r76g6fmXZWmQ/aKnzIRTdPOE9L7G0FDzm
25fBjvcazjlE5qbjdhGheZ5ZS/4ESZrMJqujd5nmnN15yyJ9AxxS1nCJXAVdqXHn0SJC4E/vJfBy
HsNvnJJEMkmv/ySXt69IfVwMlqOyogpUGbwCsYKWECyoeDVylsryz0VR2NKJlXK4CSYQAxC0Ksri
h7qAS8AJgKoIoEldU9Ju+C8JO0su09dWoncZFSxvlX0GTGhNtUnwig29ZCPL444lnkhhnT/jkA0M
7SJLeLIeA96Wn6ni5z45JEV8nZf97uTGh0WGCnF8N5MinTX3A+SCtxQpwDxKEqYCDcZ6CkNKtK+a
5D30Uy16yvkqx8UdU9eWx+DFFpbpdfwosfVBFR8cRXr/gRdJgdxQAdQ9pkA3lMSWEpMlSLNf6/+R
tJRBXew0+55mZJDQaCK+wTWFXKDo4TR3wj+H2HiM5nS+NbDwjYzEwJqQOzwW9B4PwPBZzJZc0jno
Sjvkh7nVBS0TgeLrbPyyRCL510kggh+tKm5PIRbrX3xh/qdebYBx/I16stl+Z/1b4G3zhfzmayVu
PLJE4ta/BocCm/yWz0DgUaVaRbTb8piA3vmg0R1lxE9jJjGy1EyGrgc9aPFh3t/BFOTscJrHMIhj
EX88F4MfTDuLNnLhcL+AIhOmz2xCaC46CL7oLalWW33WNXo6ylYRE0kCCq1P17LxNFVSVvaOA4k/
ZnQMYS7o9TwfHpp5NyOVhsXukbKYMsgkYuYglEuUacXgg2+45tXNx+BJJOFZxklHDZJA1DVrmL0m
ewvcSpkQlSK+vVl7XimaO5pc7uCXpvKbMJxmHnAchRvDqUUlf2eOiZ00bZhBwNcAx98sbVPQq3oG
Yc8ypToQ2TQeVPKrcD7eX1AbriBxpf3mZltFIdh0PDKEMCn8GkPfxPEUGiNG91lOsuq+JGRMSeI0
qqz6kcFC1ejz2bv3dqvfvPj0wKeCSrmzsmb5//cj8Ng3Vbyv3/ED97fcRc7r8x7cWBp5lyGt4tJa
E6QBpxhPmBRNUrk9FMfpCPVZVqSEZnBbjOWHO2pRWVGFn4v83PSczLYIw4yNlt8LgvYxmimITTO6
lG/4jQFwXAkdHXcrtJu5EBMe9s/yaFtrtDbnQ6f97w1Wuw6OjpZYdauuC9VY6QmHwFIrM6/6fImX
FsMgt0NZdrutjlc9VqtcdufkEGScbDKXSWi4jps77JShw5mZ0wGscV/rrIMWOI8VbQ1Vci7ZG7PU
jAooKPN4ejOd9IPN0uBzWp7kMycSusYfhAyJCmxBqN/7rqp+U0LUP4iVqr/aeHWlnRsCwcyxs+O6
BEzFt9c531F4qWuvcPAdScBnkMcYV6/CEdzGQsbW0pGBG/9zPWK8ofi5ony7erKd4bMXha4irDO7
Z9c9TsBlc+kFIAr36qCBi+pXE3RX3gCtgUUV0l5IOWVg/venmkeg5LAuhioBIi2smhIko4YDkoyO
R/ebIwMVJ+/D/l3EaUSXMxcX7Ah789NEGewlwoOAtx7jSSr5BwJh3Y6cO0cacYGRNjlaGwSUdqs3
3EPykFLOLGacsMMOzhFsOWh9UjiZuBTk0uVLUcGBUz/j5GeKOdjsyQHR2eOrYXpe3fZpn65sHGPA
fXgGLrJBF8MghZyka9NkUi8ApI233hrWQJFrA7rUiC85Dti585wCX1HAI5ePDaySMbME3Vpx6qrF
kqP8UC0NuXoNNZngs+M2WuTOxfWJVL3DRGy5RynzN/oTGRUdU2SQRDfk2mPcYCwlMhxvfUDDvACR
Bn5GYBW7pRjH6mrh4CNeHN7zZ2FiGOOYY4Rlu5SwKHT979GS7uk1SCxtcUD1F8wyf/a/q4bSuxFP
nX2PggDnKbCwUht+goxL/KmBsUuGaAcA4MyY/axZXeLO4BP53xp30LKwyrQQcvks7A3/VGsvtppL
7aRefy9qrM5L2HhFO+0idbjoKVNKdhVdy4Sf7iHsrHI5YcOc/OmLkvbMFhpNnzbtkfi31iRPfl4w
hZ+x8vx0nXD+gqLGfthx3N/0yJvxM9273KsjLCAJBfBMLmTD/rz8aOLJOJctsmkSWv37lIuf3QTj
La+MhLiuDKwLOX/8jZZ5vqdOGPj0bFxeEtb4rgIyXUm4pTePhdf6K1T25WMYSQUiAJ1NgCxtlx0R
PW7iyD9XCrXFxI4ilIin6efT4TJ6Of/tJWfzdRbntDiwZ4RsAwFpwu1Qirkm/1s9vahh8ArBPBTK
lUjKYKwEZE9mVa1i+vQAHfEakZmj7cN98VvJEEyTJ4oGL9PAvVcL/33f9tF6nHw50PPyt0nWViYp
S6EqnBPq9pqJvDkR0v172VviclJYrpzmhsW4G4tupJyHKIiIjB5s7X3OZwC3nxYnMLSF+wVEJlCP
A7rQDKQmSSy44NUKJOIVEIt8Lp/Hrlt8A3mPaKvuQU5lg1k/a2LE+5QPxcbZXbW7N09dFj/p7KmM
LlVGNlvYa+Cd7WvY8sMZ1N4dGBkB7MsaOKC6HienBYMNfwR2HFklVXhU3xSY46QyT2nZNdA0UpnA
aVJXG7Q2TWatR4mRk69uWEPGNmDycc+7oRu70D90vxKiIrULYuJocBaNUst1UsgdJAFAqDYBDj6W
kx6oUME8AWdnj+H57AZNCrqioUCNR90D5QfjPdU9MhbkK5HEgCUCaUlMrm4XdM9iHmcO0tNOma1a
mWzBJBdbcW4RNtMTSHzMAty9LGTpkBwLLz1b7TSOavofqOVY89VYnoJCTHnvZm1Q3/hTomhxlX86
O6HQs0yK9Qc89hTy8x5xcxjZ+xNFj/ugLNioNL5cH8Wv07EWgo6AN1ubAzT50+JC3s+lLZmwqwvV
AO+pR8e6zd5gCZcHa5G10OKKA2PiXZigUGtYgA5N0QWdzJkmqQR7tO0uDRNy9bngak6NFQqLvenV
1sHEgpnu0xqvyi7m2y1TBV/Qnz3VJbISUn7pXG9HPs7+AGW7ZWDcuatDHQwoS1rpqD6AlNJMwtYh
mwkUnxZl/bZ3nRTX6FcPbKBaJ0QeBoFDyCfLGD48/xQUiK9W/qT7IK0ahT5xC+J+f6F1Z/IOx7xB
nxlGCLqCFpXwamVc6+lSUyat3i9VGe7zBQMUSjzep66b8T+wPJFEEzKH9IxljDl9TO1UA5vpCF+w
4oExkgFDFyIloyp8YEjtaJe0QZRYBXasTePUpifAUwmSIkL9E0HG5E7bh2uPQgbkkvd0Qpkm9IOj
t3l1O+LU3BRbZ5P4i9M+Qvz23zBVFBKKlMC1qdwkpGpyixQVZDBT8dM6mEZlzrZ919ajPkCwpKld
On6VnyN1TLZHB0dPkVJa1Z4kCGJnB/dhThF+ZjoOx3YidZw9+yjKySJ5sHJd7kTeJMA4ZKreined
CxqNHoHfrtd0iP7DjREo8QKPkPuEbEqeZwWJROW+js/N0bbs4IfDFQXc1ZpEe1iow/wx05vPS8VS
+34S3Dg6RwhUAn3x/2KMYagjzxRe3ZTMpq+VmfQnZGPC9lZ+mG1bp0nzKrqY9dgz4xd+euMEqIKx
u1YrV9vPcizoGwdp35fj/p/zrfaQqSHJeUzReMNQIgqmT8uqjJcH8n73Xm6lxu4wxwTLxgvSaXxU
QXU/2qlvHSOCgYQ1JmbVBBP33jCDCzSWCMuXIXWbLem7hqlDYIHjvumD4Qjlvwr0MQ1PVaoSLeA+
mzxMOVk/TGpmZvC8OgFvCaxKGvt5TVld6Oeg/6UA7u1K5BN2Nxd0RIZbf0zhyTKdkuyniLMfjdH1
7O85km9C2qFQcqiFXp5a8cYNEgNJEVrPo9t5FzzkesQp7kKeyr4FD0VQAeZzmhMJ+iPkqMH7mZLz
szHEJ+eysSFCGMwAPY9i8IU2tjDnhVnDk4bAz64fZVBB6LN9ixzKbiH91ON3DYJVrQWIiJ8TXWir
XFmzCZrcAY55ZTN+Tzw1BzmDiaARBTsARY9Cn9qvA4IoHJm4foIPvadGnMSel1XCqANoC9BGVmOT
NH/l12PW2glus0rE/T3mGCCiYc3cL8tOs0B9y1xNqgwbPCCzBc+Te2BaXMrrIMgpFuG52HeMxeJz
SvYu8Myx2mqJdo4zDtIpRC/gMKm51GO7o5N3NlZzkaPPn0RHJEbKfSLHrmI13m6X7s2vd+Ia683v
RVr2ULmu5R6NTCL9HNhHtCp/rA8AdQ+KjF0cheCmc2PSmsv65IhNDd/OyOedMvkYomExyyFD1poM
gHn42gx3kVOOkf1q0/2bynUnEoyIywZKDSueoaBmQjb/Tga5wefTwDahlo+8Dmf+Z1sqYh9LaP+P
j2p2A2N7K4mXNFgMEY3m/46R4XRwCGErNAUbMzvBkBvOOfcIn8jkxMv8MS6KGAt+s7eoAGdJUnC2
w2MapYPL5YzdQs0XLKv8jFSRQoci+Hx+cJ6fGz9X7qVzTkLS+Tx2KNpqYzskf6h3hS7hVAjBOkGa
dOfW6CcQoKBwP8xilF3YpyEWvcXw4Z8FVjiUC485sbZE0hVUooT/K90KLR7n48P33ZMCCAFsC6Di
RWdrUVZY6EbpUmzc4erBjMDS1MUybCP9ZlbQuOAjCfV01iWLjU4eg4JBLLyQpnteoxmBqjwFT3nC
ALDr7urPUUJtgEZ6K3VqdRGknBrXxhh/nS9X/W//lOBHrL6T35vwOiI5ZxiUhFTfzgUBI/23V7K1
K5L5gAS+bOfN20mniXVYxfB2QCrqoiqL/r3z9eP7irN2eDHfZJqE56phipnT7ZRQovsFb6ZCMT9a
aHnBvHCI2m75BR0yNMzIwDi5Vol+5aTdY3NTtSvT/3fgDbAyLTX/LDBgznqGs5Vy8s+MdZfVI6wy
Lni8yMMTKNBN/216kGz/VHlErPafHR5ZIQvGPVpAbmh2iVCK8p65iHUUQm+emdAe+zks/MCJS8uL
Muat2hTOX+C5aLurFpMXG/fOE3Nc/A0v0ioTJrhscFbHfYOyC6PL/z/2iISOLRIQJPF2aRdBylnA
roYrSznun32FrAQ8AecvAct5h/LwYq1RANJ4RFd4q2WOw5inzOGf11VDzd7QMGv1ZInupVy/VirL
jTvVyc2UmphJxeXCP+B3RJqodJXI9f1y+vsnjuJD6GWl+alyG2bWYdvA1ujYlmT36LkslF0rEuUh
XYjCsvRyYJiFtQn+IHBffFC7kuQjGUAe0dqgbYgpB/shTPaUix81n5eLWSx214kFDTvezHIBcBRP
AVDGbfKTp315JpfTdlGpcb/If/Nosacg0wfSt5OkCUQQUv78ZU0qWqCY2JfFup1wwZM+VpW/E8ee
HEn+i00Nuu5jQfHZLL6Sd0j1JHdEv5JdMeuVnotLgC/APXavJJGcWLFpo2zaXh4KWSWjOlWfUTIk
9KSnB2eh3vRzsAe7UauUBW0mic8n7vIi/Mo0xuTwPkXAYtYlrM/gBgslH7/f5SuQlcLJqx1NKhUW
e0saAmMqhW83huY2veergGibmdFqVNOgwHfeBK6W1/9e+MvEB9LMJmxylGJ4KwZgsvqxquIAhsix
R5JfBxA27qUhL9OyjeOinbd782V0VI+oRrSlKdrN5aKh4ZH6nxiAuT5H+Ri98ZUBPZkmgLyJHKRq
WOdqlTytVmjWG4p8cKIlO7r6xowtGBbN7JVMUiMFLD50wwr2KC/luysQ/HAPixnh8cBuEBjjzFrX
WrSTBc2W8gP2jHl2GQNY7M43XDx2jEQkObGhZacwUAs08oCbJAgUO1J1OLYzCqvx+01g1DDaGm3u
q0QALWMCEI/nZXxE/Rpq6VTxLZ94r9I8sPENHhs29I8t/o+IPfYYvRa+rMS2+p/Qaj8dprI1KSWi
oeiIsp2xw2Idpazfe1GTwtO73KxyddifLWN0Sh7xKRdNcaGzrl7EySU5lwZyGLC9OessJwa+868L
NOIMjGrZO+EUY6wrSRf0cmiWvLZTQwjQC4bozbKEYI6Ohk8I26xwJ5NutiqYelg55oFoch0Et8Sg
T+Tof3hZZvX7gMS+j0VzyhiBMmGfKQNoXsg+4AFmWkw1a0FPKCLSLXPOeaMKa4imA05ImavCngUm
hD5IMrOtw2kc5gvRZV2+P3ealzpoieYWC1AkXPclSVtaM1inYfvgYxaTzb3QDzSJbj/E6p6ePs/R
BwEZao72IEssyuBxeJHEiezJWhyImvXoPjxJtcbAopnESYw3Cs2dYfxISQxacZz1+FR4zUWWqWOD
Fosxt7x1AH8tp+NILJzqmxUejtxFRhhEYgnRFVQWU/SlIqVMFB9r2U+WeLRbxmdFYFvA44bPeBZE
N9g8SEpMAsspMaJRcOk8ols7yjr/QcHitscKjC1dcx75b2pcPskmKEFu2L16PNbz5mg3BsBcpaHY
ZWtCdJzCb0Iss+391LzbdEJ5yZ24NyDrAiWZsoEUqvCQLuTqHJ3cbHZPWJqKeAqagVIr2aL4UJbT
Iglky4q3VjZNgIoLvUKNpALszB/s4Rw7mN9n0OCjKBOfovU1knrPby0liA1iOiHHLiETgW8r3tSt
sO6JKxCUiXojYpt6EHJRTY0qgS7NLnpzp8j15Fq23Nigel58SRkiQDEVA5ml8Vtx2JYLVG0wwnI9
9LovpV5Ouj7WNTQJVh5rXry7tIg/89KowV0b1F6C4aCNA5gLgbq8RddVUAnPOZfhKtUYg1VNa9eb
XvtNqbN4jISfyPCVSzDyeNgLNC1CksfmbqIz1Fuo+CKKGtx0fufFKCnP4xcz7UNz+yyTmNFWbbm9
h4FRRhmIQ66uubUbnT7sTCSueP+wYonVsf+kiEZhPU6S/7DTZg5Evot4QE/x5h5APCh/G5XWYdlw
EW/uLDXIdWitDB8Q3oBbKNjwfxVoyrRCRLgSZMpjnMOV+TVq2Q7oWewgxL4lVGaaSXVWJ9xlX2WH
z2QY7n2hK+zQOGlBD/Cx9A+jo12xkfx+Ss5wzC4mdACKG+LQnZGNk3amloG2n/uarRUQ6e4yTCVH
mSTf3kvozrmtUsygzQS1BoD3uwbEkMG2AIoWoDBydS5WsVFTS0Z10ucLrO9nWXpQbrtASSNX2ZTb
Z874p3cpzzBNopdi54VuJVneQ09lhByM6aQukJnbrP97PCODdgxN/6rKGR4MRhKXVJJsFT7DOWLk
RgofpD4wnx9+gBoyOlG3UmQ8ixTLleIkkMBK+gB0sRXsJ0J90KPdxNRCyl8Q9IpIW9kTbyuo4yhz
9ZmOmUyQ3ZIXM45Dsvr07NZD4xI6CpYpJRU8QPvOFZRaAupbGtEXVYC74gBR6SfdW5X3ecjxby4v
kB4d3Bp1sAqTp7Yd6nEozWbcWGj1oCQZyA4GuYRUyFKDFtBDWW67oyqOGA4pgZ5QvKkH1skN4b39
wWzvhqeG9rlvr3KbZCzHgb8oKzGH43u/zAVXEE47brSvDfQj3o3dcBJtDsQE23Dl5rceCRQS9StR
i3AAmz9Nme+xDMmWNMaPNIA/pgCrYst1hgURENtS0R2eNZmz3HjH/jKy7992Xa4fpH6uz3HUvAgy
BMSZ8rNjhaaLK/LhGxxUtyClrAF+LEtbr4DlG38iNaN0os1AcApnCAO0aOuE0ojyXwVPEtdP+b+l
gCoBdF80xgwG/phNS6RZn45zzdvoUPIN93nfY1NRW9o494O3c3cNjjP8Q6FnW3bNWo6oQN6sYzSU
03tIUHvFduJOVnHc66H6yyIqQVHUMA4lnDMBZI2EVh/EAAdU2UF3fnuzsVg+cdshiyhjhjoN/3S0
e6UyoZ7f87eH3fp3mUbwlzJ7QpIR5TAEGhm8vCljWtWjCY4mFHrOs5+MwZV94UL6d2xLLKq2chtO
8iHRHSsFaZHnz+DwqdN1eRr1hbqqGXjYxxG4mn/dFB1sC3iYivFX5QRBlnjJUF7muHZJbqvOgATW
QtPIKaeJ4l2oNUt0rA7zf1MLswYGz59CrPP7WiQTHhv8J0rE4W71LLNUyr9lpkZ3FacVUpHueorH
VHX8iAu+Cr6Mn2GUtnwnhmvTY3xqMRIhL4Zy65xPFAo0kDmo16SuV+2zwyo2TVLElQ4sIuFVT9tB
mb6o0NfcA+Nxoww0YN8FG31ao9wpMCb7TXsFNFlM5xDakqjD/iJvOtdG22ApyBPD1xCTN+p99avq
llSw3kFM3ElJFzXJDdKxNZd7M5huMq01c8YQSY3BY24g6/XEd+kLiR/ihq5xm5yD7DeYF85q1d2M
jUC9XtgUgItSSvGwat5CdRC9xg03yIrr6Yy/Q+oG6dngEGYnfwOJPC6jdtHCVmY45jsj8mSbjvNB
GDyoN14b78ISRXe/sPhJj8aVaK8u3ZwcTjaqWhPVl9IA7NDC8xTohs3z7b3SqghRZGcp1kFna057
V9UJ+sVliftxXi9uEjLiUd6td61gHArTzD37GD46IARlPfLOD6iAngsDQoNL62j+7y2Vf9FBPsRV
wl2soWJH+JNnZllQvyU/V94EOvAIcOo7U/K9N5BzX080xlC6N1lWWm14mR/GLMrNKTu3rDr+7l5c
v+SiPWQJ+p9hmmnz7WwXpYiTYn38ggt0ulwmwxn3nAc9XnVoALrA2oUVXBZIQmsW+Ux0VxFLsn9j
Aa6l5YEoM1JGDp2oyTPYs88EF0R80vTrn9fmVShqdy6oDkLCAGUTXJ89UwHyqy+8qGYXEpemQKSi
yB8Ij9/+R8R+jdpIllshFbv85Aug9csqe8bh9SNt1ozuxT/WRwEX9EgOGTgjrMbzOr4ckZYvK8sw
dC5YJbfTyMSbpkUV4AkS9afJ+3u3WcxYfhdG91UDSrBC7qM3L8fKOvsQ7m6gbJqmBN2UrN543DC+
4SrsW6nfLOW+/V2jTiJDIqQ98UF09IEnjTLRapnhnFEwuN9dmIM8vevZMCBA9bclQ5IN7Uh/gD1Z
CcReNRX5CmcyxoYLiujO9ugQKVJJsB2pwQnt17s8ZfhhKqfRnZf172mV+v0Qnirbkob+fhhQcT8s
cJfPxvXnqtGgSXjZWs9yU06iSFBgvkFOAhFUP1R6GD1POSrJ0+h8MS4RijFBftNHUrFwjAIiJENt
qinIyQLtBMl3L/L+CC9chLFFZ0OEkKSOUrVpTmhvx6NI8TFl/E/bRcnglJV5zkJBwaFEhRo26Kcm
fL03np2weLFPKontpSH79Id5qWB2ZRZcR1FCV/9lQxjKywssGLH55oEt4ZXjf4tV6ZLsT91g5+v0
A76i3kJobFYNfUtrIVxqBmn8n1KNOqbBkujMYuDj97Opj6LGmmaQFLKr4G/nv+0x3wmRwGFpzBh+
ewor32oIPU9sUf5iuEvfjQ/mlokiki72fiupJ0/g8EDpu8+EgB4HkEyK0tomfLAZTnmqvPb+NW/i
Qw3GzTZZO/1fZFfejR3iqW0AWFoLWtzH7IwkWMyueIIUWOn8UZ9LIoknvuO1rZdW1eGdFPmB2F0W
+rA+Fxt0Y+M3e9X27r4yw5HwJ/H5bLNsd2riJNo8NHcYfyLFvg1KPb5+OrF0kSPVYOzfuZjob7CT
sAGItukR7rmH3sCmPo3IX2/HQwk40B2Yzh5rUjoKkDpaZ/dIzg9dz6uYCbZ+dQkRPe0cl8MCm86Z
YS0I/ZZkWtjcZTjDVGiVzAd8NipphR/3bvAaHZaABV1S3W0nN9Y3iq9gaPqKw1PtaYs/hXkQ3uiB
Gh2NQ2kTXdMfNhQxRkc9Kw1Bwxk2IgWt+v72lgWDiN2vD4VzRD9E2IgsWCIQzsjwxektkPQVec+I
oDjwL4AL1dOH2zOUkmTBW9VgI+32C+y6uCtjMvH+KejPo1zEh1Jx/Q6qZcyltV3Grj5SMmnrOnac
3niEy6vRU7b4M85e3IzBf7bIigIYE4OxIJ95pq7PGXiWvvGxBuatR6lh3QegYH5acwoehdeXkZed
lwDCbFud254ZF/A55Y4LMgME+6+TQjMEQRW1GbCzALMv8xCCa1MKSFnlMQs+Xo+f0WN4MS9pJtIB
R/iLJer9V8OfwFre7DRX7a5j9TTLRzjqzWqGy977AH3YEjCuygA+30AMlvfruLNp30+L3yM0cKpx
lTcV75e0xTS6cbcpWHlcVTlPLbjsdXM2Yt1Ad90jbBGygg3h+BYC6TNUt4a58Y8i2kbbCJZLlsC0
o1bUcdvKKtYpkFB8oqP1S8wbVjKDIRra55PuEyma8ksnI3d/9Em5okTxkWDjKP5Wenz+3jvtg1ve
PjfbhSVsVSUcVQ+pDAQKtMeQz3/3uQ6ti192BF9of832/Vxtct9iVozLx2kaZemiDBAuICak+9ky
rEAsGL3KRuijM8eHka2lCk6TscsulInrIitafnFHyaw0W9DnbELJo2dOg7yzFltnqYpX6Q6+2FMb
X7i6nH53iSz6VrwbnQkKljgTdVeedeVzeKXdTz2HaHuklQXeVtjPlN7DsfQNTDTKB1kmJ70ieGF3
n7CH4hCTPI3K4SZUKdgKm+HaItl5FwIoFUq8yjXuXsnG92jp2kp+oJfm8SO4t5QsCulyE6xCdPP1
vfdUYigd1wr1iGWZiTUN4pTfs4PVEYFi8Dd6aav8a1v3g5IPb7urhqbAf+tNhHmxFFp98tOVtunm
80MHBRSI6E6Ar/elr4gKD/QyqzeyXIME07aemW0Z4H5MII3mlzsOjY2yyaE/CSsiRGRNHPkT41Gp
R4II/hE6uCKQjfl0C0r1hIiMym1DGk/WzLlTg41I7eELIIKMgQvoO4LppVPgBSdM2rgYBPWaE4e4
eje2mNI2LLWt/v61I8G+iJaShFNH2aTSmIgqqY2Y7oAcpbPqnx2YQ0rKqTUrUNvdarD85zQ9mFPl
tKKc4z4JL3PZqoywgqPwoiTJET3I2BBArIBHpmoq0gIC28WKt98YVkSXQ7IudlKcyscGpIZgmcF2
Nlx34WTeADvwwuZDe9Bi1AXIsMhZm0N/9pHP7cua6FnzUX5bvBwvbY+TjsBrDl4nFelbZpkluGZz
Q5OX4f8frD7KCY9ZAZQFSQ+8LO6B6aZ+qdQpAcggayYX/zyaIEXRKAhLnTKHGd7Zlb4kSva54CXc
mpUJDqXIFBOjd7jLyT/FsHwgZr7DtNNPvNFTTlLuaW85WwmFLm0r1SoN3mjQ2bX2leOBw6GFPmYG
zZe7KTTfX/HlYWtiyGzk5Ix6DyzU7PkfXYVjJn9cKlWlmyoo5FWDqUwrJ6wRs60o2VlyRHmUstPu
bePwV0rR/MlpkH5+PtFX7pidkHxJ+szeo3Z9mai507foCJve74MKwhHFU5PnjP6ObLY6XLAMroHs
Ryx7KZ5Xh56ZWpqTta9vPgw0DyB8J2YzJm/5Dqx9ZzKCPOwWb11fPfP+f5UiEDD3jQcxh88eUyRO
vT7EdsRVLcIwfEyKxUIp5ApVQilKzeBG6coy2PQDO1M6eGdAOwO+tAaUEcYIAlp5NHBEwg+CHfoT
QprKW/aHdfdMVoTxKnHS0ZCLCfFFFJ88K0owTr7Z8VPmWLKyc+mjZtdBsThBRH0MaRuvVg3sLpaD
vSc1+VNBkPUH2svC6Kuub4sUREsOVt0VTsTZwy3Wpk/vQsF8EVbZsyywLa+S5iraz7LFWBDJtu3y
HJARF0Aely9Q/j5sRO457zyX5/3w+s7ARIfVDp5c+tf1NnDcCuHtxqTlmJLnSpoWb87Ziar2BBTm
YdeXcTwwI5VwhUeKfLgUqCLxdx2dTNBOR7QEecXW3SkodYqUMhcXhX4+CEgk1yt2wWqNZvum7XbY
bVM7DABI5oCChJePlWaDEVJIu7bg57um+MkH4dCjutY61sIOoj/ylRUXqI/aSzAxRO5koAhu2nYQ
qHczd4wu2bgHFPToCuK0R/9T9lpIrExpomtqy6fSiOTDYNmEdCXqWAFfdVjSyEnDZUNH9JTIRX8T
6ll9lysW2Z2lFfZYjUn0wHor0Hxqs6It3uS6z7LWffYU+45IJcT/YuUKpaswPZ5lg4JpNFn0v8BR
JwwjJJPny4xOHoXQQ+AyKkDtsA1ooDu52l/uzzJ7mfZDOOahtUmPF2I4DzIMBEjKeOEW40l30Nxk
cSt+Df9IzabL5aSAhcun2CC2WFrF/4MgXiBMM5k2tV0YIW+NAPL05Z6Rt6h1z/HAADsK/DCzg8rJ
pZIsrphlUQ6InPUVfox+1I/PzWfDpfg/WrNDBXwcUQOIPdfj1w2udti+Yf5K0iN8Ipx7nGC0H+ZH
4xzoylBvqMt6LNJCOBiA1b0l380b2cV/aX+siAwtZxceDnMtPopWng5Ttc3kwGC1CgIUvK8kNpbq
LAcpnDGohsgJnTO+8H4JyLepENZz+bnhdx79vEoIMKjBxkKyv9TJBsjZ7NATDCHw67HDWOfRpOD1
FT5VfOTJFw+8RGipa9DHDTHO645iBt64PcemdHH3wLeIZ/US5E2Pqvz+Sz3PWsn/rygD2zw3fYtR
JAZMpm65JqTWzck7Tn7AN/JACAXMGsp+PZEzrzRNh1B/UA8wBJOIyIKFkmrfCbPedoZu6b0RcrWz
U7oWgfLWTEQ7EycV+ePYsxRc5jw8a9D5gVI38NrZE+4JRwe9PcfpGiquj4gI0zY6AYaKLzTgL8a5
lnqodGVbXr2UNaZCAcbVba+4ksGWUs3u5tz9cO32mHkAmoZW5vj0nS8jgRW/1GPdtTBSTnTAMTnD
AtgnSsGUUEYvSoCC5hP9BrZ0YO7H77lfBkcgZz23xr/WQc31KVhJe3dvpvcB17z7I1MwOjacCRex
jTQ+uey0/BnbYvuVJuJ58j/Uy+ps8YDIVqoitnVPcqgGrjZk1XRVKUnpzMkVd9uxgSc5ZeLGYa3x
OUiybbibgAlklJIikEuyi5IYxSN3syDOz4d2h5+UtiR65pIIiGI7Fk/VOcqR1OPxbAjeVUwei1Ou
5DT3YO753uOzu9e1f7C9xax1g31K342NJkyhBcHjMIWJpCcqHGpDjBI6D9pMY6eKTBhLGAT27In7
88eUeeAcLnsvUb6ZTxMNDn96Oz2QIVL0eLTmLdMnvKiTlBEAOAjCub+REhRmB5bPrFbLcswa/y7V
UWH8geBUcq6/6b6NQuhrttsWR8ctjW2biQbWtu0ZctgZJB6TjcmahM7Ek6TEvqK91dG22kPVPqwc
dxNDFYB/gQSlBR+TV3TwzHMHjoBTxtANJ8lVVXEggOOnvmd+rNFxIoq54zNkE8t+M2brcbYJ3Pr6
ROyz/Ft9NqfZfzqnQryn17lRPcP1O+ylYNIgivYHzHdPv0bC2tF3yKrUWraTU7XzN1idgZbEfNKw
OkPyv1EFQDS6VTe+g7RNFP714Yr03Gm6P9FLMKnZ4TVZvhJCrxb2UvrfgaE+zJhVrJHh9YwmOhfj
1twaTunNB3MrjqvkSItOP2OBVnnmQ6XKUA/ncxvIQt7VZl71Lu/n2++9J0nVVhdHtNTQInb5pIYz
41mD9N7xh1oJQpwcWvn4NJI28BQsMSgE0MQbxCbh/NGRXRtqABERIdwB8JGmX2X20umC79sHdiPz
0NQVpC1H7021Y2ZCHv3xKr7a5dIUkqZc2Gpv0YC0AMRFnX6rYrzK7uKpkEbvrLkK+GCduBuVnM6L
JDqOy/yYnBiInBbFVQLfXx+E25yNZ/YlphYPCXOy9KQ8GzJvUt8FinecyufZY53qBUzqFS1WKsj3
oXD9oimHXxyZx0p1TrU660/3jZ0m9SF6af2GGoqzDZlmB9YIhjAUuc7kuF7c3yqVz9VfOrJJhRC3
3EcjdbdwMeDdXyTBRkQjBDunIP/wMOCrZMWlk1fq7bhCQoMkN6a/YTm2axtueDKAC9LH61TyeLxV
N3Obc9EAnp5ttqEPmdVwhX3CMH//OfUjRAp811yz1Mj9qeH6+gmCVO1YHXMm/E6qvn0Ny07v2PXU
v53p//S3O1JPcrAexWbNs5vMMf5BvEG56ytBw45ZJsTCFBW/iEgK1ayz16+xcxDbAOpeD4ZpToTD
5MY7iC86lalIXwoQuQmhnlle8STgH2saZHmeVypj3MRXz3+W79brY+6n6IV88aG4O+R9/JffBqxB
TUE6DqKiBZVqJwMqg2z8flwiUsVufc9ezbD5L5F+e55NP2Isf+NNbeS0LOavDrpaR4g9O9Un3JZR
XvwAeEnVJSHtlOtR+pzuYQGTieyRd1QbxyxRnnXjgeWp7KUNvYEyFDKnr6P7+oTqJXDkaf6IA7KB
Br0zF2ifiDdl7VpsaT0EOZNHUrkKPEn2UKL0QdVXt7zKyhZoZoNH4KMUiB8aB3i3hINwbnp0s1Iw
6gtwvGnNigat1hFKhenwpijXCmu8YEM4gIPkHPNECHF0ufKxeOzATP8YZYwl5VrtbgTxhqTizr4p
je3rxkYoPJvz+xW8+28zoRhdSK8+cHUjjMucnrojcXRK0F/pHYxWrjyXSqupu+Oj0JXDT+oRK0FG
itOUQktHNvQUDCFRc7jWpn0xlwK/FSFxZlu+43u/O3m36aNoegWY2fALceYeJcAWhnUvYYUOFLuu
uLYvFlrf7PPTaqxEvmjFu51s0PLjiEJy4Sn6vW+/eTj22htfnPdMk8PnLQjbbP+XQMPlb63ZpmIc
fRkBLC2p4XZD+ns2xi5YkysIRKiRegRzJ3KSq5UPGrtpKIXmc79puyth5rm8Zm+gFwps680JtxH2
OC9J9SYv48OYRjMp1WV+b0Gyic2HmaN2hpjiXjAXlrL50o2LOnZH0LEh/h2Uvaks8lbfZfzLQd0r
jLmx7eZZuUkQDMHX2FrJ4jymKSAOjqleYanpsHW+KulZfE+PUAeS2TLG6rqDe7mx8XpWpG6U15Ae
TvdlrUbLgOuXd8/hTXvK43ODOhSRF9Rxm9IXSrz7Tu4F/Tr9WQfeZ4YQu1OOxDAyhNA6ID5ap4DB
s+DMNyn4W2cXdSLaReeILXprtXuw2tnmEZ+c8QVk0kXpsWg9SNnCngLovhSQb62FmFttP6y0wozb
AGati7zUr1Squ1H7kVXrH4SHuivWoU1PwapqeSv5y0LBFx9UpKBEIitAOIkO8mnZEk3/zI5f8ZgU
EvXhHN82GefeA47IbYvIl+wLzt/XvGYqbAOLihHhhIJQGlUDmEz+99yeBGqnniEN8FW2RzJwQNk7
lsXShyYZuCJo82O8m8v/3vXY27FsGQvbMz6sZ9P/2vcR8iS5nOyq0x9Ncs4v8AtY+/nh59ZjN6Li
zI7sM9h7k0Dsy2pbO8sUkZu1Mz++BNx6IJo08BH0/S5W7ZwgML2bsbUcsv7gQK8Do6b6ousjmA9n
AQMCVZSBXnNOOOTFGyeOVWMP+UFyoOrurUUlcmj/JIhjO6dNHJiqK08eTv4oAx/hGvDh7thqdoqK
mzwi8LaWbbWFa53xOenRklfrqQQ3H/7T9FQfKkVzLDuBhJ4nZMqnSUhHNFlKGP07o2XoveUw0Eah
ex3aZgCzNmhbJwmTUaKLSHxM4qEuRyxQBOlSe0+XriHfXb8+97RVv1p3bJNGTPzyp3OdGk8c6VEf
JPhSBN6IbjlgRo1TacCiZh0YqqJ+gRLurz79Vu7Ex3CViRdi5ow6MDhWXGCdcA7qhyL7mlwtffKx
3zaHBelTgMEQooaUCGbJRVakweKgjtSSd/9skJba74P+SfRuE3p/FQ+bBnnNRt8xqJF38CE6KfPr
aKK90O8zAm4uXsoJ+/5zxkQN8goqXRxiAaDq8YoUQdS3xYFY+pZBH0P0ikbVJtvEri5RmdOQoIyh
ljC+6LKoejq2tG0BsmVbf9n9lK8VhZKRRyqVIlUSZnW3/6PHJMRpoGzQxcfgOBTEJumuawZqNpOH
GMdSti0ullnQ6L3eYupePSlgZfhhqVgTkn1pcGG8m/JIPIEnAj0gMjjh+fItPIQx0msAXXsqLeYp
WJ88p7XvH89mbU2THxB6g4BwbKCu18dC4kMjYDKU521YtPGx4MLMgWXnrL6e/QEYpeetO8j0/y5a
4SKT4zjQUHwWoa8ZJmVNoZEcE4gIgd5HIZOCBnAD6S/TpoyakBcfyJZ5Ro6i3r48zoOdGPR1nBnn
4MFSuc6QI98YCMfCky8xJ2UTJVDkbD4wpBSDs1wz2dEg00WAt5CDyMYBsGDQqrjVzgK/3d+y28C0
I/tX/W+r52Kt7iQW13PaNZduujBwgbkxhbVPnisFXFGU/YyNXuDk7unMxR43IB3JrM03Qx7Rn3kS
0FMr77zSTyZsohEyKUtM67cD7ip31mS1l69NpHrk8bLWkYtulr0V+RFFh1gGZ9pcceS1s70MKfeI
7QfYtzpw0T7ZMgtSa8thz8zy8iI0jXZ8MtO9h2eGwU2/nXcEStD7F++zA3uIP+HlnFC7SLkD1Q88
5NgPH7XTraoGa2hP91pexD2qvhsmUTD4xUaIAmz7LUpUWadK7nhQf2LE2F40d+cQvZErgQSo+A1z
/80Gp0kCWvQwoDpsjEwVsq+ZrqoF397ysKwUw1mq3J3QxEDBLoA7bNhgWLiIuTOcuxoqvyBaEIar
mvHJclASh0bwTImJHPpTFChPtLub0P4kBHYy9qQ3R9aar7Um5jZqlYIEhNhdDSJ/5+QE0r1TCXRT
OrsKU7ObtgW/8yklM6+ReAkXdJ6XZgy3l9ihwU0BCTT320Pq9xnsqRBU+cdX7323uSvAnEon+sou
rV48aR/tOPyaQ7h8oJvVqrpVSOKT8J2U1l8735Twi24CvOWhShQLjZ5lIkaEizjhm5oQ9bIRLF/k
HEGLSvlwLh0dizUjYLFDOiqZqYQo2q+gAO3goHIi9gE/AKP8ZHVnx9t3ZID3L7DXaqfzgLE2EJBm
EQIXNtcsYgGBQHcQySRJFHD1Sm1SCWhyXfF0LecT4Uj88o03AJPDX4hME9aT09FfK8olZvCVCtuW
XPBJ4AILR0tovm5cv0NQhTlyMMCrH3BU2BiK8Jnt/NuuPB4eTotn5UMLQsltFQp85DMqY4EM7vrC
keTkUJOPio3Y8ETaEicWVJrifZ5Vw8cEsOzG3Ff3NE27IJ13OgsR/1Sx5GNpODRWqi5yH8dIZZ7U
jO51wc0pYd/F2rA7cOtlRZgjX9Bj2TfGz2gJ7KsD3VHop3fbEynXXOMQiYGdz5RyXskJR6In2TGL
S44CTgRXbet+wOyXvlGxRGDBbESJf5pEaEDUxiGOKWaGOVPf5R64M+tgPCma8IZhYFG0QMHPO46C
URrdEz6ZxED19PdzHbXHdIcVLxMETQ8ZBYhqvk2IvUCAzOnP8h9G0cqjdT/O5K/g6fcosj/DtOk2
5juGDuHtDBzo0iLZs8nNgM9Orws6AHnudyXZAGdqsGGBNhU2AGi/7x4qMpGG8NZ0X9Vje16o0vt/
sgaIBs5iScRT06O/WApr/wi9+P2QIpidohBxy+i0SEJQlVF3YyDC7wTQAqtEoGllBohgFxpgIS5i
wkZ3qvGQXuse+PU9Gm+UpXw1xL7ZYJbl0mFF6ZK/INI+O+YEQ59xzjicAdOJGoPC3PGQpp3myy4f
tDsKcVWAaCq/cIuuAxd5WgnRUugATI4eKycXIBRQTB71/dFhILLmL0KtE4amGVwtbTNikEmweB+C
+cUFzZ07dM+oGzUOV6Av2eqGmEj5cQWRNHl69uIEDDbG9RpZcKwqxKw0lksJSRi8J3wCoLZpgoyY
PmJgGz0p+1TV2+50BHCPQw2HJ/SH1flD2bYi4nN6FGphF66bjHnMSsVs2c5f11PhotAlDzLof1ID
ibYRT5r12Pr7QPE3BsWQdZSys3xKlW0v4n6dWYhaNZky5m6TPVh//ZGTY7gThdc7dJ2fnLkekG1W
xsBkXaKwBLQV6IrgwSomD6Zh6rP1rAA90u3xYjnCTs60dcrwph13M+UHyx66b2UsWzdUwUdcMAps
mGFCGPqEC8k7WL04PJlzdwpTc7xyEIZeK8fDfg5gFJOedFq4umXL4gBcFpQt55XZLhdy5a13iIKz
f4d5xz3I9XjE/etJemuSY+AGAhBLRNLNK3pcFWkulAv5WgNYgZeucMi2h/jZE+AZKr4+sIBRZM0p
UpBm7EVyisgtWK56hKKBm9BKBNUJunipGaGKGJ2A3v0PxNl8kn/BVBR8s2UdDu+fXGJNOJinKnlO
TElnw7N4wsi+Ok//6MARdLINUeE956VaPt01Ozb/a8j1nS+qio/J8QGV/y2ctQ1z4fXevabrqq7O
vk5dteUPxt/laRVcEmNzSKhAQ7qG1A9oTZ4pezDUAtnam9uNEzx04eM0u6Gy0deXS8fPtFZOT2an
l5CZc5XXGOSg1uShjvac8pW2FNjpMv9i8/eaeOl8k4TDzstu3fhhNLQz4PNoTbMzf1JDPPZUrzvB
EBH8xD/aDgNiACW6TJqC+FVxu7c/hSSWGe16P2qLs77WgleTry76i6MwMV8P+/hLEhBFBFxX4qWg
idg6qi824srWEVK0UvFd1C0a2n0uqEVQeHfNEkmPClsW/B70MVa+TyQROT363t2kMbIzcq7qJolb
ge4lSxX+kPNpPWPVKq7i9tluau0s50wMpZXGRxn6N/pbhS/iolPotKDWyBfk1zFkKOahvxNdk129
2iHAhvpeNbN0xkOdENGxqHO6znMxzvUKVHF7wuSzsiPMJdmLxNmzhNa+SIDIfrKavqDwGQfMnyP4
afYMW5xiTvlv+BRtGNJTTSh9XFqdQy0GPUgP4Lm18crQAWeo78ssrcrMsA8HRFDR3wDvU/a7FJu+
n+nTHhWbRfwjLp8bmMRSc8mBxpeDZJyadXHGnzjS2AbRY6scqG8hTicH958XJN/OCHMREpka5Tnr
Fw3FHtLDksx7smP5v1r0prHPa7pPuHEoZnrwJFyVV9sxe8+3JVUwY/3CR7CFg+NnBjn/nttyxHp1
rkSMVBB9/cWysW/s/igCEgLstKzNZ1NtP0bFBch3QdzTlpJ6W2npY87YLpZ+q+9y4mQg1D+yLNDw
Z8A9/usr68prQXw6LuAUVlM+bQW5REVlhWJJ7qaDr1DTlRDVIGvRKQtXIt2jTvg5QRh9JYd70AOv
CKebvpJjrWaozCWNqEpzxIbozFwgwGcSswuwdGPCnPgn2iYkRN7GAReLRgHIyWUvdKjfr/wHgTcI
HXS0Y+OvgKjA+Osoh5USLISWgUD36lbeLDLlm/WkQZVc8G1HphJJQ/vPiYe5cz90wNYM7wuBLS3O
sO+sbM5ZgQiO7OAEshnxaygr2f4WvhBUeDzxYXSi60THPTdy/KRYm8fYCgMig+O4cNuX7eNtW3uQ
rCNPEedBMKXJpROzpPhvrYtFeiua/yFJg6mqjdJ0wiCo1GULpbiQKRrIeQFSA6BySBk3Pjpn1ljW
QRgXQQUMcHa83GNDDGGfn7NibS2+v2h+VVEYsQLZf/gY68WOvy1wMZcpM8h+y64bCN1ISR1XaDrj
L1Op8X1TpwWZrsJ+NOS8ueFO1uHrO6IGpIhKgqB52QowFPlvj3tOC7EEJIgb4JiKgfArGNYbndJh
tyoiyITv8+BGzqnmsnGWk8i/9/GLuLwMlpQbafQECTwTCH1jzq/AhZtrz1k+t2wL+y2Jho0IyYSw
mQTkG6C7I3MG9VyKsTicj3rCdsiFdB/E+uTl/gnEKi87NNJkWYmZdifhoE1QPFXbAndjYcu6wUZn
t5rxz/53iOUOc5AbxFjRqbGE2X/vDeuP8Li1lewuPlVWBiPLdj35A8vqfSY0AhvRFgeQvmtJpxqs
ti3Oy30uxsSAG6OAW05n8X+rvrMH46t/y3vrt7mXW/FjpyaW1Gr5riOvPG7wBhFfGtHIlyTG7x5F
mZiLkVIMwBbpu3XkS5aM4rEyNh46YO9fogf1lBgjWXy6Y2VmdbL+E8V6ZN/LLdUBDFLNa7kRvat5
PZ8/LRZjcyHZKF7PN4vzCrt6zKCTU+703RCEpj92BPSqPFKZkTaASQ5ahFcJ+QEulhGstNUBWKd7
iyxfWpd2zTJ7SeJLh7eQj21NsxBwjEJ76YNVdibOa6ejJt91ZM6zCdHwmJ8jJX9hKwLbOxjOyORD
KVhJ4fyJvFvTX99aVYk1shIhRKospE41SosIzCs5MgpcyHFJsjdvS6B6aT7gzc6Eiado3SrHVSdq
G62GnZ/oej7FSFXFcF98+ZylwlYE+K9mKD9jgDLFpDNnyeLtChWK31TVeerWUtJtd/3dBm536obL
kmUaicXGvX+SCUf7By1uaKjuA4eWTHTeLmA49Ynb1/GYCAuHnJYmij+P7aXsoXxyy8tdV1OSvl/r
3ePHUjaoDqmqLevofN3tRRSeVSgBstbKDmpGY9HFbbjgGTHmDzL9gF+tn5OBbq1m8OGt5DM0mruV
XR5qJDvFYDSB8oDdriDLl6eaROI3Ew2pHOTmfSlDrwJq6t0Ivw88UFYZ7AgxSelJWHs7Z2RoDsNX
cjCU4s5AYpireomjyZ/EWzT7iI4pfexjLPugesEGR5Cc9wwQHquWYZY22WdB26viwuXbcf9qPFTQ
oltKJXiQsMziYjv4OQ/StXS+/i7ek8EDrXwiACMTE+kbKrSIHAxE4ecsLKqOZZ3wv+Uo8rtGAEtQ
t8/bbs3IINWel1THbZbIXEcwCmLldjD5wOU6/tl8TZTCg4deVOy3zlrNOF/Xowx4SBO0JtnC5iu1
9CyjKWcbWRc6EuSW8000jTL2mq2dROWhSnEGVRStjsqDHFcaPzeaxYhj6gjytxcD2PabJn6wqI29
9eK6jkyfuH//i7bhlGQkeTxPO87gkhDak8P0SErqv8bKcUXeIds9ONVm6spJLmHjVeRtJ1oJnvq3
iNM8oEuNBPKId+zqwmwvmTmW/r9S0eNIBe71mIo4P29MzkoM00d+HEaM+EKgLGNipUH+8/TkRTxc
mWwwPqTR+J8mYO2GT1+KCWvFmlYYsPWjLBpRXXTDiEGOnupIKff5jJYredMH3irT0ZSzi0iZg3Y/
m8wZy5oct5DEun/NonjKqgmbS/x3BDVLQMfEvsMYA3aCTv+YJRDDhJU2jixLeH0tc7CLHTvCe7oG
zJXOtgqvwX2bp9kCBj8hRuFKGfEAXY+6z8tIn8uyZxP2S1u5VdSCExQMyHztHxmSmQsqWQEmz790
v9kbnYqXjztmSbpwddOSHGijxDOxs7n7hlI4Ll+UE+/LDVLx9ZHGCeF0zX+3Q7k/3SzPdByo0k+7
nsv2/aioCEkWlxpUSE9yWbqqU1QcjzO8ULlySF3aBYrq4EKKXNGPP8iwWuhM6fSpYmitU9DWocPr
zRVZFZ3u0KWPjk4Sul3n+tqgGU9jxETO51NS0GJRtulTdl6Z4YDPeREMBiqzQRc/7Cs5RsW4cx/8
CBwSPq+BiWkf4B8G9hZ7taPUjRl1Ox8LWjPuiAFulZwLPsvjsOmlHDxuibLOR5WYpfegjjpMrAZo
K8GiN/chBVVDWSx5wJv6J80zBiojGScWdfqi5t1BRaFja9wNW0tljQGMBoNvr4LX7LvHQpexH3XC
2EZ4YU8fvPLVMjTFE6fyzNXrPblQWWTFpF178cbp0WbDXCEHndvlF3G+nYRGdb2luhE0cWdKZyfD
y+mEvid5PtQSB5fiTx9satFcLH5jjfV5Tp7nMKB6BTg52KAqhahM1MtElrv3VbVXUTvetFt9coeh
29q7EW9zb2kxY45bUH9BPOTilKoTd3yL8gCiTtzpWgRfc7jUoacTMYT/z/RUchY43nBfGsnXWcaT
NV7szgJr7yYSB9lRqN6Cd9/d2MIRT2Z22U5jAhgi/5b+30xgYl3EDgdZpruxrNbrTw/zgC4CF6sj
KAbKJLoFtQcXlDwwUmBN9ZVcJI2+XGBnUFuJZO++JbhdzcfXQpbO7HlPuU9jLqYD2gmvvRfBRywJ
XgJ7kVimklu3A9z4jSrjsoeGbyhVI3FMsCWI/h6r2LPb+M2qBebX6PQqP3+YGpPXt2uohRqDItKo
Kwa/PDmybI4prlthWpsuqnqrSZMGP0YC7PDu9NWwalYRu1H2Ge6YsXxLRx2NzsbTczA6P/8d2ELB
2WAflp+zifa1qmFB7dnP86X9uXXJXgCu4yhkfoqxAj+s7q6j3xMQSI3I34G9lrm2S8j8mUb3JHLw
1kxMW5Ew9j/TIaWx4moG35DDrkW1thwvTavfdhJd9gPEsPdo1YWZ8h46ddb+MRnhm2iDe2jbCaiK
G3OeCDI6qc7uAG6jF/kmeKGavPn9oxOgkQo29MmGW844KVKjpUNifp/z5JyKo8RPL2og4fbEYG6U
OVP9/YAetglMP53/+Sou7n2uNORtoO3ae9oRo/nsl5V30PWiNCk1XNIMYYmWDBuSAvyyA4d6v2uu
yTeST7HQN4ddNirk0DJu4WnWnstwdBxti/bq6iNAAQWGi9ji6jr4sfdfE7o55r48BALegatxMfGJ
btWyIzrtv4jQ36Q7VEBrPIrfpbno5yjIfxCX71wHVdKRLBzy8hkC9B5rBOxd8l7XeG0M+Mg/NQSp
Z2RdN+qCNAdSv4v0zjuI8iiCYjl1FGaQyHsm7TPJhEW496zBRFPKv5BOh1QwMibM+lOi6IlK9uol
hjb1u9LapZPrzuAn0Vcrne7JztQFwVCvMyTdqKF9hTdgxsflVoyKM8qIsOg3DgzKP1DWvsNlzREB
edMeQaX7YetVKdmCeEVxRz8Zjz0GrtRg1sWTF6Rw2nMPravoo3a+fB2AYp/2aWDXpy7SFVkTK26/
y+zPhHQYq6m7wDcOTaboepYUHSImuJWGjRD0vLJCP8pBmGQSoAf9rTd+1vJpCUaeJ/zUrx7MGxJ7
x8t1UEv79OG2naOuDwDCghpTKyhNt3n3BOh/+GtPyWmUEYfqTu0o/Q33vSU15cGpBXj4LiuvFIiB
jTJQs577ozU1RFGpB3q3E8WgCbhFPAKKq9b0U+DT8gOmEPFLu66WiCAP0XVYTQ1kD4fJQEe5Xu13
806bGHwlM4Mt+GdA7bV6+KZl+cJ3melsDTnZO/g3ul0ZLmq2wBd39zzzBv8uUx1IljsgsteJ5iOT
O6zvVEB1XMYR+36T8caVs1JSsitn8YxLoKKUGUAzUsK8UZBH5XwZMS6K38pSl5DVr4jwYcKnibOi
P5rmJX2fjikRZ6/lEnZLusZCzOm5olOErFvOQ7YEmSA0yJk9n5ak+CKJHX9cvFWaikQrjDpgzyZE
l8DCoTjWrWB9jVICRmOWOxxj3uQXfc4eBZ45IEYYmTfKHWTGU1VBQQxuQUOvBLA1BbbVYqSgMHmS
bkjTTwXXYJLxbETiI59CRiGw5hRcgvicrBVW94UsEW6MPmzw9EtGQtFT2ygexKK01GuHY6rd1/5b
9eicACZ/RXpGBFyOh12okWq+4j5b3H5Qx/cqUYMYzQ71UiSlysHjl2B69bKeai+bqP+5KsGkKhtQ
mo2d1rnvsPNyzKdgOFXvWbqAqdurh1xyvZnGPVA5Q6intrJE0U9kS35TZOOHMQdRb9OtHoTDGCDr
ttbxU+1vNgddXUNLJGXWjppU5gmJVYJh4DBnABSRVs+OnMB+cIo1c/EwfUiuks+5ypFykUsEtBmM
s5LnTW0Nv6OFQ72+/0xwvGF0LvPO+Ds5F6dqXNjqIPOeOYhQkzuADV8ORYMA6LRRVwEXG0x57PO6
iLpj1y6JC5cCjZ2GO094lH7F9JV2ye/CkvWwMSZn0QAE+Pn/xn9RVKp8vcIhSqe9IePqVAJPV9E+
N6OiFgbllyghAzdoyKd/dKXhB8vIevjQTOMMrnKpwMEmmvQFW/a5eB4SDRGh+EcfyhAUNcPDFZQ=
`protect end_protected
