-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JVaOiK9ZYTBAKbH91RPN8M2bUf3TknjedXGb+TMvD5Jq5k2o8GwJrB15td85Hql4daaIsP6DVT/3
d70QTRRDcGTF0h/pdrMNYPpK4He3E1ljfUHhKblq7nnPN2hT+Rs38c+Z/Ih9+SaCMMLT8va5Cko4
so/fjRXWBEcwVDfh9MSgcqKSLln32e3glv5Om3xRyLTAkoRB8MHvwFj9R3Xb4pBtHHKgUhZfwOF+
Tkj4xC33he5k2mGOHhmSeHiDu9Al4TExCs3Gr39Ky/J/uhAKyV1kzHUkKbq5BEL7erT3Ow2UztY7
I+pfyqumdYtZJ9tYsI0EOOT+pvj1Sjmanoq6eQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 82048)
`protect data_block
unktjuL7XE0XsmPV8/sBPte595MFulD0YSZ+GVUamE+Jwm/rYI5dG09IlTiux2xoTUM/3Nm4B9aI
VaWmUWXEVggh/Wyyjd+xGmmaC0D9KFIt7H3gPYU/NJt9r7XwgYLVRcXnY1+fKDZGqiOUeCSeocKm
a90D+S8IK9J7aq/OoCByPeIr297aRIkYPTfy60/vIJFfTpHqQZ0a5450iNiGQOb1um1zIt+H5wqV
89iDGWOeDnsikJOl33k7xmQD5MwmbGtBlR0HtE4eB60jvATsglvoJLpbZtgb66u4GoBTr8ExsXsV
rHt0SxPOoPlT+sNLX9765M5xHvSHX9aAc6ovH5MwAODCIxqysFjTVuDvlD88TMlKVxXe8THG0UF8
UgrFEeYc1cbXK7ypyJDziRngjUkno5vw38gPbFzzcm6Hx6Ra29qv534V/H5Y+enZ9GsP77oAEShl
raKz68pq6gHFRAjHaWWEEOYTjnZZ91+cz9uN6fkWPEA+RvVNiLEnJ/mF+o2lMrdwN8x37vD0Vybj
P+yiuphsqHKzPgPl7GXnVfdL5nZ31QYF+k4cg58vJbT4e+EM1Enz+ZFG3eHqCICe2UZgdzxwawY3
Vsjo9rvFbjKsNyw8fQDrsZcpGzNEd8Gddt1NeOqebICRumkV+rDzlkZJo0NAuEd0fPPV0rk5+pZW
3VGEHMQxcZC0ShMqRF9HrP8WjqvVzr4aFdpuwsTIYa4qcEuowqE6PdE686Gn3nOj+ALgS191cjph
NKiWlvWJlRCIkvAskSkHGssasmQSySY4tgudss+DAuDhDU8ksn49vUfIc7JWIHSF8hhQ/p+EGWIS
lpVxxRKAl96KTmPVF2ZGTjxUz9Jo/ox/w3tZUr8L//lheoRr5tgLyCq8RE/1UlMoWO/O2ULlCT5A
an6aREoH5KLHVKIRYqHWG/B/05rwlOeIyqPWnKMuiPpurxanTSPDwc0wYQql6qSlbLOa7HRlcGr3
R3n76kCWk344SoY5YDKP0XPBvCJwoR7qJAJHA0gOsmGumBeaoDKziRSUz+UQPVoKfAgSy7aB2o6d
rO7gSKOwkSANasBkMuXSY02SxTlsJ0BOAqBDgwNcb1gXh4j3LAYMVVVkA+6JXR+OJyV9yY19uWvB
6MrevizgG690+uOKzhA5OJATqBdNZSVj2LgDORMkD/21NRAoSobLG89vCeDz+LFR3ymvS1T55+5U
u8MtVNUd5wpydbpdzl7vB06Ao892K5gB+xrBtzo7hQ9D/qXJI0jiHSqrUgh3GFm9euxWASJxdezp
sV2pjDRcK8eH+E+qaDjUtyAv4zMQZSTbR62+mWbQjFcTkeExYXCvTQtZiToN1CDqr+nwgD6cUFf8
EuSHIvhZ0u+NrsqOrT82vifqQOR5Lx8KpqFY9AHgsDJNt5Wn9okJjyfck7oP6rhuABZYZPXGNIMX
ToNQjajx61V2UH6Xmc0zyGorV8IpSP8sb7XZrCcmVA83BIZJ4Y3pFOuHnpHyDDET/rQeHmX4/lqI
8CWL9HrO7YeNlxY7BruPRQHazA750TdR57jc08IW7j6+nMc53H0tL0vEVy0sUvIrOLP7JSd5e/4g
CLDW9S6ElRqgGzj/y0N2ya2DTiiGxebwCAut03LuGT2WRHYHHJiS6tKWAFf3Jw/VSsW5SKYj0URJ
776jsRDONKhNYL+dioanZoEOwY+0BGXQscLec1DhrGSwcyOGL5EErMLlEWfMhO+eAFHPvbpR8rsq
q9nU6XYu5h8gB2KxXv/9I1CxB16kbR9vwvKOcz/IZMy2ZrjkkKgdZKLEl38zNYXMStQeoHsPfL/r
LyXov4cq5geKfwJcmVhn/FBnajk87mp705dkecvIxM02YT5aZzfYeYdFQEqVl0So2TQj2AnZwvlp
Gi0wEIxEYPvq9j0rnYK5bolXqGHfRayoFi9GI9AynoxGfDpX4fGn0gLtsBegRU4u9Txu4urY6kVF
BMVgVv6P3QdzJybN5Tb3sk0Ee0XAs6B5/56vBFVVB0hT7+qPhs252cn1AzNiUR+rvMldA1V3O+vD
fjSq8oo+EcfBGfw7XeTVq3fNhGKLYmsnKWvBb6mVRFhDRGlQkSvGxHwMegT8m5CqefkPMcshsSev
9xhIss/N19QquZZ9OZ/E+JpUKJfIs+lLrvDA7eFKoxw6zn4q7aNpCcTc+7tZGy3Qd3ck2821tQuh
46u5wP57K8zbaUhxfv/jpB2zLzYa6T05YR9QPNGfJuNtwzivj//Rg1JQe+HVpylBKtZtKd3cGsW4
nOeeNF+lk2+kevPo4nRXp3olj+9BHoITGaeLtAZpetpjECCgLFxmNK2hDCYAwsMpJhhtdFM/76uh
/c3egIGo6uvMNBkAYe2OnZs6YqafF4zAcV7K0HnsH8E7oDxQYX2eBi3BfC3fj7lFoRopYzCHzoX2
xbnn1Dcwp63KF0oLL1uv3/T5W3yYY1YQhQM9wPSl+4vdFbAGbEXj6m4+Vrijn7Q8FTm5wR43bkCC
rKdC7VkvQ9/+/9eH+JMPgccx/itQX1SjDI8ZdfVSGiNrbGR99allKg30MZH6KQ9f1hEYR+1x4Z20
n39O79PYbpqfcRzqM2CCmWXNCirFnUG+bi/WYf/IdA3iT1LZzUOiVfAZdstY+6Jl79jdwc+f1aPV
exT8iPI/efNZP5CKf/7FRHq27ppeJz3tGEI2xAE7v5d250yf7a+ALvrggs0xUG1GoMpvZw+wqtPV
+BjdTN1uLStqr1vdT+s4602zgIp9rGmHABrQjsXur+FGssKGQp8tkLw4RkbIgvmyxuUsOaKuYE+A
5IsvPt0LIDCCxYiDiSqYw5CtElPMyGllq1uWMbFXreXHs+BwUsQYwQOnozwbZeL+U+UJgOxiivI4
JSrs0myO1WFzH5uTIag+309HewX0noIsfr3IKe/HCOl5KgNL4h8Qr0uFa27eSszellHZi0FPZ+L4
jQ89NcWF21NMdkrEr7/DzOS4CXUOD0QtTzcz72g3l/U+Y0vl3PWnqq3J8FQrUNU211yDIhMj/x3l
vPRw/QLne77fPMhlR1wlpvvAX2QF8lyUmelP+9S3fhRnPrVwdzDFK9GB0K0dcRLQGvzQxrveA7O+
6/DtXYzBewScVVto8n4eNzL7aZYvk8OjnylpaorJl+ovCc12qTozGhCwZ/asiQiGgw1/oNvDEowN
+fUGFCo2N0lnt1cmphwJLF9vFSdmIEnBxJElTu3T11mXlM8wvzf/xTBhLO6oVuPVs0+YTtjkCOGD
HaaS9vSV/v6f//PD9Y4WriIpLNpjekVX7+AazynejVZ/WX9Bdxk3Gw/aNTxZ1DVe+EqYNmVnxIDJ
Gs/iD8TTQPpL6birvJ9BzDuYcNXDBdMrdEoNiveoZnBjSJpY33bEbK1wsn/4s5i3bqO9BaorJ6D7
9xxIdrCpeCTzBKZHVOzT9BfqYIZVmBc4UOAcoVysWc2ynDFfF03lpj6lOtN55zqZZGK+TWsu6/jm
5MaUzu045ttM1ourFHp50eJLGoriAY+h/9/cyHrBneYXdQE7ECR9of1kvyrPscMDrGEhxaxRGJsx
4eUR9afZm/m/gzxj3F0yZV539yU+6MOZmzMkZLxniT/UFmGLIEjcazq7vI6CtlI2jE0C1xdz1CnP
/dFdBpc5qH3VrlsJjn6HeyUw3/CYbhdtLxh2X5bU1WCcw5nI1GTeMvohfCwYQlyjJrCOGEUn5xL0
oYzkGIcI9Ok/LzgcqqSOluWoHtt0FvJdtmvNulhRiPvxSI2N5mvgiYwbMxkIUp/1VzVuE8zsygeK
dDyy3W99JIxeI3ikAVpa3M3qbRp9dz01104wxtLg9r+FxNSajxVxQGcUqhxKkAC+jyw3B5wlDWlM
0B4X94nXuPcswvF0oP8a2ceYmVZcHBvleWux9OESJgrgP1jMH700HqDO6WoWRlFbgENIpNF2DDd4
HchU+1nixhIFYyKh8p0jTuigjyG4GzcjNVZouNI8Y3VvMwNeTDOyzuHJ8LzaJWP/kpixTTwvx6fi
PKLsQwOHR94r/1EiDzVMJraZTprpTkcUPm4T+hTRCh0BFzPIMKB/dpRllpjvuDOOwAIby/uoYU5w
KFAKj9niedz9nZJb2M8bI19kZM6wBnaPmbIdjU+kODNpZtVAwqqz5pQojh/yWbFG8RYQQKExiwwi
Vtzf8YHqOBW6emM9gON0fse27JfIx/Vp/ID0qknvMUiNa6QJRf0FOvt6sqo5mgcmFcIGuNy3fe3l
ZECuisKDCPGwV2sN1CNn3u4Y9y+8t//ZDyNhiC7uxn/PL0KQSkJnzyjSFK1MGfVKbW72mbOU9TTI
TB3nfxvwGNlIYBgeGCWaWXWG8oFMr3gNxvcWY5IZuh51Qh1Gd81Zawk4ghCvHKEtYKZbbGuBYZj2
K8zVxWItt4n3vwJRtBcGdVbgL++R9u+6QK1bsSx3GxgvASWLDhKdpSzDXs9WLQFAq2A4b6a+cUko
d/yqyfk8/YepxbLnaw71n9Ia+69aG+V1TayQd+FiMKs9g+8SPgjIvi89/ycbp4BElI7sMR2PU2nG
OppCdMzgnQGoR7oBucNPSbW+J0PXaRiTd8eC0ngyDiO6H4mIsdSq3Ra//yw9uX8EUyswq1+ct+tD
NoGisnjSdfoY5ZHA1oMpd2wr3OV/4phhNnenBA3O/2u4vo91yIBe618bXwNeTHJMnW5ZyipQx83q
b4+yD50Un/0WZxaeB7b+okY5QZN6i2/PVWMXq6tuZfCJI8fLYuPwpFgAOvUQgU1ILPPSBt80Z3MF
Ue9BPSSn6ZgZtOLVK0m9kQlqIKQfkCeL0U5SNNZSm1gqJyNxh3dqJWs1KQagKkR+sPnmKlqh2vPh
+w2z14jDA/ZzQJm2lSAIQ3ltucAd7qDmIQVV1qBnevHUsNL2DOTTKonBlyrOJV+06VScxG7iCe/V
OBDwxGIChcQYFkAnQyHlGZflh+zUrw6uMKkAGC73z8Y9H1zaOoyTVDGq6d7HylrAeJgDcvpfx3dK
QothY93qbU/zKspAWaoNkPLwLI3XoYtXYzv2HpZmkoq3AesUkC0QYqIUIu8YGnu3yPbNBCS/1tel
4KoIAJqD7vGerMNHtIbkUHsH3yi1NQKsCmYbPmNzGPRaARIWK4kbTMC1qW9jLsLUFhXMVQJi4YHu
8IcjcRyaRfiZ06vgOBih+aJJpCSm8Vc3ltfWJXrotNWCo9pVjkgS08vgmNC8ghEpfuNUAPZiGT3S
3vCiRIOj3sP/ZP467uDjcVedmtyI/EOVsz73nUIPRVUKwlOvr/VTbTEQotpGGkhfV9ml7w/hb7+8
/5r5u+xLscqvfFJdjb3nKczvlF9DWTRFxgEgbBUTuuTcmrdmAk/yWzAia7wFQOomSiCHRliGvvUZ
6Snpirs4UuFYALa38A/oYZx77IACmQA12+/U653e9rNKg3xM0ZvMxi/7qdw586wnF2JDii9wBqO0
l/gaZTZlD9hb5opNZcI8cgDZ8oMNwJl/hUgo3brgkGnv4Aia6Cq47y5AAKRV/kFqd6dCW7fgPGNB
wX7DxVRFtjBROJuq9HBYGSzr8ErVD1/pcRAWGNF9hUB5KD25VgGKoRiOsQk9hPmIqj1qOG6c7y1Z
Hq9stGLsZKoHcoeBOY0u7kw23DVP6/XnC4jq4ZhbRK3Qbdnv50FPAU2hjN5kRHBjr7dV26gsliTN
0hNapw84m+MvrWUVi0geKHWTSn+GMhNJzCDyCtuRFHqRsJr2TeMdiKtyuFmevh8+3xOqfiWpuTrd
cYWNC0EyxHUZQO69Uyyk9poaXX/rg1ZftTgwFh/ceLRpfA1UdmvQ+CZV7lxDHuCPHjbp4FLXL8e6
PbsK0qMgFEvge+JkCBCF94EBaN/XEu8riTXiv6D6F3EtuyfYUeRQI3Xtihy8/UW81nmb58iWKiC5
cwXOFJxUhzeIAP0jX0065bDK1Q6saBFsopBOBdGDNRff1xY0/9DCUku9qA+n0/wsg0DyHnUmueMF
sNU4Niu5T1RS4JwCj9QSl1NZP50CfvgK+4QjrUL1+5qMzI2OC/mDqymLzoh8IJENcC0l/LyNArxa
bavRDtCZg9EuyzwMhlD/z/filRZIUOWS+p/1igBxOjtFWXJE2+7RnaoVL2BqmNEmJ47l1DJET2ZM
klj27oU2YqWgmcZlGczf6DreCx4aRx8CnOQ5Dh39tyfNYtm8Tlubw6HduZMpwCPlBVnNg1nxbEa9
awvJJkNIPhd/QndIwkuNUyvTT99Rjbnss59gG25vgHLscCLe4FKqgkwi7iEz6d/UYmE0n3J5kXjM
zOAf6oVqe4kGO5ZOr0r4dtyciA84Hmfzr93kafgqDxee+dMgp6uxpRSxwt4jGgCPGOwW5vace+ZS
RLZVooTRBbYtR8pI09IngnNtZJaOBVMChNIlIauvyavweTPYIp/+zAkTqTF2l2SPdLHD/14ezkP4
m7EpuJNnsvt4SJXXy8G/RbrXMZ75MDy01cY/H7YlTkPrcbWMZm9U83Mb9rPudDq8jwC8/ddoMn9c
1x+IsDAoAH+fCoJT2rFsrQ9X7cH8SOQjnO39/N/bVk0s3ToAafmwjrZF/WmYT5n2icsYXzD+QU2/
KIwkbl3nY7cpz2gvnBxdC8L8InI1bEGf4oZ72SBRfCRrpD2cpjQYzQFKq7UgdMh7V4RZocWsRljg
U7ih3p/6nxyLZBPqIfbNFxPdmbZTIxCEypNnMsCr54JbxHbgrWYjMgms4UfHY7+P1QAh9Z5iSIGg
emf+nf3BFyWuZQXfrQukHQqQeMvZMKT2shMhI4P8ZbqRxvX66lHvXQZXvFALF/bNuqAdZjg4Mjge
f7QPurQTIdk36TQMhSBgVglk0AYR0CnVI4CQBiSMiALCsirpt/WedpVPUJy2oCbgPsmoN9tNBCNK
2GNf8AiSMkRAqEQTl+JB4B9zvM0ilX1NxPK6KqgZpDbOAwBDGtNyEK/bZZJgs3FhqhFz1G4ix14H
Lpmq45HzLAVkbohwhgwoAS/LYZ9NCpjNcV93kChC4igP+n8LCYuQDrqLmQr+orhFsdb/sRB+tSXL
nfvYGG6lTw/lZaGL0egY9KE49i8V8T8lqXpJaonZ0M88DjUqQLmjnZRvdoAqyLbkHpaa9s1tSDo2
hdjd8BRW9hDPEZvWpDZ2K1AemseZcTnaclMmIf9A0afhAs5/TvIPi6RiKEH4NfPDt3YuLS9Yd0gk
ghinaxIjx+H2g/8LKLHpcHJiyCcJqbcAgObg9/29VKIeyA+zmUUEtI4JUPG9qC2/TB6HcuAUH/OK
kTj1KS8zOuAsBDmKpn5454Nkhk9wLGNzIddZwuoCNNT1yicFBcrJsTIbKxnNsMGgm7vwUL27Te5S
jJCJ7YJktmBkc3mwZNM8V5vwN4CF3JNmGZheYppvnxNjOYbBGkLqTakcvtDhYO20ruChCPUUa50c
Tq7YzuGKB91cvOCczd/Uhz0zm0XCciFv1xfmBmJ8Ax41rA2HhKQPDIN4S4L3/2c8rK4WU/QbZdL7
e9Vr0IERZd5Wb314VDu97sx9WwhV7ZhmGxbbhDBThEHNt9FfWOtpgzsAQqV7fHIghhOHIYfrQBe6
bw2FyAGh82OZy77dvLLguDrk9mPd+evjmuSxdeg/TULaViaJbhyrsvblsKTDDL5jbpDm1iPrjkNJ
PUp8GAsBrBBCyLir/7ujJACB/kI0iDxN1Ovcp3C+dOQ0miW9NQHWySkgm61HQu46kM0yKw+h3msi
2hd6hyT8Fkhlb/vdvCXVTqA4CoTEYs49j2ovgE90Aiga09gnZdxIXyF32mlRoTbSacVGtPPoF87L
gCa3hiPE50CE/L8NxLb8l8KpgEGgZ0rLL2V+wx7UJv+rr+gzv8hVyD9hGXb9y5IOqubAGWF9n0R5
kg71l7+0JIAsTjVthb63GmFeXA39BlJa4sSNvuXVm2JZJQLCfHvlUXaAknGSaedSE2lR7pa5Il+/
GOi5cMxH+psuMau7k9kpXQUG2Vcumz2RZBaoUWc3WGoiU99bXYBKAXtszEqCQc8Zzk/LL4yzS4To
6aLWNerubDg1qZMYCrrPvJmPQlz90gc0GtYvJ3i79Mzo2vT9RZeGfkDY9Jk5fFfdsV1HMqNvaiHg
sOqLEhbV+dvxlgBdkU+o5ObiXYhlbq0sFQISkPrV8hjBEtTInfOTca20Vq++juwTy3JuT36h4Q5H
xeShVo0loChLFq6mLpYWkWwMGNYoPYYmBhAcy2okI/1euQK1kFLAynEsqTiKDtK/ZaECnc4QMaXL
SZKonDIKvcQvE8l5gCgkbbo2WzlhsXqwVkLLLCEQPpJg8X7FPhTYPU3vdbpJjQ/SAyDLPdixXc1e
W+4wdhiVTkBzGaDd5LVmj+zHatl4zFbpkrrfgu9Ekzcb0d6w+8CnUZ0sRivBu4x25FkKpJkASXOe
UdkUFQIRLaKJSROf25PqEq5RT4uvwLHyU2LTHXSz539bzH151FZ4PgJBWD8hfHWmzpo+ErcACQj6
mzTh5eBXK4Tn/sBjswJAJjPhZLFzQ2iZgGB5IGC/OgmGr8+i8UKkp8vnMpJ7VOMd+1K6uHnVVIEE
KMoFhQJ8vYZsUT5evie+xGqIKYKsjLTvyKlkMnSf1CKp5bjbB9h0Zw7HUH+zfRBRa2pmPrfLLV1S
RMtKTccYYgeX72XViLRXOoKsW2x3ZJcC0C8UVw9iYyZHT1HjEFEQg0Gv3FGZUZntojDlqpCIxdKC
PzBP0H/0EyF5671G4PZxxK0+q99YTgedeEYcS0iC0zJZav+VQwTqVBSXMZ2qUw/6GpGpg5gbWxoU
I18owrZekGwtX5iVG8h6BGD+HvKuu8gVKZd0cDHWMCaSRVontXk5qrDryoTQf3sj7C9nw+fQG5xj
Fr782u5kdQ5wzuTGDRUZWsdTx3jZv8Ioc4xc7ojLeRXdtUceDeuZqAWPJsWeNpWl8Bktr2u+ErGJ
eeFzrDlscJ4Bo4BVroFrimrO4YzIhdooESWjEuBtYYF5BSpA/Bd8zQzG/FMHY17Udq5dreCUw1XB
UJiAV8g2zE/hyd7efGBYRMlyX84idvw8eWP2Xg6QgqkhmPuRDrUDjXdGxajrWdf2OcvgACj7Qvhl
SUjdcE/a2I45aZB5q3T01rs55guZcY65deNZC/pdbTiDKs3tPnlUwhhr5vGllSHnUsyBDfybX/cY
8iYEElI0kaQNpGK1eCp+pE2/BHXoXFsqB4nfkpiUUn+evz3VQBIOSc/vOjZBZrcxYl2R1HtIhTOo
EGXF/VhRihvNn8ueAhceKig4YgiND/bXYpaVDdvyNgiDAND5w5TG8j9HbD85DlO9hZyhCzoX/JCp
T6cR0A6HRMT81Vfr1CouZw23e6wWxfTnx59iQp6fT+PG1J59dJBpR63Yajs7QpKOLUtRTXJXCsqC
a+k4Xusd4r03u0QvywmvDS0lzqAYm8LaMr1ScOfJkKluaVJoVA1jUo6tzVHU28133T4kHYAaAfzI
+EtdWvkn1e/luru8iE7VY9vPJFmwN1TqOdZRy78pEaOsl45JVzsWnXtBJO0hY1ZQEhmmTdkIIFrl
DMGZJdqKB5/kSo7qcDdXJVPUsFIRSHXvQ4OIu5bXxuogQa/b1LB6wH+7gE78nOidMhN2CreVNsOk
jq6ASxnygW0Xp/0r7hcc6UXYvEWQiQvtp/sqBjnwOAEZVTmz/fxWaoPyw6nry7qu6jNgGwNM0q/2
1nitVZBUY3vDgdW9GRvParGGrcwDmi++T/r9/XXPs0GscNJ7FTxy4/JBoIRls3TYgBFLBayKeRcu
lJzhcY9DDzNqX7i01O+UJH51qzOyhQhmHbZGGVCObDQR3BpVdV2caWP1EHiiroHevH3I5jMTWxCV
mrgpeCluBXl5zXTWrEgXHeH2fYz4UHaIDpga0pbZR+Q9gTYybhCid/7cOAYbzm0SuTMq4q6zt7ax
XmQzAPT8ae2geHiZyO3inWHyAUxcgHXUoGHIBfrJli9Uzvo+MgOOLjjTS+EyZrKsm8fWxX0sRfM5
QR7ashCZbZq8c5lzlKY5s2HkR6n67hf1N0VQoZ7afWab2QS/UyNYOfq2/JbWMwDkC2PAZqT4fJ/e
RQI8w8ohJtMQr/4b4JfzWPwaa1OUu+vxgH2fkenGtfTd/BYMjzGIDK4m409Uh4p9B1S4ARDc75Ek
JYjvM2V5HoWAW/KSf0qLuRLTq+4MVjb0zfhnDB19r+BHtTsnvJvPmzIogBElfyyBaxCTDlV+is3m
bPCbGW/Zf1AB4mpjDidInlgJYEfiwF0SqGZUpC+oYW7KyTiBlCyDYWyTISKFta3Fl/0TYOF1Nnfh
gwr7sZEo8/cJBqWX8mQN2BAAVvjUL55rzolmPWs+Wz14VA2lEq15LjvTYB5mH4At4m7az/ipPSXv
dWaDPThWrPWLoWbGbR2F2zBqsU2+mRqSYddilTcdlqASW+BV9VckIuBVcwnRhrHJhb0p+GbqOoSd
NzWfsbGm/ZytV9DXgp1r+LDqxhbB+G3YGe8yz0AUlp430Y/B9ABe4hT8qu/FcSbLEO1keFC21Zsc
vB3cPf63yuRFDe9otpwV+kuxoXujoySinAFl21DLhMFPo0NFu04hDoaiHUIdFpn7Ppf47RPgQp6z
uXjCSQMg70ucfjJ6lkIHNnymYhtJX5Imn8+CMCcVCyYFOxgcZtQEtWO87Yme6sY7LLplo5VD9MCF
DixCKI2q1nCdJWwYviIV5+hNBxUnJqFADRA/JNM+uNwf8kwmLpfN6xVJWnUYz7IUsay4zDgmzoxt
ESysvH0JLx4XFewjWECgPfWW2XIodP5/3D3ZQ9iXZczNaRfTSA6HYKJvtqKfu32IRfLT04hkXAxr
iwviYJh4vTbBVOimQGv6O1Oj18ppVxez0S8rHloB/L1GEJNawoUfpNZMyxANWrxG9WkBO5WKEjEf
5AWqwhHE6u2kSgrIUQc8yU59eFan9VWTurAmOCgCmIuF32bfplUqBsMrvWPQz2wlKy0Nl/7KkjyZ
vDQElW/vnz6UeYeiEL/xM87XF6OyRu7uPZ15wRyyiSjCpIjzBGqQyiyRnE+LE4VkCToE1EU5qdMW
X04vaOqQd8zWGTX5dF8vMoCJWYcRyJNKZthNa7haNn6O+ty43WeHkJq4Wp2/OD81zWqVgE8Ybex+
Zw8lwQMv2edXz2ya8krc5ntY798wQUIEGDtJ8+WXeBAElbtQcny6XS24YTaaqZaee9RRt6zSd0s0
qDNz0W+QpmHLoMG0B/5gLYscykTEUeYCAcYnarodGqTrmZqHX90k/FNqx82BUUnboz7OXgSUx53t
8ctnquR4VpsueVPy6tFyo0vh1+tL/Vgkd1ij7tJrPm3RomjJRFLb8TUVtfUZUwLYbcap2LQDfxQh
AqTd2GaV06z8hnwE1/blUGboWksflYz/Pnjl0bKtl+JWsHQaDeOQt334QzJq9SYte4e2ZXRY3BQO
9Y4AK3g6wUWGNuD9gW5Z/tyQuXlwZCuuYDJQKOqjEJR7ndZLYc/3X1VlwaodkIQ5dktTJtdgbTaO
RFqCgLadeSOeManhSvRcRVPdFyd4cEaKC9dLc8v41MgxbLEPYLLnQLbQVCSLdG4FUsqkGKo2ra3w
iSipExcMp7XbYFVr1MNpYeOnOh17M9Y2ug23zw+I8vzLX7KLej87057dEbJDkRRaIdHKqe9AKVQQ
Nxcnn/hNbAASK3CM34sy0QXh4j7nZWNzgMMgRIGAJD2bAlkO5kuuXt46hGqKi5KXSvM9RGVpGHet
MUmzVXR0y/4tuDDjnAx/6RILBALAX3TmWWPjJnuqIlOKbwSYGPXM/lHs9itjLcCzFdAZUcS7ya6P
F7ZFoewczQgZyUebluFEByBiecDxuGkspewmhYgCi2exFF/RGjdo217BsFgxNqKS0WzXgkUMwQfb
7Ex/voqLb27glRKZZrDVcxSTN+vuc2FS1/ncxesoQzyJDRCHx5E90n+E/EVw0rRgMQMdt4qZu9hk
I4va9Ff0troDYXWdcyqTKhDwEmuCeGccjAilA/hkeLCSa3EyuGDNTwLU4+F4Y7Rhy20JT9d+LR6O
+LVlepI79xpxaxQRGq42NoaDVUFAGdnH88Ml/bUxgM7v48fl8yQkG1WmYsE1ImFw8eeXhYvh4LtA
C+XIqv6dVak1gtWvXLO3boHe1SqW7Onu7ogSVR6DFl0vfnlRvHkNOVIblpTxsFwcByqNv4Um/XMH
19c3BV6GgvkkhZ2ZKwANtkGJrN+AZSqTMIVf7WiEojRNqh4hmm7lEEQNJ1bDMPJTwSSQkXQzzBrj
AEwthUQyzsTWtSM3eX0EoZC+MZsQhCUWp2vNL5D3zwVSfYzV3eIzZM17I/x4q4jGfmW9bie5KxGb
uGJ9fnmHe2b48q2+ejMdtwEnGgusPlrb4a9p3gStQtGR+NSTq12t9UrhOouIvrDL9CW+CTofVxcs
Ogk4mMZ+DFIWLyb7ycOvGG9ixSHFOcB4ipzg+PDK5iH8SFj7MXnGSWb3F7bn+I4i0wrJtb66FXdL
9rAT7TA4qt72BvHEJrfaL61CAXPBBUQwtOAB1np1WdBRc98OI6swmXxopEYbjFUOI7rmXTyhUpuh
0OebojF1Xh4Ucxp11Hh8PMAOXyPajcjOeX1C58jYxeLdkX8v2L5zynkCUyN3eHeES6Zz+pnZndFG
GPCGnmPhcQuhFq/mZpMxRYqRMsCqQXrBgD9HXhhmEZhF+6TqvbZSAmcm+Ithbnh49nmvi1j5FKQp
hvSosZUMLZ1Z1TgnSO8eJQMvXnk2Qe26nS18x97ne2tXp5PowhsviYWGwLLC71GNcz4JbRIQ6bJM
P5wHAhtOfFHS2oC7Cqem3MoOTWT8WvNLKu9jrzlEJq3KXy4pn+R+E8zPVSyl1fxH380msjpdzkAa
WBSh1PCCppC+k5hBbw47R8Kd36qOdx2ZhhDSOmci2OW0lgbBhPM2oR0KME9rjnIWj4TPHUH0v5e/
ArpWsLRxthP0H0kW/kQrWXJucxN/ZIBE3/wD7FeQvlObZeA+ASZ6PNu4g2sHIJ/jSeGmn4QwZ4sm
a8wcfN9GsECik4rjib5TKnKVMdgR1dmmo/tNbtX4EvxHqh2i5uQcyz96TC8LMa90pHc5APT8ONLM
UjigfAyB9/GsXatMLiYZuJZMG7UfpvC3WdIkqdYYnSbwasYEcK0cesZVykd7WJSUyG8h3DZJI7Wd
UZcE/hXBIsXGBKCzvYMQ9Tuq+r7HdMEv7bXKYyD0BhOVyvQ7P4HC3LwfIIGYFdcFNXwyX7VeBICo
BfHwkmn0RH1MFKPRIS2tImR79LnvMnHnZhoBMtOP6UTBhdKO65BCDgPkhZdjlsrAMtqv4YXwvrrV
LUQNsoiRKeh/WhNXRYA4BoX9gMNfEaDAI9UHaL5GNNTE9Tke+WvKd1IdeOuW13oWl1vBzSL7EaBu
9TE8drugHQ0aMv+D2LYOcHFSt35IDb+Vj2JfEhj7iDmURegnMc2IohhaU0hzoZ7tipHKRVD0Wqbj
ISkieWJ3cOV5e1lXIJW6fRAlSgT69SyjEu5W+zt/mwOp16WKMQ0lvdMBoKrHFfZ/EJQa2qPN//uY
U66rFMsqoFrflwUA73b//ozo/kXWEZhSAaLFBVYiDLWPeBWLTXzSH54zwRGmhEyz3JitMAuT+YAG
FojN7dJ28y1sanjyz9EBWHybUMKbwMINkJkDnkHeoxRTdj+jevv15PbSYRS6n+u9W61lTZzx4B2O
pKGSiiBqOLJnuW3w+mecGj4muqazmPj7zooF/VdyVuuemX33z64kNWwp9mtSqcLHL1PBO1O3xEsO
QmLBAiF3rrE4nz+Pj1HVLtKIsAaS5G1X7+oj++3+7gBp3j+FZtMDJhiMQ7r/vIEgEx0b8uBdMhfM
qSL99EENxFw+oX/zMldUO9/oZ924oNfa4M5YxUC/gifZiEt99GoFdkzsPZ8Pe4mD/g1IPBW2x5EX
/UrlyYBIFgeAxjUc1bnkYN/nYA5ydT/z2Z9dVJCgP7UUJXsPzpGBPkjFhbeF6n8uWVe4y+NwojK5
VxADeGTT+rgRSjgPHDH5NNL+sgZly81qfISiDGGTVRFxLmQtxsWvdxtqJ8+Ijcl7Mk+zZqsJDbWb
CuVnCJ3QyNUcezSdYDnFi8a75SJDMPFnwUv7s9JXhB5RM8WCrKyW7LnlrgsNReE3O3OYVnVYtJ+V
iMiOXFCT76oDgE/CNIu/OOBougkJyQ8cClFgxau7EYTrYRhDvIO6lc04z2iuXtI6GSk1Ofh6HiK4
WsZZzY/V3wb7LDPdrf1RDoVRwL/GQgbIBLChNGvdmXawC7DiG2UB8IJ/YGJN09wEpizamLFEkNjf
VREtRCEKBYo8FONFhth79c6+S1cTfh//cyCG69COpexw67VoG/IbCsGeqqjKy4yH1bZnen10SW5s
Ia0GYeiNwlHTkg1OJQu1JHUBBDkNZxIVNtleKW7ahDlR7Oz0qEk8qihu/aYSBizAqpdRFd5X2xYG
/p1NkUwD+hPjoZdLTVkdTRtS7AiqcTUGm1DL2NQCV1z7cpsQpRM1I3cst93nIge+W31xiJzDQ7Dc
H/KvpxnwW7pBlpxZVeamBELnR50GVLYNA/szqZbl2LqYOCEjcqlEr9SjN2G6PaXGj+Xbico2wo9P
1Iit3j+TNx0LMlwhhUyGoZf+hrBQSM28lIa6Ber1cvencl2oJ4EHIulSMTdyb+qJLcOjNeHVbQpb
nSeMM8ooJhplFrgF9za0wmq94rzUaSDUIvsE0hH/BSLn1hLZAHn7gSV5L2Nxx4JU5HyMb+fVKGD3
6/KdRlTAfRv40MTKGfZ3xQre9FUnXNRt03hiMfM1pGMgcyIU1AWv2ysCGXUzKf/ScEppE4ru7T0Q
FiDO+ZvUFBGVANne/YzDl15GG5hH/20iaOv5428ILY3FPSPEjvs+ertfUFxGbFXNVARJl9stuh63
YGXkTJvU8Qd+BqB5kWoHyn0fSZgHP0jxEyFhV5AkxxaREgr5gUuj9q0XwM6gqNH6vuDw/TGA6T9x
feN0DifZb+ijXMq99C3xEAlnJeJL8h3S1zFr2+wkb6a/TbeNgP5/n2RWErLnH+ULdcSsd7Lfz7p/
HgMiAI4efB4ogGdymBe3PmSDioaF9D52VI2MLWdce58WXTSoqRjIi4gioi32Ywq1lTydAOQvyas/
SH5+MuW6KF9vfoKCd+rcNi3VBSpF2sF267aArKDE0TbxoD7uBwtfAzvDvOWfSVA3PAGiE/8SaDPc
w+N0U9Y0H5C60/LdX2dBJka7gSN5+UcN7zd8aT1U/hKqfF8qZ3Fiu/rYNbPNtJ2C4++3Im1GMoA8
QUcbFB72D/JSJWVwqcsLcnbmhH1OJ1GDgOyShrK0u+tEg0v3u2n6lNyFZ3XYkd7cp+BCs1OsqFmU
RVgKUqlTyJTmPoteGrPCsrRCXv20SI7m3ZFinjPmjAvV5L48Z4OW0+mh3zEzyIsEMk2VWxUi6yCN
/tTY+z3KkiLCN+NNuoaIqy44KYFPGf7MNdNR4RhtZYci0jVDIlv+VRT1jHQavkZwn3nf0AQ3fyuc
CV1UqWUoX1JzT7v/S9+Me5MVuzq2tC0H9B/0y3+58BnO9uq6MT7TWEGS6T5RjJjqub8B221r051v
i+NytEqeEQK8yU/dQLF4v7aVn3sWJJeelVWeDkzhqxlCBMk2JzGSW31iCbHZtKzWVvcEFk19sLyY
CS0/EsPdZGdcuy2TsFZHuL4Mk+M1jQllKs84Y0O4GSbQRLtN8MALUkZ+isVD5qaDgKreb1fvwok7
ONPsY1Gj9nO7KuWKsVl02PgNBhYtlrLb40U/UZVg83heoBZcoPUKqXKxc/7WPRI5UarmbPWF2KO4
GheMUiwmlvDz4Axe4l2YuAzmH+qEoNSZ3cjr1/HxODmtBhfqRX7A1glxQXOEqgRE92mL6f5Yx3yL
sEkXdM/wLXvgXToC24dGITiREefrfMcoQTbE3P82t5ZSpz6h2RhGyoaqyyxf7vuZCryPVsPMi90V
2CRbz+2SYTSW4emkAWYsybRF1FSBDi9PFs/KR5kIjxRES7Nvg/UMHibwZuhUNEBkqnNKWGj3IN5/
WrpIm99QTWT3dD+MoffeGy+7cQ+J0JcuWl3fqtTZLs9r5woTJbvqqNMc8lgwDFsYAHqgxP5Fk4JW
97T/IT2b3RUygJ8PQVrxNmRNueJ27c4mZOFUk7sQ8Tu3mLa2GELMret0hR8dbdOFuOud/zQD9BdP
bHmlKkjQJHvgF5GjGu87fmYiUMJQiYLJA+KsLjrXNvKXylwRy/LsY8FBvQhP6ChiZA3T579OcbfB
L2OFwtVqqvjo4bhvav/emsNy2HWtMRCoo/mjX8nmZcv40+n3EB/xpdFe8y4z6TYH5F0wdIgxVq2i
FSxdyby3GKn87FA/3z6ijqxefxikHAZAlpzGXo4f8aAYFrp5T7rI9F75TMBMPEAXFkm94WQ87k1i
W3lckq7/dgiMESJNeexoLUuy2iExopWFKDK8N2QRoXoCYLHExe/FDOaMCZgFCWQy6wDNtbfMWu11
+IvKlpR7/XwNtYlpi+wta7jTDUak7DQvhGTVK+HDmoDtW6JyKNj8ubzuNXpIpUlLDHhoJkK4Jc48
HOIzdjDDTg/lzmJBQDZ6Ca+K2ookbxBaRJ+k8YcY6c21iBfUXP3JkmkbkP2dw8wjCdgT/1wDnjGK
ieIGIrnRqaQgaAfNeKnsmfGMKEw20RNHKIrD3BfR4TXN2IU/uJLzCCgQAUSCPtQBtJlvts7PODoF
MnFBPJbw3mpxCP56GJhQk6bSE2wbFRfB10cmXIT5+0aVIKCiv/GIh+snl17G/SdTCF514OnnuRbK
eoIZ0cYcKMvBZiUaYySuzpwxHfKNgEMaV0fftLFzBL9edMXJOcb7/IUvNmcBtIHCkfpnFWRNhF70
ua3FU9wfzipsrWB2uSoTtiUbd1oZyJrdnUr0xjAaVqthPVS0BAa+dL5Zhu+VMO5nSPM63MA8p1s8
q6D+Ht4yTHjGF7j3tx5V86Jo+B5Y5ZXqlOfI3wUJDgBxYz2o8UApe7nDJlPWkQGl2Ket3CQVsH6n
nFrm0+ytLcOhaO42xqmtrxWvf3wvMpNjrPZS2z0p8LqoHZPBaMp7dQihQvVyvYpLnIrkmxdAGgGx
sy85DhDNpvcD5olMUXKCNUQ0m5j6M9bC6igtFqJmfLHHgMAl9FUdd51Tam1ADx3U+/c4HtYJtqAx
uybtDOmnp9/4K65h94HhanvpEV3hV8HAPNMnzrMYiqSWjTdDr51OwMRHig6Syqmx+Jvq/xtdhrdn
ejbCS5z1nesIDqFuth+TUYfD7WEZHhgPS7XnPR5Ap1I3jlQM27J/fKUSF2GzCKvb48FZQ0pXC1vJ
z88KXJKCXt0j1oWASSqIpgyV0VrGORFoIExsnZVkDXRx855qCrvO/xObUtRCVowXtE/PPo1pVdVe
fIGJkUbULTbja1uXl10v4S2cv855Damb1784XHmAXrrtULdZUXZrYHeGAc3j0U/LFYTeGS3OCpyg
rnji3REmcYXymcswHKgFrMum82mtrsOmhNsuXVFDePHDfiKMo/l9hefEBGAA0wzpNCRNyPqsIThE
MMWFOOAjaN3dM46r+kKuA1zn9YOnOzrnpHR4QNCaf9foCgEyH32OrSns080M4pRdCaiJ7nswMblr
UIGp3FjYzVdsHTQAqe949HdJ603bT9z9VnKpUdpJWlSkIRKGsUPJA+49w1+6ZDvQuWEV+peAvYVQ
yl5kBOtfHEkt9U4XrGOfB41ebiJfw7nyLzTAQTXFRwl4lI4UX1mRtC40LrO6A5alEVCVjL6OscXC
RYRWB9Wic+AxX/dz2YNt2r4X7qqvl7yJnIJ/kj6Q9AFvcr8w5Ro0LnHXdjSUEHO0Q1FqSIRPcpiS
+XC1/5o38pIK8ohiuAfp8MjZfnpaNxAAom8R3Wg+kCdd2hs1t+yh/Qpn2HfZh/pGZah0Ie/xMRLf
cqkxdNvdraJULKQ3NZ9JBRE0NZ8Ov1sIxp70Y5Bt/9ClBBSPR8zrOZicJQbHdXEBWUxLlD5lig+d
v4be9Z5EoE6CcXxtFLZUOtiJXQ6Af2aQQuAvy5iulbsGTqKgKoB39Tr1csRrzapMnrf8gGcZp7CL
F2uW5Gpe0E8cHfRvbIeMMimF4E9+SQDT3p79xzdhpbthZNnkIxfnRJUIJQRop9J2XpzYE9wAmqhg
HRKnRcCHhtCmXELDeHjkGDmiBX294gVgw29j2KQt6zEmqCwFVpErUCg8waHWbto2aouLX/ey/2ak
JDFsJTfftGNcD2r1O5b88HllKlnc8Bz5SuWuKgHpKY+t4hbG20IZFW5P2nCej4Wi0n9MRl+zL6IZ
iz9MXVeRbiu82jTWSPRqF4dyqr4stWZl+0h4AtSTFQkfs8z4pG7BPawWxU00EJdj0a8Jpc7MPzL2
9iTDeFqsOVcqIUoXwnZrF19z9GnWFbKKGnguoTf9AV9KVSTwPR771uBA9J1ct4TNXryxp8ZRG+Ty
cbxJzP+iIBbB87Yiwp6cbf6O+0aZrr8my4zQCwoCkYl68X3gO6BdqsG7x21kiDxQiAolLYTGDxh0
yM5TikEFaInAaPnsTIxks37YoEzoipy+FqGknT17V9Rvjl93WoP9BmelNFdfR3ceyMzRbP26gFOL
JXLc2pcbXcpLRhdRbyx4fEi89VXKw7Ku4tp/I0UuvJsaW8nL8KuFa0tccY0aXLc1R2rian6QsuMs
X7v8agcWGDvQ4IJ1URWIBGnjDL++3FPU76bf99Xq78F7sh8wQj03yssA1+h8V4BFrIBrwAj8b4ax
GbidckJ3SeVFdLe5y//6yp/YfFbuImiwkwyjmncBmNPjoHSPEURV6TYsaOey0m3noA9eLWJa3LZI
2VBOiZON3XquhuouX0Lz1e4IjvXCz77Yjn4Uhh+z+DrTVyQmB2thHCtFB5KwkdJhRxVZTHw+YpdW
G+aaUqqNFLZuFYcHvENPsPFFQuQFUA8RspJ/zFEcj7OK2FSlAFLlMX/e7SKtNBuNxgxu457Cr3W4
uzVdD9xyNnXxojC1QxOUNJgg11M2TM1avlJnZGSCTRRk7uNmJaYTXzeE1Skwbt+SXTWpMLVGPf61
QRXoGmj9vWtKXuTIXFedfhDzl5SRVABfOnXKbmdMQ7yWd+VhiLuRYD6URJ7aeC9TCCWqW+GDfqVB
b8HgJWhTrT6U6wHDSIbbCvXT5ZviBrfOZs6SZMSu2+H3BojOFljN6WWTYmeaNXdTH3bR4ajIKBLb
CBKZKIOk70JhVajeIcALMG64eViULWsh7vwtzAzkn5zatS0c62GVflraSzxm3NK6TPdqC1OVg1UE
4ZlkPB+SH0dD3fv/qsSYccaNoR1/SiEABsGYAsFjGXx4UdXViD0HcvwZ6FW31vSaqW3TUnOcEQPM
lE5t0VsQmH6DYMYPHpacmWTEfb0zbcc7Fylg+Wo+EmFN+H20U66TAX8lSweOk8P6RWKAHWuxx6ju
FkhhvjbXw2yxI/VODHHOJ6KGlmT1WKJCW6xZ1ig7mA3Jq3WPy6pbldtf3Bn2w7d00wBYf8Fr7M8M
qdQ2DiTPikjQlQxeXXYHpa/+6Ib+OgY6pU2jxIGIHGPvOla+10K5AeZlb4OrDuz9Xbg6M+uvWFW8
m/C8KXZA3M8Djp6EmgV0JLdivXLQNGbCWUuh9KNmU9tTmYbRqCtlFDFi2bbKGU1lC+6F1yco2kRH
gQqyadK4EoBJy98W3lBlgzPU+dGQI+Qxv4j+zC1MMIkuFn00hAjLmJsYvDyVscjYP+lALx5S9cPl
IFGzxNu2ldahSNwdLkUAt8kis+MwDqQPmBLv14X3329p4z/DsemFKjV8juekV7/Os499820AXwv5
h5cXDzeItvMMZkySHGRYJEUTCIVySZfpRgUaL/rrVykghlEL4r1IGph6qM3Ol0pIw10jP5nFuIFX
9o33Sesbb7c+QK6BByyhx5o5pzgnlYHZpTvHmuJzfrf4p2dVtPAmDgTc6gCtNyToY0GJAbQ7VV90
LcKxxhGjkzMdGVwESRH5+BG8zc6giAJ1VDtfzWNbEwOV+cur6chCM7i8kqXMp7Wldnv8T7ekSHZO
mxPX231P5ONC60g+PaKawTy7EzCVsQf2BkPIU30QA2bK99mVDYwQENKT37DFa+Ia0szc4Mp15lIP
EuZiCJHgUJALkHez0ClZVmnP+2Om9+2cYsLOhHVwJLM3FZ0swfYnt6vIIJqxgxbMxP7uDxDrFwB4
M3ia1PLhr/suTgOCAFUGp9FLkx6PVMB9nvc3R+xhgJ7+MKohQj6MjYDuznKqtFWzRHBAbRM9cIhg
/JSLRHUmNtOkb9mEWZR2K+ZS3nWcQ2LUj+xzY1t7+0FOmneF/3KdQxHS9Bic4OKdSn9enIhQfI7X
U5N/3snLCu3vLXB8F3yuEqsN23agk27/oYn5SbZJwCuNtPFpbKuWj3Y9OVpxSHQCOibx0EEcFU5e
q1ERYflWG4rbfQnqmMlWAbpVFNxXqoxJHvayH0Jv8gmXmHky4HFHQWDqSmzjZaaqXcVLd8cusxEe
ec9ZDfEnUptHm0i2m5/1KXVnqDFt4blZU4WQ0PMWQEDQk+ffVloIdjRpu8wHAgCIDhW/s128EQV1
ESA+6JOa6CR0SBvX+RGFFc8c+stP0AE+IJuTM7cfVAF+AhfMD3yGkOQ9Wb2KPb8bGP8AzR5FtXRb
y5+jK+8hifaRo5Wh1pP+tDcFArm1lfW8wodFGmlP2yHtPpg3jeu9HwHBEbVTtoMOyClfxk1Cj8U6
ZmnxyYq2I8lIxYod/AEMAIzfEdk66rs3hWk5A3itKvcIidP7HBPky5fjNtZTgcCnxWq+CCQQ+dpc
azy5+ooIWwLET2qmkLMXAdu45kb7BRqspT8naNW9eUfLUaZ3s3F99dgxHdLJ3HgcExvrRRpS+phc
qVT53Q/dJipbrnyIGkd1zxuRax2zQqHjIB98Y/PD2t36nUVGZ2rZOHGvfoUqGbSvnkhgIoy0k2gC
lZzHzcV51w08KGHSlLBewdpgtt0xvuDGLhVJx3oVv3fTIGZvhFt7QzkTxE0loVPdvNKqJ5YOj6su
ZZgpNy/1ArQLFGRZwMBrI2jrH4+lbz9gS+JGTssayMd1JPN+lyPEmykRHw71Dbv401u8b5PgMcbq
nF8ROGHYLTegROxBj7TxxnMgO4SPVuoHOYVVH9dGTHLKBWG9b/JgeH0fzjjokFLACBLJbza2UuXh
LG1nb0NnTGUrN6ssxS5/7VwQob1kukkAgH6VrloF4IYeQJynSlGANkQZvNkczv/b4zycEO1y6P2l
P7tdQnO+m10Yy2MU6vJt0vbDJKlzdpVM9X5XrhvX2oe6lLJ/EyFiZjNwjmDHOdAeb0xrD/IUmSfh
f74z2PAtDnMk8n5ZvNKQ7LkDd9QapV2hArZFKsL52YucTwcu7LJBu+P41mmzV491bW+JWR9PNOlF
0JsK/4c70ATNF0CFMP1Hr17rSQenOfD2FQa9KTlYUg9ihpGvDUS1Arb7G4co2+YSTACI70YrfCwT
dyY15F9iKGCjMAjHch7d5NwOqybO6iLheN/ftybuvCcEKX7/GBeidJyp+uE/7ITHNWrQRF0eROg4
6oW9YOSS1Fr7KlcjLVB+eWQTTeMsmrE+PA3+zx8KA11c6uXVfdFqQSpZPAV6Tg1gKZUG39flfEjc
vXsLqLL02LCpXuyyB1TL0lbuGvfFv4Ztl7ZT3XjQQ+bLqyy6olZ19jyAK96APLa1NeA4jFgTHQ8l
zzTVcjVBX88T1NGjhkeOG3uc1GYMCPXvTxTma3BwwbaQAm9saDw6JtJWWRf6liQaq6wWVn3PT9IS
GlgZ5x/VNKHn0k7XVsCBSl2tKZ9wZNbJvaDORv0f+s/bc/MpYvFA2HpOeTOpwzW47roq+jq/Fzpn
8tKG6iLds1jf2zRcBQkZKA2pd1/B/1/AXRGU11+bEhCirMymScg6fS9Zf5q7E7zs0KNdXd0DtOTq
5RLDAKm3QzaiJzOyZV87yNtwyvg9tEUO+iMeHAcVufIcdz4StPJ6M0VkMB/FT43l6wzNtNKvOg71
DJZOlzbGGtCMQfnNE7cwApx0ggOrjcEKZPd/iZHznF6Ym0PqCgqKk8pT2Y30Cu6Gw82KArskXVnS
BioqqnldKcAKU/+juhN1ggbf0fnxsX+1+8wWzn2qvy8Ljmea6yApXRYtzSF67QBXfBXafBXXDWY6
kFWLMb+Qr+NYKyB0inxa9obduXA3Xubw6em4zPDNGtT09qT3V3DLKq9eZHMQjrdCHIpMDCcrI13s
HdiY+IUkZg0le+ttul2FRuANT84G8BUGq8APEKzYC1fNxmD1VNGkJzive71GeAUZ7r6BlRRaNnah
H6BW3pdby4e/66/goccJWJyKgCcUbqWUwqqu3tB/VwG4yIk/+0C40m8gkgXEve/Pcr69oIeC4fKp
T+ORnio3piGRcb7jSVAxRbLhYVAiYZPV/zqILqot3Bb/cuUs8qQYhmh9CaKLQzowqqANY9itV4UV
jmanK6OEdtSeZ1ZrUMXou8PEVSVTtxoZh0SDxawZmonmPf32K1ZoQMnwsFF3kybUyn4Q8mmFJgS2
c1NKf9l0F0ng02cnQJKjf2JMtFymWixVRlyu8Ag+vdS2/JO/R4c61eXrqL0GL3uMU56rk9bAN2gV
p3eRRhGZ6Gg3m2a7KX/DfdqXxvqzNycg/xxF6E6ABd15K9p/GebQId6P1ksX1k5otPHO5hXhKs95
4KRd9H7L0KfS/+Ena9a8x4ByO6hJuAMFT/1mPccPASZCKZlHA9rOg88hfNScTu7jEt8aPsY83Ytb
16YbX6uYk9kbTI0JuM7NeP/h4Ujkp7T1kLlGU77Kfr+TB4VOTZX4jUDSRD9InGhSFs+JaIb7NqEX
gWl+v0hgRDIBm2NLUSri02kxj9GTPI5ARzisf6xbYZY111EGqRn3Mj449xyxomTsEEoofOf8H3IB
ctVlkbTkM6Q2MHvnUIhJkqhLSK3BWgvW0zt7Jr/O7yxZWoFHxZz43Nn4yk8vEow7XMAEsLWDPQTA
GE6bDIlbMXf3Tffv38atG+BRziDiQBIbvt1zEBGrZBAkl2HSRwmtfoGgSc3yKZcaICCByyZJrXVr
yMRZPxc4IAYvib+6H2ZRxIv5OVs9G96uUVELTqubFiDIVQc9LPpojXePuK+vA5ZnrOegH3RV3nz4
hQBxBua9foDjTa529XI1dMDFsW6b1pXgVze8nPutIkPg7YIDhKp1ITSycpe/Dw7lxcr6jww6FMfb
rwLbTA1K17427ElalCpgRXTY63hR203Ipe+LFKsfVEWd/CsrpOuCejwQa/P7iaxegKbr2m97Ot4M
oiPynnXRwY8z2mL3TGTUQyqa0zMdhnrfAzwD+KaAOoyqSOiAD0QroJJP82fzAVLXdHrcxEELkD4Z
RxaY4aaflBHNL8P0W9TyOs4y1zBzZb4FHWse4MSLYfCm5tGLmg4gE94hmHEGeGre+rxFncSBydZF
U5+djr8vJ4nKTsOV31XFL+m+oT57C+1Sn5FwUwQHUBZGSyToR2si1GAvuE9dPo4L1D2lZiobl3Hd
jbI2FZf1fsIXe3y+vveT+5MUcs5yZ4Yc4giit9efLTmXYvW1A96pEH5a3tIy1kq26cZkN3TkRbUP
rOKOAhugZp1dXbXsfx0oihm0mapUfsD7u2HtdFiWZSQZhm097b6Cic1m34KasYakKkPZ+vGzf7dK
OvXazR/QA99GJjh84GR6eooqnRWlwV1nkSpwNetm35r7UQDdtwm2xiF/BH0ruD3p0ZoJU43kbmbI
DbtvIZtxPxfJQ+Slge/y23IAimxJLRxkZAc1s2kifAOEYqqnIzDZKfBhGVeEBDtgMqupbtECVYd5
0liitRzlQBhN4MxnHQGX0xH2AY561apehrPYQ7VSr2QrEm2b+bwHIaTbk68Lth0V5AXxmcpE0lpA
zvmbmbmFHp/K1NtmPdlNEf0aGm+DsxTWxLv23Y0a8oAJVzFuMpsU19F6Mad8XbXzbN2pRyaU5Fbm
nlIcQOmrsmNUgbMYWGh99gc8lLslfczCJBu36MXVuzjymJI0PD7h1ZVGynQVRy9iIyRvrT3E/TV4
IA6s2vU5E3Kpl2uIbYN76iuhsIRhLiMmn5foHJLqHJG7kyaWMumn3KrccQLQ26BiwJYLubx51AvK
sUA4b6TNFntFquHq+hY4ZlvxDkF+8egim6XVIQpluN2XITYdbm8FhzSnrSOPAIIowbraC30F6+Tk
VlTSVIe4GBE+rgtJJrXgnnHwQyRgyxxMCEO7xDS+dgQQvrUsPGhdfF+JUM7FLye7qyoPURFQf4/i
GEx4qPbVMjqQImamyH/vQ6wqOuDXgYjfBleZbCjWWjp1T72PTko6nb+Ev7aw2k4JbcjC7YfLpwTY
PaT/FuACi/naxEFYnSKZPuICsC8o8U0nUZhycsu3VOwF/42CUyQ0nkV1sDLAQk7WglFSZNwMH2pW
Ys6RZBh2yCZ7DMh42Mi7KpcmbjsprfN1Ex4sWGM49LV3UubZAYhu9mrJJgqasZWPT9TO5/nus8Zd
J0FuEqPpeUXw77osbeTDKQmfZpNBnqpAciF5+YCqpLnHsO8CA2Aju5uBwbupAoTrKBomjZ9AfDVo
d+jO2BE91x3kV9M5rYaP9JESJKl5fRhZl6OB+JybijdCnlnw8SO+5MuQ+XY488acAcwJHEm552ph
FONjdE3cW+GrPXMojeL+DLNWlQOJ2M71OqbRcfZQJHBNfR5UWTPgKNoZfEU0PUFULFtMjVCLHMqo
3TKgL+oJ6nfZ8h9FgypfvpksAkBXxv4IVwdxdh6teQ45rFVM02sPZdxfLgc+u1aaGGASYN0Xqtl+
2U+36rme4MzTIKdSvys4DHkownAM2hzuxVWZtEn25CHtE6NabjFnuxdove8FnG73yQB/TCV04lDb
gx61zmSoRrrev7Dj2ZdQLa3PGFbPG++tg7YBIAs+99KRyUrTXKInj3JVq09Fs28NKd67Z/LFpyZ1
beq3IfVu3Z+2x147wUTE2HN65tUlidHeUL8/eMKnCLJG0PIn6lB2A6izwFWvp6O5vxc/wuPg4mRx
khPfXtjs/5Q9ExDbRY5dQb4ELJ89cJcEkejpBamO3bCIAaN3je7x41CO1yamGkR2sxf59a88AVPQ
2maO0NDnuPzEQQ6DLM8Rbm4ebAvuyaN2V5Vjsq/y9zqKdqNbjYxETzx0lny6QJoousVcMCEys66H
nH8RSh86wzOOh5PLdz65q9qQ5plveCJrMlRvfVBTCHZaM5r5hI+kop1YftP2QUOItNqcWnMgUuSn
XSFSNo5BO+yImNigPkVF4Sxhy+tpcjwc5CzdujvsRWo7dzXt6fFK+laWnXymHxf44tL9+Fz7VpPs
xchWLM/WjlVX81Xkmisnli0cJW7XI4N5Nf09iRm1ekZZY3HAkEJI2C3OYqwp4RtayXk+43kcEcGF
EBPwrf/9i0hQIs/XZ4iLfpjopEZ2D11VXG8whnjwbAF3UQoAQTW9E6lA+6bmPJIlH2wHVQ2FuiGq
URXwK/5koP+qbpvYhkAD0dSe6qEXG7DhlYMba0SDhfUb+3GzARp75JGO65G4Gvc/Jf1ciC8xzrOY
/itfNpRg8eSWsIQ744OvjKeZZjUMcQt1o5rzgKfdZ+uKIXHmkTtOpWV3h0M1HkPY9bgp3vJt6i5v
Yt6jixWfVdMv9ZdcnkFhbjoz2LToiIoGVz0ub+o4YtLiGq/ykOybtTrNHCWNM3VxXJR4Rm2OlhJO
gjN2bSbjD5rJMUKVkMKF1AmTssVBegkkT3A3G2Z0ZHCZpbQ+b0Mc1LQoUmkXm7479cvmFoN5N/sf
Yf+yc1Q52ncEZdfhHMOmA/UMnqYmTbRA8rVjKI4uPfWJGSVxgODIPXoeXcKk2/OBk+oWHx/kBlhq
kPDy583zlCFs1fonJKxu3/6+P4OnlQgVf0DiI1WsQyiwwhkoHNnW8okjoDhxcqz5xBavTHpRvANk
CfayPfehIqCQS8qm8D2n/aMbDI1K5FkLZCSxtn7gDNhctg1X/3HGXNc21HTL0qOtxUbC2cq9VxAB
CeJ87An4vpK36iuKWRTKPYakkwT1PuXYP79Nq3++oB3F3gf+CenPbOIszfiojXV8OIQD69BZ81bE
7zT4XqxD3jTFX4EwjYwO5cYzdrfO1emY0bvz3fYIttT9RQSdmgTqHKZRbZORkryJyQEatO5zeJjt
LpTQgoIex1JvHcpeg745+e1lCq+mx9d7Sm1bXJ1e1z6V6pTN9n/tFedOopUKbBOo383wQ/mhdM0m
MGjnMUXrwH50+JeEgWV9iPyiF1kXPs4CgVWPrwLtr87gKcF/DAsNWhcLK8fX4Dz5gqX5i8irwrTq
pvHlDBCJiUcRQJU5ATjZfEsOV16WvipFmedHPemTq5JhbTrxT8t7QZ0uQmp7b5rtauq4xpBqd0E2
9kbrMSWRfcNNHTb8BpTsH3d/RWC9fSlbQGBDZmkWlEl2SQY03JWsbI5mbE6OrkowRWA9KLxiYwYt
GfcC/LZt+HcNAlrCv85ZYcpFMRXkmyQlEYWfY3Q7qYacyBtEm5q1a8qP72ZrylHEeIrxZffFiEwt
SwAbb4qVtU6A96/tYmn1h1a7v1uy4DzyN9rRhkpjeOloVg1LEHNRCWrW5iLGRcmECE/M4BILdGJp
NMwaJIUTZOQKfXzZhwAD51dVm3E9hZffYpQ/M5f4wEIhmK5ROyHLSLDcjPMPWppakHcD80GnTZKc
qYQSKFQEkwlbIx6HFrGEKkDgFxJO+/NJmuLu+TCn2OBohJ0WRtcINTboBxRgwFR3bINkqH7X14JQ
FZGdB1DUT7rQMHdidiDMEtrT0A8vDWniq7Civ2Hazurqf+m2L04VPZgVfmpdWKfArB61NVlwH/oM
kgFd15l9l5SRFx6SAh/aH0ilBj52dz54/Edh3UttaATkC/FksNp2Fohv+JMJoKdzcuh+TBg1QwTb
Ly0s+4V9S8seNN7wjiJlaJJKkzqldCV42SnZubY8tET886uBy+BBRiX4mcR9iRF2ezvbp/Ag9Px8
/VTZpcP1hGo7k8hM+ye4b4oeK1Zckj5vXo0XpKtISnc7gZXj5IbYMKKlQoGZBsgFk6CWqG3z4Bj8
joRxDxfLLpm68eHbXWCC9R1PV/N847w8B+HNELNUtD6KN24pguUVOeuZSNbdvA7NJL1A0DOv7o1z
0Krfia7x3zKwtcFf4NwODKfvTYcpApDju3IZ7Ptbpz8e7JFEZJrd5tKLHPJq1ddYiN9I6y2B0yoV
RIx/Z3FHGMlF5XTOb6M2pOH8HgPFInTRXIWiIPbLJh/p4xvaLu0aYkOxqV+aogCEsBB7skchrQ4o
7fsrs+fXYXgYzU7iznCROU98SXua1VvA8k9itdD5JA+ykFNhWk42+tdHxkSYYZbRxdmU+RBdwSBR
QT4wc204xz+mSuMWn16zyp/W9cpgpWWV42i7Ub51WiBiOHCLSrbD2h+4iin223txvyJ8qOwTYClT
Ats74haAGBjcsk8ls7eC+fZ76lbMvKJrNjYziktP5jhH+9UG137V3/QFMSdhjahABdxxurFiHQYi
/XafcZhCiRGMxqrGAGfrl0HjJqVwULqKJck5+mD/MjUUiGXsevxuWYC7SQJxT1dNPSBPp0L7yokz
LwWz5S1ikAAjhCT7EiZIAoWSMEeJbNPqPRP+gj1RZ1fy0aUT0SXWYTRWI1bqzZbtLfLoHtJlOHYf
3RPq+SRp4cArmBwPSd8uJLV9Q/KBZzJ0zk4jiKEt1pVyGhnhPx1KrnPeTxwoMLybqdJKAOM1QOvW
xJ2uZm+HiKdNr1I9emkmRwmO4i6NrVtjxbWf+qpd8W6WeqJdRKjn6idB8jh2WtxOSq2krvs53FfO
AyaGCVC2kpnjfe+0vXkd7iJLuLmPL8+og26nuV0cd+998PhuXJWu84HaWzLBHMl8SrWmxbwUJcdI
L6cPIzkEobFcSrgl6JuL/YrScAwNXzfmL18o+pYqQlO4uttLLz4WabVd1WpynfX77FBsHJXquVXI
vje9dbJqk3Agur6mIhVjQi8ozB3oVQGWIdnXxd8rqHDnr1smM8AV9kFrt1Xxf04HE5hvrkKoxNUo
UL01JpkRv6tBAkGLIKxd3nPrwl9sA68o0k8oreZkFrJLLMf8BiKUiu9AwBLyOAf+H5Fmxo4M3YKX
EDx0074TKkzvBEIE1Lnt5a+YMW0yokqjcoXM/X39KZmYuV4MFmrmB1QjxlYIE75SZFoX0h0WA8bq
WRY0lSjui5c+P0qc2sox/l1heHmV+vI4V7pGRuXx+vZD8EnAy5jAFzEbbCRAAfkVbAqE6ipwcFMv
n4g81wmPHj+v+k47trCQ9TW7r229wUgNMYqKumfEwUaxmlfNDeQ8qdHKWmhonlyZgD0s117LbgJ/
2AKqhelhIk3DkXM+FPfx/gV131rwJXv7X3AmtJsWstRuiN7Ggme6N6wpldhgno+GshBUdvgzFZCX
OptwIDQOsNBH0ZCFwd+1CT63/nZu6dpbaM6lP19dLxJgjyhWoxCYoLUHGMpO4uq3uGn57JanIAj+
PA4RK2jVC1aQN+YGQmqHfM+Pbk+UpbQB2TDxbB+LANZlny7MAoJT/7dDSLMPQ70ID+1ASM+YKXoX
1mpoSzIT/1InqP0wWh+9t6Z0cxVT0XYaawwPwwHbiHx8sCGPkq6YpMB+Cpbn8lejshijM5OE4zRx
q4e549yXnl89kFj2d5xBg7tFoOVX/WLhieBZjyBIz+jcPSEo0D6vwkGUIQyIoExy4z/0+ELIA4mc
zF9VJcmign71ml7Fg8vswOCiZBhC3ROY4lMB1UoGXBqSJM+MjOWi/QNHA1ZXCxJWH3iVAUQ35VR3
ui1Iwh764pUj8bh0U7WtgCPA0cHshDAfQq2sDmJUtUJNODwE39SkYvVDXuKJN4605JQLKKMae1nj
vHjpB18xmH0dAH47fjI9XJTgmnVzTpXeYkSPJrP8ggHAeMO+T4W6n04+l3zdlWAYIRFme2CvdMo1
WUHA1gWmQZ7Rv++wMzNLPUYEMXUfV1ZAv4wp2n0iEZgF/ie+85OdHqfcDajtGyoWiLAPcUB1X0Ym
BHLMiEjgShrXSycnWD8JBefMFhwPsGlaG+LVXtr0M4amR8iw7VXdKpPBAL+qedNXReqsiSvkNW05
lIT3485JnThV9CgTheJPE0i5HIVcdjzk/J25A78d89/bUTwrRAB2u63ErWn8R0fBbgu/AEd1e3nq
BG8jEiqpS7v9m6XjIS7ux6cOZ67s0Avq9ZYivZwB1qPsZAajQaYhTquZj1gV8ZZjxBvmWL+3Xp7Q
JbnZR2gLggz5765jwjr0SIOK2ESDFHMHLYWApo56ChaoU4nx357BVgijRSCJ9gHS79r2e0jZzVSO
6NDu++xKXP9HmlePpKPpGr8uldc2eVBm2Xwc3FoTEY86TqRga8J9FEvLEg298jRYt618oJIfDz90
MZZPUt87qlMiANUep+qg8CxcDY94DBYpm0zv1NbXF2FG8yLdA6m8/bvmFn9EwmrEllDh1squnWr+
ZI5YFIhnMOvqjbbUl910wlBXNKwQjvKERK1fupBtoshMDF5MEI0hyVMN9CxWkaYPuN/+d2Gq32AQ
Zc4Jdi7zk+o4clbnFryoHisik12A28TgiPYBrrNwji/Z7Eg43fZZQixBP4ET5vd3O1TVbSw1nAYH
mq+KH7S3ekgtCq90X3/9CPdyjnREOH9UseqOlVmUcQasIZyn6cQn7Wat/0URn4Tk78oPihOKvd2V
taUefQiaKcmYhfxkMlRlRQwTGrnrmLWLXawq4V3juR6mwbp5Te0As6RmPHYTskIrytq1JP9u9f7e
Paot+RMUMMo5hUjDPlPhcLy2xMpComiMqf93e7K529213piPUFIyAJyvaDWnse3ZuYoTzy4dHiXa
nkbWs9DJmp591VH3E1zny/E38Y/3eOfiQHiXyD1a8D5UedcQJ876BzISLYhf77kSan2AqaHgtAWz
yZMQdQOBLgjjEwja9zJpBrxI1BWRg86ckN2kKdbg97f8JNhVUq8dvHKT/7NzXWw2XLttIEXEsVbH
5usLF7pMY1EDQoq6XKsUsU+3RVBmnmgM5EKM/AJtRt7r5rfHyGcjm9Nc2mOta+aMuz6VPC/l1ndC
55TmL44WybEEEywJVIxfrpIBH22TQixv9vDQu5VnOj36/p84AaD3aGf72KlTX2UGf8WqWOcovGF8
o32Ln6+OadL0awFy5JIcKylsyz9b6OMd1dlJbIMh6m9NDByFujxoIwIVfi6tROsNurMdXM+E6ULZ
OuPfCAJPxy3PB05U30eByY0I22mU+mGrXlOP9fa/gCzCFcaJk5W+CFt2g2UXcUR4fR4w6Mn0SSEy
krzheesXh40QQpnzUxFZJkQdVvnrGCtBGXocGhoaONJSjWEKMfYAbtKJucWz9ngcTWomnAGpdckg
wzlSqrCVfX8JISFqWo96+gpOB/wYehaAFvSD4RoplbYtpjme08HawcrvKk+CRPgdIVO6YdEOhRQq
Kl1ceSwo/S1kFz4svgE1Zf0qpfvOv9VgDe5j9S53wH4x0krxRhrJWFeDt7KkJ2AGTzIwUm8JAmJU
TTa1gjUY8iA1S0F/z02GKOK6yMRQ52V1YZqZxAglCuh8pLUtBdSn2WbL3CTxQqEjPSmRA9xUTg16
C0W9OvSYtIY9v4wqLvblY4mQ2VDzER5KvNSGyKqjkzszD+WFYISi8+OxKVFCkbt7g/oOjOtdASke
wJD2VkUYWv2IGMPUOSn4nP9XqZAXat8IQma0SSFE2Wo22o5H0B6jWvOyKTFXGGEXKV1aVcFoLYyK
tWm61T3Xm11gJQvJ6tskRndcgP7tyVh3oPAlNR50il2jtl4F8j7i7dD5LugMLt9YABjoyqOdsmLx
CUJwBgB3yPD+RtceR27P8nnOpq4bA2QAOzQJr9zNjCLUQbnTdGwgiei8PKba6wj03rhsjsnGPKHa
efyS3NIqLAd3+c0XnRVQcfN9SqJDs25sARxx594LRTIkjIZLBmD48Apa18woZgxHaiT317EqcIQZ
WL/FZIxS+BKHUCPRDDH66ee57BRTb7W4Bux32ubr9i6aw+aMXN5sV+yemhMqkdon6KiPVbgkh6bx
FTCi7GP1Sntl8hBnD1UxBeuLDUP0JaCLRTQPo1WsJYUO3ALp/AE62fIy0TTZLvmIOD3OomYxUhsq
G/7D1OED7OAazHA6cO4qmqTFGQSa8yt8SgSTpHA018ZaE1nsglposylbZ8n+s+KsIbm4rWHIjw1T
O626ouOTA+SrpLiNr1J+JmBOZ3mwaMkhHTEgOz4DPZknmtvxqB91czS0Vr7ZhEVAKE96fKNFLo9A
nH0n9kf7/PQRJsEmanf7G53ZsVnCR/prQMMEsYggEBNw+O/DCSePqAzYgBwVSFtCvVA1UF8Jgv63
H0XJfUFofF4wYwHT7qhfWLmGFzpdddyXaGSuexiQEmMK7xh6xZNMNGtqpN0ZndieSKVc3plKjdHk
zQ5xl4MMPmiJZm+L9cRUlgBMoyWOZSPJn96pNecVq7xmD+SM1VCjO7G/gtiuG7PiLMtjqrgyqPgi
sI8cRdRRg7hcYdmyMlAEbNlLsfmiL2zAWe5mtjgUdCt9IgIuol7KIrz74qIIATz4pQxSI5EyfQUQ
7GtIOMaI51zgdB3ZBbm7IvRGi/OYQIkDmNSsF7E76pM/AcpBL6MCbbJaGc+0Wwj7oIgdDTyo2Y1z
aRsYrn/E9eGxhkA+ecLoS05QmHUkkQb1VWQTd0YGBSBLxz4+orkOHZxsLDGmW7omhLgtJg1oFaDA
wbzA1mQ8RBVbSY/FpbI3AHgxI7HR06oqrsHxtLS9V9sZ3PCwUMyTq0AjNX9F5M13ArfMOO2LnGV3
tfMvcduE4Np7C5o9Fa4CBMHmaPGJxDwSoG2ePh5tqzm9ySangAfoCUXhoj494iS2aLkdeD5qOVCY
tPKImVEAy6lSHbJSyCzBOAKH/nn157nWp3jLCgCL2iwQkZ1xLKyaKyTB4W+AYpSn751rL8QUYbZI
/uAiA5zvYx/zUNMPLQro77pOgtY8iBObKsRKhzbi8nOKZkbVN6T7JaM19LHNEhABr3xU7hlfcDRO
8uz8fS2O1YSkewasnPk7WgJGHShQj3QbpqSDGlh7UGGFhiC9jltjraFxR6lclQFyeCp6bluYnNLM
uLaNoOCKqWx89w3IrASgV6FBU84B40PO+Rd0S9ooY26wRoVOSinLdeZma04kV9UbVoTTlIMe4hea
9oPpaOIYbbz7K16iWOKaotdgczXWSw9kyjPaKihRr1O9FXxMbF81IkeHE0kDSe0PGS29wWk3ybVB
cjTHTSh0eDV6vHOBYusurd2nwheFDvxJdjoH8Gyy144vD5oMItj2oET/QWp5ZZ0koLbzycS1wxz+
iQiJnSORIRVcl5ne1fSI9nSimciWmco01aqqZedzE214IXdQfIv+ipfZRI2GmsI67aYGqVxxLf+M
NbtvszauiR4Pz+nGx4Ugx19T/E8U2F1ZhxjWHXYPun5PpUDv4G7kqYOoWPy2j/g8UfG7gNYhoUs+
1WEUw5CyNg15A1gcRAyVA4mMK3s+6FUHv8Up1PXYiXjyKh/BAz3KkQcmMWdrobuIlOxDMZzAEkcy
hkde33hR9XfccSvRz4w+FZYHLcE1ZwGXYeK25CheGW7a6hTauJNUyJWS5d5+Dw3zfDBpTfaehZMZ
sYtyUnJn9mo6q8BPnVqax4KqzHEdacVYVhUy7GivYSKs36PlS34cM+qvujtffiECxd73u9sfaj94
wfg8s4cGexQwaIQKJiKuQVu+Wz3nSXWdr5rRj+EuduymWTVZjgfhifMYgl1OiNsxptMUeRo5/xFK
F1rOAfePOXngVdRouGygFUlGQcv/bKhdT+2TlnCb7fKmomcMugi2+7Hf4M59wAFLYuqf5xgQyGFO
MDVsqNi6mUavL/eoWmSGzeCt0mA3yY+crE57M6ZjsFOtfKsEiORstvm4w9FPuCvUK4FjMdvHGDXX
sRHnxh2RZJxRQpTfF3zVWO6zWty23Uufa6xutL/fK1EFHiYSlsYZ7byaQQkBS/RD03pZx8oOxdJy
GbxdBGLElL5pIDFKDrHEIcvCFnC+s9OqB0woiCLmF7PiM9uj5zosrHHdrbga4bbJb2yZuUFaH/WL
VgFJ2R+Rqb/QfEzW0M1a5YdYnBqsi6A6x6T4vH3vYChaSZKW4yLB50eAJ9whyUIBDroAwhR+IJaK
DUZb+3YXHVvUA75MprKta37bZDXxKgxAFpI0XI5zJtZEmZ6HS+/0+p3yjFvw6IX1+g5eBYmG+Obs
9WtEuCtFZXe63wwFzVBAGyvwHAPiduUoV/khFor/ZNl+khNyr1wCCsL07oPf4na+f3kGwUtoVdVU
PhCCkoIItOsApm1eZ7Uh7uaXBQuPZIzzftXC0G7e9ZOFl/utWl0Sy+b4H3CxZt+iviFvBEghkuhd
qCN9ZhNnQbHRH3tWpWzWItV68b+Zi5xr9F6spwoBQXvr4zcKVmC8pWnYLTAYpUux8k3j+VSvaSUD
6RqZcpggBfcLCovB1BdQpZ0fUxiHyiSI7IDNJqqlzkfFX71LfTXahnAvASXhuYylX6oWs73frlwk
5HGK1cHPz2+ZENkqQUt1GssPj2wtjHr0Wgx+xTvAswIrsvrPftRCigXuIR/Zh1OJ1YHDh/IrgQvY
5OkUqXcnsNG4FCxCPyDK6vIqp2Nsja55wfUVm6hU9A1vEz3YhVMTqdytpoWlHev8/v16mAA+PZ8s
0dVZHAvSaIlHGpRMXPX1DV3L24GH54iPWVPadsfNuGgbse7GoI1fHQAmn5deV1ndFpWACWc31Ya4
a2r9IC1si08CzN8CiIe5E293iNHUkCj9kuYFS4tfZO8Qi8tVrKa1564zzqthKo7vZJiunkKS5sDl
y6/YF0ZM/8qVvHDPkPLX1MRdXY4cYWGbhfF5/aOl8N2+H3UfhSaqv6EWdv8JTo/aAco3L6/k8jWT
ZhzwXMIhawDnFPOQOWOb7CEsMFZSgg44EwQd8uT6jBdvcHkf7JfhD5R/nVp6+RdQarFANkXNpryx
+qKfcS49hqshstWRoXonSTfckUgFCCxZ71UMKrmA259lnAvszL27ibXLgFTKlsKJJY5R6lSDeft2
tcGUXMl/joxLa/gTfqNR4Pr8fHmq20ESeK3Kmw7Ow0mbQHGdHGMcirLcpmVMi7kOtFuEy25LmffA
d9O93VehmvR18vkEHU3GMRkDrc1JLv69RIqVHvQTKiCWlfPtOcg77HKTtksgy7o6UFXSuefYeHUY
dGqDMnQAR6dl51xvVZ5MeZj+TQzcvSNuET2wEyYwy2Le/DIz8UE0VtMWfxu0QeNcs4+ZDI0kYh7V
By3jH8LO/7EYXFb/yz1rvmgJ9nic/+VOpdNHUHNn36qRWIsSX+AYE9kwJt3t68Vn8lrhbR98TRmQ
lOn4X+lOYuRU1t5wXBiRElLDug5DpO105iUrVwZsh6qxgeDNnDN+b+2T4uM24DjrAF52aKhwVesp
8fQ/sY+2iyBXcVBrV0vHP2DOkx7phmHfSU6K2UmX4zEjPmasJq1VFdO2d8IepYEGWL9ujkgKgZSH
WhLg96sSyFWEuhOqwFYYrfAlE/4trYhsb0XFVn5AN39gruN3RLYRHaIX7yRG4sddVcgAMNPvOMnl
VeEHIYBpMQZShgoH2qfz6MIrWVp0g4amkjEhf/Bed0vPoTs/Ivg7ok7+tAfoiV/7vM8ipxY1ur/Q
/YKyYfqoU6uYintmuwHnSedhKdXHPrOHHf+Q5T46EaT2bW5fMnI+pJ7rsN0emkcLDT/h5lDXSsRR
mrOEkrIeXr8xnV5yj52cposv30ODLwK8+5Q8VNAR8hWXMP7/RptBC+Kj59dW7tnA/QzSqAq/TPGK
wXgAUDK/1dxsMsDU5yNWJB7XYyKGmNbNr6+y3irmaiCrRje5TjVSPGVmUiBH1v1tc6/kANSIBUuB
sLKAAnbEoHpHhhx7nMGyQ8PbgLPSyDUHC7FfLzCO6qpRhCj4l1AdQDk84vZnqUQm0K3CwZwvba7G
t1KL0LWTa5vlnVifwQV3QVRROeFRel6CSvMQJ84hszBrrEH/y/rQ0Ro07dLzruzL3DN9AI6dk3K6
gzL2dyAUtvxF3Md4JXSu16Us26k6ix4LY5Foy5G6Rvj+c8G8Nd/WYvb9/kWswJurFOunEWRT3TIe
n+YAMXFZ0JIdKcQsDJS4nGiV3esflzcwNMt5mmlFSBW/6tHgHXhM4FWXrJbImhBsOJrF2ZHHE/eG
GpYUx3ee8x6QfFgci3rglUbuMOu8RsfgO72kMCFcEISflq/O8Q6AGHAntp1OYBsynyPL/YKQRbAS
9fMhykoASBWXzukNrGaJUriPE43h0fo9+TJUBeDfTkdJX1eZXn7haA800vaPeR35H6nH9Lk+Xh61
dKOoZ4OXYDOrpq+h33kN4QuE3rQjBJa5Yqpu0Fc1TUTRp/nAGBBRyTUCkGV2iIS4UAABGF4shWcO
PodE18+hXngsxkGjTcJDVbg+7mArTAEZJfJfsCltpO+iEXF3ZrGyfE8FaTXiaCrxV5vkG5ufKaxU
PoMU1tKLkZrOUO8FXq2v5MxIcJVxpJLEyVpVYpZ3RfcAB4ALDjC+mBHub2cx2CoWutmzpoHFT8Mc
wdWl8N2CO6XKkTitY3PTMDA7sIo1jqa3RIuxo43ZUzhfSo0Ztr9blFLH7nWoZzTrz8Q1jyvKBIUJ
LbFHQTuiVuMG1Ye1TaXd//av9MzM/WOd/SQCoAvh1QTj7Q9KD9TLw9nBW2h4jRrNT0BopxdoqiMu
2K+TK7wrnoegDotZvJ6dyqiOgLk8HAeIo6eXdLdw+NIhusPauJ4IxCancSOwogsorGMN22MnIH12
Wgl3TFl4Y0PNx20lKzuMWtqCQ5JHazMz8wASbewYIaETfY0xRmcDYadg6dqkmOepMUEGLFs15E7C
fpdN+k7HijNhtMD+nblNKglWvxgApSKMD71+JKwf+P0JdRvi1qIZI1rv705LjZdLzDsJKh7Bem/k
OjSv+WkI5Sa8yKQebCb6dxCo0E1OUJBlHPUW8qKWA9I7DRM4PNlTz1MA0LpDLUZ3jfrhOCjjOXIK
zKKaG+BqewCHKj/xcIK8YHWbFXkU4jQRmq+d1ysg15lmIjxMR4yawRC0vmN0RH+u32K4nQkcj6bp
s5klJhIJOQgSTpDG1ETh95xSZwBQro6wGHinlSmUzmUd7TigKf5jgls6yIK7gslX52xTR1KVfP0M
1BGRfBPJ9QvvF7S5u1X0kZGyDg4EWz9RSAkuTqKKo0HYkCDRBbjqvf4zRQgFLIFJrHr7iXNPhtNd
Z+3TuFqLEhhKz9f30LwyiJQi3+MNIsJ8yuxLbj7NoRQWoWVNKo4le9FkfmDyU2hDIqRLrGSqi/qN
neLiPVkip0tbp/M3UPSAWJ1xK4gM8ijTEeG3SqtVjKpgRyEn/bvaDsVORSjMJF4UiDd2aUKQxH3n
1ZOr+La9nx+B3jIg27Mc37ahK4b20T4R/XJ3F9DROydvKmwA1jvsibD/CXHYbjfIjskROCAJ47lw
A29wNzq+Hw1OZI5b0filahYBqW/Aa37IWau5oMRapQ3on537oa3YkXdAmZgce2m8embVz53v3mun
DjDDdHIa5nlx86wj9CGXrIEWWR3WF+FalXXXEPnJENZX4wBEaDacaD+myk98Oh5zTXgaFv4/frS8
LD/n78ykuwzBlIqSiTpLX2IMcRFs0sBkwTVJVmEsd36C5L0Cq9mjbIMhknVWOuYPs4GSdiRhKR+H
59XtNMzbhjVV2lGJOiGw5Wj+ynBnAGf0YK2fmZyTyrUmefc0KtsUtWtcWh8a1gKhJsYzPUQJ+9ZF
LeEkOitDQMbEHjP+NrW9JvqjngIlDQhdT83QtU56k0LaMx9Q0QNUeH8t9Ddm6vgReec0nVDE7O9e
nFq4M48X3kV9Bz/ysq8tC6dckHwOvl3hFK0eAUYN4jDsIMAHWUrFjEtV6MhsDI/X1VeVMj5HaE5D
CeNHbkMDHUbA9UzCwnFqZfuNx97yDCFp2D2q4SSRFNjCcifQFWOrd1S2jBEyq1wjX0rn3E7PgS0m
W6+PxmhaopCT/Emgq66AL61PaN0ROFOS/tF0IFSGvipcsSF8qO7Y6xAgxcHXHMjJyowvvyJvQ9M5
BpLziiFULca4Q2tfb4DRL8/v8kA6WX34/tFiSe3ZBHdf1iYX2dfZ1ACv54UddimCpONlVMeRNOW+
/EogxgHOAJfPdlLVNA5Q9XS0Uin/d2E0CIOD+N7a/HgrPpNpyEMks9XOJZftyVxtCsiQm62LQZX2
reKZU4OK5j/QhHI53dpMIKAUxNsi90oP7YxobVd00jKl8DPk0GIwIEDQo2bAXZmhKpsq9D4OM8VX
W7S0aov/OtLht7mh2Bf3rqdON2nRSxsi1UDDEL3bMWAXvZkyoE9mH8x5wUHkJ8yJTovfy148P4bm
HeAdPOsHoGkMQ2aXu3lVFIUvdM242oKApZY38tS4ba7uFuumIHot3kYJLNYpIVLmBqWy1N7dcSiT
641TFZb1BSAHHGYwFsoTxYvZkAYZLDTlSuG8SJWDbvzmQ8xA2mR+jbk1g9h9KAy+XZoHFclXCyn5
mY1CFl2nUvHlvoIThI7cFKARzqfnXWh+jpBt88IOa11ULGtPYTrbKMTvqPWB0rdE0hfXb4AAvGVA
SXnc7Uzrr2FP45hQCmJtjgYFb+8ntcMuQqtmHL3oypC2BtMUjavD5u7LqSLop5+Ar0AE5omrdAxE
Pd0ON1qg9a/Kz5CcDJGkxJ1kGgRqbp/2nopQbDyi4stRXzoTsaIWApdQKS9v2tlg5xJL+OlE4lce
4EO/Y7fs59q0V1EP0KaqWXA2MPUbn6ifdx+2ZAOFi45AztUAKyfKFP2AJwQdmW/p78Il8vQD+VFH
s4APZaAXR2eu2RZcrXQB71X5YHn9rE1UBV5UK7Albq45tGq8k/lgmdCDC3z2V7RrOv2qiRTwARcd
KKmZM7ey5QM3kMRfk2hJt2N1ulrJfDcJnlNGbosyMAtzlrb/ZyIpjDCPBH1X7nUm76BRY6wKCQrK
Bg7yIPNT5VMvnY4WsxxmAsQsvdjtq7e43yyKqEPH2Dn89qY7OTpuCZluLaZqZR+3JOTEEwBFvMWI
Jjp1/GN9LyTLcauYKWVI5NlVLbU0vaJgOnP2U8hWNDlRJZo5/35nSEdz5f4H/x22YrkUO2iNisxp
ZI6tRpg8jIpVuN37US5mPsT1/gZl0MAm9sZY3LoBwHUJeNYTvKtjePqkRibWqgNo4wCo/OySKZa3
CLnDBNI/j4fQNeQrTzEGxH67YI2EVOrWtcpSLAic/xrDomnWoX33DyvNh5auit4OuCablNOCb4rX
SzSPWyNaRYpV8SLhPe9eeva2V2EHpV2w+b3RMJ5o3e2cGAHHuOFMw2QovdoIC5hyBkc1JWtYGGjj
1/QD8BAbS6hdLgbefk9RRfBWcAfB14me6sPUQmPnXwIUaCd/ZKZBfaKfLrGi0O4RP4FHh8J140Ms
4erWWatwgy1P0A2n2+TqYSL1Wa1ke7m0Qfwguis0t/7dsoKp8rNF+5jS9Endqta7SRYiLK872lVp
/swg0zwUWg7JBOhmnGWne5aBm84NeooszDJVhN+oQc2NSbbEcBIikXD5sqyLs3L71EVDmNk2qJC0
q0SI2dpxygiWA1SaX6ZxgV3UqvJglpM/1j5TVkSFx5mYAIM2mKv2jnMwz8/rWxIA6C+/BXf8E16S
0i/32xVLBdBNZiikc79zAK4w+c1glQS4JcS0N+7Nzcdgn0+VL050YW5V0ThSzQ7XJhFrEW7pE3vv
H+23+16ZhF4W7S1Due3kSeV+ulIRSApaRD1oBPNQkCLM7dHFxySxy3lHYc1pWhhTgE3E96i8H/Y7
RfSwh7DBwkLpf6MXEQpxm8SAO1GXE856j91t5oswh+So840pmzmK56bhkf0zWpRVS5en3da3ZMdN
4+Gf4/pfClU8Jjumn/zqZxXjKCjVaZiTjDmRJ5p4afyH1J8qwyV1UllV9Uriw2RUv2fNL/vP1nfA
DzC+7QU0I/tsTut3ZU98PyvpFddmIsdt5X3/Ze7lmUF56+qBLKNqN1vkSaAmKTVbgGr/xSLzOpS4
ic0SqlcruqhLgLJeEwJ4WBQYDEQqeR0D7YgY9SZEDgl/mqeyXI/iNxQXp6hc1p20cav0IsSRxZQh
bJi1i1v6ncN3pYosmbjT15lBMmqZh9XeQI9tvDPMCaLk9gK+u4tVxqXEUUQBhXVaGmjdtlJ/DvLw
SXRucdpEpIuE3pYIRGzUsp39AwS/rrjKMCfCBUu/I2oCT+lKdGmOLIXQGUp9DIXcwXlAetnhBPrx
WPV/nchIaEHKeV1eOXKjsWOT0UUxOyMde1Xo8pB/bIl9ZV13dQjGH+23AI6vuk6zm1hLsacoYuQs
bIMv1HnpsOwc76mtahevHtxVkXMYCDF3knBwj1Ie2VWCwuUKi02+lLKEzV1kbgjsl8FY12M5tRZ4
tARH+Zte9efnEM5zlK8JuRyZW+2omOuc5C9hA2B7VXrL9JMU/nlFsjFFYKS0scPW0n8JYuvE5Z+p
cfwgPu9oZ1jfGl05Hy2sZTKLYUyWAQUOGAupqITteOBNafGJvhJ8MA4aHkds75YeY/Nqjj/zY8mB
QBa/WnfUQRqCEltWZdAXItRGPGslVJfQlDCkkC4G61TUI4PFHdQLqUMW+eFZ9TLMiy10NnjuGTKT
JnPmskHYTWsC3uQjdn5uceFIGtc3dhwgeKjjav9FMKrTqNdl6NQsiwqFAaByVD/1t3wpalhSboMS
Dq2CKqDst1RN4DHC6u+5UBetNtMPEDMi2xWsfNP+LfVNxj45nPf41OLyEYKIFKoyABr10QTHBO9H
6WE0a+g60zfEwQAvATFJW6c9o6nb+vC5wAcGwcw2FRSf2YIYJeD9uce8GCylWjRtadJ02dUVQ+JO
eXFHwRNnqV0W+RHTV9GsuouwhVcTukErNgfk3Z26EKQpc62TwCf11gKiyhL4iskmjkf+/Nmsnt92
VbllyEyMMyxJ4PzqJUenBblaFwYfBI7fwuJeIy5yLNBVERb6f3/he2kjVcofWmxFaRdfQaqsT8RF
jj8fZAl+npj66MgZWhTzGPmlhCi097dC5JCgL18xVdNZFLrjs2olJelRDc4YsLYkNoRTKmoZwFnW
OBgBFzxYITwaW7xwyTFsnr0B33aSCGMAxrUerd4mlFRnsT3++kq5sxTB0N+QCRIq8WwV8yMAXMJw
GDuM6vnGs/ymNecchEhPeqpUxAT9eSTqS6HfDEf/CSkFadtqnUSoxV5eS4x5F+v2b/JRF2hEknbM
HHq85Ovsj6f7TpBl+zIEkQl0s4LfMwqEcAIIjCLo99tILL/ht5nEjibvFFy6ZO3oWCo/zfULCXsN
b4nn3Qkrai6gB5p5P0myYA70TSF2Pwas+wVcckt6rWZnvSJQW0lqZQcqCriAqFKh5n8AlvVjb1RZ
bMPbQle7htwftBD/foej/zcJ2YDA3msaIuoN1qypwY4GtMeHVTl8SOFMU2A1buYdboJMLr+3tVkg
Ckx3mj0muJWoY6AMRqy8lSuewGU2d1xpWwD8cMsgw2Auvztkn8sKr/YAf6GYbAVy7zQj3ZWVM4q6
1PG/FLteuIpyGbsdZ+SVS6LukaOocX4pV48QyW9dbP9pQqt2/KCkpOE/XAXoo0JB1v0nek7argaU
LdYLh8gbmNnZwiI3nDYe0L6dAxA/u32F/fYdpjVf7/4MTuxY5CxdMPOO0cH5J97bkyRxph6F17tO
cex02MQkO2KLpwZs+nPuGgSrImENGl2IiNp9DFLIUShNkGWwSxRdUxMNIs75aONHQ2TLpKx0NYjL
EQAxuiIBaeXojHDf3m0/5Dr0dXxKOwTpw1+3XwDZQDlA5Y8tC+hF+dpcuCnhkULcYMd/BUbapfKZ
cBpervbngC5G5HTa7ZKqkkwgehmRpaTpIAuh4ZppRiB1506i4z32/szWdmJeT7rP+xibtuj/o7Xi
twdGo+CA3Djupi5MRb314mvFauf83ChG1gtovYTHygs2JjGiC+ckilOlJpZd8yVT4yQAjtaBdmkZ
6TqDhEOETwYs0mGU0otqrJNDptE8dfKhwxTD4b21rrsJ/JDbUtylN1NvKB3FnqrOVOl6sNn21F2d
SEuYFNpWTQv2lHLKrPHccFijjRPGN9mAUpb4VkFk63bRa+bInLMcdEOEv92bRgUjZXXwMm7l/fyT
4sF8fw9tSEhIgKnn1gYS9KPljIGUftLLc6YU1UTYq0FO2GcyCMCsjXq4T06X/vUYdQ2pXS420o1P
e+H/u+0yD0P4AOj1bYwsPnwL22szF7o5CcU4oSyycfyL0Ork6g7CswQ3XEd5qg+A3SeBcX3/NpMc
ZS+0NI6AvIYtj9nVk2M75p6affeQ8Vm8rAZIf7JhYgj4ZcujkkBUATZwSxuy4+zwvFshiuSQzatA
WY/ibUjKuW3RGTdgynhhDKI6SaIHqDbdqkX88o2ewbJGbwMr+tzWWxLY62Voj54GdnqDwcwoa5VD
9kuJJZYa/rRBdNxVsXHW/UyklVvjOou/8cue4dsUu2LvDULoDfiRz61EZlFwnYIqapntvGgKR/6e
Ku2Cu0S7NeG+Slag95TIfLJQ4Zit2IUP46Ulyge8f3UrQe48ujCGkUnJYX0bKOJDJp+U68Oox4Gd
ZlpFcEt+cifO0WH+upTiFEGTBWFnsv//P89YQnhD+iqtZBqK61flVcOTwPHg3CibJJh3Rbae8T5f
9MUG33MwSrTlEfKmTnabTKJ1ibMmoHGV1biyx4zjjQX/unh/45T849nbsRKCpDVwHT0GtOT7T95u
fRh6TQZAeoWJ+PKxy8IA0PoWZbmcfYWGr1FOKHpn8KIP31zLMtTYO9wi8HFS+jIAnqqsLxBcwXc3
kHQU8/BOkHhbE8hI+BnzfGF652H0aVioELj4Vb9h13Ozptsa7Rz0YJ20klsE37roomTmo9f9QuUJ
8mHXrFOTNEDkVau0CehoIVDPhpfoJzLointXCYAFyuby2uEFTEx2ydUO3dYXCv2o/Qvn9taMVkJl
RwbJAR5lHd/GcFaxt5nqfCRUdNaOsRc9GyuLAdnbYZo65yHsbNllMDUSOzBpiAPtA6NDld10uYdC
pdNFiTu73lY1UHJGtZU/faGkps/ecQ1R3dqMtOCqX//pYFrsJGWtq8hVLkAVhFv3f7zZYLYa1HNT
zq5Yhvf/M891oSfXZiTcuR4P4B7Pq0fM9xcPUnF4/mIaZJTpcUpojMIpFSyEIpQ8bYcUJBxNUJ5h
hXojzDr7Cptr4TmDSy2hO+2LsLCclIbuYBDzFY/NVvUqvpCispCSnVyvLpQSSODUV9CvYeDls0/S
a8HnZ1npc0+jIRgo4BUkfnwWAEjdGyBSf4Ycm88xa1XjvapAYZpD//A1wWVi2q5WFKXeOgcBQmYE
kjKJxr/IcBB7YL71ymKA7tw/eMQMtuNeVeqS5YSkfuPnzch8k1VnhfUXR2P8oS/7IaeflZBUysZt
NWWTLtsRNXjjA08oqHKdQ0kjgKjRC8BeE9x4qvPjVUfCepMSUPI5vnDyRKczJrL8yz8wUpZa8uUA
Cgcq7Qca+qRq5YBnKzpwacodmzvRs2kFdz3CYcy+SdLm4FYjYNIMq8sB/MsQTKjs0QUyPozocfTy
7iSJxXo01U3IgZiiTROnYTiP90EuD3SvP1dQDLOjOP+8UxfppguLmfj2SaakmWIeqjDJTzcL9ARY
carwQLi6dNr4w10Ha2dFpyHZh5Tzod6dxBhIEw45w+ACvO55MH9eUQnVqVxnZZn7dcZC3rmg6JLc
5srdaxJjnrhL8CIpgaCIQv9vFcODTSOtVSA7M4N3839BMmQVaAmDtn66+/mHyzWPEynuRYOkhurg
mcgfaItCP8djXsTZP4V9C6ogg/LZg5wHuSi8+77taNEy/0rR7PkjA5oaYCnBRrpks+fq3VvfzFCq
M/yUC2alCCnjkP00JtI56vASL79zzPWiiHKT8JBv/ngGTVGIISE7UY1SNnogkMrF/s1hHKQV1SnT
eOx3ZPH5CsCMz2Es7wXx4GYCbQjHG5P37GeB/anwN+mlKxWTnc5pOSizNXhTiPAzJNKkWFJA+AQO
CzoF62k9udRxDVRIR/YcOWY4Bg8YmUAHnE6yKkh7qCPZAWjKGeN51hm6X8Bpi8kY7pmOa72QIy0u
L40y8bH4l41o6MbI7E8T1Slyw/jopyrhxDenbQyt5he9WdcBJSuUkaSrXqJsmBPIrek5VD4Zcu9w
2pK6zv7Wz8XuCDvAVUqToOG4SdBEz4zlR7JzgWq3JVA2zWgFSsMdMmcb9FpywqqUyKge6Hci3/1K
E+nY4eak93VinLPCDUtxM4rEJPkxBtZ39tumKH1G6LSLn3Tm+6SJCvMWRt22MOih59oCFZhtyU1J
G4IMQmqhZhr3E17TLzXwk7OY8Dzy2cwqhQw3x522f3VrxZo6r1vViIJtrPM6970WG1lIiP1oSz84
GRdvTiDTzhfd8U7LrJcTj/DWREyL8cPQyBEhuExzfpL4eoOI5mG7q+/vLVR+m9ixxJvHlXZW13J8
GkrVpJC2TzRtNuqoRssIOVCc+VS5uTzeG3skDwnmgDuVV3I6Jd5hQdDpPXHEwwR+NK8h6JYcADnC
MFGw72hi8kbaE/bgXMz5P4UV2wOvqj9ZYo8FVFCE/NFkPhF3gW7jGvRjl5XcB8dE+B1yWZKbjllv
r/QGCP7Qk4ha+qrEaw/PmfD/hseYB8LqQ34VWHPg+B8zYbWsMTKdq3+iooLYVx/t4diEI3e3O6tE
3FQvgnQ02JjUsubQ4PeabUVNznbP3yGN4fboO984LtLiGvyzH6fnxFNpmQE60Ki+YkVw4+sg6SfC
W31VyA0Ud0JVRvJF4j0oJn2sRPnphdvd0698yaKmykSI5QbJ1JpJuWDUfuqwAnfyTbEZq1E4+bws
VaKeWzj71B9JKaCAZKrWpuGxdVH5CrbEaA/NCbvAYPvhh6p6PLNp9VpzTJo3eK+DnAidsqFKGewa
cFoc0UFvcAjFy+x0NsW5zb/0HVwCf2zoOakOnehHUDdpxcLsuMLa1hR9yVR/wGQ8G/mHEzzHHgyq
/e8O8B6SZTk0gfwQFu+rSUuh3h6B/iQIgXMDU5yfEVOnoS5ugx5wyzgQIHuxQns0yjwPZw+LnQTG
qOrI9nf7aTeae45qpVjqf4tlgsSIzuBNSJT6YC40xyx1SkrUNw2YZAmlEY+aZuXaWKQAYyz4sOCP
V5jvQE1FzYrq0XJULdtF40t89q47uWawO19CUkPeQfwna8oczOWfTopBlpBWlTa9fHhv5KsoMMmC
wh/hzyr9DcOzDuWopE5IwouIaLXX/BNkI+pKu1E4zhvKAe34FYVx2nezsWVh6c3tco5Z0UnRD0a1
g5fGvQ6gnCjRSr5m0TztHMOvBSKJdSWRm4teaqTYRfAhKtSBNFJFfbjeNMBZMdBbb6zXqr5Stm5d
ajX39RSMA6pR4VaIsHClnmaMEuqnD9hNpeZdZ8te4yW0EtMoSUXDNzf0EdFASYhxwIoow4BTiIcu
uQq76mZtgXeDUBxwjxYR5XWfbWdXOVxaUwPA0nEv9opAnpMJKk24G1X+mu2akWGliMVlxt5a1SFc
3PMoklEUe1/DdVTAg0PbBVEk09NSly3xPi9KF7rgGN2o+859U+sGdoYh2rOZP14wtm/pabjgKOye
pyjSi2JUp4CELQ8SdqP77YD3dvbS3HELAOfx74Xn7Cae7rl27cXrZ9Ynlfjvj8lJD6OJH1GIepCR
vskQnfja3K9h7RKGzrKtqyuhd3+V8QHGdaOd6/EbEAmdvqsxdoBwEFKksUuV78RFW+YVxbygrhcs
l1KEIeJ+Kfs7+Jb0zBWeo3ctHmJGGDHja9jokvRriblpO66JAhSzwBd8pW1A3u56FWlkMiuYJx+8
iFJvBmFroaprD160gUCFzWlcgNBlyJtLmNg23XmoCffgRbux2xGbmrat9dgJIv+Fexics65Gz4Ao
PpRXp5w9TlvhJV5vVSKItvDccoIivZI9I+Yt47LhRwOsS3kkmBLRqKgVGhP2Nmib5C6BzJ8qEdRw
kyp1L/Zp2QG2WGp+RKRCYQQoVEje3Pip97baGTP9mBMpEnQ8xb1uk/WL3AbszbJv1/x96yuTZXsO
nxV/0XKBeLHmQB9TPSqh6jRpsWQoleKYTyRP5JjyycPco4mF0mzFBBot6VP1Ac62o+j1dLtPZQ4A
mAP91dMjyv4TyKjEa7voSxz/1NKHcI2/btsW0n++lqJSrbBkUvTla//8j4WDNeQgciOIrQvCagcA
jaWZ9MHRwU6i/aJrN0JA1swiQKpDZtqnptnps2rG3K4bBeQ8l604wJnTaGP2WatK+PrMGZpBm6Py
jWz2Pd5Q2WcUGrcd+tCLilepIkVyhuOw6vYWDd3vvoipWsc+tvddCx1VhaiJLToqUiaduDjuQ7AR
fJzccoswkFS5YyzNaG69dD38FfQcjIu4DK+qnUDGmK0YviZ7FX7LLoEFjZtbCm/RziaG1VsDn0uN
8U32RN01yZQdo+WWE15UET7/CqN6pa8fR9VpTnlEispKcwLs1nCUgfV93NADjRU+oX7yLvH+cJ1Q
4hgZdP16xf1b3+KmXyGySvxPjQN+vAAQ82uagoUrdcaZj3JbKh8dYc0tk0wzzl+1xjahx+vG8bEs
243mDV4VYrOYtB8IVr3JTy8N6RhlbpdF5o97Vf1vt7bQOjDV4bWB7aTky4fT7oC9U/6+Zi317vtF
3wmeDiE878egqSx2CpY0nVxJwH4Iq+/i8BpbouJ9dkiYvy2A/pyU/jBKKNghiPYmsE4RTJFMhwkE
GvT/eUBRazA6PmpdTZ3Di0ygTXpHl8uwQ0ggbK68sAya1pxaCoXgMOILulmagFkaslpPeEJar04r
mO/fPj76a/GNO1V3p+tXxHcS0gMPZpgjfF+eJmhGAC8rIGwm4uXk7ldIC66pbVlq0C8/xVucvnpM
0s3GPPKJE3rs8vifY89fYACfFQNweANQhj1P93kxxN7bcO6g2NvnZGyXNQmvULgIG3BrHKqAwiuE
su7llX/v0AXQ0vWsAH7sR/LiAm2z3owcFD2nIe1CMHrc/zIrDOVCmWzQIQcO/gEWsioiIwUqwX+M
ofXFhZKyh5Xg7ESZvA1dfRR3a3tcDpVWwq2q/DmTNtdCXxVou5BltPcT6aGsfcNBDijPvp/6ogiH
HqCeqgILzIo1//tfg66YUcXhYoFqW3AclScQ2nGRMRFX5pySqTrk8+p9y98qglH6T6i9mSeR+eok
GOlBFpMTBJCmfa3e4UVrVFuamvhNE9DpodBJnhevzlQTXU8dB/T7U7MAufkk3JzBG6ZzlefC7Mcr
ZVYGxXZqsJZ4gVy32bv+iq87BGQo2gE8JHB+JI8HDper442lCja1TUADqqJjMy8fAbZe8NShK1ug
2bhkdGms5/GKlHW7AmPc4W1SgXrB3LuXilb1mAW+RH0TGy7rvSDwV4p9eMJunL8FhSM4Y9Dal2ja
J3YLYCVGJbip/mtnsxNC0Z+HuHVMrj+47MfIH59kQa4g5Jukgi6SOiIhAC+zDMPC0/mBYBEmp+8e
rmUWrabnppwcAShF8AzdfSqC8PSHBpkRFASloz91whOnzUH9R6bZic/cXGCQfjJfRvzW89CAiRc7
CWqw1jR9wAAkKPx1Ct5cgHbE5Dg3Ww6NwdRGASOQfArNK3FrxEwJfwfT8rC1W9nEcpAQ0zTRlHYQ
As5ELRvaCv3xvcBaj9MydrVxZ9pnXSXQh0RQSdCxb7xBbYv12jXsYidqvt94jR/AJOiY2QOwBqm/
XVcJCez35P5kDZj0QFf0lWXhQ2ddLpKZLBWzKtcZVksZ4tXJ4QbPAgIeTFvO/AFDAEAv3SgOYzj2
UlQUojlpxmLFmE+lKSQRZ6SfIw+HIqvyv9s4+Rq3KjQKVaUss4J8wtoa0yjWQei63IdKmNYcUZov
+Nb2WTnmGhZiyMrR4CkDdong6f7OI05mozLShsCpF0mNUKKbo0vJiOicEa35iAtmOgDS7ClRfO2C
0qOn63jQ71Kx1HgYGaJPe6Y7xDaAFbWuffCGjR38QiN4CGVcUR0/+W6ee2mQqICHg42KMKVKlGh+
25rPF/I8dcVuqnsBE50Td24ASujnMduMr8TkNkDFAY20rIztDIf6fs30eOtCzrsS4w/GspgsvgdY
UESLU08GAZj/8hZHw+i9RXaCDLE5kWCM56hA3pTisCOSegPbast4AZZPiqtd0QutAd+v4sAAoJFv
wWrSwDRc5jNKtV1vV0aqlit0nwdLTjgDSt3UPmajTpHsmye9WaOkLtpfpl2ndkLv73Zs7VvTxnGZ
wu0SYn9WZx+jL1MkkOWLYLRQWi2tT2KHJUkmEMTEV2UM2SKZKi0rTy8GS6HDwfW1EdbGE8b7vA54
hhQT4e64onGgj3C8VZVjwLBmSqBOAoU2bDTy3OZUQyduaPH6XsTYPgWDw1xViu3San2fXU3VDxXY
xATQsL9F1dgEHCAq8jOlAa/0RadjTylG4414W9EUEaxQGMkdBdLxvC2B6wW1+oJZ3nr0wzv9aa/U
O4bjiXNKDj36Hu0AZMfIp4Sm+soSOjiMAAuysYpy2aHfPtnCOE3MIOYMZ2hGZpYIQzWnrUGAyDx1
okFfXRZsBgiZiflgpwIDJXS9voTJ5pbaVCLIeN5r94tACgTKHpJs+E4DXQT2RHImvHotKd8a4Pf4
C05u1iWcHyJV8hqEs3N1HG7d2kTbw7+g2upOmTferQinWKYkeZjCT3ilLnj1EUaP/vzcuJfow7wM
CStwuFJv/ghLk2H+gQeHPDVOhheHHbqyHEh1WGROXOxpHh3YQHvKKh05CxkwjES/yiY7TgsO5xTf
25sQkFY3nCyIvw5fdYM6KnlOZiz0RLQNRH4El88wprpY2Lmp+VU5ux0EhDBzoov5LfPPI4zRKt+2
Z3Eg2YbsOnzMbQCjQhsQEnmiqNFaLxIUos0hgUGiAltJiGHN3bJIlKmWziA/rrnlTaoPPmDF7oga
06OjeO0HB4WjGeO8vdu9a6gcnpAwvpAKfgQwNCEe/HEK7jy8detgsZ1uncN7QvxzzepNSnoGCsIl
okdlMn/mKBJfqVSXT7v63XGMBAYtGEhtLhDy/bpNcjufJFXPIGTRICgz/RUa4GbNlWjtmL6E5MJq
Cql+qH4BLw2ZtZH6Fo4kUPJjqgzOPK4Z2FBcmUC85n0drNilw5NzGTJd1HmNfGhYQs0mN5f4H55A
jYc+A7AX8YHzOVz12FzBHDisZ5kpRoPzD01xZ+9lfjyxtzmR9fgvpkA6dBQBnMsRfPE6jOlSPrBc
vwaebo9yvIGefO/OGtz5dGTE8Ob8W4nJWol7w+poo6VO4FLsL3Bsns1aaRRN8qsOFv00ehG3YkSb
HyIsHTgSlBsvJAMqUzZ8bUkdDrpNqEWx4QUZgPcazTqz6W3cxIQhxAY5jXya855vIJMruv5PzwkY
9uS37IDP9wxDCKDhY2u0YitAr7rD3NV9U+DX2EwNIAj0+OX2p7bMOFh9eNes3g/ClZcZJDxuGzE4
YPhigXAImSTtpsOqhZ6XZeq5mKUWOANlgM3Kkk5fMoQDohTNQMHkfhjS5N5FgnF97bOuwRsN6nz4
yv44JRhcqcrdTxaDoqdszo2nNc1UdRUKRhUPktV5+oyWZkVzTGOWgk3DSlUbZJ7ZLMB++Z8kJYAn
3Yagw5NQFtk9SRs8rOplut/169+WdVnqsxaVFDRjLMEsWrFL91LFEM3hLddT3QFbNyh4crHP6ftm
UW32vMjxzSS55ahE/IEZHgzXmTVuaWYoZUitaUa2GM5FvAw/BGsPazVbI7XlAG1vs+gEUDViijq0
tjwyRoOSscU/KBs3nduEHTsfXFfgpGkte14eR7tDDrEdAdrrltb9H9ISCE/h2DL4Rk8iQlXC19oM
qfHudfLzTtfF6D2Q8J9P7ggAKNLw+VABRRolImdqAG/vCfkWMAGCwcjAPk6oOKNtHsGdKKvNb8LI
Ep+VL4j9IHsVuis7MEiDsxa4SSVfuQ37MC5/4+FYfUhmhQOEvRlnGjeScyov1dbuVI5wGBcj9VhQ
4Gll+qHgyRdssPE25DI5ncZrDXwZ6RATKinkmO6KebvWHVMp9If69K9RKhqFyMZ2h0ALcB2IrMEH
NaAs9UIXNuDAEl5P23nzdvxh/7FYmCy2meDBkJ20aQYnWSl/2s6GpHyK1s0dZOre/yhCIIXVbGVM
FVTGYG1yY4d8Qx4XAy/hWvK2/BIkyn/GyCy0u+WS1nXQBF0hf3nqLBu6RyV1itbcMD7Pwb5XxxEf
rVizrG30mfj5DOq+jhqo/arUDIs7OkxPFquz+h+um0JFeiQxG90Ssk2ZKi5ccC9R7ImXa8f+ereB
DacfyFivOAnsUGXxscLqS6I0xXka5/pUVbAt70zq7gf/WbzjVVl8wHMJBkeptdME6Co+/VPdmW6h
TZppn1BYiV0hFVu029xRS8hNORnhKUHAyB9GlZ0T5a4YsVpiYy/iVyAKfr/MO6elu0KqyIE/a1vr
pB0UFVJl8q8fDWe0zHtYwxcUBaXsIuMHrT7/shMPCmWRlnfNRDddPAcHXDSr59VlHZ+Mo3XPYfm2
CNEa5X+xRJrK962mYdumPzpV/a4O+q16I6G/4TyO9KFS00LQoChBKwpANzZBS4tA70OKuuk/CU33
mF0O5Z0S2GhaQCbKDzQnpAP5GK3KZ/z3jT9Ib6Nz8hVIRfzkU/4ol3dPOUOP14CVDAp3w6Xi5tgb
Cyo+qZU8rSLKorHHF04389SRY0grXT+YCW6Unqf2R+9O41Jl4AuKPy+xYabPItSZHKao4mlZcV7N
jxFgzP/KMACme+X3xRUQrb5+VmY00BwwSQUEHWZD7UmeNX1ek61k9pYL+DyJl5f6nn2rq1izIekD
3ZIf69L+CeM3d5F+0wlat9tWv+6FmAwbGnwKXlUy3kPWA67iF6OtywyXh5we/g0d/G0GtoB0xQXP
nH+hgmi4SIR2M84+ViX9IlhncyUo8ha4CXHqMB2Jro0j1Gw694ymwjH1MG91xIYznlWdtEyBD4TC
4b7zAQJuIFo412cPuT/7XIn+yRsRCB41Za/x3nnl2IUesuwW1GV+nE4Lq2gubEl0xYLbCTTZXQz5
amH2rM0DOlWGkrJyyiuDmUubvxt3gtnAuDHogeu3WnXtGepFaiDcJrjEx7xOORNiF+vZ37Aex047
jr+JfuQLBP7xqJ7pz3i5CS6+f7/iYFAT8b+ooB4fLvEYOvZ2EMN7fc7vkRWUA839EQQNlnajhMTE
936TQZIwEwtoJsxGtppEDQaJGCZTywsfrNGVzkzI7UkWNsCjwoeZA4jIPwQe/jRrCkzkrJOIMBWV
6Ph4Ci2mUeyBjf4FEuazCbPSKpE6n7cCtqbOGYKQG7mSgmXqRtxP0gm3dhAB5aXPZYwmnHBn9z+C
CNPgNgrrKsbgbzs4hMbHTTp66Q/nSN9QG20RxsRY/Kd4VHgev2B6XC1e+ZlUBZs6/xArGNMmJcpj
h4XCee0zH3Fxlrlip8nBLaLB+KH18C54QD/8+kTrHZOuClUZ2205MLy7llk8Q/eBB6v9Hzf/gAZE
CSHKrKQjqWdSQ+NEJnIIvF3u2og2YdShWFf0dHkwNNBZ+qaEBPVKAP4L9p3jKZC1OELmomrWB5RI
O3UrGeLUndJQQlY7Fvl5PQ78uEk+Rjaegu/Rf+Gi+gmjtcAFeq9vC5QkapdKVl9BpQRsCOAYt3ab
8N8QoyjniJE9Fw8AE+XvwYaLhD0kZ2hjUx3cNCQ7km176Y7evN0FwoOuJVfvEKN4iO2MNg+W7air
k7DbSVvhPr3gyUY0Xj5wgqa+zyXaiAeV8TSTV+aCw6v+TGcRbh8bqnn4bfbBHBLZp6fbF5oEOl1Q
3y0XMhKvLCbW1nq6bUn2DwetllOis7hA7p083TiXCjZ77jfmLSIkbuLc7iTnyR1QyjviYM9KyjAR
wajHPeMxn80WY+mS8ue/jMcsHyp63GJF/H9Y4ZeVg+tabwD0WhjCEynFLFw2hGeoWKvBttDybSTt
mvR0Vd55AlgxyydLuLDTnYwThbwVcjbOL9b3l7Xd5v++3DHhVuW4I4Dq/50TbUyvvMfCNGZZhsef
WgXKuDgqWjYTZ0MKyAHlaow5A3GzkB7UMW2xE70TJmu4AweK2mDVepVfpQM2MpyLwt2PJ4F6MEPN
Wd/v17MK/rIuslU/duJYow6mIaWgK334n3xN4C0gQ4RaEBfp6W/5eh1Vyk56dRMlCrIavk9Jcos8
S7HJSNGIPZzwburk3eC+yvjm+GCh9QP5/IpiQ0Wb4dIXg0X9mlQLXAW28oLNey5KPbQQ8P/UxjQE
1dhCjrk/8yo9TGuSLFg7cHcas80TZaW9/zZdlM1BI4tIyUQwKzeFnXRgvBgl7vGrHUeR2k9Gf2an
ZkdVdxSpBTMJxI0Hc9miq0S7Ynx6X/usuSsMp2aCxVTsJu+lE2Nd7q7VkUFjD3AOu+dg7UIAJUdx
TEuhPutK5AWykBuhIvtdWBNFPwza1B4rg8uEldOkgL5tgkVuhKadTr9kddO1Z5nuoFd2/oYeUxAL
slGU5WziGq9UWOb+lwy+ADMGvS8m4Y9J6BxjBdArXXtu1/eMtW+toC93qPHD2hMZKcxml5+gaEnv
/MB1GUjDzGBRWRiru5oMlWR6r2RAmAcMESJO4GcuECvqfBUd0ITIo8tmEFEjrhvjcLMtZZYIl3DM
HwPKWJBJnZU7keXyp0c4xfUhPvTxyU/1e/qA3rLxRNCeOjIa1QpCrEEsPwRlCYNsg8GiBQD9EpnH
yz+fy3f3jJIZUmDvXQecw3KO70SGcCrB4KWYIMc2hTrU5Y/Ghzzh8Rh5d/zyZ3KSkt6YjemsY40O
1xAgYkwClI9nxNr1bkGNaFrlV+7W8P5zaYTenJFAScCB1PBa90FCvSPtVhQw66qnZidkhNX3JUpY
Tfz88uwR8O4HPaLBSxV1hcIfIaCfQfYJNOOdEZptEaZkfk5LRnGD0/SkXEtqL9c4rGe5mmzIDuho
8E9Ibi34slgwwc7Zp6dALsqy1faY/xOomulvW5Q/33OluKWFUv9TTQ20VWT2vSc79AwCe1Gn2Fsp
bmrDh2Xaw4eLE9Fs9b3CMu/cntE/8yatH4m+psuVgNo/OSPKWb8rSt71Sq6xdKHCFE4ih+x8hkex
/bREnUp1A1+epCwoDeSkPPlweTf7S0s/E2tjA2ilkHp4cWL123o9FStjjqobP3sbXdqvHYiuA62L
EWu2SxXnRzD5GtYfDR9CHsmskXa0X1TSl/LrbeFPXY01cv6Q+rHA2qnvD0liOdM6+9BxqmslUNxN
qTB4CqUi0tRXBa1lpcwbaRlCXNhXAMosaSwi+TVUmxVEoMhhyARtTs3IAoim1T3n8H3/nbOdSrYF
GXwz3uU8L2jWvhYgqGwRU2Zf41QuY64egyu2hUp1EKC9Dzxz0+qYJ1lNJlXOBBoeYGxleN40mlop
kLKTR7WbLo9R3ELb6WhW4oLe/A+pK9EIWxFfC843bZTPFiVVPFMWac1PZfW+Z5K2l4GQGFrvGxky
9tHp/yZFHOnnre5fDkpYLxOYDfh8JTvyOwgNztMAA4Fg4+x2bMJf5CgLE0o3XpOlbdD1uFeWijFk
KDULtgIII7TEylyY8VFrfRBQoqI02WO2iiEUnudS25FM9ce1HTrmpw7FcPIFhyCa2SSyhCpKcuQu
tzu/aPRYRRqlG3tOt6XwN9DH0DXPwLxG6t29yXOs47CQKaDVI/2vHMZi41LGi3a2V+Erky3JOwtv
hwnWp6KTiTHeq5ah16tWVvLTXN8TFGJybcBweQqmuuzW+rWzv46axZxm1zdVywtXEXzrxncYC8AX
maiYXp13kbREf96B4vlaPCTP4lO8AoFCQF3edaWqwDr+fJgG0GBfFUfdXmoEDdkvVVdP/V3T7aqv
n8xeF4qKxsxDYhnCrOEl8FO4gVRoVe4d4QkL+EAos3+tbStDd37UkSQAOvqSQPtRKkueNHF6gWMn
+GvwlsliyAbbhJTfXBok2RCOltP/uJG966JsUFIB3dusZk7lQEx/rLmwfKR1VhQc1iJMc9Jcevo+
8w3a7ccAQfcksshTTEQ8jany5OraLHv7hr15z4wD4FyBCGrpSURZ+3AIUNZFE9OhZ2jiwMQOHJI9
H9iJIqTeFtv0zkUyn0BFkWyv4h+2HJhXA0QYPvMS8rQp68/mMntQjLzafVnDpzaxFi4sIo8VkxP8
R6OrcWydbG/9xwMPhQIrkSFZSc2uJGx5T/2akuH8G26W+47CqRS05oU5QW0ZOKlirRsaausgA7tQ
upk5HSrsNXKKbfFZ1y3Ivw8pP+dzM3G0SFUisxLy2Xe0m96ju8M1cgfAUv7xvvRlhqA03ErlSdwH
g3WHzY1bM4ZduEo0tJIOrkqLvrbyM+KuHDg3NxRMfcnyR/wF2+At9YbaRJEkrRXtebYUKPcOJAAl
hP8jInXRLqX6RBLxMzggfAXpL0kaTVTTDxwYERU8GFh6mkXeahdLpLAc+M6kTYOzCZGNXAcmyIzp
37CQLwPrvTtcZs6EIPjasv/RBNFIqzYLBA8vxOtyTAhgxFAc4P6ygw5YJjLhJMqzxYvKLPyDX0J9
2mil+XTCHqjiqDHFmRBBrSTpQSzGHZy/SF09Bq/qW9xbLZ9MXxOn+kisZMNvTCwJX9lU8DqW2cpc
bh7RWQCauN9/GL1TlL7Ge4AO8DlMPBrV82D90Yc/BrLTNN5YH4RipdZ9wkY/WKvXbkGgMbiYmQgk
6RzhYb1Hi139/cAEAR7Y5jgYBdXD2+Zt+5kEHOEztqhG0QFXHU5wX2TiEBAjW23rPp7Kt/hPk2Rh
zTFaVjIFE+HJOFST43GNodRsLsuSilzxyfgzPSnCc+80SgROah2BoXAU2iWmz/eptB9fGPnhOKyw
4YsRbUEEdtuaSZpYTFnSwXeqZNCYcA9nJWrB+36N37FLQ6Gs3Ldt+N22NDFp7AoPt+HjhvD6l3F1
eN2ngphrJikBdrGpiMiXlZqAH47m46PeNzmqeYvQefsqXQNXaM4ACdU684YDmgmK/g7zUGv+QNwB
/WusZ1+5wowQD3Q4jM0IbMSvSbAORhN4LdpZoMftRAViY2PaaSpxfMuD4bZc1fnQctWAAbTErx6c
8HNtQN3QdbEIvi1n4jHEnqJyDmir7rYV5JgGcZEawIDHddnkWFkK90SxeRXuqu+hQKL8p2JQdS8u
5qIx+/tQe+6pUWy+StHcyv9r55UPIDokROF/9OmAbvGnD9LSCFRhFInLXIJGsuAC7vhPuX8Y8Ykm
5nMrpWtrK7qaIl9+wwJLXTKX1ST3OxqTgdIaO7GNFT35VK0VX53n2asGQTa8mWytKhksc1YQXDND
5qPwra38h8MhrdaqPKcSMb3x8ZMaFankfNc9SX9YDdvUD6dWaPP8Tn4vrDd5xKOcZenXdv3KFiCd
8cpJ9XN3wX4zmjzsMzrbuLxWedCb7WY322yqHDvftbEPyx32DED1BeJUWAMM80eLq7sMWt6bwdRY
6eTnnANnSSXtDYeu4ycdLCHj1RCzUDNNB+ts5uWF8205dtAGgtwC0piDivhj/QYiVxnpYu5w4d56
Nkw6wMHaDhi/bTUKTuEuQapGvcn+qxABZimaD75LPAt3Bwqo3nXY6CiZTzsqcfz53KbTRM/FcTwW
Lu45eZ5H7TaXlLQ24z5r88PbTEgvhCzuEtdXnOBScfosnObReVJTcRRml+Hi7e3N36fhlXeAXY+J
FWkzQHIak94WcT/z7oMe+cj61nr77uEUM7VSAG403hhSzTJ9RTYMMvo4InVbm+GecFEC3mwWNuco
mb1dq71PlPxfZAfAJ/gbqYGZmJ5ko5g6qpAQQOCOADTMROZlQQOljnx1HbHRK0ryjF4T7ci6O/vv
9WYN0DOFAXLJzLav/JKjpYQAAopfs3NYdJblImc7JBZVlRpZNgsZcLV5haUHqLE03qmJvH6IfSEp
Skg068YMPsEO0y9gCdsoGxPnu3sNp0q628cV7u2zlQmLKD0PmVXuC4rsSIHCWHaRAKoVqV5iv70e
gYFwdDqeWFv1cuC4DQsKeK32thqt3Kst6w8G3eIL47Eum1F7T0nATmCaP2D7SLk0/Mw0BzYS1tVS
zYwtXAD3YMR8y02j8B+55da3HO3Nb4A07FtnPkehmUK1U6K9LfBcL9WUoEyDI7g2AC4HdnZlEe8p
Na/Yni9kYRplDYzADpUEk/zDADKKBmHqdBlsgvRUhT9zZSWx54TYl279wtnHl1ct2d2ARQeNyc34
znQHe4hIwZHxuL0RHxDjX1l+RbY4ow7QjsTS2nJsChTnO83yioGVPGoBvBceBndCWvI9+R46nlIA
Mr9/PubeZEDH/lgMn0c3lOWmYxqPm7MTV0x3zql23oF62jXLMwOr0fjgGoxbGIivjgDxPG0Wd5ZU
VmNFw1sVvxUFPv0VjoCKXBq6vcHakXVD8ztvt1C556U50JFzSuAfCxNiYYoeSu+VNh7gW3OxYUkx
X9xB/c3P1C578L/eFljgAI/3Z+RnbuCq9EX7WMy8rdUnsbSVnQtylPaqwhLYD10hDCFNffUKMz4+
dYPL7qET8MS4NDsl+A+50zG2blVOF7dizYuhzDud19oCQg38gd1X0vxON1h4HO8xjuAv9de9dfX+
UV8epB5KGdsgaketsCepC9/XVux9LDItqCthD/hOlh7mX7BEoRcZz9f+YAT/Amf6YH6X9yFaKHz/
WQLd7u0b+GUYp74zZnPF1DtTdwIY1nx/t/PD/f1J2EGlQIWPNYNQ9ALgbKuz32/4xaJsXortJRJA
uPVoWW7PnG3Nt1wLu+LsZipVPXein2ev44hYAcLQDrvlV97qvC8D4tiT6yaR3wiDtXiQFfGqKdsM
3oIvKQv8WKk526JQ4ivwUGkjYgRIzrDhzy4Pu4DHHW+bRnJNbzhGNhYE3Ut2DIeeygPQzdBtKJxq
X/RkD6BeXzy7XGdfIRnmz29kMmKHOLqbbFHQpkv/0Z84/Vx2bUQT1aXR2oUFzwlp0xUqH8Qaqzsx
x+GbSwVlqxuWGnqjUVvaeWpAHoI+DaaGkFXMvQq4gF29W07NoLpq5SO2SAXWyWzAJ8dRrVdoRsLh
fNP0WOdicQeHk0RrLy2Vku0NUtFewMYbnrl+QPgHZ0OwrcqHYY405TbgQOX8SAEkv86NIyT2LFz6
dhKHm8zzm+II+Ip4EfNs/wuLhqJCHGUZCpucjgocIr0GUdjolQwYLfmyq1966kEkMpsg02CDv84d
lhDVQuXM7tRPuodVMvR4Y2v9N3TVJ1CdyQEeZal2TgJxD9nvn6lSAGPecphID0Vze55SZT1FvboZ
hXiKbL1YnI1CFbE/g4eVRj7O2JAwvsVa6m9UIjUQ1GzoigOCx+pFj2VXFmHOGnQ3jukWDxahzjrR
3wtoBV14atRdRhy+jyve2vG+6lGpn7XIaSfux4FIoaKCcM+hAjavVn60AiX6pT8SDAm8B4iANAt1
iRz5GUmtB9r//SMMVR9eUdft3AJl3/Cqeazqiw9Dbklo83ogqnkxd2tw0QkJnhzl54NZhDtcu+4s
l7h3Nulr6PSjdHfqxIktzuSiDTt70+5YTdsu7Egjv/fPWgZgFutFbw9XF9Rl+6gLm+ovsLYA+itl
9g06jh5kJM1YLWzKSosUfuoEcH78LdvQynocQQ1noKNUkAYHRplMYbYWv5Sk43AjEAqcF3YiphpZ
ABCY0Y56ZfxQV0Bo0pXPYYsFAp8nWF+oMgET4FTG6itCflbF281z5EgEAfcaZuPw6WAYVdmI5q13
eQGNiHUbFLUb23e/fPJzuT8OK57aC2pMPYkE/1onRZbGfvVbcMvujh3do6vvG6kt9n10EZRLlNrE
M7M+GgQLZzoqBwnW7u8QqpOgVydZ/PXMb62CzpoBCm9BnEmhznP1Hf1pXCTItQwtv4NMV8cKRJz9
TuwkfgN6G2ejAk33XNpkdriBsPzHbnfp9FeRIjnfEVVXNemdnYTwfuvsp/OAvrB+0RIBUmJBSpE4
CzR/HjTxzjdr+UjsmjoNsStds5vOYrvYvZPgpB+Clpbduw1k6i2mwSTigmhfMBg82ewvJJEbcQV9
3dwc2ZTnzhSYwyow4IJ/nELhPYGMMjsSPdHe+kuqAhL2k39LZ/4xZd7VnFPUVDkb0kk4/VGwWbbf
P3OFCrPqeOy7GWb+V1PwRpWHOm+yOANif3PySeiOEmMnSJnR/E/EZjbEZGLU+4JQhb7QD6PutiMz
DkyVcQNDlXAVtwhBEHess9DITEeT3SL0e8XqbC+DaGSQBwAIPpRc7SKkPTcvVv7ga3m1HFtsxRaT
AtHwYsetRItTf8dwMly0aVXwONzBRcNwipCX55xv+0CTXAy+hJCHhrXQmfLu6r41k5xuq7XH8X95
XICQnIAuqgkOt4L0CeRWu1fjlBW30fB/62N9zVJxtWJYuIFZQTOUkCQI6Zl9tzvpy3f+1CGNWBLV
lX4r71P8YQLauCy+4UdbvYsiuVHPhdJaiJFP3+c1CQo05GW8dNjT9xkyH2JEDdcKiKhmypCLkWav
NQ/pzxfpr0+0Ox+vEN9LngkpizApZQAkJ8qfqTJNY5dG+iwl5tCxpe3Ih6gay3fyXb+6iEvJRUll
TuB6w5ZItKp3k/GfpWb25x37Tl8daw0hEX6hb5oDevjFeNPU82U5rt2wo4lFW/AaLAjD2Tfoz513
qlFRT7s2pS4C1fceGRrGMo0OFaQaEUDVmGtQmUtxtsYgvEnZrnr0QOqYvAxs9+v0FLui+h2l2cNT
EG1g/khCxiW83I5T1W6beAEkMv/0ENmuI/0Gd+oG6/occSQTQKPzKdX9OBXSraNqkLz0bQt0BkUe
i79rci01nnl+u2vahq3RqAK2/Pl7JpbWt9PWsvxpwjIc/PazcQwpFQBr2xulxsZnGJxrztry+606
SVd+zX4OcQtL/e4HE3aAFCpMJXf4kS7kBCb/CF58n2H8nlHsc/go3db+8MCO/HDwpeKmjmvcbETJ
YOSfCiOaXlLNvpLHJeClI7sZirrnYw5HWBHJ3p4R04AS10Nlq+nyuuiWiZL7+DMgSvCH569aJVg4
g2BVK/KIzWW0zkEUlpSAxbmpFVNMjXJjUb4jAUNVCXz+I3pxNE0CEPTWh1Fb/VavRyUbcxNYJ6+q
WZQFJz05NHJIWxJ+7VPz7cRxRIlV5wN2SrYmCLIjbosPydQEuufnf2zsnAOEb4MaVFg//ZP0L8Xb
rqk8oMf5ebYorKBDnUgVPHJ9lmDx2n59wk+g74dyS+JOC3JCntiO0etOyjsA97KyzolkLXkQcapP
pw1klFq/cr1xLLGhLMknQMczdXSWjfXmBKLhyLhkvtklJ4tTJ3j76+2NSFlvaprqiGhayr/RqgTE
6ItfrDeweDZptvoroZDWFNkV/+MsnfcGWBtkXk6RiKG9/zR4WNTPiGnCdQr5YsTpCvHGLba1jafw
4UH+HNKM7VLVH98RVgOxJzruLPEeQe6xYD5OKmJ7OqeKx6vZOMRgPqRly880pO5egpz5cPJzpqzo
DvgUhJvia1UxzuKMK1sC2iHiMx7g4spE2aPlwfrs97OHqDE0BlZ8X0Xb96zeYElNw/i5VRNM44a9
kbzl6EU7Uh6Z/LI7nZeK5gnyb5NYDv18Dbxmwayi3zhP8QINJ+iyCKzrvWmB8b0tSXh4ZajqcLgS
RKps8/KvWH80eR6jObKEK73ZXeIe05X+NYcsoPOd9SZfPGd0i00M9vQuO0IYWxLZ1O9SNNLzMm4o
NDDvRSMl3aPLGRC8vhzZ5uU8dA7/LeXeJzqyu3adEtXtjKnf3uWbWBvgTHQlN/z/P2LlphWf6fJS
7pnBmNyJb1azyPJT1pfDZxUVbWkjxEMw65ThZCybsZGDr5iEqrnmWucwOwPmgZscoyvYjydcuXgj
n+f9gb9TazvktwUBnyn7xJFSadQAq6d8qOfbn5xOi6gE9qL6QABJHK2o2S4ovHaWHSQyoQzTeosB
OAH84J96WWs2V4ACoMBgPh8eHckgtvM+Cl4lkGvxJ4Wm0LE4I0pTgNnmGdJj42Yrv6AjnxRx17NR
QnncH3mYwPUozH+YRZ2Sbc4dUF2cKlmSM5bPjmSymuX9skRUP5eYtqBL9s5RVxALtPysz/VtPq3d
UqANsN1LkdoKb2pIP6SOZn/UJ2FMui/IBDAyDoxoo3kmabcDzi8qkXQilaEdEFit0MWBwYU61u0G
ND1mqZNe03lNY47FPKsqq8C1L2PKEUDGEz8pgIXptTgbempzw13BBaG2tawCTPEZ0SJIl0b3BbGk
MU4y1lvFTJBDcTq1lYiklS4HU27TWxfORaPnEbCLixJprSGByeqG/7B3pUnVBR/Ac01m1eOQWoNM
zVRSy5Kmwt3/rFx0Ygmc/2V1CFYOpWFpHdv6uqRP4c7AZZ2pihLnuspYc/JVIgHJvTMD3ITwYLxz
Uz/4TXGhttOQyRiDvXK5A+ALFcC1I5inI8YkTN6E4J/WBOz62k18ws5g7PqtaCZR7PVU2l5+Ak0R
SdzrOKzpmw9OHT4Id7Kd5QM2TjHCEqBVuH+bUSASZ0Oq4XkCAAInppDXhaZTyhAAq16btFJ5KZ/N
PftdqYu07jMCguaei3daDFk4hNzFZyRU48NcT46MQ1mhvWo5qQU0uSvuoJJ+gVGy7xGz/nvaTN4k
djWxWnprhD6AQ9n2WZplfJy/ixzknlEifdJjX1xHx3MvKm4P40T+mIBtLYryQI/7t3QvnoHRPIx5
g/WgFD3HDcLwEZ2hmjpPVVMTgcuWFRvApRFjidGdf42aEU1rzdD32BQGQEPp2ttw0hOflB/RyShQ
/Cio8DgKIrm82HLBQSxH5Sl/kqXeu6yUjPYMVBOpKvaomvJWD5qZQok37o6/OFYd0y1YOneMSOS0
pEV/EB8RC/bqLJU/qUL35X7PJrmnVjIYynMkgt4QJ3gjcPMkhq5WVW2HBuBewvpv1+s4k6IraaC6
tBKCvSd4Pmz1tpqmqiFasEo5EOIxmcNoLZfx8dPKChiktSYYdrXKUjuO5fHFpWWubk3qKJcpnjJ4
KKelaFXCTkTG9atiKo6GYu/95KQ7NYQSKSMfPUE5qAGAN2N2XlIpge1Ba3YruBNUxr/guKDiP90B
E6nRTxbK2PLFUw03q+LOijitAUyOmEBZ0+L4AbcU9Nz7AB/fGBMdE0kIOdIBlxkXNV1XnReimnyZ
iP/r6YWF61uww2Hcfxg3N4EELkq7lYe/Rk9U4q/3hyLC9H5xK44OqmxK3EC8jUsJaP3GxRx76t/G
XulrLbpQfxHwGQmHTkCilbPbzV73J+N908RIq0C6it7byc8ROqjnJ5T1T/17uZf8p7D1dHA8s+XV
X6ADhiBp/wnfJnz3djOlrQFMYegNiR4QpJF51Z49gpg+d6IHtx0o/L3eAMM10iQ4CDgPIIFx4aIr
F2NevGBCQghZPzRAJg/Rq2z/V2aoEcNrHFsgLAJ2MgEMmNendsaSKPrIr3r6+cXSndJb3SGHimDe
sxLhbnM5HGiodDmwQMmXCQbsxb/0WC0X3JDokljfmkCO+Ysx5bQ68k2vWFsSd2q/Uf9e55DvvDX/
tKXyKwfr28zXyeW1o3gJdlwV0xvalNIT/K/EmxsUrRvUbShrSZDDjOW76fub53sWxXj+olHP/eB4
oY2yyodU3rbSAJqhful+EaLCSO+r/aEvJLdw/yufF+75H+HiSVZtaUFXtaDOFJBc7oP+1xdzNraZ
NmZ48+Cbbzj/QHb1L9NwH+IPRZ4aAxtATcjOYQHaBw8lUNc/Qillyd0/b35LDOgUkGpdj/VRChPA
t0VWpFskE2E47bqVCqlTLgI22sD+tucsozGnxfna8k3N0IBiZyfmus6lTbfn4z84LR205IFujUjU
MKGJOye2moj4wDyGvGn2jZHKhc+cpd/XBNWxOCkw0LlkyyvcDbKFLXV4WwLx56/mCtuTTWF+P2eB
y4zucmYTxF41HxeWD94FKycB472irjSTUQ2RnS9NdXf2sWgG6nkECaf6EroxBGLgmKLTQq8Z9PIv
Nv/CEdj2xBaq7UTgXQrjMhiZBPEDmsBXyu4OmCiNKrQQx587dgIqmoTsbZb4VvfvzkbofzNnO4+Y
shLvZvbW+WiAS7Tmrgr3dy+Ctugx48+7zpH1NpVzBT3hc6rA8uvni4WIn5nTPoZubTgDVw/vqItk
tMXcFL0jo8TJFoOyyiER72rbyGAzziIxZGjs4ba8Y8MkPfkDEdQ165bpMmUr096mxMiNHTiuHPdm
uYNYzEsfkcBcyKet4E1qAchKo7R2PMAz0LiEtLQ+BWK1fuaMzj9gpsx+gF2Xy07a71Np9RzNKssI
aLsVzNlTf4ovoqBLHJ4keRjuWdHVI0JeNOhSAB+Vv6zuCgjmbufLHhoMB81xIz3R38qmtl0pIaIh
iFi62WS9AMUiiz7UI9XQv8eRW94QDmU59fbM9pJQdHnDMZrYItQBd//ygKMx4HcIDSsEeBHvImxN
HSwzY9WuUkFZPvLUj6mnRTWPqICCC6v/rwLvwiLeUEK1OxYpEhC4ac7phcZsGiQqbMHHG/jOj7EB
8b9tqxwmsSivYmIHAly9LlJgl+Cs+djCPg1GmX2L8gsUe1oBCn49gKhDrsjGkzimie3cYsmhCn/p
gylbqwLoOZ4bVeqE/fjvVcss1ifmh0mhRDk0DR5alZmMxR6ZdcZdXe1z4VToGLj6j1h4uaIb4Apk
bJfLDi/Fl0zu7RU/b4qQ8H2SgVkksxPyI1+MMdvPjacCfk8BZBaqnetwDA77ztRmPaK/VXJx52SA
c1R+Dqdmaey8eqQfhk5ixb75dpck+DhFKwoAtw3iWb8MvTemX2jazC9UjVxDX9O6/75L2Z5wd4p5
+4H5kpVPjFtNoJfCBiaXVu2ydbpp3kcS8kiwfmC43PUSLK39RDq/qutdjziyBHS2q4kh+3TPGAdp
dGvEGtCKBtVsqX1JL0KrO4k9TMUOAdqn1HCMFNJaTgzLZR9YiLsjg0HrzZGJmixTsw+69L/1b4Nt
q/nRteodr0N9Fxt9AB3swlrOfTBxm6OyuKuQ9TLrw+m8/HGRm+eg5/KJYnkK/d18VnMO0dIfO7Tf
OMz2zMW4TLo3NRzzJ2rxIoZcvNwYp8vXcMJRd3w/HXYhPyu8Y2VeeqFPrdlJddgXY+RAmH74qIOC
4puuMjGeOvyCsbJotzu+sFdWdthPuYHDpcpiX+/XKK+VI0Q27qvUjJX8RydgWzbRI6T6ORtnf66c
EgG4r6uHTt18hyu0YxaQuditj6JUmoWsk9ET+kU3HghoBsToDwhVIK0pT10XCwU30YspIWvcn7kk
csAh/kR0WA6ntRKarKWlVINwBzzlFKFmfacCRzlQ2Ine88yPN5Wo6sxg6wbNt38Af15I5iDt6pPh
BTe7EpEyu/40DXmJJCBEK7oMkSQLeIv68tAUqwsi+cdHDKZhy+21vJB2uUwm8x2pXsEVi9nSPCeL
lg3sqJ4BMU+OzdbU922ESfWmgqMg3LRbdtWFqOAV9C28C2fYSzxE1jyDO+XIpEQ5zRJ1GrwJmDGk
8ry3eTJL9yljHF3xmu3r9Oro29fKXX5OdLKOXINPrgZMhtp7ZwfiPdRwIj5CkthGU7lgT9oEuGCe
m3eNnjDYrMhNub48OZuhwZB8BQOMTm/86xo+56kof47QkqngHCgslCaUc9rDvtG0HLmjf2HcT43a
/8mUJD4dRuPAEFlmnDR2latKwYHR9p8qKb6Bxe/zZ4ohUPaWvaxSXJsyFuE89lDv71bGSazGpUIK
HNDoCmABwwNwITC5o34bmL9ber2Un6lDAs1dOznZhCX+IDPyIFXmBGR2GVqgO+PBRclYHgQejApP
mEyhDwnE5mtjxdevhsK3UhVhGkp6Od/c55JtQqmUP7WPYSM2ouCDZGCI8YAFMisyb9Zw2k0dkciI
Me8Mu0W/DnVK1HwDg61Hp/NKOtBdBVAdOAhssr8Q/IY375dyfYUPxVRvSz6YsKqJ6nH94BqUSbht
se21wEaXg3YMIy8E/ZSechTECNzP5lK+a2vkdW3Y9qUIFeYDU4m42zCZIF8ke+ojlcLYgi4JrARc
zL0G3I7HqPaJL2lBm2doGgGv+Y3yctFBOKW8k5BNgCRitabMLzDVu8grzrCLh+l31bozeGHiKf0N
nX+Jl+W70pUhIZcZOLOwZywQRqNG2EBNYDkQa3LxPLR463OtoGioQXwuRtIb951RIClsh573mj3M
wUl6vRXMzn+lcgI8W00lUf5b+zzR2DknM3pj5EIqr/iyAqdStKBaueUZokOk+xv2K1sLBmRzh+bs
jVAbv5PblYd6rKKZ8Kijkz6i6zF6U2hZEYkMM3KICM4osFF24hsC78x8qTKRrIzPUx5bgAyp6m5U
mdC7vPWPPZ3v4nkuOJIuLuXUX3bGS/LbGgM04sIcG+E613dAgwuSgm+hpjlEm8vTYiP87jc8WNM5
Oqnc6lgLr3ba9W1ruIDuZGmIyc1VFOxMVpTXQYlUZyptTquCev+IxCCrQz5xDCw/33XQYrrzIFjW
j2oyO6mU56NvbE5lJfY5UzxBSIhyimfTEORa5UI7jPiK0BRA1tOX0Nw4dKFAki0lHdESHgL4zyOz
WgnFfYZNJHFT4x5hSYQEp3OYjOxR4tEglWY4MMkrKPt0K0jrIMvNhLFzg6hyxHdtQELuAU33UsEm
P5naXw9HOk+H4Waj/X5uIYozUvMS4I3gtkhKtJtqy6ZqQs0/sDkQ1vIjkLBpcqrG2Ac70ENjlJS+
MxU0XdN8Bx8flXfwwHJikCy0NWgubLormua5Ypwp+EpV0sPuy0rL5+df3TNyRGf654XhYQzVTYgW
uCsOnUx+nBoqpH48Bc7l68VxZDGUD5UI8tH6pE94LL93TI6TdpKpi0/g9V1v2zzmNTF1YLT1WSFE
CMIJZSd4+9vlgO2Z3l5PjDuLId/oMFbwmsOIgwclnj1BqphZrR9v2s1eEvml8IWdvv4Mm33y0NXE
PXA838W7pS0QN1MFkt60xrAqge23SYZ7ODb1GBIZXq+VBpwWPB26NinLprjbLsklCn2DlcbLJNyt
cjWUK27Y8GjYPVxPSiRtu+OqqVt0jOYt4qoAy1X+U9qKS/xfrJDExdWWJXNRahNqd4Hiy43puNDm
vtlgv8vGObVW5KFaVml30AFKZrOK6EIdZaYN2B07oTakR1mo36J9K6gl4kXhLP8gJVt20siaJpfY
eMfnaCEM5895GmsaBWnibttipvd3k9v46qxSiUqA+l0+63UcUkxejT06xZ13h7dInKrhp2G8tOX7
AvsKKBxoouEokYOCiGSOx/QLY2/zE7DfgBzuGiuTyT4xWWEQl4WxjTtU7li/DvURmg6x7Fg2XeMD
oIq5DK/Z1/MUgpvSeb9fVL7jpz1Nc5QlzYeQSuCoRiiRgZ7sHynHe1qpoaVG+BGknLKp8pD8jtZ9
GCSuZ9LcjmJ/ogb9j6bPxbFFGx8RbsKCd9hzncA+6T+pemkOY+Utr+bOmtCxPsbrp2TCA1YN+0Lp
mT1s34wSm3Seb8Mh5VUzgIqFaBFoeTflRr+2Ch8a+jGe4g7lP/ZQu/tLtrmKvk6EaF1S4o2k74sF
hdBh+4s5SQPkUrtoQ5BYGZKIpzy8PkidKvGqwj2fpQCU6dHh1Z3FfwJzph/sWt//lrsO955u1Acx
kCvPqeJQzPWvwxcyD2gdvO6Q1xDJnmucsNnm/iDopXq1YbJNlTTqKZOraZ386geD6hYkYrhbnf0P
DP1xCsderjOLK4NmRJQitzE7ocvVij4iyNM/XsxXV2LNSSrGFNPEd39ntufT2PFF5XoGW/J0anOD
YqQdCrTPSCs6NjMrYQnSgZhga8TxMD86oysvw8ajPYBjhrujkmyKw52u2LO8PwSebq0FozLTMxMx
S4ngrMP2usO4Ddq0rk1fjSi/3eGgYf3ARnuPpK1hxbZemt8x65MT6kvNowVm/9TsiLVblVqEwatW
LnklIZEkPIa6NF2cVooemV57f7XmVTliu6fFWdNSfYUs3RngY6f/kGzJhzN3TB02YNfJ6VXE1jXx
QO1Jd+Gv3cQZcJQNuCUXxznEnnuYOaIA/WVesjpFXO/xfpsg2hq1NIxS+Pc7SOnV2qRiDL8sdsJr
N0WtsliVRrc7yxFD1uHK/qJaQTgmYB4d0fYACDw85ahDRF+br8irqV/tzVdzASItYxp6kzNwvPFP
gYcJDmmy38DmnRSdnjgDpSajv7kjTfZVxzxXpUHwhc5coWw4CNukMAl19oz0ukvM21UlR4FgiX51
sIvEq3+pbJkQVk1NatBE/ti9casTDuZALHmhWHtzLc22tKWeAS+qc3a1AABkVojmJ/eD693bM476
J8/TRiSW/2wAgqAELrwGC+CcuzePVto8XZ9GechRTIV4/DWpIPwpZH+sc/c1ofmpBaZxpOO1kwtR
QsuWIdRvyIdSMwQ8POXjHJiA7lw/ZG2q2cLRLZDad5uEiW+IHVbYIZnh+NkekIvZonyGFTUcB4Ui
pWxDtHVSQ3pQUVJZwDCjW/3ZbnaeSvgquj1U9Ih0Jgvbcsu8NrRbqryoFRaQujTCgK/yASZaaTm3
prN3KLQQJFsdmmXEIM7KSqnvZC/WvZlUwtbaJC9/wPtdHzxNqSW9DQDBiOEWiiNuD1vuxCZV7tq3
fsNMAQdmvro88NqtHQEE8Mfvw33KYuy3RmhglPt5NeSjTWlws9AexTcA+imkatWx9n8tyZi9nYQz
yAp62O22OM4exLfYQft8vGymr//uMp8+BnfXJtMhEyOayAQ1pEFJXhvUrN+d/9lTfWwglMs5ji+v
/0aSuc3vA7pyKEzzJf2V21GDAww2qItIs+yVAYESY5b8U68jt2S1lwmyGpliYyYMd3AykSwGCfld
ZpmknBDh2xo4TWP44/PheI+RrRUHyM/xyn9adTnu/WAkBvO/psDBkNV0TLMVnmPSkNw98w87yCYU
2DM0Vw7B+173L/ZBgZNGccdlcmVmtnDqgGfZN4XJWf+Gndn/SqmHaOSlW0fAEPdnpdwuBjIBfxWG
4yMRMe6h9/DQjpsAiBJzUwv9eXNHVqJ44etLp7Gj2TKsY/ZR6DCAGugy2m5fXbL4q2yl8V64RM5G
sz7HSI4T578m2iqg9pd36Zo382Bmhu3gRf7oU3W7ybQiK7jy9/ob+qfjM6owAw6Ssv3ay3bzqx2J
5D2wtwhivl1XFOaV85U5msRI9EU8xLLhx1p/jCS/LIgmOG1aSa8za9Ddo3OjN+M9ODwD1CiGetQv
axQCRg+OUh3OHZVbdbKV7lnTh6OMPF5lblaCMC+CpTL0c2/TYhL3hyBKcyckRZZS3ezUOyd/dJe/
p2dmwlk4bUB+GkAKqCUdChQ+yYAGA+s2aSp1IFtsTUSdZwptfRFWCE4JostqJidLExK9vxz4I7ig
mIaBtrvHRS2dmKHpL04uEXMqMZn2CU/TX2cHlWDC371H1ljSVZAGwJT9D3s8pDqTCjOAN75kb8UC
XcYM4/bX4wSzhZ+eAB/WoUaY2nWHrqnhTO37Ey5v3Rr0nhtLbdr+HjVwI55wMdlRWM1NsQXQvxSs
chJhjmo/ZNBR2HWUATWT9o9M2NEPs5isP2WOQgIR6WRChgAnozTbP/0A5OYyXqT5bnruNQRL9j/g
EpAjjs44XjGLYCxyfqA0YuvuQB1rh2APcG+Rtr6NBxOxLlHxtYM+X+lpFHMfOYqz2XG/NfLUuoLM
72vgDVUqhlxMm8ns5LZmVF1hjvw+7OEcKmONCqGOI+EXn3eUZ2Qu9ReU4A2Kw75rKl2CKETxXIUi
98PfHzpZ7L1V3hwBpYXNwL0xIEA9ZFCNohZMPIbmB7/G7UBxEwBEetkyGiSui9XlxHOk6e3ajv2S
vNE4bzVheYAI65l9LIVQDprBaTZgP0LR9c2Eh991M/ETHUBHE5dm55GLfVKmd+nbM+L6MHw42y41
ppnzH0o4w+kiXVKLVYibzLm9oZGVCi4ABXQC3a40EOScWy7NsFKEC5N3BC4cGy7okAj8m/LIwLay
sN6SIcHdYbYIvT3grGyOZ+K30jeHRUnrCkHMSQ5Wl1XClC6yuVkfwhWgt5YXrzkNewdEuyQoUBTY
NhN02M9Dss1PURfHDnFDlv/wcFjfFHBM2pKQXkisOBRjM9CGQ8cYDDcYhiGl5bXL5PjIuhzwhNAm
08lXw4/7Y7cHy++PKygXCiwqVY8sNURjD+fm0/7nHTLG4msFTuNHEMayArx/aj80wLVNYSx3DRt5
fs+jjo/yutQzgZZAplJXmNKuBsZp1/xKeuTAYoQhXT/S0nr1ceJLO/o8hyYGf/dvorVCaAAVzMPw
9m0wlMKgo3y5DhuiR3YAygfhGN+xTbb4Wfj6HSjRQcqqRQGcbI6+OHJROWBS+52GQJOF4UM6j5jb
zFeFNhYc0ep7PhpP3Ex/qEXI/Him6BJsxKYA8MIPaA9vxrK8ApOCQx6Xx55dd0dxaxx6qEY6Lvto
dWZI1p9p7uRkz9GxToPWTciK5bTBDEHCw4XjwmG7MryI6Q4WXxnnke0UiAbL/5bEyhKS+ZcJTmvQ
kh9WdRT4ZXNrdUaGsUoZ4MY6co2BQhJhsZglY5ATa2rzu6POGcRppVyqtKmOVW8xt/TJgnbbJlMI
693blcEjzyYhHTWPQIJnFGFrh94iY5wksqwVbP9hg9iinqB9UrFXBHK/JJeZkdXRrswxrsyjw86U
XHu9BUETe8VW+3/Mbisq1lx62YHaZODwPIsHaJeEx4ZLV7KfAh+R9USTVy1xIL38uD6Pd5eWSxJa
NNr0d9UYWWKGNTNxE6tG7qXrxYXb959yLzun6lf94LeknXPUjNjmGcJduUqZHLJ91ZQaJBQ3Z9f7
RKp1P/29b0YLgXc2RkJjVKIg1D6NMCkFW4+OvA6LsbFdPUqX25JnFYqQmEFOmXTwIE5NhpMsvG8B
oIUsN61QLUa3n5wPatf8IQzrSvyx2r1S+g7BajsFbxM8p4IVtOOfotpvtpfkIgMFpooAgvPzX3PE
YSLNrYCI22zIRIqN9BFQuCf/S/FOBOSMnrz9M4zUwnvEFwGX6sEqfQ1oKDcF/KEItyL9ykKeyKu7
P9yrliVzQX+0DOCWR7O6vRxxe0Xncz6oPNc98o+3ONsvADrUxh3LIwl9JCCHAcPxamWNbDjkljti
V2FAXFskA7Yx5p/D599OsIOcDjJ3oxSvlr7wwozhHGd8hq1LEgMk7g1YsxGwSBWtPwbI24Ix5sx8
UjELF8wRwh/dv+v/ET77XTDCpKQ74EUOuMPv33xPT60k62akJ8Bh0kYf482B39nd3NDrX9orDe2l
atrHpyLL3sizS5rsEhjQwkfrenm+ptWvcKoVawP1v6OZHuZ1tPhkSlc/JLDsIclY306QsZCwf04G
yLEdRLQJ/7C7bAvpGywWAUA92tBXtorU1w0b9l53RlHsPiSuAspWqxPMMnwEqkU/9olCDJNhuBzW
HQIFwt5vu/5huiJSJSp+yASHxCRWWQjuBxTnt//IgSLA/9oqFG4uFtz3HCv9DtIBjTzgRqB4z9Kr
Rvqv7e5WHXGeKBdPo0efXURTC99Gvs/OStkFx/2N6/GyfpSQUFF3Q98BvnEz08QncXMpUnGvb3By
0KPti2fgADtrDtzS21yD6iUKmPCM8c1mvGBQFO7rR4lbwzJvq8yVFaPhRWNmpLR4nbU8n0v7k7b5
AUaJSWQY9dxhXOgyq59qSnZtrBsCTOlB7X14nsBpTaNJp4Z1op6kSVoKs3lXQZfwGweUWpwi2cka
WuAO3p3pSLIQk/9irZlkFWOMbu8NEnwKsTZJtFLM+0Sh1/+cw5PUWWZKqYboKM1zbmHt2wsl8iyv
tVWnNlcILspZdz5EViV8CcHmBaC+EGTLIzQePNxa4F01gbf3cxe/Ef7alpxKJgZ5CMEynxmyjQx+
3hIuIhmAUm/Vcp3QyuR42Vi4/NqK60QmOQcT5kJiIu9X65IjYXUr72s7qRJWcprGtn2VQdR7E/aJ
V8uIRhveF3b9w7+pcwBSXhaGqTd2ctLo7O2HWmhO0WZ4fhhiyLC0neGf9xWAnrxqSsobEtW3+dhA
m4pKWE4cFQ5jgebom2F+/0pkc6ZdCA+3nX3rhYOnXKhiT5cN1zENh89a0V93mnlPvvMq73tShKmG
K2nw2hQyI114K9BActg8c8lqzClNe10J842hAGqKejLU93cNd/LmkIrLOE87I9QUBYii7hBSX8Ac
47dbIIM8ZbmCY/YoJHiht3byYKMGqZlUtDSJCIdxBPIpG8E6SZ6u/Pc56zUa/3EJvJywzD8qWSEv
z5lmoDgX19yAyLq4xzns1Fj474nrG/lsf9fb66HWoiOOTyMSzzwa+vSLR6KLzLokob2VDQTpYBRu
sYydUOC0S0BGTOcnMyPd1boAHIX1Oz3TyJh2oahgGldRLBRISfeHZnJqo2QOQq3jKGn2llqbMZ38
+2tI+OdhdYQChEMWw9vUPdWaLKu96VGlpgB3FkWRkz9XNh9witocFDIRRGKNARGwTO85TLUaR77t
D67gwNWbCgoOMM3u6JmUBZopaIpz7d4ATXsp8vx6ox851ekUWn8zmSfBne4nyNhS/zqOFcyRhCnL
YJS72/sEL1c2j0Lu1xvv8CYSWUP0VUZ18oUwUZIMZhJlJ4VMf2y6pmMMCiHBEoxJ6hxqCcAJkb5M
vFT9bPqUUq8+T0EuJcEYw4iaWlpLm0LxozsK/6G4CZSkzbOEBZu3VCZEi0dXhghiAvIQdztJC1pU
kkeYEXa/KlXSQqdQQt2FDYHS42gKeDPeHMZXsMGAhBxmpevbYbItOC0Xh7vFCM1ZM5eaYgIMMdUK
qvftRHNKfFH1d5ETZMMfqeiHounCfB/eLZH1VVe9yYrj3a5ik5ToUynGj+aYuyuum6MJ9FtZJtNL
98/wokmEJMdvuQyb72a3IjnfThtXrg0NFzNFfT8jDbIZ6ljjsgi8XC3J2PfCaRm/wH1NgFq2vn7M
8K1LO1VZfBGX+0IYwqwUjG65cpmBLhOy/kyy1yGVYYUJjto06zpvb5qHaQwd0xlSWBEQDapj79++
bBO0pRZZDxasgs88Khqcs2AY7zaLNpIwUx0PYQKZkUcbCIJ50tcf5AIlCrBGoDt9GnNsASH53jdF
xyb/KACrSwxVxdS+zUtXJeHRRv9RKqOpdnmrOM+V1Ctrrf+msxWDD8DdWSbo+yzmDQrtDE6sdpjz
teYx0ifH1EL1Xj58qdCvpYn05JwO5iS8a+9RKjNk4Mql+IBuJtNdrqQxWGBMSQiYZswWQag6n1dr
hwy992y+oeue+1dwRSa0Gj9Uys5a5Y9qA6Ghis8siGNRtDVa6g7ABhX8ypH8tqCWTPO3gVjCJ3sT
KQIxpcmxBrDEwEawEYt+GcGty0FFWRIyMcY1u1Qm2EQLP7GHPt8swnAOvAi6Ql9tnWvgP10Rgc+1
r26nDL9wXrsMcpzJXGGwkKaB3A6DoQKZZclHvrBAaNTrKpWk9X7ZQeieJzXJiU3kYpV7IXqqBy1f
REAv7rVPVLNK5zgZrAkeiwX7Y44YfUcAIRdIPsDD2DzXtNt/nP1AleGwFal88llEtQtNp2VvRvY2
y1hqexCuzU0dsxY7kWi1kSR3PgGUM/4sCfzoMx91Ll4ouCQIO945gdT0qPw6btItca7vb+FGku6n
GckhBlH4FTlzgGPoW3I3egwW/+U1nEz/wC4mD6JdIJ1wNGAieBiBFb/F/KOEeeU/gnZ54WaHbBF/
4M2MbDxb7/5klY+bGD4z4HQizWBbnN9YLxoEU+vGdXfRwCWaq+suGgh0CWcnz8uNbdn378VdHn+z
AoI8xWyRnztZ/UhJQBJnky2FByxk6f4Fhjhlice245dkiwzO2jjapurKa99EnhyWehu6uF+b/3Xe
CBt81wPueatVfoL3XZRDoOXfHo1Vml1KMf3KBKgI/NDgqlFYJpmgCFYfVrM1Yb5yfTxTnwYBiQxm
xXWLpwBYv2PfCSWI8n8eyp2vMNqeTvYYU36ArP51lZQmiPDP7CteH18Te22XN/1b/0jnDxNVm8fz
Hc9SrCIOaMwvLrO5NRM2Od+58YIc+5Mk4GWOOYxc0u9Lo3p7tQkFlEDpKHGdgAKGFyQ2nNO2I+rU
L8NE6S+mTDJF9JwNDYLxXKEJBWivQ7X8oW4li7ylEhKJXytf468KJwfARlw15t65WgXWlHf6ztxZ
btKXWhmcCWfO3h4sd4fikJ8omFgSfOHwgH8GUnrCxg/wUjgNuduEm3JUYd5YhwDATEJeUVCFv3a/
tJAGlqTw0Q5XvaYhRyZT6uHIwy89DmNPR20FiZtGZVoxrzFpJsI6FEmHi1fcbCSyNxNbO3k5ISv2
s7/lMUushXszPqpDguaoK3H5oRqURFcV8zdNWGo2CkVhVxHUK56fxlYmH1cO8mIe6b5tIqdj1rRG
zE7PNfgQgQqXAlidJU4y0sosUbrIYlHGObeZn2hsvvRCNaeIWXoDY8Uf70QKecBjNJx0eR1Ydxky
yaFdjmHDUmpDWfwknGKpw2TNdzRHpbo04ZPsnnePKwUniUIPZBCBOahdclBvG8OF2A+yqeFvtdHX
zqrOXJe/gdpWlSCD7BpCmpyt5qMPizqyxQKkty9Rd531RUsw/WY7aeZq7H/BJCQb7FtN3wmC9WvF
HN0WcgSa2IhiCbUiD4gU+28QSvFRprTwHrJZxV8Li/1ST68Xb4T7Yl1+ZttMFcIxKqVU6jhybqBh
GQAjQ4oxUC4nBpEsYBXVohE9lJ31MGlik3Tu66asgsimCImq6w1BFVV0tH9Qjnv+HytuOld4Pl2x
m+TF93sA/dbE3Vo4GLNIup5Lsh6Dr/inP3+4LUPMTmg1vD0xmAtj/A9KXwH39KM1vx8DYe81BfJH
bbe6Pgq8FcApV6IkVGtfRhxfa1nfwt2yWijoOtxs0/wxaXhBINqosf+Gjs94o6AXB91kqSRskj3T
SQlAjEyQ4ssakMT3PIPMnmxMUcerW8gC8ysO3Nwn+X9A+NhYYgs0tuLsdDD1k/105c65AT7Gykwx
fRd8AR2ItL9Lls7vNxSOgc0y51bTh0H9iHHpWTiPVlREkzIIcSzVegoySaho4J7OwMRkdZ3NMHrU
SpoE8LtZoRcHDNrzz2mj84O0Y132DLihHm3puZeaVYx/8ql+a+VpDYkWMjVXnef8oVI2zD0V97O9
6KqH7XRFM2/yP1LNwLXd+HKRILfWtFLKSCGRC34bPwqavZd9v/u2jKiJeOoVMvE9Mn3zy595oXc4
s7dmQgsg8KnGiOc0xHQdMz7rLd3GCbafRNr7VGOW92l+ANLyYLqxh21qiwWKnM3zudPt+1GhHBZE
uRMUmxMLkR/FoP8dBVHTxw+YcC561NBVIOkX2i7mjzh1cC5aADaHbbjM3IWcpyu7QNRzz3T3muua
arNhJWuu0TiqNTaPiyWpu4r608kUnswCM1of9+05ZRrSKbTpumeGAodIXVLrwqH7roRM0SNSCMfM
43If71+e9nYIvWapg6Z4UxB1xDkCVwlOnZmKYaDwUbSbcSlxlVj335mHHGkPz+y66natq1OYT9+9
PseYN9v2fMsLCPaMpoyxiaFAVbhn9rKGlJtN4ckR5hUpLR5RXJDkF4kuP3TCqla15Wb9m1VXiEwy
oTYJyl9TEckZLqmX1opPMe1aUkKQ+i0qv0ZcjiI5ylyTIMZ4vkBDaAzVzk1NyBDrAD5tmenkce5w
U/mnRLjy8lKpZtuoodvv1DOPEKCIbtSVEtYuBnorZT7c6U5WjJ03OmdCQjYT4BENMVqsuOu8GJ3u
p34zGL5v4Bv2G4cy2N9rIQ/SBWLLBR09UfHpLi2rAVysHep2k8sc/X+lliMyL39Y2V/R0lFuENYt
YMpjmtVy8znGWGvdqo+UGGgDapHYjDnTN91ohWkqAz+4aOkySWkT5Z+LQY1D5EzZpYi+VYceNUlb
YUNe+dV8GYnjC7NkG0PAJUDyC5Rk9a9xEZyVTe9lSKht0qEXjJ7MvIeHtwa+MjCPB4XAQ3BVQ3aA
FJLfWxeoVHRV3XiOK/MCayHgp78GK1LZmBX5nMhvm4s1LTDBEgpwDii+MFgug5Taosjt0F9ZXtay
9b/KEpQbBuxCpWSLZIZSePx/bGv32/DUSuT2S3dRV51K+O9Q2WWqLtylDhYQMmBP9w+3d09yKnr7
45r7StU/H55TxthCYnc8RBuuGctSHXsPzOdmBlSGiwv7jb7EUJq3D9Z0OGsgyHlaWRwt+srHzLXw
b2rBwmwLthHwG09okCJWVRMEY7lPkw7mvI1TzKR8qMzxuXGfpGmP3Mt5l3D4Bk4oGNjDZU+prDgT
R3lN8rWLY+kvrNkUnJGiU6JXmhSUFBWp/aa5NnG6HRsxJS2PiSuILBCWRvTOVBoZfQikEtpJbMA7
0bm6WmXOv9z9U24GnMfOzuq330BIiDn3LMhO1uBP0X5xs97zO2zw8bRS+3bkTwsDdF46Hov5NwGL
TTIIxVu2qT9T7GwuPF5CkzPncLoLyV4QcwDdTzE435nJgmmHSbnYBJlnKliVwToBJG+XZRevVf9g
MUa1cQU+zikXzcw1kVNqtJFIGNxTNLHmGyW1ULh9aey/JRtb+bWwFDWAQe0Y/jldcRHnZ4knktW7
nsXZbShOb8sHvK5b/Z65y76Q1gigkcQzmjuYwdc17DF8VJM+0gjSSJhCpqMtbpMOj2P4uH7Azp1i
gjdpN6o/RgjhXI5t2u4VCmeGivcJZDPn6CgaK7nGWv0l/5QOeywx2u7CuXJHAyc0Ob7Nm19bfg7X
m3t7lsRi7BmKFy+Dwwr/HX/zcBqH27nZXvQo5OE4rEtr09lQ/EphY/C6KzpRafxoUuAdsT9IYJB6
hGPAw0eBQgnYPNNXxT1xUxwFPwNHZ7ma1lCXD2hSYTRascoBwetnuCco9it4sbO9NmNNBbsDK4Hl
A0T+N/roSQfgPdxk9/j5yJKQ8I+kTJZvpnh9qxM7Sm2krpxl/+bwUmyVX3HH2my1Jwdngk+y2ZIa
uJ8YWpmjVYEJt6BiJX6rA4Z9dj/ePRs3X8Iz4iFa3HsBTM4vgwDPEcYO0Et9DK9NMf9gvW9Co9Ah
oBWOMMn50+exJSOMdDhCvpm3bPWTJm2qZcDb9baM/Xfaq+j6B3POyZ4XBfW4GXBOfk4jUuGwoBDx
IzI9qV/TSR4GfPlO3doxlIlDlpfeuqbhL1yugOEk8KcDJmt7vE85J0Dag5BZ/ysR6dTpEet5srzU
0qcbHle0ZOj/oEIFWzxSkFdELe7LOaRMXHI5qsXllyOUi0KR1rHBsQ710mlg+wK7WLCdGM7IAJ8M
vLpDXtiLaqYHKP77nBizRamUTQgDdcEi4dFl2pPK7k7fkIH6CudQ4x0I9jpc+tIqIg5ZWUCJPcE7
uUCWbIlHcALB49wD5k8y1A8pBonzkxV2J7YP+NmHYcbVsoI5OpHscpgP8NoYFk3frpg4BfaEqs4m
nQaOTKr/u4PZC7IMX3mJngPFo5XHBiyVm8kjUosG6JIn3wWaNhPa36W6wX9qdYFOKAaD3sZEQrIX
2zdS46fWe0D/6DLGBwShsL+Og6Rog6HJeCi1qzO/3vU5ApGJgtCpHc1+yo/Xw5+QU3qmZZo670RY
q+aDU2Z54TBxA2kUhltvseUFVpxl748wVv0z8EJUnzHJcSGi6ugeZb82qPnHPFZ5nMEn+hDFjAaD
ySXEJVn5dvuuu+Rz2lrxhRYkCR07Y1DkcblUWOpTRY7r/XU0WNvWI1u8d0xVBwOt6jgcTlMALUoy
D9v9/LWsaqLKhfT90cdKV1wffQ5GhfNSsSBCW6/TnNyaqRAp7mWc2XrBnvsMMFTzdzjZ4BZ623E6
WCSVdQyP5MN4idFEU/qPjSXhu5JHAQgdK/cR6WpQ/IJSPjfJb7JypxLJlpVr7WOVYZ3HDyku+cTJ
dgb2SBRQtv/6Y5B5pkIbeCFjbbCphXtSqNGimS2ZDTQ3qvRwlPOnS4Bcfqljkml+G6Kg4jFlYLEv
xYGApv/S8ng848ixPTtuin7m9QQIQbyDNw/a6xPdPV21hJV6NHP2wlqN+iFk2+MPZpLcg8LSphJQ
zpqpTnLed0sD62DsdWwC2ByfSHf+P5xMjakxAHNHaD+JoTXXfX0mqO2qNnFoc5VHXKz+skkNz4bw
ggGFFH+dhyof3NxNoU6AAjtAiqjsJpDS6vzaOV3TeIitmTGjiSGWpzZzPnVblAR9LFjTO9OkdzkD
s1fgDszEoHWEl9gMe6GR+OJtoNaaqRDtaXip1B4B8sVnbHc/cBUqWTS1/9knf9fdrVl/gvQznQ/Q
iFUJ4r04KehuasycQhut31H+ndtbfZyOVVLmLxf7bbVgwqlBa/yVKETyg8igMGQ05Ae2lP6oQW6N
fwUSKVS+RJl90iX/MUgk63UGE+Hhzu6H2Rjk3UlN45Vj60Eb9ClidLSx0yvzmlz2hFdnHVVkwYSC
Z6mv//xaC9MvmXO1sc+CQ9W+u+YScgQXQWx+s4O7P3fXQE0fVHGVXhQNzcmtw5iSVC4BTGyWPyDt
ZYuDZV2+JvCuNWtdxke2Xf2bsUKvIUh//ou4DfAEDm1h3KpjsrUUyMwdaUjChvfyqVEtEBRJqx8M
2r/gIVeJk+9BTJVcZ/ttjkC8Gzb33GvDXkMpcyexqUPDpdlYxcPWe6zkgTOzFdGjVHqeEWgbSmwb
wjesQVaqVkBqjXIqStyGtR13lzNxOxNkH2H98MbRROlV7FVk21fzKnc13EISX3MXkC0bR+uaUVQq
30TCkILo1Y9kvj4b0WqauqFhkCCef6JbKIAeVUJ+oLcmhGoBsZr1dC0gJYSZ3LMW12Qn/E1f/eoe
Kb4p2+1dCZ7GrqOUMKQ6+gE6UNyr7tsodVl/k6xskLgapJ1gj2w8XMcjsGjikATKlRs6cXFqUz8f
h9w2sz1PqgYsNxk6TmZ0WkuF9qSVnu5Lgbgx3hjvezCm9L7U0OkoXDD2avfkUF7czxEmtIE913fB
6B9zXMonPG+mqxIT0XPnalZe0BfDk2krDAzBGaMhzVp8At0/wUbhDkta1oluZWLocmeQDhz5j744
3tHR/gn0V7+qTS+m3N7R/SDc352SqL/NH+qArbctBhUejxyXLJGjmMyVoOZrnnVzPeHeBDBPoYVY
YYLrNqQqVXzM01XXXv2Drce2VgqyxOPGab6mRnb8/hfHNH9D2rgPfIv48Blwj3NqM8WmYqtek/j6
xSf3Du6tsEPXuBI2HqiKo56TUMFMOcMgnIDG0333ehakmb6tq9SjO6liZs/uL4W16QMq5IsPs/79
RUp1k+CuEOFDdDSCt2O0Tey/+opd+6UZE+Wi0yctiZfrShjY/uBk6BKaA4Vl6YeeEjhcnStlFMz2
0ab6lfEeva8XhqxX2EcbyWhaKJvVPfJ8wfJnhJw9g/BHeuA6pNnjrgKnvQoEmcz2eYFzGHGt2sXs
x/D5Rfsyg3UYqLkPD7mU91JT/NCsiJRvG5v5cgGytXNaMW7wDsdkwmthmh7Usrpyqs2o6FSwhJHR
OIQVE1XqtdAmb+5jyTAEJQxk0FriLpXFgL3skzPGJVnIAeQTkjTecnt2qU+bfe2xMY7Jms1nQkuw
hxOC5Pd/OAjQCrEk3JKafLRJsF2wlfpGcdjE+K3STyWvL5+Vsv+pjCfAL+uP1j/++N8m8F1D3FLa
SEqdvllY0GtQEB0gjuCOIGMMxxKdFKskFyRaHyKARf7xJpsCtLYvw1au6A7oHT8/X8BExebHqQfD
VkS7VaCP0lgGXNUY9E2Ywo5GIFYHIDnymteNN2p0H9ujm4DMlIRJ8PhIPOcs516ZVTv1saOPk/x/
Wf3Q7F5On8d32bwNxu9clCkNYdXtHCWfLSzbc509jOmXtLYAf9TKoNdowAQ01/aguO3sM6I080C7
+Leuys60YpKYFUVvdF73XnribH5AlVO9FG5wg5+6JP+xEE9WKdhO4xMEaD5JOHjwoGK7C+ZEzpg/
tdgvxWYGlxVRMsvE4mh02Uh7Bo15Naz8hHJMIMK9a7GgQOnxtlbcX5nbLRe8BVFVk53017rbe/aD
EBnnEnaokLOnZh8VWqo1ChzFCClse7UYQXPyHBF3ewQUSiHMT5TzPhQkh7tjAC5Dnq04illtkhAF
kN6CjNSmCzplSmUaildCr/Wa743y+pngV7K9pWDyJAdE/6t7M0V8lLU1vjK0tirGCcAFnr1jjoXk
RLTEU+qkl9DqBlTDZskheM1R0K/BL+oZ3alcqvc5KtR8YPJIeG1Ex1AhBVEJFfJL9tYVM6YEox8J
knEC+bH5SeSPpzGjli1sR1MH7GgwuZkiO6173VmCrFNpTtJF9ZhOh2t06osWaWEf1I/7iaHov95D
Qtju9rcJKRgP8A/txCG3H4zUhvNxqOy5XE9YyJ+WbTbvMTu4w8d3gDb/M9H0JrF+xKKylSMogqzS
nSqVf2w0wxu9FrNkg1oXpuEGMVeJjkaAQfmzX1Njv+XcRyHWzVWYviF7VKu0wdWKKNINdFlFOXh3
ZqIhbBWNIPNUU9fH2p4OBdh3fShgylJZSJWIOj8q0NyEij2n9yUYmjUA/RFO/NB2N0UWDGZyiNc2
qKVCstN1K8cIZw3TVjw5mgrlCDh5hC9AXKaW14cYTHAzUx2VoryTsxcimJN1nK9v/65vwp4N7CxJ
iHwDPEDeifNqgSitIRQZrTpAifx0OaKV/qKhslxr/zjUl6g0pQbFGNG7mIaJFp5G4SpV9vEzxuUB
G+E5ZkppobI/OVUaoe00+L4wEWv4Gv/bMpjbxDR4I25ryMJDBYqyzjyZKBFQGCA7HacuqiR6zXu/
ni941S68nKVm2Je6weL/L1lENjZaNT0lBnJiWn9h+r3w4PY/TOi5uQBopa6ebO3yUxPzPp5qAitI
r/tV1Fs9gJuOlTwucl48gTmMiTuKZxPjM5IDBPu1LMWlOx7N3Zrs8x7P6bbfzPhyO16WM4UFiYUr
KWF469CFkeMr1S6dROSlZpJ21A58TT5UNl6HM5bWQPmEy8axs9PKeNqBfPb49ljBB6T9IOgT6QB1
NDoynTvn59EBrk7g14/lrIOg4CMV9llB16HvhBZ3bpltfHb9AOLq7qgQtLDfPl/8UZAyR5Tyt9BH
sr74KMLw163hUxY79AmXcalH501YA/WgBREbWuogpE9tS5WJNRoLVYgdcuN0MlNeXa390cZiz68I
E0cxvTSZlU6vMHDkASDaAU4mxgTteEU0pfdzhM9PL82xbJ+qPM88yXgjSGoLTaASuefGvdla4ZhV
F+dFV0DwAMfU46Osy0R8xKgPUJ9J3FSljhf3/p0QHhXnsh5nMsw6JBppS43LK5Y+6PiqXPkNJ9nc
Wrl5pl7jIg6wC7oaLslpWIA3DvsFzSCU4mSs4E9fKU4NDOxKlnbCR45ptRE3JuBBDjMJYmb8wwly
ncmRhALs0D6nMtX7dP5fOSKbccFELs3lkas3TVR4ZK7JvXw5Sq3iqFgB9bgliZ+4QAoXJTjgh55E
k1oQH7L0dsgczk1jqxflQp5edpqkJF/ZfCWeqwN5xd7Z/YCyneLbZunXAqzdFQzQsZz0zH9VF0Tg
0Ttc+w4H/gkg++kg92Op74sNqBpgvcxrHb5JvEymNKOzp2RhHxCmDv3z8J5v4m2vk+DwxNdiaTVo
AFNnmLpwPUvqhmEjLaPwYV1WIfYclXH22v8cLcJeJVN9pYLYQAlluztls0MN3GhjXY7eBS4mMfGT
rZLQ85p9SfFePvIf8Yj8pYfL19Lf+Lac74tbWmTAZ/fcyyUgrcI5/eFdskueynjoo5YLqChrCuyf
DsN9XythsuyLnUEYTHH89tPI3CDTAJnsqP8TxztxPkMkNIRY8CaaNB5ELrkzJRTEuhFnn70dGXOx
4WUiQk8zN9yAM05NmX70YF5E+fgQQsLGrOcZajzx6km6nAc10MuyEz+MPNet88x4FhEjCfAMQXma
J95WPpdEPiOX9tnFPkZ58mD9PruOVPa3Eq2YXaNCjxn/rZWJXDgF036o62tHwk2oN5WurjiAEUB4
A9cCrJwNfIaikekoWWLnSrF19/S8/v9lGIj9WP4FjrXYof6vtDGoCoGiPoRFL4UejxtXMMFueFZw
2qUMHc0n+EtSF0zYHsjWvNRS7yXUyRoBSw873kKKUXimQhfWuF+Q7JOyVGrtrp3ExjCwlRg15kTp
cAATjwTLIY/wUc93Q+9I4UxX60JdaB+BKRQpz+PyTy1LGZovPY7MpO/4zWpweEYx0bsN//owGbuv
Hsv7JfB5x/3TL/upqLTqW6egsPR0v3Xtdh5l8pTAVGp0bOqRhZho8VOPcmy5RRLZGXvaq8bnvpnp
5///kgxb8DBiji1NI8wAbcM0U4f2ZwBlF93Egf0O3w6hUPnNk1eFYBcbyKQFvcueauKgE0QjA8gx
ur/xp1D4EjMyAO6eUPbTu7gUm2zP0/qUXStz+ddZOqCqdt6SnuRxRmkOlBiPiqrEhGsRvQAPnB9/
KMMmthFxDhSi7/Xr1QrGiJHoDA7aNtEpo4jb75xkwg1v+cZ2XA3orKw8r0Mc2nVWvPDrL/8zbAnZ
Da4yr08Quk7x26blLw6fz7Oh5mE2tIAjLQLWBPKlgZmqZUyK6mfVrBqPVIM37/w+8swNK3meNQuf
BXvYdwD7ORcaZ0f8EMDXrvkEG3ZOYA9ykcn8944EoV4V71yY5toGlPmFF1c8d3A5Zmfd2qZLUngz
wNw7YzBawoy6eiMLNbtmVJ9oUzZgfaSPRdqpzXeeyZl37QkUgJ+gHA/pis16DtXG9H30BK+BTQFa
Lo3j2HhMtj4fwmgQMd6yymG8g+gdcw39Up7lpnB003xqMMhMl4QboPq4P+Dh6qfQLXoXXi6ZGlyP
EH9pmKEmwRpp2X11xpURnGcUEbfw7XlRGNDklWNBQVOg/F1H6L9T4Y0aziJiDZdHWrb7yKaOiZuG
+vZGzOKxu95hUH/jZKowylWUU4SeWyy7yiZH5QL/OYqrXYLXAO4pWZTdlQreiu3dL7t+81nt+IJn
OyI2AYUOcf66+ijEwyZwUzK309+H0Ed+dM89wc2bJ9LZEG7vAyPKSdxaPvNdC3lT9nMzdya2XCAY
UnQVw66UUcqPdbta89w2fXvLhLXL7i8a9ogVUj+92EoUHNM3eiDUWf2coNECg6ewDiiJxhh/LHw4
DjURc4vIkjA2RBuFtXRno7ucsUEEorcJi7/MWHmu2V7MBXQeIDndvdnEKmPQizHHv3ysXtryIwz1
YvjZdH8W0m/8YzSMdq3C6WlBmi2lBrdPElDd5uFHK7qoONPH+R45brZyspQ9zEPJ7lIVPQzpNp27
eTVUAoPe5SumcY/qaqCsZt4IKPpICu6pCvuAzQokNQHHO/zXCBQNIkf7foru8K9f27JnkhTn8N19
SRvTRqFth4Tv3ZmZF5R0kpEPnSBq4hddU/j+xaunG0iMzY2NcCmYDLqi9hYJ7VcstNANPMX0hg2Y
DjR3EPAxka1BSTPBAVzD6wYocLxGAtnJolYPf181klkZ5/FNLsg6lcVsPf01jzVpEVSPD3DJ3Dj7
0uToaSXkeONhdLYvkOpqywpDxK80cqqNF3ayMruKoU+Qil1D76l34gRxczTziPOgIhXYhOb7xifR
X5bWSy7aIywc5EC0oLYzMDPt2szvXDTakFyd2qOkbkcuQRHwbR6HNTNEmWO6s6C5cp5ClM8NmxEO
bxSMmMDKs3Wt4efud+1ygam7JudoRkhTDkZrO1nW7KuxP7gtUMDzxr8rNQBNFyOwvlcaR4l5yWSt
OTmvOjdRbbdPzlyDhU4119nISJWDAXt3nEibUNTJZinJ4gsIkzbtxQGMyfRnJ79sDinW3AlHgNJx
Q8BFl9Rt0e4BnyinRHKMyqgTzobBGgXHW85QaRMeMWMUEcKCqV0VgKA81fyyzWUcuQEVm3lerU/9
GQTWGbcB7OLlmfUIo0WmraSfreoFzDuP/kcJVoVjxpYNHISXFUGTDngYQXmU3ISus9WApp30CbYh
eewLcXK3N5O9yrH6oz+xYtHoAdWy4mBDSt2QN/TeN6Hcj6eaSwAbPQi4mr4jHMzOEewzerskqZqa
jC0I4V19iV+g9OW3JNhLfM8yHZQFH4F34yuDV73jnydTnStO8OCyEK1oqdgWarJYukX3JX13B0w5
EabB1rOUNucb5IhsXpn5eC3if07c2U4YpCzpBMe/P2RwKGIh2J1w6TGw48OcUnh68TWelzHCWYkg
zLoFVee/g9353atqdn0axSp3Ei7/CelgxpVXDrgoyOJauJxuFLQ2BgTL404lOOubgczDLvB0ySbX
o6h6ErRUdh5yFOGImg0TLDoO/0Bc3KzimgOWZhyrO3iyC4V9zU8JWead7iKq7V6skFRnE+P4XCrg
DVZRCK0nuOR6FRK8YyTi5FrzfJfAYwTtNtDYmY5gVRCj74jq+T9SfUwwJYdIZHovdZLhJxwQxOeu
vSBdYIFS0OtolNNjenRg/uhtsuOIM96oMl4VW4lj7ZE8/X5EEoGuSYK8GHRyiBswOxURVZOtOhpo
+I+/UfjzfQ+YUJ/cfolHB+kHqXVrgmZSOGjEmQ+an1lg3/pt+52qIvojDMDe9xNxELfZ8AV2AXqK
p8taAop2O7IUecish/0Lp14Xdm5NTcDoCW12TTNM4sLbKlatHkUC0UsQC+kEDY++AzSyf9IjMrZb
EOnzuozK20RYcl20BmVdaDqN8AFCw0AH2KT2rVd2yiNHs4sYSkqiJYGwFI/oYoobQy+hX3n/WNK0
SrDnPalDecM7kyNMRTM8I9Yqvkn3yp97WelZkHBGuaicfiKWgwsEs+SqJw/oY/1tacB3GrJjjLue
++CGVCIc8M74UI/tGe+LXS/NOOLOpkrcDgm52LGLuf6a3p0sZ2f3Cy6bHRZcnh67hHfUOLEX8kSt
Ecyqd57ikZM3M+jOTaBEye6bGtN7m/vmhcw4ynDNWSZgQ9FCVyumvMEf6wmpNuBuCztPM+N4lGjK
+UORmR6NbfotF6W/Y1CowGd6NjWmM/mEJLecTLTQY6nzGLNAHY7fBYgT4cgF60vyqlZoB6vA0Fi8
Nq2iZpvXRj7RSNA5+fllBPVmydnlq+SI55A7OrXRKJMNjQ1+myk4IVs9BjqAfyOmtOVs64TSYt5/
pYLKiDoFuDWN4tQIDPDJHV9tT0Ls+dVM4dv0alMXQZ8v9MAt7kDImu7eRpaqsEQfsqPOjOvlZLlL
7EMkXwUbkNl0FG2rJFAbrUfGbqR8wDHlrRPP32UtvL8eNRQVpAxAbV9WNh6qjXFYCQLe73RQujk7
WIZtdNtpdz69UQNg7cfC49VfEH0UaufIJcytMFmzTYByHt0QxSZKXQvcC+uWb+qzMjkoHhFbaSa8
a56IoOhFmkrKXo4S7SuwNys6Pub5Fu9RRotISqTQ/xWpIV7AmfLS1o+Sm9RHS6mg3G+fSbGhxw1F
GKxqXEEpH1kCaEwNvv9E+ihUEzcniIRKKYZ+mbZrHmg/fNhDmkw3SIuTAD2HERVO5GPU3ACF/ki/
PGurYmWaItCOP2estiVZBt31GGsvoHuFB9sF0Q84Yzk/fK3nw/Arf0Bjsd3W0n8A43qEsPIxTadX
JlZYebSkPcfHEInUzHOsPCDnHW9fFCVsTfFjNGD4fROFK6weDfbWTSzt2XufPgOGgYedU26Tecz1
U93aTub0TnT5V4Aj7h/vvuO/1cbrI8ShvgEfruIla71ObhnEVVuEvnDCkdkFGZC3NWLQ5EUk6yi6
Uf10/TjrzlvrCGLnbeIF94XDrOpnl0/NG2SRt3LtZNnCXyl32iCBmo34HpGGJ5WytBD2X/bxnK7K
LBrntMxAc7kFTmB4RxVC1GPKmMVVMbkIg2Ri4b+DCrtg0PmTmFz6EhHtyfCHtm4/LrqjfE7hi4Ni
KkLzjdh5azfYAhzbd/U5Fn9OSSTLdtPSWzIZ27vDZpAP9F8tRxKJ4mNg8NnVA9KH/mUsbmc7Dkvn
YlkTJwpq8HJqfQ8EXxMSwu/BI2+I7Pua8p3n0ranKNYvSKfQgMsGq2r3Zejj8cjwScC4t2ewK68b
JPYioFPf4VsX3PrHhUcW6jvHDjjbxENrXvLoOIG81DXAWXVwRmnF/1QMKMUJX/yOeaDzOZFEax0T
3PQqlHn9RFqI+mI7WHbtlwnGB7KYgfgbAep//iNQuTZfLh4GA420IVWmcNVB9fvp/HYyDkp4WmTi
O7nY7VfS3gXOvePhs/4d/KvcYMgKUkrYML8disMMpZLgTvxyRDm96IKsXnEMVv3kvY3/C1a0DDJi
4muBGwI1XwThZKQ/CrPYDMUnitsdic4xbj/nGyNYVNjrMHvGMunixXItRQmif4deTXCLLMNt5da1
9vxLr97qufFp3EgNVSDOwu+nVJi8CFPASAxQDY5aEzzh9Eia1gCS8VZ1/nMCxAOWe+aqraa6FkZt
h5U3SCV5M0iylCQWFTG0pjKSjB/wHqu3njJhAC7AuKxFUAhpqIyHfgMPcq65Zflf9chDu8UjbZux
24nfIqu87RTsfy1joxBSqIUJbMrIJldK2MTjXOlWMyD32TTFJakqy0Zh0DTZpOPkaYK5xkAsmspW
bx2Uv3o0Ns+z1pQuk481K3dSGHUG2NuYRl2tXBlZ6vgWWNVscK+5zfpcSIf/1P4UY38/ILPF6z1P
Sd/NQAwz4mUQe0Bdfa7VssK6HN6IKndy84XVO1dU3Nw4+LR1i2SyOwByCtHLQS0s1h2Dpil88yIQ
CP2L0Ak9UVwxztXegNGRlTTfCHmjnDkX6eUC00pibrfhVNimqQj1Ykaizs2Ptu524uJtYkU8RJRR
q9BCoGErbe8HDfc3WS96Fy2epRrPEfLCHooyGZldj53zb2TVVMRuXGyEdsoHxRWZhLzUQm83UZO0
WdGgG1Edx9t2vavK6Oj26+DfenQWkRC0LeRIp+gVDPll6/t+mIf8vg8lPKLop5XVsnjDMDpEPEvD
QmnUVJaORWGByYXn0xqvVsLq1Tc1FgWH5gy1d+nwb91PEygtYiK0rBnyEKlLrSh01KqJdMpqHBwt
Psz8vwcCyJcb8nfIwETXQhfsznOkLRr3vpr5hzvSX/pN5DZM3OmAVATQMhtxAgRCJ3qOLCitoVsh
AlADmd7RBW43ONQ8rZ/jIe0OKytMpQPtNJoeG7lQ5rbbPWdPmWF4ApjqQdDLl9CXXeu/dSP4Qy4c
vqG0u8CXEhmamXFL9g67buSFtx3t/odYfelsdDBSxyVlM5Xt2ZYpR6pVn98PqgKNx1RJoJlxcZ+C
gOygJHnjJ5HnyWV784Fw0Gy+VHhcsCD6+JL/xatuMKlagENyH6FW1zQC1u7+0eQSrbZqxmDyhPTX
L9iSdPNtn4+1VCOmrOkE/hvBRNsJThGl2ny+LDZF8KVWXVC3aa+p26RLIbA09Xu4j0JCcTfir6B0
Tf0TsHGYVTInQ4mitoDGc5GUbmWsQgM3FpLm0xMnpBake/5qo1XbrbYX7/IU2e5axaD8letJuOj+
GVCUhWj69j+wd2kalGNRcTQAsAsOgPnNF4Ecd16357xIkoGsqT1bWlr3pHBbGVpSxDz3bUWdNqC9
2zHmyXv5wpjOfR7f89zTCWZDBfls/A3t/o8zKSYtPQ+s+DqqZ8CD0TX8DnFDqj06jw/lX6T3OIOz
LHNNdJq67yvUD2fstz/vbh57oQ6dSMiLStvz1nZCxpyFevE/AxeIWveEqW97l5/owLIy1X9wFgLn
zCCaraYG0RN5q11t1l97NqgNyIAkDZ66r14EpZCAwWIf7zMnPNYKLlSU3ZLcjA+IdWF2yU2xwBb3
tpWUW0GB1zr953avAP1+B2NK1yeT2mrjmK5TGa4nOUSYOVbZ7elW8+z16cx69cYNtDye7EPmabzf
JUEfykw0EBPls7W9omIhQ0Xq5j3zgZDEx5hfeBdWM15yYLQZW3EoKN3ETbAWERdIhd3JQnJuzUXi
ZExramkEY4DDPi6fbc41Vg+zIv8MI7MhPnsrFBTf9B1N56L0pgshx9TY+1kG/CDP1n/ef4B8mV6Q
OnYqX4U38FqacHFCDRlYVhoK2HVQNtXvo6ZBSekCxNOkk6R+Se8gR9WokQ+RE1TknhPnD7KQDx9y
cG703qa5S0UlLF//p1JNqLdDpl51xhfR/uYdIkPKWbwq92DrjajdXKo9iWpwx+aESxTq0OpNNvLb
b+2hjxn8UDrX+gs8kV28Sc1O39/ummX1lbf62EK/UTL2U4ZggTO/DQmMDCl4Dla7CgfKohzicPP2
vuyhpug2LAv2tqsgNZrV6+xMP1oHN017I1oUQh/QNAWZ9qHDyDPKRs00ZYuoiMI4YGph1rsPoi5u
CaeTffDLX6cgKDAi/UD2VuoSxEqRvzbcgoQkbXsBXTSFuWVYocbvqUA3Ziu5/M1TVV8wwC8kzeS2
1agzjSnpzZiuqtMNoUQRlmCnMq+IRyNwFtdvKsL5Ar/CmUiqONvX/b9kmhtOEUBdTdLWtGJaMe1z
gF1/82e9huHQHs6y9rM98zEh3hVYNGfEYk/PrH4mS65xkAvZcZm+RjDzyN24OeOB/Mxo8JouxUc2
L9edbZGMvkaGxmJLR7Ux53WlwrHuBBJguT+vujEz4FlO5VsMWYSTvxuggVuwTNdWD6PGmfxTA88r
CaKFZlgfb6r5KmACSdCPN59qe0l/5ZUdPB3YT6UdXc8tWZRIofxy8+2KBGMxX0t3DMgjvTBOo9ZM
LTHr9oB7saOpr8jlgN0WrobF0M/onrKwmCOW18K3jjaRZzcvUAB4/kSLxacYMMlvEEPyS5p381Uj
zHDhcvpe59WUWbZFm/68QmRdisS1VhHNguQY0FdDkw2dDOgi+saOMKJnmdBS7Ci+KJGM8Zgjx4+g
ozQih9WzVCLb1CN3ybyJ8hVBJSk+5wnxFWFxSFNJ/bDnmxyi98AymMg1irpQleWvDlcUzcJLaY9L
cvUeAmp4yIyaXpFpOeKZR+6oBOQ2dBElkv0v0rqVBuBqsU+QT1J/0FDMT1TnOX3vxpFXrSkWagp8
6EQAavpk+fotUXljOPCJYC2QUSfXE6HPKjuK0nLCxS4ppqVmqUcl/kO6srv0Npw1WNlkYEgL6M2Z
Lz+RoILUJx6JixcDyVpgg2RHUoBb8UWYyqNmlMJZOV0/OgT8o8HuUGgCilkqTGn1QORSIkHSdA2p
M8yBexkSEgCMZn62t+HhLUoS74YBtPXdjCb+yIOuUZ3GdAryIzXE/ux4ZA/u94K3ViHPdtWhgFxy
fam+xY1fgxmxFOHJ26HqsDsa6+oypQ9AKYeVRaY17zxnddNYwUrHRnwDWwmWVu7pyBnUgQYEieJD
goXiUHb1/3nMozaD4QoLx8dgHxKKxgr0Ru+J/NdyCEVmt0JvAnvGno+rkqtOYcrqq+byUh60ko16
sOgYMYyfNKX5Rikr4ZKoG4sXGczxyWo/+WDreUQgnIZRE6Jo41tgeYFs5vxZGTLyIKl7phK61S4x
wRLywpuPX57VEbyNZK3l2UxC7b+iBMbcoVxVLDdzVTzgZMo+J+fCAPvPl25/nXcaK8XnJJWNR1rC
gaf38uhhj4J8Iz7Qh5u6qxpBC+fPpOXq+I+TgiWlcRFYkJS9DjVxnk6o+s4DtYYuKmT1sus/9glu
8jgnoGKpW2FBzqdhOF75YzcNonsskEhmuNMP3M+OB+AEF/uGGGwe3kelfoeLfarE4JF6K3WyrCDJ
1FaEhE5r5uUFUHdSkWFIcg98AbH3Ele1YLvO8riw4SlYrFZ8FlouXQkS4YKKe81YzwA6gSTL4IBi
kmd37c09X1ThRehDqpv301e3jS76B2RJV6jRjQ/uieazZU958SvdOdHSEtJsGyvUUJKFHo9/kRBR
D/jHQkTchnqGPB/HSmrdxIqO314vNN538T9GHSnIQAwmBEc1BZMKWLc5es2ztNTfaiAxuFDN5eE+
eFTQgn/zK6rFWy36bMwesHtK/P1YlVCGPHyStlWvqUlPNePBGEqbWPouiW1Cs+HRVRnYGdpV9Hej
CLqEa1T5YxFlGSXL4ox7Meh1zJJbJADHOaKBsFXta1mamQQvqDXD9yWd7dAjULepfZAWKyzeLbky
KGYvulbthJfHCZpZ+T6EzNlIHUHu79GXv9jh6v849iPO2bqQu8/0WtVftLzSwGoyaKNWeVjHrM7p
X4oS+ebzd7RyQ8QCgwwX2rubo88Q31lsMtHCGI0rYBF8bDdiTKVKzwuSfQnPK3ll4QoHGP7AIA25
H6jDhNqG65uyg5Pt8kk8+cYYkOvoazZs6o3zbiD/9NOsEXkz1D8W9aiP8ymc3BK4suOhwOf/R4Oa
UZoCt4/FpaH5nsL9RzQeCJze1F6SUtfjaoqlo5W8DU/MMM7k3w/7igcZ+RHi+v+Q7MgixUCBhC8K
ao2PzVOkxXN21IQT23S0LT2S8jXedLZYqOIWX60HwwalEN8WhOF1J6o1Z9G62Y5oDNuEbwR6IrpR
rBxxR9zwF54gOlKJJSFsXhoSKFmKmmhtG06cfiJif9HfoGYciDFONYdaKDFjfiDdKDltTSKbXKyH
kcgmjbcQ20qoSCLDCWo+RK+CkUPc06Xo9FKPxALh4KjkvoPbzFSrki2qzEwvlgcQeZ7wORHLozmZ
83PRoq0brY7YwlQe7UDmlMucri25/uBCLZcsXwV4CmOMLjs1E5yePvQrBpP6q4Nfvt7JzrnTXv3l
UqZJgpipE9sqmf7YMvOhe4xPUMyZQvT/qvjEL2QqLq1OTFocCalPcAq5ANYDq2BGIBYzV5v761iI
XM0sggY6dIpjxt6kD8xwHY3QI5FWgmjYxWVYJNHVMNwtoq23AGIyQg2Wgakm+B6NEoGTbIni3HiN
8CuO1wAJYPSgzf7Ua2LGrq7p7RlkwmxrovbZ+51u172FOh/t7gW5D7haQ0tfy+6YMfAPg592iR7p
TiPlxNybPOt+JC2NQ8p8aMkf1hgOIJAjcXwgEENnA59XdtCulYwb7fblrUmnB1KQ7bvu1Bzqi9WL
UTFQBxli/9KLDb+B7UODIl9u7shZ+P3TPiL4enIaWwoOtoSEA6rOITBspWsvfDL/OVLYDdf1QnOP
Rq0Oip0rZpGv9tih84SL0dfRsL5Tn/P9GI5lid71ujRcYPAUSdLZ1xcQhwvhhk+iBK4a8/J5/GBY
0dQkvOMORHs798YzHaIR9iDQkbJs2dpjKMhRv7xhG4ZbAM1C4lOP1nRe+H8m/6treONDdQLC7OHL
ty6wJHLORtjZbiDDA+JXwTvU/suCQ/mYbu7hScmca32nAvlipXgcyZ4G3+OERB2QMkjol1EHJe/z
Ym7nuqJHvjvBYc6ieDrjRF6zgyfuLk/UZ3+8SpXaVxvrt5RS7USQCBFbp4ZJ8AsxgIRSh9Zvv+Ka
geTxeAqzRG0bYvJEA3B8bjTeIniSLLPy0uMVOcGglTL9WLcAGORw08L041LzgrXfwyD49G0StyM/
6viL7oIdnnOMg39/f3No/TyCaL76vB/nbtPrLMewpl9sk0dPKuyamgRCGEUevVbhYwnzPq+Jfedh
vlPw5cgdVlpINtHF9VH45LnsRi7Wpfu9FisodAK89e0C3pxIWQkgrVi4KZQ1vpzAJ0NN5c8NAWk9
/19LyCPTqhC9CIgOzVRmWrlNE+pN/BUJGfAq/AP41M0+HhiQCZmpMi0lqSA323WsIHPFLP1VGpdQ
CRoU6PM2BD0Yf5mUK5i0ETP0RPa3/iECVIeF/iayL64ar4vEd7+s82A9+w3GfKudE57Eq4KBMMV4
Fu6MF8+ckGLsT8jKOq0ClokoDBhxoke+TLxd6UD/KPUBkfAt4nSco3VnXRFNE50cX1KiKYOInDae
MHmmtUKQvjNssHe1iNHkN7A78K6Bsw/ARaQdJFrD2rVFPw0SpCT8cCKXhHRuC8WhdQGYXNlEc2LX
PYNQT/EFgn3T/faP+MIcRKsk1ZtCvchughyBvRSJtuvHKRgPys0B3nSCTqcWa4RrGityrJXhRec3
4AeHf+CoDtoIKJoCmj3J3AyEKvNqIeSglYuyqxb6QQQux7fzoWZnsI92KBG/dp5C4HLAPwOgRJ8H
bIidrABwON8hTGbymXPVbKvn9JO1N2/6K4gP5x6syxD5Kbuh9z1V4LImHCC3FiXxHNJ/WH9gsnN+
N9i5ZlXAlGsHXKZLFZBpKozwlGujGnBsGN6TUM7gx+4zR2NrogZnFF4M42kRVKxi3/kYY7HamxzQ
ZcHd9HoWQXA7OxRfIGYtvUc59E2uRmUHMDom3DOGTq0+tx3d9b9jJZMSSxeXONfli0JdL3xsfz6F
YF+DQqMe7smSp95dxQcug+qX8XnZOamqeNUw+WkkunnkIDMUnGXyyb84LA3lbwxRbhPkvKz91Wv8
hUXAW1pqM+jyejgesV1DFt/W1OPUP5MtbdeOFM/6o0ge4aUfbc2dW3j+8/9ofQfYcDXj3EtOvw9J
x4XNsESjCAxCALka/bM/v8z3lNJSbEpo//Ee0RSzNVrANHvNYDGXwSfDnSXSLchQWyKo3aMQWfxp
GaHbBlJCYRGti4fB5c3WCmGSKcAUN0kA9/3h7INLcz25I9SkZx8gY1qatPHvpfVUibg477NPUa1h
4dSMN7tcmiN3pMDOH04XdDazmO+IDki2k3ewurWMfFHX0iC63w6lNrD2QpdgzR1fU42RvcB+J/k2
xtnjB+kD5pN7y46RH/sIOjsO3IQq+U3Esxe7Bz86eOi0nTZ3SFXesGir0ym6ulpC9CQf6vo7O9+t
zSv5S4m6JLs4yOqByoulpC4KFAoiyRIVshTvFG77h9L8MB8OGTIDj9mNRCIZKaIPCaILjZAZDg3x
drv4RL8r3NzyZL1VXxowDts7l2w0bsox7U6So0OCOlNywrIX56HGTLoCzMqwH0Cvr4Wl+zZJuz+H
ch3fTfghRrKzCp/8VKDLEuK9kYh+tO7dxn3f0bc9XU5pBJNNOievLFHjIbMKMZlQ17/gaxa/a8vW
qmhmRSRoR9Cz60FINgsYTUku7U5OcREjBHD0pcEdqwbWbGxh1qUy/ujCZhI9q/0S8oy/eLyV/9Gm
qVJlD6h1EfOQ8Fsv109kBTfH6H/QJPtZumVFj6Vo1HTnWJqayFa3AV4g87P3jY6aOw9r/RTsPKpA
JOIWBqHrDM6pGvTXGB6s0TPT5QKcSeGBDal6p19XFCVcAspRykMadMjFv/ulDlxeR4AF5DzDy/n2
e/I5ECuLSQO00+gmtOLy5ddh5H0wZsRca8wKl+O8yjJy2p5UaEReEBT+gkNhekvDlOa3cmtgTw9I
EvzpkUdCS15/8yHfPQIPagSz0FO/uwQxpNrhn5Wqrd5JqYsZEFXm5dKawfCKygo7Tebb1ULzumSL
X33Y/+JxH/ssuIxaetgsGFPLPWDf+5AlmL6DflKnPhuBFxI5/ZpauZFVia8dAADvJVcO/Hf+6G1i
uqVdFhSGrAJVVvzsJU9bWEgeVDpcmHuSaU8GfGxMnyepjqNRte3ax/PWwftZnkgrG4ZJO+gsAvjV
qvNQKAQMkLVEY5BxPvshYoi1wK8hrHY7VsIicVkLVE0BYO6YL9iQ9kxQRtWmeEAmrOJ0iDT5wTc9
dxymqdOU8pkKlOdEo0C9RD7MowSrlYeaDmacjYkXgvmFAe2y4iROnjkSqyoNPNMsJmnSByk+f4g0
7yeBd61lXgCqCXkqo/tE2Wm/aJJsfsDzO2jODm2GK49OAg3vi/2DuKxRg3X1X7oRdvR40/XfsBwJ
OPa/nO92NcwzFFK7rhbpAT45aXLOTdd/u1/mkfWdGkbL6cGzOnZASizgC1rW+u1ZUTVcs5pxwXLp
wIViLw3UYPa8DqVFttH6Tk3ViI+GqNdhZpt7eY7kmf2DNBoOmJ47o1FHnlTOn2ffeZYz1naiZ890
a25+2sKN7SyAzO25ZIR8k1ima8RyLRMufPTVoCbhS6sIc4CHsbhIVzbTspPWjFYhIIiLP9uI5CPg
9pB8ZWVkRojNNPiSIP9aFhnfLvVdKLtlWWhnDcne+Iizfc9lcPqFq2VOZEOH/mCqzIpPOihQjpmh
SkgmiSlbYM1uU8E0oUbC8ZkGi84hbxr3XZGlX9fnvpCKLE1un0Mg9N+gp/mUZpQ6LZQqFxy0iMeu
6SJbWxXnCVxoBR3OOuTksOiNSOfhJ49DmYbfagqFwY27nb2Z1KNm/X2r2dmyhI8XlO7UcggTTmjv
6L7lAhedRQNUbOySlHWjAZ+ov+ES2Lvj/DSs+jh61JTUR7QBlY9J8q/Glfj5VS6hPiMt45NBdX4N
xdm6Cy0o1ioA9kutJlFOs6Oq7niSd6An2hjm99i2XsDw+TK2HULnDpM9K+cNCex2rUMGeLMFG+9L
U3uI1qCq6pvmFURmXPizzEJiLFj38KATknh7RXn2/M7xjMjdFTPU1WVtwGhAwWKJk7DuOPwFEyrq
O3cAzWfXLOLlPgU1ixboV6T2eEsOIapl2gy9nWLwhSPndNk2RCp36YxWsMunukZ1SO4PNiR93VD3
0wCvtzqU6P4kcxdiFYbdnHsoj3iDHcyB2oZscIrKLqMq+jPssnEYU8TpvOQmQvh37aVMjfuuathV
I7+z64T6aUSd1sXdwyuXTCq7DX20IjUWL3iE5VCvgvCn3t/MxNUwkFRzSPtvUuv7XSrRo5pMe0qf
7ywaqejaMPjUVLJxAtfrAjQu2h704dPnxpFf2xjLfRqtLMbHFXzf1/GdldDqNXVdRXf6oNGLYPyR
dp+pDZSzw7ycTZkmbyZo9Umxx8QlPOWb4cDfXVE5zRjBpfihjUhaqKl4BqrXKiK99lbGsUKW6gZV
NYY0uxrdMjV1vn0qrA7OrzUFX53BnVJLADOBHMd/ilQ0WgBlHe21hpLxYXAw8nnFLTKM9wSoQ8ox
mnT+e6PoP6XPmIraFUHFezLfTbo8f+DcVemIzLz76GErrPAWay2Cl+Z1XXI1p1W0tmRc7cCT4GJ2
TDyDA3MMgxapVGs0PmjYxAjM6CHQqasfMLRHXSJ09NrFSBoT5zyPbMTpR6V2fhPlVXAvgZm/y7M7
ow5yTZOxOwLLAe5PsbGqkAaWJv11U4FlBZP9fZL8sbcddzlt8v7xaHJ96lKXXAUL0k/Uy+4sQDm7
BlymM8J0ql1yJgjTtleAJGVqxVOmElGmpoZ2x5RA/NS9AHSWz6VsiKvJwKVlIOpw/yAyh89znOzb
+R8OohPhQfZL7wkfgp/5drAkyCgXQ8kUeJHqEY5PYxIufrXGo7BVMg1xTwS/5jMmHOFAUOUAysOX
nJfw7nBxbaC6nrYZQ//UOt8HxngUT2MPpG/kaCDxNbdKgVun5CPD5rhT4ev/kdQwMa7qVbT9dEVJ
TEUbWB+n40LnMs5haeNI/9z3LaQjs1IzLlyxmfWS97louMAZFqVFgpj3AU6akByY82kcyWw8l1Wq
SlLDJhphz2uCJdHQAqlvUakkSytLjGk7Ndf3qsdSoUXjhQlsNGbUy7qljp/6JSMri+PBJxGgOqiV
GkwmMYwswMrOFxPz0ms7wi76SIK/EayIvsidmHHCw5zJPssQNGounxH82y0wmbr927gYfJ+cwm0j
CV8rQBhZ+Q/0Xk/pM8Rzq/r5UhdsTqiM/b7tDsFAktOZT5CNgPBzeA8MtFlG4m8sV4bvR3F6dibX
Onz+jeHK+2bhYfRhneuIoypnDUhwsgHrPuefg8n5QBVFsBT/RSQaG01oi/9FUyNDfA/8dpK4X/iS
vwiXg6iGZQ5ApppVYJbGZ3Xpt1Wte8UvajCuzbUldEDvjoq9wX5zvMV5iu8INAppW1ASdPz5jXcj
AgmVeTtmqHGhRXbFSfrVhDnS+/LoLPJh7rujzPkpM4v6EraK81ILoAE9AH47zzulU5NXGPfOLhM+
cbUyGah9DcRc2RCMa6GwFkCMmqBSZv2IBMY0zUVeGvHfHkmyyDmatDXdINQBvWepkWeDbqqktScy
UWaxOVppfVtotQ15MCmfInIygc+L8PjlYCivUX8VeUbj8t38LxXFqEytCVIyotnlEynDB0JHdLO4
BvX7y+9qFeqxyoeEB1lHlEFnB7mWin0/FxV0IleuvrXjcFkiyo1fM2IbHZiaMYkYieLj+4KkUs9b
Gb4+xLpXKV5uhtUr0VNddlvZyuIiaAtj+G+57h3K9L4XtYUTJeGDz0bxij0PD0eXirNeWQHmvr6E
v7RzcFO6P89ohprk1MEs+l5Xv4UEibv+aMkreJcdNKOuBB9JlRLi2UD+U5kKo/tihbT+roftxc/N
D4sOgTrfqLLCbRhD4eCUjEyInz2Nu207DI3g1aX5ndu1a5xgHFXBOMkDvEWKzwhsVlSA3mWO2tti
evP+kfVFh9dty15/nEG0VrJ16cpFYagHYP6P+cEtqmktKRB2mT2AeXViTBMajacHAkCjMO5FnZdq
DYkNw3IjdLpA8B9q8eQx8C+w0DWysKMjJ7URDIiiKlXcHYVy7PfZVfjRJnLnIc2Cev3XQtLFrr3t
kxP3iqa10/t/LWOpT+Q14mDrM4nL4xoz3KbqTDhmbNHRVysb/6zAE++BtH4N/sUM4nRx59MzemES
WdGgipc3XaMD0V1pGjJCXTil4Bh8nUy6HfE8azGUaek3RW0GoV9sKvc9ybcEAl+naDDnvnabTtUO
krr7D5pCir9clP6GW7zwVh7mwY2wg/1VotABZQCyTRTjSo/AcsGThoXYiFj47p16l0zhP3qIh9dx
YMdbmS3hueKTLpIFX2s5Q7akDoNXcrfwPAn1C3XB5RmWVy8343k8dUmW7dPC33RbOCo0R9+/goTB
Gsyxi1oHv3Sh/k9CjhovHzbJgn79qrbRZLo0wCJLQYrRh7+T5QY7ZGAOGtfLbW6zTdte6tmo/ZwF
RiCuNg+GUFGmCBo/ouE2Mbxa96WyiBTGFbCq3qsidlEQUSm/8WNvBU/qe69tDAPS212SeercL8gx
3JQRMg5Lm1hJD+g8aiPaX14jsZbg+KTQgiBBZNnHYTGAD0DptSjVIdyZEw5eAz2auBRosnBcsi/m
5Z3mQuJbjyd0UtOZNthukbF/vLX7S/273sLGVIBkSAGIU08mMQZa9SXmbUg4vUFc45VB1bgZxDpT
iiyc9QSkXcGkiIeLsCqkOdUUrGDEZy+4/+9lydyV9SZda7MY4wVO5T/UffqYiQKHTG7naFFNKwFm
8NGZ2Ohpttofyn64v7hrG1GZBkDFfcTQNmjYWtcbYT9wphXJgTp3+FDIs7N6ptIjXwjo++qRUoqb
u20mSeMp2H31WNLkg0ZYUU+ub0u1VaG6Ho65bHj6R52sfKcJVRFrI4YBLz8MSmm7C/69P32epfMF
W+1iKK83QlIDRo2mC/f+CsBO6/ZXAGta1/I9DibPHi8IvwIfaKh5bsxMVK8uHyI/LBw2lortKOB0
MUUDi2VuWjZrofS7A4Cc9dEGkWVXlPsQnwXuoR6fIHEJA2KKzb+BGswpSG7X8ptFoTZkFKuDO0Bc
OaH4tlwYZ91FCINcwG3xnPksg9m7T8qpx40B+QbwVNNvDGp6qfarO2ejKxr5NShE+X74R+pP5nWW
ZCh0wxw4AAiSr2DSVkLSTKqLUij1kHU0nK/MZfYSkvuuUslUUbPJvnlENiCaOPLRzFrOMbiCo0q/
Tk8eXuFdufxwDmKg1oBr27QcQc08WdJtWQ1Y0EVe5CtxaKyd6xNcZR9iS7Tn6u2gKtD9O229ufWw
SL3aMDCh+XrMnFzMm6acJiV1u2KGTslKcVfYXJcB7e0tPIw+XcjqQ/6p40nbcYHC2d95odjVR+ZY
KTzcHVAluWfJr40EdK1IVXoCF5+JNkOvgfZ6SBH+nscw/hf09V/0LBDv2BzmcUivb/hFYHrcwypJ
5q9SRgFSBxQ5UFEn6cQMuDt33elYmS3O8kLKDYHj3gzpRuoFebt7Nk8b2t5DlIlCmDdW3ki1dUDL
GG+Saxv38+C8qP5k+q+z+NIeFAEfinPS/66RPuqeLoIEaRjVQQcBJTP81OluKy9YtC1W0LRwMO3s
wrywGX5DYCj0Z6rZC/vxMTWaMKXzwnbP/rFIcJd7PK1+d8JQi65A38XprU74+e/Z1wGjj9nodxpT
adGHQGpsm8KCFt0uCw2qS9Chajx6fX4BCk+QeQJiF+N+Iqed3B754gjVsQoAQgwZYHz3qaT6Xqfx
DhrcDiz6Ys+AXnsMq+rb7VnDR+ZvKpAKg//mJ7v++vKmXWWRO6Lls1oi15br+6k0qyefS9O1UvXg
Bknyy3ya3kmBfw/Zxo2RtfObYvc1IznqTeyAWsoNU9tY0H+uaUoV9oZg0vuO0C7OrG/dkYMezvzf
c4Ol9vDtZZZtek0RhwBBvmGwKv9glRRn0u2pLDKM37bHWHzYV3+fkUJC+ShTLzGpukK4IkeAYHXQ
ko7CnR7DUE0nNaHbUFz4tL8FIJckdUHWQ0UsPybgHg6aB2f9yrK99bXCiF+7miCLXkzdigt2JsXr
VB5EGV+K2+RvKNjmQrQbvYoaGYrM2OBtb755s08dI2CcgPZF1yuS3L1xgJ+x3yMv2amK0YE0NTwf
21HqZ7IiAStqrP/ZTsxUhhONSr3zansRfsM3NK/LuTDdM7gDvKuH4wIIyiSv5Gqaz0elO56Nhj3L
CmZhy1n36LxQhzzKND7qi7cbS9yl6R/Q3h/UqLPwwlEu2BDvfMjoNLDu9VXzFoGSBj+T/zAEkwSZ
9qZplKcR0TZRpqU3xIuwDAB7yTbAWHyJCbFQp5Oj41QpTLunswf8tuJy0Z9oXe7Bgxf7nWw0DsFt
svktXd3goPEk9PxCBmR69b+txDENesgHQtP9qwnuo2RzoniUVRgmbhEBnWLJ+HRKq2K34PhT+rP9
XFIdGdHr5JT6kk5FnzmtEPypzg7wFf86bsZ19dYvgrr3VmH19RxRrHMvktd+VQBGiSiAksv7czJH
OwHn1b0y+2IzVzVks8kWDxRCPTvHdDBie/chYz1JKlqO581I0CH55r/r5lT7lG4qHdfC4Bq9hN/S
5h+AjV/+jN8y+GL1BsJoPHYw/ZTZLKVssmODLngtM8AG3fH00VkRQafuf98IAZqGDhkXzbonkiOD
sDMXAVFq+KB1SP8q4zbM6utcM0zOCIiItFXcD1SupEkCWiWVXa0+Nh/5/sb0ekODwmC6xTrj6hso
Yrxt5CfgpSVKrQtZL8+0VYHyFSMlqPTTGo4WvGi7jyY+K69kRLSSy5eoDvpq9eGVhGJVaabBaBdv
31d9ZCzsPfD0ruBektButpbbLQKJlpiBXiIuUplXGdbG61nQmDVZYVpYtjZof6qe+mpK9YDhfGho
xqFjcYy1jIHT5IwhtugAveVjiwnqKkOjRo9mU/n96ZxXoFKOJRCeKrabYUfcbJ9Cf3wmWjryanKH
6qRXzMqCa9tHH3+APeTCPNqwFTQ8NTA4g0tJsO79ZnSJayl5AsOhROq93Ms/+VzWFaGuIPivl59w
X9zGL81MlUDhuZVIYZaPEhlbkrnq/2wvx+hocrZU+2asBuEttFqLeclohVyH9vqcMpQTE4Pj2o7r
3Qrmhh+rKlQwkoEWerrai/wfQRixuBf5gFOJQ9Frw4lusu9RFyaSx6zate1VHkIiucaTPxMQDMaU
dDhPZVodrG3FumBI/vMOB7XH9yUxkOdeHOqzik6d1o6/mYwVq8oDWE/wiB3zadlopTketUMEjIM+
F0zJSEW6/UmvqCgg/bOeKHk2TJ/6dddIiRozzLC3kFzD0tyB87hJjeO71u0zytzAlTpkAG4ylQpm
fy8Jun+swbNVEghRG540V2xMLFqbJNUQHXUSeggf4FY026rBJaV+eVe3040dCiNbNf4F4P8F1rg5
jTxozo1viMJ35zwn7KEn8ipjjpC1znlFSou7lsATasoK8IsUhG5J1X6vwliGLLY7wDrjoTyUbVZ1
76b7o0la7Et1rhhvIij8a8szxqNDXNuS/i7El8RWQy0MoKCAQqqPsfYTtWPYUBXctzLPoUosjQvv
1PligJY03KKoT81ENFZTGOjfFd5x51RXGuCLnQLtRW3vnRHaDfQX7tzDWpldYVGs3y1cOBDx7nJ1
v3xhYHjLXQ7t5viMp0S/hXog0w3vFN+IHu99WnSBW6Gk9JGTSAjsC0zeGbNYr8PF1bo2AQkirltD
q112+PQcEBdEITGRBSbw4dKYStAKUMgsAuWup5juDaNcPkA08oeuETJ6vqP4slZZIRvY7onHqFOi
h5YOkZy+3LOahOJqvoY8j/MK3bSIsHz3h7iKFlraM7QtzOLA8s2psRgTtjojurwJRGpxo4IrObtC
6pvWCkZNQkysZ4B4F3jrWIHGuirtpDErNlt7lmsTB3hgoXkgEGdFK103xO7o6LAh7WHGFqAT1PX1
XldoYuD+1RQNGTkkTysNv7XTkjKXN3DTdmFPU7p3SpaumYTLlHCQ8jufC4PWypSE3h+Pp2Tzb5eR
1usbZZ+SL9sKDbjgQXHS9oIXX09HrAJ943oWxPAt/A6WKqcx+k3tCHfnxdbsRaAsJkVQZNuRQrpb
sseIdl5Puf5ys4jPvVSRsTc9Fxr63Tz5j3qVJPwyTu74Dlwp3reZE+3RvAkkVCYkbtDnd3OSVYdl
z9KiTznEjHC+/EakAKq2GV8fEZIuRj75N+gh66FSvmNfnxs2+h5ELZavGXVijQ8tkN5L0WXuR80X
A9OfwBNhBWOmfXRkyzK/69leW6kbyRvB8pCwMHmshuqVEuUakSkTho1mOiYRKKohvzam930zLhX8
pY1cNqobnt65spj4EYh6u10lLAR7AjjYh3Q3VOlTAmRJrqFHAIRe2lBFb/DirByV3ddyck/9RnUK
bKawc6cNkITWHeMnBcZNkKWZhYei1dw7P/VuwjyfL87070YH/vbA4ZqTNsxOhspklJleut8LJKbX
Chq3JA0W4EhCk+omm8Fff4Tt4TceHnM76rYjhPDVVknmBBhPKy6A5CefsQgvJRm09Ufcb0ndOHp6
XxEW/haFUZsLvb7APiFK9AbTWF9w5A3zET3BWW2cOCuIC9nre1x6EwxRJUuCkrAAt5wqTY7FKs3w
Xcwym/bVmmYhp43gwtBcj4fRr9Khh0j5AQ9GvwulFKxJ+9oBHeQv9Or7k1XwLgxDkEyCUm+IuEZM
IWtWpYMDQyWZF7DK7gsKSzfRmqVNb25KPG02Q+ckW7u6EyPUafl0Jtz3my0IRsFCzOVTDNOkJ587
Mot6HJ+8b0SLzD82hN9qoO4syIieMKeWEzr4VOIVR6sFmmAubOXv6o59c2UXWMscVX6lfHfx4S4T
I0zqCYcQCTBZdcFs5sgud+JdFTZWQFuo97TVQvwscnwlH26BFU8Ucc0FLcjQhE6eRQeWN4HpSLlQ
tMoRwcE3Pt5LbCmS2yDQHPY8D/VTMDLMAtrsIq0v6OJQTC0Au4g/khyy2VCK2ne4XXEEbeOi1Qry
kidQoWuuqi9f6JA+vjUyz7cqCIeWpcsbv4QGvhFqbc341p8Ym7u3jknwov8B76pTGwrt1UR9nitm
fcme/nFW8ltm14DWfni0zIodxkEMKGLLl+5bieKhFK9qDp/m34Utwz04B558ozFYVmVGmbxwjeL1
FkOBtRwO+GwaFpmZGhXnyBuE4YO5byietOGGkgTkqYZJZ0lAt+UsOBma5oalekGKQGzL4XjJyQ+f
WXbqZUmUI7Hd3TIK+OxUFQAoI1yax5WGfZfF4x8ffTbOfL7ZWcMDNjCvJOLwUQu6M1jotH4iACqo
S1gnCz8YOz29ImFWaxiZMLQNnW650vUbFjl+W/bnXWDclh8Xusz/gMPUc9SR1TrythDMk+jXXp84
2oIJruJH7kiM2fAWcMZZhDlyR5CMHJmxMud7zoPjDIXdgNEMe1zbV7SyDK/SoXTbHu9KnX3g0tHA
U8d/UOIYgPo2Sd0UZqkhiJTjaBOs33j3wfwAr61RR1QDmXrYavNyRxmrgoez8RC6Sz+5NhSqcD2g
ufzoqIZgtv5mUjRRuW1xs6u7BOxDaKQXohht+l3gDqppHQn8/EBjByO2NxWQVBTV/zCPYH4NaUjV
OahPnD+3tJqyEFhj+OZG9fESzyNRlFt4AjNE6WbJk+SzTUiqscWvGydTj4mcn0SZJMgB+kiNUL6H
72pnEcI+dzm73HiONnJmM8ImXA3Nijlpd5Jvnccr+yEzkVHPpzXUpZldItnbzAW0z8fgt0M1sx7d
9285ctOFbIMkrDHIsZ9t12PFZiyzp0vIs7VEKoXh/L3U5R4zPNatGotqdFM/nJmDnYTnVveYVtv4
AE2EK+YNYvkAP/cBuwoNJPxWEW1x6EaqA2bjzAJcESoosK+OfjSC5tavUFOFbKyVw2A6DUyCeoOg
3cqy8NeRX7z4dxu2bHA3ADwnpkXaaNOsWpuncFT4EoZTv/LWSnOYohgE23/TLTyHrHCuNk8AAyJQ
f1nGCnAEeZ7iNCzURpTEXbfakS+FKjwpuIAjWcDYEB7RBm2eq15OHAfzCC0ni0OU6X2vGElR5agu
zYD7uOz+N6DyoOzzZDQsr4qOx/DSvFzlvwXp0/hxIFZsWlwiWnghCE7lppuxwdH6UK7TP6ZLXydG
/WZy/yXWxn0JBtfPRfHFEIRy4+OX/Dv3RgUb7G0gUcZO8LJkdiskBJig3nUKppgXiieqoUd2PJFB
hvdhLHrbLmy3eZQO1/98GfiYJvoKKQAft+dywv04+n452FLXGysWClsWaN/HUk4JmYTiyOGl55Ul
17kqxY9TYT1M4zd46yQAuzCSRk6ARojHvPkH2kWNxFhSnkRIdMkAePxLsNUIpGu0tD6X3yIGLP0L
3QL/6xAEKBaozu/yE73kjky9D0oqNBImOlah/kwQ90kKTW/HSHHKBBvGtAJoAK6UjFANMDImAAAW
5cDWeMmUdazXNT5Wt3WdE7IKlVfr0g/ApcD15OKJtj8gcH2IyvbRIvDuX3NBUib5HqhagX6Thl3P
6TfSGmTtljXlXNJRa9SUxngSHk5nFAI7C4bp+3/KZeCM6HXlb14Nch3r13KoC0+5x0lKojjtfXLl
o8y2N7cW/i41Q5tDO7eXPcLGM2hrLXjCZCsmgEm+6bVDzTV8gp43gQbxErIRZVVBHE59AWD3icvK
RLwt5jn7TUIz3q/95WUBtefzoz94RyU2nUKMP0lRxat1HqjrLyQXZrmSqqua7sJLZADdPksGfoP9
jf++8m/tazi0/H4kBKGTMrB0iOR1+APcG2N2S2ekLEjzCo2rs35OoaMoY60Vh/tM6x20sZ9T+VOR
LJqLxTWfGE5u08jd8qo0vevfLM/dei/2Sphl63avOMDBDl9lx77+UIyyL5nutdXP4+v06YzjgL1p
Wt0aLlBIQKBCK2ksUb4DY3RyctlkrR5h2sFguKYuFLgKhZQyJYzQf0N2m4A5gRdaRNeqzbkhas8q
tYTS7RHG2COkq9y/n+I5f/1T5perWVKOZOzwFEi4+Y1aWrPtcjhSXCFIWCEaPdbOxLuzYdJmVWUo
Gb5By7xE9cb4yDnXTsxKRm3cHRjJZ97EIMdJa2pcICURRZosRdaFZ/h937mVA25uRA4DmGFDY0JO
OG3UW1528rA8owawXGcQrhGuS8fHYlPYnSi3ZBWpGYMU0pnYnJnuEZSSFJdhhiGBWx5rxlj7xqn0
ceW2bdLzh+6wo0h4nia8A0mLoMRhOBL/hvP/SZSpTzU88XjQwh/GmTIdAaep4xOgbut6Hn2+a5wb
mH/zuduCSly3QaZky7IyubiQ6obwqOrPtcE6tO1Su529OA57Z6aD8UZgRY1SOGP9gxwRdYHliV4w
iULsK0vFKOoNfaGU8JGDSPLoewyF2e3IQHyZ/ZNDYy/mAbGpOH+oO9uP9k7G9DTWtP3aYvctMQh1
qm6UlDFIqfQs4MvMK6oZcRebC3Nn5hnT8mnRSfKOeowKFydk/+ymVkg7cOhgzfpnw8PGcHw0jJIN
6q7wX+qZ7Q0Rc/Far5cgExAIoWiK6UlAJKj3j3720j7zZ2TkTMhbNqLYfeHL6Sfw8e8oqrFWOkU0
M5+aWcRyVTGaCzDK0ENTVZ17V1wcd4TswvbjKGcVLn8CgD1T6affpsobX+nQHs9ffrz3xzEgfbxC
tS+e5iu1IubaVVH1fKbwSnBtMPt5zlDiZaNkC/V/lFI3Wte7Az/qXdHN7UzVwjHnRkgNgHTE2UZ4
BM49gZQ+gPX7unHjx7WtVVruXtRBZASN3xwsJxSTni485wKLF7RQN+XTGDs/KG3Vas/jh+2GlEpv
lvBUue5QdSnnN4TnaNbOOURZJ4Y6ajdRefwCV+gZ10KY2f00r2f+0E+uyXPrm3kBboNgGogSfzzI
ULakgetuLpzkqbrxrd2xtuy66uSAMABhWOuShwqxF0YbP6v9NFHIBYY4yQd542MjiDhq3EXITihy
EBHeEWR6sVDiqN8eT7iwM4/rtCmGcOOonR0eQcGOBzYuuSkhgM9D0leCNx394I1Se+08Rr0KhBQE
i4CZbWgHlpNFaMzAprMdOb0NeZfXc7U2b1PHoF1w9pyGeXusuH+XID1g3w/wq9P+NUP+gwGHqDph
o6oiLZiIaEeyLUW4LEO5XvMMu0VfTISS2skjOjIsMAc5zJ/47nJh+gPwc7URpWYbDtUddGM99yXr
nS25xvQ4a9rhWkf/nvPOoD+5nHJCOTp8FQNKNLQwCB2HaBE6O/f0KMsSqhYIcgZhV3wSUCp4hmqk
O4Vf6k/CQw57hZBGL+3Q6j+U1mkQ+WVlHkralZIBAuOeBDAo9lZ1nlZDoZBh8UqDjhWA80J5mSYe
xa9ukWxY9jt/3qEoo2U42e0jKzl77VkkzlLEkb+B/Xh8D++/fS+YaQgFrCREx6JbnQR9hw92DPkQ
ulhgnjevNtkja+QqQ9Ldeko0gZgIwMJ0FSKZMAcEsjuDxXrrAte4WgelDXavdyWYKrs2TeXqptko
Rxo+xwRXPAqid/L8HYs4P3QHgpa1/hLH3+uw/kQQFbELzXJAyd+UorlH/ICxEWz4IbZxsOp/pa3r
a0JXWJsi09tORE4XSLA2XwQ7QqQk3+zcDGIEA8f6LnWEwhfc6LyyZGTaojIQ42ERPq7i4g24tchL
ehG1yO45uR5kbtg9Pnv1EfRGIevr7GjLY2cTMpS3I6g4Auci9d1EKcbiS/mbz1FacfAFCFDmKNlO
yiRYBBT8dGaZKjmBUxT+SgTghu07aIyFAHnbsuIsniuZPMyEIjjRGYWs/ANFdToStNM7m8jplViV
d7TECLUNiuCCyaN6qtKTrwdUlpeuvWGPu3cOcrtgD/NFi+ZHNfHwIwQrC8tH1DhH7LkXTYG4+RSJ
UvjTzYInWbEWgR7GeDYR/hr8po6ckzFTZUXc4ibct8PuMA5knhJgd+ptMEn5wPDXToTLzqXwRFLF
UqX4PunpWrohylcIkW2wgocQZguV4eMylZBWhyzreHSzjkLQGRTgKwnO48gJTtPGEvolQlbjARCv
g96LLfXmEDAg1NrSaaFh1O2/OgNKv85D8+JwDNRiNu5VhYAvjRsBJSyEHe/5Mzzf4BAh6srX43D4
G5SsPmzrEQoRz+V1KbzH1zCYdU89VfIpLjDEEByXdtPln2iS2ZSIc0YDL+goQnNecQ1IQUK6UjRd
+rHzDwy/Ah6EzkbMT3yDeYJ2uKXDwJofQzFw/5sEALUqWSd2hP3yeWddpd1/EjeT0f7t5LvjVUEO
6pqKOKmy0YlKbqU+pIgCEmJcr6u1D34IxNpqFsHVOS2ZDIRXwggs7WFi3eQO13m+FGmjC+cz8fJY
Atn54Kmhhdko0Ih82KziW794rEKBLcHILGHoF98Ga2VaiorvU9P0bRhGy2cckjOc2itclcXDZWyU
mJxgWe0nUm6vm9IzDpPjCFxL9/vZTJZ75LeT903bFmYjXg2zRvrCLqWoPm1nB3J5OWf544JR7Yux
HP4yHVhV00Nl3y9yhDpRJUpNizeo/f+DNgZe5afzsVFdrbK4TCSUrTfx1xaGWDZu6oyx27YWhYWD
b4u4KUtn+cTmoCMSpKjiVVFfNIDlXY+I2pYNryL8GxYmiqdATq2+46nL9QjwctkMOWtsFRTEV/Jr
q/H9AmgWyen+rzD+8keF1LMzNMAgham0HQqFaBwosSpunUKBEcDUaDcLauzOaBf0b085oHKfV+vh
E0F3jCepPUVqIucXERSrmhkU2fNZC53LHBGdUcdcjekcchaNl30aMttJ2ErxIVtb3QZCiVW/b1c9
ggBDWfeCgroiBKpYRNZryOFW4MtExdCKpNtExPNMA6meJ4t2xDS8MJd0b/ZVdOTl5RhAp2AdrCQq
NqJuMkEH3HEg9gH7yrFS//RgfgpsQXhvHlZ0n7tZcy29uXg9ItxpFYV85WCQZ4ZERfFKx+Bm6/CH
itNK9T5d1PNK1RFJLTLkbwLFUWisNVRDWFmNtgzgBVq0hGPgsBPKh+5FbdOqg0rA+7Ie/kNHqP7x
E8CzsRLt7iBvJb5tmH+4jcxXHeQGQeooj//3xEaepQRGw+pPVdns6JYqzay8ZR87OFJDfDkcQi0i
3dI35JNuFfLpDFN3x1tfR97KBoscW9bmTNhLswKsEj/XwlQ/IRvRobu3hjNM554nAvZ9+nxUIUxO
LlmJ4pJQ37ngGhXfpMPCyB7Cy5D/xyapLGa0bx0elcN4vULGqFZT6NmEpR/jljdamgYeH5sMo8Bi
5tlQtGPZQqWUowXqr4EoruUq1+X6RdK9YDH8YnbM8JOnsSUEqmlVDg+AI98U7WeRg+JbvbDRmBIV
T8sxwuuj8ghgGNLxg8ecQXL7r9XXtIRo5W5IEBkhkxCLx7jT412akDWIbz1B9t9d1Dvp0oZ3FDMG
EkHhIm2aCexLwYJ3RO8KnZ2XkP09Uvk+EbcCixVNvEVfkoB9rgVJ6biDBeC3zU+0Jw202n3c3kZL
0IlT3SihsiRjO0B/I4mgKW4mnNKPPe68qIfpiIAeWwmMNLu4z54wjyinWaz+ZTJJuW9B1+qel3oU
K5eYHjOcIGzBQYqWsW54rt7OZ4FAU8Bx5Qc91dedTmTdZRhtuPKpGJyCaT4WihWdReOs1CBooVqE
BNusYtuO1EeIcEsY5r2oHBnt5zMkkd1PgMruIQeERvQWWJa5ph6+u7Zqon+Y1sUjSB9q/4qXpGdN
q2ywxnp0d19LJTTLrl9COEvT2BmFwyIRQfvDizUCMxyu6YB2BeFJ5BJ3FYQLp6CK0u742VZ60D4v
lbpBS66QIamy0xv+bizl/KKx9B2iEQwxWxxCWooK6RpKCRsYsrKShqJ2XpXhTR6vanx/Nfsg/OuW
CFFWlSjSCnSbkqXxmcWd3Y7veNoDkFF+byyZ/LfGTKCKsrVKqkaPp+ATJyi28ZRLP2c+eJg/ZENj
bf4/PdIyo2YdMb+Gyfpt5qRoJih3m1FDXI/HBE5E5bIiDs6bxqWWnJ+l307Z0LWabyWg0ryEUa1k
ezHkIrQEDcTEaggvphmVxHdg4c3+YS1iaLPUXhiMmcvrweaRZjCLkExWvO8x8oZbEOk1H2jGHQo2
fU5B7idaZvHnc02BTA3JHJ/vqSh8o/qQc6g8JTfcLmXKU+Y/zmf/U7YbluIPaltn5Q7XBvVAYJgQ
NpKbVAf/Iw5bNHkumBHc3KqtbxOKocLnxVtHI94S92GjPk1h1UtCzxYw16vELAVGsBMjEWfb7gQB
sVLlDTLhmSUgnPjfD6p2wq9KWeZxVvLFu1piKj2fU4g1/c3DmdULSZQuHyLkoSdD0F5ostkRbKRq
SMn+5Za26a2aPvXIH8PL2XTFofE+8gCUOwYT1l+6rcFxNEzXdq3Pzn2HSo8zcJw9I+0q09I9NKbc
ZA0SPEpDHl82xFgPVS3DaKnpXfPmSQt6bkJ0eNkAARpvZyagFEMnk3Ss8GtsZxV5TS9Fhkyixgkd
isw79UY2ddf1q7kj9WvQJt2Y9jHU5OHjF8ByIOy5+Ci6VP7Nnc0k7FzQGvxv9H/TH5ajNxMODtZN
45Q1t+wAa0zyLmHhzGIi8mpuh30iUbUqHnvDYlgw2/A9gwZDuEovaR76Osik+EcZ2PBgDGaI1pm+
GrcL+P0eXLm008c//wQuKq1fCuksu6m9FLYvM/9OnjzwAv8GhEapSiX52mEyMe0c5d28kRvBKjUG
lvInzXaj+GSLf5FADnEYo/9s0ELLQnG9SVvcahI8l8+HZjcOylOLqisaiNvITyUbXSQxyW2CJFP/
R5HULrXoAH8hmgxL+JtBRWbCdcwUN6yHAxhzgTBiL8P5jtHpOiYvLbuOU9goqR38vpYdLsw5zpSu
2M41Zrt1djtmYxerM3e9XPwKsJ4Zw3cuar8T0bCl1iVpG8qyZzhVpJMviHjVxBAM7DC4N9Y2TwR8
8+O4rOHzrDObDU28I7MEdFq/QuB3S2zMZxZDqABmwAoNDDz3T4hL0tcrOVW9eEcx8U0SRt+tEEbO
wMVL98WsPja84e8gn1svJcTywOLwAfJoNU8wqOWzxOMKdxcOH1QSLsX68RyF/ROFRXA5LvRulvin
W2rDPHpHenSQF6vajH+utbZ+e8ZG5eE0v90qm22F8FMRgkJcaPEbaYTc7pEXgt68He8wm05jr1qx
4hg19xTFdFEmSpdkzEPWDDAmwgNAYidwdfU21S0nj9/BlT6TfjMnzH9K8/1ptLOBM9h4tF43l/Pu
X9VbuyvNLXVRCj35noG+b9Zvwa0qrqlRUc8yZPkbDrmvB4tPUCS5Z08sQbHN1XbpMm2n6m9uGxB/
qsQnBa/ZYOstKv3dtVAtmV4aBtxUqx6S6kW9J31KNaiKh64Komnk5F0ZRFhLQSk2TGhlYpJKjP7X
YSKShpy0+j0v4KB8T36opK3/+iQJqn2s1dqfMQ1szmy73rGdP0zLGIDm+JL5QsMWJ+eXJ7ufnQ5S
Aq14sZ3pyYqQRGciBFvdPlmvNy2SLa4DYqr9FZ71E/u32vdvRpLZcLDIJngOrMku/jw/v+cvUJM0
9duxdsTcc63h96GXSc2OBPrEkq3j4V6QQ7BEOFYwMXecwS6A/1uV51157rd8InQgntb6hOabRQxV
TihbcwAVil1CMjazNEfcuWA/YarGHG4OmPqBGjH9h5MrPX05oMARTFL7tthQnPUHm74HBP4ek6YP
23ePLI3IMH481GJ1jB9LlkL7o0hRQk/fwdwaE1Ujd5PQf/blUuKuWBTxMgyMMRXaDceyzPgzQaq0
ve0z4rj+B5fTws4vnpKhr3JhUZnZuXu9Oss9Yp/N4lpeTnxJED3pW3YHGdtgI2x0Us8VMBfI1jgD
c4DN1so8UckIchNeQ9uyDUT+fnrvhg8kNJZysOD7YFBoxn52Vn3AA0Cdx6M3/7gjRlqqSADCxLN4
FIhEBBMYujVZ3y6VN8vlIyUONo+6qZKS9JAJqVcr3oU+B8ARl5GWTg6VVMBabVhljuOEl7oWRLHK
tgthXUOQgtohI0igs9uON+5RxidU2nBI7rGIdNg1CPPSwnE7/8ROoQEG5BTj34OC88u2a9ZDa/d1
TG0rJ8OovLhAfRe05TMp5uCoZYg0RYV9w/bph86P93wuVBB+R1hAb/H4wlxHo4cipqx4VxXZWyJm
3niCG4n81dDfgqnhxnu69y2l+EeE8Wf+uOWE6P8FzzGV7GQQ0HQHXH3Pvnwb3/MZumAUbF4Tr2mL
WMldwcrfFzhsslu9Ym+OqO7Zw2rIwy9cq7bg8mIL+NCM6uLfPl1evWBkm1YCWp+p6E0ZShQoZpJI
6qPBUymwExavKOEkI2dClIQEK19AgTkPKo7zsKReKj/lFZQmtHcQipxqiGOZEPjky1Tr00ICwh5A
e1Is4x3DbxKMP8briqXCkp7j43qPus650XFxa4TXgh4AMChCai8iOc3UqvkQMgNbWEor1d1LMRbf
TWJpRwbie/dyZlzq2FTaN+/mQ7nFrPDjTds9NWdZvLgruPrfl0auKSlB8r9lBINyTmVFOAilT1zK
xRCWddOh4zJ3S3D29sT6asmhROOXXM3/4McruIShqgeojPH1CUaN9tOZ/q/e69eEIq7TGUsqsOrv
Y0TInLeNpyC1lODH7NOCW6bCQDVCw56LSE8Qw+OUmm8J/U/WpJYUonbrEGyZV6dIZyzA4ZRLzU4O
2tZyBw0Jyak+3N0/yRww6VODGQAx+giCdu9F7lnViuGf8a91LSJ13nr/4O1KaCKcfQy+CyaN0p/E
c7JUZ2Xh5I7SYa9u3qjz3QovbEKt0tMHwL3OOQq8kidTZVHc+BSsy2VQFposkNp5a9P76yh7NZCj
X8aOLZ6/tTkrWiD2ZGxV+CREak699MQSpcr5c4J2/h9ygm4kNYcvBtsPNSvvhEtPXqAA/4Uwalol
5MVvamupo00tQ3KwztgFUDCKNuFJuWrQLJyZcYd/VcSmK7NqBSvk2D4qYqiLPbErIv8RD4gYeZDV
Af2v5GILnbyGaVjh0axoG/Jf1FoKbmuHl6/316ndBrg8uT3+r6Jb1PZkfHVlMpbHVwRRv707Upfp
H9E9uhQ2Nt9bf3ReGgXZoS3617mteEgIMQuJ/CSzuYKB1n2X8+86UkRkitUYO591On9EzRsgsp/F
9j/yEa5mRzLsgtYA9Ro49f7fTnyH9Ysr302Id1x2uGBplj/xfNFZUBxWG19ZqqPi7pdUJvySpg9+
l26ThmQl6HHJpRuQuJXGwAOgwOoBLSaFpbCxuBRe3LjmgFBcFMp6DBvOTAsTvyPfHdYNn4calyoE
ajX2vWcQggVfS6j6LDTobJEQoIYe4tWrczDjIfkf1SHPFT4LeoBQGcF/5v9J3/5KDgqtg2oNAfvZ
BvxZ4GXz1yf4bKvq2h9pLka0dU1HJAvuYZbTZj3CCuO8WP8+y7He0SWKmRBnCwheZLVWeR9Rizjz
Tjyqqp3/UNa+8Ho5AbUVJ9jiNGgX+9jo8gp8t/RoRNag9c2qYowDvSXk1DbS/odX4IrZqGdYUeuE
FmCdfNy6u6UcmZJBvtjG8xnt14qBpvIQAnor3seu5oTnOiqyN/dF1HlizFAqE5wtd3wAGnx3R268
4Z+R2uhod2af3gCqURk4rZ3JsXdPYzwYboQWZV9drVRdcS/ocBRFiG1uuZMwbJhHb/KJEUbXy2sZ
jH0jn6pMiqGGd8VhkSeLawhUXCwZqzf94Oz0nVMOuWWSUKZ8KFqqWGfHDQ+Hy0HwUO54ZsWLacBm
VdxTw56gHEDiHSOWIUnq5286tVQzHvPQ8vhA5bbxWD59wmKNtqrwtXkdsIHzFGmxc3q9WDv01X7L
FSWmNvVVQ7mirix4FryOpRapZgEBLhlllLE8x7+KfNwYmEdHBVlth8uczmdI05Af5lO+ZSCwAnqB
Xv71/nhZ2GM92FPhru+BjaOOwAyx/73HYMxgmLjhyj0wseaajx7dXzkMt1ov3o6BEMoJy/L2NTyu
WcAIAiA1v1HSBTn9+Y0RFWHiPzAtkI39afti03PTbn20AC1H8Wu5mwZNuNxU+hsTHj2PwhGmenJt
fG6MomEeLJbqdCehDd4QUbQTNW4VKXRj6JHeDKkRPEZM7YwT0xClKFIrC9kic8VBjYUELD9vS6le
td3AwcPsBeT7sUnZH83zRaBuLX16hp04/pFotXR6alD10h7yFc+YIg3TS03fJmvK4gHeNZVJcvEB
tgluzi0dQsZjDjo8jqx4BQQgaSEFEhv0olaZW6NZ7NB94K06GhHTMQgOPBQjUP0Pg9Ue3T5Lyiap
Ydqn6wyPs0J5E1wx8UUVM3z7jiZU7liKyxzIlWGONIiGKpP8NLoPEfPJndP6om3ZDu+kioeuFohC
thwcwHxpAnLe8LO8ZO2urpGQH8bMy1S1i+w2jOEAOnGUcoMNjgVrMYFY5sFQ9sKfwz8UTTj+8/R9
XdgHHVNy+KYU+o6ECbPRptFXYlIIBQ4XOUfC6BMhM48+au87+1a7nqfOKQ2n5yKrn6xd/K/VrmSR
0xDwKHgVl3ygL6vWE3+9L3Kch4J7pdmXIA00N6pR6rMhH67gcywkKe2EKZP+eeVP8n+aBOlbT4f2
72AndJ0kw0sWYaloyk7kFV6ShHF3R0lnc2Ci2ofmWIb4gHfo/BqhkrXV4xVrxrvitt4KMxFFXsia
JZLUiG9GJzPv25IhgsrwcUGVzzbOywuyXw==
`protect end_protected
