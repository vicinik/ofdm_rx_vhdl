��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@����ә5D�yJ>��ɬ�v'3mj����7��BgJ�����[�mK�Wj��k�L�U�$b��}��pz��Hᡬ��\�t�;/J˟6���PGLD��?|��G��{��Jt����ּ�
O�>Dm�Dϫ+�'�x��ޓ-��E��.<�nY�cc��+�1��K�;U��X�4���+oւ��h�T9Mj�Ғ�$z�����������uJy��D��k�B)E��ԫN�-Nܮ�*�<�-�T�Kg$\�ǿ^�c��O�,�N��4<ܠ.��JWӷ�b�$CI+�&3�uB� �d�u��cf���f��5Y����`/$�.)��T�-��v�	�i���KV�ۺs.<�~:4��ڔP���6|�9g�'��d���/zǿk#]ɰ˸~�]�8)I���bd�^V��y��;,�p�|�tJL�v��mM�b�����l��獩O0ZP����nڪ��+ e�.�s=s��j�R�	v���PȲ�m�����J遙P�:KG���+�7�ٕԟ�6�(�'*z�s{~8�� ��o�)}<�M���%q���G��0��z���Էx?��xp����?cJ��a������ht�
���6ҍ�|���� x0��>i���1ȯ���Z}�� j:Ղ#g�MBP2����Փ�$�k�μ����'s#Mڸxa�fh@��+�@�5}?����R6�'e�\7� �n�k��(~�!;ZO�ƣA��z�'��ZfRT��O�a�cw�g���U�/u,U�@�P��6+�:�5Wˏ`#�is�����*�sS��/�C )��z5�q�B�T�k	�@^}�|)��f����)�~r�v�-6�C��_�b����=���oO'�as��Hm_����ӯRp
a����ͽ�8�X�/n4e	+������^p�:�����%Qa�#:���V�Z��۱�Эa���5�|���+��s��WL?���9D-�l�9w������R;ix�Pg���tIE�C�!�z9��4���!��:4 �L+X�7`l4M���r��vR�u%��|��0ǔC$�(IH/�𳼡���0R�蹽�~�=#P.WX`�X�$�zHi3�
wyQ��;K��E���)�}Y����"8!j���=;�`f��bϐ���P~�@BB��RX�$�n���/+�T�wK��2`��+xA�y/�³��RÄ�G���y<��6ܜ|�ѿ���Ԁ="�#����[\�8�P�`�Ҭ�^m"r�v+-z͚�x���>�4pC�l��M�b:���>`���1�"忨0=8.'��Z��㑊�x4�v8N�L��D"�Z=Y�b#���g�n%:��xہ��&��_��YN
�}�oڬF'9&%�a�o��Y0��}�aTI�B_�t4m
>�"!w�m�):gs^����ӳH���. ���s���;{5��lUi�C�v��
�h��L+=��_~�k0�We,pJ�-yJ���� Kv�*la;���P��T��W��<P�6��h��#�K��<w��^8����M�)X��Wf���,,�y�٦ON�����vd
 ��c?%��$�.-)���t�4_s5s[����F� ~�ߗ�;��V!?b|�"6pOY�mZ�M���w�e�9�r�^�<gp#���]�Գ���<��BL5�PU�/9{?T�T��-����꨷��+R*�+܋�B��7��a��W�v�����\WS=�T�Oۄw�b9[��^��؞�@���F�|�G\[aBaPs���4�>Z�Re��A����(�,7�����ꎦ�5��C�{��l�! /eKm�]D��?�V
q�A�����B�4���Ds>�H��SJ�X����mEFN���읞F��gNK[in�����@�5�<���(���ώ���C�NpTԃi�s�Ť�43�,9��܇�h�9Ȋ�U�ḵN��l��%G�l���l��r�4O䯕��Ư�yo�D��Aju��+����/��Y,�8�5�����Z��b
��E�֐�,�zGv��ϯ�v�L�R@�ڞ1x�Tiz���JJf���Oe�եkr��'@'���z�x?���1���xoU���sb�O�����Vǝp���h
��2ݷ�m��:�Ǯ����"�N!;���C�͟�7��@μ�l%neC�P�sGX7^5>�0:�8�;huA�J��ǭ��_�>Gi���~����
-ܺf�!������%��!W)���k���9����
�\.ZY�iytD�+�_����޾m�0̱)bwm}����z?�\G���?�ƌVD���b
)+̈��9�4ct��Xw�)ִ�:�/��haڵ8�-����vI�����{�|�۲�qr���P�Mc��L=��~i��9���nZ�q�jJ�y�(�U���@��op��c�dKe�G ��	�tȋt&L��0��׮F<ܝÃ�]�S�u�)��s���)�z�+}�g����y���5n4		)����?gY�M<p�A�@�nA���,����$�?3�5�T<���h��,��xg���L0��_ePڄP:��-�C�h,��ʔ:�?u�Hh&>�$�ag`}ԍ�\9��6�˼�-��~A�u�u������L"�N��F��*�#�����YamHt�]�ޜa�q��:�Ga���޶�'��@��il�F ���[���Xb^wb/�I.� ߍ�Ñ7��dWs%2t���I�'��%x0o�S�O@�AN���F�/��OQ_n��t��v�,�����9��Y�[Α
r��ׇ�0U� �ߪ�QR�kD�[
���rܸ]7m]v� ܡW��c{h����ݻ<�^�g�$�c(�I��]\q{�k�u{����-��dY?�c.G�b���~|HF���d6�㴛"�Ư<��$C�B�a�c�"V��6�c_�����7��%1� �v1���%�����@J)Њ�)[�yh�/�(�ēz�cS4���`U��)*� �:T�]<Z�Q����X�ۦt
��Qz^����Vi��qޏs�@*(x�VR��[q�
}��nS�SW�]�Cc�)�%�>�x�4(e-�^��I���Rz��
6�Hw9�M@�5k2�[cy�E���xr�Dh���+r,>��A��6���z�2pt��n!��iͲ�?3Ql�u��Z�R2��_i�窑�K�}勰T��g_���ň>(@���┮�����8 Ƙw�?��D�o~����>2��ks�>�|��Ǣ�u��k1�0/�?�Z$^B�|�3�*�ZN�u)=|x6�����f��N���AC񶲌���uҧ�k�ƿ�6a���j2���.�hj���&%�lc�j���;��^�N���7x�z:$<�x��	7������9\���yN[{\��C9�q��k��_�af՚_3�������'��K����N-4�|?�z��;ּ弱��D��[�fX�~<ov~�,bJ6�=Co�;d�mBsi���Ӳ�H�3"+Tv��4E���f���3<�-eTv����xb`��)�������,�P�����w�p��Ԋ�T�.�Jgg2����A�4(8�4�a���6<�Pf�kU����>a��}f�k���ڮ�Ճx��(���ÚG�W~��� x�f)�@������Gl��kșI��ߕ:����1�{���%�?�R��o��if���!ځ&4��4cx�У�����l�{�H����yЀb˸���U��?0[H(r�;�5���Xc����$}�'�dc�y��G�+mYH�q�#Q���:��ǀޘ �*����D�i� �ʱ&�K��ʡ���Z��>"�=�&��O]���\��OBT�	��hY�Qΰ�g>����KK�7�m'�k��i!B����]V݄������P���hm�޾���o0��v�imtif:Qs��8��P�K��%s�l�R�a����̨���1�V��9��>�f'����aG/���F��Y��W�b�(>:�cIrˁ��	��۝��Ҙv(�����M�F��OjX^��5ۧXshQ}HzJ�:&S�a9�z�cd����;Xơ!�*�rh��lδ] ��7.o���	[�(�8ˑ�G[Q��%�%�8�5��O{y�t����������p�5�!��L�Vƚx���VB*0��!�25���X�� ������-��~��5���>�.����ףY��a��T��l�H'�玭_�KO�*yҞzd�wѨ	�l�u&0��+	�Yߎ��H��z�Z���pR�*Ĺ����z��j�&����3u���5����LR\������;n��C ��/	��h_�a(]�())<c�l����gK����#����\-.(=��r�����рS�PH)�;չ���S;~<4S���Պ |`Vi��6	�6ɰ2	�����"Ms�2fa�I1����=�'1."#W��M�C���qA+��������2�����+���z'�;�;p���;`Om/HE��O�E�����o[�VDʚ�"bK�Vk���m�[�>�Hw���*���Y�NM�[�A$�T�f���#��	��~�|iQ�˰��#ۦ �x2XA]�8X�DQ!&�/�b:���i�q�o���c$E8���O�Mi�Ѿb��@�s.�p{ކ!�����Tܾ�_t��/��G����fj�\!���.>�2��n�XU0ɥ����q0�#��G�"�r@���:���C������S}�DX�X�ZS��K��������*ؐc��h��!�"eDP5i&�St#k��J�l1�HytQ���b(�\t(�%f����c�1�أёN���MH��E���ŗ��8�Z8=Ѓ�>�����y!x@Q1���mM��%�.�44���x-S)���L��2�آð�;*z�q[p3�B��Y�#���nP4�?P������͌"�3��77��=
�	>�V3�0��N��)Qe�bT�@l��/��)9E�T��ly� 8,Sb�^�q��j�� ��X팚��/�.�����	�W���KS��~��`3��)	�X]LR0���J��!�"����3tcE���i���ȥy�*�
t�Zn�N#=/��S\�Z8��;K�2��R�y)w�%��*������|ֶ)6�|0SY G����z�;*�	�f��I*ԙx}x>����&�!�y�o�L^D��K�Q�Y�k����'��죊Ӈ�G�n�<�$�r���ɒu�/��
(�Ƴ[�(��'�G�h'�}35կ��4���>�b8�U�U���XfDrή�����<�X���4�:����|"3��-.׸jӂ�mϔ�I�T�b��[�{fVЖ�>h��E���ŗh�X�@�:h�'��	
��K+�D��2D�A��������/��O��f�؏��t��]�gR})#05QX�C0K��y�{'�4�VM���^ ���<(C�+�FAW.�kM��J�
�F��p�iR�Ǜ�`��wמ����\���O%������ɗ�<k�1d*л�.�aS�Ʃ4���kQ���� ,K�$1`/q"�w���q
a�W�_L:�o���5Ix�~�g�%"_����5��&�^Zo�A��8"��9T���������.%�8�G¡����ȷ@N ��K�F���"k	��%�\B�c�:��"U��bm��IN.2R�7lN���w��1ͰO ���l�졐�ݦ^�җ��_��kNN]h����{���+A���FEct����J�K1�l�uY������e���
 7#�b��mK��Vs���\p��[ڠT�E���y;����x��"���p�E�!(�q$f�3�Ca�f��c�j�!fm<J9,��7����h��2Hl�.<r����|���.�ж�o�rۖp+aMǲLe]D��cm��������������{c�>���Hc���:��4N�}�����(����$W�s�Vp[c:V �r`�t7��j�ۙ�z���(0.���HBj��y|�T��)7Ңt�TAs>ZfiB�"�S[<OL݅+h,��������B���~NO*��A�ӜV3#���V�ρ�rF�Ne�FG��"aBm�c�;BN��!3�Sv���bH�@Pm�\Yػ�A*�����˻�ϖ��B��tq��g!���y}�c��C,R��Ҭ@Pd��Wc�A5��d$p�-@p?�ld�V�Z�=�V��Ft�Sï��&l(:5xӕ8s�X���"���?!=�g��M@��h����:�JJZ�Ǜ.%�O��AG~o{��`�Z�(��`��^;�o���sms��ʙs9� �^5ep@Ia�;��#���l�Ŧ�31����&�� ab�P�J�������_K-�,",}��"�����5��g<�b�A�Ѓ����AU��Jo����Z�������L����/<6�d��	��$�F.�����Ŗ�����"P��P��L3���8	r��������v�F���qm���姇����T>DԈw��b3gqO���x1�x˓/�M�$0�6<-��tĠz���^jn�{��G���vWMff��׶,h�������R�2M��A̱��:���5�����ҵ"q�!H2Bs��sqY��V��T���U�	�#���=!�m�.9*��-�A��9($=$��k���`�tBت�Ԭ��W����	Ȉ޵��L�� �j���7�m�	ԣě���ZђE�"��H� Z����d*JZH֢F�"��Y>O���d��R�4]^ � {���7��8�E�!�V0�R���qT �|�>x�~t��y|�	,>%ws%w.�#��S�b��p��*��3��#���n�z!7ȆU|lj�f����8�y�^���I�Q�w��B������$d�]ɇe�	h���XY*֊���'L�T!n�=U���*���~[����"�? ��������H��I/�mz���"k�IP-��C�v��^�����pU
[y��rמI'�B�C6��"��	���l��u�7��v�4�#�k�:���,�/�����S�Tz^q��g�2�<+���?kĸ8p.iD�{�����Bt�t_���B�TO������s���!.P �Osu/u��<B�8�_Η�7 �r$�J8NX�]Z�X��LbK78 �u��
xB���P��QnL�#x�Sn�N�`'���6b�W>����2�;L��Q�'�&a��qy��B�Qg�dZ��B�j�Ѵ�t�Aj��sj@5�%s�G�3g+t�d|.A���`���BuAЦ1�y��IS���D6��U�?�]�f˃K��e��>3jc`h��!�֪J�8����8��c`�t��2�Ҽ�z��\��*����w߽���g��ɟ���G��<V��pI�5E�o�[�b�ނ��uc=13>���~KO2k;c�1�|�E�7���>��c���1�%��?:�Ͻ�bGB3'ֲ�4,����">{������uB_�&-��q��9���ycO6X�^�_~�zI�}VU ܀�ɧ��%�,�Y�l(E�{���*�h8