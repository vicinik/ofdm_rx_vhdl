��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�@�9ڇY�)��R��]Fz2�n�fӮ��p�� ���4¨����,�o̟�B:lJ捒�{^y�J8�mm���b����O�=>k�3�]<���&�b��p�3kb�e1/}�'vPL �g1�Ni5�+Ƈ(�(:����	>����q�@�P��w���vc���3�����+�	*��ڙ�:oP�T���T�./
�N�P,q<s}o�R�C������Lgr���&;7[
t&����zz�����x9[�˩��3҂�qƄ�V��8�_�FSt��,Vj�Z��"},/�:A8�o/@Vw�y��I����ԡ
+7$/�a\ 5��I�4��^���3\.�8\�71�:����O@ d̞L�^���Y;�G���>)�7ۃlY��b*�JL�k��^Ӡ�}�@�,�g-kj �E�U���Iv�Z� *#��!F��X	l�fݿxH�Z]0J�|krr�Q�����������8�E�vpUO���Ue8_� T�i���'xk�ɧ���ǀ�,L�� @��TU+�K9%\P�9�W���Q�tv�I��Q=g7��黯^�s: �$Y��,s���q���Rj�E�4�����z��r_fs1�\��l؃.��T���gw�~���#�-������%6�@�m�&cH�yJ=�4'nޚ_�*�C?�c�.x���/�A�*�T���F�N8�o7*��-b��uٶ�b~��eQ ��N5�y�xjե���%�t�/���1Du��!%�\h�F<^\���C��r�w���%/s�]�I8q5��w1ұ�,��$2L�GL�Rj�SQMUY��� �)%!��&���ͣI���:_��\;ރ�����t��Y�C�SDNT�[���e�8�d�^��x`����>ۘT�{QD��h�"�=��(�*M;����ì��	�5e�"+KĄJs*z(#^���@̛��C����`S��&�1UI��
p6=\̋h��LI�)�.!���`9i�0i�Oc��D2���,��I�r�R�+��uu7SKƆ��rs;�	&��o���Mqq'
�S�����P�ƒ�VφҺOS��z��b�`�t�N�X��m�Yc��m���&�a[�!���_�D�g^G�|)�)�u�yL(Y@�I�rw�����.�a��'��2Zf��?�V���hc��{����f}��2�rwI�(���� :G�����s/��p�(��!�6nՙ��k��c�n�����V�.��W��fP�����9���`I���M�F�P�p�� 7ˁ^����� ���YX��9��6^��_�TG<��|�=må��B�s���W�O�O��{M��9Q ��������N{"<>�yZ|��gጜn�O���2]��L���@Qߕ4»��DD�<*K����F4?L����d����Ǧ>M��cy�@p	@��!ېϩ'I�1"�5�@S(�J����p�a�+.��l��'���A?��"� H7�\K L�2!Ot�1�1�&Fʱd{}L��)�y��=��������{Z�`کF���x%��sNw����Z��C<���
/$aZ��ٱ&Ky�m�a��/ehM�=<���Z�S��6���XK�R��C��$�_œ���vE�Ei�=j5b��v��`��E�����d�܍�=U�8n�4�	]���歧{��'ش�<C�f�\���>��׍�H�Y���E'�by����P���?�iX}mJ��Km��"z�j���ۜ?��+z��nX��O)F&̀.(:mEf�qcr��O#>�Ŵ��ǃ>�6^�L9�fm,���V<�v� �'���t�gL�����X���*����D~rգ��=)j.���Ԧ�|f��0}��Y'F��/$����4\1���yQ��J�&�@�S'q]���]L�Z���������\��9��4��. �8�C�*���46���q֤Hu�Q�թc�b+����wG��	�����%������Z�/�H�/�RU@5Y�(I�y��CF����^��6{kJgw@1��2!��aCF�ϤG��_��hH@a�W0���)2�m��H.��A���)�SCP�	e��¨X��I#���+��}�t��Kz|hB[�:�'��������Ù�� ��n�@�k6�����B#�u�F�T���`����;�h0�*D�-DX;�W�pez�����������b�)[�P^|"=d���Lá���S�z ��$��p�_����diq�ΪReR�i�dSP���å	^Q����d>ZV.pډ�����ر֏��XuPd��Q�>s�
���	���r��	�_o�t�����Q�ꨑ>X��6�-F�p����焾_�鞟0[���w���c��m �  �i���=�zĈ�x�ɕ� R]3����+1߄���D�*-�7�e�8,@X�]�Z��	g׮6W��#D��^8w�ۿXbsN�,��G$��p^����n��ڔ�1L��}v��a�7<��UJ3�T�\a��`[�G��\�!�ewi<oVZ�S��G|�~���+�Щ51���Ew��j��I-./���X9X>\}�%���Y���Ӭ���
9�q��~8�K�0TTsw`Q(N�6���,Q<���{R������%W����T�H��o;�T9�d2�� ���v9p�6�X�k������o�o³v�L���͇�E�.�⿍ν�5��
+�Bh^���P�u-�c>�y��t���X�F���3QC5���r���`��9�rϨ��s[����٘it(R6��JV�K��l��H<B��.z�]��4b��E+2/���k�^XΕDD��4��K3b5�"U���,��8b'�L�-�(۝�g�&�up{p���q����GB�Q4����rl��fK�َ��)��j��G-u��
�0.�.A3�`�N�mE���}<b���F���U4���U	F87��n�2d��'T�0�?�@�BU��c�tZ�VBMP<�^Z3&��-V,�Hǵb�
�t��|\��`�]�o͸\��9�0d�;Lc�W���w���m��#��Kg�yl���q���ʟT�3��� ��<>��h�ܽ��<�O�D���}O)/ur�{��~����q˫vd?��G'����E�6��m]7!#{dW�i��Z� ��~P�j�`ȉA{hy��T�Y}���`���a��7�{�9h��<Mu�h��j̴FӤ�0.�)����6�Oz�n���<,�@��7��p3Xpע&� |�G����:�U�
#)ߩc_�qѐ^��`��1o���s%"My���.9���(E��u�>O�/<�Uq��YtT��k������I�\�p>"��O�-���B��E��d�a�y������{�x��s�����V	]�*������{��W�i]���+N�H�.kd!4�4�J���f�bB�ȓ���
����U~'Z�7��x�2��9sYmQLN,ɯ��5h$	+�C�AuJfOUO!ο� �X����r7�-J�qК�g�I0S�'���]�
�']O��g9�Ł^�/�eο��&.j�6�\l�7z��
����)�0��P˹�eK܎|�"ڊgᄩ�u
���S�E�3u�?�N;wS���4������|�wd�	rp��35��%��n����g{w�ro~��c�r�z$:^�d��a3B/M�ᙆ�i�Ή8����?Ѧ�_���N=rzMXy{]�d���zO�[�)2&����g��7�5͠6�J�P��Ң�5]$S���H��q����*,��o]g���3��]�)�g!�����θ �%5�܇�w,�D�7�N+�f�E���;/�4�����j^j��E�Z�����'{��R�8B�W�K����-�$�nT�UT��! ��CO�W��-�rE�����=7��t7�ӿ�h�,���i�T��~������j��<^��c0�ʊ l��c���z`����]�on&�+O�7�0�c�x������fgT�?Z��tO��=!l�˫y�Ux�na��� 릧���%��]���HP��S��>C�q�{�B����k�L�odW��5v�ؚ��u�f�5SوV	�)��sc)aҤS��ˏ
��A]
73?���{��CI
5���(`���W����E�r�<g��?���䇆�/��Y��h�EM��]m�ϑ�I��W��ժi�,�1K�,p��d,�*M�����\_KY�8H~�S`E����������m�|�;�8���Z;O�R
`�'�p���HCԽ��19������;h��)���W�L�6�������3�������+]��#��\ ��o�J���R�k��wy��+9�񩝙BRb��å���3�Ã�|ƴ��x��\�E��2����ۤ�n!XEBY�.l��P�XB3�O�~�����V��h�2�u�t��h7d��Sh�&����e�2}*���t�܀h8c�-���r�VǼ� �_�S�2���T���kن�y�22)c�F p��>�G�: ĳD�t@�d�ㅳ�h�
�!��ŽjOcVq9>��Q��!
���}��?z�EEc�+~��,��g���Ήh�!�) ;}��"�P�w�l���r	,0�z�L6p�$+;q��J����j�Ŏ˭8�W�G�%�Ѝ��� ��L���$��>�N��j�I��m#� khj��g=�x�i�E���q�z�t(��psK��|����0�ٸɯa�H(����Qfr��?)��o���g�q�V�1Ɵ��:���^J���DR�}E9U�&;K:�,J����&���8�ݰ��^��]�>����Fut�9����R�q��'��*�e���<��Q�31@���R��)��:��ʱ��N���>U\g��/��0Hks�Y��T���f.�c�
_��B��V�N��1�U+Nm����_���b�^#j��0H�By�Z�^�X���u�X:�����e�z|ĢO U����^�g
ҥ;�� ���;�0�1'��47��[�B�;9	tk2<���,����Sh��C>.0uރMa��&�cd��R<���=��z�������He���[�Q�\�����P�:��Z����c-�Q�"���לr��vk���K�L���D�lH �!y]�A
RCNT6b�����'IX	� 6S5:t��V�����W�{e�Δ�$�[D� 01���s�W�O��P�|�&��:��'yC��5.J����1QP|��_bUY.�������Xq%�,*��=��	9���9;:k��j�A��P�0��n�;�t�$������&�/���� W^D� �*��m�֓[U 2ӧj�b5#��b���i5�NA�Ӌ4�H/�h_Z3 9Iti"X�B�ߗ�?w�ܶ�Wؓt|�1E�C����X��ĭ�L�����T�K�1��d�����Ed���h1�Ճ"ީ߻�E���p�+�&S�#�!/x�%�6�h�m��:P%�ö�*� ����+=d��N	\7JzB�q�$Q�=��܁���V�ڕ�Nߐ�X^���"�� �j�T�Hǉ�V�7Պ]zH(yR��D�=��Ԟ���'b���J���x���累@��=�Ɉme.A�3�~b$�)JT��}����!fQ� E�h�o������#��_��x���_�+�n�^�m�+�'�T�h�Эrpe0��1�	�y����{�9���o�<��Ù��q�o%p����UZ � f��T	�qc�5c,뎄��e����")�"\��>,��̳v�B�5�>z�ń�:{{����tî%��^���+��'
��Nd.�6��GzEwfT;8�j��%��_��Z*XT[#p{��]��33�F$i�� +a$�m+9_��Jj��H:/ym;��#��:�+�*�������F[�^z�֐s՚|������~�u�d5R��L�Zm�����߁H���c+�X����"!�s��ֲ�ۆ�E�Mə#�C\���K����1�d�V�V(E����0՚q7}��#�%B�i#���_7GQZF�Q���l��~�G��n���_��z���|�bJej4�9����`�!+|��79��sի�W{�@v{����<�Ciz*�ϸ�᏷�t�S���|�%���K��˓�����J�H:��7��h?�\.(߶�h�GG���L3���2߳Qt��Ą�R0wၘ���Y_Q:�A?��%�b�a�c̆#��^8	����l�6M]� 
�G��TMs
B��5Ï���M������bs@����l�\��q��u|�M$l�;Pd���F=�
O���ٜ�B�g'x9|Zw�PnDպ{%���T�3L�ޒa@��`�v��;ȓ����E�u��>!u�J*�~!�G��Խ|k"��S���D�c^[cUm�r�4�nc�(\���2����tD�yy�͔����K��$�<�[�y��}q�w�������ʫ��qA/ZBÄ(1���̱^��8(sK쓼��je���^Lk)Q����sp��4�^Лm�R�������V��QL�H���oOyR�|�8b����#�K�b�EY�mA�];qph}\0-�S(Ԙ6X�B�%��bJ��2A��[�ŴU2�%NWĔ��L2c�]SG��������κL�5z/��/+*Cbb���(�׉�6V��&+A�7�zQ��_�o%�%��ɴI\r�5[�8.���*�0��h?���O�v^Lo�G���'~[�H��?(�� ��6I��a�W��I�I���>���Ce��p��zg�hq	0j����Ŕ"1׬7@#��2� �����w���j�|��T.p��?�K� ����;�1 Z��\��9L�8�" �y�i���U=U�ŀQ������=�#)�j�Eӳ��m��%k�h�@X�r�����:f2}]�/N�	z��Ҩ-i�_%a���߄�<�ʞ�dzr_8B�M��)��~���K�{U&X/N��y����x�p
EZx�O������1��7q���%>;KTǛI�}t�����w$j��Iz]�G�����(�?�ʈ�R�,!�#:��e�M��F'5��b�+��$x3��Z�臫�J�H�<ui�N�ѥ;`���f�X��s��A=6�_^�|���u���yj[��T|kF�C�g�1zq�������)�<��29��t�/���:簠�*7m��ֶY��;�U\��~�=�ED���!͟�l��(z�x��.��ԓD�����:���0��g������!IC��Y���Wɥe2�T�P�-�����]v�l��k�lϭ�����B��^$����7���٘��H��þ�rD�j����-Փq�hYzP� ��W1��`ߧ���G�Ǫ.�z�qഌ{�̀���}z&w�d�U���6�F�d�i��.�����«p!<�M��%�s�#�����]�n�x�v�J#��(ՕD0���/J� �qd�ܬCTm3��U���zI�d٠ ��n���u<�A��?�D��ǁ��K� J��3�Q�˅oD��SG�0��eɿN0/n����qa��\4Izu�ðA`m�"ی-M���?���H�aGu��'W=��I���
�ЖѶis����S��˒B<z��������TYm�
]>�t�r��p�����J5��^�Pbd�}"�`�U�������3�v�s}�j~/�XS.��هɠ	R�?���^�oGtC�u#�e��e�r�O����K�5+�����mj�i�VR?���_XU�5.�e���\���+�<`��<�l\�{y��Mh�{l����=ma�2��e���G�쭿�C���/��6�R���ԛ���n���<^�\����ĉׄ�b����v\���#%�ns}����t�+\N~:4o��N�-yu  �b��@�h+T�����m�:��ڊ��~�Cf��f�Ϝ>���'�O
���%�<���e(��#�Iˈ5���5�U[T�tm��}�-��g�2�e���CлX�k)��G���r�"���aX��hS��7��}��W\�I�	H{�%E`l��;�7���.Z�YKC�0>T͜`��؈�	Mw�K�˺�/_�*]�W��n A?���Dp����V����M5ۆ̻���� ��/Z��o�����cq���B �0��o'��2��0:�Y"�d�� ?8�Iڣѷ��>��U7�>�Ս�Z�Md�K�,���~\u j���̈́, ����o1�n��!$*p൚�q��9o{�s�:�#[EH^�c��u|&��!�bz,�R��C�e�ŌP�__�,~�y+�n����gm$T��0 �N�}���f�@����O}�.h��$����9��r0k�����ε_����L<	C�+�~/V<�8�{?���/޶R2Jqe�����29`��Oh��E���ѷ�L��q�T�Ϟ��]tg=�o83�ހ�f��
gQ��1��g���T��)��P�� �dݼ��5�|��(��c�܆�g�I���槻��k��54�v�����1+`Y���Ak�1�l)4i�}Z4��{�J�Ggjú2 �PX&n�r��y�ɪ�(��9�C^��?�%Wi{���#uc���*�zɘa�<+�nux\ֲ�;g0�eGDS�ĸ����Oq����A( �ƕ2���n�����ܓ���)�����v��u���u�m���l����$�S�UkCl�!&�|��������/�-�궕�3�H�}��/A͗����3T�^B5y�=�� �����{�0G�'�sQQ#��i,��
Ü6��?��'9��>�`�f3\N�L�Wْ�P��f��r܇��W�ʧo��a�7Ma�iW��K}���W�ObGF*HX�v����7Ȫ�q���8LO&S�S�j�,�U�aF�����> c�!��3��=�C>�X �.�V�xt�:tځ����ap��)uP�f8G�X�b�����D��`�ԃ}bQg��q%�[�>L��X�s:��=@�(��|u���1�[�5��ڦ����[��3����5�Z�f8�Я�ajdI���x���ׇ~_�����)-�"�Gyu��;�[�Aq���(���sOߡ6R��0K�W��KA=������>���u^*��$CJWȤЫ�G���4�ȸ����������7/��z�^�b�L�X�|�wU3��c����e,(]�|(�<{���uDcy$�5>h� i�g<��x:jV����Ti���@���?^��B�RM5F�x�љ�=F�>:�z����_��n�Oz`*&~�w=M>���6�k�rS*�!v}k�v��H����J�'E���>�F��2e`�3y���k�@IK��\��gܐ!p2s����kӨ9�C����1��_V��S�W���YR���]a��~���.��W�	3�2�˼�#M0�H5�R �{_�d�5�7��f��H����ړ���:S��S��v���)��[��.B�0PU,|
�H�����=m޽�G�hv������wFX�j̙�O˞^�V�n�N]X[]H0��O�b��I�J�hj�p����tLv��@Z9�B�i֮�f$VK�\�B��������W��OK&#�Hj�G��c��w��7	v�a#I"tϵRǞ����J��w�����o�Wk�:���g5R�*����Y!�M�ē�s�]B'�$,���z/����Pay)������<����d������U����h댣D��[j�	2ޏ�/{��� UAԃ%��dFf��<���g1��H�%o���]^����M��4�_s�R3�5���^~�n�7l��5:��(ƈXhD�h��;���f��Nh�D�R��6؁��ʰq��[�5X�q��-z�����`M�4֪@��DZ]�2ĥ����v��E>#�@�do��/����^�u�$l�㮂*g��H
�V���Z�ƈ�j@�l������� �N�w0Ş-��l��Oq�
��ǲc(K6�!�ey��� K�3�[̉�16Y��h2�!�f��ʳ��0��5�2״s�����^�PG���.l�.���n���v��ҍ*X��m����S�T�/��l��IJ10�3�㤿$�%3G�Xa�.`�bP̘�)T~�'�ej�D�����F�T���Wà�>h����ݦ�ًo�T�ZZE��|��%DD�8u�>q�ě�^(J���/��UDe���ӽ/O��BC��K����������%ŅH�=S8�c�JNg�4B|�~�U5��P)?C���٩mC�خ@�
jˠH�SѶ��� �W�ǻ��m��������k,��Ļ���]���eor�[�|��邢��V� ��^�s8,yghk�D�#v�B6
�I�E��Q��;��H��U얕���@g�{˷{[��P��uFJấIH�2�u*�`8�
ճ\�^ "s6f�# �va��0�g�Bj����V���c@���L���ؔO[�(~��&�4v�S�v�)�U��	O� ײ�H�y?�8��q�)�N�����*<�M\5E`�ɀ�ͧD�|��&�@�$�ku�@�f{�l�D>^��d�e��Y�I�����󸐻��]��P�8�(���� ����r}�8׌�J�i�b�v֦�_��_7��T��?����| !��l�ɷ�fI�c�n8���넘_����e]����YYN?�=�3c���$Ve��u��B��z!�@����"�V�u���g�o�T2'���wkwM���Qнe2���N_�B$�F���/�������I�?mR��]���EN0��׽ɏ���>��� ���3HqP��L� Od���`]�T�C�GPW�S�U|�s���o lb��E������~(�{����n:x�"o��Dk���͝��	�[�S1Ͼ�|�˦ĕ����߮]8 �@���K.�wy�O"O1��c��11�|ݖ���,uZ�󐎼h1�\dG��ݑ����<���:�V������Հ�.���Ю������1��U�+,�4O��j�G����[R�����
��87�}�Oc%m-$�=z ��������,�܁%[����K�0�N����N�?P�$�↱s�{������CP�f�d��Ė�'�q���t-��F�W*�ov�L��PuI}�;��*3^��z�A!��N�xm:��(n���+��dK~Vȿ,�\n����:��_�`��@�GY�����PvCz���5��!�ε�r�����D~i(�4��#tFnV�Z�	J�tѣ3f�	̛a���l��,���}�]�l4���,W!�\P�����tH�Em
�4��Kh�@�hZh.FZ���9�����	Z�J�AS&��=��_���ϥ��� n�nЦM��H��y��4��n~�X���?��>��G�}������ҵ0����{��%`-�^]���d��yL�<��JM �-�d�n�@ӊv����K�A'���+H�_<���y4n1C�`���UC�gP��Ā|���`*:#	�����QsL�|~���$�0,̲DLZU�8g�`����tF����1�����d6D��D�	�y�G��bɍ�Y{rk��6cU��U��F3)w%��� ���`+ʳ�:��AB������R`�وBJ�Uy6-j��T�7�f猡����^�l=�4�RT��v�K��	��I��\	�m��8:�Oc�~�i�s��͝���:RuA�Y쁥q��UO�4(�Lح	�g)���`C�����y�=Ri%2�ؙH46��/�(+��h��J9ډd��Y�ĺ�VW�62d�Yk6�,`�#I
p��[��W��ifup�ci��(�Qȱ/j+��2��6�C�uzϬ��X�ȩ�@�Kʳ��Z��F��ݚ���y��"YS�o�Չ]�)���@�T�����_]1>�9�]��d��ԋ$ƿ}ߢ%�4�VJx��k�����&c��X�q�cO�)��'Q����T	��>1 lw�b�|���Վۨ�3�W���,ɜ0����4H��4�R��x6��W��3}��a�e���ZJ�Nת�켶�����1.��*�&i�bq���n|t��6��$���g �)-Q��A��"���eo|dɹ�����������*�:<N�}�c��]�kLG5��L�s���W��c20|؁��}w�vF}B�:L��)���%B�*s� ��K���8F;��{w@|����$�ln����R|�<��iG��38;`"YZ�1Ze��6�[���F�N��I@�]p���K���C{�5����?�$=g���n��8�*�������@��_��ZYq��C~�%%��^��I�j`��/2���y${ǣ7e���� �[I�vS9���׈�xk�K�Z�XF�##@��
����	�}���:���� ����d�6��>p*�V���G&v�мx'�	�1#.t�%3��ΜaPQ��x��n�[�XX�=��>�B���W�ǈ�TY���ڱ��Zw�v�r���IJ1^�:�
����%���=ݖ����U&D[�����s$�d]����n���x|#mHTv�(`*��û�.G��l�A���_��99��ߟ�>�"�ʯ�=��b���������_��l�{	�D�9�8~x�Z�!�A����ˎ�M�J&$�d�ܿr	/�e�}^=08�jz'I7�z�,覡� ��t���Ǌzn��zD�8f�����Wo}<�B;w�╂�jW�iWHE hF1�1�]�<��/@!2�i�nډ�a�����%V��rE7��1�B��^m�		�"�%�����_�SR�qť?�P% ��Q/��oB[�4���J��%�?a#���1��0��$-z7<��y8XPx�8C8��pD���4�/���nhR�u z f�t�%ĝ[��xR=�4�a�=�j�z���ӹ�X�?���<�b�͍}sW9�~L�Nd2;�8�gK� ƨ�圆Fa[? �)�+G�K�)��R7��g�Zm�ﷲئ��C�Ë˻V�����#Q��C"��U�C���]DR��Z�}���W�	�#�8��)o��X
ȷ�=�>q$E iYm�]]��7�ҭn��R[d��>=/Q��3��GsYsr)�W���S�JZ%?=Q/S;�vv����y!f�*��'���+f�O}Veә�×��)���s����P���9��DC�>�=��T�[��JVV�j�n�/�vj���H���˺�d�<��<5sTsX�����1���H��Ontd�*�̠��R���s	�}��Ā��J|mav�_������ؑ�pg�|��YxV���Q�ఛ�7��}�3�����9�|�/��u�r�_�<X�N�kc<�lٵ��#H
�x�?��B��A����>�M h��C����� ^{�W.Z_�M�YLb�Q��}����w�%@�Q�E�%�I%�j��8p�U�R�䨫�q��``�{~�v|Ŵ<Z�&�l u���OT9���7Qp����_�w����v�=�MLfcbm%^��[+�3�](���W���}�P�V��0��ZFϓ&��$���Ht"Ў9P3Lj��apZ^û�m��� ����5���(�"�{��"L6�YKf���*BHH�5�dw��]�C4T��iU�o��yw����t��E���9��0K�nS��˯��v�-[��Bp�M�-T��h	'����(b�_Y#]�
����f�' ����vفU>����=���N����X3�R�v�L�_��2���t���C�h�F�|�<��֒�"��6װD;<�Q��{e��E�{'�
wNc^%	��cm�dIج��>��E��$��}st�A+V?\<��b�7�,E�}�CD���:@��}�@�R����E�0T8�G1���f�)�u�)U���i��aW
�O{���c�'�?�`P�Z1�:���=��)��!�Jtc���ͩ���}�Zj5��.t��
�s�Kl�h�m09�����{�8������F��������g��}OF��mLҾ.:kb\�`KbM����wd! ��j^�z�J�G�bh��F[8t0��L�
v��,\���]�MȖjv{a7��gK���6	�xV,�gA���,���ޭ�w4W�Q(�m3]Я�~�Q�p�6tcX���C�:�H�<��L�<1$�UtɑR��3wC��� �a�u�2z���ۑ;�W�WB�q-Pi��	��2����feh������u��k��v�+�k��� ��`�(��Qn����rN������9U��#��?�i����"�(~�U\��b�U��.�b6�;4~�l'�E��j���I�Bv��׹�t���׮(�(�������u���?hA�7�$(_YU�����m�g�^XV��˦�`����ZR��h�m��2���g�.[n{�I�������Y�|�K�t�˔'�Z�����*�;]�Y��)Oe�\kL#M ai�ջK!�W����y���_��`��+�uW��Ξ2�*?�w��[�E��u_!R﨔����Y�G�~���,��*�:g�/�:���8��:�Ԁ����o3���s����{�j{�lx���&l^7��Q�?���� ܋n�c����&[}킠�3�UC+����I�o��ӑ�$�r�<%K&��h��i?*]3�n}�FP�_I֓�X,8���{Y�Ёz�f$?@^�D��;���m�~D��v� *G��������`��(��l��G�O��pqt(��������:���ʰt��5@(֑�:�,x�D.76���(o{t�T�E�xA�I�$��d'�:��@xɿ)�ҵ�Ǒ��z�U/	�)쇅�a��m�bs���F""=�h���am�e��}�9�+ndms��B��aү��a���Rn"�o�j7�d�ö}���&��^�3�͡��>��fT������}���p�Qq�V<���,�6+n�D�G�+9�K1�xĈ��VoiY�а Zu�3�� �X���+��#�g��y8�'��V1�;�NAJ�"o2����|0�z��T'�G�i��e��!��������G�ϋ' ��M��Ьp}��v��K��0�]�
Uε8����dw	S�3#z#x %Ƚ�2������b�N6�T���J�}��wpA��GlN���SE-ʦ�5C,��"0���I�ՈYLx�Q��%�L�\���{_��j�@FiL��XVs�_�h���A�\h�T1����$�NU���8�/�D灁�Sѳ:��.��s��u���R�A�Z��$+����3�Y�y$vb|)�����E�$����q��`�6�ͨ���$��0Yd���g5i��X^D��?8?^G4��TA�=�@� Q�����o���y=C��ּ�!I> �<���Sh,A֣xd�
�>9R�mU\�8�������]~��A��0�����$��=^�m�c�dmUyK��Ҳz@/����Y7�Xkω��A�kF�@�=�&�Xj����N^s�|�i��J�j��s�i��4�r2��K(R���4^e~ K(�7��B�G~W��!9R��V#y&t��8��=E��%�O���]VY\z!�!t�{��c����?��'��:�?��=��pe��n�(I.,��f,$��"z&�=�z�;�J�-m�%FL�H�����Gc� ���ot��[LJ���ok�@{F�F}W�j���9�<�N\D�B4lf�M���c9��x�7feɄ�<õ�e!
�}u�mn`UE��MRr��״�(��\�ϛ.�#IVk����53��v��
WϢ��a���1֨Z#4�!�94YU�uzZP��*�� ̭�:!��	�ļ6I�!��u{� b�Q�[�O	�'"�Ex̔��`��S ����c��#P*�H�`�
�̷�����m�J��3%`�'Na�^2�Jn�P����;�D-^kkwX���3�>;D�$a�T�����M�[�/J�s�lH��z�����Ξ��`�X���T� >�����#������zt��	3�p-a��Me�m/���ON�Swkt�"�Ր��}J��S4�$�H��j2r�y��Ʒ� ,2jx�c���F�o�d�p�ܢh'�Q�"&��k�2�W	!�4yI3ڃ��ƅL�c�rO��f� ����Y� {�Z�����ֱ�.KG۰zD��ym�>��۽����t� �ٳ����"E�����'�x����£'@u�f��P�5h/Α�X*Rl�ݪ�SKl<�*�~�ꊘ;@��B���oQ_������O�)����ɛ
ڛ�Vf����w�vlܘ�m��A�p��f8�p�n�s#��ğ��a���q�p���!!~O�J}/���9;|Y8�+:�9�BO��[x�w�(z�����7ل�L�3��֤�d�@�*?�����"(������e�=�_#�3LC�՜؂Ӿ��G����q����p&Hu� :�ၲ�"q�Y7�K]�'�ļ�=W�����g�6rG���._O��莉�'P2�[x�ز~��⌸`֔jn��Xy���J�e@�w�q��F 8!�Zc�xo�x�v�J�1b����}��**�����ɽ�YX`-r�hq¦cI"��]_��'��@r���[�=�񕤣o�~��:�1�H9g��~����MZ�D<�H�)9�#�j�P�bJ��:X^׶�������Lx�nm���V�$*{��&���
�B�
�z�,�p�"��o ����E���T6���D��6u	�;�o&��p�N�톌�8l#9@�O ��-R�R/>ǯ/Uڮ��o%�#�20G.A�ԏ�}A�ȗ�}c���;�����a$V�I~j,/�
�O�ݞ*~%_�2b�R��ț{l#Ԁf5�&����Nb��������8]@�`�| �aD	J`���Ty��Ur�V�K]��N�k����,�,!1�i�h�~��_�kIs���/��[m	�S����(�<MkE��9�Z�դ��~��_�N;#B��x���!���ֺ�/b�ͫ�,��C�jG�4��3C���6~C�Ha������<�Q�����憘heD��-����	��)�k�V�r�:З����Q�T�p�UU5��$��/z_������h�EhI,"�S��Ͷ�{���$0��>À���©�3#c��#��h>t޽W�-["�F������ۀ;���$�``<���������d,q=.��E"���,$-_\���}�O��j���� �ba ��u�%�7?�?$D�"�I�wl:?���3fK��:���҂n\/R��?M*x�(�Z5@b���$t͐	#bӗ�o>��n??���̍M���v�����4��]*Ta�݀r�����UЯ�	�)�.
���D@Q���0�Z�LBf�J&����PiA+���Gzr6!W��w'f�Jp(��L1���@ɉ�",�y�P��jGe��X˘�p@��-�F�ǯP����N�yd�����P#���ە�=ʱ��A�ɛ��Ʌ��g��QäIl�a�Rs�>�J������o�4�K��lׇCU|rQ|�b����l�z+Qg7��g��̡�r�N�$3�,��TIZM�у��e/g0�XI2~��*:%��w��t+�,�I�d���hAKމ{�2��T��k8�l|���b��Lw�G� �8[��3&B}�^͌�A�2����%���oF���h�����a+��{��
[�����*��*AHH���"�|�W
�r���_(�Hf�pI�Cs��^~F�9st�p@����J�`�]c+������
�3`	G�v�)�R��Rv�N-4�$O�v�
D���ި�6�cgCc��kD�8�]�(�i��g@�ix]/��,
�K4�s�t�meY�^�mP>eȾ��]�Y�������>��<l/��z�*Jʴ�E�l���£շa�=�ޓ7�f��_� v7J��^J(?�#��]��n@pT�8�ңh���?HP��q�<jɁ�j��O�b�U��c.E]�{�>���Y����O�4����V��V�t�~y~�,-�x��HSsH&�Fe߄��0}��/��Jl���wԁޗG+�46[���b��~��ޒ� *� xGϷ�bIN��n�_�s0gW����,��Ł��OQ1��^K`;��r��?��Ἰ�4-e�%�0��3Ѧ_J ��z���o/�I���v�I ��p~�VZLdJM1�ȡ���|�l�_gڎ��Mt�i=��zH�!���"@�U���B�/�$ix]t�a��v�1��?.����"���ּx�r�Zz����s�t��E��P�n�Z[��s�:x# �b�Z��V�s$6��c�,4��3���A�檇��*����P����+��%O�*i�p�R�D�v�"�w����㠬@=�&�v��� ���M�|��hζ�X_ �� �.-�\�Ggn���cj�[x#��k9x�3-�<�ֹ�fn8���1�σ�Cu�"��S�a�Oh��������2��&��d\�@�^�7y	�Ul-R�`��H D����bT��Pj\H�F�:��x.u8v�{&;��g�c?]���� C��e�]�|J���@7���S�(^�ʊ/����a)�ދ}�&�[�<P�L|�u|ar����8���a9�����h�(�����d�o5��I!���$H��<SQ�-���R�	B	����t��麘�&��b ��>q��G� ���8 �<_G2�J��)��-�BtLe/[�_��1<�G����д�?��ҖtǏͯ�3u�"��0{ ^���p�f�2�� �S��ޛ�ŭG�ѵƇ�� �^�
���Rx3(�_Ctl��0d����f4t����?:�B�4|ә�Y�c�_��e<m�$����p�]��4����}�a;����>с����01�rLJ８Β���2Ю�?��e��%ř���V��V�-��wJ9G�j�u�tH5A�ޮ��"�E������xy8��>nw6/C-	?��)��gx������m��G\����Iàhs�	���O�8����n�e[E�-u�d�G)�s�a[mx�������B?��vr�X���HbI����0��=L��_\������c�l7z�K�$���(`�7��Մɻ$~�ar����d�(<u&�r���&�H�/���V[岿n��1��s�Ӈ�D ����<�s�A�]F�Q�jP�Le�C�d�N߉�/�)t�ڜ���=s�5w!@3�6<�o&,JJ5Ocg4�ja��\8���L��D�ގ��2��mba�R���r���na\.7�Ԉ|y�����x���A�u)x�����>��[C���G�z"��~��#:������.��"W0�������r3n�Ɛl:O
�l�
fB�~6#3���L^��l����u;_X�T��+|,�uM��V��@�T��=o�����t+|C� xg���b��������&h	,�;����d�ހ��W��PwB�>��@���z��&�E��	��Q��(�Jyu�uxFo�#�p>ݳ*�a��Lx�P��S��	I�{�E>��X���hY�})�D�*;jBB�g���F�	%|�AqXb�?�@g.6?�OI!��}J���8��f�� �#`��� $3x�oa�j�n���b�M�� Ȃ�	���H�a������v�.��i�*��{�|KC�#֨	���������e�]�OL�2��3�kSd��\3�O;��,-�^�td�y�,��~"��iٲ�6������?�s(�D�������(	����d �����.����[��e��'���3o�=I��3d>~.�V�:Bz"�8�w�2ED[B�D	qNV虍��8G]� �2}��-�@�:	ؾ�&��P
-�N}㿩k3�Ʉ��8B&Ύ���~c|&� :�M�� �@�<��Q�ry��26G����T^��_5~��$ì�rGgj=�3���3�H��|[�:���#x�%ꐽ2_j�"����C��"t�*=n���M�v�Z��/��_��
���%�IX���)y'=�C�G:�p�#����Ͱ;�q}��O���w/d}5�Lz�CO�kSK�b��t�����F�F[��u:D�"Q�q��~�&iY��|λND�H�_���Vq-?�f9�_�Vg��Y��J�5w�,=�'�%pP���f>�i{hK6d�q�]��&�6��dO���ν�ܮ���<�;��Y��[(�O�C��G�Ց1��"�+4�0�4��1���go��e�|i�a���UR�p X�Pb=��}2�Ql"�R?����|�����!���xF3�����U���Gq����M�Lܙ��Z�с����u���'���n�̷AU"��Tn��Zb,q��̦0cǞr�㌻�.�a�MV��fu6������an����J/��L�>�~�ˌDw0D:�9�� V_٭8
^j�鑑jT�I�̹}�RU��h�ʜtP��?��ӥ�%� ��BE��C���"�����O����"%�Z'�a�k6�
� ]��`�xs�X��_�+���&-�h%�����g��RѺY��}��B*�u`}]&��|�ͅ�i4�U�zZ'K:��e$}�|&�wL[����x�4���к4X�L�&��Dԉ�ֻ/�EY���JXG9v�(�Kr���ʼ��G� ���[�I����$�Z���.O�����|��6V�x��[�l"��j��i�R�oP_�)�XG-vȞ�~k�h��}���lAN�:F��78}jT�[���x���傍�M�MۛU%ܝr�V3��M6�.�h^|�q?y�����9ly~>x�&�M+O%9��ȑ
#��{	%�y���?¶��GM�������+�X:Mqf}GiK���y���4��S��P�#�G�vo�G��0�l4�3�}-�Tl�nB/�u}�~�̟Ꞓ[Y����'�I���s�0��03\5���`O{�nٟ� �'5��ti�,��h ��k���Cu�wUu��)\��i�!�5v���{����������鋇��R�׸���߁��A�4�=�����G�%� �}�.!160a����@��};�@|r��\Ty�h5�����#����i�)s[�����"�o��i�/����ޑ��8*�l�g��Z��S@��o�oʳt�ܲf�]oh����T��<A��8G�5�\�؇�{�x���g^>�e�o�+0�5��:�<�S憳�����]�K���ƑE_�F�m��h�+���I��Zi���7���av�NM2�|����� l��'����l�^��{aуh!�lU��wӻ}�rD��g�a���Dn_�x�r1�S.~�B�e���C�����(��� #�{Z������)0s���!1~Egզ�TJW^RJ�q�W�ꈼ�AѺ����*�
�{�x!���`^�"�#�g� [�5�2��^��0z�ω�Jf ��?fj��=�w���'I��>zX��|j�3 P�m֞>E�l���`�P�b���F����RfN'X����s
����� (�����F%���+�(W�n�7g����J-yt��Ld��1f��Ѓ3"��Cġڤ2��|�#�L��c�CĈ'�l���p�M�;���#���]0iy�?�l/p,�R�������i;�~s�-�� �v�v�vO����
!�#�w.x�
��(l@�[�5��d�b�m�b6QsR�?>�2wM
L[�}6D�m�o�U9!���l��Is%t�p��)M�O"���f��MTa{r|��qv n��/����:�d��^dg���KoL��* ����`C��WcءZw�x�|��r2P���b�8����tGbx���H����AL[/t"��0:|gQV%�h�o_�`��'�P[�����)����k����A�wh����<8��n��{�`�B���~M�X̀
(g�|@�1�6W�aH�x�{���>��Ч���xjR\�:�H7�F.������*����nxY��ͻMr�����R8�6�k}%�%��! �CNr���b?���S���*+:����V�R���D�J�T
G�z���
f�����gWć�� �[�e�b������[���&�Az�a���u���riAi����"ɯ�>E� *��t@��E�a�5x��Y��䱈�&��>�Wv��z;W�F��A��+x�v��Z||F6�YB%��2,��sno`1��P\|��>��.�=ޓ-5Ww�R�	�]*�)��D�b�N��ʖf�(�������G V��o�ؚ�kV��O�q�޽�1����}G
5;�=�,�P@����$V2
#������+C�����$��~k�o̖N�̛hL-�`��1�5b����^Y�H�4���R�u|�xƳ��,������u�G��n��,#ȯ Keiz����9u��>ѹ	�h+��r��]�N�M�TuvX�	�9તC�m�<�g��i��6PHkj? Kf�ˣ�:i��i�0�{�}VG��M�b�����2Yh�}��Uhج-'�z���:��:pp)�.��,�[���������\�["~9�����J�}����J��f�KY��P�@�B��w� �su�����n���Jd]/c���\}��.����������u�0޵P�;]LP�V�/���#��	{��T�:���x�9'.�{_F@�1�����N�����d�E��� �~�2��`�K£���)�7Nf;
0MQ��s*���Q�E]M��������27��>���(���!��V�ا[AV^%
ˏ j����Ε�S<i&	W0T~#��_p��FϠ"0������SE�$�c�Wb�0$4l�Gb�|�ћ�x�3��ψ+� ��أ_c�Q���uq%fՔ��/h��r�T��7XH�����Ǯ�w�G���{Y ]"��6<�3�}߱�v��=��ry�1Wl%?�M����@{�<!"֕��v̓��)�ユĭ��н���̺Jq���QrY��4��C���6�.����J�=lN�#��ȵr=��Ѯ�8�`�x�i�ԃ����.���ZxJδ�ѽ-�M��T��6������G�rŪOr�V6��.J��tԑK����;H�d~b���Sm����?�����l����8�2{2�� �3.p���k�yD1"r+�4 ۋ%"db������|0l�׏я��m3��?��N�������(Uy��K��w�-uI�	�e�N{�|�蟀q����m}���ԓ��VYS�{f����N�ꆡ�t�c�{�+�$��Oͺ{�!?M�����e"�_��:_�8��3���f��+u��������n�:��S�K ��i�o����Ie��|5���é-[9�ά�>'���m�/5���"�4{�<SUF�Si���;�b�j�8�JF�>Z�Yt7R����a��N��"��h#������Ss �n`A�$���V�Ő���z�tp.0�S�ƆkIH��C�Y���ݎ��7�q����~9����&wل�F$��=�c@$.-s��}���˓�|`EȀNQ �>%ϡ4&��Cb�X���%��oRݛ��F��OJ� n5�By�ɇv"> m�Z���n������n.���*aߺoA���8�h�DJ��X�,��_�sf�`��K�r���cH�.��@D7����Ә"�#٣�(��R�y�	QxK?��Qk���If_D�-D�<@�Jz�!f���a�B��>���#���DiQ��f��X& 	kNs�utJ;8P  ^�S[m;�=7��]p��7j^܄w&\�x�5��e�8�0  �������Kjo�tr�'�b� `r!���š��$�+�(:,�$]� ׈����<�!��QS~m������8�#��������֐Z�g��=�AO���rY�#���K�����k��!��Y�|Uڰ�3s���#�W;M1��D�
j��(b�M ?K��S�}'�w��h�H.1|��'��:ܵ�(�ۣ/X�e�&�<�͇��x�=����dp�T.�����a�t�(<�<�i�����_�������G�KH�+<t͉K%=?�A9/E�.���1bg���Ҝ�����BJ�G���Jg��y�r����3�p�<n �h�}9�̀c���-el*�\�[7���o6��W��.3W#��$��Ǐj�i�	4\���B��b��0�!�k��>5��1#/�Z����Ll�I�ɥ�C"K�L�A�VC��k��L�~m�d&��,��9P�`!�0�Y,������Q�1��N=�L���U=l3Vv�_$`�{��%��`� �Lr�(�0L��.Y�l�7�m%,������OB�nBa����>\�f�x^ߪT?Q*7�XG��o�j�Ծ�g0�[ ~��f�6���5��u�VE,�?�u<_*�ٖ����n�D�^��>d#�h��0֤{wĠ7R
�0���/#��X:�@ɏ���n2�r���ƥ��Je7u~�N#��^ݕ��XF]{�][S\��hҺxټ��~�|E=g���:��W�y������P����c�tP���N[�^�d�_�9�A��_Fie��#[s�7��y�;7�/?��FU��\�����3�,�ɚ{Y7�2FV���]�8�^����tn�b�OB3ۡ"v��
�b��}�a����:^Q#��nf&�_�ER��&X���ݗL�5���fd�u+>�t+�����{"�VQ��2�/R��Ok�و8�:]�c�����ûk�?/X��^瓗��)������I�فW�<� ���0��t�(
e*S}�J���+~A�v>�ح�ۧ�i5E�'@�,U���h������]��=��7�\�Ъ��6Y�b{	"���.꿲~�4kZϮ��oJ"R�C@_�b��O?r�x��T2���nJ��q:ID&�0ǟvH�
e�>yxaXp%S��]�vb�X�]c\���ep`��hΨ��A��u �@��ٕ�F���&�W܆q:A'�b�H!x���] ��j��[2���8���}� �T���j��NP��CɆt��P	�� �ݫ>�b�{���J"K�^ _������S%ˍ��]*����X?#M�P`	��d����H�@�A�,���δ�GZ=O�;�jt`�L������Xc)�t�>��Q6����1>Zc�x��t���x��Y�s M`�7���c��'x/0WE�׻��2���?��	,uL]�Д�]rx�Rӗ��j��2s'�+AÞ��'W�߃C��F��{Gl�g�Ҕ��;��B��֎	h��B1���� {�5:ɳ�����~��3&t�_���K��,��N��g�T�\Hy�kPw�s����:ʐ|J� &���Y�:/nJ���� �ج{I�
筑�]^�ͤf�>>5���r௭M͡E_Ck��Y�۠8��\>F����)o ��P#�IB������;�j�w�lKwe}���z�q���]�l`~�9��p���NZ�/��
���(A]�jݺ�H�t��w�3�Q�L��WZ['��� �Q_�$ά;�?DĖ�Y�
�<��	7��گ�~ac;E�+>�+a�X�p�C�=���|Є���ͧ)�g	I�TԞ!U��;��D�����M�X������I#�ŶkfO:���4�X�����8�Ǎ��Vr})����7�p���p���f{���e?5�J�5{��|n�u��q�AӮ�������	~	�<�r!(�:^�\�$xW-%��q��B���j�&(�ܐ�h���DG�<`;�_�µz��a�$+�=���c*C��q�*��W���9���xY��2l�~�q�$)ᑸ/>Ad�/��v�.���:﻽!�G!����8<���:Um
K�?�*�U(����xδ��nm�e�󌤀�u���W�g�u2C��o)N�yi�E`��F3h���.���	��:��j@Ou|)5d��S�	�=+g�[����s��C�f!�v#��������F�}���E�5�fƚ���Q�����9�{�@����\�&���K54�a���co����}���a#�+xf�\�� P��6��Y%�	 ����D}�iC��(��>?�{F��'��>.���ь+B�ړy7����>���u՜�H)5Ĭ_^��L�-Q���<��߫���㣵?��:ͧz�rt�8���,��_I�y�!"����H4���"�qI݆�k�G��Z�IK+��{�CN��Ѵ:r�I�%[�E�Y&S�t=�X��(6Z�ѱ���S�t�U��޹��y�"zm�h��|)��%�ђ}�E
}>1o���z�4 �)�>��ҾR�HS���h�|�li�t�r��U�+��-E�s�-F"�#�����7�y����	���8[�Hlzyoԧ�_|м�
���q�5����
k(�<v��Ƒ@���xՀ%�s��-Uـvɮr��	�7�6�)���}���1+:{
R-�)�8v��ht;;�L�-? ��['�qEyS~沢/
S>����ܔz���@�ɱp�ˎ*w�y0��0�0~����:�� �̽��f�qm˜PSi{����޳*�5��Ż,x�%No�]�W�̎c�pt��-X���'[F�	Ȗ6c���Rջⴥ�pU<�h@x:�Y@���]���Qտ�Th�Ŗ���h�Ie�F�����"�j�t	>c��3U�,jr7.ޛr�Z��+�q«8�������;�pG���<>�_}�;S�U����H�yRq�77�P��\epmWv��:�O8'����4�U=j?�b�LF-�f8���Z�4�;�4f��4��D�\
�ے O��Ɉ����(4P)=��OA��U�X�E�dt��C$�h���+E��*�J��L���/��o���������z�*UA��a�V�d�ggLL;��[�rgv��oFR��/�Fj�|��=���;n�:�8�� �����У��IZoa*��<P5W��B�4�����4���O��m��쁆�� ��exH���r�~p?{���_��۶�Mќ��~�-�}>v3
#:������!�Q�>�h���V*KtA@X5CZw ��=�D��f*��߮#UO`K��ٮ2y\+(x��o=���y�|��G�-�c���J@:�70'y�81�nY�;s��"{CU��sS��W��
�|j��Ѻ��8�{҉� >�A?��c=Bͬ�e3��1 �s�ny�"��ZB�ٍC�Δ2>�Gi�z���Ka֑�5]�u�e�~żz0_�/�f\N�wx�Q��_�9������.z�cb��͊!�j� ��y�P�a����⇢$��Q_�rP�[ţ|��9�|��1�>�C,����B:�x�&�*d�&p:�OX��<l)W���哾��y���r���r��Tv��z�_��H"Q��ۼ�N��<�Qsy��ky�_X�& T j���Ȗ���!ռ𥪢���.U���� 	���V��<�c��ǩw������MR�v�r��'����+rI�p
ɻ�E#`����Э?��=��h��s⡰��9�Y"��g�xtf趣>F�����/3u���S}�LE��ǁ=���ø��D�P����
ɡ��&��fӜ��Y���02�2�A�qw�ϫ@����_Y\��a�H���|�1����Il�1<�niS0ؚ�y��������p �b���O�ҷ�k8����e�L~߫��7���+w��E$���\����̄�J�rZ��+�j��Z{�0/�=9�럛a,&ϪLV�'ad��/�S̈jsټ8p<^�L�����~Y1����K�'��"�<��1Kے��M>��W�j�}I�弲a��U��	G�k8�7m��J��z�'�VZ�s�^���4-6��:�V���o�S��`�� c�����6_��&���T�8�=1b�I}�H�*{^�'����d�	T��p�� �\�		�+�󒫦ƖN-ρ�oҙلl7�tF��U��ͤ�
#x^Q�����-|S�<[�����K��m9��-l²�W�o��O6�⼏ո36��z��}�p��u��Dh/�]�7�vA!5������3�$fh?{�3�p����(��Y�y6<7��*��F�6���|�֜�&שY��͙�'�v�m��;�0�M-�T1v���;��a�sb\���̦�b��l�$&������d�rb�[�zȷx������S�Q
!�>r��B�Y�pQ>%~��&�/�v��ov��ls��.j%g]~U��!�J��$���H�p#&�=:F-��oFw��:x 1H����Jj���)�!�U#)om7�4�y�;Q�ݶ�K�cʟ3�R@ձ�e !�ςY�ٯ��wW��7�-���Csۏ�MN��؆�����EmmKn���⃣ί�Z<2m|0����a%i�����]�=h��y@L�IbR�HY��×��{��ߙ���ZHOy�g/�٤���h��g dk�iG?� ?�}�'��Mҕ�^��!�A��8	�g*q>35�&�����ҀMXy.p�e�3�|&_Kk�� ւ�'��bm�|a�Kq�.�,/���J�"��-!�u'�F�����ؐ��?g�����Q2���<���c+!f�,��uK�Wr��x؜U+j�ّ)������l�:]��]����y�]����qmM�J$�}��
��NI[�`�å��D�!Q�C?<�X�Y�� ���~E���_W~�S��
��/(�-��n�T<�� L1D�},k�!<"s~�wS�� J5��$��z��ON��"���[������O���ʫ�$�&��6��(��a�S��L'�	�f�ޒ����Ʋ��֖�/�w8�p�C��x?�d��}�āb�
��1+j@��>�L.j�������C���y�c,/�z�$�k葖٠m�~#s �6;���+��:�����'�pD✪Ix�_�,��˭�G�:P��(w`�>�{Z]%[�޵φ�l�uú�V��v̴q��4��![y���i���y�e�ۢ�m|��J��myE�R�L�����'x-���D�|p|��``��b�V�p+��c!]�L�M�W�m��{�f�)�����%*�i�r�o� ��b��K`-�U���6)�H~(%�: C)�񫶛i
����7"qQ��rҁspx��3�	bf��q���������E-6�-�	V�f1�ҍ]�A��z�n�� ��}�|���2�)֡&��~EXR��\����:7���}X��l	&ݐj{aRD��Ö;Q��K���U���*��)]j;D&H ����7^Lb�vuyӯ�� Ƭ�e<��j'>�
E`�;���AT7x�����1�a�_� �:�A�80wN�p>���G���};�8t�O���U}��r���*ݻX`�>�/H(�R���%����}���a�{���u�;���c�j�YmC
�dmY���L<8�r.��MrÓIǐ`�����d�vfA�̬'�9X�U>"��p!�c���"�����B	�ox����[�ˀy��k�(���{��$X`?ؔQs�t�O�YPXe���iWi����Wb��p��u�]���/UVx��B��@��*�,s�PD�J��V����l�"�7��R���7�`&R]^f��w��Ud(�/�:�'e���m�ڞ׃�9l����Sb��=o�<�]�X���q�S�5zn[1��C�����iJv��B��d\)?�
�ph�g�'��1�VRaL�*�\����!����"Vf.xC'������I�#K���� B2|K���[&O��e~p��)����V��'[`ª<Z�+���&�����[2�0v�_!#�6���|NX5�:�3��y�E�į��)D���;��K�j@ǻ9Ri `��M��<�*��%\�J�.���V������&|D�v*�$�pX�&kQ��馲��X�<�İb4p�Aan��̀y���4L)�P!�7�Hk��H�9���,-�7&�0Y2��G�UK��r7R{��5�l��=W.�t�(�,"��[�&[&}\ybO�]n$�3�͹���r��_�����aν���˱�@��Xj���I��Oe�d�(��FL�TUVS����^8sN3Bƨ錭�f:�K�$@�����sۘ�\In~��vO�N�t ݴ��*�xkZ���l	:�O���.rn=�ujB����8���@Urzہd5v�xV=l�����1wgL��#���"C.�����ԕ�L|�5_���n �}6�:��r�&/�ǌ!X8X-������粞��!��/i���/!�MuűY�.\��b�X0�>�����c�kB�B�|C��%��%x� +��,}|zmU��H�)��C�A�����+��1�hhk��8T�H�F��Rl��"�@��W��� ���0��*s?AԮ�ɬ-�݇)�k{B��^�3�M��:.�����xG�5��H�9�����>�m�E��]�/��fż�hC/�}�҃��2<������l�4|�l]&�� ����a��u�8�|o�z1源�N�D�����@`/yTq��
ժ6�Dۢ9�jP��N��I �"=�������VɌ#����빋�[�^�^�R%����[A s�0's�M/+:�CH�
���O�s�RپhJ����d"m��z|l���@6mV~��:�4��T���,?�}����p��bC�����[l�O���|�vj�_$��S��F��O�&s���9��BW;L�fT��T����LoqR�Q�1<�R�O�|�<�E� WC޺�R���z��&��(��ޕ9������K=~ۏ�b�5�x��P4r!P����tjz;�Jk��(�s���eHwu�=@��d����Dc*,�#���)yO� �*TG!'�M7^�s��	�����1ͽJ ˺�w�k�Oʰ%��g�(�!cҷ�Z>L�Ƽ����Og��� �D�d��問Q��1�@6��!Í��+4�� �|�۰R���k�������]yƶ�D�Y�Z���"S�YS%f\��˒4�Wx�ci.ciꓭ��}�x7쯞�S#�7RlϦƂSv��u+�Fbd.1�6J��ifdم�	vŮ�q�q?��wiC��^ʼ ��e�T$=�0`�(�k�r�,��tZ�ܛ[l,�uO�T�Ռ�n幚-tb[���b��-`����&�7��ɩ%(��v�r��3݇K��ł<)*cqO"�����bFQ��/+N�zY8�E�S�@���m|>Q��T�}���rEFޔr<��*�f(�2T�6b~GJ���9�}�AV�~��@M�QM�i�L���  N5��9�Q-��2h��WP����]Z�a�Q�H����]��@����������j�p���v�_)���GܢM���V��	 �!�t�#�������K�����Ei�]$oÌ����^�V��v�O�B��&G�en�=텣��7���G�bj�͐](�!��v���t�(�˪�O��&�	_�J�3@��?�r��؈�"�è�E,�y7t��e���<���	N)]㽻="��1��Z;Q�]�1�Ua����F�r��E�3�q��� l��j��9&��j�M��>��j��e�����`]mH#��6doJ>�֣���^]�jԕ���,A3�"tn0��p����t��mr�����h5B�yY���\�vn���tO�w�t��S��j��������}�a�y�o�9����`�Q�1G���c�.v���De�o��so��țƼ��P�*�q�=S�~o+��q�Q_��{�6�Q����Id 2Z��V������C�bU���a��]��������#!��2�l�Rtۈ�EF^��FI�o���0,�$�)!�ln�`������]q�H��q�ۊ	{G����dÐ0��_������de�_�K8�:�:���p����蔭�o��Ĉ�����s|�ȿ��*e�)'�?�G|�ł�Cr}�|�����gg��i2���������j#�6C@ :y�n$m�g��1�w�=�$�u��H�xoM6M�هfiE����B�v�(~�������q��悰���� ��8�aJ�b��gbTk��;[�1��6ѠpL|C+�L<w<7E\n�]�[� ��g#5�Q�g�v$��W�3�	���oY���;2W�v����(t||,�
;G0�i�k���)��Q��1�\n��%E�k�VO$��}�ܴ�ɟ<ȃ*6�)S� �p ��%�k�~�!_��4�_��]�A�t���qɻ����0�md4��*���ָ[��AAu�X,�Nʑ��h�#�N�֖~�mLf��U�N���虁�Z���e(�m���^��殡�5[F �WP��O�?^C��V���hv�7M��1n�{�73iJ�&��mt#t�e����;�`�go�N�dp+g�����ܔ,�c�8��P��ݧ%#�������=�D��q�����FH	n�9��`�����fA���\�V�tl�m`(nކзU�g`��������@9pQ�Pǈ)����!y������3᝗�yꡓ��y_Q]:�4=q�}�t�7#�A��
��\�)�te�]ݗ�B.{�E�M���U )�2�H��g��qp|�v������Lo�ݣf_�ّ�����h�0���ZU.:c�<ָd�c��͊q��֜��Q?Z�hA��r����waҐ�n�����7�E���'uaqRM{���0� ��aC��Bss�]�8�ͯm�eE��v374�k1�O{q����vd��Jʑ�X"���W�^�Q��|c?\�5��*��A����Tj�r7K�{��+���N�����Z�q�B� Ots�2K��U�����TBi����|��$r���=S��	��u1�p�^��uy����Muj4���������97>Fڕ�F��RĿI@-��,�ٔ�:?eg�Ъ�-Wi&5����������3-w{�QL��"��a��v%4��⾋�5�'/���/��4"�-��)A(! �E�PY��r��e��������{��CꭼR\����՘�T��j������A1���ph3Z��4vͲb��cL
Oj���J��Y�gRX��Gz�7xc3�@��ʹ�v7
1��iE���td����JY
���w�J�/;#�K���i�z��=���k��������z�P|�d��+f��|�Y��P4�S�&��n��z�
���b��s�ik;ˆm
H�i]챐6�/Ӑz�ވ+d���Dfw�4+���uF�x��B���UY��Z��&�~�n��)\⮇����'ޕa�ݞ���@��p���[��\�"���%٤u������t*1����t������"~FH�3�{$n[8#`'�2�����Y?_1��=.�Ű4��X�^<#uZ�_$�����9H�G+ƿcC�9jT�[��Z��>��{~�XY�J(�T{1+�M�q灜	�Ԑ���S�$�ӷM�{���d@�����5���taP�|"gC���c�s�6��B�4��ǽ��A�ū�.|����ch�-������ Op%�p�[L�[������7������Z����=M:�!]U���l~[jfv��c��6m�}��%$����.ը�'���{��q�GW��w��c�8���T ~NqP�܏d��N���z,�[� ��]��ͅ�<~)�&몿`�D�B�Y�uxTĤm�"��;j���%9uH�c�߱�
N[�uԯR�CI�/�!��P@ڊ�1Y[�1����h���A�Vw�������Ex��;5ۢĀ7���\ߓ{�p�1�F�.oy�fq2r�J�4O���|x��Vk%�1b{c����w�]�Lhg��׍��;]�bn�]�)��poG���&Ev���A�a�[�g��n7ZS	Ds�f�|C�[,�9X}����zϚ`�t/l�"%މL?�#Paf��w��@ܫ=.;ˏ!.��)y��\S��?�(��b#$���$�,��	X߈��%*�P'd.�����r���>����-z!���0(�g��5�Y����A�>9��貳uX��o6u4�?ҽMJO��v�1��dÊ��y�t�ٌ�խ�wBA�qW�:ߧ?p'�\�t7?�;R]Wh�O��@�$i"��VdU�f�9��s�]�X�Xxo�~��<�� �Ӆ���x��Gi�7*�������5]W����K�����1Îx𒟮���u�z�ľ�/rM_+$��$����,P�=����֛��C���?�{F:Xvo�.M��Q�#�����7X���W�m}��Z��_,��Lb���5خ�V��?82�f@�Ę�=f���?-���'K���)�Vد��e�^mB��YpQ[��g�|iFRZ�J���������=+�0�Z�������~����ZRf?JLR�Z���v�)�5_��2���^�4{R$
�E�QTkxk�K��?n쏍Ғ ���A��MJwLG,��E^z�-�T�/��=9�<,�ik��Z�R�4Q�g\��v�u�i� �h(��T:� ���
��]��T���L��U��_RDٓ��Q�&%�X�XT�����f�P����Q�*��(���y��<��X=��(;�l�\� �~��;0��D�R���2��!���N!�����%��h<�nɔ\��H�r	A�ɕ� �G���}�WP94����
,�s2~�F�5u�z��FNs�l�������b\i�"+%x,M��R�%q%��CuÁ�6�$\keS�1��\�����,e��q�k��|k��:� 3���q���?�_%�Έ�q7(�3mh�5P�t*t�y����l�U;��v�yB���F����Mk���J�T��"��ί,+�hf���^ՙ�cn����"��x�0s�VO��(�}�:K�AU��tl�Y�
��dzYD��ip�R��(�|����J�kg�Քo�)��*��6�S��jm���9�,,����a���s◉���eS���<�[	�ucaĎ2j�C��_+œ��6#w�|�l���-��Vg;�W��M�UQ���$	{���J˙�N��.���TZ>p�'gF��UVtZ��y��@_��B�����)et՜MA��
J��p]9"�o��G�p�`�A켁%Y������^!����d�le٩���{�E+�L�v6;D���ybxoM�ڔ!�}'��I��8��ݑ�`wbs���&X�O�\n3ή�bP�V
���0{�݀a���Z��c�}�P�����4-�4W�81:�QX�#"�e
cm����hw�N]0�n��ڠx3��r�?;׈�U�u�����gM�,�eE�rB#-���]F���T��[�lG���Y4��t&��ܱ:�^���p!l�A��?�Lk
��4��R:���ߚ�!�@Y�/	?p��4�����5Whz�Cmg��NMMm����K�T��4W`�l�6���/�v����m:��*���0��/0y+#����`�!�6V��/��U_f��K�1z	8����g���V���/��s����kH�B��3��]Ğ��~�e�qsTP]�f�T���VgW|p5���g[�	�ffT�p�Y�*L�ЯG��XÜ�'0½t)�.�:�Ȩq�/�2��aikoo�
��'	 '�[�L��(<��2��cA^E=(�VԻ��3��ߙkw���Ӡ� �n���X[уb��y�BV��D�WTҭ"Ɨzbӌ�o�.T�o-�+��>;E'���M�]�j��:^����Ąo��h�ȉA�����h��OT\?Βm��{�I	�z�~h�?����\�_*�9�:���3�X�	5�Ö�:3��;:������۴@4*m-�R�#6��ֳj����� gǧ������"(�����m����W���=��Gv�.M��7V6���:�N�]z��N���1��X�y�-�q���z9�JbiLj���2��ec�YA �ͥ��BT�u����v�;%8j������zݍ���U�YQ؏��$˄x��d:�,�0]�p�5�$V�q㹢�$[��b{50"/�g���C��!�Kư�ߡ:	�~dv���&�	"m���i�dyc�ȭ;Ҙ�{�N��¾�R�=�c8����;c��>&�f�M--�胞�DS�@ ��'8�cgC@,�O�0ﰭ�|RIW�Kn��=��O�;���/�$����@Q�F�Ԋ��'��q�w�k�2�<�i^4�r*��EV���&-Se�#�q���jv<��=�P;@dJe��e�u:M(����v_��b��5?���= ߳WOW�"hP�Y���V}(i�̞/��N�����η��pOV:�at�^U������5-aY@�$Z�ԉN�
�U�͢���tR�`D�܋s��ay/��Ru�#�cUM4jH�4ܼ5��TI�l�_L;v05��b��|�&vC�iB�غ��|\��)��\�s�TwZ�.�#Is�b��Ic��ܷ�!�������#�ŵ)\-�
� 7`k1�)�������T����x�q����a��_ �
:͌vu�1��5��Έ/W�(s(ԟ���%�o�����?%b�;G,%㊠�@%�t��b�*l�C~>u��HзZw֜e�P����2$
9NS����!P�u��+Cz�~�O\�6����J�gЋ���a�j&zS��D��<�Sh�5������t+x�)՝>q����C�7��L�?�t��M���Ak	��g\���ʲFҡ�����,L\��z�j��5[�'�]g�e\��wu�e_����"��fbᠼ^ST��}��T~�qTQA
���f.���5s�>Vь�?p������[v����'[P�:A�Q�^��q�s�n�D�CQ\o(�q�rY�o�p�W���했�+�dя�����g�B�EP������;�Y�ĵ�ȥ�U�^f0[�����J7�u������B��|\�:#c� ��r\`���sKk�e�ӐC���J�r���G���V�l�<]�nC޽v��V_�w6�F_6��{gׄ�3S��	��7(�$ԩ�%}�EL"%�Y����@��|mh��u����@{�qvʇ�\�j0C����.�j��"_��F�p���=Vjx7lc��*L���|�����I���f�<�y�y|�]�aA�kL���c$5���9����r�y��yJ�$����Y��?��\�)��|sk���^J�ovGϝE>[�	�ө�����2�9z�18#��Bn��)>5,̓�=�hڨ�0�RK����9��3��mx�x)�t�����)`/�u&fP���8י�K��M��;���fL����lrFB�c��o�#ښ۶�!�\��|����D��îb�"�w��Nk�O62X�@������u^&=�bFo�Wٗ�e�'�}����
=l;$��J�7#4�|U����ih��L��0���JJ��s�,u��\��r���E�-=6vK�vO��H��|�ڍ���n��$ڶ�������h��P�>�F�ˤ�O��YB�Ƒ4��?�M�/t�v�'�7FB��ϛ ��gc�Wӷ�ݽ��^�M�X@�<�������M?E���7�q"��a�q�� E,��\�����<�ü������9���y#;RygXw�VK(��w�h�v3t/x��J%���$�}`S��[�u2�F��������v�cug�z���3��21A��a���@�֯>s<`Bd��T�ل����^Ϲ��4[�ʘJ��1�!�B	�
U����+ഞ0����p*gP�P%C���zO�#&�nW�U=�@�L�r�H�ӗ11_�y��y�,p����l�����JH�YP�.;#~�� �[��R��J�F]����4#�� �] �r�q���O�4���E|c_-y?���b3��kT�'�n�{ ���^֧��9�J�<'p+]�)T��X5��,���X<	�+�RrILo�l�f�^�nb�Z+J�۷e�$;,|�h��%�k�g��%�	2`��:ɡ�,�K2�q��˽X#�]���R/��M���I��D�y��-�����y_m#��}|�leo�-O�x܃0� �EL��P-=WV��$Н������O�1< <5�do��.}����=ˁ��� sruP�P��8��db���>������A��;=��6z�o���#[i��m�э�ġdMO�ުG@1���ܤ�S��ݮ�C���s�L�k��'ݻaF,��R�~���_J�Kk�Po~qc�A�Ow����u*έ���Y��z��ע�n�����o�_%�3YJ���*��|8�k����L�]�}q�	�����dEb�+6�L�&�ٹ�g(��YSs-������>�Ȓ��ݩ(�gV�W��[mt�nV�����/s�h��`ͳW3��*Wj������-��ʜ���>j@1C���_��AgZ�x�ugR(�5�����CFiƫx-��!MB�U)Q #κ�ɟ �TP%�^v  �ݨnDьxný C�vNb�� H�*vӥ��������OP��d���B�����:�vBP5���@���蠿� p+��ְ�wP�u�$?��d�"mL�C,PD�͖���T�$��,.{���O~�"��=ִ.Y�`n��g�#kx��J(�4��(��,����j�jx�wvp/@~�|��j�E�o\t��lSyR���D�~nW�#i�A�4V�f�h�!x#�8v�2�2a�� ���|�sDĜ�8G+^���r�.��if�5�-�f�-rW^m;��=�V��^Ӻ�cȡO�<��F���XJ롢,�J$$� �a�Tή)��~44��3R��Q�F��e�@�ʇHV�^��M�#X��CFW+���⛚�!�H��Ƞ_]Wv�: ��7����+HX�e��&��>Sse�� ?��O�����f�d׿���������&�U��R�#o�:���m��0D�G׏0}W8��o�ǃ�n��[���z�i:��N/aݥ��F�5q>��g$u�3�n��?H��p��7_��0c��#�o��� p�������<�L'#��\w�i�ջ���蟿^�Z���/���]C3~D�|�݋�K{���vx԰fFZ!��K���6�KF��A-��I8ZJ`���YNū'���v��T9I�"�AT��i�|x	�����EtI�*D�ۨM�I�i$;��q4�ܭ*�V�;�GE��
Քc�׼��t,�Y��l������i�.\���)Bt��ε�2e�=9f�8�*���'��
��7�X.���s>'�)C�������k ���hq�]G��1,L�F��L���n�D/�ј�R�̦���N<Z���4n6l=��o�����[i���
�?0���z�jųс�.��!&�ߺ_��yYN������h�**�[�j�}��B+`k�a���}���ll�8	˳Ǜߖ	��a16�o�f�	�K��
J�_+�q���mxj�O�7���)�v��b�����#v����n�g��>�ؤ�&7c/�غ�J�����* ķ��o���߆{Bj,��0��ݎ�5��=6�jKS�0[6��6�=�W!��l��-a���]\�'j�b�h�Ѥ�n3x�9�q%#���3�3��0��:�%�Nm�=���4�(W뤏�]�KX���M��ȍ?NAN `W�	�� nFF�_�:�Y��0_������ё3��D���%�D�S'�;_"��k�{��8 J���=P9�������mr��%��F�T�ViV�k�ich�	}��RӃ"�����Et��o8���m�X�e��~	ȍ����:��f�ՌɆ.b1 ���U\���\O5[F�]c��T��(��L˙�J�s,"HÊ(Λ%PVH�ޭ�0$E=<�>��A;͌�P8#�<B�|E�<u$xs��r�|/� � �m�AC�C_�����,˶�!��s/ ��FO-}�r��'I�K�� [n�g����̾-~�.O���"� �� �+�x4.�J���-j�A�j�[�f�)�b�e�pj��PWJ߮3�?qő��� �%>��H}b��'HJW��.��k[��Ni�������ߊۦ3+���:s��>��č!L�)�%�;d5E���:g�9�>�K��z��F���|�X�I�<!���c9�q�-���xat��Q�e%�\�t{�!#s��\�it�F��f����^3��"Iw.�O���5�l�'E�Ҏ����b��k��
�m�.�����H���O�?s[(W٫+,Ɇ���(��7�fW�	� ��|LI7�p!L8�Ȼ�P}G�����樂�� ��ɣpO�F˙�_O�#1 ?�h��Ū-�Se�%�6�Q{���COe�ܞ�H�>۠Aa���@�Tz�T�u�&�ZRH_��=\7�����I3"�S������m��R�ǾN�]M#�Ck�c���,��\>��"���t$#��	.}�9��:�]�麔��>B |1�F�6l�����`lM������ej�M���d!��N;i�d�<��خ�!<�b�yo٤��?���C��)��絿��������}kۋ�POWi�3a��zUj���+�t�_>��Y�?��aݓ�4(Kw��V*�6�`��:7� ���qS3dAQ^qVkaut'��])I�-�)Y���H/���25ҭ�D�(;�/�����"��.x�I%�Qj����j������=4���`�v���(�^N� ���@B�њ�QyS��E'���ҫj��[(��5��xBm���s{u8�&��h��}U�Lw�!�|���)%3ў�~��Կ8���	�����Vx!b�"m�p��P]�}��4q��o���}u1�\]I����p	U�	����E���A��d7E��X/ ��DQS��d+v_�.Q���&��?���|n"�F�σC�����l���mP�Թ��{�5�s�?�X����7��tHD�����}.H��<�N��3��(R�î6˰����d_��+���˧u�Ĺ��k]��Um�K��Jߡ%b��@����܇�|ۘl�}m~���a;�#�7,_�ܓw�0�Vp5]:�	)y+���l�㯔3�ᩗ���O*��z �{$�?�$~&�n[�[o���ef���e�x�ANB�w%p�[ԡ��z{�Q�-������ڢ+���Y.sYD�y�#
�����g�mĵ.B�%t6�#Vtv�Ǭ.�8�:t?���ɶK�M��3G��Ba�K������X���/���5��N�^�/X��~nx�D�h�HR�Oqe�y�5��lO#��g�Y%�7�LD�`k8�.��8������І��ڋS��d���L~�yb�`vyd���^�T�L��1�l�օ�#9��g��hX���C[����fV�r���bԉ���i�
�+J���)�+�p-]>�0���!.ǡ ��WHf���h���Oɘ�
l(����Ci�d8��
�Av���������� 3s�62�=Bb��?��O��o�Zo�5������ϭ��䢁n�A���.�0��/���+���78O'��^�Ns{E
�N
!�E�N���dI���T�K�2�����nR�a\٘�����0���U�	S$�y-[���WQhb��Uիfֵ/��;6�*�):�%t�_A���?R��P��L��]�]�1o4z��Y�D&�\��v��QT[��qi��c�i/q4�S�k��-�V�νց��!!�����������mFڐ0�S�t7����@��l͘��8UQ�4��ϻ�󼞳��&����} 5�[a;*�F����B+�������S6���fk�����+��CǓ
`��~���T5ng<����H��S��C�����w�ʘ�y��p$x,�h�&����僚���cG��1�
���*�������u���J �UO��'w�RD�[9���ܓ��O�A�18��V~��hK�{]\��ϵFڷ��X�˜I�T�#��x�JmO��]��
r޼��c��kz�%�.	��յ{������bG�ֻx%���k�x����f7k��Ȏ[Hi�L����ޱŞ3�����d�}_�[�Z������"M�"�q�W�����UJ�}�"R	�����!Rg���T�:� g�\�߰<M��T.�]B�������
�07���[����-�q�7p�~&)dD���N����j����Tm�Q�/Ǒ)����ҐJ���#�"+�}�W�Q��$��rEF���on�
���-��W����[~�QIf�"�r &��\"V��wOUj�l��@��Q�]�}�zНg���/g���U{�CWd��" ��	�f80��R������)�t`\�o��ܺ�_�P��55����]Cr��֋�5���=x
�T�e��(=��t�0d��i��:����Q�]g�S<��kd"�ć��0h~2$6vbE��D��#���*PU����yN���	��L� W��Tlu�|v����T杮{v3��3)�Y�h����Dg�~�4�Z��zWҜک[P!�v��go��,�;C��D�>�lG�'����M'8"� �eڔ6�X�A�����*�OuF���j(��0ZU�P��1������#�0#F��	���e�p}�i>�s���e rs��g�7�׈���-�Fø4[�m��?&?���>�J�>A��m��g&V�1g)���33�DGQY�h�[�����t��W��R�I���^��� � �~�D�6-#^d)lY����$*H�ݮ�C�M��)&JP�=���B��ك^�KH+��>�oذp��5i�g�P8���'����bo/��b^cu�*�C���L�(C#�\ ��q[>5zP(99�L�K���&��@>�7U
z%)M|�F*[�Q���^y��wR� O��4�U�Bm��H	't�\����:4����&��`�<��p6��Z@��rئ�+�0�A�5 �R<+[;x"v�lf)X����$�{F�n��B��;�����,�n���0
�f��x��f�f*Q�8)2#d�?&�$X������E�r��'�=]t�C}u�7`�vcٓC�������쐀Ar/�S<�1��x�t�Nq0<�>��Ϛq=�},NUk��P�F.�\�N�/<Q�U;���^DK�Rz����I�(BBeN��O<v��Wc�@�E�M�Bgro'iMb_���.(P��@D����'�S�ջD20�<}@��iR�/�H�u��;�I��rB�t��������l�Ra������J\��4��<��v8v��pyL%E����{��=�`	���==��,���A�EH�>p{2 q�tPu��F���6�vN���˙	��j����3��Ctco< �����3T�@��pҏ���W�7�e���``i-ʸ�.���H)��[_�6_NW�+a�i=�lm�4��T$�g�t4L_$�G>��M'S��j�\&�|_�$H��4�e�'�i�2;%4J�+�V���3���3����7T�k7'�X�H3cK�s��+�Aʥ'r�a�w�aM�!��JS4)�&3]���b���1��Ss-����ݠy@��!v?O���1w�Ҹ��c����G��(�Q�>��F�J_���)�� �=:�E��P˽uT��
@`�[�He^���o>�ޚ� �~��c)���e8�2�_��*������j� 1�-�{���[��)91�6i`?���.�U���'Q�-�1����<x�x�^^����2�Qd�(��S�d��
`�0#@|�A�ӸZ���сT\K�k-����\R�8�A�ʝA�`�u��-�"����
ޡ��z����ay?1�g��]i��2�pT^��G�!_Avh�e�3ܯ��o#�O=& =�H轉�{�c�b�GulY�����h7&N��5s���ph�2�b�~�Ca�hD��Җ|z��������3{���Fo�����z�0@�����C�e�;x�4a�;���Sf��/�;�_���'��8�]*��2TI��)Ur?������wT���R6FS����hX�KJ��5^.�WnW+�>�IV����f��%!�[�a���xj�
�S���b4��a�b�� 7����H$GFR������׆���C�*KS�gJ �j�ju�t���C�m��t��VQk�E�h�,������M7�G7�W%�}M�q`kk��=�UU�}�,BJ�0�*��_I	��0��'��$U�q[�oH���U�eX�c����D$�f��b������F���2�/���:�8Y(,����1�t�*|&�̳�!����ۚ�Ǎ���kmя�5�ޗ���@���,L7�����Ι��w9�����ax�G��Q����Xc�<Z���������9�+���Q	<^�>���m9^$p@WB�,��9�y�uFݪ-�����';���������&m4���:w�qs憴�\�<�>l�`��󸹁�Ԗ&�l�R45s����Ơ��%�Cɞ �%�z��_�'���=i����S����_@`~��3~0��3O���nuA9�3���V���,���巃�0\���o��@5�2�0Z�1wf#(���b�렍I;��Hߎ��av6:��s��PH5y��zHT������]����PRU�%�Ӗ�Q�>�n�NلQ�{$g��B�-�!�3DƲ�������I<yF����N�
�FDS���F�\f8k`EW]s�W��({3�3�*�L����׃!ncs�}�TAKRͥ5(lV�3-8v��Bفp���#T���
8���V��6�`C��c�l1���m�A{·?���p�7GdH8�h0�n�({V���J�	`� ���X�^�.�r�f�����c�ꎣMx��7?��E�W���?x&�+Dd�I�ݱ�f�w'���H�Γ 	8n�dZ��Q��L��j��빘*��I�t���C����G��nꕯ
���ХaH%�el"eKP+���>2����iM�zM�<�KI�Db>�1-1��}K���h�=�dn3e�e�D� ���pT��Mr�k�á��8��ңJ���@s\H�B}�5&wJ�v�Pk�Ga,��l�0(@���<�Z�]���=�%sS��y���t�#N�������v\�ẗ����y���8Kaޏ���B+0J\�f��Q�S����l��}�f�!"����K�2��=	��n��Wd]u%H�T�߉&���!�9��ZGl�7�F�$KͿ����א%2���`�1#�R�W���i^=7	K�w���b`
C�f��]+)�ʥ��-c��Q䠛��+SF��h$`{>s�&]��jj�nAY*=j:��6 L��dA�����yC[��ZF�����"W4�F�i��R簪����.[�L��8G�/D˳�po�ǫ��g[ߡlէ�#���j�'6W� W?ެk��X�3�u2�J!��҅����6ՙ��@y��)���^��r�bO=�"��b�f��ED�v���zǃi_�������֤��hl���/���<o��0 ��\�.�^�b��*Ej�_��#�oI't1�	�9Β��� EK�.�أ$1�R�j����V�oq�$P^z{�{�Qlq\i#���`��kJ ף����=�������>�De�(��ٹ���x$8��V�t+��N�A��4�&��r'�ݎ�_��|)�*"���Rk]f���'h0ؽ0參��T�ɺ�������P�G����)N�#�Z瓋F��u��t�L���FR����$����9%�Zm�ȥ��JK��D�Le�Q��!T�(�m[9K�8��O�˧xe�h���=�����"y�T�I<�Z#�$�)@lX�]��g��U��;����v�	F��"d�[��8+S��� H���BP�r��O�V�N��ͦsbp�]�r	�`,$`o�< D����t�6��M�š�fw�[�Y�aq?�F�:6�ݻ�:�v&��@�M���`#���2���&�m���e;TEP!1��m5dO&��:]�#�����>�����0�R��d��`��[L�ʮB�zz�>K���~�Y���IAF1�ʯ�T�o���ʬ� J촘6�p�y���V�a��Q���|"'t��FC�H4O�/�4���x�ѕ�#3T��s��ݷѺ�y�$-<İ�{�����16��BĚ���D�I�x��� ���Ұ
Z,_���X'qf�E��êC5u'�����L}��AX!���P��!NS��ʹ"��������@W�w�<�/�"HgA��d�LIb���r�HTRb�g��ˌdە�V#�Q���v����C��ANiDs)���Ow�h�3~�a �d������b�1���L��N޵Β�s�5lT�m�\sBik���K�0�#��.���7ZzLyV=������ϡ��b})E���`W��R���A��rO�^ߛ�/����X��[�7�q����5�|�u@ɲ���S���E�1���[���	lJG����,K8��6,��4�뀫��d7��VUM�J���w�[�3еp��l� �^�@~H,#�2!//�&e��b��1�G{j����4�������� ��oޒ�!FCS7�A�s��Py��!ń�C:���1�O�t�`��+�0�IS7Ai}�2|�6�2�6�QN���L��N��úw�,"8�u��`͏
4:")GA�ݱpE1v����"d�#��8�����k=4�̹wɝl�6 �>���]l���}/�{o鋁�a�������xR{���#I�޿��8��g�1�C��lc~כ�^K�?O���[�K�[7���]��f.��X�'��F �n�Z�o�C�T��s���R�3�lj���m�G�'��'q1���-��Z���-C�����fU�nQ��}��'��	1��Ϙ����]�Ro��#�幆�E���;bܘ��2׬�
ɯi�0-,#8'�p�~�qI��9H�2��E�N�:o(9�: 3VR�elt@Ga��U���� Tޚ�b1O�����T�(�Ƈ7�r?���;WE��7X��}�]�/�R%:UW��y�y����R�DF�M�8�+nMW��B?F!%c�����䀼x��rp3�~���j'caf(��0!� ����B$3U��e9�5_sȜ���E�f������y_�Z�bT��,K���Uv��d�t�_�`��nt
��鴆:4#P��n���|s>������
�;l*��#5*cC��i�_�����ׄr���+oy r4�Bڕ�H����Ӌ����QJ�
��0��L��鰊 ��L�##m���2�5�MR�����q��RT����4�-��γ��|şW�wʦCb�k>]-�u&����C=��-9h���Kl�<pFY#a��ڤ�/h��qD���̎����)H!_���/[=:��#�����Fy�%�8pvd�00'�<t�:�?E`�g����␲����XG����hUUL|
�k�<Ӫ�z�����0۬|"5�F�C��U����r1G�����u�u$'ߥ���qe��@���Y�mCU��(!yX/ӳ��ύ�9��!H����7����X�8�k�|������nX�� O~�pa}�K6�%
��]����S*�"���ET[(!G��1p�������i�x�͜$)��b��y�.�E jē+tN����rR*�+(��)������!h����H��}���rׁ��k��Y��Uiٱ�@�!�W�3�xE�˅���sx�	���-����A���u��x�p�����vQΎXw�oVH���o����T@�-�W�6����R���,�� �N�<��
ח�:�����˶��֎1�N�PΝ oM:��TKS�Rv�N�g�r�c�>���7��	+��.�h��Ǉ�iW��`mT5��8�-��>���v�?�λ�CY�R�����,�[��D)�����t��+���	'B�Y�5'��j������8ґX���]�d#b��g̡>zx=��p��x.�dK��Jz�E����xh�?�}e�5=�T�D&Q璓t�^�I�!n�aM�M�v�z���	IcuFb���pr�5U:�~�:��}�����*��X�9��Jh^��:�9Iz���NV�:���s�)#5,ر��/�D��W|�Ohc�����ݏ�r%�N��ʝW)�0��Jֹ��h@)�"��k(����'(h����,e�FZ�����FV-��T�u"�!U,�(fcv�e��
����{t��+��!��9}�B>�U��K���������?����JS%<V���9�:�Ȏ�-����.VP���T(�����s����F(=��+�%ܰ���!\b`r��`~ܰ�|��z�:uWvaW��Q�ü�L�,K������_^|�ꮊ�i��C1)Po��Ԫb�WzU�2˵:�A��#����?�+?�e����S�e�����if�3b+Q����>��R)��w��_�,���h[� '<�54���Aǋ��c�����
E&�@���Mf��@g��k�L]E�)�R���5#j�!��D�?:K�]��~�+�	[M�����v�� �P�9m$FR�L��'W�k���G��J`1W�+�)�y'@�ռ�m�9E���iJ��pY���>f��z�y��^<����!Lp�����4�y6�-X���h����X�BTh��� \nJ��!�����kG�vZg�)s�'c�̜�Q��گ� 3����|�=x�%&蘏�2ZX۔__.�\�6\�ޤ���L�wc@¾��G,`+��K����X�nN���5����bݳH�wU�WyU�6P������O˂�q�o��EʬVG�iA�ꤥ9rgL��U�R��{
� �.�m���g}�	я>��::�s�0�=~�B�W��	q2̧�� �&uZ�����B�W�W�ߓ�!�zwl-�\��(׬=���uF���.9l���o���U�02�g���h�O[���6���+0l.����Xd|zN��r+���y�vߪ��4o���̕:?�L+��zܭ"3҄�	8h饅�rKte�����-����Th�I�gF�
-8D����
�o��F���~c8���{s'�d�v'�l'Q�,$�ì<o�P'�pH:�g\�]�vۍ�`����̕�)v]��*8	#�Lh��=�u�8��6=�A�(�^�l#��M:�5��)�1g��+ o�� �~#�_������1H�=୘��%#`�?ۙ�FZ���ȸu�$��J�I�tr�]<8x�枠��i����G{U�K`�1>�wF�N]ߴa�g}ϻc
c�t�V|�N�I(˝T������0 �!n4��e���?�;E��,3Vw�*�ӵuS�n�/��|�`���	���Q��s�#���;�N�'�f����H�3z>#� Zp��%%^�,�$>�F�_�:���sӓ��7i�� �,�<����}=u���dك{��' ב�_�ڢ�J�v2���P�����%�D;l��݊r#�|�j�we��Q� fo��9�>�Q����-�n�Y����yN��򶟗>"�Q����F@��^T﫵�GM1z�-��Q���0�_�I�*WmH�&�N_A˄�Ŝt��G�~�c��R��`��@z>un���n�^ϗ�8x�Cn骈r�S�'�Y��X�:l`��� �3�-2�$#��E�nO)+�̐��a�Glf���Fƙ/3
+�Z!� V�YD�l{Xt���
zT��FU�Z��g䯀`��!��L�}w��	�Tv��φ���1�9LR��Cm�9x��ACE��d�y��6��P��%!�pj��*F�&!��e�<~�~�iW�t��4s]���S�����E�G��x�6��Y�#7w�*��pc���X���c�=���5�[xm�^��|�웛DQ���65Ԥ�@f��=�ot��n]���A��~̉,�o5�ue%L'F���c!�w��t��И�#S�����k�P=MO�������z)��r����������8�6J>G*8���)��ld����
Q�uM�Զ2�"�{5,���PNc�l��]�����g
M%O����1d��m��������Y-,�ߋY�	i���lFD�I Jм�c.�-����0����83AW���Y$R�=���Y�8+�+�����*�^5
F�w�t�_���Aav:['�ϥ,?� ��ķ��V
H˻T��e����Z1��U��k͆�ѥ4�</����'���DQ�а�H���˺�Ȫ�H��{�����UP��V�L$q�t����b��G�Y�r�<�9~����0PΠ*���M�	�GڗujoEB�ˡ}�b|�I���z� �39?�����`��{D��U�5�m�I��j{pjGx��R����i����*�k�ut�Rz�$-j�bT���^J��ί���j�S���;�I㴀��c��-�W=^}����_�ݒ~fm��o� i����n��Kc��������c�������)����|��U�.?���oT�%�Hm�ލ:Z�AYz9n}(�O.�i���`�jJ�˕Ç��}�5�I��n�����E$㽈���n�cO���6�V�ap��rz?�� �ɢ�vg�Lo<sy3]s�U��0�?�Y�O3���)�]^ʍbar�ʞ�I4^�[��|�?��i5E|�bΊ�^�hmX�`�s6 ���l��י�c,h�{߼�:��)��_F���Fs�!�5�L��ز�Ӣ��ӗ)�:���ǵ�J2�����m��sdT�Ё�j���)X͕k;�m__dIT�~�����L]�XTކ���y������U���%�~�s�ƪ�.��m2�Y�&���[{�����ߵ�4?V������I�qV��˨��Ç���yhK�c�S��
�G���@b�ڒ�>��w�*7�^ѣ��ӻL>ؓ���.ӱY�|�|�,b������흲U~�$�]L#\��1�����E`W�n�(_k**۔����;L-Ӏ����̚d�7�$ڜ�b�:r=��Rh�L�eD��f`Ν�#7D�$R��W���?/�/�R�;I��A�k�he+��i?�(,��WN�N���o�U��Ӌ�X5t�Vy�7p7Ԏ�TP��\�����N�q��d�("�K�߾�FE��g��$�v����*,�Fz��8� ��t��\���EM��ϩ5ˏA9WW��~�w�=�|�U	�?_�q��߽;*���#).4S��!U��4�׿�(_���ঘ?�Yq�U�D� |�C�;;U�~t�M�p7mj�!POP|[0ń����)��O �&aҀ���MZ<���r&y� 	�A��)m�L�{P����a)�ƫ��?������}�8Eډ$��#���g��%'�=pᢆ�g���2���;���Tr22�p����_�	�(R���4DL�`��SlF|�E����æ`��/#�\��gm��׹�]"^�dث9E��C�y"B�o�5z|�;h"z�������t;�?(����Ѣ�H)��7Q��y��ⵀP���L�8�5�+�HD\�5�;�u�(H-{gShs��ɰzE�B����
[�#U����yl�L*��yUE�@������UA�kw=����7h$�k�"-����й@΀��r����j��B"q�����W�@+��bՉL��LX�☳5���Yk�A*�_#������N�Z���Uta@6�������,�a�H��g��/�RH�Sa�������9\S��跑c[yyo<�|�P{�>K� ~9�� e���^����ܒ�r6]�C;���$��7͘�C�6@z�~hn\b�6��>j/vP�#�����}��w�
�a��d�2w�D h=j�+�*jZ�	v��z���6E��]%�R
�`�V��U�Z	%�������{��ц#O��a��e�>ϥ�R5� "v3t� FO�	�����t�C-M��ɗ�5xO/6|�%�M\b3� ��X/C�E�&��*t�NW��s}$X0/�LU���*�	Z��ґ�/Da��F�o
�e���&m�m���JZY
6�'��
�����/;=Bǫ��}6��[v�9%��Q䩖������?�\�cM�Kٚ_��j{1�o�l`~�R&it۳���bJ�����%C��B�u�u��3�Z�
�`�	�EsMT+c�gwY>K�!�]������h��ٱa�]\��MD�_%�ۮ&Al�I�#4�6�^s��j�R ���q[D�f]��Z~�u�*�����v-O.DL�g{ލ�tL7'�����j��[i���L�5c��q�[AG��j=�t����1��)���)h�x�B~/w��΢��ҙ'r�ןe	n�d����n�va�ag�Je��a��t�͜��D��o�!F�[Q�฽�`���@��F�Vv���.OӅיn7|�1��p�M,�N�Xr辋^Ж�MԍBS�e4�x�������#�q�P������E�^C�e�jOIϖFئ��dQT�h6&vzᜤ��q���q{�TMH��!�XE%�"2N3@��B� ����F�n��z�t"�p��"�8P¿Df�޹�h�%Ư��|�'�t�5�Kqn?�0��?'%-9��k@O~+P�t�	%�Ǆ��-�la����B�1qV�H�7wI��v�L����^��4������\^������C�ң^6�o�����Qj$����(f����}֣-�F*�V�B����<�<d��m�a���y���sR���zZ8��~K��*����Me9�:_��q�}JC
���U4:a8
�i��#�JϠ&��a#�R챃���S�0m^�J̀J��y������U�ų�5�U&�ku�s�h> W��WՆ��0�]�Qf��OQ���ɕ��iW������M�j�+��͞�X�2~��b��=�)��������[�XI�ac�R��8O�E�R��}l�,�hT���+�:D1��kC������ϻ&���:~���)�N�f�x���P�O�IŶ����;�`��~IB��������s~%�Vi��YP�gXɏ����?֙���J:690�X�ڇ�ԉ�?8/��_yO=�$�9q��U��V�`:;hB ;��m/L��
O�{-M,� *}�k�����
R�
8�G�)�|�m�܆\޺96?��Y~ M:�[ȶ,���;�7�^��`ݍ��jZ��xG�[��2-x�a>x/k���4�K̻N�VX_(��u�8b���qXC��}ހ���	K7g_p���a�ax���%cO��	�Vx��C�e��f	b U=Ib6��ON�W*��Ro���7az��O/@M?�>�`D�'��x��}C�n^���?�HUOK�}{�zDݲ�ݜ�Z��DiO^l>AL:;[� Vc^�K�TDl*�bpnb�����@V���;��&��I�fB�f��-���C�s�����?������~�:�S_�tM:N�4�e�� ��51He�8�6)�����a�cLSDI��W�����'��NK�T`�QC��6�#�O	����-�@ʔi����qT��c|ߵ�J:�c(��SR%��U:#	_�y R��n�\D�����%�|�%rvs�$�L<l���*Q��p�j��.�!gl�}S]#�a�q��L�n]�l�:�l��Q���.�\2Y�e�J�:0��7ql�A����X��t����JVh�w��-v���x�:�l8����q�R�oۛ�pR�h^bR����_�T��#1�Y-�E���l�b�&���Մ��^M�~�L�:�p��:<P܆1�ᩔXd�MQ{R�T-�!��f;z�(f�ߧqGЅ��ƨ�	ŵϫ��v�Y[oQ��:�Yn��;��4@Am���A�˦F4$�u>S��-����d�+�W�foC�Ȧ#��7�N>r>�	�8-��F�Y��(�k��9˅�P���������%��&���,� ����@�U41�3
��;(���4�a�������F{�̣,}��L�?;���K�K$���g�'Xg�5��L�H�3�.�I��?C�Ҹ#�p���{g!-�����o�W:#ŏnc^���,�iKE����UrFz�@l�:���)Я�s=e�Ji�:;v��)�ރ���	�#(�/kM��9m�~i�a�����!Kꭣ@�yB����XQ ��/`�o��K=������!��8���2��?��Ō�1	(��j�(2�9�`1�)S%�Penu[0s�U{ϭ�,��fw��4N ��8�4�$�pg�~QV��^����g����t��ҦuM���e���]��w��R���(%�\	X#�	�W�D��!zύ+�����ؾ��i|Hc���;&���2��U=?��e�]7p^MP�X���>�h��|���%��,��x��C\8��8�H�9'5�a4=�`yw���a�@�6卑K2����~~ U��y�[_��>\p�mw�?k�Sǃ,� '��A��PP�l�L�� �<��S��ݶ�]@���� K�Џ��kr@�L ���[b��2�yb���-��0ے�Kt�BZ0�3!&d26ު �FI�	�NYG���}{Ej6��?9�9&^���Iz�`�T��3s���fi���|�h�?D��<n��Q��1]�)���c���Uc-���̛!�L=rs�sB��L��G\�9I ��v��jR:��j��1��W�SP��l�F~��D_�v��b_�9�5L�1�nAuGt朥��rXY.����A���F�u6l���������� >K��c�&���hk~�|g[����W9_!.��ͪN�(׺)3;�"���E1�V�ҠK�,5q���x���j��©�X�^ 	�Rd�>���C9���/�0�k�����pI0��]��7ʚ欬������0f��{��_�s�f������,���V��CGyԡr
<!�K�H���-��l�)���-y��.\.|i��!���+��R��7�LP�.�S{M�
:�_B'�*)ox�t1����5��|�gѥ1����V+�W�E \������Ƭ�B�Y[_i[ �2�̸��L
l�HH9|�ݩ�P�n����x^�A���|�ז�^���_��o.�O�D��������:"�eu6�R4a2�����T�cI�0��2����H͘��l������J�[�e&t.��'�0ڤ�x$OL/4v|ph�΄�	T:�D�OL���(�o�!��RsX�Tװ2�􌐎˼����S����g��E�4��u3k��B���/�è�[[[I~(A˷�ȹ��~���@�[��Pt�A�o�R^��c��M_OՁ���x�#(�\0��p�f��.W��&e�*zj�.�	!P�"����ܞeE�n�\2��B�v�T��BL��SUsr��S�j�y����Qp_�b��2:|�!�Kct�7�(�4�;Y���2��|�d2�]4��D��`�|�FO�77�`���A���6��U8�@�3`K��#uݟ�u�����ɩ%�k�^�Cn���4҄}�,���?��T�\Z��*Q��+�i��NQ��ؓ��m�zrA5��~@7JI(���{�-���X����䨔��.���e&�6�7�Q�Ԑ2J+���u"��f}Q&���ɘD8��J[q+�b�ͩ��d�$���!ͣ�g�z���D�kW�Ĭ�R���I��P $'���k[St9�F�ғ������h�{��3�w>j9������4�>�.)t�r��Ivڋ�#6�Y;����2�g5�����R�:L��v�]�}Mj@V'�}���{�J I�ȤP��Ѳ�*�!*�+���+/��Z��z#�㫶5��D#���ծx[��n�_���5H�L�{���3[(4��]��x��zՓ�,Aui`���.8Qgj�M���Uz�M��ì��t�`<�\	嘺Q0���0�A��g���́_P�^�y�  ��4�n�|���n�p+�M2�V��<o��c� RU�=���-N�Ax���/Ms��`'����w�������w�G6�f����c+�AmD���%
��b�N�ߧ#���q�ʥ5�^B�$Y&�p�G5ɾ4��L^�����e1����gNG�N_�f�X� I�%�L�8��8����4*	]_����n�����9�c0�7�t�g��!/\D 4�s~M��� p�1^���!!bE0�o��I��Ǟ& �n�ņ��V���-!�:mj�uv
�Vi|�>2-���[?�i��1p.�z?Ez2�_W�d��K�Cd[,`o�ꬋ�a���.ܣѵt�a]�2�Dc~CÞ�1�M>@��Td�It� �-V��W��ޱ[��Ha���Aq6m�7T6Z�p��s��N>�,��[���X�H7�����X�V�ޱ{�;�4ߍ�i����}/s���ߡa�^��V�����q�5��U߮{����y��/�d�~&m�few�3.2 ��]�E�j�$L��\W��M���G���v	�>���J��%K�|�W���"���9�c��]|� <�Ε�>g����yj��(�6H�z�a�O����@k3V�uV ����<9TQBqf���ˉ<�u{��qũ�U
v�L3�>�gk�a]�"D��B
�H�-x��c�`���w��
[1Z[�dx�J_x��\�N.��h���+�6Tf.h���n�&V�߁(��h�/<�C}(�(��Wy���#a���	ɸ7D�2�M�=�~p9u��>R
��"�7��Z۲�W���;&�)(x�%���V��B�1S<ָ���U�T_���v_"��83�x���H���IS?�d�#w1�"Q����a�����|yY��O8�62SS厧ܗ��T�Oy|��H����L����]��#��%�*� ho�Q"M�V%z��ۈ��f,s�/����9W�.2?��qQ��;������Jt�t��gV�0���a>���nQ��R"4Y������-��ب5�A�3N,UO��ܖ�~H��i]�+q�*Iӣ�&EF�Q��P�� �®H@�s�MX��H�׍�a�}�����D�_6�]پ\�" |������8J���g���=�~=�e-��p|�Cx*>8�<xRQe&]�'t����'�t�&ƭ��w�v�����>o{�h� Rl�ī$��r@�VߔǇ9@Ԡ��.;�v�mi)M?��/0��r��Ζ��GpI:��DI؃ :}�j��:{C���S
r�''퍙i��J��A8��!�{gh|z�e�b�!
?�����v,����	����Uh���� �C2�m/?��h�GPd1g�9kt�')1 G�Q;�h�'���Ӄ��
X#=����v�r�0�����0�l�F+���qN��l^��?32�f ކ�%��Qn5��TWM����ҭ��/ʌ[�v����|��h}`?�7Ȁc:u7d�S]�/`�Xq���+��\���'XB���hl��M�����밮sh�F�U	�R�@L��)S6�w�܏%�a(���D���g �����L���k��1g����;����cj��ӂGd�0��;TVa��u�Q��5�R)�|ن���aۼ�wuC�?��)K�Q#���-��։OS�RO��\⻔;��I�ي���P���7�Lk�s�d��2��H>�{˿֙��`��-O�l�BQkQ��j�fV���2��h=�-["�ϕ��7F��)�r�k�1��r_�U��f���^q.��}���S�T�b�h�N���E���q	�YA=���$,\��j�>�c��-���e���!T1>Ψ�Hɕ�=m�%�����zi.�3�m ��|�eW�obw'��owlc�ٴRf×��i�#1�ڷ@]�Y߲[L+�]�K�����)�аR辍Ҏ �n�$D���Qw��|1=�A����Z[�{Z��Ȃ�Y��r�`Yv,�71o:�鑎�<\������*�ϣ{�r��u~���9�2���0-��X�����h��#f�:n/����T�6�+�FW����}�ݾET��U��)U9F�D��O
s�K��/�H%W&�C�0E�"���l4�gl����_@�)��hH@��3�6EG}�$�Q���<K�6�y��=�=�])~����M7��
���tmb�H�ES�JaJIH���dH�7Hq�NY��o��O�)d��]5��.�����N_:y��j���`��s�����-�ӫs���ڷx����V9r�G`��J /�6/�ϣ�gq������Q�K�����n�����e��)�eCɰ;��z ��~潉FYR�E����z(�M� �X��[D�<�=�lś&��9Dl,k0f:��dA����D��U�)m�ٽd�9~���������ŔP~#���ӊ��d�f��`�֎,V ˆm2Q�)� �A�q{W���5����b;P�^�*iJ"T��h����f�rYu�pW�g
L���] �0��i������z�B�0�.�����̑_�&c���`l��Mֳ)휗�n_ۺ�V-��9����=�f�x6e!/��&���k"!$)�V`*�=R�O�5�Œ�C�to�B�J���Uƨ�eb���������G�����~@H��U��UuB���C�;�Dc'��}��BQ�U�c�t�%�R�;B�F���"�1"����0`Ž�7��0ĭ����j<*�<�kH��i�Ei����(�QT<�W'%|sck���*�P[L®��T��1ζ��f�)��|�-8k�$���L�ε����Q��4��]4e7�y�%���@�ĴPz�W]iʝ=b�"�hHr�>�h��{o��k^�B�=(h�E)�fɸ��\.��_x��I`�����
[��b�%`�J@߳�������89���>�â�h�b��մ�#�Z&а-:v�"�'�9�Fl�������.�N��G�������`�
[��`4h]/[���j�\�w܀���-�10�'�
�\2�p�HrEW�ND��� ��m�컱!�шa�:31�]���u�4�����!-�D�@�����mp1��)��g�D�E���3�i�����3�3�nSex�خ�^n�8 �i�����=�q��(Nq%,�����9���9=�F��M�#/l�C_��zw�����=�Z�^YZ�[�vsjf-ɀ��b��f���zmY{uY���	��(��!�K���Q�#tȵ�g=�)O*���lw`:D+(��ɟ�';�8DJ�f�PkJ��O��o�7o+S��8��B�ӛV���Pi�����q���[b��|<�bj�q�Ɂ�~$��c��֥ui�i��KEC�$�qu�	K�,I�Y,��J��H �uY6{�M�^�<���km*ʶA!�'���NZ�0C,.�l��6�������������S���p�O�0������B�ŕ�Fd,t$�M�dҀ̝�	�c��v{�S�Wg]��0�����:��tx
����;3!�yl\iRg��,���aS��U�ν5���t�Bs����_;8H3�{2�Ʈ�r6��`4zWF��Gh�˚�(�sL���GC3����-���Wï�	+�cw�:'~Ad�Ywnޗz�����t��3[8c+S/�)ERg���^6>i�Q��t=3܄iV�\��kE���J,kw��M9M�Ȃ�ѵ�A�._c0$C�)�g���VvÓ�8g�f[�KV�֖���h�I��(����>_��w���+�^M�s	�W��;�G������W/.�!��""/u�.1�v�+���E���
trK Hvf��%���h|�W�nqk��L��-�yie�p�7�}�Z������K?�o��8y�[;Gu��?���������M�/���g�-�,E�5�1ؒi�p@^?��ud,�jN�`\�r\�Ya��1���AI��A�,Z=5\�Xq[�nԾ+��V2S)��LĴ�Mw�k�R�c�i�@mN�R_!�I�i�\��I����5��I����\{F��	`"w�  �O�8Y7������MP�C�L����={���J��ց��T���ֈ�O����;�����Ag�b��y���{MOц�^p+O�ʵ�����"x-T2�|�Ț��1��Z'\�t���x%V����S�	�%���`�tj- �@~H;�ԣ��Ъ��y����k.�I��L�~aˮ��x/V@%Sg�>�aǔl��oXؒ�Wk������7�o-�P<�`|�4y�T�^�r~��ś�i9Kr����<�"m���P�8�ge�a��r�^ߩ	Z�W� ���F �1fr�Lw�rkN�H�V�
�����[9��V����$�^�6]����=&�O�Q��^��3�x�)���N~�N���MW�ӽ��p���2����z�����S�8�nc���-}N/��넡������3�6t�F"U�����ѻ>RۋQ�ڝ款eG(D�U���~�8s_���̣�P��ݙ"�c��	Кfa��3�@;�rx��D�t�16�!�@�&��T�1�	g��5��M�ha�O{�2T���]o��j���9�>�})q��6�(��������6y�e)ܧ��+��o��ɒZf������� ��x���ܯr���A�����ڦ�)D�ԝb�>S�Gz*0�����r'G��q1KV�G"6��@;�l.���(��Q�,!�`u�eU�d6��������r��6:S�]�g�G�#�hv����$\QM�<d`h
��\�[��P�Y����iS4Tc�7>鄜���v�1��<�v��K��^8�Ŏ:���p�l=]�*������Ѱ�"S�KH)P��T��V(`ڋ�����$YPߞ��(ѭ�M�d��$Lq�e�����s�{�������vc��Զ/:�f� �,[�qg��^��_@��C�*|���E�$*ݓ��j(�\��� ���9��-����[L�޻��+9��/��G�^�J���0]}_]Q4f<*�b�؁"&Pv(ӱ_��\�vn�^9�����'�TQ��2�_�X���i��������U;�>Y����M]�_�4�ִ�ð�3�;L���$uh��e��l:���KV�,�Ƈ���A�5�J7[' 8_�JP���$�4�ʐ���#'�D#(�U�P�[B+�#�);H�C�ld�Ę`P�G07�W!|e'(��{��@i���}Ƒ@�5�Ei[����TI.Ɨwi>m��~s�/���*RWŲr1�f�=m�Ɓ�6B���W�`dB�.p\)h�
�oY7��O��2�x�9���x"-Q�*N��!&�^*�ͳ�FWx0@��빭=�
��:>�U�ȴ4�4�����p�DBA�8N�-F`����0����ڨ�ՍW��i�y�1�sR��ik6��D:����T�p�6OmL���x�څ�<�Έ� �]:Kr�,�f<i�]:��e�[j�c�n9<�RV�<h��4�"-�d���%�-��a��vM�}�b����$p9�W�Z�5�z�<�@xI�^|#d�Cӈ�d_�KX�ɈdW�~lY_J��x�;���|%��IJ �-���Be����|�@TERT���@�h�s�7�x=��}�h�G�b���ہ�o��:�I�J�.!?�v�����k܄�wNל����+�-����,,Q�h�J���{�3os���,2t�L~Y�r��aD�8���CC��MWi y�Bֽ���➻m���Ap��&�&A�M����ׇA���x$��G�v:
Z~�s�^U�H�m�vV�9|�� s^�����"j�f�LVM��oV���K-ነ)_���>����'�{����������'�8~ļ�D~/��.��k��:����.y��o(�#z��xV��z�m�\/��0L%��:lW���^|���)���K��ͬ��̔��Q$�0���.�&���<�F�<%�6�ß2�u��2�����p��0��1��|�ɶ\>7���I��~A�������k�=�[b��u�;�\��
iߠ�3/v�,۽��4� 1�'��e��1ѵ�:%�%>i �<4���(���+��m��kGq����_9�V7�p�hȠ��ki��}�����M �L}��ͻ�҆��276P�"�G^g��H��4���w��t��,-��X����H����2��~�}#�w�&i�
�s:*�T��D[�O�]
�����*��Q���R]ן�m`�[���]�p���-xl��\5u��U1���ǣpiN#�TR�Qa���F����z;��(>!�f�&�	J��+��V�
s�@�3��0�sb\+���k�ž����Y�G���Q�v�/��ݒ�P1�ӀI�� �ԗ�?�#�;)�xɍC�x�*_�X�J�����;��N6L�z�hi���=	�X�#���Os�k�n30^�����;w��RU�^�N2��(������F���TT�a!�jfF���>��9W[Up��1��Q^��kRF�]�[��?�c�e8t��1�!\;�����}��'�o�َ�U���o6��ę2�����g�I�z|�%�6���1w�l���3�l�^���V��Є���x~5_��^�[�2�p�"o_�)V}�/{5���1��%�MFZ��X�*b�� �}������J,�и����`�)RN���'��IT�Z�趎l�K����8S�N�0wu�(5���4J��8�>$���;��C醧�3��Ra�� ��m�\A�L�|��0���f�G��leJ�v���xk��������j��CT�}��5�����o��	�\4V��s��N�Y���������]�"3� �3���ҳ����*5U{꒲C�Z)Z0�F����Tǹ4�rgp��(!��Asښ�^?��Bd��R�-KS!����^�݊�7Ɍ� �c�n�e����4t�P�ԼW����\͑~��.�8A���/��Df��%��Bh}� �x� �|+�t�[:˴���@����y3��C 3Ox��<�:<S�m�����\Brk1T���N �~�Z�[)G8����O��v@�b/�W��I2%��� �j�*�&{�M,�8B�ۮ�
��v\��Dw�r�
[x���pe:. �e�n0��)/`��]���qmR�T^V
���d�Zh(v��	������r�ŗ��v��\��+��x������Չ�0	��3td�R�%�Jo�k5+��PzR� �Ŏ����n�;�#��2q|TF��&cܗ<��Y���
���2�ޢ՗��d0Sv]���:8�7JҚ+l�R�kDn�kV�TK������@h
��zb��9\�R ^b�����ޘ3�sM�+��h� �ƫ�h��R�S����#@e�+3_���6�>��Tz�8<����$�aQ)@����$�LΎ;&�>u|1m�iеo}YV)X;&�%S�K���ג}��(O �Mo0d)w�Jd_H>g<�9f)?_�BBM��R��!}md��[��y7�5�A0�Lӑ��U��Ϊk�0W�n���#�p��MS�=a?a�U����`�*�H�z(a���8�>�6��Q�q�m��3(ZK���ֳ]���pmiۑ�e�@Qe�����`5nў3Ǹ��Ś�����vs��� ���,q�����kN)�P.���D�r}'Ex�� a}�J�%C
d6��C��*���f��٭a�1=3Dl�ɥ���8#NG7�!J��azʑy�����~����ɧU�T=r1�ʟt��-u����C����������C�]󼵟�QW�\��0�q� ���ڋ|E�O���#�r}�?��t� A���x���θ_������3gNIlƃ�Ӌ��n�� �!�\`V����a4�8-?_:<DT��1�W6�(1I<?�U�~D�g��ٴW����4Hz�b�/.f�_�t�β�?c�Kk횎<z[���Pz��k]���L��2��hyl��&5��
�"�8	��a�o���à>+������ao"��x�"ۀ&V�6I� �oML��̬ITλ��C�g�S��b -��4iWwYS}�% ��i��^ �z���qĕIfO#0�`;?��lX"��9�DQ�����[Rs���c���SF½5ɁJˌ#Gt����^��U��[��Yt��g��Կby�)?�5��tf�޿� ����ڏ�)�YIZ��P�\֗��-y��Mtx��M�q���zx8�Z�M ȴ��Z�!�����$�GKl���������?ڴ��u�@u�[�hzg~���/MJ���E�N#�B`�ZNm����vc/�:Ē��k\���'�bqƦܜ�z%B����'��WeN�y�@�a8��.T�@|D������8d#��z؟����+[0D�Ul����\�?/j��@��Io|�h�{�����?��3��*7^~���ݓ }�e��њ�
#�(�S�0�Lb=*?���p���8k6b�*�
d��N�q�G!���4�T�����.%&���y�q֞�S�+D�edE�u����sA�3�	u��և���B����!0�sL�[������Z=�c�ˉ]PQ��{Y��Y2��\<�S8ON�(�[MO=XE� ��)[��v�|�0��>�PIfy
"��\�CQpØߛL��J�ޤ}�M�G���9&��*��t~���6�2�ʻ׻
�c�8�.�myUr�By�ft\�Hc�
�ϱ�uSM�����w�#y���IȪ���d-�=RI���&=W��D�ˍ�`x
C��J�6����m�����@x�(��h��y���tH2��Ì6����q�rD׍z���<�WML*1C�IX��({G� K�u(>�V��d2/�·��cUu�y-�:��I�Su���,Vt^a � �1�j�����+pcN>>�C7���1WD�1+�N�ϧZvrR-���L&u^�ݻ�A��&wO��+H+)%rI0d(nGIQO�?���,X3Dp���&�1�e�N1�C��oAQ���oh���$�9���� G�n`�O� �wS�e�c����~xAHy����(�{��1����n�(�hh�V�F��L��񗉣���1I����G1��b=H�5���X�j<�w�:b�<$2<��K��L��_C�D��(�9�C��>��H��#�YB�8�tّ,r~s��U�S^#ß�-�\�=9����઀��֌Y;��#��*R��ָE�p/�H��>�
T�4��`�34��?�D�zؤ;�n������Q{(���	�𦤲��X�.��6��8g� F�����(��L��1����qqth�Q1\�\�`�d��^JR��u��m��� ��[����^�l�}�u��!������ʩQ�c1@c��P��Ĥ�4��������όqrVt��^v}B�9W\��.ky�lS)��!�b:�qG�@�b�U[
�Ł&a�ɮsq>q)o���4�����G ݩa�lZ6���l��9��WS����l�k����S�{�+$�JC�k�*9G�5j�J�eԬm� E��}>e%�#��]�о�wNmŰ��x��//��3_-��L;]gS^��^�p�L��L!�OWn��x���7��8���K��@T��U�5.O��$f�4�T�A�!�h5���i &�jI��bpQ,��TR1I�M,_�����t�&-(�45&a�zs�/���Q�wA�/l��A���`�;Q�C�D��
��;�^O�X��-�m�z��4�׶�,�|i�X7���*~")��`!q��Q/eך�D>£�K��˽�a�%q�k��v��F.C{��Sٕ#�u��ϥ۱z�T8O�؋�FJ��E贰궇	�d�=�w-���i3�0?�2u�o�϶���X����K���U#p��M�rL� �&!��Yc
��Ѿ)�ڒm�M2�r�p?�l�"#y��]�g��*�%H�G��^l�;��u��I^�U������Q���Gk��b�N(J[;�q��7��}�@WQ�e��L�z���݋=�x8�� �N���,,-�����	a	=�K���4 ÑaFbmJ�Čh $�g
��W��)]�R��~b���w)ñ<`#���MLj��5N7�F~o�}��BQ����)Rb���>����4S�*9dΥ�h�F�j*�:qI�.Q[Mο6�oߥߙ��æ��f>\���s�&>�)�
N�9���m��؆OF >V��!��(��d(����d��i�m��;�BKf���!Ń����9qĞ�V��e`��d�wx�Z����[��{��@����j�
�N����T&5)Ǉ��V|K�o�������~�K��5Uɛ��u]Oew6�J��Пc %Bd����#����a���(nJ��;#�.����3��푞�r}���r��=��Au��Rmc��d�eU��� �Q�{�Z$.���y���l��4^˝I�E�?��	 ������4���<�z�p�t��w���)��b��������1P`��$�ҚOe��dzEI�\j�'��܎�.�Q����ŷ m��r���=R���v���~r�������� QATJ$q,_���t�K�r�'��C�`����Ջ�����p�z�	�rA����o��|(�F=�	��B�2Q�-R��P��d�vv]��c���ciI� ��O���	���3�69��%VO%�:�j���æ:���3$^L��-d��.����Sbc�@f)��j���|lB�)>r8���>�	��4��;���wf�U��*��\xϮ�Y�Ь�����"R{����Qw��9M��Xó��ěb2F�^�r���h�T��*��ٌ�#SP��������E������2S0yWsv]�RGt_@�@&�;�$��e�A���M�QC��#�]��u���A��ߝ�I������8=^��� @ֈ�A���3DS`�ǡ�i�_L:U�w���vS��1\̌]�!���f��D�h��̔��C�=�JRR�Ҿ����}~�,%2Y��=܁k�R3�g�[@�Dގ�K���mdj�%IU�Ѳ�r�8]q���yxCpgy��a�C��!j��)�@���F��U���L%�W��se�i�l0ȕ���2���ƽ�qZ�n2[����T�E1+M�V.:���U}�	pY=�F*���5fj3n�@�l�{�����`�8ÚWQ��T����ʞ_���)���E����xHHz��.=��Qt��b>'pȰ|��9���ч=s�;<Ι@	pk��������ӥ��7$�,`�8&'#�v6#X�4Y��bڬ�����N#�̽��$y*lj����H=�(�6$�Ɗ�x�$*�}�����1��g���p�uj�r���'�>{k=��4��G�xҒy����w��c��-�n��p���Dh�	,-!1��>�k)8Į�����zO�c[ep�fK����0l˘!��C�c��ۈ��c����P�o+�;Ǫr댼6&�����b�C/�GBP��*X�iF�.	����?8��M| ͐4w����<�(Ğ(�!��u�5���i�[Tpj�J���l}�.��
-j����>�L��rX��O� W�.�T��Gͥ%Y��k\)'Y�S�OO�;���'�s<)�q*_Ք����%n6�b���Sf�2�"âF���� ,��
:]�'�MŽ�\�����s����`�L��M�H�xm�Z,C(��eر�ٜY��.����H��5�7,��a`B�~�=��3���پé���1��2����(�^�xV7������:�1C������X!s� ���y��՝ y���^����SQBSH㡤iA�kU8J����/\�x�Q������HA�|����,�s+��Ksz��	09�.���s��
��[���ڔ�B�'�u �1`����R�!kN����ep��`��(]]�}$E��q�Z���;�V@��^��#��H�A0�N��7e�H
�@;J� 9���9Q�7�9��߽�����|C2$4��u�큃�����@�;^$N���c�<=e�m4��ƊX-�s*=Vҳ�?Qb�Z$�����Rt���Ib�;-m����[D�X�r��F��c��d�ᰏ!�����h��n�5ox�R-<���, ��Ku�}�B�ID"�H��� M����G��Ğ��hJ��YG�b:}Å+�t$�����WG&������8�Oh�B���,�TZȨ۰��&�AG��g��=yƳrg�l�2�`~�%L�������Lџ!�'(�N0[������ ��3=����<��~?h!d#Q���,���Vr��T�a�h!|���)�y`(�̥�g��ҡ����<ֶ	��3�Ђ�D�c���
�a0��q�H(M}
��#L�����ư�ۉ4�MC�h6x)OWd���.k���L��zMa6�>�Q|��j��P��Y|�@W�>eU����u�����;w�ܚ�}I�nl�`�:�&B��Zg&m��E�g'$�UH���d;�c��+|@ Һy�oTgJo�6���T-2�q�(5�Ad���\`�
��g-�AMߔY��b����a3,Y6} + -�CM����%�[���[�x�-��4�1�U�,!�R�su�e'�cw8q�qή1{�,��	摐!n���<5�S�Z�+�\�����s@���C4��)?��vd�U�x����E(��u_�;�Ґq�p�ױ��U�E*!�OƀbX%;�D��sGl��pN(M����5!���|-���=�4o�«e�G�N���5l �!Ck�8��� ���Q��B]Ey[��(k��\�]��%�̷b��5��f�GQ�����k��0�	���Em��W�Q�=��'u�m�#r��{�+z��IU����2�r��Ǘ1����0��t�k�M�\".p�/z��p|@[z�~B�ss
���~����tL�U}Y�U�MX�o3��Fڌ�ٵ���񹱺�� �b��OD�*��ƣ |��.���^I&\a��nǁ��Y�D�n&� �T�vZMQ(}ŚN�k���'s��p���X�&��-�	]��͇�^�Г�k���B���H����zDI�(��y�?Dv��PԌ%K0V`1c�{�B��.Ox��ؼ|t�4�R�Rrkz������uh'�Е�,E��}�~�۰eK��\r��+[$�1d}E��l��Q#��v��ϗ�ʖ�\g5TY�s�"�&���(�9��:2��2� �5F�S#k�k��u֗��0�t�%�d�(�f��/[�,���;Їe���Ht��:'����t�a��p=6��H�6�lq���}K��Ux6yt�Y"[�|Z�v].��FI���5��د�f�x'[�P,�[LB]��~�aZ���D�?�F�X$x�����U�z]����L�(B�2fw��^}�����)ʩ�sXa7����Z���R� ���5f,��q�h����%��ƕ}��Y��Y���~GL�=GJ��/��Oɗ���uò;��>D��3jNji�	�,X�ˁ�7�|��?޹T��x<_���f7gd����S_
�צ������SU��I�ܯ��i��'.��,�)��\���W7ٮ���!+i�<�`�2o��v/`�޷�h����(�X�A	ܔ�Uh\��MAu�~�K�ׁDBl,�Q��C4Zo�y���;�i8�EF&-G�*�1�k�*�+�M�2=��õ��;g��W�	=A�fA��I��2�GB�� �@��{�lq��M����	��|l�8#+�|t?2��2��)Q+=�o.����YN�ӝ�j��^l::�̒י˯JS�_Xwi*XN��ݶDO�t����	����J�ܳ�c�7����� c�N)��*(cF�8+��7���isa��5�4��� E!��冎�ʬXN���i7T0m%�r�y�#b����^����| ��-Pvk�����nÿd�ڲR��!�U���҃�	5�Bt<f�4Q�/ȟ�_�9&w�)�2�Ǩ0���
��0���Q�"޻n�#��\�7��
NR�e.�+���E�^x0�l�ى5pi=>�;dl���]&�ˊ���UE������~�=-���sjx^����& �)���I^��WXV]���Xp�K흍�5w}PX�����^�Q�KÖ�X��3]����Y#�D=���#�[yC9vw����A��a���7$1*����D�:?��< �&2rj>�$���d��PZU���:R$��d��0�m�� niuu�����}�ʉF���s�Y��_����L2�����7#Kqj%�=�G�0���-�O(��R��:�v��(|_�-Z̎���Uq�i��&cA6�٢Pŭ1X�r_[�]���ꚙ�â�����]K�������:���l%�s���N�|C�L�* �3fe�(8M��8�S��_���jH�yxV2g��0� V����/`����t%��b��v�UQ`6��U����>�z�2��Ϩ��5K6&���o���Y��~���ɰl����j��;�L��=k}�t� �C����N��� V< :�/b(y/�Q�~kfǠ��<�n�*�D��� MlV����}��ǔ��8	2�V��S��-׽>�/�Z�@�=��ľ�������k�2E���܊oU ]����"i���rEe�X��|81��������Jm]ې伆z)"��X�O���f&1�vy�j�(����c�'ړ���&�_����O��VjWӽy�id(�xx�1;��x�,;Z>"�کc��I�v��!��a�KK�L9>����&���[\�Qx���ڢV�c5�HrBaF����d=�8�,�6e\���s-������~gž�H�Q����nt�o �8�������W�x��z��ѯ�ڋ�|S�)RV��wO�ެ�_�xt*�A�N� g�1*���nQB\�d9�Ӽ'�,��
���@�Z�i*��u�% �!��t�\�{^�U�'�������4��U�6�Sx�5���C�����;g׃�,��$��S�9��H�+�\rx����^��k����S��@�m��Q���{`Q�pҵ]p�6N���4[��{���`���82t�e-����[8���w��@�<��hV����Z��G�B���l�����C^2F�-�S��}v���u�?7���>^v��ca-�7򺌕�hm1�)����h�����9U�:����>���.wP���}�q4~r���(�!8���%�?2�H��� ���Z�2&�g{HE�?q�J0=��u�/_*�;����%��_��'���.4a �}�&��X ��Bi����/��y��by��	�(V���@Z*�H�(�z"�2��( CHR9)Z�_h	�ʡ\)�F�o[�~�B3[H��U�5��`+E�>�b�p0��.?F�!*����HT�[�è���|���Yu.�;'��f�*NV5g2��ٻ����˽{����	I'��i��iA3l��0�;(��M��b�z�������0v�t�ݩ�!�i~��Ѩ	�NJXf9 ���fl��j7���+Ix�!�^1Y}ޣ�`�i������Ed{Y�q���'UW�z�CuI��>o)n+�nYo��#��أV�����U��a��I�$�fc���:Y�mT�}��l��l��v��%�q���=���A�G,���
 OJg��y<oU���QtL�4���C�]I�'��1U	N�$7v��Kߤ$hS�9�AM��fa�a��o�r������;�������@�Y�r|u�ߎ=��N�=Y��{����wӲ��g�34�
|�s�#�6M����^�͗^�U�쬛��P��8F?)+6!�9іF7=[lFp�B�:�45��k,,���ƾ+%s?�b�jr4#��\�5��z�-Z{dE$��iR'��&n1;'	�� ���9��\�)6��a⠁��QN1���֡��y���@KݍB���Ƈ��V��N���>��?6�s�L�=��1���������F�Q(�s F��d�<3��}9�*SAZpo^a�9��l?*�U�E�0>q5K�|(�Jgr$�-$RCN5����9���@�ֲ�%��9���|@��Y[������M�M�[v۾M�/1�?���x��B���'S��;x̀�����d���}IT��G&�Tfި�b��M�3×��0SժThw�������*��3v�m��]�F� ���5�R�!ﻇ�s�Ԯ`�~����ÈN|���_I��˅MQ\���)4�$�� �V�(x�ɘAd��Ta�V��	X�מ��0'��,vM�9�L�7$)oU�I������
S�w��YCƑ����d^%����i<�#�I�.�k�5S`��z����Y�y�����#��0����]�r�pP
��R�F%�wI�B%�!H�\��cN�=�J�ĥ��)��q��g�`����N�#���;�sY����24����ݻ�߄�%0HN8�z~�@�Sv��fr.g��9�Al6	>�E��s`r�}����6��Q3���w٫X�$�7g3�Gק�j�ՙ�M��K:��A�$H �'X�\�zi�8��w���9e��W��!=����Fca���΋�.�׽�Vh����XP,ϵ"�o�fG��77����	ؿ���	�Y�͹/J�MA�d��l�ׅ�	�����HZc�NV�>y.��<���:>|�kx���Gn�^������� ������ n�y���̋l�r�ء��}@��Zi��)��X`.���_c" ~��Vew�@��'/J�2��<ǉ,TO/ڤ%�(;�=�llxZ�3@��]���#{����笠�Iz�
y[F��;x��E=ʩ�Z�l��A�wbe\T�+S����;{�X]/I����T�O��u�v�0������aL���@��S/!�`����Y	�w��A�ӊ�� =����Ĳ!�V+�[�O����������HR��P8V���.�"^M8��g����&z'9�"�hl��:Bs�v��
,��;a��YV����*����Cx+gT��m����"߷���8+��b�uMߖ��u�0����:����ًY�\IN��|8�=��V�.�kԊ�t9rw���(��h2ǳ��vK�h�z�<�Τ���6@,�7Ї�z���~ìkF&a��kJ�+	�o�\*
��^��l�B&���M0�W��jMR�B����]I���+�#���!�t�a7�hZ�P�9"��ό�OufH�D�x�,�����Z�]��-�����տ]Cb-%8 �Q/��i�z�rJH2�M��Mww]V�r(�A���+�/@�GEE�G��9UɄ/��NK��vrX̻1�����vx}� �e��<���"3K��.�]/uЂ^����^�TJ���e[��ζ���BP�83����̺��%X�+U)c�7Oz� �f؎�t�P���Ɓ�U\ep�/c������g4�ݟ��тJ0�D���Bt����{�jn���W�	\�ذ*����P
��&����K���w��{С�L>�<[Z�;|�$��2t�3�oO��D����o��뭗ߠB��*/�0W�Ț�	�J�6Bؚ��޳�9O�)��F�'��#���v����x)���t��f�SL�L ���R��;N��c�|C���h��|��z� w�H�[�;���r���᠞g9�_�}p[�h��K����o�io�֍>7��@���H��Z�ư ����COvj5/�O����A��`���1��4ZYU�q6�E���cȋB{}��Eyy���|��̌����"���|*��fd�D�3)�*��D�{m�]g�$����0�3��E�����9/��|��V^�_�}!Q�d��5���yt��K�	�9/>D���˪�i�b==��z<-%Lެ��� ��$��f��w �$f�HrX��|��>��E'�N��:J��å��R��m`^����Ba����҆�����b�����`��~�"Q�T���Ni���h`��D��g��N�!�a���F'V{1�����m�_g�aK����5������K�jٔ��AL�`M8/A-5��'����Z���$8��_n[�5��hĢ`�g{�N�!L�콐�,l�o7��}~����Lv4�`m}C��t�w�vJ�[�E���(�@��UIkR�����gO�7٦@$���yЧ���´-�F+cܡ��m�YC89���#!�Q` �(2�[���"�|�� �5�@��ýA�����n�V�����t�+�=�xo�V����v��/}��gE���G�ԫ�����]�pfV��"i�nV����*v���g�b\���VQ)����S�G���D1�HI�Q�����mO����:�qb�,';y�@�Ojktr�R�e��0Z�(��]>b���[����$�	�����b�h��o�B7��g��ד,���d����&dR�|����>n6lA���ѧ� �i�>U�,���E�gw�%�E
�h7ƨQ�N4-==�<腳�~5p��$�b��Q�G߱_x^>9�(O<ه���xS���G����;��O��M�@}�dӹ�87J[��%b�{w��JRح��`��[��H�E�b�m�(p�R���,��+ěp6�׏An6p����Ӝ4�Ӱ(l��m�!Y�'�b�z�����Y�\�$
ush~q�cA��ͅy��\R�����`>�F����J8ÚN�e˺�Do�	˝w�ʑW�*�1�\����Ѡz~�:~ �h�ßu*zM�M0�ʟF3&���{@f�J�e���3w��,�W��+��$���N��X[�PqwNn�J�E����)������5�::n��c�wT}��u�y�t��
]3=u!Eѡ:L	톽D��v�v���ۮ�ï��C=\lk���y�B��� d|^}rMM�x��ۤ�%���٭��E�)��< {o�Rw���SE�i���]P�B5�Zl���ܩ�ْV�0���Q�F�]z��~v����S�Uv	:ʸ��02�������Sky���.��d�䕽���E�C/`(��>����r��1��t���K��?=V�6a���yh �ڵ��FdLm>J���+���40�T@�/<E+u��¿�=��+�`!,Zyk���>E�aeD1�LϨc�-B�i��秄ό�D�e���B�]Z�X����C�w�J�/���i�	�k!5��-����!��Au�=!q*�֜yA��,h�i�	t����Ӭ���^"���='�Kr�P�G+�� R��B�v���HD�)�siģt>!��Km�U7�Iկ��M�P��̊o9�p��{XBѡ�����?����w1�*L�~��Xl��H�ñ�L"���>eP���b'ڢ碪�0ǔzO��{~���ñ3&Ж�)K�{�G�эeϖ�(��jO��}�aO$�v���@���K�\X0Ӌ�fiK�M��I��G*v�
'�1����
7��bmh�CYW��ɣ�ϱ��^�ЪL:Y��:D�v�Z�\_̚f:� iL�AƟ�@�����R�B����(U֬/y���/��J��M#d���-V�x�XC[���
b�Pf�я]�Q$��,Di#܍,�O�B�T�%Ky�sX���x����Ƃ奌x���0
��8^�E:�ʅ��R7�
I��F	k���b���|~�%1�1nea
L��������yZ�f�q��rh���E;}Np������	���9o��!/r$+)х}Z|��c��ABEep��v�}�o�����}	GeE#*��E�i�0]��n�{w�-l���W�C�oQK�x�ɰtI������G_D�iꐯ9R�Obc33l�}�{��yP'��<� ��{=�i�0�z����BѼ�3VG�0��
X�b����9"�]�����z���Z<�ͨ�Y���$$/�6g�jDP>W��+@BR��%�4y�2��|�dpw����Q�M�h��9Ñ����b���G.��h�<���@�̹�OdlZ�"�v.��jv�*�v�U�b��A����t�_������IW���.�[:;����_3��8z�-ڷPT�1������0x�)׹Qm>�i�*�]�5��4���M#ڷ��q����^��!�^����_�M�V�� J�:�|����xEY��5^��IV�(��T����#��?���w"7$b�"� ��E�a��ީC'��B��R?�I�A��q)�Fb7�Zl�����՛��NR9������{�����>u�B��H�;*��D�b�r8�t���qv��|׷x�;�v?�6����x���eP�X")87����޴�[R3ٲ0����2�� l�
�E�ZK
�`�۾�*���ja~jǭD�=Z~aq��M��-x��,f�p&h[k���0�5uAٲǰ�>;�4{~s��n�el
�ԆU��(j1��*,���x���2�XO���8�c'�T��_������+��)6�ڃ�s}u���vVg�qp�&'��b��o�G�J�[]8>-�/2L_,{�6 W�ث� ��,����;����y�cS�}j�=֬4�N����IlƻN(6UB[��me����'��:X�ړ4��U�T�x�Q���{�j�+Cy4<>��p~\H��[B�9i�4��z'�YW�n��0.�,S�0&w��?m��BwՃ��e��.��C��8�=�hp��$�+��$`������Uqp�k��2������0Bi����~K�{"�=z4��&^����X�eUh���Ti�Zx�MQ���Y	u�6�6�ʵ*`�,�Qs=_�����r}�Fػ��X�޻Z�g:l��Ծ=g[�T�1�)Ċ2�����{�SK'M�a�a�V�ހ&�d�kB^ ��Zb{Eɼ�U�Q@��O�����[r��!���[?�N����d�@��{^6�<�|�1��{}}����W_Ory ������t���Z�c^B���Ϭ{���\nx�JԨ"2���9_�G�&E�~0Is/AI��M��g��*I�Z�(���6&X@wy�3vf _.yX�Xѵ� ���b#�u�|F���zs�
X/��L���7ein�J'pZޛ������� �N3��{:X���IF��V+|�a��2��ѫs�%����^x 
�������	JE���g�D���]�L@�8��	YI�T�m �$�d�Wk�:)<� _�:��Ĭ�'����{Z^No'r�J������h�.�b�d���e�i
+t��`E*.�iV�ܥ��%�<��/��qA/�HR���g�k�Q �$�_ ]��(g���0�'�Z�
��b�w ����F���K�>�WH!����dD�g�bw��hm���\~?��;�3/��3�\#��!�x�s�/.�
��J=`͂���-j���>�����u�<�geW'4�s�2a Ų��vQ�r�i�t�V�A� �@��>�w��@&@�zX�
}�]�t� u����)�L�i(�	>�)U�I��1&
Q�T��(�����޳�����l'ޮM��9��5�՟=��V���:�H-WZÃ����/���q��姪X�^��a6ᅜI����h��?����>K=#d�ųm�?*��F&�B&ˢ�-b�I#�k`;���?	F֣p�Ǜ0��� p\\v�7<�UO����O+�Y�zY�0���-�-���l�M#||�2>�����+1�8��D��ɫ+0�����/g��oV!��D�F�����!׸� ���F�g�y��>���u���9����H����"��⮻��Af<�'w�i�T���5��!Q���XY���6�J0]@}��ٹbu߯�k>B�nr�B8_]�,;5Ei]�6(|ROz��(�6V9����,C~y�����%^��3c:�V��&�@ ��A�
>u��'��T���vxdJQ^m��(c���w�s����O�Z����/�,��gм�G���{庮*s�!�<�l�"TP�����M"�d_�K�\�a���U!�d��T�9�t��Q��Z��eEEJ�%��"sB;}�����S�)�#n�_��V��Z�l�YP���-(��L�-�|�"I���|�8)�v����u��|\�#*|�(`w6T9r]�Ukl�+C~�+�R�x�j�����-�I++N>y�0b�	[)&�aԂ:L�ԡq��{B�Q����)y���t�lb���y���~	K�l��"�l�s
Ƀ��V�/��&ܸ ���؇Ѯ�ԫ�;����R�ʙZk
��.ȼ�����UKۆ��Uu�f�k�r�'�x�t=PFɟx@��^�bC�/Y�ķ�G�B�. �9iyY����1�a�*��j�7ϔ�-L@�\�l�'�	��@Wi^�bFw��|��$V�*��J_ݜI�$�݇����������m�j�F4�/�4vk�~e�=�qn��D��젷E���%+l�p"����7���%���Һ�C'D.i�ǒnD\' ڣ���|\HI�m����%g5��sP��A-��L���m�]9W��퇽����@������ϖ{+��<���Zx��ʩT	� �'��P�<�`���O=��҃�ʳ���Nkk2����0�B����
>��G^%٠M6 �80`x�V�����O��Ia�޲n�sF��qB�V���]N�=�5�C����k7�	lk�3�ׅ�Ҍr4N�r�v]�H!������vZ����E��u3�X�u��%e/<9}�콃���
����X�dW�2�Һ��{Y����]uƃd`x���H�.��d�Ǒ'>UȲ}�|�`�4�6	LP����]�;QK�P�RLo ����S��'�&d'; ��A�S��=�K�Pc�skʄ��0��O���*w���|x����9�����Gd���`zvss!6�mN75Q��+�.���|�kU�+��b1Z�f:B	�4��gp't�d�1�p�3ŌS��%�Ǘw0a�^�B�k�!]�U;s1,}P>���O���	e�"0�tCx�۪_h������g'p�(q���yV`�Ef�J%]�(7<�4���V�:��w�t��h��]xU2<���y7�����W���
,I�%֕cA%�7��V*> e�����J���/�"i�ǃة+�V�"dǀ�	x� �5�z�����&�njH�Ի�`�e]���P�nJt�9w:*֫�7��Ni8�*c��\1iV��>��f�t��l�vM��،����iu��NwG�]���e,�ώ��`	ӹCx���,>�@m{t<��<@sh�G���148��9��CD�Iše��(�� 롈�1	A�}��7 ��'�B�`~�F�A$�E��@T��KkjFn\���8��b�-�M�IК!�h��-w-9Eo)1%9Ax��f��آCV������BN)���a6���X�qe� P�7Yz���RMVf5O�۷�^�=a��%>��>�����E��&���n@+uk�kt��
�HY�e_���S�Pa�E-2�"��bH�ifo��I��VpЏ~�'ⲌN���X��68-��f�sN9����W���0"M���q��M�ں8�5~�4�K��ՅF�e�᧭�U5�óP+o�E*)!�,
�_!�Skw��ȱt7����_\7q�
���U�R��	`�#y����sF�)����'6A���r���~���څn(�� #�Ų��XY-���� G�c�a�cߕ��k�Yn&�G�U���1����=�0�q�4}εL�*��u@)�I��HQ���^�`�1�������|�o�w�P�^W�;=��jM���J��U$���%B�n�s�ȕ3��c9���-~C��`�ʊrZz�<�zh�*���Q���~bMi{d#]��Ə��6��zЋ�}�W,h8j1��n�h�����keA�A��Գ3������F�!+�~�,�=c�-��E�/�����Ty�k��л��	�'
J�ɳ`���
	�-��RA/(Ǩ[�9�^����^��^�L_MY��Ґ)g�bl����\'BC�|s\�dn�lg>�-���U�\V�E01��H�Bk� ��`wZ��G�EyϦ�K������;1���[H,���
qc5�"Wx�x������+���4m�Nj����-]���a�A
o�Ԃ�\i�ȥQ�����4����N���&�Q�C�Ŭ�k�a�3ޣ#��֨`���X��$������e��Κ�ϝ�!As�4�^.Q�~�ќx��v��>t�U�n0�M��DM�vڕد��3���jM�A��Bsm3�Ҏ3o��k-�7�_,&����y�׈�A���^쬤w-�)��)\�6?��&VY�,�3"��\#Vb�C���e6��R�-���B�J�R2�]���u<�n�&������=�D')�+1/n���KLM �8�&�.��Xz�nN������� `0g093���<4�c�p��;#E���D�km�\Iݢ�p$�;��2k��i5X{���ḃJ��q)ZE��k�y�h�M����j���r ��+�L�s�
��H��E��>�HU�Z�s?���^`�Bj�s����O}�&3Q^UI��\_rs�>f����C�f �Eq߾��j��j���[����(ܝ�7�@_�8Sh(�eQ^6�B�n����zNv0o]���*�n��ba�<:A}2l��9F��q�-����{"�D3~����. ?�ʦ�G˟�lʤ��Q��24/����(���IM��A/�ZT	IH.�+ ��>=m�/��H��U%,�Uɭ�V�Y��{���`�(�^�j$}m����($Pg�{䷡���ə��eq�/�bU��Q�yo�;U>�7��
W#n<c�*j��mJ-��K����;�)�uO�]P��~�C�=��!��}���X��9ZՑ,oql欁ܥ���L���WK̭|`W�����#��p�z\"�����0�0�|/oێ����h�R�o�p���7�I�q��"�����椆�vf�I��bfw������}��������OW�Bט��V�{�\l�WT�y"�x�A�p��M��q)>���ɧ���(N�0ֿa����R}=F|�ض� ��{��Ƹ��ص��s�l
�ao��$�zR$4�(^�+�c'�D��.�WBĞ�� c�H�4B� ��#֓9~��lt��b�{j`�A�N��D]X/\3f���K'��6��CC��p{�
=�Ȭ�ʘ�{A����*���n�W�����m�+����Ay�~�cҙww��*k02A�&Y�MM?�Nf��MV����G���(P��B ��\a��6>�pp:��wfmr
�,�Fe�0�eeZ�W��P>@,���v�bo�*�L~.�S�+C�6����U�) x��f��f@L|0��E�~��/�fT#�C�9��n-�u/�؅���7�y�ɥ�o{�K�]�,t�i^w����W�t�
w���d	o���:����f#�j�p���2��IW�4N|$�nFv�y�Q�olT����!-����C�6���{���������3�PE��.�K=E��&P�ސ��U )s1��f�P�0c�>��'�3� �.��+��M��T���hƯ*��U���P��
4�tո���@3JuC��Np�U���Φt�h[�׵e0�����%�7�L��`E�R!�gg�/��J:� �؃}Jw�lI�m�̴V��~�J�F���3�����K��[;�d։˒k�����
@���P����6��,�_���L������h��?!A���rO ��_.sa�
���%4�1��V�yJ�-���N��G�6��@��HJH�5����se�Vf.[�
U��UA�+Ѩ��cP�I�)�5��,�K4�Õ0����a�uc�qj��H�k�ޗ����usʒ%�S�
�(w��M�t
�G	dɑ�-*����͍(����pl�Q!�v�$��n��-3�F@���%��^C�;�E{àe�[�a�n�:�����?�)�g�n.L�T�S-Ý���y>��ν��U^�%��Ȁ�*c�I�\Y^pIcHR��y�� �7�k���O!Y���4������s3�f|����T(�ò�ފ|�μ 0�G�a� �I�����񉙲��S� �h3_���﷑w���گ��w��AH�l|�8+����+p	WBau�&���T���M��"�9��U���?�h�މ`�e�u�.-��8�iA1�[�aQ�+-2h�?�.`ԫkZ�$�R6%� �E�m�n�B��y���LS�k=B�a;㍬N�?��:���<��N_et��B=����J�H[6��.L�օ�6y�#����?��ߧ���k߉�/?�A���b\����IbfB��Y`@,n�ͼ:�H�/��_�Mq:�=��Cr1�˫ʋ��޶`6�Z@2�t���ș��r�֫���PCyoH�m��l�e����و�1#e�<��'�2��g��OE���D.��T�F:�5p����X�*C�#_��t�Q0�}PM�5��A����ƾ�8���+��ߣ`��SY5m�.��jET�����E�>PCЪ�����I�
�>�����F�����t9�^�(�־N�hN�5N�.��y2F��_g�0}���hS%��Ԓ�q���jUx�t�0/7d�Z�m�֞�Z)-��;hɝ���a>S�����b�0=Ȓ�O��%��Fz]c��#�ľc� ����b�A�MqV��*�C�P�X.��΀y�(�];&`�]�.��� F��Z�ψ��^�~I���0�Ly���)�����~��u��P��x��[����_.kߺ}�����m|��R�hϏ���3}V}:�\��" p�ovO��I~�j'�;�2�,]	�cI��b"�N"�/8G�}����R��A3<�r�n>�SS5��0��Y}C<�#͵\Q�i����o`Z�n��U ��JhO�e�1�'�-:I�MĎ�7R�	w�
X9���5	]�7\��v�i�-��w&�'<�SV��=����FPkc�2��m�/�20R��5�r%C7�F�ze�����E4���<��;��]���P�-�Q��z\�:��������Y	���H,�Og����L��i������P�r�O�B�X��.��eU �S��暬�}T���届;�/������y�d\���gҩ��ap+���k6�(2t���⪏�����Љ��M�BNzBJCt#�3��2�J�ؤH8�����0�Sn��Lѻ����ۘw��H��?{y���+�_%��_���:���J�,3���L��V�P��hB'1q�1ǜ�T��JFY�z���;��2�ph��,c��\�)Y�X�^~?7�ƫBe��,����L��N���:�n��=i�a�C�݉<�763�lu$g�0S+`�Z����]��{�w* �߃4ϡ��i��_ե�������~{vY�Bsb�#a�+�9�N���8cw��A���0�~q���em�To�F��.l&�W�"J���fSd+d�(�w���P��}C�WӚ�5�r�$�/���tE�n;��-fF`�w��?�*��>�!�gļ�GQ!��Z��������0��!>�����"b~���GC#!�e@���?�"+�Ձ�ֺ��>�/�$���*��:�����Z���N��Ī&WK�1��x3��=��xeb��G�hH�Ժ��$.�x��\����F���ŁLs������.�/y��,��3�f`�=�-{�SusZ�����tMS�=��7�ndA^�ۯ�8��-��<dK����h"\N�C�F��vz�%���8L� o��R�z����m�y���&H�����I �f(������OԠG1���>g���[��8�r�f��>���Ύ��5��c�ޥ x�}��-y)��YBg|d�~�v��Jx����S�rڜ�(]ŽϻOzg���H�h��E;�@������8�m%F���紓�	���e6�IEܤ�*� �r�:�)^a��g	���ѐ,lv��A%+y#��ʉz���h�:�\��W�1��cIIG���-�Tl�=t5�5�%o�up��s	��|�{P{�ֱ\EV��D	��b���;��?D�fS##W���IG�Ԭ�R1mb������i�o_�_i�cܩ)��1���ԯ�Uq��:�:e^��>����$�G%}��}G�7a6/Tq�B�ҷJ�<7�D�)��EOЋ����o�H���̪U���������D�㔊e�j��y�垜3��KJ��C2���%$<��\�\Z�A�Su:��C��K!�/p�*���a��Fl����/��F_�i����R<h���א�}L:w�+mMf��4'�Р���!$\&���,��jeq�x[zn��9W4(�x��\ƅ����>[�; ����dv�gJ���]�W��RB�!V�*خ&)]����OkmD�3��üA:��q������2;w��Cbڷ�a8�5�W��q�8u�d�C�Z%���[�*��쿱�jI�:87�Y�2���HV��{2��G����j��I��	��!���B�ߊ�C�@{Г����a띧0M��y�,����Ƕ1�@�ڞ����I����5"Ɉ*4*:"P��V!Z;O�A�%��hI�9]m���=�J�0�{��33<�w:vK�EZ����v��!#�Jp����|��p	��Z���e��U��J+"���I慄�_���h����u��s�3)ܕ�	�c�F(�le<A���o�x����T�Y-g'�󀙂���Ew�3DZ� ��^~a�{�R��
�D�X �h�%��KS�U��w6�B!��I2��Th�Vs����%
c_���}OX�]3'1��;`�������Ժ�_"T���[�{�Ƚ�f/����Ƃ��]��hr���m�B���>��4V��� ~�d���o��it�L��A�c��U������]���/jiδ\�uL��.��� � f��xc�W4��?�aAz�9g��3v�S�T&���o#�I�<��t]@0��At�ʘ^�+�_Bz���u�=1I�BZ��0���w�B�
8/N#Qw�]�z�bkJ=NI�O�nߙ{���l��P�w����'��ao���O���Ɵ�6!j��Ɋ�R��2T�~3�h�--HV��M.�_@�q� |}]y��W�����Ls��Xo��c�-�f��A�=n����h*�4�>)˖�B��a���2JR��F1��;�-��V�D#R�%��F56��YM�j[��¤�U�����9��v�k|�&�#G���)��A���o�-�q2Mܱ|Ar!Uc#t��ܬf �?����أ��O�s�h���m�R[΃y���)&�]4+R��5���r�9�2A�(�w;�~��"!��V�=���C���!� d�]��d���beJ����.s�P��Ă�3(f�	QZ��=L.͐zu]0���������¡��<�/�9e�U��6�.�׵Cc��M;s۝��jE���)�z�$n�@CxL���9�m���]<J䯔������̲�ד0�5Gh[n���.��]v�U�E�X�������gѩ�z�v���G-�-��2uS��0��\b�ĕ������UD;�H��%�����z1�>4���%�j����'))�\-��Ś*y�&�c�M����)Y���R,�Żl�+�= ���N$QѠ�rqQQ��hU��Dh�ܗ�}s�G�Z�u���ۈc��∣)���/�]��$ �B?\5�<����o�Qp�qzZKe_�%DĚ�S'���5+�dgW����M�3](��w��D�n|�2��H/�P�/���߭S�*j{�� �7��j]W�W�;n6�~t,�?%�K�(�ăA[���O:<TΘ
]�:ۍ���|�}C�P���$[9�7�0��C��|) O�=��� 5��u�8��Z?�٩қ}�x@=�y�ۖ�*%�,�s��(8u	�Ksw����~�9�������O���`gݿ�a����c���8*�B����ַ#�� ��vn~��sD�?������Һ��u�?�Zy��ل\�U����C��ɺ�I��Vl�:ʅD�����M�}�ً�@��i8/���]��]�V���Z;�RSЕA�����>�P7��z��
�j��c󠂙8K�8�B��gwEhW6�Q^�*�B^�I�U2�صB|f�>0�飋I���j�V���]}#������?�p�c�8��%A׆w�P;
&<)]%	�/8��t�R�Ct�L5����B�]�k��IP�&����L����k��ڄ'Z@�ՙTw�f9����jP)�HV]ի��t{,�η�E��ILw�]�Jw�XX���om��ۂ5KRX���}p�P {rR3��N_��^^x�n��ϖ�/��/��&���()�K�Sh��N����`���4�. �\��oõNbLC�	2�%����3Z-�n�8��3��_������UK���gpN4^�d�[��u��|���zL����g��An�D�7��#XO�7���v[��a�<q�H��q?�)7R�M�A�L��%�G85Ʉ��I��Umc<G��U��3DC���'����P)6������X4t��G{�Yu��eb#ữ=�m�lU�<��$�W�>������oɡ���;~hqtq���\�K������R���>2�k��z���,W�O�J�
{�'�Cc�g�� y�Ь��S����	=����!hɏ"8v:�r���r���%�4�6��쭄�����N�-�t��(��1�$kK�����wO`8Bv���q�����[6�E�?�'�-��b��È��/�G?c�9�x�S;.{�rJX��*���a,+9wɖU[H����6� ��������V�Ȱǀ��m�&v��L����;�!ɉRU�d|�h�ȔȊN���B��܏NQ�n�ю�(t����h��Ep�f	�<�������)\_��bv�(§�X}����i���_Ϧ�J�����4&��n�����99�t�eY�R e:�rQ+:+$G-d��&�W��H��<�\�΅���d,&J��;2�ww��hz撅fQ˰㐱�+��#��M���Eo~������oWJmTC�%�[����ը1~ A)|���9[��v,��q�u�q�x�Q����sY�b�Y=x���*x�qL��-�pl�r�Љy����$���m��ul$:��s�z�*X�ai[��O��Vmh�6�N9�Ն���2�VL�s��8�����&���p�D�\(��0J�ZÁ��M'�P������U��zG2%?j'�YO��5���]��MA��M�z,�d�o�IkA_$�0���~����4��3��������@��(ڮ͹�먻�O��n��lʵ�h�ô�I�Qyx��%�M^��E����=�ch�B���sgR6��^k��FdT}a����ƛ�p��W0R��V�� ��ps�u׮q=�&�X�,cϭ58*���X�YI�`�sh�EPz��Jw�������^��[F�����i�h��#�>�*VҨ�N�u��Φ�m	V��.�e|�I
 Buw�i&vsG6�kwAXfZә
�n��=��Ftl�n�hH�8�,dW����R,GX�5#��"��Ϝ�ׄ~�*���*F~�T���&�˖�m���5��Qv(�2�H��׿��S�,'�ڷ%�u�J�^N�y����H_?^��)ay?�+�1WurrQNf�k덨�C�;� Z"�Å��������~���,�!p����oc��X����*���3����0$Hz���:�r�B�(���uU[C�Cd]ц9�R1"��r��q�u������<2=�ֈc:����d�����Q%�`��m�]a��(9�(�[⁘An����i���ۗP�+r����7c�'I�p5o����X�������iM�x��� ������\M?#s^)���[}�\�,���6�>�t��3����2
|� |�6���Qxq��N\�ar�+V���n���M��"I�0�~�m��H�Z�F����J��@9�4��QkDb��K���q�]2�R���M�J����'7��!J���һh_�a��`K7�֒��௃x�=�˪�|���\�]i�b:Z<k���@_o5�%2�����$[*c͡H]�6�Cxd�Ά���II���U�+�[�O��k�=�2K׬�7���4Ф��4������ː�o�7՞{�D�0{ul�f*lQ�[$D�D�������/���.��i��t�?^��� �tC��#ɺ0f�)B����2N�.dM�K��	+Fo0�%��V&�j�JAS���dџ��Z]k3��Z7Ew5 z��d���1�+4&58��0�JW��Qn��n�ш�3<����ޫt�wL�2G��e��l��h�-�D�]|�cwX�9K
�Fs#uwlã��aX��Z���@��L���1�B�ɣ�|"&��P��dȏz��"x�b�3W��5bB��u��朂)*dGk���_�������H�4�,Ĩ���j������m��	J��!���#���2J�Ď�����0OX�ʇԄ����*ІY.��C��n9YF5��(~q �8�+Z�Iax|��0�.�H\&`DSP�n�D�5��٘*���^LKb[U��d�}�R����F�ǂ�p7���X�\=������pP���R�s�ip�ֶ���ݘce����Ȳ{^}*U�I�x���˭�=���1WPǺ|
&^/S���a=��Q�:<��@Ǆ� )�(a{'�2�Hd�r��jx2�Z�a*Q_0cY9���`�Nћx���7H��tX�L#rZ��l�X�"��rrf�yԱ�xzB�
���-mş��%g���<I����*�M	�1�͖�B�f����?���y��h�!B����܅��d1���V`�R�J�^����	C2�1�B�$n�v��J5)E�O2���,��������%�F�uA��,���C�/V�LX��`_���B�ҭQ�¿�� $���wiL�i�Oc��DɭA&��"�u�}�}�W�U�� F��^����c��:�s� �%+Ϧ��|��<���1X�y.6��O�Ij�ص�gF���4#��%@���FF��{9Ol+8�7f���в4�w4�pi�S�Q��3=�<����C��]V���ub`�1�jA�#�e.�>ȩ&�XɁ'�~��L��Fw?c$
%��a��M��ԥ�C�h���=D:�e�.�Z;j�R/U��/E����P��<�?��ũO�d菀j��a�����J��	�b��(}�Nk�o��yj���7��yj�E!� ��0,��jr���̜�4��������w��������ƥ��jS}E�D)K����c��#Z�!ij��Z?�9Yr�V��m^�SM�@qE�!�Y�1��J�ȡp��a.f�(�,���6Q%��B���J�H������8���ٕ�F���y+�n ��_oVC�l�8��g��SiQaKD�/!�~�Zb�9�5�5x�4�U����Q��`I�{�����B��nC��[@�wo�B���л
a���-<I�5���q5��	���r�H�[~=��.�%�+�k	=5��S1�D��t�R��ML�E�B\�|���9l|ca��m�x;"���+��
�������9ߺ�n�X[����|9��Q����z�����ա��G���h���lnc�8R}�?H�G��^{H�x�b�q�T^眻�(��|�&���5<��;����,�N�y��	0��t�n&1�������1�)�&�!��>n&���L!�"�Ҿ?�96���S�������9;��m|� �=�$�G����&��cz{Ɋ�m�3�+ش-�[�R�+�O4*���?�)�xЩ���&Ѹ��i����/�CSN�o* v��sۑ��m`r��Ǭڍ��յI�D��tl|�FND�)�/ޱ�m%E"*u�Xȣ%LLD�~[h�T�+��:3�Jͅ���^��K6#��T��[ɍ����>Lľ�Ḁ�|<_v>�3�xI����lM�o��K��`Br
��戙���;Ēi�G�q��r�02����L5�ep���6��k�m�ٮ�K.`�6�=^���CH"a%��j�Cn��i]�GGx�~��~-6*H��Ks����x!��*H+�N�MF�T��`��#�_o92rI7���]���*\@}���O�U�nPzi�l��M"<�<�s������m���{��N5��0_�!����ʜ	}�Z��|�A-{�U8kݮ��-[����U��0�&��;�}���1*����4��8?��L�a� -�E�P��#L�����9�q{E����@U�a�	�lf���N �2��\;g�c_��86N��G���@����NJ�l�xu4T=��O<�[t^���:�z��Y�8u�#�)���2��� �Bb��~���ƶe��MV�����kkI6wl^����:}�!|�����:�����ãH�� �Q�Ƕ����:}�L���Wy�k(W�U]�O�e+��ۙV�Ê���1���S�l����l�/�I�8�}tt��{(h��H�m+!��E��i��W�|@�F��WD�4�B�z�N�[��T�ͫ��^�7�c&`���&�VNb!l"��_��hE&�9x�^��z� �m��Ҙ�rd-�Qo��.��`���͋�S�d��F�O��2���v��m�~� /x�77rdi��T_�o����o��x���Ss��A��h'f^�<�
L�;��}��>4gE��{8Y,�OA(N�f~�h�
�Z�{P�?Q
�R�(�ҠQjM�C�j�?����H���2P���qioF�OY����gu�]`=��h���v���2�<�&����3���K�C����-���"�g��9	���|)��hB?�;�>%�O�4��4�wOj.�)��b�S	�\�	r��7^,��9ᦦqN���JiI����]��&BGy!@qW�t雁9����W�rsM̰����D3,���ڧX���B��c3��������2��AŴ��3 ~]GJ X+�)��R�é�S����,��U�����0��>S�gZ��˕�[֢�*Z;�]Ez�m�^O��Ĉ��s��ŶV���'���Ɋ]c-?�n ��Hvk�۽j0���6C��X�2f�D��� r�k�����J��,�CSM�y#��a3�&l�`�-/��Xo}�B�+(pDip��%7o����6���%#iCv{����~&�5��Nf���G9�����8͇�>ZH��+Zc��ޝM��Z��f#7�/ \-�>��] ~�I�g�m��K�M/�w#G�r}=AQln�!ao�[�`�L��l�{��P���%�<�H*�Nb �W>d�d��k�_g����G�K}}ך@aS��Ғr�}UA���Y�fJCA[�pY�3AH?��K��x��mE� yR�����s�^[����i~q�PAbD`�Wk����YA�|�\�
]�.����Ԥ�ݽ��/,��k�]6XLn���Kx[���^m�ƻ�[2Z��	���	i�CK��v��!	��/X��Z �n}D��2�%9p��F�ԂL�b�9=���S���m��r�X�?��9�@��S/��!�O�f�{'X�F�_i�آs�C	ǔ8`�]��&��N[Dl�_��{�V��Lf���[�X4����D���Y��}S�;�h� :�Q_���\Y�Ȅ9{�� ɾ��g!��ю�V���leMp�	/�u��[Ǵv�%��+d�J�7��B���J�eE���n�WMҜ��thWe�[�~�R2����E�H6�J�o;�G
��y��'~��������� ��z��b]�[� �-${X���G��/%�F�
o��]���k�Y[�b���y0��b��܏��Z�MRc���b�Z�S5���q�d<6&����x_e�a5�ѿ�栌�(ݞ��,�E����^%T}��D������c�w�z�v4 �2����aG2К���4#���T��\�VtK+=J������.,=���U��?���?Rĳ�2 %�G���?�'��!�[a���d(���b<��56�Z��F�r)�gOL.'���2qs㭩�k�����e�`��;Q8)�R�{S���0��0a�d���fX��!����Z/�VL\g�"��!�����jV�u+�?�z}�O=����^�d�O��.�܀׸����yKy:�u�$I<3&I�0YB4�]�����>.�F�d�����N\d�$���ڻ��'� �϶��yaZ���v�S����/�����>���H%���^�Q#^l ��ک(��c�7|���ݴ)��j��x�xɼu�{
�}K>��ؑ��{�y+�U먣�; �g2kއ����è"��A@���H�\��2	s�� &�P�B]��r׈�˨H��B�2؈f̦;!� �3�m��Hn��!t1�_d�'`��1w���]���L��&6���18�!\���¬�V�=ts��T�Y����X�Ԥ㯍i�z�,|Z�
"�[����q�a|��חE���6@h-��V�5>��߃�l∊V�H��<b����=�xgz�&����
���U&�lɣ��_g*  ��7AEvi�R��x\�l��O��b�U�uZQ�R����[*%���ȋ�gIա,�к}��FJ�`�$���x��pPv��+Y��ry�Q�������\�~�f��[x��3 z4�9�! ]���h0|�M�آ̭�����Ic����H�@ݮ�dO֭�ď� �`n��Y0��9%)x�K�	� p�I��	�����"�$��i�
�WQj����NNIT�1�lN����6H��N4~�7���ot}3!���?��/��C+;0@��B^c�BB(:�86�Pf1)��rL���@T�*-�b�[ѝ��ҩ�6�LV�l�����M߭�����1� �-H�w��S���Ii/� GGƂ��Izt	iU鮤�H�\����1}�F���]1mmB�$j�?V(��"���d�+����?{r�O�}�r����o�����X+1`Q{�`dr���r�X�������Q����lS�6H�ƦՁ9�pz�̽��AeKBv!�gd��Õc�.��"%lC56Ϟ���	HX�X�R4��Z���&٤��o��k�v��q�}C�קK�W@W% ���=��8a��|/1���$}�C7�-*��*B���yN��H}f�&�b�+inH���Yw��v������9����J���;Ma�;-#��D�za"�(�a3<��΄*�Jb�����~�g1��>��Cw�v�]"Qe�1(��ʑR���B�ҟ����O��v����*R�r�#��Cod���5���b���ݨp�Y�����b�A�Z?TR�i$�+�&"%{�Jw@2�xU+���]���d������&W�i�F�x�ԃ�/bx5���3a�1��fR��#�T���Ÿ�����fz��^q6B��˒�:%�?�LؘB�qt6� |��y�˅U��Sy1z̥���w�F\�oy��!F�;%��!�=Ju�oK�+(��Q�����#�X=�؀��}�F�3	b����O#[��¨X����{ ��0��HC3W��<�f���w"�CU]������=f���<S	t��io<f�&�VuX!����A&�M��Lp/%-�5�d�2�&h�x!����Z�'�@���գN�ٛU^��ܿ��n�yi�K�6�Q���f�DdD����N�acI����W/���1�}��
�I�y,�g�8���V��f}���Q�=��ϝ*�%��g�����yxf���,��<�=s����4_
���j���`n��AP���c6¢�-��;�IW]�uN�h:�^�t���-�Y8�`�$����ε��������<�$52�:J�� ��"*L�w=����|����$��h��:W�k~h���1{���I'ԹEc�~3��=��vԣ)�~9<o	��*�(���6��ő4N��1h9��N�pa�ApM*�O����]�D0�H���G�K%���0p���J-����%�x�"-h��?w�^����T��֜pD᳋���:�pW'���>��I���C�^� ��C�>�<����2�ֶ��
��b�*/u��*���ֿ�}H�5Z�fNJAX� ���sd�x|V��;[59�6��*�6�V�7�$Q�\�[W�u��j"��y�W�׋�1 *N��Əo@N=o<܋�#�eB��T��}�:!�ŀ�V�_�ʿ��&���_'����<Ϥ!�G�W�E���}�9��l���م��U|:�ܧ]��X�3���]b��
���4+u�0��olH�������~G�Iga��d77�z��'{���-T�q.��4���Lk�H�����q��؏�Gd78�����feVn�?�뚱�-��"�{O��A[z?l�k�^oM��������	W��#ۦ��vU
�#<1��jq�j������������,���?0��HO/���R��e{��O�Ţٖ�8��%�M�?��-��/5%�[���3�g+D�,C����@�a�Ğ��d��j�A���e�ۻ��bGf�NwԦf�4Va�Ct�+��PH`ְd[@���-=<�h�ۑ8��I������Ε�S���~�H��s?�?�+���sZ��SP��B�����Nn���!��&=~d�$�����},��ԮJ̍Q��X�q����n�;ч�.���S`y^EsV��%�T�ȩ�ե{�*C���;�g �4*H^,���#^�"�i��3WW��O`n�@�g6Pm��UJK��Rc�!۪%@
MQ�����%��dS^/<}�exk���z�Z��|j��y>���A���QHY��Đ����;��(�ou��lä� ko��Us���� 1��Lm��jU��J#C��P;�8����|��?f(�$\���)��$T���Ss$k�4)��$2����yFK/����u!��ṋ|=�p���P�{��\1�߲�>���9a��!kDX��g��s��ͦ��p�YH�	e2F-�v>�-rsp�_�����%�����7�5��w%,�GՑN~�m�.�V�̝;�����������cH~�{l[�1n%�zu�=����@<O��
v�E��D��MC��C��@������f�a'�m�E��"1������e�ς�9HN[�r��r�
@���po$JgH"0��9���y��8�w��)+�kFY=�Ѵ7�rR�d,,R�ӄ+*;Ĉn�ǄOl�e��v8,�X����NH�¯j�WrĶ{j�d)8k�{��;UfۻUd�fG��򨵗��l�:"��x���~��d�ġL)lm3�W�q�<}��,�|��D���u?�Ե���^MZ�h͜���pfG-76y�N�r2\"�5y��F����W1�4��� ��U�� +!95��|�8����Նq/��\ڽ @_������␸Q����:�2	���l�JcT*R�Mb�\p����~}��j��;�uc�2���| )���<��~B�E�������ؖ��)NT[�DFEn8�Ww���K���!0���"*i�|9��B���.P���-��ļ��r0$Y�Iǋ�Db&��uϤ�T�����(���R�$Vҋ>E����[ 5%�$c���4I1b��x5�i���`t�X��b�}���Uav����s�E��ǣ�-h�G���6A�p?�$���%�+c����s,@���4j��� �\�.��Ұ�U�ffx��~�a�l�%Y\�e��G�~�/��G�����&U}�0��fV���nTc-5�Q�6$j�k�8�D��HZ]n~]�X�&��aT���jX_%&�W[z����N��k�\�vٵ`�#���	��i��<���C����E�����Sl@�:�]���:��g�J����f�V�5�&�8E�������)V��aR��b�D`�*l:�$�P}k{�-z���XK�N���V���&�2��@P�����-�c�z��jؚ�9�L̶҇-���!��н�j��KGl�IKf�Y,�� e���� ���oѐ��J����R{�v��$��� �¸؄w� p���A���J�R��O7�ǿ0��������ͲX�M�sr\ޓs�k�r�k> w��k9eY���M-
b��p��������7��^��x�Y�{���*����H�c������b����WG�nL6�LB=.^�{^1����?�kcx	�64�Ǿ���ˍH��!-����X��]9�Y��]]^H�#+7!�2r�8'n��xD>�de��li�URk�D��(i�6mCu�t��s�y?��V,�U���C:3��j��B�'}�pIz���1qɬ�O����Q�U�m�:��$SƖt�@.F�3L�?A������-�zr�_���e���c��k��Vl`�2���
����J�KX�&�� �����;.�)��~Ye9��8.���F�}o$���_iZ�l�+T^ǋ���3` �{���[G�Ik�������̱�E���fU([��9��iÙ��z�Q&��j�P��!�tϻ�� ߑ��vV��1B0Z&rw��(qi�%��_�����Ê�vzͺ��/4ҫ��x]H���|# �G[+W����9�|5L�;yC�X��
Rc#�w����'I��"	��r������r4�F��5Svi3{��_G�����,_�F����k��xm���A�s���uOA��xd�}D�ޝ}YѫW��C*X����ݖj/��Sƪ\G�9	��iG5 �֓ӧX��e��7pMf[�q��ޔ�!{���$Fe��G�񷨦�ν����MYlf��}���*�w�s�ƌy���z|�\�T���t_ ms����l���E����
�5�!Q0�;�7`�
g8łh����<�[�Hh0_fD{�>�!�J�5Ņ�]�Y��N{�(���|���&
��`�����7�IJ����u���o�zH�Y\�����`�$vC�]��&U�j�y�L	1�ǀ����/~i�ߔ0��J�A�V7����(�[�o`0��Ӡ�@�ا|�B�/	쀩d�7����ʴ�d׮}بǉD�I�@�7v�l^\�GSQI���[�W�����3��n˒�-�b��/Jqn��w�*}_����3<Vyp��/��/�ӶK�]I<g�5pT���ƬD<�n�A �#P̛'�&X_�cQ���%�Z�";<�'����?�����B�M���~'����o۩��A��=�Ц�oH�K� ��T��p��m��PY��G����$T��;�Ɗۚz��|#�/o���EЀ��X�p��ƣ?�
�2�g����l����I.Mi%�u�e���?�A/�[�s�O�~���y2���2�{��T�C�Q:�����&J�.�펞_�o�ᒒ��ǝ��b.�^Sw\��o���Q������s�$_˰023�1�!��^�mN~wU���k;8)�x�W��9�L���f'�?1���Z�~P���a�}3j��MO[?�����
���z.F+s@{6͒vk�z�gܻ�8��8��bhx}�\�'R:��/�{Q\���˱�͋Vwr�U5�T8��`g�YUx���a��MH|�1���C���p�r�CuG7={.#�Kq~�jMcuD�βY��7by-$i!�l6�U��n)��D��@?�S��6 ��9��h�49����p���,�ܭ�w���	�b�n�yz���,�j���VlRz!�_8��l{O�I��I_��/��V4؂̗d��9/I����,�F(�[�L�H��ʆ�;�N��N��ն�
='o��Ԡ�?u���!dFȞB���Z��;|�����`Z�4����M���qd�0��s>w�iՇM���i�����G�������Y�����NfS��Xz=oLj�S>�9�-܅�cF<-�o�)7����풧�I�/'ܽԅ ����mG:0�+��18�U��ǾP��)�3r�TY�p�A8��`��]ۅ��	+e�>�3�� �3_[ s�E�cG��@Ԧ���X�
�-���N��7��Y*��O<�hK8@T��D����b93��z=<S�A]Ɨ��6���z���m��9Ad�w�� ͘"�`�������<�U3�M���"��[|k�f������Z� �.�́��L�0>pa�s��Ml���G@D�9��� gFf�AP�g~������M�k?��$�
�vy�Wrx��>ଳ'�̚	Oa.��S��f7�q��\�(�B�L��Ua�&�b��-�fޅZď�C �4H�M�6��e'���t��~b�h�I͕Ip�?W~���ɠ��}��ʲxr������1'��|�b��Ĺ&����A�q�O</A�qL]�9�׎N��&z)3R�CXԅ�5[Η��o�8��W���4O��v�Wأ0���䃩�<���y�ڇ"$N�o�n�YN
��F��Cr|�~���m�� R@��t(e[FM��Uv�n��ė�K��R�c� ��30����nb���I�P��)�z�y�i	�ks�d�f d�mLd\��K~�������kU�\�l6G~�L��H%�u��n��ZA�c��"Y��I��ǎ�&��ٕB}�+�S1��A?��X,j8�P�ôo����ޮ�'����2�;�� ]�F�~�f!��.\^�C���E��.H0�LE�"Q/�C��wT�$�2ܻ���P�-����`�Q��Т��*�z��P���M�\��P�N7C�%���1��Dq� <h[/�.>�J%�;�4�Mr�	�Eǧ��]#ש4��k� Ng�}�z�����7��ۜ��+qH��؅��dz��A�t9̯\�>	���������;{=Oi ֲ����O�2��跾:@�W�,��?6B 9*Ԗ�E���O�j��=:�+s���}�F���^�Z-D�;ן�����Ϩ���0m`���ac;h����|8�u8�Q���*{��<
�Q�1��B`uJ{3�+v�a]�"�XD1���gε�,��a�wE�9�@��*�{�����
M�	IG��s ��dwK�1�M�B1����j��߈�F��h���^kh�1̞�%}�:�,E��woI�M4կ��w�>��8��OC�	�j���]=�]O�l�6�����V�3Y�m����_*h!O���և�&�Lr�H-v��,�*GC�iڻ~���73��v�c`V{?��6�>&�p��\��與ŭ���}e�(�f��1_"���<�K�G!��rCn�$/M�p,��rdT���97ˏ�Ӎ\eF{oL;Qr�Cjʟ��%����vψ���Q�x�%B��,XO��v�V����tb�dʮf�a*5�.C�?V�.Y:�ԗPe����Fr�~��;��}z��$Qu��dRoE�S���"�뛸ς�aס|���h@ID�c�߶"!OMN
2��l}��[��o�� �X}��ǆ���}^D�f!��}��R�
�7�i��v]yM��R�ޅ�ћ�I��� =Rh�M�=9*���0�*
���L�徂w���]���MJ\��`��B�U�A�]�*U� m���35t�u� h~����@���h���S���jk������� ���s�QUu��!UAH\�7k7��No})�>���5�v�ٱ#�8����"���U�ʪT<����xD5�pY7~yh�i����8�o֬1�T6QB���5�aɖwfJM����$��b���_'�]�����\�賲��WI�jE�����ɕ�q4���������Y4��rM�6�O]p��7�{9�D�����7�l�l� �l���},�0[+$	|�����u��@���
���<[#��ǩ=����5���V��L�!WMk6������=Ru0�^*��K#m�ygx(k�V�O�{8*)��=2[�Uٵ@�N>��U�p�Y�h5(���Ҿ���&V!Iռ\�ju!�h��0#E���Y�ฺk�ɥ����jh� �ı�����7��5Z��N{�N-���\	�	P_[M��(Nm(���oZuO��7-�Ш�?����|M�.G�Y����63uU~�6t�e^����i��M�|��Euhnk�ZB},\�}�'*�p#��Ŭ�^g�}�nQ����p����~k�Ky2��|{�z���Zgul΁�� �s�tZ������ѝ��vWm�1�7�lq`5�Y� q��W��ӌg@	ExCFu7��<
���m'����]L/�b�]3��g�|��2�jG�F��P�J��R|n�@�V�Fv ]�{�	&]�f��K[:���:��űe#*:*�����K���OWo(pe�."�[}�9���u�P��{ƞ�]���~kX�u�Eo��ý Y�f= ܋dα��C�c��~�mPJurC��&�Yh�ϛ߃����O�p�F��N�u�š`/�G�������D1�5i��M��0���˼T�?��0�`�2�ư��e+�Aè�,v�<s��N���&T�6��7@X��`k*'�d�(�K��/����Wk(Տ\�����.5���l�o�2�Y/����^<�i) D�Gp��,��N[	A�O:Avn�HM�ܬk�?�B��w��f�6sߕ�[4����5$b[�Ov"g��6���tZ&�sw��;�h�Mr"gI��� �܎�N��Ed*?���9��#��5;��j(�۫��9��a=uڬ��&7ӵ���2�y��	b���|�?c��>���&�.�\qVZ{�.x�Z.�ED��"�&ħ9x�&�SB�y��ۜIR	ܑ�P�nGD�V^9ݐ��L,���遘z_z�iK������I"�%	w�$*�K�g��?����O��J�O����8W�%C�w	=���VH[���U��^({O�+����F�iz�+��e��fO��N5�l�U��ty����\Ƕ	��l���jȲy�^��@�./���\��Q|uO s��%X�C���Q����T?b^��&	�K<{��D�r�b����G�`���.}0bV�\]�J�{�c�����c@]#X��};z�(;z/_w��̀&H�5�v\P�Q�_���l,xҳI(��6�eDSK˃��"��ۼA����Ga�]�k�|0�/#B�=��^�u��%�,�3�e�\��X^\%U�\���5�(��8
���I[C�Y�=MM�o1��ǂg���u�2	,sϙ��O��H��=��z���-9��!EI�/�m���� 	u&��$��dVqO��8�8���^�=>���v�<�#D��9�&U�WT�>�ސm����+2�f��Ǹ� ]m��q�=)��/�Q��-�Pu~�b"K$l�co)����z1x�|,br�
����D�:T��.��т|U���:�^>�a��S���7}SG��I.��1�O*��2~������[_����D��З�AP��}��k���&1�.�Y5a�@��R���Im+jRVr�&fxPͪxo�m��
�̲h�l�44��_C���|_�1v�����Y���-�����Rn?�V��rJ��w�,1��f���p)�]A�m���pD�(_��������l{��=�9�7��;z~����b]#>HA$����]�I�@�,*ե�+�-*sjpDS����R��!�n|zkE�}�!w`�|S�`b�&�e���ϹX"�vh�4\Y�NLD����������"�D!�11s�<�e��۶]
��n�Ǘ�A�s���?��&��h�1���4��������;#g��
k%���������,+�2it�*�H`r���\-����l��z��Ϸ1���Î�����L��{��s��Mc������ߡ���*e %%�O��ؤ��aY�O��砥ju�|����*ܓ�����i���5���gݩ��As�I�x���%"�����]hD����bLM��}����!wO�扅bzTs|��A�^�j��"��ky�ΐ��jܛ��w�B8�c]D{LpT\�\�Y��$`���[th�R�xI��>F\b*I�Ak�!�0z/1�.���2�m'�m�~�u�^�wn�`�����F����О�Sz����c�ԧ����g���8 �ܼ� D��Y��6V��0a��	0�Je��������h�+ ��0K�\r y��$`m�̩L�g�����*-Yǐv8��(]
;1.�uo�s�����D�����B�DݲdE�#��W��L�L�Vo�}Ů%ۙ�����{�t�c�݅k���c�
�z�bѷkI�l�9lK|�Ku��Ŵ���٘�޺�XxA�,�����d:-�,����%���E��I8'Ъ_�o��p=�$�"�i��ttڤ�}�Ka����^خQ�,�cX�*n5^r#Lă@�|�XE-/����3$����^�� ��Tܹ���
a�ú��hT����|��k_|3�ͷ�_�4Yb+(�hJpEQ��(_��P���.d�Ȑpw	���Nv�/T�
Y����r������@c[�����c��~�:�Hd�^k��jZg�@�o��	��-o.�����qH T�.Jv��>Œ��Iӭȫ�i��E���o������λ�X�*���v�Hf�,�T���U,P�	&��K��Z��\�3���j/����-]��>='RG�!d�`%|��]�Y?;�.-S�H;5Šq�k���t =v b�vb�ė�A��E-��� O�<�+�9��˕�'G�.0����Sec�;vѳ"8�E��&8z�S���_ �asF��xs�`�Î@ޖSρ��>�o�#E�b�>!�|WxP��K��RzJ���=�*����h;��'���ׁ)Sv$��8qI$��d{x7��e�:V��<����#kyJ��b:��q�s�!��� oSEmȄ�RD�%��B�p˔|-�7tZ!�G����4��pB���hU�~p���L���o��fb����V��щ-���V;�I�ͽ|���b��������bo�]H/��=�d�����y�ZV?�F,�br�~�/TD�E01�{��|8� �)^�w��\���R�b�Xɵ�I��d��c��qF �i��hطM�T�Et6�%p�+��~�1�<�֢�-?�A>Yp(�4�[�NK1V��@����Y߇�[*�#l�7��m{l����M^� �91)��ߍy��8ܱ�1�m�6����+�x�3�7 s�₄�72$|�ِ�	��;������E�p�PBp�q��.1T�Kb����w����x&�,��-l7�G��#U�'Tb	��I�H�6��2�6s�gO+uK �h��1�p�sI�č����7P?�°���I1%�z�H��n�T�`�;��҃|���,���^�A7	
�,��X��77�
ކ���JH>�{(�]�c�a��,����7�\�m�,2$Ð����*��ۉ�|Q4�;E�!ʓ���Z�G�-]�@U��o}���b����i��}��E��%xk�}��E&NH�mo�v�` ���q�R���qL[mʸ*�<���!c/��*F�!�Q�C�Ƭ%�8�z�����&�����Q�����Ht� �m.)#��l"�	U�E�F��-P��;�4}E����v�j�F�����^�gu���	8Y&��adb��Q)c��AQ�B�A)�#a􄣓�+xV�^X��=�lO�B��w���I��@c�)�j��\�0����]�i7#g����p-���J孧�[C��}����@rv �|Ι��ZY�1�/�K(�m�A		9y�@N��H���W"1�����Enw�ը���QfEJ���^}��QL��[����'���&��u��(J3L�_�C
�,]�����Wf#�:JV�������Y��2q�Oh�C��� ��q���;����c�\��S@t
�a0�*ܥE������w~��
�Kߖ��<�-�VY�-�V�F���!�More�t�`k=�,�Yl�<r�G�Iu��Q�g�
�3���3'G��0{�E�˥Ⱦ���Ŗ�:���^<X�Eê�Ou�9p��ClJ� 0�N��B�>>�e&:�����7b��j�����_��fH�@ɥr-I �*�R�O�>������h�wA��Ov��gM.$?�18�Z�Q##xCk>Zs5�G��p7L6Y��o��D:=�u1d�yWG/��>Ey�zݿM��̸t����E/{YQ��.�>M�'��(���H�_�K��Y�E�A�'A�@<��33uy��%��g]H(|�ߊZR�ϫ�"�K��*�y��e�¼�ڪ�ЮH�҆l�"uݥ8ej��b,C��Y*�+�L\��]6"h�K*SM�.qUmͫ�X�nl�2��FNM'���Vw���l]*�an��{��&�k��b�|���ds��Њ�ƶ��ǆ�9C_�	��i���"�&"1���b��`Wz ��^�`f'u�v�����<�^���O�(���g��̅��c�y+x�2����׿:�S���s"��񧬳mS���0	���V������<X糠�7�h���\���6���2��>�\	�/F���7qsyB�k�w��h�������j2�'+�
�ưׇ��#�ޮLD0���M��h7�?ʁ�l,j��m`q�B�v:�dS��Q
�f�Ra<�#��?�o��8�[q��VlN�5v�R���`����D�+=���B�+��p���
��۔��uqv��h1��R�2����M,Z��ȑ�cb�1z����-�qE�Xc�!M���C#}�$C;���B�}ؾe��:r9���;�C �b�*J]�XbS�Ne�sd�Z���Ԯ=	*&7�W�H	��	�*e��������X�����cQ��T�Fmk3��D�^4�,����Œ��F-�=���bW
T�8�*�*ȃVw��B@�ɧ�`|>��͋o��wQ��&|����6�%lTx)0�3�ߦD�Ti3��E��
�ȲO1������B5���m�C�F�����]vj��8
M:��/y��ѿ������:JdaW%�p��CtAA�$J��>�����ҵ�����aY�^��Gd�؀�b;���Nka���"��N_�i�0����Oz�=�Tϴ!:��׭� �0TPȶ頨��t��E�>՜A���A0T� �:��Qn5M/by���bE�O�_bY�,D�+o��qF�M����N8\{闉:�1/lx�o�e�S��э�8�]�蟦�Tke%�O�c��f7���VZ�M��%^���,�H�D�Ckx�O�»���	�?�G��'20ʊ@ε�>&j�hZ��4��C�C����hm��8Q��@D����*�A���}]'0�_\���7�(8�Y��'X��ڛMC���+M����h�5R>q;�z��"W:Fw��C�ڮ�dq5)3sv=��	9�
�&��W6�>��P���^xz���#s�����OB������p�s��s�֝	F���ϊ���*��$$�~U�
���E6+��n+�5�:[��?w�x�'�R��Wr��:.�}K����x͎�ukt���]��΄��:�U��t���
(Pc�Kv�4�`I+��. ����E
,KwoW����J��H,�
�H*�j]ʥ�8�]V��4/K�VwF뺋k��!9��˯M�����
�W���e�{�it�>97&`�	�U���=���r������ �51G�`��7IG��F�R�! X��NH�3z�ţ����D�d=m
�tR�e����x�|t��)��뼂��z�˥a���e���8��fK��A_�>1�|��� ̃�y�`�G��)RB!�i�M{���5��y?l7�I����cx����&�DᅎRA�u���P|)�2e�篪�p��� ��Q-���٨��} �<Я@tE�,����_	6#i�.x���Z�h��:�L-Xm��t�Zwz�y���c����0�jz��:-�r͗O�I��a����'�ͦA�]ت"�؊o�$�Z��}��.�C��E����T�n�a�1ш/�Z�[�j��I��QO��:����V��.7�qW����W'e�8�Nb���p��1�q�
p�vYo�5��-?x��A�C1��.L��F�j�����v���κ�F�q�m9?��r��:�t2h��hx���%�~!�[�����-HN���i_�8���'���yw��ne���v%�X7��˽��FY
����K�T�#���X�� lg񦇱>h��K��� z8W�i�����Y���t*\Ga�l ����ҵ�����æ���T�4K�V�i9P�U|���(G���N��ر4�L�6���)*H���,�DHG�?��1� �2X�ޒ�p��R2��L�K�����4I���a��S!<O��V�U�3�	p�Y��jp>�l��y�L�������2d��S�ڃo�v�����BNޕ�O�s�vR�<��>�~-��ś N�Jn���OAfe��:��gp�>o����y�ֽ�:�ޚƫ��t�IW�pq|�]2!\����4$��NO�9���'�ײt�­Q�n�W�14߀��Z3�2X���=�����L������?�'�rQk+l>�s�N�u�,����!sҖ�Jf��C�ZG��.��,���)��z�б��v������5���(0�q!���jL�|\�!��T�S^����IČ ���i���a�!�_NN�-Ѫp=�F1��jJ��I���
s�"߿�E}�w��4Ԛ�aT3�x���P��$���=��M(wc���;=��8�SU����§��I�l*�u,A7�&3D<o~�8G=���.�|f'�O�]��|���?�a2�>�`�pK9�
8o�Hg�c~��BpL�>9����=|w�`���3IZ������:��J@�]��tC�w>��_�y��*��<���܉�/�4
�*��`[֩��/����f��.7��0�����e����5��}�2f��8*���-	��9$4��d��ͪU��ѧz�0�zA��?8<�$�L��$�d\�ݮ�W��Dsg�m»E{x�w[��&�G����1{��5�L�M���/�cQ2z��zI��o��c/@R�Y�U��3se?�E�1��8��L�"�3�0)#�#����x"غOc�/���X,˫tkq��>48i10"��g�S������@D��\œ��Ǯ2�v9�^�ʼ�������	��M��_:J��¬�d�}#��I�"7����hs �PG	��u2�>������Nv�LM�"�~����RT�rcO�3�,�0�{��6�r΂FhUoC��LR}]���9�Wnڰ��n�B�v��F�~q�} ���+��k���(���̺|��������Bm���gIs�Yɧm;h��n���ro�6���l���K��sx���Z�H�o�[Gpk�R�
ט��[�7(`������������\�h�v�I���F5n�g�Z��A���[T}`~��Q�ӥ.*�C@�u�x!A���"�2�)RJ�&��ek�5�CiI�4��)��1��o�����pZ^�Բ/�&�"⒳D��Sq�i��A�N�C��A�@�wس+.�|:��.��GudH��?���r�"��d�m�t��C�j��S�&7��?��xQ�ZaG���ݲ(#�`ʺ@"�g��aT}���I��٩��h�[��tg�s�dN��kՃR�Q�O��Zv�/F���'�(ʏ�h;�u�����}T��ߍ���������D�J|��-|7B8f��7}�Ezt�pK�K��[��?��&g"����C�;�h�R�|��﨏��vCc�N����`1M�i���or`4e�T�?Ets�Nꖛ��������j��JA�L��5a�٣��p�6��tذ���� �[��|��ޕë�!��%]���W��\��p!���2��0�9{.��_Pf�S�!��p�O�lY��@�2E�~�q
��o�^X7�;d,��w�|%�d������=\CG�U4�9BPޘ������g.qb�X�W��`�F��
!:��i��i�B������_F��	���P�O��Ru�P���'i\�J٢�ΣXG�Z�K�?�}>@��}�����+�SY��5�T�nw
��)���o"����zO`��J�d4zq]��
�x�|�|"Y}M7/� �'�3�P�t4ƭ��tL+`Q�BL�}���^�9+RTĮ��E	��U�Q�;7����xr�G�������e����?�@Ϋ������Ȋ��i���aP#ht(U�i&�^�3�
��� ��h���������q��
�YL�^�[.-<��Y�{�3�`[Zߌzg֬���v��/ު�w��=n�>��`�x�k��Sz���s�1���+�M#�����z�f�Ky��r��>(�]NW������P�3���m�WSЁ���tMlyϭ�j"�G��Y�F:o���Y�`���x,-L�Svg2�� ��Lx.���@�I�(�C`>��� �:7s�������>tp���}
}�T�m�����UͶ��O���s�{�����a��}�Ge���V�Ȳ���#Z;y� G�b�=�)�f�s�Z��E�ju�>;�0�`}��}���؇��Hh��ly4b���t��^r����;�y�����N�1��vՁ괙���s'�H!iK�s�b��m�T8��7���X�%��������QC	�ob*��i�=0��~�ǫ���`���y�b��Ƨ\Ӌ�s�c����9F�1Gml�c�h�žM��nlm'�y��A��L=��X�l���X�9�HxI�Sd�L ���]?�����p�=�%���`�$�U����mWbS�H��b�����j�b���<b|}�KK�Y�"%�u�ܬ� l�<C*p�#�Z���OO�N�[xj��,>�z��Ǖ�F�t���4��`[�x���na�ǡs���?�[��֪�g�u����Mw�>��#�͞/4�d��(g����m�Hy�O�o��}�}\�`c��+�:�Ho;�uT]�7��U�K;b����ɢ[��et�s���X,˭A;KL��!/?�L������ܚ��1�9_��$"M�J�yN���a��l��8B���;/�2s���L���U<jە�X��P���:�X{=.yI��:Hd�������-�e�^�Y�&5��l�@5��EZѤ�;ns`��E�[��Цl@��m�̼�X��!;Fp�5s+i�媈�S�3T��c����'ާJmd�UŤZ{$��� ��u��FfuT�:i��3LZ�7�;�-�#�8��eH��j�sq�6&`�"���6߅�� ��@3o	|�&m<�l�QWX�`eΩ�Ⱥٰ9�~i�X��z<�b�]�g�[���lb=~l���h܏�.	���mz̕�uu ���vq��;��eR/O(����	:,��j��l4�����x{�r�m�a��O"b�E�����GmC%�֪ԧmCݯyV=s�Č���̴.���5���_��:�Lm5!����1L�8�����D�k�?@UY��ż�Q�:�Kf̈�(�giͅLZM�1�y���> ���'_�g���N[FeA<���+�և�^��������T!˸���pN�.�\#��X�����d?
V-ȕOt>���q�;Ϙ�5�z�av5��4.���F!;�5~ o;�y^R�Ԡ�M�Q"(��wX|j��H|��a�K<7�|�6�
�@��h���)�:�ILlJ[�_V[����9��VP@���cC�/C}�阀��m��1�}�_�p�0����"v�׾�$T�)1>�}c�]����z���`u:�ul��h�*a*CҚ�`��B]i
�WY����T=��;r�b�Njdy����Yׇ�� �@J�%�4����q^�C�%��+��h`��=��3��`��D�g�6:RS�X�y��~g��a8���|�0�}>�B��d��b2�F��s11#~)5���a$D���dΉ�~<y,A����Ԗ��k��7�B�v^qf�y�2�5���Y��;������V/u���7ٰ܋.���L&� �a6��a�l-�v6�h���u����5���@�B�G�����NN�{&H~2��Ce',[��Q)a^��_�ƛ޷��\��p�g�}fl�������%	�`Ɩ��� 2�9��.��In�m��R|�d�g�O,��+��%}"��(v����ZP��O�?��5]��l���T�`�� x�l���x�l]Ɵk
)ww��/��՛�>���3�,a�c*"M"�=�^o���z�1�*�̔|�tXӹ�젻���Z�-h60		v��O)3�]���i-A���Cj�����7 ��_sV���h���H������|$=+��%(�����QT��Q9�fP2����V�.�:�z�p��NMOWۋ�̔Ba��� ���L,ʳ���-�c1�E��勵�[7n����Π;!��V��C�������(Џz� m�Y�*��]�f(�<�`�S"����b�~�=�u�P^�f�~��,��'��ڥ����j�*�_����e���X�2�ܑnu��A�'��dY�H���WZH�wm��yQ���d�<M�I�q���
�)�U��������*pW�VW�V mP$`�PC�$��q���Q�^��`ۑ3�����VM5/�}3�<"}�fPc;��$��X)���l9�o�h.���db��U%;�$R[�Ҙ�6�h1S�b�X>{/[��g�L�cUv�
� Vw����Lci�I�߫�-/��P�gl�<�Te�?'��L��e��J�0�' #���,�0=_Q�	`O/�ar@��R{�B��eepϝ��ԑ�����<��[M�Χ�f������v�- ���ݡ���O�?:�^�M<��<*��������Q�� '��ܺ�)"Zn���m6(��
�6�1����mh�G��
е��jY	1�i��ZgB�]׌Й|(0.���u�ø�0l\0��,�� �"�ݣ�$�#0���h���l��y�|���@'�6�Lԫ�p1�~5���/��b��R���C�6�T�߀��8 �kO/I���V���5;��#Eq��;X	�׋��Za���M
�cS������L\e�t7�G)=�ۑ#��� /M)LX�� � r��^�(���6�[,p�|��\���ļ�<��=�,s��Srv���,�mТ`^ꋹ�H:&��#`����c路�vC�o�ql�4z�rQ�a�]��ڴڰu��0��Yt��%�x�����l.�M�n����Å�Ñ%:��k��ϻ�@ǫ��@��S�2���%���U�O�G���_�fMw�+�\��N������1��ej�G ���[�>�F0�I����ҢL�C����+���(ōe=��8|�U2[����^-U����*�����m����32׭}^�e]ܣ����ӧ����j����QjڂN�˪fqڽ�t����+�7?��H�����L��]r#j��ڭ� ���[����Y�j؉iu��D�eV(Ee �q�
����Fi��+�Z$�$
�Z�F�BR�]��<�ڢ9n��?(⮄6��[�xPz�g��m�{��UAs\�!4�V������llj�sd[u�ײ�/��sq�?��q%�$��}� ��
��4�"�́d����P�9��c�4����c
��Q6�����9���Xi(Cl�Tp��C���������W�"+,�d�:�L���H�:U�}��Ƞ��Cp�ø�7��r�DOs�/ckS��� ��o�5Vc�b�(��9�ɪ�f��PRW�ܡ��k�hxĨ�S���Z�!�wF{��Ѣ��O��ˈi���&Ow2OQ��6k�y�>��&��2���q��1�&-l�"����XfJ~����ˊ�����fR��S�L?UB�<�^�km��Wmڝ����w�`4�,�����/&(�����<9P:>����/-��*���2$��{:쿯2�E&�&���fXV=�["K�����r�2g[\@�9��#�- �Nr�.5�^Gm��\jx��%��&�9��I�5�P3�/�a*7�Z��z�����ʠ�$0���X���8���N�Jf-$�ET@<�J+����C;��2B�m��d#lW��fљ�)�'�ԥ9���]�s}\��2	�M���>%|���K~���+'���Nl��o`��$~����O�s�6^8��ז�	�t!h��yT6�:[�؏M�8�J.����4�	����w���-6���6�s��p���۟��'�`�y�@4l��r=+�QԭI��ƍJ�W��,�����T �"S�kWy}Oz,��NB�=h|^qz��漌@-k�)IK��:<hr�$h��o�$�!���^=Z0��ܻX���vtr�k�3Jp����7��^X0�o�2�Ú9xn�A�K	�j��Hצ���
1m�L��.����$�ފ
AC c�
�i�J�Cm��+�ٜޕ�+y#���ξẂ`�"�yG��=X�����Is��}��εh�O_���V������M��qD�5�#2�ab&�-Q��m����Z
��*��@���ы�G� <�H�S�!%��q
G��*��fC��á4�ְc`7�?Q&q��)�k������O R�Jի�8vUE���GtW~�9'��?an0&����w+U̵k���,�j#+ow)��`:h��B5��r����C4�̈ۙ��:�.���rm=������k!E�]����o�}�����%V.Zk�U3� H���ԎC^��A<ΰT�ڲ��۩�6�nȕ����o��-u�
��\���A��{�4��!�������X��	(��hO�g�B��r=���->�7�D��e��)5M���s���\�#2����}�K�/��l�ժY� 2�R�>���.V�s^����f��髲 L�k��h��>,ϭ��8�<d:[�4��TIL���ҕ��� 4h��g3��R��C�"��6ϱ]t3�!t����nSg{]�	�N'T�C�E�0��+����|�3�������S��8��3>*[�Ȯ��R�L܏Q��2H�;��y��X�'ƈ{�9����IꖝӴ!(8���iы/jXT��G�TT
W�Y�
VD���z
#U�C�"�������_D%A��i5R��(�9�gd21zi�~�)%�./Vq�es��=�'�*Q(MJp��逫NSI�̘�xkUg�Vl��+��F<0�1�&�"X��l�Q��K��Hb0�is¹i
�T�SM�]�Q�8=AÃ���Cx1P��ܛpT�T5�e�P�E�j8s@"�$���N nga�(s{>�����Ih5f��g]�O]�0S�l�cy3�~69���~~��.!� Phm����� �i�1���>Pӭd깮�<si�,@?g-�+�_{P(��l��}�KsDӲ�ߙp�RS�e�z �F~ͱE��F��JM�M��T�	�`�#]��"ȟb���IaO {�Oc�n]����3>�����#[��sJ/����^�q��vdCr�0��9�ȫ�<�i�����(�͆6޶�'Πg��b��Z��v���:T�O���P��{@�t��f�`C ��O4,�)��8�����׹��b���0|Si~��`��J�
��0�V׆�3Uj�0�Ӥ���ډ`� ���Y�Ҭ���s���h[�b�kF$�V����MEQ>!�c;'��Ο����3_T{�e�ȂͿrӷS������cb�#�%yKep��
R�_th��w� ��#P/��VA�:�������P;�wE��o�M�:e�JD�=���;\�]�����Z.f �3Rt��J2�e���ɂp���N],��@zT#�����+@�>��t`ϕ�,�fC(��������nU�A���m3�/�_���\�S{\r޼�<�����:s,B a�`K����O��)E�&�Y�LR~b9C�c9*X��?d|��5l�j9"��6ș��p I���㱈�׊��b�F�a�9�B�uQ̨1��w!���c ��G8N7�;y��<H�s�X<ϧeQ(��f/Ցҫ�"�D���F�W<�����`�����&F6��M�;1&B*�*�st�;>��A�����0}�3f��dxQ�m`�$ 6�{ b�|�A[�q#Q�x� Nv�d������l��zG���B5��`���p7�jy��R��Y�9^xr��Ң�3�ޱ,�AF݅a������"������&��/Զ M��y<q�ԟ]�k�.���0\����5����9��E���F����J�I�¹&r�уK���%]�P���k�JK�����G	�-#a��[ F6��9$)��G'��"�[���(�ɱ�	�V-F�1��L��A{��^����
�����%�}u{nM"�&#���/w����-~a��gU�HI��a������es��Ԇ؀��^2H��/�؊#_���w��xlv��cr�  \�$c}��ѡm��"^׾H~��v�hdp�,��'<*r�,�XY�.KcLag�e��]�D
��B�B�~�2�}�yo�	���Z�oŶVF�VZM������P`�֬#�ƀ��\��s_���jZ���_C�ӌ4h�!+�����U�#���MY�����n�:���yn3V��d�`�����G�6��O-N����	��Q�A{���)����e�؟M�Xbk�GX�岕�hU<�ڹUH�F�k;���=�_���j�.m�V�W̒��D�mv)��#��gr�r�AX0,�>�~��T�H
�+�!�au�_:�|0�9ٔW��{�溡h����:5�����i��$�rJNxG���������
�A���(��3S�7~���Yh'���a���䷱l���Be5�X�Ef�J�fj�湧5��싏���j�^0y`az�>�쓾�iVtls��8�EK85F�;T��!E\�1ZN�p��<%$e�c�z�+�G�Plv6��k޲3i���M��^�V�7�ٱyP��Fw��m11���]Q���T.�0����CN? ���hO�KC�����C����x��J�[�^���/�#����(��o5�e�Y<�{�°��p�Ff�w�Hy��Xw�����2���Y����F���|�H\��@ p���X��	oN%�9��������mw*��$#nYaC�D�YYr�w����@�	�5?F��c`�n�����LӍ�K�D%��y��S�-�\X�k�'ܽT��
�aDk�i4���^o�mRL���o��fo'�A=�T�rM�8�����/?�e�yy�?Җ�"�Dc�E�(���+vZ��L9RD+ �XV5�!��80G>A@����aA8N��z*��V�F�N(4f�b����ӬS�θ��-bH��s]���dv �N2৶��ù��_����zf�AU$E�ޘ1�	��J��3I5��QRE2�H��#b��b��Y�ּW�,菉X�e�C���i����£�R�=�	C�A���8'*<�/������Z̡v���]b\"J��#;IUiwQu�Ҧ�x T�悓c�O>=H?��=�iK�f��Eku��ΟTs2��w���Q����?~:�՗ye���VQyA�I��D �qmdgh�s�q�?}�/�@k�{�Xb���!NV�kr���lIe|�� ��ĉ���\z��H�����^��7���Ɖ��od���*�5pw�#�Y�����ܙ�X��j�d|�������G�3��2���Ų�c`Z�Q�w��V�uAe.!�@voU��fP-V�f�̔��X\*s�Y`"HP��*x�00n&�}�X���(�V���ER��$�O�*�գpǐ2�����V�7��I��0� {3zs������%L�����K����>c�ť�܀^눨�U��&~�@��vD���9Ɏ�<��v=t7m�Cc��4���Ԝ4�	�؎sPg�}����{%�\Z�R`z��,�3Z©���-�F�-O�������W��\]��xIXju5"��!a�+�ܙ�ߝ���@�g1��$��p��,���ED�n����-��d���D�Q���X��Х&|���b���L��-��u~������ ��x ;�4.� ��������Y=�4����K݁X&:��xt��l��y�z_���Lj��T���:�����7P*Y:)K�5���a�$U󡼕2L�tA�T7�7CY�%�h�)����ƈ�S|km�7
���#*ozj������ �d/qH�t�8���(���d��U?Us�b�c�Z`͈~�+�!/l�=[W\b�$�tn4�Z>��o��|���A���{_DJ�I�/n!���Z�;��P�g���Hp:���60{B;��㽍���5/S��%����t����������p�<�7�i��v��N�x�>�_vguE	g<"��S8j(]����+���踕��c��>�2w)��X��!Le�LM�����wK�6�Q��	�l�n��J|5��/y��|��n̮��dT_v�	_j�c��-RU�TNj��QA��l]Y]��9[^��������`�P�zL�i���J�G������Do:�	>�(����С/��jc�?��@��[_/O>��li�dP@�f2U?���J�:ң?/��έ�`��x�Mm�6>�Rr��[��4�>�i1� �9��i�ol�N� �q
��s'�N	��l{5�I��r�ft� W�No�ɖ]�rG���꺭[a�Q��,�Z�6u�n�4�콺㼖`Ըai��-@����+�~�*�`m�1�SS�Mdj��.��'n��vy��
�'���t�V���Po��D�F^vy`��Rw2�zV!h道�'s�v+lt;��%α�
�x��FT��u-ax��>e1b5�-sM���r��ߌ�@��T��f�W8��W9����ȗ*sH�6�U-��?Ÿ(,{�B����@�L`7,>2��XBjs>�Ҋp�m��@�t�9s?�H���23lG �wkw?������)]<Qw
�!� ����-������Wo���V~6x�?E�.Z���E�-��).NJ�{x�`Mb��!���)R)��;����z�V�*G��rY$�mֶs/i"���Z/��3��)���"���g�
�CY�j5��pΧ�
�1m9)Ro������CO���I���>���z&%ך�AcB@���A)���e�-���큐 �I���2������TW��D7��\\ZJ�6碧ʝ@���H�N�$��p����d�z��ɬÌ�Xi^�R?Ƞ�)�nyB,�8�%�t�~����9k���m��S��Ţ=�X$Z��pЧg�$ޒ�H�P�ۘ�Q5�����YM�����O�T7z���Rp�aP�k9�z��p)�RgT~K8A����]����x��,��2?%nXZ�*JFl�%/��*�1q�\	�=�RUf0��YG]0r�;`�p��r�k0��.��Q6v�~�8����$
�-͚��H97mw��I�:��b'�s�iAސvc����:�T���~ ������ԷF4�%�CT���F$���pgΒQ��.@?M�Ǆ��M���Y&��~kW�v�������"�ٻ=<���2d�i��׌ ��	M�4�Z��r�L���QR3��\�6ͭ*��	X�ZvS-�(? -��Ƅ�\�������R:�Hg�62/%��#��2~�ScС` Q�M�Fd�SK���r�Aj|p��"6�_��_�p��5I:�����3%��ma��'�R@�u�D,>/8_����k|���$�`���Q̜�7z�� M��MRB�@HƑsX}=�����2���h�"���Y��O1@}�&�nѻ�?��B��h�����[Ig2]�L3gp��k���\VN�ABxq�Ds*�D��5ś=J� ��w���g��+V�q��:�cĴY���[�}At��M�*Ii�*Ӑ �iݨ)��_��,CK2F΁�:��Ó�|��ғ3�I(����,2�yDr��io	SgKf���:����t1���O�G-��?��*��0��HR���Z}�c&����n#���YP��fq��f���z;f1DC��9��m�P�%LO~�y͖�z1�c̚9&`���?�F)��sfk�0{���Tr�ˆ���q�jO���)����Ǟ�5\A�B1^�+E2Q��˴C���|��FthLl��
���ժ`�������<b��j}(=n��<"F��E����*��:��,I�̔x���1�eA��D�������4r��t�¯����ƃ˪��*8p��8�hGo�U�U�O� N��2�,|՘:^ӳpg�.�Ը��e~�3�w:[me��a@7�D������n�����
�XW>�>�Bx,�ק�G�8(�e�'o�)��B��"��-Y�v��{$��T��i��fg[�Y]�xO��V�H�V)�@!مj��j�^Պ��=�g���2��F�-9xdcq�^B��"⭿�l,
�u�Ӵ����������{�v�,�4KD!!.�(�l���qe��TVէ[���:w3�L�q���b�+���<U��"X́d��?~��`֖���A��:�=�I�k�%{O�f۫	���H[��l��%�I��k�6aD�YK���~A��C�f\=��i<�0g����T�_6�K%�"+z\����`k�,c�nC�J��U&8�S�l����S�����9���ES��&S�5叔Z~1x=�{a�	��wG�{��T	s���̞�d��_w��mR�!9r�L��Ȗ6��`�SZ�^��;c��;w�^PR�@���Ą%�8�g)yo��sD����p-��
�C��Dhg�Mk�ߛ {����^ˆf���OT�dF��؄/.%eeWv�Ĥ�ǆ<�I�.Za�j��x��Z���_�e(w3������ԹT��!�=ϫ3�s�3{�
q�ܝ�Й,h���ґ�͑X��`��d8z���'�fb6S;ܟ5"jv��Iv�yl���I�S4����p�ն�vuY3E��7hɮ&A�,i����J~k�2�Z�O\:
��� W���JBW�tWA�e�T�����MeHU�����?t5�/�U�r}�uz���E���L�'�`-�*)��}Qj-Cȧ`�ɿ�-��KX5�0,C�+n�V�B+��ۢ�
m2|�x��-"�e��S:by�y�Ha�;�g����.�o���2�0�%c�+>���7ӥ7J�y�+��!�2 ���#��
�6펴Ԟ�A#A�mCfW��/ٮ���ϐ@5�4�+�$�"0�ɓ]�3�:�W���QZ@�&�=�Q�^���	l +L��Sa���/?QgF�|AZ�O�	�g�e�9��w�o��{h�X:��@�*��6�n��8A���]tי����)��H�~�ڃ���/Ğq��
�xeR��4?��N����vU&HZ9�%�lస������L����F�Y�E ����A��:'��x��w�W�K��nt"����R��9-�ccZ��t���Ԑ�&[1�ʘ7�~��9��t��w%�*��&lHMR}�d�h;Y5�w���xq��.�|y�l���1>Б����.������켎?�b/IN�Sdb��"�8;�d^�7eΣ�ei�6���"8��d%~1<��}��+���-4)X���s�ֆ�N�6U���nM'~�̑�̍
����_�#Ҳ�dӦZ>D�NA|Ȥ����bI:5��5�.=~�u�V�I�t+��'8 �$QK�䦡������f|=5H�`C��e#WC��]\��g�X
9�:G���c>�Da�ޝ�"������y����D��Hb��uܻ���L㤘G�B����6�2�;s$4�09r��~E���X����[%�xa2��Co��\�+*�,�� �h#<�>iT�Z3_T��!�[�p`��XoJQ Fh�U��h�,.P���[;
n��(�_i � UOm#���f�	�N{B�@��X���E�e�HM��{n�:'�	|x����D�hu�){�{\�����O����������]��M-��Y�Y����Ys0�&�i�����R($�n�"�;t���M�z2���d�m�-�N6�Z#�\��lW(]��oaM�q�%�����uϷ���~��>�xU/�0�	�.�ü�G�����P�b��,U#Τ�*ɩ�l�� ������߶`m4��l}���z.�-�u�C�Lp��<PUz�W�J>
k	�;�N�x<����h<�Z���ѭ;|2�W0�ǗT϶�zy�1M��9�o�yx�ja���t�s�o���=*�JM@|��W�hH4��{����xF�45o��ԧtZ�j����)�[��Hv��D����?(���y��:���Qs� ,�N���)�^�%@>���ۍ3�YV>_�EYm�/fj�Wƌȗy���J���Q�`����8ULd_o��k��!p/r\���~�ET��$��A��q��*V������\��c�J(��|K�:��n�ûy��N�աV������mh��9Q>A�*s�ưJz��e1�ìxo�>�;~������5i$���Po�q|�8h���V5PR"p��\ya������
��Z�J�(�s�׼�{"��n��E��6 j���i�7��}�uQP.�F�s!fp�Gs�ve��ם
Õp$���(�(��t����R���/��㰏�8��"/_���2���lT'4Ҭv�c���������	C��Z���P ��]�w�Dƿ������9�D�@��b�A�b(V�&OO"yb�)��=L��;/�����ͫڥ�*o�%`�(}���[��#G&�Os�$_�*��'�		�������mM��F�e]��x��h��!�2
ro1���	���@Nl����t�4<��ة��F�������̩�
2�G_jڲ:gd�����q�JT}�S9�դ�i��1~������A^��Z_v��zeQ�N̠�v���2r�,{i���[���A��8(jl��%�B*��>�cp�����Se���M���(��.�������v�N�B�<�A�8*�Մ�V6$��֤�{L �	�J�����L�EH<��5* zM�����|��)�򪷤��"�t~�%�=�0��!��/5��t�O�4�Mɖ����x�ܓL�)�21o��c���v�*�����ڷ�9�f?��:���P-rk4�&��2�����G���0=s'�T�(&��j!$�
��d�;t�""!`4����=�yRe��Aዟ�����#���J��8� \�>�Fa�0!�q�	��C��H �e6����˲3�����ymmT���{0�[�)ĺ���`=<jka����XBz(�*�+,��ӫ��n$����z�ة���#�����񵀟$���������ۂoY� \J�̸�$;�T�}��*��Y�a6__7�����jP懒{�xD���΋��x��d��4��������j\�(j7<X�]up�F�/�Qs���
##�x�s�4��/y/��h��b��f&��7��W�g�qm|�zK���| v��>*�q>��j��3%#���n�d�����x��6�	p/R�M�:��aˎ��uY@gp�;{}�p��i���^�
�o1w;B ���kri6�|��z��d�`1c�q�x�Izg����,��CS���w��vX���>���T]#�VN�2�_��)³�b\��*� �8��b{}-��j� :H\!���0 ʆ"/F�ԧǼ�KD��Y�3���\i���
�q�@�焁���l�ݪ;QFtQAGθ�?�4iq���q'����Y���J+g�	^����=	�r��x��}~���J�3I��ٿY*Yŝ�e��?p���ǯ=)�X	��E`]��䄆g��\��q�j.��ӈ5'��.6�eޯ��������
B*p�;�9�������H�Ck�eQ���zm�i	�S�յ.+CN?No���x_����[E9��Ln�Ȁ�����g,�@��s.ۆ�hk[��A`b��#�TA�4�_#F)_+Q��q�:��]����
SڠE���\�S��J�:b�ӄ��:�(�#VW����f^�r�Q�P(IŢJz��6�M�Ex�Yn�ވ�3��#Z�3�1����oGeCp�+�e�%��0�;=��8��aOM�!���F�����4���]H�G��s/Qɲ�S�g��u8�I��䶆Hg�����p���y�r��>���J���"N���(��(h\�?6IG�Z���A'�8��yjF.qV�N�ǵ~�M\�Ә��%*/�9O�x`��I�hT���I�c��Xn�k�a  ��bHkĹw�� �#r�,�ٖ�^0Fi��{�/���3�b�
�Hef�k�C�d#�+���5A��+2A�f�[ذia�@*�.I
b�6��'�%�Z�5�1���ce��l���)��`����M�ɲ�d�A�"�G��=����q-jm��iڹI��4g��_�!k�Q{@��h?=�Z�4�;p|QB�+���<�v��� T���0�Gm� ��H�l<�o>X\+���͖�<#  �|Lnw���%(-�5x	.�7��(1����ܶ�X�6�&���_��g��� �1Z�Q$��
k�:�|p�O/ɱ��2r���f=��5��J��>��5�� L�~/7K;�H��ڊ�$���@]�P�SM�+�ȃ|+������EgvZ+���i��{��A�x����<��c�հ�E8����3T�bxK�yQ�M5f\`G����G����D�`Q�IX���'���V��r�dnD#OB�s���۠���*v1�s0��{�������'�+b,;��u���_��`>��P��]&�o��׆ 1��Ub�2:�H=�2BX�P����0�+�"ʄ{I�ݎ��G����o'�������Aы�"���1؏E�O������	�5��M+��T��z<v����M⿃�����'|��xD�7�$��
7��Bl�q�rƣ�:(Qи�yM�H�r]w�֯��?.��L��"��kkPYa(]S.e7S~3l3��{)���U�	�	K�������vb^�G�0����
�Q����B�#V�yU�%�2��������ZJ���wp��O 1�����,�^��A.�}�B�~6�f�M���������.����ٳC�޿9_"��>q�=���2ft�졟�S4�)��G  0w4y���(	��	�o�����c�F�������DK�D X��e�8�����aB�ϙ.!�{��͝T�VL�i��!6f�k�Ph��1	|v���9�����T�G3�)�y����R�w�����_Щ쿱i؎�w�.\R�?s���>)��������ƹ�+�oX��2�`{������f�:'��h��*��
��*��iF�^�������,v���ɦ9h��N��.�h(�h`0f��X�hK��ȅCp�5ԙ�/'B+I.-q�L�f�S�4�

Z�����#���Ӝ�]nb�ߤr��"iA���d�Ld�1O�	��Ó��YT�^�Ue��U�oK��4O��B�m����|���`�TEd}փ�c"{�o�5éI�L��N�z=���<�c�4Q`Jކ�iɚ�J��S�Xˮ�$������a��e<�U���W�=ρ!�b�R Y����k��p9�jk�}����^v�$*j��:��_ _��b�9��]10�;�9d'�� 5�p�l�!��9`Y,x�^���s�g*��N���שƵ�=ҟ��q�5Tsi��^�d�	ߟalpo拹|366,X���j���2�R۹���] ��j(z�~${�kl���m��%wI���6
��1�x����gPh����eSc�խ�BH�>M�Q�S��a���KP�<�6F�d��&��zb��Mh�q��L0�2��e�`��״.Q��a-�r��B�� A+��ăT����R�kщ��M�j���ܼ���P�����yy��e <@�d�eK�'�]�E�g�8�ةxZ����B��CHv	G�%��g�s׼Ƽ	����OsC!ó͙v#�	���e�A�ߟ�|����;�������m����fF^i��x�,�s���hV%��� �L����n�Pb������|��� ��G�~S��O����oKq�m��	�n���S��R���2��'+�O1���+ѻ�������z]ϛB,367�xY���n]��Pv^��7��q�Eu�xA9��q1揽�~mE(T!�z�qV��˷�P!Y!JT���|���X�DG�3F�8P�����>d
T��H�1sB��3P��׺����C�"7b@��yV�"��,�M�۱
���J+�����1�A�N7�w�^����Đq��u��I!�uw��exS~l�Ar�L�
>��
��������+�rp���*����m}U��e��]V�fAKW��ܥw\,�j�LぞcI�e�^�Qu�a�R��u	ۚ��q`1{8�)5�N��Ny�_�18a����;�˴��:e�0}��2^�P��@w��0��`3�R�y�s?ᘤ>k;��/��Q:L���O9Z��Lّ���i�:�y������c��=0�"zf�E����n����:��[�y������� q�)Y���3�̭5� �0�W!C�l5F�����O��ș�Q��e���Oh(��os�Ӱ}f���}��D�	)�)�s�a^��-_ ڱ@�z� gJ5�P��/'7������GHi@�Լr��E����Z�ҷ��H�x�Ž�[	�p�|ܖ�8S�'XQ�i'x�{I}V��?�/u>h���+VY��|�l����.c�S|��2'��C;�����	7!L~d���%'���e����W���\��,Ʈ��mԆ� c;�p���F֥��B ����fH:��m����ZL��WX�y�"j��a�_�����7�������$���K���aoK���v�ەhv������K��e�*,�B�M8t��Z���Ĭ�K��
�f�+Q�<�!�tcQ쫞��|�?�2��V}f�W��&�Q��L�(����%�lO �L�VV8����s�(v��zw�sÇ�{T~λeV��9$�U��� V�2v�d���L�)w�kd�:�f�I�E,R �����5,� �N& ����U� �����*~���f�q<���XfKH��~�)��>�[��w��iSs��}��
��0��&A�P�>��yx(d]{�f�L�X"��Z���$���q��Nt`�F�n���,_ pkS����O�ְ����>߲ͫ�GF�P]6�$e
������5�m�����Qqg>��k M�?���.�V�6����K@7 ��ax�[D�O�����e�Qථ�
��f��&A� ���%�OTi���'�/�X�n�Y>\Ǧ�>����7��)+O�vu=Ax���&���k���Jجd��!��̦%Y!�M*`�"7p�.�m:I��wuv:e�O����2 �v������)�E��7_H����Uo �'Ϧ��Tghx�8/��iv}>�tR3F�7/�x�NFT�Y�Y9��c��6|}QI&^�58�1of��D����mh�W���ٵ��*f���q�=]��#<���7����⮤ˌ���J�n�KǶP��(O͘I�"/�A�^|�(�I<�kNT.�8 �,��Ω&�c^��}f��zD��`O��}&HCW���h67gy�^��OI�\�C" �T�v?��U{�y����v�&�o�%�FM��h,��wm~3��]�}�IJ�����;��Ou��u5ڍ����]�f�pu����Aё.��ˀ�x��=o��b��ݗlDWJ�^^������g����}S=ǨT��1p�/U��)�rHے�����l;�b`��qr�V(l�~�,����k�ODa\.�,Cid��H�������-N�Z��e�k�h�̆@.R\��H*���,����;�����*y��
:~z�!^E��bڔ�Z�#urE�b1���&l�:��5���1��/~�J.0�����>��yέ�dQT'�v�0��B���������N�*oqp��h�ק��,���*�h뛐h	�G
��mU��Y
أSNӪ��bR�R����0#6����I�����|lӘ!�����c3�����w��4�<<�U�r�,R��ψz��|�D��˾�~��p�-/w�4����9oJ�d��=h����=\3��9���<!�M�H󳵺���ߢ�=FpQgEj�H=>&�@��qe&�s&�k��^Y�Z��h���#̈m�%źL=�.��3p��E ��q�Y��?s����μ̴n��x���1�uW����;�o��&4?p?6��7nbRG
B�|Z:Ae�>�����:lN�E&���5��^�5�#J�-�j�t�mw��=�@Y�k�l�x�b����g*R��K���CS�^�� ;ny��k;�zޚV�eu���K��a0j��ۢZ
�2d����;RGqs�"��K�3�)PG��Y�#���Uw%F�F�Y=��u���5�����.�ƻ�h/�O�U���2i�֘g�N�! ��̰u7X�%��$��GmH,uߡ��9Z��9�|v9�����)#�Q�q��
+�N����j	��Qy���|=H\��{��>K�a�5��I���r��#]��Es!lXV���Ό�As�q�[�cr��{��~Ӓ�|�mP7c��c�7+�pɦ�Z4�A*��2���0"SCP'���m�,l�9藑:�N/�7Ԅ6�Ţ�m�__�B��sZg*R��ʰt|�G�p���\A��ܘ��sTy���|jr_y�rˌV�l������a��`��c^������v�@0�k"ZE$�P��.4y�>>u��2�������Ƿ-��G3�<ЮD(��}���y{�}.����\�S��}���D�VËE׏��s�M���R��h�O��F�.�c��֊���v]�^k�V��&��>o)�1?��߼�ChP�)W��@e���WЮ�/g�.�9���>�d¾�/[���wy��0<u��Z�F� �b�O�E�YL��Bw����o���D�J����f��}��D��n 1epyA+���~���V��_�EF�aHi�a�]���>"��-�����_!�TԬ� ���s�zWLuh��i��l�c����|�qJ,6�Cj��#�Dĸ���U�k:�%�Tl�汊�ė���M�6Z�>���F��Y�e}׫k���m���<�q���߰X�u�:{+�.CZ�mlC�>��MZ��������.���g����3��nw��d�E�'\3)W{�E��臛�'�)]�p�SN���g����6��4�!��,S�`�=��F|>}Ƌ�ܫO��J�@�kC�j�i~�-N��#A�7�j�Ԇ�/��L���bY�	`F����^%Z=|`+�jY!�&_����tXJ�ϰ�7�A	͒�a�rM��!���eu���j�P������1U�	��S��TC���d��4�D���YV�>��ZM��p�.뜃����������'�l�ƺ�ju�s�c ;{n�tǣ���{'�a������X��b���|9�]�$�_<��JmnL{�+>��7��dG��|ĭ�i�a��)W��n�m�U�'Q��������Y�7�h���v��3枌�3�mw��ntW������#9��~����7�{������7u*
�H�[A���:�S#$�!>*hUg2�h1�U����f�p����-��Q/��P����4���pP|�ݥ��6�� _��3[{N�t"�*�h�6�d%��r~�=�J-5@HYj3�Hkɯ�;ȗm�.2���,H.�G����[,$�3�!Z�ұԟ�G�qH�Jz�*&�,3F�?��V�~O7�WU}r�Zd-2�tÛ�����������.��E�>C ����/�gFŚ��g�_����Cj,ᆧ�U���2��uv	�m6����h]/�ڎ�<f�0��0�j&���ya<�G��/�qfe��r6�_��:�kD���u��7.�`+"�T��]9���P�@�[�%W���L����Ȗ*��D���-�s��*�9��6��X}���[`��nE� ��-6��i��sX<�g����m�Zx��/�3��&�Vܞ*����'���ڟ:�O�j+�;�=�ˤ�����ߦrOq6��|����1F4�pΈ�6��[�[�"X��Q��,��(J�rw~Ԟ����f
� F>~FؙT�'Bu=�:��s%�|��A
I5n�Ay75�q�\���|u��͜��@X^�R����r��)ZbE{Εj
�\�>������B�_��!Bbd��|���$��vVҜ��D6�F1�!�X5(����U��@����}��q'�%�b�(��j��V�-8�>:��`ep�/�>����΢q�E6����"���^��b����%���x�Q
 h���b@��0�4`��^w�0 i�>������7�c�nPcn��qey���yy�>̋C�)_�َ	��Z�~b�%���y�����c6F�R 0`):v�6��(�1�D$�2Eu����k� �I�n���+�9�;-���U�z�B+�ig�e�x�~^b�9��0?]����� ����,3k��k�����ƒՑ�	r�N�8�f�Gy~��C�}���L@�w��rh�HY�����%%t�ۚי�Q����	s�����O|;���2bGk�v�}�˘�m�+V��hU��F�:��7��)"Sؙ��sB� }�4�V\��w_�S�Xi�jn�@O������7 ꊻ������R����_k��Bש��ĂA���4�`�v��<E��R�,b��� �-h��,�}��(���"_�9S�	����t�:]]�ĉ�Uب_'"w�{��a�	�j�0, ���l顚3u:�/����%[�^���9Dֽ�tU1H��_)ڢ���gQ/����bp�8���/����~�7���kq�'#A��޶	L�ˮ�����g\.��B��A���k�{U<�(�r5A�˳b��X�S>������+[���Ni�ɟL�Bv���^���7�>R�����>�If������^�I4�����!D
���TXS"��U���7��J�g|��ޖ}c�z�!l�a�
TVe��K7�)��g�
��8����C�0io6���رݫ�tr<&�w�"YNXC)���g�`t�+l�H�y��0�Gj�lP����L��C*F�C�L�IK/�tmz�h2{� ո���⅃>��Xb��P<�ybk��9!#{xY*U` "2�L F۱X��F"*K����_�7��4���`��ʘ���xf[�D������S>Gw�Fn�㲴�͞��"%O�W6AR�)�W���+���J����7�S�N�;xU�:�Д%Q�Yw1s9����8s/N�������5V����tg+Dcb2p��P��"��8����������W�2�*�`�/���
$[��C:Hq��@WH�=������|�'}$m����r�"C(iH����/�*��&}*.I
1�ƍ����oU�V��( g�[{��(a�s]|��x뛗�(���N��?����jr���n��^Q�	;��=N[��,��Y������������A#�Z7��%6'C���NH�����"BDK�j�q�讁��C���]��upp|����@9s����Q���}���_ߜQ��8d�r�]���k͟F��q�n�r�ȣ�W��EF��Д����>��v� DQ��u���D��"RG�x����iYuG=�J�[?��c��Z/"���T�b^���N-],@�z�ip�slҙ3�>���SH�3О�>�A��W�x�3�����VB������3���^�;��QA�9�M�&^��θ\kjќ��ŋ�����(���|�O����bǯ)�N߹�ڨ�Ry��:|=��k�r�).i����,p�M3<������R1�4#g
m��gsz/>En?o��4M4G9�%=�}XW4"��<�e6�w&lRkX�IG���H�׌7���&+?��j��?�z��2�	,%�����8��:����G#i�H���\�Y��[#�o1�0��M��'o"hP��G��BGO�C����xY� ���|u���m\"6)�=k]؏,�P�v�G#�vJ#��u}0���~��PH+?��)�aI�1�s���tS�۪
�
h�j�š��O�l�B�� y�,�*�ɨ��G�_��a#^���1mC�iYjFJR���ex�>�Sp(s�J4Z��s���]#�2s���y���+�S es�>�nUf���X��aDI{�ӽM�Rf���|P3�g����`sVaJ�3|���&�F�d e�<�	��<b<	��) ���Q=)��#�4ą�+A.���O��b���fl��,�d1������Tj2���tN��<���)�Ij@��L$��H����pik� *Z��r'/�GҴ䠦��h��8/��0��h�.%�o��6|{�y�G�DW,�$2�0H��|D��nh�y+z�8�saȾ:��C�}}Ϲ)��"�r�_*7�\^����*%l��p�X�K,�O��\��wI<�43�Yޗ�n)���(�����򫢈X�F�J��|[j[e�����1>qY���"3��������Q�˞���/��L�'��T.��{�~}�seH�ZS\��j���[kPc���Ə����KAf0g�|��Zre����A�փ�'L�m�E��1����3`Z�m�F���7ep�*ߠ�P<�5g��vSA�w�*��<��?*�$N���n����� "i"M�FQ�KzS%�4�P�p5x�/���Q�R�k`1��.�t�.%}1�����2���R��h�t�a9�=��gI;:�{��{Tޙ�2	Eb&���J�M�V�]�x��S�O�+۸5����^����w�D�ɬ��9}T�ļ���O&3�����'�-9� |jZ&·�~��>��Q�)�d����)�r���b��t~E�Vd�^�
L^@����+�݃y�|���ש�����qw�*I�M�O�_�O%eN\!�1ޡe�P�$�q�������&�a�ן:?�p��>�AQ:]��u؀>���>"^���_��_Dwd�B�RQ�C4�ܪX���#�c�E�\9�-M�]�J�4d�;�cg�?���گ��k ���Ȍ�����ɲ:=�Ra�U�??�8.^�m��)<k'�bj�QH�0�{	MS�썥��w��mW��@��ձ�2+]Y���9�B
v�����F<{O���\�S"N������:�
l�@� ���R�k��fv�nNͫa��7�W3���u裥{m��1�o9�ya��/��"}9!�uF��炷�r%Oa�M5�����,��+)��\���n�
��u�R�HY���r:%;������ФO5�k���P[��e���%��
w��C���mw�O�"��y���O2l��V�ƨ�T���<�,#))<��*eg��eB]���Ĥ9ǔ`�h�:���;��2o��D:,x���:2�5�Ս1[y��5�֗Jg~�N	8n�:��]��x��{���<��xyC���Š�q��~��ΐBŎ�+�I|�� �����]92
�xd�875�R��-���)>l0����̶�'��sG#��'�Z����bp9,�17횧P�K8��w�V���{<�r�T?x���G�dvsn�������j|��q�'�U!,g#჊�M@���̿6�j]�����awj�FP0��k�-LJ��B��	���LѮ����D��	��2Y��@/.n���|�fվU�$���#V�P�O��H�u˒9Ǥu�넴B���B��4���>��_���\��$�1S��<�}�Dwn#���5H`��h�"��j��+#��߲HV�]H��Ҋ���OP,������X"J�j�CW[�:�8��n�X�.r�W���]�=���%�;f�tgh��B>�7ᨁφ	Z`�'U��vr���[F<�،c,a��k�~N_��buD�([�q�{��������YztZΒjE� ��Mo�E q�@C��78P��/��˄��	��Nؿ�d�=O�;��kc%BܵƸ�����ٙ���n E`�l���䘥+�wVK�XD��Q�}jc� �ka�����+�a��S���[N�<�&�N-3���ٙ��N"Ѫ����)p(���K�������0��/E����y�	O,p�Y��?Ow5	��v��n_�5��4�O��O(M��9�5�s�,*�p7�FaZ�;�ܷ*s�}��@'�&Ғ����G����I�Ď�	fB+�~�oGN�p�uQ{���s��M٢����S\���B[���($�Z�;X�׾�6�,d'�f5�s�)^0M;�|�?���U�R�Ah�^�T1a��{�$�թ6#Jf�u[%^�Q��R]��z�}Pdo�(NW�T��!�XM����&�:g����oF#���0��/0�	қ��ö�H�4a��zɛB]�(�t�"#D0+��؄�`�F�Ɍ�U�nވ*��Gvm`�8\4�1��P���Կ)O	����t:�&�z�H�����5F��8�m���Ӽ\RV(�-�qћȕ�~1��v�O1�?�E��%�x)D�"�*�8��ڽ/4Y��,2a�$���%gA�b	�ąY�xiP�Ah�ǽ�P�Z=궔< 4��K�C����d�K�!4p��@��W�	M�;�(�B�S�/���h�FlQV��$}D�W���K`H�[�
�ס�&�*����z�V��0|����ۦC;�lh%+��P4�?	^����~7�7�[ס��ݵ���Fo�F���U=�Y�V�  |����??@��ǖk�{`M��o�ꏹ��o��ù>M}]�m#_�@m��O'Z42�	�h�9Э����r�����C4�%f�|#b=���~���H~?�'�C�C�K�ҟmI���a��0�w+�m����fF�� G��^dY�'���v�e?Aѳ"#S���x��/I�2.��՝	��U�4�2���O�Ϥ�/�t������-�Z��@���ݬц�e�ڤ!.���I���$ݱ UY~����Ԟl<�O()���ڷ�����sN�#�V������}n�kg�iҡ�\A����ڧ��5�K�+�f����(��EY���MA�X��+L���\�#+�u�@F@�;A���������wu2h����h���CX��o!�?��L'���}b�RyW�C��G�
s@�0,B���4-�Uv��#�*l��X.�I��T�:���a^��D�#* �VU����-=͗a'5�d4l����	�7c�QNJԖ�]�lr�P�<�h�V�
��S�@UKj��;ٜ�w?�"����WҾ�*�.���� �`-����B��h�$+�p׻!)o�t�u��qv>ڽp ��Tzb��<�G�?54>�����Y�k;����W2�K�B[�9SJ{�'�����E��k9�D��
���Vdw�Ѣ���P�6x���{O"te���3H�V����`��Yش���F�>�5ʕ�@�L��2o禟8�n��)�L*�hǌ�;v�0~B%G�bn_`�Ԯ��g��&�Կ򤾒tFy�8��C�W~;�w-������'S:�����"�����W(b6��^_�]�MVD��0 h{�9�g9�aʪ+n[���� %t�?$����N��<9i��bdg�Ƀ��/��>����L[+��D*��]�v�X;�8��Qd�B+�P�0l�Vc��
��K~�E�L�&�F��y�]����G�\�v3S�5rO�������D�T0b� ���%x���\�:nvU�~3
Xk̇�����=�h�gC�I����S�����R3��|�����N��I
uA:��]����CĤ�`D��B�g
 ,o)mfA����qF�FO�g�Ch��83���X��n����xX��z㱅ϊd*��i�Q�K��;�N�7�k;��
��Y���>��A�_H�OoH_s�P���:���8(��Z�,���dT�)F�.A�"�Bȿ�:I��ӱGoR�ߝk�]�"���]s�ׁr�+��Z����m�;�����8���P�g1@��U�k�8󆀊o������&�)R޵��	��ᔞj��4��GX�#�zݴ}�ηg��A�Peqc��xƏޗ{�,��\����镑S����k�k�r�\���GU�����Ę>;3 �'�׫���4<V�&��x�O�i���cDm�@��r�iaۡ��{���ȼj�bU�d\�=�SPz(?�>�9�٨q}�ë6����_�;{+~��Q�b2��/A0���6����*���85�WU���Zgn�2��zL.�>?^/a�KU�ȿ{��^��A�ε
|�kk�f�͑�*���i������{�[H��2!���h3|�l�I`��\�n�L�ذ���Ķ�b��F�2t�k��c������鐥+�8j�H�x�ׯ�t���N��B �[1�d3+��Z{O��/�>(�4�&��l�Y�I���$V�zQ��tV{����˩֪�bl����w��� ���Da�V	��jl���F-����"�Q#\Q�@��ŷ��ᐫ�)�?�@C)'Bਰ������Aԉo�,�\��s�f�`�w�{KNo<�|1˔�~v���-�����P��w��V������
���%����>���N�G�D:�����~?�DI�sE|�scѡ#��J�5�&?q���8����u�SdF��sjtbe��uo���M���Š�J��ӊ#JCnv�j��؜
kcta���dF�^��me�\f�$:�AO	�o�WS�ٍ��|�آ�8�6_a�Η)_%���(ޯ5l%V:�H"տ�@�{���Ōlڣ�-�(�C���,���y����+�)?_PD�t��K�Jm
�>�"*0�������|��T��r��S��l~}�}J�8\�m�So���y�!�Y4��t���i�oL�+��Ļ�E���[��"�ݖ8�C�}�����J	>k��ɀE��@2�}����6���lJ~~����Q��[gG�!`t�}�.N�2�}k���2|g��[Ӝ"�>�=�W�n�6mO�&LTo��T��@VY%��?��;�&�]�=	�U��@

u(NJ���Q`����))�7��j�E�\ox��&�&x/̌g��nd<�Ċ ��x�k�܉��>��@�n{?Ҩ+�Ix\?�x�_�>M�n�y0��Ԕ�!X��Z�ה��]��%���3`iO:?_��Z�.�D��	/p���R��#Q|G-�P5yΊ{�ɕO�qL�?�r��2!%��_{�E����j����5��x��J�K��g4G�����*�L_�O�պ��=�Y�TyF�LC�Ћ&�s�bYYQէ�i��\�Æu�����y9%.�E����E�/�g�A_A�)8�6�/�� �����y�����#<C�yɞ#��ׇ�_��ː��`i(�N�~sr���"�z�q����-ʪgZ��yf8C�!6&w�����(�P�K3(mi�/tE�hraP2YȲ�;d~Qz��S��50��e����A��1'�HD@[Z�裉"�taK�-����N>.�$������gX�s+�/aϏByH;U��M����%[ 7
c[M���{.��Z���:�Uނg�{v��/�W#Q#R��PJ��n�=���`@<-|��u	�G6|�&q׵]~���Kq�<�H��6 �W ̫,_K[��U~�2ȚC������w	��(�����~���K�U7�͙*�?�H�y_��)P�@��1zR����@�rc�),����T�Oqү��"�����{�����y�E���������g|��
��1��H0!��qn�K�"8)�53L��$OY)bY�|h~��L�OG<D��|:����]e?;P��l��7��h��@��%�u₊Sk�]M薇�Ć�9���PkE>1ڼ�5e��P���Y/��j?<����?/��Y�2����	aayǊ*(�L��5Q�«�Z%I�����c�W�W�z#�T��c.��rD�(�6��ͧ��KB��RQGn�6v�Ŵ�+��c�5�Ď1��������G�FcL\���N�A�[t�n�q��c�v�X�� BCaJ��O "��c���{�sE�[�G���cј0�(㪭)�fU$��&��w���(�V�zq��g���l�0���ǝ���2� � S�9����˫C��id	 8Lg�����z�e���f*�Ǐ#g��Q��7��u���5�.��s��<n(S��/��
f�E� ��F��r�L��3A��%�|j��ڎr#_��ዂ���u�����[v+�<�}����A�r�L��監閻�e������"Ռ��,��O�x��0X�Cr(
����2�Pv�=L>�E� Ӂ^���y*8�#�G-�a �Z���3��:ni�cczSFP9i�����/<nL��cq8넅h�Cf;��H��[?�ِfV���d��3�<R/�L��6��kBO/ʤ��67��>ʩA��7b�������X�B�Ej�����2�Z���X��Bx��8�I-�ƻ��xp���vچ���C�&.��y@=�s�i�������ӫ���m��פ-}'�> 
ϩ2qϤR��je�u>���+���q@��0l@=�������On'�U٨i3	�/C�/�f[IS��}H����/�:���.;���>�o�DL�kaQ�$���~�:�*���QeJǮ{�nD(%�2C��G|6�C�\�|��H��0�����S�`�E‫����`m<���J��B;
V&ɟ7���w��y�&��4��!�ʅ���*ߕ�}4ﳳ<�U��+�O�5�3�.լ��V�TȒ�x^����jr�D- ��V��o{���8���P�[���s(�vo�ЉF�p�M.�|�A�$�1X�+�I/�� �~{��?��+���`�f�h|�z �O�Dx�Hm0�ڜo���!8�='S�o}�1�o^W$�9S��~Bix�M��u���mP�]��4�~��m 亀�@t&��ǟ}B�_#������.(�;�T;�=����HB��{�ڱl���h�R��0���c{iW�0[x��s�O�/�"U���#�>�K�kz�����Z��,RN�)��*u ��qR�wቍ!�:B���{m=$W�mץ����85��ϐq_L����Fr2�:�*�-ٮk����}:��r9g����Z�/z����Z��b��9XM�Ů���w�H�Eh��*kl뿈?*�d$(�}l��,q����[=7fVh�v���v�6bQC ���K��;i{��Q����̂W�=	�ȶFޫ.z�-�½$��/`�h,��{ 9&ฌp��8�T�NSVg�G%�ؿ�=	�X�����yQF�{�A ����_��.R)Q�B[���(��i 5��W���i��u�GB��;����ע�s�Y�g�Ѝ98޵sAs��K� �w��� i){34�.���.'[��I���5/��co�G�
�T����W�r�>渣s�;V 0
�+a[�ryQU�t���lU�kq��
�����Q���0#J�Q����,��{{��k�蜃&U3|�*1���t�{���!�;�
��3z�r�oo���ƥ�2��V���'�9�v>֝��J��&&��=�xE�cz����5����������K�]-�k�wؠ��b�'ۜ�uA���sl?�l|�H�����0��������r�f�|+v��xWY�X�]��$�?�Y���Nioۢ�f���H�~h5*� �=�]�Z��_R���������<��8.��j��'Pq*�v7su9_fQ͔�{}���X�R�
��j�b

�0���� ��sKZ��Y1��䯹��t�V�Iw��>]��|�D��%����Z<,��(��!��*r}�vzc9{8�]��D5���qi��Ck�� �K]�C��Q����A��z��Gx���!��͊�I�d�7r�w�2�1�*���+�ّn_R��m����Ԍ~��J/�������LӠ
���L)|�'g[�X�ހ%&H��H��>���,~�&���}u��г*�eo���wȩo�Ӧ�@�MkM���5��x�`rjX���`�����=3S��(2N^
}$&'X "9��γ%n�,*�^���iGC����+j�w��>���Mp�,�J�����X(�X�vܣO��
��E�M�/|���C����*jX��P�5@��|��� ��3o^>���=��ܣh�߫�][��� �#�p�pȽ��[�	'0��eؾ#\��{&��4r�.h��~�ٚ`U�1�Z*��,~h���ç��c1�$���	nՋD�LX�(Qm�� ����%[r>r�"VjM|�]���G��wwo}��p��=���
��
�3�.��%E�/j�����5h�����
���7�- �B�� �g����lr=�f�� v7��lΘ��%�N�̲�������K�|M���o}���U������ᘄ ����>ƏP[��؊!a܈�`��Փ<_�J<n�L�_帅���cl���Gͭ�5����[A"
o0��2dÔ���@�]���� ��NB�9����)!�{�/sq\�E���g^�ci���:xA�.:�b;�ͯ�]r�S-������?�2�s�J� 9�}�{g�|܌��#��I E�a�Ò��d,%n׮�[ǃw|�.�l�����&���[�G�7�I����cj�#o5�)�ߡ��*�37��s��q
VSvӠ���W�<5��("����f!���<���0o��f~�r�$��,&g��x)���O �?R��^����ʟ���
��4��Wg�'5oRj��!87`�w��#��y�������ѣ�u8׍���6��ؾ�rS<+��n+<�s+&���U6���-uH�YS�"\��&�j� s��Qe�g����Xw�!/>��(��E��Y>�ɻ�ё[�v�&�9p��`��*�a&���݀�隕Tm��%P��y9��<l�`(�e%<T� ���Lˠ��L �
�%"��0:��Q��JC\��J��s[���li�ލ�0csMI3�R�{Gb�I�>(#rk����.,ȍ_43�������x9,��������Y�m�re�=.��']��k��S ��a�r��67���9'��"�"�u%��iWz��z�Me�6^��O{nAfw������eP\�?��,�-"�?z��I��3c���K�Ďl��٣�q	�p��5)M���Ov���g��`������弲 F�B����l�,J�O�؛S�� s�,��\t �*�>�]��((!�m@ܱw}-��7��
����-�P@=��_Gھ�U�d��N��;���2GX�Ϋ����>-Y�n�h�9���VF:�'O�J�����b�le�oBbLg?������j���'^�������f�_��E�9�0n}�+��$��c��~����5q�z���������~�濄G,\��|���
u���n /�X�	Ꞷ�s	��v�������u���n�y�s��DO���I��a$X��M.��m>��*��N��q\YWZV��]d��B����'����$?�Y�u��E��@��Ž�}�|O_�\%q�6���D�5A0,^���Pd,�`m�wœ��y��K臭�S:}� �:�3-/�������IW���)�j>�Lr&ڶ����ΫN�_�R��bH�J�n������_~=Y�{����0	�#�N��r��X��U��{BL��	?��0@v�{N6o�%	O�[��S�O}�۰�?�u+��
 q~�YGa�Yf�9����iQv���:��E�h�[��x;����#=����L"��(�K�'����0������m���u]9���SGb
d$��C�f yz\ ��i��!����S����[��$#����]ⵐ.зn+y(����ڃc��ؔi6a 6*�=髩M��I,����!�h�!�-���'�K_���>�1|@X0��Ջ�Y<�PpjA՞EU�6���qv�r���#5�!���'ϋ����Z���/����"�:�X�6��Li��_�˕���⯟'ċt��S,���_j���C!�A��_�?�_�sZw�P(M�Ŧ\XS!�?{�J�o�9�Ch�Z�L�c�j��o謹��>L)=���}S�e�;	��*����_�@ʠ��b��2`�˄Q.���:� �-=�2�z�=Wt~"�� %|+�����ÁQO��i�:��6�7
>�}�%0��7��C�T1IW������a����J�C��0\��J��*ޖ˝����@ɲ��3����K��'��u�|�E	Bs��6*k��$��&]�![ߟ�dC��S�st��m\/)��݀�fr�80;;��C�ߘ��#�� ׈�律"�a�QJ�,�)� �㝧���x�3a��9.@����գk/bM�l��В�Df��ޱ��Z�V������QtR3(%�Uɉ�	��i]5���=��j�Gp�
�i��s`�]}oe����''�D~��������։9��0opd�0.9lp����d�����%{�+��$c�	��e+nr�P�h|�1���&jB�ܡ��#�b�U��+�ۤ���'��7h���O�4�h������� ���m�g���[� �ki=Wd�P�Q�DI�����"py�..�7�)/Ō�N�UN����R�e���%��8��B���.��3����9&�ߛ�K@}dY9�ȹ�pѥPh���d�7jUDnr9ylr�!�ûXm��͸3�-^���3�@X��4,A�$R\��2�nȾ6i��~�ѵ�{���@�������I�~[q��}R}�)r~-J�@[�v����o
;#)ǘ/^E~�Ma���mi9��O @հ
�j<ӏ��D3��.��D��*)Q�kj���	#��LտH�'�ï�	�on3���9||�<�'Q�-�=B�D]C]��ip}`�=��'�J3�&�5�����ޒ��78<��`���Y�}Z]<"�F�,~���n��_T)��V�;�05�e�(�m���7�g,�1�]e�r}el��F�\
�[c@�����5�r3������ x�s�/���ٔ�?X���)!?]�^i�m�X�����2�ʐ���QRY� 8�#i�R�?�f;J,W,O�7飠� %0���Y�{�)���<�M����e�.�!u���>�˧�S�i�w&֎M/���ۿʦ�Д�T%ܙ�8�V9jBU}�؇���"�Nb��ewT���-�G�b���M����&�LZF{B8�
�ۡ	��f�:T��ݦ)�-Ҙը�1���{'��mA�?��9d�k�v��
Ͻ
��u���8C����Zf(zG����Iy�cFF&�D�8�i��"��5���������o�ji� 	�]�]^�F�C��:��Ŵ��&���}��	<�N�	1~ה"A�
��(5�N��#��<4��F������@����D<V�S/j�T �~"�4��C^Rœđ�4ӝ��do2b��p,�YGL�O����l���Z���2�{Fg����S� ���ԟ���y�Q�}v-�g��k�fË�|�.F�>��.�.���l�)0�!v�b�Я��DGڳ,��K}ѣ�]��B���R�@�gMAeŢ����z^y��k�[/�6�Q��&EL0j�H;�V��n��]�)0g͕hO[j*ƾ����d6��'��|�T��Bk�W:��m�=�+�r�:~#�7h=��^cO��Ty�,/�t�&�DG��&S�&a	�[l�sK�LկyX��X � >{��%fbzaXC�/�6�3�@�Fy@
�͇�8ӭ��#�D8ӎ�����s-���d�p��̅�nDe#~o���<�M�<c���YG�&�LG.�*���=�r�ÊU�^���~�V͙��ב��G.Od��֙���u���$u��P����U��6�cT[!�5��*��BjAq6�[�c&���o1k�ܷ̳�ŪU���2f�{\p`x�" �ۇ��/�I�uN�:�-��,�R���}b̻e�s�K��emNK��^�\�8! ��j���G�5f�R4�����u9iS��G�R��|d�R;6���UOx�&t�~�G�Q�:��L��*S�vt6`�]KRDÓD@��4}KⳮĊ��E���_�@����@&1_fC�Y�6�N�e�U #���#�5�i�P����.�oX	���< �I�'��8b�6�p�_�ǌ(���0�x�����݆�7���V�"ޛ��"�q'Y?�dC)�j����1���<jc2���U4b�cx�r�^\՛�?���t�p:��y����n���,U�l�^C#���!e���^��6d��>�߫a�)�H�U��C!�w�F3��35=i'~���1��,�D�� g� =Q�� i�O��|ȔJ�S'�~Y&�Y"@�>;T�]�����E�BOU+bR��5S����q���O�	���т9I#4���:pw"Y�R/��Ї�~�,B���u���lmDO�ԅW����i�I�?s��O:�?��`��'�A��s�6��漬�$#.�0A��g�ڃ���`�\pJ�R�A35���u��v'!j��x�QXbhpr�%��8�RB3�Ė?mmθ��TB�ԅ����i���Ɛ��&)~��2�;��͋Mq�Z\�B�
Sߛ3Y�/69Q�FE�J����˰�Ρ��r2���d��Y�_3���G�Ah��%�L�_��`�;_&ֽL���h�(ɤ�o���&��c�ܑЕ��<���z}H�Y��0�=�ؖ���h�o�C)'=v�P� |����԰�X�0�� ɰ������cH,^�؉�PQ�v�.��y��Jo�8��4��(։&��ї�=\��ǟn�H�(�����_b��␀�Zcke�Mw_ s��:���Ia!��-��B\h�4'�^}N�}��x�.�����/L&"��+�Pg�ć��~���e���1 �XfG��9׸�7��G�~�)�;]�)I�Qp�w���"�o@F/6��	��P��]���D�b0#���������0%��"�|�La�	�M�e.toB�X�����S��>oy0�m��%��;(�"�Qw9�\Xۤ+/�����h�VH16W}��+̴OTD> {rR�ɞ��!R���"�Υڑ�t�1C�}�2�����ݷ�̔�Gf���� �7�A�sє�'@-�~9�ao�e.՟�f�[��u�F���]B�B���nur��#�A�c9��M����F���b�[��#�|I&s��A-���kq(�E�ѬTu�M�ѕF[�J�o#1�h��3���JI�I�g�U*j��;���&�4�?����m,1�!�������7�SyL?��(��To��: �]��>�<=��<4qX��u�5�2����R{j���:@�@��p����)�z�'3M0�
��wXl
/�����r_	�	!v���6�-��Dm>�|�m�H+�1�U��c�b�i6�~��`L���2����5^+(���b?��b�}�����zG��u(�or��m+xT��kFy܃Š���0M"���M��r"��*��]�2t�܊фay������b�q��+Y�[�����Pt
\�C��K��|��0L���_=��IBI�4��]��\����PL�Y�W{��y��1��C	�F�y�X�]Er�*1�Dy����Ȉ�I�>�Ш�M&~]�f�R���X��u^Y� �/��%��8�'���s,u������CO0�L���L/� �p}Q�IӇ�	��2GW9s��O( _��<�ʃ04���3B\�4f�#�;p�*�P�#e����z3��b%�7��NU[��K��c�!��cu��	��~mȽ�#Tz��~��5�i�Qц&���P������8�i&�5_��#z���h�7����D>�=va�)���d�N���7�_`�{��67,�|����f*�|l�ߔ��K�U��+u�2��s�:"�䰄�u
w�OB���D&񳤽� .}>S�w���ff動69��.���y2�xB�!��-7Ք��3��F��{�7@z�#Һ�}����um*�:��N��i ��H�iPh�:}#��t�!�94IC����/�]
�O�t럧�:����%<������1��i��5�̨�r�.����Z�݅�	���*Z�]N� �?���t(�2w����dme���MJ֜�!'S$�tU�_�'��ԆP���4��2lCDk��OX��V�<���L���A]�[� �� ��|��ބt�Ȃ��u^w��?YE?���E�%��Ƙ%+�Kp~���b��Y>`�X���S��� �Mj])�?|��dV�S�GbVu�%�v��ԏ9n�zA@<������I_s�P�OϲK7�^�(*�d�Ǉ�jгq��SVi���������������_�u��A.N菵�!�z}�c�c���6�r�GXm̯8&�|]��~���(��@p2�b�s%T7,���Q���Is���D2��Q����p]zئ�xLׅ�k��k?�����d�c��{_��Ѭ���C����&�T�eP�L�dUoMϼ�P����-�$R*�~�p%���c��� ���;�J�a��3���Sjs�ֶ>�vx�ͭ:��ⴼ���$Y��
��7Ǯ�����q'�+�,�^���]��a���d�c̖J�tCt*��0�Af�]�Q��U�K�Be� A�"3�Q���tð���k����!#�A	r�F��$��J�C(�}�}Ӧ!T�yM�S���'���~��e\��ܛ?Z+�;,��o'Rb�n�H�n~ڵ,h�&��G��8tЌ�Ly�����q�YX!�k�9�lϥ��ŘɪoZ�D�o�X�e;�q��rr@��[�BHD	���Y�������ƪ�qO����p+Fg���/-N�߿�f��Aj��r��S_�f^�D��a��F�;e�D�D��n�a`��E6��Wb`��yNDQ�1o0�ˮ��a�JE
#�)���U��s�ۻC��V����Ya�އ7�zL� �cN� ����U1��s�&X hL;���������-��3�v]�lb���,1��;��s�f�6�f���휀9���r���Ξ��Y��:�8����LO�5�I�W���F�jǈ����/K-�Q��!��Sn�zΥz�h���h���~�mB�R�J�M�^DǦ9�ѓC?��ݾ�d��>{j�aHm�����S BA8p������{k�o�hL��a��s����`�B@~��d"߫�D��BI��@����^.�0�?�
����W}[y��W��9�,xﴉ~��u����ֿ�����lǳfA��P�?��o3�W}e�&�;�?�JtU����840?��U���G�_'����D!O�ߑ�����F�k���#'h���{H�	�b�3��-����l��![Z����eW��_���ݝ'pݡAf��P�A����{�y~K�^~,�� ���n�Dx^���9���g5�?�%����w������y��=������W��I*,�^a�lf�H��<P�jӐwk��ϛ\qvmt8/��ղs��:�πvx̣��f�"8U�xE۲�4s0�n�s�]왎0�j�uW�]����k����:��U�@��Zӫ�3�x���!�߲(�<-Vk(�Չ�l�3����/H�K�u�vh?�<}����u��#�. ��*�,*	4b�?�����#9��[�4��5ް���h>WS��r��Cb��Lb�fHRG�w=	�秿~o����2@��Ҿ��yN[�/�-���ƅw�\b�eJ�I�<��ݰ��~�#Z��gl �X���pq���'�C���x7�JK	�Q��Z��av�L!�%�~�L����j�J��\v]n�Y&Y��MϲgFz�;��])W�`��eR�����f�4� w>��$}��6�����rv�����LA!}ƒ@2�7�2e����v�Ỳ��Pv*��<c��6 >tj����+2�ER �>_�=kd�މ�����{��X!v8j�P�Fj\����փ�E��І(�O������2{Ӝ���E�SPtv����a:S�Zk�l�ģX vK]A"Иe���q�fT�\�M�t���ȕa�)c�țm�y��u���Z���̜	�~E�ˈ=JJ�]m��q<j�y}c�$�������R��B��2m7�g����wM�'��$����;P5��L���J�~��V�ց~<��U��.�)/qjo�N^OF%$Ѷ䘬�Ͱ��:�d��|)�������O���Nu��fbH��kh���:0�Mg�
Ʀ���7�V�S���E#��ff�f�Q*ƒ R<�Ѷ��&M] ��rcf��e���HY��-�j����7���*[l��I�P
�8^5���6:��*GE�vؗ���0�a�֝,�L�R�����:@��S?|��6�	^�>c���ڌ|6ϞEg����5��(��I&!��FRq�YѾ�U�`&��M�U��y�+�ʼq�(Ih0h���u��>�;�_�D��-؊�֤�T��665����q{�Q.kb`�>�Da@o?-��OC'��φ�(��?/���I�(N�9�dF�5tU�{�c����������!��IV?^(�dCsb��|�U�,k��9s��"��,S	_�h�0moŧ�'�Ȣ���T�o�u�����G�u�b>���Y*fO�9�&Ǯ�`\$˷؊��{u�X��*����~R7���A�X�!ɯ�ә����bಥk�l�㢑!��Eb�}k�_��]�b�`?�}F/m2n^���<��6���h�m��D��2��O����d���'�|��l�a�ӏ���tk����%��?�#���L�jDALK���r5�u�<�p���-��� H|dwK��%�|O�T�NkT7K8�3	�,�
G�I����i	Y�k*����)�������H��/�����X����}���Td8%6򳍟e���kp��QT
j�h��}��| Ĵ�>]4l޳��μ>���D�X=�z\���C݅i)�?�
i|�Ԃ��g���]�P�0<���f�]3����͘��=1�r���UT\?��o2�92U��y�i�@lЎ������6�����H���;�()A��t�/�7ɣ_P_�c��ЍL>�AK�o�4�KON&���qe�;���(��-�V��#=�ޑb��w+�T@�����|ZNo�%�� 5�D��U00oSN�8�<��>b��=>�5ە�G� �e���U�s�{�}�]�"�cH�Tz9�"w��� ȑ^�̼⍞Bn�2��Wzw��[?�Y�̮�2?A`�:|���o���`�%
�r�x�BzdŔy���\_�����s��� 4D�2�Ĭ�r�4=v���,�} ��3��	!��B���%��-�&_;\�4
a�%��r0�	����+H��-�U��=+�`��&C�O4������Q���u)%���������G�LB.�����{�+�#�Qr<3����7��7#�eڷ��I�Qq7p)��+>/�s/3�Zl#Wz�ð�^ؽ���xD֘�]�Q��#!�G�^7L����:*�ds��<�.<_�Ϸ�_�9�Dӣ����j����=��=�o�^�<:��m�-gzO��/�
&y�����}$��>�j�4F��=
Ad�}� 5m���������-E���ЂF�Pdj%l�4�I�u�ux�����
��.4#Zi�wk�����7�'h�yu�MaY����uX�O�j'�,q�|��\���P����H+���]e�jL|�g��rx�6wE�7�Ow�_���n/��g�� �G�aЀ0ȧ4\�2K`�;�Ep�Á۹�� �4���!$����q�s�9�X��]:G��zXxE�f|)|��uq�&o���i���������[nx�~~ ���YV:buL��s�V^Q�At0�r2�7�8���!7"� ϲ�R�2�tN�����ɟ����l[��35NeA�xZ��4��Ĳ�Z�#n0F�����2�U�l&���.f����_!2RZj�@N�X���'(͏�&��8 ��2��&�`
ε
���8��(���N�	�[��gT� �lm�g9��<�����.`�����9�`W���������)��fON:��;$����8d^���?�؍%s��7)��j*"�I�s>�1��_�@����e>l�̂�Ƅh�
�5���w�g]h~�)����8��M�4'�@�
ʢi��s��xR�S_+�d�?cLf���VN��2�3�ߩ� �|gb�C3?��]�
�~{fA5�:R�J�A������E�M,9�#�N�oi������yUN*��7��.��>
����P�%t��k���LIT�"���Bw�i��sԾ[��8���vcCA��]ͲY�8��2ЈK�Z�Y���v������W	0�	�^�����E�ַ�$��8���&vx�k���9��ΫN�Y3����� ~��LJ�S��V N_f�!#2oq���6�K�����ս8�Y��m�(�)?	�7K�Oq�,Q��:!��ds�� }�\l���4��Jm)3�tni���?V��\Pѹ�Sn���+�p+��ew"K�0�)�ϻ�M�9�"��#@�i�3����d�	��Y�&_���:;���,���w���ec�KνLQ���>ã��s���d�w�6�7C>�9�hT�����s�u���Q�y��<n���$],Z���F.Ѱ)���-�a.M��&k���,t�&w����cAh��++�P2��z��g�i��uߓV��o�4�Q�-��`$�uo�����'����o{��$��S%�&�N�T�Q�^a��Y�L���s-`�J�~~�w��"!PX��6!^�tvW<+�	0�lv���R����?�^����+w�]وk����C[�����>E5���;��CSv~�C�M�.$j1��
[[X��ү0������	1F�Q���g�U��ВԽ�Xtom�E�����'��:���A�xE�V� �W��I��?�ęn
L� ��
]��Q-��]g�ԔC�ӌPxo䤈?!+�x�Ͳ{9�_��
�/��ϵ_%,+)�;t�!���ڍ�ш�q��T��(��w�q��6KD6��y-�rAT���O|]�ߥ?��}���ͧ��q�Զ���g������C'm�y�M���x�U;k������If)�l#��-R?ɴ�Wg�S�,'�(��Y�S3�?�j���m�� f�H$f�-7u���;������t!J '���xNr�U���k���f"y���H�j"FAZ�-�;�l��B�%��,���������Y�K��st@�u�E^� U��^��w)M���>����,W����unT�	F֓g<��NT���ѽRd�fkd+�;�;��(��j�]8�^�]�Ȝ�����Lj�6�b��G_dqT��3=����`穬�!0ZD�-�=X<-�]���'�֠Z�\s��;���]����KЇ�+gv�X����Yڡ�K�l��ϽƣR	h�X�hv���.�S)A�$���[�?fu��N��D&��O����(�KH��s5��"SH�Cf.�L"� (�����v�v�:E�7qc^k;���?1?�y��W�I���*����3eq��R��_D������� �J(.��	0p-�V�x��r^Z���
L�C��d�r�~/"�u(��\u!i�ty�4�2�^m�g,�V��c� -��S�A떱sGA��C��/m�m!�S�U<]A�v)��#�x*]�;�׆��<�RQ��xg
+�W,��(j�e�eaq�U����~A����o�ǻI�?(F���ƃ� ���#����&���2��?c��f@3d�>�ync�����HzY�gFQx�[6��K���.��}�u�#��1�'�G��YXbDG7]F�.��4Ճ�,{)��<��7�9� �~����M��bA��8�>jK4A�G'!T}�`o��E��G��Cl͟7Ц 	�,�5m�s�m��W/�c�@�R���+�c�Q��[����ou�t��x{�0��df�m�.�K���3�1C!�	��������F�1�+9�����Cn�8��W�î�L�|�v��#��<%ӛ�����	/@
z��p�vq&`駶g�^៽�o.�v,�PW�7F���x1׹�n����(v�hօ���|�����B��*���gk~19!�8:k�{)cˢ��AJ(�ͦ�|{�*j��)Im�ޱ�+?�8:�+�~�d�����t���1���Э�{+Z�6��t��~iC�q0���Tw�o�l4�+��V6�*�a�8!�pRq����V�b�S@c/�n��\jg�؜�0�kja��p��y��,�*�L0x'J^�
nt"�x~@E ��!HN���V�%���8"����2���⠿]Y2��rM���
M�ֆ�5�Tf�CW:���g-��2r�]���6�^#��蓎�Ŵ�ܪ���tҜ[g���A"��<  �eC
1k=	��u����xk���؈V %&nU�h��^���p�����_�M����y�A��G2����n�o��2��&�ed�+���T��[X5�s���.�A�0|����;s��9fђ�*@����C���`#Y��1����v�yj�j+�5O�S-GQ ��z���aD`������5�w�{��b�.�����Z�j��iXEx
H#b���N��SW������P��)��s��)�GL��-1,��lS$.�^���%G0�&�T��u�we 9�e��M�(\�\���ݏ_2�@�m��{�ȩp'~^�w�Kcֈ�,�1N�GN�|�j�O#ӷ�F������s���gZ�ҏ Td���n��E��lc E�@�ۇ�q`Bm�C<�e�{%G�T^L�lm$
�x�x�A�](��:F�	"�dڭ;���CцD4*��-o�k���X��ذb�R�)��fi���2"�Y�w�T-*����鴤k"�t`ʺ�vx�Rj�C*é'�ӅL���ׄ�v�0�z0�{�05]�����ќ�F\k9�� D(�� 9;ŊsL!ӑ3��.){�ٱ����`���km��������VDo��Zh��GEU�����:9�M^����Ec�d|���ɏK���z7	�ĳ�A���P�0y�d��"pC�П5'D5J���A�0C\h� ��f���;&������-� �ᷡ��ʥPpU��I$W�My��[h�yF��VA���`p�������~3�e��C ����A�CZM�� �O�����H���rp=,��ߺ��C�߅��3$�($�FD��KNP�Z��f'\�'.�6ԏ!�|��A$~D���a����z�2�k���Q{��f��i�z3����6�z�&�D��Ȯ�a�R,u��߲�>�|���Y�o��ٛ��	���z�M�-D�P�=�MZ��A.�� X33�)ԁ��΅.��^2���P�V�'VGE���eD{RB9l�1X�s蛓�+K��-=}65K����7e�����@P)����dy����c��@o�Z/�k׏���Tl�oKԞOa��_mS\�w�
y���]gQ6DA�]��p���ߘ�Cs��f�y1�j��T�2�뙔���C8^�`�& ����,li��5r�|�w��,-%8HĒ�׏�sx���v�L�M��*���-v��j�Y�=7�����}*S�u��� s��3u�N�L�W�u-|�^"�|�u��	6�u���4��b��mB��NǦ�)?���v�x�|q, iF_��J˖/�Y�1�l�B�ʷ���3�b]8��nf��n�A�t5��i�$�\�A���c[�ȏ�����cۯ��9�%j�'(��އ�{J8z���b$+�<hw��AX�d/R��+L�`|�/�#a����d�!i��Mj$�(K%�l[F�:z݅l_<����Z�wβ�]�ة~f���{�f��\=��܊����w�DD�p�G��TK6�èݠ\=�Ĝ�����M|�S�0 �p���J���R���@��v�3\�uT�ե/[E�x\�heǁ���@݌������ᡆ�g↤ 4hQ�3���F�*sqX8�0��UfV�ҷ_7�BŬF�2տa��Qq:<��:6�̍
�Q��!��pC���2�y)/AQl��Z����W�t����{9BJ�q|��A�N�P�<[��$hV[Bz���%t���ַs�1�"�cN��j��9K��������?Z���_5�.hwA8����r��/EO��lEG%Zu�t�~���8��
�{z�~�vWY�j�I�������w�<CXY%jۥƨͼR����)!������3P����w��Gf�m=儤S�b��̳�\�h���Ä�F�o�J��b�|G���>.�R��ׁ+��Q���*��PA����`x�$���9L!�
�d:� ���Sx�Ų�{р��%����7*l�;�����y�ѣ�.cz�:,�+c<������@;�c��L�4���=�!�7JS.�\0�d��;5���ͨ�����V/��HK93`ߺU���".sCpy�u�>�ֈ��8���j����Ԥ���n��t焪�̾�H�]ܢnj�que��S�&����/�G�kُ�m"�u�S<ԧ����r�o0�
3Ō�С+q����ٜ����vq�#]�|V�-=NW�s@�#�\�=�g��9���4p�V�i_*xi�A��byE������_ҁ��ǽ��F��[�	*�����F����.�j	��U���h~��hc���7��x���J�8M;�{���)	2W��{�o����MltO�{V@o��3��f�#YQE|j]-F��QZ��$�m3�j���ÿ�10C�6>@�q~X�z����{��V^bC;z���ZܐW~8	��sTJM�2���d�.�9<j�D":
�{�y����z�o|�9��S�Xز�Y���q���0!;��#���a] �)rM�gj��9!7�gAJ�oZ��ݧ�����R)Y�C!�f�M���+�/�(3a��P�⎉~N�_�����2� ���|!��}I]�n���}X�a�,`�kmM.��x�3��q�VE[Qk7]#���V��+1�A2�ԑv��	o�����&��Yv�����z� l�f�%�8Ŷ>�q�wfe+7��1Ǘ$��ߦ��7�U��;��X�{�b�#��l�T&S���{ �dh������,`O��v6���ms}��C�e)c����aE�:&�*i.]߷��W,��T�@x�^��L!j���ti�>��81>����]�1E'T����<$�Y?p�O
a��i�U_d[d�)��09$t&R۔#��Ha�M�w�O���u�,��Q�d�,����nA,q���H	��ޗw����z���L���N���C�S�>�5�U3��`M�m��cS�����m�}=Q��=ש(CĐ���2Ɩ������Ϲj�X��Զ޸�]^M��?�T0䑰�`�=@�m���ӎ�c��F6 �5rYo��a���Z�.���E���AX8�O+��Q���t�S*|���2��Y�&]�9�����ޞjA��]�}Π*|��c�k�l�*c�|�0]�,i;V�b@�\�ྫྷ,��1���#8-o��Qg=5��w���Anƻ��5(i�����ȯ d8�N_�y��	s�v	5e����,k�69Zm�0��t	9/�8�6ZypxRL�qXn��~C��Ys�=�$�~�mo��D�1�	�
A\Xqo��e�W���F������
�[~W�k;N��ӹ�����D�	,PK�H/`�z��Cc�^ 2$yƲA�u��na��>��)V��OW�����A��a{�9~ޘ�s;�Z�y&^z�NCi؛��C��q��3�e��ͨ�0T�f�#��S `�/:�~��P'
�:��ةho:��{�4��e�K˃�c����e�b*9���B���'M	��x�6	V���Wd?9g�`�4E��u׋����O�\�N�&/��\e	�����v�rf�3�C�J��۰�$�i8�EdW7�E���?����G�,1T2	��-L���Q���Il>�lm$���Ya�=���zo漖V����gLɶ�[qU&'��/5�� �!a�ըNz���������ѣ��{+R��~;>�s���W�ł�OO�"=���Z���]�%Qk�۾'D�؎D���z�s4:��&�;��_M���w�����R�̞�N�Nlo�z-����Ü�tbU* n�t���_�ty�j�����KS<�q<mgR�W"�]�\��A�KK$)�|T6�깽 �����"BE��?ڼ�K�Ey�Hl��O�g�]�P4���Eq�MV�����s���c�zK��l�q�,��xO���{�f:��N��#�J:���F����#4$#��5�
�]u��o���^�KbH�Jl��w؋nf��O�WUq	�2� ;�� ����⎛��ǻ���e��*����fk�W�0�	�(Z��C�ed��.e!�w����x��^mv4�ٍoﲨ�ߺ�����r�!�^K�JVjX�c���xZ�[׍�|�<4PG�z��o������_ǀ�d��8<�{&=��ZIN�ׇ�jdNtRR�㻬�җ�����k�	*:�Z����`���s�ʛ7����G���1x����1�I���r��/ΓҊ�f����Sn+>S~4�+g�H̬A��^���������;��/[���!L g��"�y�
��1��n�����fʉ� DQ�+T��W�_�`���n��
f��Bt	nR��l���z�9�x�٬�Q���ܯ�����
�J��"$��u߱#��Ԩ&T���ڵ �]�`�,T����aWE6~0�#�H�9t
�>��-bMM��}D4��"��5���'���_K1؇=���ؙ�]a��i�6\V�CF�[k�7_��s�ޫꞙ����KnT��-U񱝌#��J+���',�Y�&�]���@����lH{H���w�a̡�����>��)���=�Vrg��#]u�Z9���.-ف��8�F�UnXta�
��캐�`�1%��P��/{.��bpI�i�|��ע�����󍗰�|u�Y0 BNK�d���k�@rBOb3�����.]��~7l&":iq]���ut2�{��r�W�ms&�v�=��6��Y̔j�����[�����N�s��X�r�\p�"�yT��T��=C�>ԅ��k]��#��l_ʝd�k��Vr�zG�q)��C`ZJ�V&��N��p�mX����� ů���ER�RH�
z�7&=>�[��×��C�)˪<��\֛��U���f�"�O��k�i�u���;УJ��Х�B�3�ϵ���S%�"�Y�Z�T�2�˶��OF�L�&-PQ7�6�I����%!�

���>7�b̐dd�1ibB�G^aƿ/�"�n�B�������{G����B��\{�^#�uL]%!��ED�<�6e�k#��n��,)n����g�U��<��e�B������^^o!c�*S�C�G��ܦD����zπ^a����Y��%TE�$��wM�v���8��~،�rԗ�|?�`y��-4?R� ��I@�w�RT@:�Ø����aQTvB+�lG��}�w"Ǩ)��a�]�θL[!�q�a}f`�/�BIS;���QQ[����5v5�+G�o�x:�ʉ{҄x�W��^�P��������6s�qW^�{�np/9�x8���t�Iҁ���Y7���B������1�N��ݶ��mN�c�{��qy��ѭ QP��f.em�������y���֋���i,&��>'[�w�V;x
;U����WS`=��AoK�j�zpF����1Ż�O�MiӤ��� �	�J�GB�[��g�j��N
�`Q�KE�۫	�6��W#�R��GsL���P��p�~�|~y��="UJ�IV���
���?���b	 t��q���
	�iJ$'eXeZr����a�ޠq��E6ߌ�gds��߁?��f�������b���������)�;^�.�fu�	L�����}\�y~Y8����Ӕ�R:C�ؘ��t�X$0΢�/3�4��TB�F3��u��D��#�~,x"8����	N1|x�3F#�"ϯ"0�[����*��-�	!����f�K���n�%��"�/-��!�.*
:��p�Y�vS����aap�akP |<����r�����3�XqHq�N�`c��wZ1�_���V�z�vV�T�P�f�R�x���C�Y%�eX�2�?xV
����s9K<A��?@�\�9���w�]_$�d?2�۝���,J��jY&�SD�4%���(��B������N>KSϥm�Z·���ފ�{��|@"F���_������v{�V{s�tŦ-���/Gଖ��4	�K4�ʄ��9�W$+X��;�v3�>Q���ۘl�u[�8k��)'�H�MX�L%I�ӝCڛ�Q}��m*�!��dz`��	h3��B9#��ҧ{(�c`=�f�4������rzg��m�ڧ��A���l��:T�"7���v��8����8�u�ayu �[��k���:�>�/L⸭vW�f����~�p�T�A��9�l	��#�e�$�����]�&�J_/�yPT`�Q�g�O��.e�ߘ��%z��Q�ūV�	�������G�����m��	�P9�<R�eҩ���S>W��F/���s

z���L·�eJ��� �oHF�hZPłW]jW�}�T��g3�>L����ksx�}�s3]u�G��>���z;[���>R�(�����kVVU6��%�b�d�ȑ�7R����ӡք q\dG��$�T=t�I�����aN����r4m�+{���'���р���~�k�nݝ0_'�Mв6M�)-d�"ui�QJl ��BLfa������9����r�p����>���e�LK�y�:�y�V��JC�S�<�)X����!@/�|d����1������ ��Y�Z��iYw��(iU:'5���^Q뜟a +9�m�>Cwg���R��o��7�Յ�_E��c?�g��Lyj����8�B&"��r����.
����jK�K��z*�Pv�^��3�su�����Ɖ4��b�3�U�F�+�3J�@v!���/esBOگ����&^ņ ����U5_��[�ﮢ�Hk1i��iK�d�§��r�Q�s�8����	���A�.�Z����Q������ʙ�����l�c��P-Z+	ۈ�t�ba�%�/}2����r⸄�K���o��K
���ۅ�8!��g�e@�:�����i'����M��eݿ��6�����G�M
��M~���%��3&V��r�/z��m�����~�E��t����<���EY�1aI�U�F�d�`�{a�*�ON��y�GK�a3�٥�Rg�q���_���P��7���i�KޤO�6(}]]�*���btq= ��Pf�A�U[�wa/�8�Hp���7�)���s'�ޏ��]��ٱW�Uu��|��ּɧV39��W�v�Ok_���.���a���o��O��o�L�+����2��ij�ch�J��:��N�����-�ݜ��b�|�0/���yU�� 7bc}!1L�
��BA���3K
� \Lb� �A76����4<��%���lD��X��,��E�#�E��vnz�,1*��W�~�)�6ͻAV������ZKm���5��ԥi(�k?�W�l��6�։�_n��D�[-W�iwpUY�!Z*Zӥ2-�\�;�R�f��n!��j, E��uuF<�l.V����U�n��L*����QT����QE켐���^O��ћ��5׺͹m/�ԃ��"�L�8I�6a
����HdGt�/	Ź��8��:�T�_��|=�NG���⣪d�	U�Հ�~��� f���R�1X! �a�4͙x0�GGi���r�8�/��0�WM�k�YȮ�]6L/N�p���s�"=�	���Q\��fq�e[�<B�6�4�~(H�j��<��NV�lt��{af��
�Ѵi�Y�9WtH��-���<x���Զ���:|����;f���Yޣ0�)Ć!6����k@H��_4N�h�cy�C �1�rM�L�kr�m$铊yF^D��&L����<8���0Drq�|��@�IOB�9�� GIX��
L�|Mʋ�����%���*�EIG
�ԯ��q�2��w�`sn9j��r�����Wg:��`���D@GL���AVK&��Ũ�%�%��4<�c���-�g�w�
��zu�e:C�7ZL�T��w�͈��]^ՃGD(���|���=����&���_%_T(f���$�Su;p�Y�Yz.��Ejl�%躜g��vD���RL����	�uR��y�-;q��5f'�6u�Ĭ\ާ�
xh~p������ٝ�f�"�O��b��!�t/���E�t2�R�u'��p����`_���8J͠�8��Җ��w��k�w{r	s���C54R�b����h��͆�{�痗�W׽:�����#�!!��`Ӹ�x����vm�Y����ݴE
�_�������ϣ�'��\��{����bF-����oqQb;߃�`�"��n�d̃�N�a�D�m�Ѫ	-�e��P�s�ZZ>���a���j+�J	��FD�)���EN����2&?ҡB��~�#�����q0�^��4��è�R�+��<��h����5�M�u���/���E{$�=Ř������Ho����g'�]��OLUW��E�%�4�%��T�7�N�kt,%^���H��"dBʯ���w��oh�~Uu����(���(̮��]�ݟ�>��%��K[�Y2�	��zʘi'IC�Ot��x���!�-��T�:���q=��u��v�˕�>��vY;�~{�k�I�/�p(%,����xe5Q�G0�>>ۋ��A���_T�]�f.�2�!O5mZ�Յ��&A$,�D��[�L)N8+���b�ɽ@Ѳ��fd��d��o�S0o���ˡ�wTg�Ԉ���q�)h�T� � ^h� "�`[ A0>��V���]��Ouf�\�Ë�G4�_���ԭ̰��0���F�3�dt��8g�W#��O�̒�Q�tg�q,r��A�>�:��Y4�
>�J�	�Is-jR���V�����C���*��i��Xѽr�}6Ov�#�8N��r��?S�	=�E���].'��Y�qڽ��N<�v��Węz�(N�7�,��|�%��f�N�F%�$�~�K�����2��L���H�K�a(��`\���ʝ>;3w:8\[t���;Y�ӂ��hG�/�<�]�<���o�WX���&6=��u�B��Ƶ"���IU�LǑaBYh�øBJ���ઝpb�(��LIW��������;�hz��7W"�<��Q�?���
�^� Ӣ-do��=��-�~U�B�(=t٩�9�s�yf�r��]�㵒����I�����5c\PpD������X�Y|��/�N{}����%r�Hv�����u�n�T^]~ \���W�f|�߉ػ��ў޶Ny��I�08'�Lor5��/5Ä��͍��w�����H~��c_�D?�=_ݸ��7��u7=��y����,���D��٣�%�Qsl�KIY��P��(���y[�Jhz���1���OR�X�Q�h�+qs�����������w�P�Ο
���DR���&Ke�\���� y4�)��6��I�^)�ئ11��#%�,��K�\͵:R
Ҵ�,�bT�*�؜w�/���cNO��|/���F�>p�X�U-�4K���^O��0�hp���/V[���Y;����tR&��i��u���Fx#n�JʦD�X��A
��}#\� ^'���0=�`AM���ePpҜ7UT�������x�V`חG���m��G���c���F���:��_>��wBG$��,�{;�B���	�9���~���_ZXx��U5RB{zrc�����ZoL�'�x#.}�*]$G�I�ӂ�8���*օ�э�����֭[,����T��^X�b+&�Z�販t���L�ދ�y�������#��[�i=+�`���6��E\�)p�D�!��m�p�^ Vʘyk��'�z2Z�o�WXr�݇��@1_E9��%*ʈ����G,�Th�g����R�}��#���"ܐ����-���9�y��t]ex7v��1r�/�p/�"�X�j�[����6n�����ĭ�ƚ-�,t��t3�( �u<r���d�����B�CI���v���^D��9�c�07��E��&.��`��������S��W.���s��
�D�_r��@���Ƭ`�B4Ȯ�J�ޝ��E�F�܆��'Q@� �U����r���/1���Rmn"��6\:�f�w۟���^���>:VM��Lzd��h=���([N��H����ƭ4�ޱ��g��[�8��v��������i(;���yv;b^�\�e�}�$� L�~�y�x`��`�@��g/�ZM*�����:�[Êi.���u�[�
GAX�ǰ�ǹ��<����&z�a|��W��,O���v�"�r+lƬ�~��{NR@�»Y|�� i�5�n:v6!}�YV˺ğ�l�HT�ġYu�B9j���w~���ݶC�*2ڦ:e�67:����v��@���T�S���~�}^/[O���M�]<)q�os7��*,��d�����4��>m�]h�� +ki�69T9_Xc�>0�j�k6kI<��t��24pt�g�v:�c�nĺ�h��?w���n��ֆ�|������"��U�LD��Ӟ/=���y���cǣ�b�����;��\R��h�O�. �F!M/Ld�[�̰.�I��c��<�����H������-_e��VU�0u�f�m�$��z�F?v���3q���4.Ki3����lFO�����a��	7�v�e&̆s!-!�QKFv{����2oձ��Q��-%��i�=.$]�>D<���w���kT-�L��4'`���Ju�T$s>�L�!�k�)A��5أD��Ei�reҐ��:�=>��Gv�����E�j����;?��zA�i�@�V&9�"d��:��nxA��1e6��;� (K�s<K̇����I��ܕ����6P��� �20�i| ˠ�wȶ�S��w���i��ni�S*���	��f�;Gӹ�x�T���q�2;~I-����w%�34��z�[̌�ڭ�?����h~߱��'[Ԧ�yD��"d=ϓ.z��N%$�e@h�1��sP��]�;cv�m�X�~P�� �ī���RF�>�dϹ�/�"�~�?�!&�*�7d.7�G9)���R���_�9�d��u<�zJ���U��Q.<�%0� T�_��3PR�
H�̕�=��R��a�=g�G����$DZਚ�Z�3�*�����(� ����O0�"����2��x9B������x0D c�0D+�k	�6���'+�j����S��Ϊ���,F��܆x��[^������t���Y����t$�up�u,A��Ax�-.�Zd��!	�֘�<&kҞ�/TR�� �d��'�<�!B)l�C��b�$� k0l��#M��lu��j��]�l�8{|������e���&�-�kT咲{���{j1�t>�]a�W�@M:�7��%�jL�J&�-������OJ���e�U�drԛ%;�2��yZ��Ѻ(�Vxk�n+ݧ:B�i�3����p�7�<�G0��Rq��=J"w^����i�.��5$�(�w#ؚ8$T�1�I�ƅ�������/�+�I�~Τ�$e\~�V���s&��4��v�ЛsG�Z%�b�q�G�A{Gp���M$��v��%�xB6>�F��u�N)�U�=Y�����]��#�Uh���0fU=��;�[h�b*��ҿLR��'���� ��;1���c���r�A��$r\r�~So#4lC��ǺǷ/�_oTY�yJ�6XcQ�2���Ŧn�+1��� �P���݉ɮ�A226�t�c�i���y��yw�t�!���V��`�q��(M��$e�t/���Ӕ}؏Q�������=>Pi2D�e�G��I�R&�8>,�ݜ4�
������d'�8씚|����=2`X$�\�:J����Q;S,��0ڜ�5"1�E��BϠ!MF��)��`x���,a!cJ��IrZ�2��q��Ȱݡ�
w>�dw�0�:�}�>K�����Rn�̴ÍS�O��"c+*�IH�e ���kϸ��L��▶Q�n���L��F��������X�i�6�x�@�6)}ꆓ�m �0��H��h6U�e�@;_k�7\
�x�fL�GLڏ
��+�y�h����@B)(��������껭b5B�\~�j�R#DÀe9|UX��/٤�A&LI�w�3���b/b�,Ƒ:s���j����1�\׼�7�Ft�|���=s��tLr��1��������6z�((Q �H=m����R�x3�1�y�J��0� ����T��S}�EЕ$ȅ�6Ә�\#FU�.�>H[�N��=��8t?T�?|߉��`|%�"}�4[|���iI��J�5"}/�:G���|�@���\,,����ɴLJb��Ո-�ҭWh����ץ��j���0|�[�a�NTz��'E=6o%���hT�6�>���O�z���yܴu����0q�&��%����p1�@w|���C������=����ki{) K1o�u�}�jB��\Ƃ��1�_)�9��i�nn�9���
bj����Gqʁ�>�L
}#9=�}����S�{3�]ZL��mm�U���(Y	�2Hgފ��5BWr^#nw��Y���teK�Z�M��9��p)��a,�mϤ-���������&#�QG�I�j�(�Z�k�+OP�g�<��
m����J';��"����}Z,�x�N"���I���I�dD^0�^3���]<������s����-��ͧ�P��;v�'��&���?y\�G�9	��Ѱw�N5���X*8M��F�lQ�y�R�u�xR��-�^�M��k���aJ�<���&D���"ǔ9tg��i���|A4�X��)3���������NC�W(����M��޻���Zu�(�)�z�F]gP�g/4���RỤQA �85(���%�����Z����o�n8X>®J{>�-�v��Ve�飦sx�8�W� �c��A���z�B�����w��ꆐ(\��n{��ۜ
�y��	י'��aT�n�y?$���c���:����[#j��w܁WBD@������H��l�D 
n6�I�.�V��vL�����L��v�)Y0J��u�碫��h_�FS\��d��3��vs�i���5/��?K�H�J��]��:�W�M� ��cP����6-8�]��~�7�$_�N� F���u��U�GB�o� u ��6������j=����KL�9��"�+�6�G���:�,��	ro���s�[Z����@��\�6�k$Z���{T�mc�\$��x���@x	^GN���0�v2�j��$R9�5д��[���Ʋ� Ld�d���hS�U*+�׎M�T�'c�芵�Z�Ԫ��������1>V�n���3M��;���'X�/�'Yo����ЇS����JI?�bA�.p4C��j�O�@�� LF�	U̕�[P���K��H� �go�fJ�I���i0A�1����R���!	�sRu�c�b���;	��a���/��m|�y�q��r�-?!�jH�L9���.�3�H4�MO���ޚ��C�D
W��z��ɾ�B�(��}�K�~� ��`z�����)S1й�R�,.��6B[�g�L� ��*��"��{J�6j����b��c�*�{F���5�FD�$Ѕ�m3�X?����>W�㓏$Ȣ[ �!Q�T�I�a��??�N-��ic�s�z��wd}���RKv5#�Y��;��F�&L_�Z�*ei��lp�{��Co#��X<pu��۶w��Jꋊ�gU��E���V����8Di>4�F�.K�ɽ?
?�RÎh 6F���o���f�WG[���J�m/���[�5صۻDz������/������PL����H��k�I���F��-Q��fSK��k/�Ϯ�gɨ*7J��?о쥲F��K��i"r>�9fUG3��`�r�Ɣ��4���R��0уp��0=#`��#]p` _��
#���@��έY�gcx�,\�cۑ+c$� ���T����mK5��������;�-��&��3��_6��V}L�w�q����'��Kk���^ǈ)E�l4BA��&K�һ��-DX��v%I��mcy��u���_KYZ�Vud����Tb��m�pM%kJ�km7�{hwҿ4!�˷��k�fA��p#qh�Ӗ�+g�Hf�g%�}�f��r�H�6��9��i� ���I�+\��aq�f.�v?v֨A��@Z�}|}�߻�4z��ԏ�;�,P��ƞ#`a�ߴ`�ᵷ��{�Wߢή\�G�����b�9RKZ5�w1�ɤ���qZh�(�:��]�U(�.�@wE»i��� �2�K�����1�`��Y�	���>_"qAGvd/���7�e��U�7���=���g��,B��������wi�5������"�/����E%��dJ�#87&J�|�9;�j5�L��˰����l�1��+P�6}E�r:@pSk��Yx�K��,�&�+-��8������*Dgp6@�0Vs���]��.5,��4j��3l��K�^�rKC�_%�5&;�o�e]n�c"����p9���z�'#ښ(��&���`=�I�a����1��ф 3��%�N��#
���}M9���w�-9��.�� .`A�����U�_�N��!A�!��MI�Vǔ,�� !f9o�"�g��M>�����m�2��w�
#ѥ߹`��ZHm'nc2L��T5Ct�Hܠ��8$̣|+�o�'�J�s�@_l�}u��)E�	'P������+Q�&�Z[7$���sB6��ر	�p��X�����LD*��_��G�!$�(Y�wI�[zl��f�(�Dwv]6c�S�)���iu�lJ-Y�3���1ώ�o@�<	�D4��l&�Oou�N�����s�H|D����	�/�^ν�%A@�!J��F,��oJ<�*u�uQ&���֥0���w6pCY������{MCY��ӆ(Κ/e�r6��8	��G"<��i6 ������v�CHsϘ�/%@��Xy|�Z��!���I�NT�"f��5�p�mG΂�ŁU͓��u/�+�����j����RQ%�}B�0V)�g���F����Ȗ 5s3��8�����|��/ e����$O����2/w�!���m��x��|��]���z^��gm9050���ܷ=� ��q�3#�^����a�L�Yn�Bsً:��i�G�g�k+��~��d^�WH6�ҷ?��6���ǩ��k)��);�T���w�ft��P���C1��7�\��Y�����f^s�f�<W&K�l� �# ��Ҝ�:~ю��/����@�1:zLbR������6���CC��V����'���V"S�޵Y6 �7��p�a�iR�[�;�k7��C@~*K����sT	?]a��=&�!�p��!s�G����;��c�JL`BvأsBYȄ�a�´�9�ǁSp�E�����A��2s���s1*�/ԋ��wX����n����h4��<�����w銃��Z�:�*	�l���F���Ǵƭ���@2L��?8�>��$f�9��� `��5�ä�;����^����h��ʇn_+�W��3�&�&h��+���}T�̏�~�ah{j]�C��@��0����c�s�B�Q؁���i����F�m� P��qܫe�Q�T;��2QE�����"�u�;�Vfe룊�O[���	�n�wL�I��~��m����vd���HCR�l�LM	�sy����`KJ�����or[�u���,�� t�E���2�C%�J*r��Z!�w�i�PFV�?����+��Q�s�ELC|��yD����.�X/�ē� ��g�t������a��UX�����B�c��=�Zg�Q��\�52���eV�%l���	$��m����BC��y�U�HJ�����'�c�S�{�x�-�Rs���"�\N=}i1�P!Z��q����x�K����Hig�3!���h��e��b�vYr��u��$w{>z]Ø`{#�A�=}��Ī��7v�B����%>�ߚ�^�����D�W�1\���`fx�����?S�����p牴�0�=�ñ�wE�LK�$����e�]�۟1$,6ǏC���w��T��o�=�Q�<�$袬�
�$Q�MB:�Z̐x�pnxaK�\,똒<�����l���r]�aD����KN� ��x!�@s�u߳Q?r�����`m<&}L׋@U����Lyg�X���Rh���Am(�ひ/��Pğ�8�wX&���#���"��Q���8y�3p��a�bν�I�J�97��X"�PJ6�? ���ŭ4'�EZ��Q�
���˦m�2�*���D�Db��-��n�|6�������I�u� �<��Jɿ��0Ird�F�3��afI*3ivT �m��(O`��|��W烻,�8[,7��x�R~Ahx�K���F5��<К����Ԍv�x�x\>ѭ~qʃ����"�Ĝt���٦�Y��[��6v�ԗ�1sGv��d2W�1;�v�[�����X�v�oa�Q��~@�
ख़�'��`1�e٢�u$s^�У�8A@[�$��� PO���+Ƥ{?�BW��|���`/���w;�2GԜI�(J��U���lQ�Q��r \c�C�1�M%��=~��������Q�c��5�V�\"S�~�U����p����<9�f��j%�JvP/���9v�F�:��}pa�Af{�j?mUt�P�G�O괄X��^�P��v!7�I���r��ʼR0dH��䟦Gp�%�@ؚ��
���(��{;�����Gu�	�0yKp�П�T�M�eV���"����}����_���Z�v��Y��%�4��-ܒ�|w�2�1�a�3?ބ�W�"N�a����g�����/E��yB�����3��\R5�ʨ��9�H4�����ݱ9,���T���#=�Y���L���X�<հ$UH��(bۑ����֛�Lfʣ�����-�~�.��zP��/���/��	tG�zr�8'&k��_�#G��5���rN?p��?�ľ	J�ث����[���z3�K����C�����op?�:��e��u>�,o���IP&FL��G�?`���9Piz-ʘK@�l��B��w�֞j�	 ]�b��;�`}Ɖz�:�e�JƳ|@�<�V���7�8G�yL�+�Ӑþd+��4�9�@��Àw�3�T8�q�R`��"��2����/l����!w2�ߐ@YB�R6l�=�Ւ��#4���v�e��f��)�
��
o��v+�}�%���_�*��@��;��]�N�Q�6�e�%\Wӝ�w��B�'d��'H?��bB�8��>��fXc!�q����s��4��?s�x��u��?d.9xT�=K0g9:�Ζ�F�s͏���4�W�r�L�4��A|4���ȴ+mF�;���Fzڞ�z����H^�6�n	��ɩz����4��:����h�e|��
-�+����w:��w b^�Y�P�C�0M�Pb�+��e{��g\������o��nt+����ә�f��i�����0C�O�R�**���_�L�s�D���I�؏��~xo+�5i����||`JDU�0,q%�:�����ICً��qG�>���EQ�_:
e9�*��0dCv���<K1T��p19��)S���R}6��|\I�QGXP��W��Ok-mQ�)����8j�����u�L�W�D�Ӏ1T��{����^��,�??��M0�>u?��Xu8Kc���\ZAA�cP�����%��5�p:�V����X^j�G��IQ�4����g��3�W��G���YB4�ڻ�6��{�c�����?.�_��i�${�dB�[CH���S���w���]���۽ҥ5��넊�/�]�����>!�����16\���t&�%�)"�zsG�gIz�i��$�����`9����F�U�p���-�V��0�M��^��h�(��" %�R�܃UE_���d. ۘдO-���������:�N���t��K������!����	�*�S3�ܛ�)�]�d��m��׎�N$���?�J�OE�j@z:��Ѐ�2���,[�Y���-��U_xF]�y����&�� L=}sO�|_��L���O	�aM~D���e�)�T�z"W��qBk��Ϟ'@�k��p{=�y�X\�n�A����>Q�EP�(Q	�hޭm�9ў`�,�R��FAY�(�x������@��HD��D���C�x�^r"Wz��ʣW5y�L�zwe%��S� kAm|���1�5�w�Z4Y������acu�3�m�uixA;����w��A99IO�lRފ��n~��P��}\�n��oF,mv��7K�e�Ѳ[���Je6���73��9��)�� �=�M7��=@&&۟0�.��a.�Z&fW��3x��Y�rۛ�g^Kn"�m��y�WP�������r�²v)h�e�ژ���Un�������4$�b������%�����M�$@fT
Zq֔<�|w��V��'���՝��|l�d�F1�>�esί��e����]��#º��9ą�^paX�q������2_��B,YW���j��"#��Zb�,+L��_+�A|خ��~�)�C
���5v�b�ւ$�HO�	���]K�'�38]L�R8>e�)�V��ϨL���@h�7�ä,%#&?���٠�(��X=�0�/R����i�,�P�1�u�Ԗ69�Ӂ̉#��;���=vCk�bw�U�S#�*�
Re�-q�:Z�.����X�������\+z�ʴB?��U�7�g�惯*���;��a9��^|7ν���Sʃ~�<z�{dP<�74C,��d��by�͡���E�h5R�P����!�y"B�`��?X��>�H��U���'lZ/9裮��&r�'Κ����c`�f~�;F?*}� 3��̼ʽ��6�˩FO�w�15��/��;�$a�3\�K³zk?u��#�Xzh.E�	�U��.1�d��˭��6/Q�sA�/���9��ibvr]��V�OS xDd�a=�v�_Pj/ �S�'��:��w��(9
)��Ѫ���el�$C���=�S(�o��ҺT�d�|g�a ˥:����&a��I�p�D��v���d$������=�`�mjE�1����4����8BS���S���bO�X[R��R��yz{�/	U66�g���L���K����C�#:HVְ���r�X��"��_�?��.��ӗ:�ơ�� ���(f��!M}�Ŏ+��7��N��t�_�E!>qG�ż���n4��Dc���hnPy��i��I4y%�Sd�f�H8���q�ȅ�
�$cnZ��'�d�!�w��F�>���
Ai�2�K�-~�]�W�*�b��0��MEl�<yd߁td�G\�Q�/W�b�v�åUH�U�'����QsQ��uMw�d�='GN3�F�\`��Du/�(��S��U�h�W�i�Wl�Z�X��R�ݞ ��k��z/�]k���+z��#nF#=����ur�R�3��i��̲^���2ЦD If�G��ǌUB"{`�`Y�I��U/}�=Y�,8�Ž|�g6�c}ű~�H���T������ƫu������e,;�[8����#�7��~Z�ڳUց3��ǏI��E�LZ]�* �lH�6�Lo��K�bڋ%��,�.�]���*�Z�h�S�(�#��JG���E�j�5<! `�VO	��g_-����H6"Ç�������,����2�Es�)����^�TB$j<��
܀8���qhX�װ�Hĺcf�*vK�g�-6"�W(��]ʷB��"ޓ�Z��������R_�I���Ѫ����H�l���)8
ek11�O���&zt�����!S.J������v��ُEE���CCV�$ʩ��湲-4B�p�=�>�Σ�%�²�!�b�h̊P��\}&�Z�z�����W�F��I���a���gVT����n[�B�]�4��O�V�V��"p�{ƨ�������CN9M��
p�3i����_Tm��c5�Ɖ�3Y�H���s�ly�?�.��X��%�����փ�|l/�3@F�챮��"��?�`]y����,lM��I&??UIܚ�x�6�T��ǩW�+�FR��Qn�.9�#��#ʦ��\�t���!�|�OM�-���*R��H�V�Ѹ,n�-5u����g`��8�p3����>-uMb��ȷ{8��<h�!�!~��Q�V؂�-���V\�|姝�3�[j�B8=�Tdc�C\�dq��bK�mv�xz�S��N�c�3�w��M̯}^n�W�����A�)�w�z�m�6�.�Av���Z���l<�$� ���)�t�{]���J��d���mbl������r�P�n��7��~(���Ke�-PZ:��U�B|۟��ԋ�n3�,i�55�t������}s�Rv�d|y�ԝ`����ڴ�7���]�N��TC��VN�k!{���6C�Gn�:po}<� �C������%��� D�Rߣ]��)yD�:?�6�~�d.>�ny03�;M]]�ҥ��ǩ�֤F��d6C\{�Z"�
8�����d?yꔩ�I���|,F�I �->|3Ld^��fɼ�����u9JzP��ƀ�M��R˹�i����6�p�8��t���/�-��^&�:?4.�]�h!W��i;&4�(���$q=��IC�����W�SՌ��EI�7�/�	�w+��&�o�[L���y]	g���Z�4/I{�s��I
/mׄ��H�J� ]�x��-����m3-�?,>������w�4��@�KZ3��Pۺ����ex!<���K��:��S`Aq���,�k���VZXX#C�;����KA�:-@�nR04�^����J�l�h���;qƳ�����E b���s�_X-�!��ߎq^/V���*tB�8�z�:I]�x[l�R����<��Gh��XMC�Q_k��oO���_����ۧ�g�'�|}Lc T�f��jfz̘L(a��p����~����gf�A�gL��d�!$����;&dA�y�"J_ `�|m7�r�����p�&m�U<���m�/i�܉���o	۸f?}��S�e��ч1Sr\K�bt��2D��y�L(v���I�{��5Q���N_L��"�$}x�r��G��6;���̎��)�	m���^���wԘ����C�n&1|\:�"�eJ�cԀh�T�|w��hs+�F���6-wN{�^��ꎡԖ9霋p��0.���Pf��8sN�Ƿ&N��Q��?ŐM�����o�R/��S�Y���2�c�6�=�*l�LcE�����V�g��|V��A��.`m��8�[I��>+h��S{oW����;�L�[�i�̄������W����|��(�xV�_~��a���2-�h��h�� x���+��%�ʓUh<V�(G��{iy��W|#ʖ���O�t(�ێz�_ș�S�U�t��6[�>�Ɂ�l�uH93~ �>l���)a�����+8\� �@�{��3#r�O{I�8�!�-H���k_�����8�,(��B�{��!��ŮN�ɳ@+ٳ�F�����GF�������I\o�ms���t��?�I�\��~��@t�N�Tр$X��P��A�kE��1� �\w�}q���L����WW��'n�$U�_��Y%���N�bf�2��U�#O ��χL�R)LS��)|$�^�H$�A"y}Q;�zG#K�a��V:w�C�Hov�f��3w�,�*ʐ�����YJ�2@������K��Wb�׌2sΑX�糟ɘ��W�#��;R_c);=�����4�4�$F�WYڱ��3����.�9Ie�ӺW(�1�-A���y*�& B\�6���x�_$Gnt.E'��K#2�z���︱�m\FO����--&2z�O1h��;)Bh��7�se-��0<�^X��_f_,��i��(���	 S\\͂X4V^�|B�G^���GIs������M��K��Ox�X�)�� 	��׋K[Y� U�Ha�Ze�*�F6g�\�NX5ϩ���Fev,�O���0O����� m��m���T��ۖ	,���N#D�lL�+�x�G�q0�SYot1��^��k#B�A�i���n^���=2����ߎ���R�Jf��g-Z�eR�D���)��ɟ_]��E�L6K0��k����PoI 6D��9!��.wIGTw��-�-|��\��8N,Z��"g�:�=}W��S�]X����u��Q��:&R�(] PA��[cTܟר�<[ޅ~��b�}�|!{(�<`�po��R��g�M&�,2�Ãd�N�7��ubI�[pX��d�k�u������.ͳó*�X����j�NF,E�F�پ�Џt��Q�^��X����'^A������Njd�:j)���@	�O�*�.
gb؆��F���n�<y����������3Lx�m��m�<�0Yëɦ[�<�l�۫�p�ܲg���`˞����Xc�^x솖��xg�:髃B^	/Ax��/B�6,�qkN;�c^'�o����Cf�~�O:e�@�i�P���ɂ>����94L&E�!tA�{8!m����/ z*�j���e,&F�w�R#��(�h��c�Bݷ��L_�e3�lbI`Bwn���)�{3\Tmq�J�����[���Ǽy�uN�5�D*�圭`��Y���a~��x"ۜm�{��
�*yiW�u"�s�W	�	nj�d=� �Zk����1�ݠ��v,X��$:1���%��N�}��	C/�L$�Ǳ0�7������}j�E��J�̇pЍ�6�w锘9U)�ߖLlߙ��u�o�'n'� �h�|U�mԳ<�&�p��m��*�{B�݁���"?\n�a�J�s׾���x"J��9����0Ř��J萘�L����t(�'���E ���4�7�ɡl�X�F�#���K����w�����s���p���5��]�&�Ho�s"j�
�l
V�m�6y�?�$��S,;ϼ)���8���b-ʠ�kt��=�=�̷�����;(A޳7JMM%ٟ��8��'�_ȍ.�J/t6H�yɦ�3ƛ�麛-���;�P��:�}�6�9��s�q�˹6�yL�������vETbݱ�
P�f���xRBa��DS�)��^g��׻Cŉ�C�M"e�W�k�4�J�u�u�����F���wY�_��!v~�8����/��|%wH��C���)bA��ܚ6��S%$ݒ�����ډ�δ��3n9�C����/ Cg��BU7�,�$�-!I�e�1ӁJb�������)���OH����D�F�������;���0&\�1����C�M�ۤ�m��+}���׺��I9%[1{���Y��_���t�?0�+���"'�5��Ր�қ�}� P�����)�f�<:�k
��H�Z(<x_�
�'jV
�JV �N&u8�nNK�%��YM���t�;�'+�q�h2u�ƺ���~e`f��U֔����x�}$]��j	�du���߼���$B@,����EHvi5�ꬽ�S�;{yv��b�Y%,�s��4AB{���*�3Yu�+�j�I�LH�u>]���f&�]jW�	?����U�:},��0�_!^ɪW�.�]�!�F�yK��Qî�OSO��l(��%�Ս�~z�ޥ�w$�PRb������:{re��-vI���f�&Nu7ׄ�l>�Xjf�Őp�W�QϷm�w�N/���硵���ҙ*��D%V��9��{x���A��!2����Ha��]_�@m6Z�/���'t#G�-Q)OC�"��BLQS�{��C��3�C�1�Li�a��h$x>�9 �G�VF֭?����*K���]�gUٶOЉ��K�~�%��R�d��Y���t��%)���lk��&>1A�~Α*��T�<*��y팈�]�#ȫ�,%Q�fX]nD4 
�ɳ�.�HG��l7:�GmмRg܊���]);X��ZT>F�G�%P;�1h�{�H�M?[,5kڔ�t-	��m��?��ڧILje�i�{�*-3^�C�q �l9�E�w�)U9:XA�f/�����-���7Ɣ��=e��"K��+�[�wÜ�K�n�*`��C��$^��K�q���HM�vJ��:�Ʊڸp^��eqRuU\2�6F����C��!����'��F���AM׸nI��,�Y������m���n�l�S�SJ��I�Ġ��k��t12�WO�c�ذ~���:~ս1�z��8��+�KH�=��9y���2�߰��d����}����M+7���F>��I��<��/��ZFu����S
/j���^.����.�b�SJ� ��?a w��pD'M��ݎ�L�lE�����귱7�F�
�r5�{�lR�5S�0����/NmX���D�$K�*:����DY����D�>��%��w�
���]�����Y��͌���l��w�:��>*S2�۱����z~7iF=A!�1U�΃E]��@���9�y�mwU"�QP���g��|��a8�=�=~w-���[-]��qu����Ä�����/C��g�f�]Db{��O���h�IDqV%mP[ȭ�D1*Q�ص,=����ȯ��.���/�Q�X�-�V�-�v eC�W�W���c�u,)��E����ek��A� om�u���I���О�6�L^r�NIO~��{�Ym�.i ׺>B�7c{��Fl�ӎ'|`h/���K�Y`���d�3�����=o9�r������HE
XvFX���z �\	l��������3$ J{�wn?���V�Zn삾�$�{�0�An�ƪ��i�0뱪�_�<L���RO>A�����2�-j��N7;��!X͇�}0��@����c�瀘�<���`BnKZ܅��� i!�)I6�����'��vȭ�lb��qj��s�3���֭���6��َ
M1��}�����b~÷5�v�[��H� ǀD���K�4!
��98o�:RυOӻ���&Ɩ�ttk,A%������lM�rN[+ �ϟ^+�+�X.���K�� �`z�y��Q�x&��j5��a,�� �G��-�I%�F�U�U�L\F��`DjQv����Ttw���@�S#��{��d���[(T�]��	����� ������8� fO��`-�ң�K�+�^+$vq2 ���>��Sz�w0;\z]��o�2��7��:�a�S�VoYS�G��,(zV
��F��~��U����޿� �3�:Ű�����K`4�QM@�$�E�򲅠��\�(�/�Y!A�ݱ�9�eYLe�
,�\0��l�iX&�>��Q���i���rU_��I�4���T��ۼ��@q(�UZx�)�kT��5���+L�]=^��7o�L�r��˓(��H�� �0K}�C�1Wݔ�O�IB���e�T�5x��y����)Lu1#S�ø�n�	��>h�;��:C����|Y���;����{+�<�� x��#7ۘ�Ug�*
���H⍀�̯�GV�����%�Y��ũ1,����b8S2�l��E�������X�6�UgϠ¨�m4:%b�&�2G_���՟��홌{j��_���'�J6��f~�7�mo�l�Ct�`ۥ���iS�/"19�*x_�|��7̌/k0jtjB}Kj�cju���tf��@h��� �����b�דJ[l��!_bD)|I4PQ�5�"�������b�ߖ�����W#�C�AK�~*�U�=�/K�Kj*s�̈́~?<�a��c;�~���-J�P��٪�Qt!F�x�X���TVh���؁ƹ�j]m�������k�r���WȒqIc�U�]��$�G�t�9Y�<�߉�0vn`H���M����Q�;y�3����kk4P�
�$�r1K^vfbr�Ս�S��a�?$$BP�Z)����a�͕������]�<C�N&0�x�<x+��������j�@F��*����qi�CK��t-g��c��h�<���FE@�.�0�E3�sl
�U@-���p\�SK"Kի��,=�_Z�2O�	9�=���D �BW^�V4
�bu�[	���FKH2+��Hk|�>U�0��z9/����^v�\K��?)�p�,��ǭ�$�(����'�%Ms�9@5
쿿8%csT�\�þ0��[k������4�u��q^�k�>�+k�-勬������C�il��m�_�p������`�[D`�j)��;�yֶd3��#>b��i_3"��Od�����p$���a��\:M�$:3#[&N��+R���槰,��9>��J���'�2����Si$�>p�l�mMw9Ȯ�)�l#�׸ ͨ'�DՔ^��B��cTF&c?MA����ɻ��ҝV!��DNÉx�^�CO ��Ѣ,��_>o�i�nk�=����n�B��0��]!�n7��<G��ۀ�QgY��}�ԞXgo����?~h�^W돫���^�A|iB=;��g��n
+Y7�bOE~}��3� ��!+3}*��`��$7������w�]��Ə�i�ԭ	�CY[f�e�.�e���2
����+�6v��}#.C,���f��0qp%j�&�y�Q�-�6K��R�|���:��dI�EnP� ;`L<���P�+6\ݮ]!yW˓Fd��D���|��0:�-k�	L���c��o�-�4���W<�/)M��ɥC(��t�g	N�8'����ܒ������Y|�&�X�lg�i5Q��S�{D�[��3Ͷ��l:�ұͺx&(�o���6D�ڠn:���*[�
���B��q>
�iȏ���}q�kH2R���N�3
�$Av��t���nP^~ ��'f	��ә;'(��|)"�k�g+�2��(����FrO_��k�2y����~�琢eEzQI���k=�h����^%")N/CUݜ��2��Gh7�Ң���L̦#����o&0��[�t�3�V�ׇr���E�h�B�<���'R�(��I}�M���rQE0�ĝ�j����F��(���/���3�x��L���=M�����ʼ�E�L�=g��D�9Nx�����nS�A��
�؊ې�V
�N��)��鿕h��Y��|�?8?*]M�Kc̷�-!!�<�>�#�#�lnug�	��C�[=��A��	Xb{�H5L�p#��	w̩?�9?mGk>��6����Dz7@Tg^~9�l�
� �U
��I�K�����3�4���d�}�ܦ^�
��Q���1������Y��O��^R�"��ޢWӦ_��[��~�)���J�}�D�o���;�M3������}?��l����oB�^�=�fi��3�zp�}����49�r\u_������$'��qxs�\�]	zs�1)��ǉǚ��8 �2��-0��WX������^����W�o�	;���xZ�j��	�d���V&��-�!j��.�x�
*�"Rd���V�q���?
��9(��ff� �2Ę��a�v�q���+j	�[;���(�V|�������ꤸ�UY���y+�
G��-����J�c�M�=g�"jҺ6���duLj�H����i�:��6׼�z��h�=�ϝ�1�iB�`�f�Pw�#����m���6�-HЧ�5����]�S'˽7��(��9
[W����*�Z�343I�G0�ج�;������d���-o������f�qm�\Kb����s�[d��*bs�-� �J��@#|�|��xhV���&�@U��X�4<�|�rr�R��ϟeQ=���HK����!�ywL5z�P?!�l�0�����l��[���:Ӌcv�����Hv�|��)b�*Z��%pTI��HA{��H#%��#�����/�����k����c[�1�4��4�}���Ϲ�Ð�-\�8��+<���O��`,���a]	K	���D�����:^mqo���E�m�n�a�M�����������������x����LvC��N���S|#�P����,c�{�o��v�6t�����[mI�j�;H�錀-Ʋև��ɴs�+�QwX�� |M�w?����K�eǶ�۵��M��c!�(Y�^@�WcYr�#�8���o(�G�Ny`Mյ���Ck6�L�N�z��J�Fpx8��(A�����<���qg�� M[ȑ�������e������B	�A3�����D)x>b�
��+w�7W$�WЉM� �En[���S��4n��T+#�W������8aĤ�Rk��,U}��x#xC���� �z�¢ԫ�!+��<Uw��}��L5�;���ZbL���p0��'M�=�"q���ř�4}c`�����K�C�F�R��΁d���p9o���C�=H�[���d��������x�fS���+_k����>v��쨃�2&3.:�1�@>^�����Cܨ���6����`}�?��-4zϜ��A�k�P��i��r�,�C���RҸ���jϟM��修���F�I�_������2('(l�I$��ڦv�Ƽ�s����_�}:uGo1�e�wsq��zD��h�*Vҍ1��R�\e7�6�K������!p��9i[]�D��,�g:���}�H?����~^O*[Z�h�M����V��$ޢ��M�/��!䛒P�>c��0%�y9��@�2�kʉy����E� ���0��[\��=<J`af���j�F��)M��Z�W��9����^����H��sF�	�LCEOJ<2��ܱ ��zTn^�O:�NA[ڿy��9R?�u�����̃��ƕw�P�@	o�of�)� �&��pCh@���y b��n��X[���g�oi`��Fl�:1j.���|6���615?&r�$C�`�J�lt l�`u�'=��)_��8�B�<���	^�g���|SSCc�o8F��KH�F�Vo9o����h'ݚ�|�T�h�N%Jϥ��<r�iAo]�$�=���wdYk��\�]2U��FE1�% H�M^�E�,��T3ħӝ�����z�
eM7#ivt�G:��#��'��8.�rb�"60kG��{�L��N)��vg���h%]��	��L��V���$e�21���^GW21��C8�*71�5H{y��t#��'�:�-ٺ���Z9�O=�Z]�)X �X%��sgK�wi��4g��	j.�c"%�i�{b�=wm{z��"!)�ry�#�����Cfd�N~� �hV��"o k�����A��
�w2UZN�6,9��n�c�v�NM���j^�P,�R���t��M
��J0���ܹ{4ƈ�/�5���^��7�l�W��k���-[�{�Y�ی*��L�}�lUሤ%	
,&������,��u)x�rB;��	�;�vn�
���,�I��Y�%�Ze���y��B�:BrKD�X��"6� #qٲ�P����a���DFN�f|�c�R��<*� ��m7�t�a���īTD����Wfl��H9�"�ٷY��
nȦDi��t�=;��~W�|/�ew��K��t��*B��ʝW���� ˕M10�<+�)n�e	�zu��1����C��~S?�R�ݻ� dT��Ͼ��ww��_Ū�4:��(�'�/�����J{�}N�?�)�A}SƳDtq0�f�i����^<�聞#�l�<F$���;�A����:�0�لl�\��	L��1�z����YY�|�q�#�E���f{��^�"��o
��wn6n3��ԛ�UH#�mdY�[��ON����*v�?{���	�� �^��M�G7l+C���nRX(�'$���P�ɡ�_F�q�[��Qy1��)�6T�b��>��h��4K�\�jvd�>�������B��Fu(x7�`���[��RL�5����h�D��sy�OڎBAkm� �*���I���h8�*��R�b�y��d�f8Hdk���w�Գ�����Z�:d{Evhї�b�����茆���/��q�Tߒp���6W���{,eJ���`Q�S���g�f�㥷RW
�6��������-����
*�Y<CU�h=&u�;���j��/wC+�'Ɖ����"q[d`p��}���~�XF���3dӽ� ��V�A�{��M�-u�Q�},TT�Y�jj.F%�^��nz�=���������]�Ib�S��U�)�?E~z��F��~CEg��z�Ʒ�w�0ɺ���h�@L�FV����s l3� \��I}8EuX�r�\h>���J��P� '��C3�tK���Uj������4
ʋ�x����U��4�u��-�h~��0�u-�p��'��7��x���S=.%�4�o���5>f���-��p֒�D���`^�Z#H��0���1*E 2���J?v� OՒ�װj��?0[��cM_�<�Lɛ�b�qU!��Z5T):�x`�ow~w����,H��"���ƳM��C2�+�j�Ѣ'�O]Y�����?K���+.�q�m��&���������S�P7]IU����b0���O��}�H����enhZ��)oP�{2�$!7L̉�R �|R�ݚ���M8��w;e��Z��#�dS���]0�ϵ��_��>pg�LU��"Ro�]{s��nxn|1�<%J�ҟ.����*!�1u	��I��*�m,���E��9��=��S�w���N�;����z����t{V�!�������-(ﻍ9h �Aވ.�J��LS�����B,P�Rg|�$�|�6�����X'�8�]�9������g��<���H>V5�rWߟ�__pc�DR�"�4���-���Ds!��"������8��%��j�^:�8��fAன-����繑f���a��䁛��Έ�ȫ���Gf��>�~]�h���f��H�o0|O�٠���na�T�N���Wj�5H��A;��eμ��f��K�O6NĘܱ����ZB�ܷ^�;B,��rv#N���~���I ڻ�ղ(�Z�/a]8,Pv,#�����-��?��j*}Ue;�z�ȯ���e��5�r��%�^UK�2H��a��t*�{J�����K�s;�̳%�K&���g���[�ܬ\y-@�L���=�ɢ�������u��֗Ч�$y�x����[�}� 	����֓Q�/b<엗�J��	J��.��=���}>T�HL���*m�8n�V�JӐƝ.���k^T9� 1ř��$�)�n.��Տ:Y<ߖ�jL�ΑgZ�+��z/{e�a�w��{p#7�<���p���'�X��!�M$$P�}�� ��#��(�
��D[��I����(M���}�_y�(ef��(�H��v\^�!��^�2��Y�l�|&��Ы����_+��5�ߢ�A��S�~"L������ʲ~�@G0s������)�����`�Ж��<h�-�H��ǞЁ���ǘ�>�����[�"�(y;ۢUE���V+���^4MW�q!&_�sA�{m�Ȥ����͂��+��Ԫ�Y2k�+�.s�4��LY:`6gvp�����2�x�f�-�C�V�WWTt�+%�:���ew��	���Q��T�{e���[��YD?���I�R�;��;u�4a狒�'pr�'����C��R�#|���F���8�� ��9�j�֏��r?6I"� ���,.�]՜��H)&vDYXe���fL��
�5�S �v�>��C55��7B��V<�8��_��h[�Gn>�e;�C�����<�F��A���ui���;M�Y��3��+��s�>��
 �p�W���?����˓��$���ŉ�k�6�$6>�PLql���+�yø�E���l'5p�嶮R���3DE�g��˨Q��0Zt�s3U5N�b:�'���-�	����1cb_M��E�;�g'F�s�}�O��~���|��0nْo�>��!��dcH�a���������$�(V�o� l��9����\|`������U�a����؀"s�#��-�/����Fo���}�[�ō��J��=-`�a���~7��+Q?
�>n�69[n��B��}p'y&-Cn	���9����Z�|Z��z�Fx�_G�����B����jN�b/a�md�)&AMT�ܝ�/f�b�y�,�y?DW��g���oYz1;>h��O���/Qє|�N}[����m2�U��k�,Tj9�~DV��XV�[2�m){�z@Q�{π c�}��kW&�yU�X�Ok��J|p�̽y�F	�p�Zcc0.�G�e��w+�7<���| <b ��"��}G+.�듘i[��h���?��z�+'E�:,+��w���$qp������rY��!�Cm+�<3��_+�Ĵ�˭O�� �2��c��[B{Փ̐�FpvTM��>�o��YqwrZ���&|=��C�P�2�1����C�e�C���py�p\�g����~�lu�#p�f�����щ�6�{������9BM���g�q�(���d��+5
k�-L��Saj �f�Bz�@�Mpf6��1���N������n}ժ�$���Gj��s�	��xL�֊bd�ԉ�����а�az=�tXٛ��x��)���h���,v)8��4���4k�Gy�R�^1�}���7�c�W���k��(�Wσ��qh�VPx�E]�qNc��2�&n���. ���;���ͬXT���T��#vg���$�� �E�P\��tQP�1eO� <N$3�*-����y�c����r��4��?��Hm�̀���5�bA��6H�1Ս�:L���A���~���p�Sn��cq|]����7y����\���P;M���-ǯ�zB�s�ƉxM��T�QW��tM?�A�p��DYz�ի;o���y�׷��f)t5e�1r��/V gؚ��ؚ��lz�D8k-C	���	≉��RxK;� u�|�P8��u4:�h�<h���9Ȭ��6�7D�sq��ܡ�������kѠ e��fC�z�B�J�\w�����C/��*�4��J����k��P��b�bh��E����M_m��� ܲ�����^H�\�$c�]�~B5��+��"���}��x�H�������PŪ3α�֬��0�!pj��q�����1�'՛N�d�[���R�"܆��*��~�%ܯ�q������?�E��:�n�N	{2{呆m�Ś\���2u�Э>������]��I�;Zgi�dA�I�$���w�,�`njҖ�R�<�6��F�'4�L完��%
�_@���+[������=ph)DsR�,7c�V�A̓�{9~�=��޺�b=��%�ɟ`�������f4��&x@