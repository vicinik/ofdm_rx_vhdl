-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dfRR6Y9k3Z49nbM/e+KzlrdsS6YB/ax5wTsNau8/jO0cIYj0MJKcMXuIXAPkThnH+sbU4jBuRdjq
HijUCZ7rwfSfu5PKQI3syDhHgiTuzvt61R8r6OIC054PZJWxPJ8XYX0RPZ33VrxqRDZB7J3kvBZJ
LQfmNeONbhYKSmjdy+99+or0wqNq3jGjXIxdf/aUKBq2S0vy5d8swynpLgrOrt3/F3KBi2COhGyf
PjI+OYBJw3aKM4Bt99/S9tOHsCoT8+JgNF6DwQxrGdlgyHoe350U19Vr79q8EfQRLdYTMZrPGN6q
3aLD9sUtYfSlolMG+qjljcbLyVl1GHTZJNsUqg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9600)
`protect data_block
UqvhgE3s9A17bbJtx2SXfBX5m6hO/go4pIJShHqwOm1Mxng7glpnrni6BPqnEc57Cw6EK5TKej7D
w6ueXLY66YgnnaxRNl7RLKDlSk50n55HGJCuwua+/s+KU4MwEH3lOVhDcYeMyp1zXBUwmTiSp/hS
K0cmoaYlSQGHxSIhsdCLi9c7i37Ods5vSzlqfgBxp9rlgsWGqj/fTONdTJcgCbm0T4l7ODR4Q1f8
mrEarutKV06TurB6o5T/uUGLQyG+h5Bb3IQbyXFgbQ0fBfn2xBqtPGQPtX7MsAYVCOF1mr2/1K9x
7VxeMk6n9d4iYytJqiB7YC8QGOQGW9XXt+f0+xpLIL+q4cDKtm6/jiXalV6NRIRQviC75pYiC/dB
HQxHtCnkRtSAwCllF3gltUpTI6TyFfkwc6ko2AMREslSWlmGzK3EiEkz0I6iHPG6cGorkaC6Xq0j
5XpIAk/z5EXFAiyz6DUtyDjSQeh+a8tCef6Xy3FEVCnOL1UMluMmwmuVXCvcUQRuQW9UwTx57GsK
asfeYIN+AE3aw76rOL8Q7OWrcfJK3ZNAK3hNL3HjfQ4M9iPmEjH9q8yQ+ukIwacs4ebv8EroCrb0
FrL3oIxP6BelNVwgmnFSPnSRghQcwv72WspVMgJO7M07PVVcPt+tXe61WTcYMRs9UIj/ZLL5p5OB
Qog0Y+vho2nh1T4HlPYlT+x9zTYBK1liR9TKAeN0II2sgolOCKpUkchBbi51o2FO3oeHHLPzCszJ
fDpY3MKqAFG5RFh6LGLxZ91sUAsyTcmchPzJmFH0T1Oqtkom8y+OqIM8+1k2it4jFiz+qaTuge7f
0kydAgLb9PfMUxldNHrmTzZFAMfC3OVrCGeA50K3OSCncevtONZCzC4ES99WSbVQA6A+9atyOYF5
V+8kWjFOZnJxEMNzYqRVqWuYnS4ae2Yxrvo/Qk4ytwx5lS3QwjnKZ/YCXLziakoXmTy3Ekktin9N
yj2Mirgi/0bvZOnf5aiFXontTp8G/rjAIivQBVNYUqsxyitUzrQWLHrxXHk9yEO9ksPDngenGJOy
Rl1JIFj0dAWDPiaHfrFm3jIXUR4rGlGk62Hf2MjJEEEs7HpRDOSm0KOPdlsyPbCVFW12swyg/K9I
DFws4e4PKx5xo13ajZQlUeCGTVhdyEo02oQEh3f0KaDQ2lwkGDgjQXEc4issKK1z3U1FrUW35B/U
fAYcbWnnGF1cj/BUlC1yWfB05ASNWduciQ1OtnYzjoQdVSVQcqIblPYpTRF5U6OeSf9g7cQnrUG8
taec9B20kuiX7g5XEhO/Dq8/hrD8REMLHuZ8IfssZePLI+tAxrGH12TnNDsK7/adUEzS/7z6VXxR
NO+6OkXx1EKf6e1v95BSrWOk1ZeMqRG4sXWqxuLv8QxH8XG9bX4hyWf6GqBWUjBcJbE/r5Wn+xEA
9RFrHUJdTj9OLD5/uKHdS/hADjU21RiSsLDIED/fk9IJ/octYPiRDLtwYLxOCdItAlb0evVnytK0
vHNWwgyBsX0dBh4ReYozVtT8VrUcWckWtjn5H//ueM8nBB7z0EXYgKMW4Mtpg7juTCVnPee52mRB
5v9Dqq950p2vJ423Dijiku4o42JF954Cb+zEWrtFswxR+FwU/9vT9FLbir2qHDfY2X65HOjVQk2c
6Pd2/axJI596o2JOueaWG5BokDtSyDn9neM8YVYK2QqEd/T2oJiR74svQpNxSjFutkaTyPPMn7WV
6BQHwVzUJW0PEidOh9Jz1k7fbKMRHr2UOT7/X2Op8ujT/hdpCnDXDpKevt6XEKiVVLZ/ZG9WkuTl
KErr8uQtBMbgUb1tfcu0xuYi0Fkv9XWWWQzVKZxjThQCdLS/9odYr9MAnbmzfTTADW1oTiDHQoWE
lXQz+9LFKbdKba4Irp9X/jC7OsyP3BeZ/HLAclt6m1bDeQJBmKPiNVtwdOXWZ91DBfgd1soNg22n
32GKca3AQC7YQKoYM5Lqrn8bJm83Wc9c2H7MeOrquZ+jv5NWv1y+QeX86PLEz3+Tan7BPMAI3D9b
G18q+w+YyzbRnambY2dtj4VHC/gYGcQZoRhF9FakUQ4BdIHRIhyNJ87KFO+0BszAD0hoEf5T0SCO
hKy0KvResRJHAsI/Vss/mvpiqMPoQIT1QoefuApMGVBgDTLVdiAsCdXmRbcIK5wjMenoug1meRdS
BlI9G/FZJsB0tYdQbz/uVhVag08TB0MdAmZehImS8NwaHxDVtAHWNezvH9Ucziug3Tvd5o9sVHzR
nXBwlF01gPtwHC1kGVxxso3KKcoDvAA/zYFfdAGcGLjPgAov10/AUbkylKBKEiFVqZcBCVXcd/Tz
h/W+RkwSeVBjOT8VfP1LHvAhexvkZZtk+W5EStFGo2HKeMWBANXB/zt7t5yv0ZLEz1pFMhc8Gj3j
jxSuH1L788iCGFjKA0f060fFRXgKM3nB2AFzcQfBwWtQ8B/4V3We3nSL2UpvgqGztjIRVK76PpjL
J7BCLzJ1lpU9ed0yc0HWCsh+e3ceZep58Wq4Rzkxc+EPkASWJNT6+hsGiTRPZLLKCV6sACQba5bY
AzVzNlFjo1XOjH8grt4ZiWBhwffZ5KLaAlh0p7uH+TeYBCnqX1f33hcKJMdwYRhRX5lCAT6hcOP1
MHvp4zweOoDcRA4ys5nd+IOy5wKpqtRyBi5LIpnVFwnYNQGW/Ary3b8yCdlaAJLrVfbFLRTEKjgg
k0gAE1rzltHMa3i0ZYk6bQKCAz5bu+Br3IvnDeWjg9/jkXI/Dt3kyTnzGtpgTryrLfr2zQwEa1fi
sLPpVL01Hp2drJe7Z4xFfZ/CYMp1EFkke+LUcWDn1cMENdf3NfoBHarBaYwfMRD1yV/RAhfTrRqP
+ip7B7KwV9WWaX8XJ33VIYOZv3lRpfcsj8DC31O76+hzJP/WGz9pFMiK1lLr83axETkCLYCcRQTf
Sf0xyIucl+BnU7fJ0n3UacnFPAA2ueRU5job6MbnX/SPEBpRYyzREaZ4MNdmQYxc6N1bY7ZCEqLu
YLUZBAceb7nwlzZhDHz1xHW3dvJMAQ+dbSyw8HLObWZFqXE/I/PebIKQ0C3ijZNmuAkxQYv4Rlw2
Y0pr77bxtl3Xi1eNnAKfvd8CMU8h43ieI0aOglOKmHTLAvPoz1ICrs5feaEF2y4yAS9iJXYhLnZU
pxf1jQx4gnfVb/HNSfeToNNCPuUSGJkqGSc2oi4sPI7uM5CTLyHCOwPIC+IyMPpRep7EDyyQv2Qo
BZnURPBowzJmvjgthruDItR7juJNJm0CjmPxAFK9TMMkjkoiwbYXKSZUZblM/AQn6XBM5LKhciLl
Lzk4iAqgnEyWnbceylElre4V7di36Ga4JIw8r1AgzQAUjovMII/fJHlX5icUdHJVJ3v8FdK68evq
Stve2sa+6ebMTwJ0zhERJy8zE1yyuJTE2enb06FPILDSohSZnsGH6zy/xnlwQ0sZyk9oPk5GMGIv
qVyUBmFJx87rvIYkbDixLKg03a/biOROHMRYFaL9YygGKi3LHdKGxf8P2hIsedLonkVuwcxuoMUA
c37dE5e6OS12GqjwXK8W0IUSfz9XkPRNKpgvDmUgyLw7B4YXOCAqTFHoP9A0r8emR6QPX638lf5x
96uQUwi/IX98QEPbAe5ydVdjrlVrB8+r9zE8lauHdEIVsxrYxQ6IpNp/LpkRALo/Aj/RKXLfvIOo
IL+fQwXvuux5zuUs5BU7bum0Gl8c3UteDeVQBsp+VQEz+v3T6AsC7LVWo7HPcUTGhnktWrMYAAsH
/SJgv0WwuVkOxtkBj/FIa5s7VETAxZjBkeBL8aCiPdWO9g5Z8A+ZHZAyQNBqsW5fu+mjCVWyJa/r
9MlacuQSwXLgNZz7QXQaoEhxaUmLQErCTMEOnUYwwn1RZE/mF1ujs5RUDW3HXgrK7EFGZgCZXbvd
KEKU5YTH1eDPRBsrpGRhPuaZt6ZpJ1dKyVR6PORf+qTFp6m7j9j1cuLZdYJ5RDIflBMJB94IT/Ae
DV0eDilZoO+r3uzP7mT5Kf3Hxs/NgFHSw0Liz0QZVY7NGT/dsTzsnmur65ujdqeUCTbbvaH1NjWm
ej9hzCttVO0Ik2aQdAUe9P22EPFasUx5ia1GgaffGYVHPKKurjh2gNeMBiw4q67H1WgrD/kuX9P6
MTOEaT3POY+piX+6vLAY1TWArh4Wrhuz1NBlQSCEZWHrSWGlVe1BA3ZjTG2PeIuoEpHygMzVFRKq
Vm6xcFG8J1cc2yXqf5aNRcTH5jw2FrD3ilArznqQ2MpEOFed0FWypNoV9dNTLJYgnBimvloMEH/p
H4nHATOu5sIdMwIw/PxV1QMtBt0ezRT8yXWgGMtoBD2LgqroBlK98CovhgqJEgm8+Tlyqq+naQSD
4xZhHvUCr96/Au9zKAf06H7GhMJDbVup2ipff1kJIexIdXumRv1qlRwo0MQRW3KIey8d4HnSz0CR
fMIMy/GwT84T4rT/UyQpqZBU6crDeTmvBgwloBrKAKCJSKq9ALO1Yv5i5e5mb0fMr7EWK14cVUWJ
adcJQoPlF+MtomQ19Bkpt5uSgUn+nwc86DUQ02jR9y82eiZv14d7kiYWhyHd96NP+pmPhJ3ySl7U
P73tH5h58ClrZqvDEbQfh9BGzE6Ey/9AlyYxXBTIVIkqQ3GS/5jK1j1OENTetuUdYRvHpL0Hf9GR
6iimszUnYH3DcW3Y1ySk5Ww+ogljYkw/MlZaQZolVAhbjaru48LMXGJLxRohGbTVdn8MvLA/baFT
TYqF0AEn4+RnDiKkPpm1FLL+ObeEOp8vu9rA6SIhCbbnWvfPGBOM1aXqC1v5xDBQRhW67+iS3tYB
gD5j/dYEbJPxvbOBJYxbPThRM+pJOH8L2/tQNWL6UTimbo58A+ZazToIIfSJYs6+tqIBGwVYdwbM
mJHj9kC4UGo03AtcKiPQq7RRF/BCDd/Pb4GDDRcbHVv3ovGJlDUEFFMphjSnDrR08V4TN9Dn8513
QD3d/oRaM+sZKqZKhBm7sSr0qjvjayG60Sa/3ixxmTiIj5vUste4/U/lof9j+LVYVWem+vznDrVw
2CORqhLEb1ik1H9/FQMckg00k71ahwq4/x6WDEA2c701mbnWJUrztzqy0mILmb1Qr3VRzqs5IVM0
/Muw5aGUGKsAWuaNY9N/USe5gcOLsUxVJmABtVzYvBJe1yLCu5yzMy8acehmOinhqVZCzGb9XVSi
fmH5enK6j2azG03xbMtMfCaHeddUPGbsXQP8e6uxECGPph912oBMzXw2IVz9kqndEZoDJi1ZWhoO
QrjuKJ+PSCvK3h+qHsBGg4OXj0JiH9k3PfhsQY0z8w0lZkA7a9yeuxk7phN2H9zLpJJaQUoy/Cib
ypOQdQpW/AYmx3jptRpXmw2RmzXjgfcLkM5OaLFQoT31NR8Iu6kZI59erCvy4AtjGc0V2aX+sSU/
hWtY2ErXdGiZUbTk4eD3KBufI5v2YgRhW3/5LO7hwoWWvP0dGxwj+lEfsFtmLmjGNVWed9HtYtVX
B7svNy2kdIHTTwfkKR8Z4K/AZbkvC6dk3OQFpptCj2n/TLFt4smd0xfgGpZwW8RK2M9A0inVwYBr
L1p8pveykYwvss1KQy3gnjgbAayWMoxSZFO97KjcB+oa5QAzAhCoJokm4HBTlA0nRRgV2K5YUD0w
tBirzo0nWFMkjPnC6MFenGXU4/jUDVuxSN9BSicH3nvgZSoRESc9csdB31ocZYgv14yq6WII+MNb
cz1o6oG5mL9a+WRCTVaxBLN7QpP4fXXcgobOGniUHZUsfCfMBfP2AqWfUO3m/UphQWlfGRsRPiaA
DLecKztGgAiuY2ETd99UT76XT7gh2IiN/WWWUd/JFgPfHeYUOJiXvUie0n59/B2Hq8ljbPoRIVCc
lyqqeSUrExATHwlTHWsjBqg25bAQm+4zMFBs9/dzAIso0PnRiGhtfHsTbt4Vgt9a6FN/RYZBN6EY
mBzv4Ekp+7TjT+9WIs+MaG4HIHRcagLPuI0he8UYSKvzKp8ZQVj2ApWZ24Y9oQ+mD6o4HJklI3CG
wR2x+LVBtuPVJ0wL2J3dcDKZLAIFyRR9RO+HZJmZhvMP2+MCrARdzrINOg35jAqHaEud4ksEVNnd
Z1IQwTQEapCHHfLzs4vBhy4r/mx7j7yy3Aqw23M8ji1mjE1M/1rQUIY5hIf6Iv/Cel8jzHfIPrRA
ciPyqF22hOoETdj5ldFGOj42LY8lCW9n0iqT/+n28mz0bsVOAxW7MLJSj6sbWcudwn9TjrI+Wjnj
LFDVwsfMIr+r7GlxBKCazDrOS1M76TAo7oQRoBE3jBnwb28tFC2ioPsZvE1yyaKfi4PSU4Jp41Vd
RHbrSryi3vKHZESSrE89j2wl4IF8gcbacfWC949/AWe7sKO5unk+4rXKwXqovNwhChNE4tiWoX8k
Hz1Ysl9F/+PPYWj2nMBJrahDm9G9Hkd0PuMxeWzEKHFJ3CLt/12u7ISaXTk+AJM5FeFDttlj27WE
CT7dyVB+BHU5ZZCsD1prOkWcDD0lPvMHES5rByVcybK0QovGfasg5tjv4hfaqtykNrauCovj3FTY
JW4ZsvVHHg4WEhKVe2VmDCMC0Htu+87SSEJjlnX136IY5VaR1oYsFtO8wRRzI/R9NztuJWzUS9k7
4qplrSIQnLrcT70vA97XTIHdBqEE2TwFTEstegUNfxBFh78FTZz3O31gRLcJ1DwRCBXsIDMXRwJj
Srt5Uu6PpPdtjs44ce5Ecwh2Ogr1i9q56k2OQ5OtQUGcacWpnG9p0rLHG1knKI56dU15mZnt74Y6
PIB/uQsbCzH6G5YL4/t8JtJtohetiQBa39apn2ETRTNH531sdmrsndkLtjbmCa3MvmEAymGp+MNa
gech/kvolCjw0ogF1gdBmWI8vJHllqOYcOa7cES/3W3rZZuUv7zeEnbJpGDYC4sip3uwSxccWphm
tTc+jXXBMk4UyK61IGlkZaduAIF5bM5OhQ9hwy5H9XH7GIoSXeXMSZbRL5ZP+O+afDwB9uQch/k0
in3C7AdwSV3kWetue9432WxotQzWxvm8TqHcMKaCZNpszG/ZePW8RbaWpQa7rX51MbpLUxyAYDdL
W+Um7e3D6+fS1+h/I+lXrmlLAQBXpRjdNIxHlF8dLfQtosuUjCRZZX2+dWLQ3PuwhcllvrxgOPwR
ZBzRmtnaeyaNsyUl5D06+YT7CKOVcNB3hRP6qjGVknJ33ABNL1LyGpciIW+ArhnMV5r9qdPnlHpu
jCzEwUnA4bKad34iae8Dogs/moxH+zWXcBEbOI6NMpkKUcPbX92ntbaspQpkmKCw+h9mqd9CoM3L
Jp1PNjV17ySIEIQe/vZKOJ8+GsenSY13R2RUurepPrxnp7AX0jwndxCF1M16Y8Y9KEO6aUXXv87v
+WLYfI/Zbr/2ftEUYRXlxFf+MVWf8uE8qf8OQdjk34dY45CNLaZ20fiNi+cLn94hqLemY3yGZc43
e+5HefV+sdMZO4XUnyhoJbDQuwVBfWDOH2rLdLUuTfUzM81aKqCJCP3Vy+bF9WAPOM8fx6yd2Y/m
oJXFEoRwBYqGP80FnaRNZD9FI5WTpQROq41w9J74J1G/Ha9j9nzmdXvsHDus5KsDgONA28BGpjtd
PMZGrfqUeoTFn7heBopJBT6BPth5B2zLP1WzbzpYp9P7/xkqDRM19Rw/9RRj5f4ZU/dybAGoUglD
yFIi7BymN2+hdJXHppRnNqfBFfhgLJKrRstLnZLDlfG/tcdLpBJL4PtnwGhecN9CepKPowuiOy4p
cklMgkE4sxI0zn98ijIL7yw5S8tgmX5K67GXpWw73zw5JYxU6ihIGg6MSILMKIAuODsWU08Ma5//
hknNzIRjDGX36Y24sepMeC45/kcvyOFgGx43CS4GxeMrH7iAntVDdiw6iIMF2Usy90/KqbaGeaBR
hkzSJwI+lTukWoE56Ge1lsF9OojmmqUBNioKRMzvIigzkY86kgfU/xwgw1d13CQjOxKpny6IiiVx
Fu+bWzpLHoner1kWDswvM4t1jMKhJPHD3GyESS2sK9uTSi8DdWB41zH6pwloSjMBbigD49wu+MQg
RnfwJ29gi4L/5zRjg/eed1S2EJgu1LW9frBrSe3FH3ChGiWKVWs1g/6eVFMCiByPF+RZ+SP6NAwm
rkp34Vy5XcAcp9rgzS998I7cvPTPfNLxE5tCGNiPf7tzv/GAlOmyLxQjhsnG8JT+BhWylYugH/3W
N5DApSXwmuSgAcsHtc2noBacvycb+JNFDQRn3tOHXQkViQwS9wOS46BJT52Q79//XrvuuDIzbR5Q
SX+50LrbyikNZbrqiSVO3EvBPl3GMDzPSgM3IudVo41v4obSGKcQnvr4rh0OvivQfjKCFCD4kdd/
q3KWQiZ3eqx1cxw2Z1+Hl8GpydVGQYgy0Q1pk8pe5gaBOv2n4OsXYpz4pFCehtaQ/X5sfcvVWLQ/
XwNrjJVyoGDaXnAAiwa9bY+BRNs4nxpI54cwEMVNzb00ytri0ICOZVn0J2SzeqVXum3yV7REv+mT
xDasejqBJo2UfS8FQpEHFj4cs0oC4VkG7BQ6C2VuIWM7aCmQFgj5rCwHBBFRc3KS8W6B8lGH0Aoa
XHo0u3OerSYDVG79nwANmg3Cl6jzsjxNnoGPf8jZbxKAGtF3OAdAeml80CcoEeH4VLRIsZWMEJ6b
8dUH8yM/4m8PQSR3CIeODgcn/cWGRmRkJhlGbg7EPFMHHMNgzpjMGUSh0/CTUU7YlVRqKa96Rf0n
Bmmy3/J+xFQpxLuGGv8KTit1XA3tKTsEcJcPu1GoN0ir/oSqidunlv95l88yLkihhu9nc3B3wRHv
T3AwavxTXxZHDDHfOVq1BZ3RpD49Egxe1HU+/62h7WOqpO6ASMdnbV+uWsLxprt5SGK9VjmsTV2x
angKTSyEQiqTM3BXyplibmbbo9qScUu4VFwwAs21xOt6Ns0s3DQ2dO9oXZ2fri/thmGlyxMq7O1X
I4MWakJurDeFScsv+1QUzuXjinxmNJqFpHtNMTwkraTIXu78JCxxbLNIPTAK+59h08oyQ+EHppz1
rnIhRwR4lJFzXMaiQKqKVn8QdmkSGHzoomhxHJw7H/2aoGIOZ55oGXKTffmpNSQUDYH02odznC0M
j1R1Ut1Qxmkl7Lm0TOB4Y8W2cQOkpNW50T5nQQKuKluY97RZwuFG2NbYeYduNuiZDcHIticqi+ND
WLsdq5V28nlyLN4nEfkivrLSsAJdGg/Pu5uIBsF67i3LC8A6CNfwUyeuWKiqgvkvGy4V0Hi4yqI6
3ntlng9I37/rZRUywsIfpmF85EJjwNQrSy2FMOGyQj7nlNwD86Rvf7yVEyLsmG3FFhVhDSRFMyeY
er5ShWwyIMz4XKltiB/QuJERMmjoQq/BNWNB4gxC19+h7bJgDdRNomhR15cyKAlDF50kpRD/cDlv
l1i3BzvK8qzua9qRG2A3IZtYaThSidWzl/r6gA72Pbp3OLTkXH4nawC5XhYpIM8s2NQt/8PoApYZ
6+31wrwsi5UrIHr9GCZ8bCLwioAjf+wVGBsAJdfuZHatniM82PaNdgRCQ9joUrhIYtqH2EieJZkp
V54qUxClDRahHO1an6cpxz+4C06sG3ooMmF+SRqQE7hH+seo5AGi7ksQSgK+BSJfSFg1GtRLlDEu
Qx/F7hTdaNl4W5AaJFCDBQM4z+0YB42isKBdNb11/VwLoJNfppBHH87bwH3jowt6aQUo92kfKthp
oZUsAc53OqVqfVoy64uBn1f5biDzqhD08aXgC9Cw2zaKDoYml/VFGzsTxQRk4WAzUTobnUeyN9n0
YEALGx+Mz0NbE8MddYOrWEh/BvW40XxRpB6PTIfbc9HzUF4XK8pfY10vjKQ5vQOO0n++p1aJZEXE
HyTvtYOorLCoIM4aNyKtxQ7TPtRkIbuSSOlXudA4AhE4DGwCWThge0uWB+ZttdSUXbKzZZs/tSfv
/YJ+HNXlT+xZJ7GRa0eb7UNalhWEbc+ULUqxnxTU6PhrXwvYqwuAkQXk349UL4r6RVM1GXSGGBOh
zRff32A9N4XCFJuQi7BDgACToipYcLo1u6E1HlGqs4WCRI9WSvC+v9nKegexToClrEiPud+X6KSy
StGy4RV2P+ExrsIM9EIaus3VVIKDImfjqYowE3SIvdfDuI6JFOzR47pQhTjs3eDg/zLq+D0lo+tH
H3swe9SLcqy8DoN0/ZE+qBDyv8EBcUlHpH0iCRCeaE+qQQ7+wC1f88cP0qfX9ux0wG9T1oZl8kJY
HsHfCwufCOCidTF6B2w8x1R8fiF3ECO6rMYCWw8rDGqt2zR1pw7gDR0Nl/x86I1nga2F0NXqbN04
P+QoB6uzR4FXJLnM3lFYHn8sKmLpexlaveiWzCjYoKx58X3BlpkGvm04HTF/d1PauFuJFgIPPoIN
WxHPnh6GHoD2XT8Wqx/s5FpxSnNW+NZ2/WZFalMFiXrLx5QXNyvaH7k/8RsdmdM34w60LO+NyqPq
001xeUfqP76rmE3kaTsTgc3z6Sm+XRnFlAG9XBdKq3HCNVFwvZoGIrMP/ULFhI5RUBCY1/AvY8As
FKPJjkz5xYvDuaQQlwwCpeO8Q3YZ693Oq5w1PVHXp90U5Nj1a9IVh4CJk5AqnTDyIi1A+god/3Hj
/X2bEe6rENn7BAOD2/AVpZn5O5/D0kVcGYMFZa+EKVAKkNhPS7g7kSmPaTuhZp42uOxm3EdNu13Z
g0b7wArS6hxsX9pi1ijmrDO2ICBRyVigs8XOQxZx/CMStpxsryIVqDHY8kd7YF9v+jzCd81mZGNd
FOPlp5aURqtswuBrZ0lBLWVrUlrmYzY7d+s/cINMofJERurksSfaBkuJi5H9/+E1mF6jQtfEslsV
1M1IGWwzr9YDXqNVDb5U+5VIbInNyhh9bMkxgqGtGUoXIOQ6s1RFrWR+oM3fEGeofHOX7RVzHlmH
xB7qjfc4blxCQeFD6thPZALWDYCr2cDLMbbi7d/ijHpreKnfoJa9MMm7KvUEwtEZ3iUAPU4OlWNJ
YwWGRZKbrRVER0ZaahN/RQGIoJfbj7Sz01kKj2lRaI/6C02F0fnvqEc/EppEUmwUP5NHVCfIJ30A
L2po4AP5cfmLYvrUg7qhid0lNzQ32hvDYDmWNWucgVz8DEzpsUJqcwDidc8tuxqxPwaQ3g8HrMZX
mdgs8WULTb/MILFPUmyDOSJhr2ZTfNUfA08pwfQw/v2HOMIl0Q+WECulhXb6BVSrZXDmNWGf44C/
rRkMqVaGYSrbA2ykEb27Fu5i10QSstbT52h8rRK8dlgbgVlVOmjwHlwRet6AoKgs7NoR49DQZ4ip
OBhKECwRek1L+xVuzITO42IJulzSGYUouz3GczjV9dHFdH4En6nSdQMc3/nVn+uWHzE6tNLwBTyF
L84wbtWl2YcBCF/UUc3jN7a4x2afAsEg1ajYZth9owTxBXdjmeEFuxSCqws4/pFCHw7JbIicRTiZ
e1x1F7GlARQ/FGuigSfHP9Qx0MYd2f8KxvNUE1dg3ZPgrm2xP82mz2aRy75MUxUpsjXcM3s3DbrF
QI8rFZjWtiOIXkWm+BqDSVbnqJ1FghMVEuPLPO5T2eKoksDI7+aF1trYHg/LqgnnM843HZAd1vQA
tLpTSAfH8G5kEWCMyVNVwfi+NpvoyyDK9kZf+pFGOlvctwDAVRGFBtGbHoqYAtbXwPvaLur75OO7
KXujh7h0Uy5WslfMWu5c1WXm3LDle3o9y8oDzPyQL6k8uQvKibaIgb9MnX3+Hk2F8slutLPvaJY5
6Qo4uZZ9mDjZuV/EKuPv2WmvpGwNif9EMHPieUFs0I/j94nAjrGBP528mGmOul1t5Q/4nR5iJ1Kj
/fTKdG5b6ShrLEZ6F/tfEajtr8GReF9c4sj9GoSBLXzwj9gTmC/fpxNOG6rmCrmQFlvwY3voF3+W
wgzob8fO3iRLof4iCZU1JLD2w6BZ8d1bA5kY91YAiAU29OqPOsHD0h+/lCPUOUI1BtmqgUSIwRt+
lrQNVihd3M1nqjqUHnE7EqlYY3xH+qXSkEV+X02UcU53xQvUo/jIZHSjgBUO5IeTH8X/DRYKdUEl
rA1SYyBZe82r0Cm4mpBNRqJw3Gfnhdxik/CrDzy5UgppTSJasXlN6oQqAG+tc6rXObCx+CAdvj/6
0GwyJJZp8tVOhB90Dl9eQOcRmP/3xgtMQF1FnaieW1wfsdtIdRiN0E4s143yFeBF9dJyFpuhlMnN
wDXcJw2RG7+hNeFqEMtKEXH+GQoXYG0y2/Xw2mDtCfNOQYmwXsqpX1WDkkAVAw/KSuedn6WgGyiS
UH/2zCaRtX8rACjXsiy1VPo7X4lR6Xx7pi4oQzcdQhSWV5Clj9KBKd6DGS8cT1lLk5jVupVq1xsI
vL7q75b/6c1uNssmmUKHHXLEf2+7ot+2s3037dpQwJWKj1eAfNeyAgWLCwL9Qh1nN5QgjJA3c2S5
x/EUHkNbg3m3mV3HU5XkeL4Z4nKVGpg2NjfOcjGQv5L3bEsaShdha44U+UsIIJdSik5BmaqM71nr
K4FonQrgiex2idJw73CD2cKZ1w0nFUpNLDMM9W7D33nh2nK/Vr4eSGauHx+hJLT7MrgUu+UN8ZSA
eEHfWW27WkkbQTeck6/Xiny9dshzCX4jQZUWKef62uUtcdMcNBSqPBLOBHo65OfQ7F8I3bdwPSSO
YSvyuObGZaDNxqFcHFnWcsYwXRQMrH7/
`protect end_protected
