-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
czYFcusGR/CifCLzPj8Bc5ygv92gGXisjeb1j4zuF8/Q5d6isjcXeiEQePjBnchSdxMjasVPRWAh
tMwoKd2bSJTqWP9jnpAb9EyNg/uhiDRXhGL4KqoJCpge3vnvAIdXETaZiI/VFlfBLBIk9iPzu7kZ
nmwSFyMFRkzGWbEX3u1ZoQmr2ZPKD2HvMkJS3IJKOl651XpyT84ujyAyhhrHk7I+126Nl+Wm/ZZP
GpLPRIs1k83SxkPr9hsVqAz9DLoh1HIh4zf4gkYCsluKbr//0tzxjwzJ7d7SC756IO9XKALBIkXV
eFoXfhuKYMh4xvocbcibNFpLPCc+fXB7ywO4FQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20864)
`protect data_block
75Q6L/klCxmc0oIoW1t0mB+MkW8uq8qTJJVurQ+dbm3JZgl3038YEcwNiPFxMURIlNHbN//yNpbP
MMVc4WGeC8Zv4qGo9jSEhi0+qHoPpAP1qxKzAqHYNOrCqVD3/tU1+3AxtItYyOADXgRVLvZtO4gt
GU99jCHs6I0mRVXlUSL9Uv4EcsT5exVhqDHZRzcJLAoTKpXLd01w7DbPz9Mwtf/sQpFEV+eTa0mU
8obdUlhTI2DWJDGMbo+Xi/v88bN08lihUVupsJKHUKm4VDtCM18J7HaqTI6CnSuw0ED1u9N2n/up
douo/KbagLVIZNlaYVKdRyFPEamyCwbcYVCa95dy1dTS5SqIAgI26AR8leEC/4HFj9MtcuNMJ1mM
iv+VLji99WXhdSj9i2yQ+JYuAjlC1C8vbHIEKWx4yXb1D6QhvYH36z95pv9+jHHN/DEEyZdtbYg9
31DV7JA8piq60OBeazqsoKD8hX2I17/TKff2C2XZZpvuolZxNJuHxfd3enMtrcYqfO+iEcvYd04c
fEcgAmgMYABEKWFN/OWj1uilkpN4sEqTDv59NylQjwtyH+ilyMJi4uMw0+Nx26djtjHmRbq1sPfe
E/aKiWBvpGrMWo4AShOhtSyBUpuhtgnsaQwdTZw9yxH8daI7G2k6QwHajJyn7Slo7QfD6uNvtMTg
nCjXbowZhDJ9Y/3JMJ3hbAQqHBVVy7kSSeUDBiSFKWiMrCEXbZThqUAB/84K4m/xkgHtiGrZ68zG
3x8+5/pZ4XLSJ5kFo7JfKrs9vb4jwNQenE+AuQGP8/pXoRrAH28m8Net3jxHzU5Et67GqqOYDG1r
GG2drbgSrxGfdmzJMsFm+YYxjE3KJO6pm5zmM+zi5OJezi1tVDZzKqQRjhIiz/9oXX8vdnJxK6zT
JPYq9qXmFYionld9/fgG7SPJvNYGOVScj4hI7yFUpgstJWl1RroOYlcuOAtzs2XSjF8AUVg1yf1/
sMjoCRCN0JL/pm5G4OUyzuzmoi8O9CeByZ9aGvNprXVpFsQ1AFgAKiqZ522VD1Idxv2UI9Ij0x+s
14YlB+eWNeDBDVKjPUekj6bLKVcXeFducO8j+iy3UEFv6ELiYNQ1bJ00yJN57rHfhbOqG56eSBzt
i6RmicZGis56cf0XYpjRmSw5WQeNbpkX9rLYyD77T84ek5ZrSGcriK1t4y1425enEx81B4wbAu20
VsxyFoQvhRO9okZdXG+yFz2264abJrD0QxL16uctz+SafGeMotVa4KED8hpUHrJF9aIZlm0RxTqz
n1oNtre8zWs7rR+rU08x65ijf5dC8bVEsqlcmau3/xx9N0zoL7MeWwauyQt95b+otrdWp8RG1zJM
iPev0aMCHbsKKF1qpYsTGREZtLKwbx4VxQUObbdZzYeDFvAPS9oj8Og9jGFV/xFwHSG97ri06XM5
z15ofDs6Q/zExMz4Xidos21PcXjU5CHWEFVXgT0qQUDPVilDef3XkZItE3sbsP7uzupVB/IsovZa
g04LIJpaxI2/35XH+uYyw8/HfdQGcW0K3cBad00BpjwJdd63APE5M1SvecIIAywI9Ja4dHxIw0Hy
JIsbqbpOr2X36w88iprxgoqXaje3mGFWuL5IoXL0xx8ixElLVisi+KEkZOmE7kh+2GLh8v6Qfiw6
HKAJoov9OlmLg5l60ngjzxBgjfXMXHzOtdHdTl3qX7w5p3V8UdLhrsFJ89NNE++iFm7Abni3aucv
HpCPlarUy0nbyT6RITU+BLVpDbB6+lmiT7b3dzXf8cHeUzt1NaI6dUjUYp2aHVdqdsv7BZT4xx1y
zOkE9UtE4cnewlVj5/b3SCGU7k2slq5dO8CTWTgTzTz+vVcMIA6gDkuPHpHS6kPbXHfmDDb0WcAu
DV0bxQRk3ZNdUClE/wa83bthFiQBK4+4/+XfV6fGw5gfeS6r54aCUtRUlHN5xOqBbisOZPHhAcsN
CN65BleLWhnlf3jO8bZwUEPoW9pg2QrieFzxfo3ZzBTAnnmSrsVVISOr9bIMhTlrVYCp3Btk/ywL
otj6fraEVb9P56aD9Yk+vWw8jX9zGmP2cnh1opBzvAgkBPQPD1xV/Sjtb1KvseKL8c12wC98GjbQ
dqmD5dfcemalHvl1XeRiGOiP/Y5wfk+KkgHdMZTu+PWS/eAbVGBhTeBrBuDs1qGacZke/X3hnXap
ZqmhTJQsu5StFTaolHgrlXc83Y9KXsYjNcWO2mdHi+5A9lXnUGPQYom466xfsBhzpTwDiRT8sf8o
1Em7YHsIwJUXmcDjXc/X7aViZCnEAPzDhq/vQ4eMw/ZnN6ZF2U1niMIusakL7y4FbU8eoCfKfcld
n74nD9Ex0r/MrUKRpweS0M6RmM+IiMTux71Lt0V8BoIma2AyHSa9XBjIX2Cbul+JOqk/rMBMTHgx
LexAvVc9SOHJ0yF8lI3qNKXQAwMkv1nhCAEJqVyrCGWebqmCmdMCV+r1My6uiZcZ8m/7AP6wfD/0
7KIRCi2p5wcBL8hxBlR91KRlKh6nl35IDHqEPQU1xp7v7W9LrVxO2XZPwIKcjMXxt9hiHiPB8swq
1pOfAS1zFcD90EaPsKl9SB4mMApCyVQrDf4Txzm17P4oFCLOvVvDAHV/jTMsfwMHOqf1o84EpS9j
cg4bJLUK4Dq3N07fp67/MRCTWJE6mZEFWMW74+mrXDG//rALGeGIXwuy1CbQ6rYIts0zpfdUrWg7
p8TymTfk1xqoUidfHDzjv+/6DLPW9Ix8/K0xPeBSvoTDfO7BRKMKSrsqrs1pRJewvpB5f0o04GHG
Psjb3ik81wxaD5XTPiAlL81mQuvPt8wbADtmpLz7Jud/xhng/9lOX72xnKM3qy1u+lrAjWrQeqOQ
KNbqX+/jtlJ4vw0UCoOz1ZKZldiv2qmXvCRSqQ7MQ5BRC6HLpaudS51urq52+Lw7zYAKpqL4nyg7
+mg0HCtD/Clmam5OYz0BQOBfC5FIx0Lw4eZl8UBE/gKXCu2EMpaPG8Q0JRtoYSLTIYEwAvMRLqWY
/ZwbmzdPRgHOXqQvT8I4MifCIezY4fDilgBEkYqe5/mBMOwhgc8RLP3N/ovfEQba+PosFDzMtuDU
dQnw21arEQH1lhtZ07rT9Qk+K/WwTWyEsTrMLpsd5B2tHe5JiZcV3DRZk1fhsKsU/MNM5PJa9ATD
nl8WfODLyKsuDIO8n5wlYag/TN+NXp6Iue+KDbtz2Qzlw6vakVALWDzegVI/Wgnih2yogNU8fxqu
WND+JWbdzoJXUCLNl3HiOF23joSdHXSm6gDFiK4tnSSFQK2T44vCI9paj6L8GZFfWJiZwIOp8fGC
Q9CummqyKHVomU2jghHDhfD+oDNisWs3BovStWx2J13sEtGGRWesdNoExrm7vVIuRFHX3n9V8Q1z
stoHXFXxJ9bADmL5mpZYaxQ2NBown1lrbEOVSmAJgEa+ifCyzkKNyUz2rNEGGZn8gnD+ewyFQNoU
byzxZehnmcvLXSsEd2fozUbkq0nfMsD+VBqkuvrvgjII8gMlyBhw1vfgImbvBPUcumbBt8QqvkTh
2HEr/u+63W9UjIriCDyhQQJY+HMSS1f614GfKLOxqoVCY4NivWm8WViGXaRsuLG+lTpkD+U0c1wP
UIy6Ao7CfIR6OqLQYuTBWtBhcKWZdLbzohTFeS7PoPzxKk7wojhY1GQ7n0z37FqTqHFJCPu5c7b5
vg1Fr15IO9L6oGLdWxvu6giEx7ysUgtv3sPDrJX0X70RfIUoVEKWxnOTHq+yYbAPJQParwbRpAOj
5VC1YdAS9d/wLcHiJT2RG8HhHjIq+FJacHkQaHKFVbQ5iq45869WdYFzGCxy3EiFXWq1aX2BbRmQ
SvStpx/k7qERhy75ODM91raSRCTFYQuChJSRnVAGp45nClcCViV76CQTLp2b3arnwTxWMO6H2vh/
1TkSGcfLUBhAaTmNNNDXo2+F1zU/QoIM7UbZELyP77wfyl/ofJ9exveMhiZF9uIJtK0YKbQwxz3t
OMllrbjqHjTjrFy9Ljzp1pSnkHlhuAS09MWk+hoBOFEb9JdaZxENgsSqhAK3QJU2bksiieHJbKxO
rlwIHwM7fcFXXPM645RkKWSv9/VJ0J21RAPv+AJFrdilboOJJmLJKfT9hlbQvQO7QxgEblE/PR4q
9dQLBEnwcNF/kIIIryoKIY2aUvI8uxL1LmNWYh1UW4fozuk+Jz6SmKzj6iMM2Le87Hf1pibOggos
u3n0KXCp6P/SoIA80q3k6xfud3MExfkxF8/yKqCDvjYKdpOAM0lodbkRmpWLGgmHXMTm7UOdVypL
coIu4onp4Pzoye3df6QiiNYaWmDRIZQqETxOhCS8XeeReDb1kIcYh4USKr97vc5XOCY6q1oKcqFQ
jKId/jAo3uMZQDCrfM4C0hcBj+HbjF0hrdZP4JuEDHrXGdmCZHqDXIWQZ09sip+o5G+yY5TeHOw6
hrXeGF/tjHsYB0KgKRhXJs6YJ59PoT72asstNOe00eI6x+Ahv3/F0g2FPzVAFR9mhMDSzBlhyE7C
rPzV6XmmdvH6v4jKsuOHoywBC41f0vJ9Pjaq3HTpiCll/c2/nsxuobBOJxrh/aQhp3gHUtzab7r+
HEgRTdsQODAEMNvPuTqAEpdX8kSzYPvw1apdUyoi0u2FTlZrlyITuKouCjDovMH7UKlKHejkWabg
xvDEKPijIsmd3foQcxgYSgkVj4gqLd7yP72i8IfWEdmwjGIpFKlg6iZixjyWsV6regoXfobD2Akn
Uq0vNasuqyM7wyl0JUpXoX6zb0fTO/jfGONe6st1u0EzfHKVFExBXvrX8+FVzjYX3Iq5Xd8JWb32
pADuRHpYbBqZXh2/YmapK3I3HWBsES7eKOpm/i1ILWjMhKUxOeVirC4qwlG2md8rB74Gjg9A+LF7
esTK8NN+vl3F3K3QtlU6ZqYtj5Flf/GysrVMAIGGbt/MVJ2ejxah6K7qYY8npVMA/UWiV84phbZ8
KmczznzB8dkyGUkiFIpkKp+ud3cDjCxcUsWV4e38X5HHL/9Udvo8zEZphN+kGUWuO2hNcrjsbXCo
jAhiPiiEIbBE0vsjfNtLxnfU693GW7QFGZQQ5EeY+81pIX+c7su5EN3ztv/O/dxlRKtPM8HgsVPX
nu5UD/UG1OzNJjxwtESgIjTMwOVX0nuWLetjZ2DH0d5Z9t4bkk2KICx/5La/8j986JN70zq6u5zm
fKKQZAYi74E8L4WZR7fifPy/MjY2pjtqTbOf6zlGiuuvqXGAZEHjNEw1AR6IhDOwS1yKpVnw5wqh
Yu26DI4UsgVXHAxZwHaFyH2wblpSPyeHuwd7wivQWjJ2W7V2wPJDOn6TBj/ya0mVsRrnF94VpCkx
pOgGwtAeedLDNvS1iM1diO54cDjeBtTJZIrla93y3E+kvMF0izh/xf7eLlod+4ufuwmju7MblGk8
OAAEnC0nOfyHc+yHePsx0JhdEz/CHm/tICIzKPK6DBi7gz/QhDoN37vYfF60sNl3xz5/K+uGqB/I
zGnNCycatt2JUDqO7J7Tqbsp30mksHS9y8cSvXRrRhTMMkO3+FmUP/gEDwTUm191Y45YzCdwV0qr
ey1KBCiGOIKpheMQc0i0a2mb/nIHbiuuPt3iz5Mq7nOQeC8YXBFpneR66Iy2CDE5dvUN43KF4JLI
N1tAhZOzU0Gn6RNVfgr3AihslpGYZMTtAAr+unHqUD6hm/DbLq/Ilyte3LWr1j3X0TVOY/rgYG1V
oD1vFKLPOXzplvOZe5VBZYluA2ZL7HGMjPN1Monz8lVYPZcrDwWwpRhZ2uAlreE8/mmgB9RCRmCY
Rw0EFuzA7qJ14Y4f47p+G/TPrTNVrdQh94AESt6Na0jAYV0D1ngI6rWN53FXPLQ3ZrFHQDbw5k1R
a+SlUxtTSZMl09k6Mk6AHuiGCoE7PhEuzYmSmYFwx8w5Xh+SOiYQHO0XiUZoJFErslGxrEELEE0p
qf2KRo3Ir5iHfAwwU8TxkNuOQDuueqW7lFlZ0KfAraH3fJt0AkspNR65l5MJGja3EnP3XdzHfDX5
m5A/g75wFXK8WEpjjO957zdtN32zCp3OOSekg8foWUk2+pzV1I3wTUDbyxuKaJjT6cZ+sLY3U/Al
b/jSIfkizjawF1B9cNYQHKZCFoE20fgxAexJpcuat0xgY0fPkmMqqkUErFGCxNzzlnSujP2cLf2m
trCLTZx5Z+99PSLkQoro7PGVI/VFjWEh99fwJ0PV4UVASrSiyH3ap3Fw9cD08NWDMTMSZVfli5pM
DAIMEM2b9lGejvwFkqzEKU3/Ff7PolCcMeUhiZOqRd3bYIMgqHlTn1pNjvqgn4y7J27JyGo+MqIB
PcRLcixlb9H90c4dTvSf9+XorBWBmFDU9mDW3Q/AbQ9Plg7g3LmAsw4GVhxz0uQlGdzgeI1cRoZO
asWqmOMZkTjKHFQw9ky/P1rYTyL5U0nGCn7cA5f1BMJnKASFdw2qpqSfjfY0mLYXt8AYu4EVoLss
UcHPK7XTigGWc1WOuCIPMK/rTZZoe+6/Vs6b4nrAluWROeBOEN3TctnhhzVsZlTsWrvoWdBtwcmA
zXwEA6XYmJ7sedliEth1I6GA2xtB8q7+7uGBy3PE9jOwcL0G7lx7gtvVSrObmugFt98fTcMr1K5p
VEdgzpaDR27sbTtz/3d+8JMjyrnRGPcfKSFi8qLdVvURJKCNDhU3SH56bju75n3jzciE/eBm+KSj
5K9EZpzO8o5BUsmnz9NXywUsVQWzTFWy+ZaV5/BPbz+Nnzuiqhmc8+5bsFxL94mYJqcZ3R/6u8ni
cRbYHt0bolMsocf9VVFo+EUJXJhh3cMhCnBNmIGOKHQtEB3CbXBrdSxeM/jCqN408TCygulb71CT
PA22rAt/qOW1O7Pu375/Jme8DW1kh5zoVAQoZaDxxRxLu1s8xP8ibNUrBJqWrPpT3DsC1dhYZ2nc
5C7qlDSwGKhu8MWYD9RfBPe/li+X5ttFjJoZzlr9paJDNmVMkHG9bn+XdIUFOE3m5T67gOa4vS3Y
6xM5W32Iat54hXMiANGvq1nFKhy9SsjpwtIILpZMXKoiUssEqSKcb/19dHq3iebPdNhQnInV4n3v
zWpqplbIPswf9B1sJowSh/tawhM8aWutoiHA/uOFmk9sKmrfUu87ThGTNzFQEXccRPBOylNFk9F5
rc3cTM9XbtMlksw8ek+kmlIVm+2NOSrUwMWXApah8yOHyjj+ZTBowy5cZG7w/foy1vKDidLerZbn
Cx7eY5obGNdDmbFUJlFN2OGQ22ZJEqAcvUP8TDz4GH+6U1604Ge4txAGvecaqMCey1YeU9fk9lUK
3zMnfNKs2ACDsbXZihWxoBJ7Bhwy2xHMBECcv8KVYT0bysl6ysKqpYLtG5Js//MhNBB1ReZG+Ka/
tL8RBqJOjp+SOf4mXXeWhiaRVVGgMpPoMW/xTpWBsj2GbTDvt5mcHEC82hQqgj8QXshdutyVVxvy
IwJLBkKry75VjZcy0xTEVOX5DuMxYL7ePv+EEXv/u7ss+sd6lr6s2CzpHYgp2KyoNXE7hAXzrSSk
UpuvJ0zeenz3RD5omrc22F7FFOdQoGV/pXUF5QKQNF/O3ep865+p9AtvUHOmVjH5VfwZx1HZbdSb
OzNBRvpfuiPhEHRLTaj0mBFQNcjPnusgtJmKp03ukGuyQi0zQrnxfHQxQbN6VvY+voBhWiOX0izP
lQSEUoLNZ7EckqunpcvjDOUzIsy0QLIrLfv82YL0fDqQzdXvZF1pGA3uTHS7YvcIqiCgmC9EMCa5
Q3BWaiuRS03GBgTESvIIn3uwoT2gK74s8E9HjRyxMoj6lUI7140ckA8dQwArtBHCC9DTiN+o5hJ1
2L4NaNxT3PIdRpiNF9KBTR16EL8KWCRKBnYr5y3wdXKdCEKeJZnVxChqUGYMfcJ8gfXdv0aLIoni
xyruhIprgHlF92MXVZb15/xBOstfP22DiiALqHjEKtddYbwSSjev9dNUJc4PIg41z1MQ2DxdPfUR
aLPyOStt+0Q2DfyCwlugeUk2BUEC452uAtbPys6YEWJUXbFKW/LgtagXJB7m+TcvCaNdYY9fNqiJ
r4dL+81iJ0/HBOGVQrYceaW0TpXqRJA+7TnG8Ml78AaUsgfJs/gH5zahPhuOT2oNvgNk2O4XMM6I
aUNIf1dUBywC9lhRNCtuGuRw46y6G++ezU09mI8l0dj+yHxPm+fsOPhT9o9cvBsUncy0fxAAjDAA
jk3CF7QaHqfg+JHbfNvDQjK0z12c0ZxpCcwOOfqeppFNxE3/lH4jgT/pvSaVDJyKwYSdNFVgbhFw
/uRtCigCaC/aE0IywDHemZpU4RQbdYVZDlwuRhdOEfys8vN4vcCBKxrXX57uec7FrQ3Rh6vuzdlp
fYoKoTrjqt4zwxfLWJVkYJZMRcQjy8/zmOKFCxcgzjmU59/k03WPvawd6nmG7KF42sLPwBme7nbl
GuB66jUnFMPNYm1heJE7HBL2lXChL9eisbaaP/CBWduGVvzMfpY3pIuMegFQntrrRPsCscJYMlUl
Smlx0/1UnvFzu81fOwx74X7NOMwOUjyfNR2ujNR59F/c+OWONeJxkxZ/+QJSap4l+GqPRbzmdbM3
a9xB3QzbLM55jcwZECPiQwwcE/LDX16T1x++iCxRtevpMAjJJ2egtmEEMlpTz1q/56KpJYiDZWrm
CYNyPxc/FccooMif1ozRlntjdfv6IOQX5bI4SH52+OFvuYQV3kFSmYrhscy/joxn0nnRldNaf91D
oYD30/eCIR2Rx39bMEVA7/lV9H1eiBVZhkM+0aOKXGKDYOE+9tgF4+37LmXBPIXQM5M8rBzPzDOq
cNs4efTG9o6cAlPKe1exzEkdP9lDvfKtJ1+u84HoLK+3RjIZnJlAVGPQEye/U/MyNzy23V/RJoWq
HitQKGitqmMmXOLbjZZq72OugFQLGu2AxE7CRVqe1VaZtTT/16WBpH3ICwuFS3eIYzxrppDW4j1L
4MskQuxU5JmUz9aaiuE+ugox+ThePLkoDZOcRZqjcQWvjyGhotXy/hUxHXfExJJYALfuJFvnoX/e
46VJPgKoPPJmSZmaeKhr4RbPMWTEWxOPSw4hqABtMy2h1Wp6NvfsQOI98R70V1NQxi6DBzsBxCY6
Vi8PmbuZDLy0HJc+5mdYFX5K4jGy7VaVuj00g8l64siLyWPFvpyAtznMosLt3+DY8Z8tu/E3LYiv
EbYqfrTg4fGw806clI5QGHFdEhJ0eNTRfBPpkGyMbGBSV6BeLfpq4Db9VVtgG27hfVZle5ZwzrDd
v6knpLHLN8khvG4hjhN0Xq8K86BDcWUKHNR+0urowaYY/d+zcCGoaZudtA+H0DrPOZHFhiuf62lP
Fd2N9jh7xcYj9WORgUpatBHpwmp9FMRqVLvHfDAlFlxSeCbcAQQx5NuoZ77AiLcSZgjBFfuUbM/w
u3Wkn2/k2bouXDnsLE7CVtYk+kkCJMrWZg/vLLYxGvxGKSt1TL64Aw6h/rFvoG/oKNv60zxV/Ka6
QPeFHsuIxpvtcxcO3VjRruaM0OBmErw8kP2ra/ZL4W8bi8YLCMWyEgV/BmXWA8VGvKhzgEYEOP/v
GgloSfMKmXBJoiwDntSdhaCG+f3I/LsouL5AwdbLbQb4noWKkKmPGjI5DIFM1v1yuhft6ldvFwW+
AX/J7VcXQUBtdEiINrinExNVHHfdvqc20X1JKOubF5j0fczagvKs/l1+wH8S112s/vuQ/KtG8M62
5wUoP0BljqIYcq+3U6bUQY1o5De7kgo49b7ShKNcJjS+QBXdqxHNoSeo4KCVjXO1KyNqv493udv6
VvQqz5hjyQI7yw8IB6slGQfr8LtI3QoMhCMFY9jP/Epky1avBOlWyDj5XxY2IGxQLLr+kqsEJbCJ
OEO9RkJ4jjDEmVfJaYbEifJM1kZYSU6sr2fNml72LG2LTF09MoyeSyDNPyIl1RM5wa27TP42WHHK
xsa0GcvZg4EU58OM1CPiL7vC/W0kCiYJpn61ypxwc+if+QzjuJ2sR79ZSr2HYWiQ3o21fj+lNA5W
8qH/KOUuFPh0SQ2B8dRtq+TS32G1rNyscKBXOiAsuj9zVDGplIYo5AHhZ/7fBU7CfYdPME81R5EK
7M9zO+9q325UOXMX1FYJK6IM/ZqLCs2Qom1Y6vY2ovtwgLedsieTUxsX69LE9PMTe5NbQNyBpjKj
KSZndSgNyJLbx0KOXFv3M6NHSIt8aMmo+IRC2ZWO1GV1CqCArWu77aVy6JwMebAufddWfc2Rr6I/
MI22cdiY6jnKbGEpwo7EpcrmO2I/gYrYSNKEAg7xrUGennzzKduW9i7EIBsWW/9Mtv79EIYkohR5
2CqZOsHReTUcyNoer06NsYvWxq9LY7DJD/g816crGPjmCYH9IDoBIKTNbXIpDwwZxbXYOn6xVZbI
WOZzsD2MdglsbfL1U1Rlanyu13oUWoeuBVQeSzDPx2R8QD5K9i0MDM6GjEY6Gzvk39wFucsgjtm6
IDo2iyzW4dNN1FguRoyZrirgOI+Duawahqbyo2JQ02f1n7o0nBwq2TKFkSEWv0HhmBj9MbtuoqJw
oVHFge9Ns6k45ZE6rBH9mQbS1R+eeFWZ+42T3tUVUrrVGyBuzNKGw9iJb1I6NVyxZmsvq4VAdAe+
LGa1mdi4Ovd7TPHQyXM0UUnNfx2nKz5a0nfc8LzayhrH/BJcvc/HqKXQ80uuDDvNiy3K4AYzL3VU
KO9Dq9Y/UMwflXTTS6/L1t36EbNDhVgZ88TtzuuE77AQTXXcvvv6z6ySjR7ZsP9d8r3JjIZrH1zt
YkA8cdAYsq7rZpaL+4n2YXvMlp1YaSyJVxTCvXvxO4AT1nSg3EDXEeiKBWBLp0jD5Gou2O7QT+vE
+xMxv+7JuIRQ3q0eFTyWr6asUslEw7Wm6t/qw+Qaez7DVMcozxEQx/bpDgQuchaxQexpXhO/vX/c
MLNem9z/UusiMpkDWqrQYmWsibaVMf/5hsalKWFF4eaxWJeJQmJYziK7Hpc2okoPIiPoB2GUQ0Z5
a1J4doMEZJINa0Rym+IoP57aOHoPLbUi6iiYXY26/AwsZI50nKtjQ/S5gBzG8d+QjTStvR4DGLR3
TLl7SvI9sEkR5molgI8FdnXWYDmXsVW+lEdrq7hsdOV/YyZiq5TbnQXOXWtUSy3YbIpy+8jrlhAT
paDYzETcnqPcVfgCKsdWaty6RlUjBXeX3b5lkZ+DNs2ozh/PrMkXJXhUqtTsTJbuKXuP+rWJZswT
Rp1bZOzCDg0+CvOnELPUGP4iYkPBqKaRJzvbfmJ4jssKD/NeBnYl6kcGySSXa4El36Etz5881/Pk
qU+s5oHnbhsceZBC5nJCG750+JaPQcBZCDrh4VS1nd4p8My+QzOsGZrLe7K7obcYO8v2fvTWooHS
9iv9Vy4eFU75B/ck0GYummnQoSIqcKgNi27nbxSBkHa/GQnHcCJevKGqnYYX4ip5REcLNhFNu8Vz
gyvVO5FZN28LRVYdju7dnROiP4U5viRJ5C38su4oEK6LOOdhQZY4ka/AqJJI6GAVFwBtFDbrrpEf
+x0TDv5xqjqSg5Adq3cX1c4eYa8Z8vP5KGjvnF2HWgS1ig2eZ359/u0DFRdwb2C9AJW43XUjPLT0
84Hwzmo1Vs6JCFQex8xj5qCk1feY0xpn4TMHACW5SPDgXcyWcpweV2UKjR9W0vysrJBk/fQ4nml6
dUSaqUxdL8QF+MW26tWsTJfU7L8ALf+FlmtO3JZ2ydCb+UdvBifCLl70HtbD9dMQC9q9eNeoBeME
FbiENbbGb0guHGvQP2BWUScKWLjUeo8e9G8J7hZeP2RGzXkED4e55T8RCZsF8AoaX9NhOEhqU+Pi
BCX/T71P9bLCthXH3H8i6/SlxstnslA2u2j+HDPWGT4aV1ok1UHcs3d6RHwk7P49xUyUgXzqCIEn
D7e5aantRDc0XfWkUzVm7lVXQh4x4LPZ8qSTxNcngbueeigG8fObQcoItlS3G4o85sLOWIB8kpta
watHS3zt26S9LCR+CiACxJQNg1uRKvy2wsC75Ie5dQu9wpAlSEXS/fyb92W/yCE3/LhqD4Hu9lAU
8icGQvrbsYTIwyKnva09McoAGarAPwqV3Z0qPJ/pbuqV9J/eopLF36JOQ9ZUa5gCBqjn3xHUNbJb
tCWuGROK9EAcIB2UzBcF9M9CN2utFR2tMTGky1J8OCt7Kn97zi7B3rJmoOKD/XYBTdBeBnbfYjCF
xCU9BRL9rF9lQ0DbMwUmx4WxzIKlFhIhaUpcEkNhgAm4qFX6SpADqtFXQrrD+CWDPNp5zzbsiv3m
7HOrwKHnqtmuTD9/+1jTCofsHfkkBjrNObXc38WgahCDk+GZcr9YgBjNTtC5rf0kiOQjBB+8lQIW
zKWvyBYdSPvSwpWtdztGrLTGDvEeI8KcMf3lmhsz63mqqqYphvjH7EUHTtnIJyI+U0mYHp+sq+jf
epOcuXzl3lnAF5qQQqmsr7gh42wJ4wBU3Uc5w0/QqVOCFYiS7bYr8EVqXZZ23zxP9OSvHWEqRMeW
+Ihn8+JNnphNNOcsNyVcKKGs0v2I/I//UVoQAkUKFWZOtwiahRLUeAAmjQdQM8FVGYKYNuA2Rvib
qZJiu496sX4CiMBKXXrj0loZeFgm8DyhEevupLQYMhCCNmgjQuGkxaJ2GxOdGYDnhmPOy5ozg4fZ
BNZcZ63SunaFCi4D5bFtDWBjJ3DLZECfyksa5y6mGULeYEFQMEhg7CD6xahJcNS11dAeGVbQ1T2c
J0koU5crds23KZhSaeUbDE3G/ys0EbsmLkhxfZcSV2VoqBtTuOUBNCfBYET1d6G0BwQUXN0LW4i2
iyJKLmEQcQpRpWA9l54Xfh66mfG30/OTtFgZu1j8w5s3Go6cxRhY8E/nD7jgMdf+gLLuKZY/i0Xt
z+EZH0kx+HfkMGzqYzNfnZys1JMMuzswUVjcvegr/MC1sNZmvGzxK7foCzerB1CmxQGE9LyZwOjS
F1ZiFmPr/2AEMsq1P6wqVr9PT0kZNyDDOVrlwmRMoV0ZUEouCq8E2IGPi9MZGDsnWp6qbUUaDlTr
YF4KCi70c2tIOC70KzDtxvArTREsHDinPZVku8kchAbSuPbHPEbfAbvzNEYbQOUa2pf6ktPstev2
OpRGRbn54uwmOwShqEhg2jV92bXBUeruLAfJAOMtmxhh7RwAe93sDk/pRocGiuqE75HKYsdjt28Y
esk+B/t/wp5gGnCHA6BpgBDjc02fc1rv8EXza1MzsaweC+2gouPnEHkLDaXtovjt0FJzhv5htNJi
Iph6514hYMM7tIOU/b0fVn2uzUXpfnqKjsx34qBiG6QeqNCeiXYT9HT6/KH2+o8qfpczne2UmSpp
CA11TkCO3BHg5HG6LnOGyQFC9uzzr3SgTC2jUh5c69M2pqZ5jJB3I3u2fI7SRmxE2SHRL34maAbi
Q7sh10IEjV8vPHUno5wdSD1gpmR0BKlbspcFaUTzhUYR7rl6WXfGaAoKQlqUWX0ngJwkOX3+9tL6
Gw0SsB1DpddBHqYS+RAzNauPlh55qwffo5eC0TnYqPlAo54BmrY7QN07q7rC0r77y24ec9O5V6Af
VinmI8SZ/N5Dx23jOp7YlhYLy3OQLzG3t18nPlZ/UsI/8ilNkeVl1VCS2e0klBu/wAe5DAd1tV0C
xZ9dg2CWT8pu3N0OG6O5OSvDyX5j9LasepEauC21ji7TBhyAyss0rl4zU4apxJpPMNXf5fB9xJUR
qPv1xp3w6W2vaPV83g+I1nqb0SJq0z+rvd1/t0AQDuxi6gzCoSn9tkDOEqD91Kx5qAbFCK0LvqHr
Mgbfq5XncighRex5PEswT03bwiE7rm+m9tWEIUKyiPAwJ23IM6Eefnp9Ci/D82qlvjPDHHGGnBiA
F9As3MoXrEUARa2lrp0rVrTr+ZoEtMLHDfOKJP9f3rQvt7F65kq7G5lpa8d2gtaDgta5j47S2LmQ
/ETRh396NB9FpxawBZn0+GucMeDa9uvFWsTSOcMg8NxEu6Ck+jNrCujT6ktgyzFkrRE2TX0khD3j
JlCOLKeBj9RXL6HYkqziAd7FB8iev72ZLMIuC1TKAJL5MU/yynElE+/v4/Mprjb5AAFFsn6OiTFU
NtOSbVVt7z2qvMkKJ0FOiSA/YXyGqDP3kPNGmYClHjAfXFMZr2v9cW1ieAfpuY/2OvCxy3sPA3Qy
3dlXC98rVTdOFwgZVT9i/yRnHlHAbZM25mWzBV1wnQ3j5hJ45Q9CYES19SGLXJjD2sMUFFC+e0si
kGcbK6yuYNJprwGWeaoN8MR5xqHWw+UGzH0ZHgWpuUABi13Q1TlXnonxB1ZgMoeWLEKKDGJQ+CpV
uFXrAzG3l5nYsdhjJ4b1ncZq6oKnmFHAGXuvYJOfSVDS9mD/ANPZG/IXzoSU0JwW5Ht0dBkRRnyF
Mb1o0M4tQE0S8R7XG+VXsbQj5w2Mv1BgJoaaUVznacz7wBQ0SUTGmUk/yIEA0l+15SXR+29iooZO
WHxqB9ndh5x8N1X9BUqBqflDCNHM6yYCGRHvQRirUWWmxWMHQSa7lSkk356MDf9zh0ZV+NZu8yjb
fb4kDeS+tqn8wDpERxkq5D9SQT9nQTmqrPI0za2eFc6Xu47gaAofSgVpyWGOD6EamWy99wCrpcND
mSeGUS5nBz85WVrDCTQYfRut0fbMOSUsw0n0gpocjIyJrIGa5Zk4lWrcqCawzLtwubJUCRvE9tPh
lGZsd2NeryHYIr6VTAwuCATcUZOlbpbQaaXZXq6/SAIt7UD6qoG1OFbebC2Njc7BcfggxE9x7AZW
OhTbI0GkwixOGwSpiEoC5ygMyatr9mItnxoG9X6n31fPm0C3EBzqVyNRX4LCUxgFg28gSfTS4pAN
6efzcOjXLaW3t2vPk7HlWO/tWtuquF8UFtUooqK3CxyAq7YuV2tvF30kfrdi3DcmmRMhKSyOh4cC
rx61PL7LPw4SRKdhKYepxCXQpikydqKi0MSErHPb+dehqgAJTNOKuFzOOivOseLVXI9OkV/VtQBE
0EFv0AaJMypfODvUec/naP1Cf6ZfIbPrJ59bYny6VpH90pkABA3/jifiRjzLbaCXNk2XAa5cvtPK
WEAoOTHpkkWcj1jgJcH5VcoLf1O5tla8Hr0Ypmap5dD4mn09uSA9LdJauwQ1SernNAUoWx8/SzA9
6OwguM2hfzneM8mJ0mMgC3ts+5NauD6vTdyVIWWrZ+W7Srv3NVwlTrzIy5+QL2Ek2+UiagOCT4z4
7JxAJzTLhJQPfaMTPkjzAVf8qiep0+1CwAgMl25AuN7ZU3Qnwjrr7BNug2XB2aOCin0YxCVJACA5
0BeLDLaxwK/aEoIU7oLqKFmJSdU/64VSg1HbSPr60XQnaF+3f6PuqtVtry/662NghXSxIWEJw9MC
wmy/UMvgDVCsLOFb3mnU3RfNgHQEC4TR6vk0GY79QCcnB78XDwtlTHkKjkgp6AR3FR6eav315eyT
zRnvLuO8MKdT3vjrfZ9fZtEzVGXQNJKmI0rympPyziOTD+BrlzhTtOLrL7+lsr/za7sG8jbVwn+6
N8RdC4ORYSwa3oiM08Uyzu+5kHnNGymuGUx6bon9upyrd0LmC7se9opj6XkKRehrHyjnkRwXHnby
dpvxLm3TE1oQRKEjlMOgYoBNQv7toQn10ydgsdGvA841ER9HrJJPIDfIbTcPZJdbiYPW1/pVYtl4
VT6e3xxojovPmmqNT5CpuicftJkcNtzg6HJtkFRGqTF0GveFGeKjNdtHEPKZRkMaAkJrni839B+u
febFF4Y6Hr6vop7XQj/M3dEkaVvQ4nFeocxR7bsvaETL5tUZSwcB4foir8DmDThTKf1v7TDFgRqY
no9QBVJWmyPsb/B4J83cthB8gtlJvAWoZL8I8+zao54wEWZ4MKar0szWBs/M5xzIWju/6J9sMdRi
iShZDYTwzXe1W22Yp+4BfUJvSkEcxsPxhRzmHDZj27mWmhAwmoPXv828Vg/vIiNpAfwB5Moc1zWZ
7YnOofbPylVAkOsGyzy3dJ6L3RUPw6aHCoxU3mApPYoeGSE7Os75OxEZnZVR+EUJ2q+L+YXK1UUA
HfnUk68FbXefld7WVhA/D9djt02ziyJrOQP40sgyVcsc7sibE2RUNjJFNctX0ZV98hBAZv8iSbld
WMgk5ey1JRtklHM3/Wj7AnlXBnbOqDxwqpQWS4rIg5ROEqd+7XLKYw697s8MUdQgV1MySrLpmVNY
uIEKIWpxz96ZVP3mDyiV+F3jjEHm9lFtO3kTE67C5v64KdKgIFwsDDs0KlIh35KRsJerRC/oRzt2
PxW0ldhuqWzWP2VY+Gm3cgo1fFNfTvjnDh+I7JaJzFcryVsGWUn2viQdZ+uF8ixFYSFMg4s4TPwZ
BXJYXIDGP6elnnySjGKPEazFQVmA8ssNeMEgAoRWqmn7ATiTO/wtBDFcuAKKVgMGECu9KKDSO6aC
5Z8O9zJIEKN3G/yaYwYoD20LwX+Phg2nuI8/W3/MMemdWp0totxo4lr+mXy6vsCK4hHjoqr2+1I3
Ghvhmk53nVFE57hIuZTgQ5cx+XuIej/rdP+t3HDE6a2tgdmP+sFd/FuLaAJJN5jlk5QQXGMJvFRl
u2FR1VcDabNHFauMvtsZ5f79gqz4l3nebJgexvfaMhttvU3hPMycTcpDcHgKGOsvUoggJ4thi6+w
P39+e4AoMrHyHlh+cog0tOslAmT26amdMS3BMzr1jk+ZNZt3oWrJHkWse7+SiVIyTbkqXKaVvLrJ
LcUlKUM77ib4NyXTeLtQtBhI3gewXDAL1tNL0WKmVvaNsosgwSRSSzcUNZjAQqol16YVTORfv+aG
WKt/hAvzHt3VeDdNseBKWSG+MDK0k82YeTQ27oi7Av+KDpimLMihaRtljg4XFubLQ/l4XxxWXJdP
qVyvNafFd+Vl5hFmAF6wIgm8s166KTchmKngcwSaPLBAYSZhVh37dsNTA8Zm8tBf1w6sjVWcDGfF
MnL4yA6frWY+6/GM0rrnA6qLruwuKlWQOkE4D1l7zch3suL4/pH8s8oIKyLOxK+IfYApY1BcbJFr
W4WRR0VWWKgiksCKtg65zBFjc+m/tAATZerLNN6qZaipOAgUiR948EtBNz6j3uWqOPdzymHoop62
tzerDEDj56mbXIzvcMhH+YKB3X+rO59xo3A90ltNnEn2SogB7o4afzsCCXo5tmxqo8w7efBV21YH
DPI6jOTT2cfiYhiNcQYk1RP6/UrfvFE5zi7oDWMSie7n68IMBCeFom/yVtA8mYDDOlkeadkZtW0k
WmuN8vhA2Ipqds53OCscjTtCx0ZuGjYsvUq/XwmwuuoFlCaT3MsriIyyyAE6VsBviKK13rRbEe0c
sq0gxwgZMKl/YCZbVQ102IgpvboPIomyIwaArjZcLR544SJIv11C8Jf3KQioqDvmALUpfwJjkb22
g6Qssje4MHUWJbmNVMur1ScVMeeU0/fmGlkS9kgD6FJiLGlqt6+VmtQycaraq4OR4M9/PM1bLjq1
82cuvgyIbq/MSxAbPcJN3bJmXc5p+C0PxZDmx7PaoYqxsa/RXv3zo/Y5nblLJ2aiMiByqeIR7NKl
GUCQ3sUW0tRm6TXLNDwS/F0pirq3H3hqO4QnTa0F6z3fN2U6x1RPnPfRqt5ba4GD4J1DTzNTH5o1
Dtfb/LQ966Z1ceoaJBtKYGez+v0w4K+MLCaXTF0uB4FgosioGpbcGydv4BDUf1mKosn2IFkM1Ovb
Aqi4fSBFCqNF4hItnx4xHdU8/ut+yxPckid4g9E7+7aPexktMzvD+cjb/pXx22853CsOR9TF2hTc
MBYpQqUFpKYH7BlDxYXH6grqGaFMfML5enWYtIgellpIDq8xiWBL8MDkQ7sxQkqUh8sX+CNYdTns
LmhqQzzn55YrnIF1q3gChX8P+VFBZVDKW5uy3S0Lm1JtUs0QD1NBlorKMv30+0/zlh8K7LKmUQ3t
/YlU7kxX0TTiFQkTNUKXJp7c8F6ZntEG54MprA4UMsgjsicA7C+4ZWXxEAcYykOicm0eu/VyaShl
cH6NRajEJ0Y2ESbEDm0RBc+T5jYl7OkYsXnMeY/sVLxEaYO6ciCBhJ/vxu9WSDo4qjfMLoTM6wCD
HmfK1ZPsmDSaabrYsdh0Q57UdjVCbrm0dXdmHMQJA62pTAYYi05GsED92UrW1hvYcEZmCBCsGVod
BZbP40wDiWHOWZhEqmkfWwMXGYaMaqb2BGY23UShF5ZPmKeH+uwQxlULLcprmqoXedrdPmdevVgZ
X1vZUE28tTjeYiiJK/Yps0t7QSLjFhIeK4Ir3Az3035tCt7PGGNbmPMG/sWG4jk6N0wSAi/8VTbP
34DyRoewBFe7C8MnbYVlvmHbX4bAZ7EEbS0GXjOhIp/Z7fRHcduZqDVILJSsK3vWg8Mdqm3nCpw3
AXa+1r07EJiKAxQGF7pJM7kUVBsrkjEZ1Y4SXOKx7O/6vApHDh2PWHQkF6ck7M2AhzE0H0CkZJEd
+XHWRoLsdLtZHrqGHtuZhYy0o0vPnW086Rgj4zBwAfoUgpoDvhaTA29SB+JspoOT3PrVY+W+tjXB
SnRr9koE1L6MLfA7WDFLJU8/WSUdA8MIv+6g/ADJUxYFS9dKZ07B946KkSqu7F3LoMGjFxtBflg9
y4JLPJoWEbr3Oe6T4szpv7rZiKhwCoNav9aLPGf5+igR/pYUxDbkD5QzaMCVK086O8qBW3v/wdAp
zyb90o4Joh1ey5N4GCM/WE998/su6zZr4iATApBw6t1uEm13Rvsswht7t/ddR76EGfqZ3OldAaWi
5FX3rAhOIUWGvF3XAokBMNek3Hh06qBYvq54eMcC+svTzvjfEJ9r3D2S8jPEGqYh5giKeJlV2gXo
F6ZID1nV8USZiWzK2/JDvkqaFnH02uKpPC2uYx/yyTGPfubtwOlIP5ImveAF0BMlibXXWts1Z2x9
P+foB5sK/z3DzMocmU8UPnmMdyPY1KnowumdygBgm5NT4TXdFhDjGLqJgRf7mSWUmdoT9UiktAwz
4hIOFUR8HFtvXNZ/Ghl3IEAkEvUxIoSdU4wIRfSrhDy5H4bpZ5ZPtWOk9QmDxGCeegdlZB68Krre
5Ipa9zgUwhkpzisA+79Y2QlLYPrB7j/bBZ69XtkyQlKufPcEa9g8Rn1GItqxuEKoUJnO2EPttU3k
6NQh3H0XNOf62v0sVA6GTZhIKKMFAFSW5qSC/QjiVSGdYL/XbBzRqfkj6x6O6nr9UNr4RLwkKz74
rLsAF5EnPuIrnTv2cblrd616/a5n/xKQxWFunoLH442SeIx+dOVQwy4hQxYaJfBhD/Iq0uRB2sop
UkIJhdJpB1we3TPoX86k0BKlGvQXvPgSW3omKoIopLLIRmjaArN3leh8tqFIVsDMaDti5L2pW195
nkp473/JmRnT3NnxNpBQ2Y4dXjdd4lt57p8CR6o5oFChZurEz/k2GcZsnC8pFfDCVAu4CPSWd1A8
O+zFO6Z8F5v8jY25I7luRPwrJLWWXCLebfN3u8omlCRJ5kblFdxzWDv3LHJRXLG0SEIZTrMIEOlH
mLdWC4w45LMKGauZ/mJ9u52ZEPnOOz0O46TKWew1oh2V+OkvGGFn+621q13OUUfCe2YIhlPRXxTt
NEH80YRurWjtGT1CsPMXlOgFgHUdcIOQV0VaF0Lvj+FCwOmG73g1TGaV7E7WQncQrCrGNflPL91d
Uc3EN3ItXADPzhRnGr5HcMtd2iZ8ME/155byEDojtbOvDIvNe2lYboXT5n6DsO4jE311BUl+1ClN
AYqGkE/5LFeeVjkB6qQhR+tHKlhw9UtQHXSR9EpbCMv0vy9PpeIVteVpBC6509FnXkWlCQylPQ4w
+T3sNC/K5oAnQ0QK8lUAn21diM4PZGhjfqgZ4rVDap8VsQHzwIRn9jytNZrdDEeqWsmTp1WTa9xk
3nYADGyL3adl9s7OfbnnXMzHPZX5+2z5rzsxozjB8GUbYtmpHUvZngWEgRH5ge9I1AisPmFPxcjM
nkjvRmrWv+YTkwWsKKjOgU+OBP7d0QWuUwMKHr5SBKUZnEnTS5h19STsSN83omrwLFi8JIJo/z3P
LprLPeJJ8FKgURwrFpEJc3i3MfzQFKvIIrOXO4ZuK9eU8g6rk4xzQ3vwZHNDZAuxsrPkHcRNWetT
7GntOuX67g1VK0ksYpS2VcXKVzugcrAA+9XhXWea5Npm8vwk8afcF/E6AluP0CL4WqWA5T6jNLfC
rg9HppwiKkBlj/C3Z6i0/SwNI00D4EbwVyOdTsrx69sX1VKCy85/TOzGU2VQxa0tvf6w785BW4i6
LAdBDIN6CeD3Ao64blY9+dZ30onlz/zpVEZ+PH/6BWScThHuVUMKhj1bZyBcuG/fSDK0Zhz4uPxf
dOdOjcjytXmTy7n2HEBFjTQ6IAeY4ae1MAEfHllM1An1dFG5prire+KQwb2zMsFCFAEaB12/rfto
tpfTJBm+ICwdkTvGLI59z78R4uhAfA8z9fboTF7agvsdLTg5D5F0ZaYIySuZU3tGcQezSSi7L+Uq
KmZnxrwliBxXWXJGtF2QDmcEEGsLW49P5xbOxAAurLqa0BW5clQEDFAbjYVSDQeWPyWQyLS8BqnM
HmJyMFwWotJofCP85RkC8Cub6yEfHhoVCQjAnq69CYhrES0iLHieiUNWTjxQTgOFw4RYmd+fXqKK
xRnhoxQgbpJ2RhTvhiG5TtioWw+zIB4o449oRG8B3e0KGdbxm+HSR6XtaJUHtv3FXjNR322r9Eu3
/BwOtYVO7lVjVKEnxuKoHqXLxQWgtLn2LHpZynY/RAZ+ZJiVYbp7RbTjFsQ0tF3X73L0w2yAcCbG
7SrKCmivkHKyi3lt4PakDFUhDDQWvSzJxKJD3jM/DKCogbJhxOntNQWETziKOBmO6QO1QXAN6/pK
faSBrJtLKo0wCu/uvcAyqF9s93oMYMr2K98Ewgl8Dqg7uQYpHrX2+TF/uI/GOUvkeM+eKw2hJLqi
VchaBzWDPTneODGgZ1THuRto5t0HW7YBVdXdgNbovePgRVoolZzyG9J99D11yHHDuZQ15srenLIs
1vB9pVsaNPwvZeAxfuUf/pTD58kyW0ny8pEbLcM/T7PPVhv7a3Cg5THv8XPW040x/TUxCt8IW78M
ACEsba3RE6eC4GpH70iXAwRNrJUk2qWoP5qfZ68VMfiTvj9dVaQhk2uH6PFKQteOLMyvbin6RxEM
6OW6CENTODBeG2G5T+5SEGXC+4T3htqu343J1MvLkLZ1SXH9B8ZTyWh385eFMkB1Cvds3I+Xb/NF
jb46WljcF5x2oKCqfM2/tBEYAyP3RL7fFyf6vLQPmFu/QmTKEl9hBiBDYGKeAIrSycBcFk2+AGWM
iIlt2NAnjd3qw4OBkIg+VRLzVqfJJ42eSJmjdO4YajK/TdtNDJIXU4nzVvUxAJbJUv40MBeuZnBw
jrAYZLXXBruug7BSVTaaOYK211L5f5eDiWfjEfqdfdBa9HvxfECdbWi7aK4xZrnujq3oUfA9TakZ
36zTTVW6jNJDo+xjeKgMNLLSH6kZ2qPw7ZK00H/h6rrQpLXyoNxYF1r3+xUVDwGEAOMbUKaOCm79
6BB7VboDJxKI2LMDXWMRilFe1a1uw6F5DKsSk/nSljP3V/R0LJjs/PjMp0jaDasXCDDu74gzXXf+
YQYiF4/KY5oZaGSemNF8HN2BBWPJf/VGseX6HO0OuREunBY9ncS3h/KVKY8/P9BQsFwaREiRnecJ
H9P0iSwSqMZyzSDefhM8wKCzt1G59WE2g7CUJCq3CtBeppOsqemiCfPFPAQuWjncBBWWoP71tbKo
pDVhmGc1IbkmhEcDcWSphunnNVlLqbLOkY4Zq941mrpHpqUpCJvyqTa4BISJRTFCbNCyQr2sm8Zt
70oAZmHLURqydfVurZ1+1FYzTI2n+N1VfjPnY/FJkB/2g9flX4wqNmtxWc4CUZ8MYargkMapIHxv
SGCwuZ25r8Q6blDG/TGGEFDCUL8ls1VrrJ+re4b4rkeN9AuSbitMKf7ULq/CfwD24FRusGLWGGsB
bPhgYjfSXOLo9oRFCRvVN9D711tfkts5ycJwWTNlTX+41jzx3L6iTKngbaHlKGnf48MZATM/bzfr
JYsybnNEbGikCTaiEPb70oa0P7q1eeGocFJ/lcwB6jv1PosbIANyFXo9+HUtpyzlzBTcyzG/toZc
JWjC2bapLA2g2cKcJembAEcHCeQdANF7lAQY8sHyCUgVkydCzU8O9ivgqnEao5pqSOMiDu4x2i/O
ZEbWaoMfMDX6WRXUMc67x3P8kFToe1TNcJcEJe8WwTlIs4VhYIriw7khgyG0dU6JPtWkFEkRTjst
n/zz2G+ilvbN7kqFEoW+esvpHKZnxKBW3ZFD7/Dg8lp7JedJw3RzwhnxuyZb5MC++XXRTbIro31s
BxWo1AN5UngMyYp1YQZaiLUs9EqgIo3loDZ/q1rT7pvOvQVUF/jPmkB/m/bX71ixbQuADWF409sY
KiUzLrQzmceHajuaKmoAgJCkKXVnW9Ws5xHKbtaPgsM4w9KQMcGYSOuEOW3WFWF6OXOtQWzuUV8Y
AZK7cMRHc+eQlq9QRHycWRjXN2Ek+6cJvnc56VdGgLyE0Ejaj6XqMOxJJMuJ1KRdAO9jPQO2v9aY
9wgDO+YPQQGZikNm/ihQXvQzBqboFgQ7vq4iRO6xVxokB56FQZ4tszSsxPXPoradvTNiMeqycsmv
FUFP4ps+RrsGMYSlULThzxj+5bL2PPaS/Ffnb8UugItz8KPxWFQzA4RjFhQZY4FBJlY4av6oJONe
6FbdSP1DdsjmwQbLzfFWdgyrNUQ5gQb3gVCktZG8RqdNZ3AR4zFwYtBNSoWFIsWbfSe3tpzK/hDD
Qc+NvdFMw1jLxmbtZjmb2ix7MzRnq8EHT9GIBT63Yw63zKjeN21RY5aw426BvYg67osoXmF/fE0U
E7kWkIlsvn9vvighGBvhQxtPnEcpxSvJTd15IgYr/skoro23yiHa5ZJ/3uJbA8ZTPAiqo3lCAhL+
/jHov7BRp53zbKqtLwxuiUNiaIXxwIy+0Jmm/I4YcqzbdcD3czBN3qgB6E+WCj1cSYz8RuKn5auC
Li08hRvxpyluzmhTpMAGZ+955PIYJpdEHs2Lq/+egNDjB6MWfRX/zwrCqE6BpyzLQ1OTRk3euGSR
ErdRUDj/KEviLuIZ40bKQ4EP+g5nWp5oHgcX9FZchqiW004U1/rev1RhzWcLU6PsdZiaXlEmpeDI
aY4GII1ICkMcpDNmmGS/fp2FvN56ANYdaKLDXjeTVa5oWzOefTNMMqU7o28WcDrxRgXsYLOkmUUC
RoPjbmVpc2SCTehaT1ptSDEC5tfteh5QBLixMSx0126dKgVBd62Q52jGhLWcwJXrSbdbqOj1ssRc
1fozkFy4v7VwhGiUUusIP3woWfXPun5va7G9nWqBjndIUiJdl1LWnAXlwpico8sRAQE9r1s3gcCT
sVXaFdsHMpADe+U/Ru23Wi/mcQMggcDiqGbEaMuWAMNGEN9SlDiQmrK4hxGVPyDmgl8/byD6ED7z
8MdhQNmjOoJKamk60WMX22kU0A4ullFy+ge6etvaP59pf7fW+04Sjmj6akBp6jVd9/SDxqbMVayw
jiQj5ut06YQ5YVXuZRw0dRmaRPLZcdSg7CB6hnk9KloNX2EhU9zllTGP6wxQcJn9Um/EjPB6Gf+M
vylpal6yez+9iIAbwkkbnhC1Q3Mfy//eHny8mtNFAVGZ8Yecd0GoNzgnAHsx7EsNQN7CuCNw/fzi
b2+6owCJLpF0msGhL4KzdMEO6rCOAxyFdOdTL+2zn9u6xaipa1ahwtXy9vEz3ydGX5OmAMbZJzbC
Ba0oiO/WFdXBkZ2TnQZwkyDox02OIC8s12TmwYPWS3vg90c5ciaO34v+8iEQDsQgP/Jlknc6BUKT
gnH8Uw3J7zciiloitj8YWSUWhUfWX/wap+bQUZvVcVkiTOc32KVpnVR7tqwyFGXh3pTKdb3Tgq2B
KttXPvKcg6U1jZsljARpKnTOFRTKALq83ygazg0lExfgdO51nN30eik3bD7LpZihy/cFVhEJuPWi
RJYT51pGAOrmamYwZ7znHjM4LaVnJTx0jG+af2+oOzuS78L7vvJru6gUVW8sFkbDGuEVFabgoG1D
EmOgKcX0IE+sXd8ICjcd7vIBohkd5QmNWp7GOrpcHsD2IG0NHcKIX1+MCwOyWrlBJgfTKK9lzdME
J1m5LLzITnGMlr7Z9n8MHhV7Q3T0aoZbzfxiSxAFpqVbFsFkkW7ezTcmhEGT/E1Ycusq/HLdG8WL
nSae0gXQyKd6Y8Px5kRkv8U2mToZFpgkNyJ+pPnitnKOmnJbsnVONQ++EeeFxylM0/CWZn5s9Kfx
YoM0H6wi/XJpYBlBtE2SvoBmNJi4x89Xuadik6Gg1zLVvoFvpPE7hK9lPjZ0cd51pyeQuft9c7GP
zFgy+EChnA14IkSLID1drjxjhy5ppU1NEJIfYu5g4D/0EO2Xm3/MKEIam/trhqD9KKCEXAON+U8w
PxG8BQ3maIXUruJFoW/n4htY4KX3L2IktGcE0TPeKakjPEtc/xU/OctEJOpi7nNYzVwG9LJBkoHn
tt6C/R189u916wM7nSWHlwcVwc/jYe74tN/8QZ+FZNR7KeABsXMsH99J6GqGkhkltdZjOnezizmV
l2jMb8I1qIRBP809+4NOJpBolGCVlxlIg3gf5KIOf5aDND2KdKTjTxU3TtOBRnmCkYMwu65Hexre
j/Ic+AVqQHtgJ7/M9lJu0gUv6Y7E7dpjz+v9BdWx81BiveYbdGq5zGGk6ma7LpkBAedgaZSyG/ka
+6kDnM9hF7nsI8F7iYDBGn26SQ0sMQdrhTgp2d4HzhJb2rpcRmxZxmCIHigjSA2KjU62ueSDPvuC
ZhW/VWcfmnEFoioRgco7kxLEJVl875PPxpeAqhb3svSAWSqcaHg25hsoVc2EYGo9KhGENO8hbHA1
3GvV1dYzFAFILrCKmhN2+68yTSV8jROBZt3YXsgyZgZrrp1Dpt0JHd7s2U6E1lZqbGtD+sGUDv5Q
hOIWOblfc9dFQhEx1vuzSBrGOsTmOUTr+DMXt3TfEfIYs9Lk7z7FIz2BateO7PKyqSMIf6jD07n+
3Ppho06Xb7A0CpD+DyjJdGsYVgJoNf9j/iNdqsl2jlVVSiIEP04sm9QX/ZeOWd6GN07c6511sGlq
Rhr2ShpprMzHH6RZKonqiym3F9IMejI3x+xl9/2JOWgt0eAGYA1vFbfgp09t8aj5wUex8ARu8iV3
/djwMHebgMHiA8PXNdOTFi9h9X1RtcMsYEGhzHsfjY47iZL+sSwDZyeEDLTbu2UcB6muhh9JKVj0
36hRRNhNXZmR9e3EqF4To36zjhf0hgR8pfj+AklOyt4IYJ96sq+ODSa+8SPZHc0lL2JWNx5iZBPK
jLs/MI4n53UTR0hhbViiMJzsAwPO9CxRxIiWWBz++HkFbldFM5lnHoQA1yDHlIE3dnBwCeoEr2uK
wB6DeijXNFU/t/pVSgHuMBA76Rz6NCcXJjcCbYnrqP4xPwuy86BC8aARSY7RlCiIY/WXdP1UDb9U
jKbduObslVPPjcwuXMhNTHuy6H/XPISWdzt8l+YuERKwTZEjyB9Hx5eO2cGCp8rg7EsFrPFtOoOp
Hgx4DRrIV2FZEdY531PqDHS7ot/bQo8e4ktS25qLSHfbUfuO2pLLzucNPttKq1gYJtKj48enjTds
9DVjeP5b8yXr5gGxVlPm4EVZgop5RY5QIL7JVzQUcdUrQOUarTFXcEgiDKF0fUHIH4shcWUMMQQN
UqmWTHzsOfxbwEIAlW8B5ej88GXcht7AsHptXOF0Qv2ceYHbP6VqjMqPnRhHl13Jy3xYin0hiuuv
UymYkgjFMrXexmUyhi0tq3IJz2BPI5nzBP2p6VdW4nnQCbLF97F0u2LSgdU9yqiHI61gvO/6eS0R
I9xP63ca68kyTbPVik31fOuRNOBJn2u/ulU9QQT8XUlDagv9Yxi98s4sg1CsL8Z9TTyBiasp9XDN
ob6Qcj3sghLSlsZ8tYaoH3mqDewTAVDayFjq9QA1RrwIGrCsHKL6q7/KLNIIADiOYimrsCSFIG59
nAsm5FwgQ/e9dLBgTJqXaT7Ku3cO1WJhdSaCnkK7ZE7CDul3gputF8hRx/xxZKEfShbzSiv73vkS
fd3v8YHIyRnGrz0OPDAfJ3SH/8MMHa5Wy7Kdjq46NY3cPk1mHXKheQZDSXkv2HWpfwuheQd3aNDG
6cVOue50vfASz+8z5/RVG443kPLa9w+SRS0P9+pKEVj/12xmf0Oy+9zz/q9JaV3q1bG/AOvl0pqA
7+/Yez4hG89c2nni+K4Ly0lrMv2bh2t+0r2USD8nLxSREs9Xp/OYTnhpbtVhpdmYSg42ehMe+Hww
mPNK2aVibCFIYReOkDf1zOKewuIBRKcem0GVjXt1aUMwjFdtcqyPY07WnIRs8Lsx/GPgtwTcRexr
Ab/dei39hHO63VsBxUvq7n032PXtjYvBayDyiIK4p1N4TXz6jzhKjZ/IlBIy29IyF7qOlZ6ygZeP
rNettGupOWbecQGTNL5Mvxg0YneJoSJSvPnM+7NZZL6orEXmfnsQY2V7gkVYOGY34pFMnvamuWhE
UHdBctejCDb3KPIwbDccqPIUg/XUfJ1kFZ6xfRzrgQOyngsYCvASdWZRLTohpey4QTfQu4Gudik1
f7CnZ+n2pmuHtR+nmKbGSmD4d2X31CDRfnWaFHdp8BcWPEyTtBedvyvr7Je4cAhTjaIAVzZyFpQw
EzDSLB1ujcZnVJ3w2pWfMcz7weaW3jTpmQEuZ8ElzpT13ByqM7fKvhAALFafOCUddD7sVFsW9l++
RDvd+JEZ/sJakZe0MlVnETmLA02zWir9T1uAkxncpOWxPJHszLQD/tDbL12fjFsab/WQV/B+ranJ
sMxC/wh9BbGf6Ncp3EXFWTJKNEhhsBhs9cK4DmJwODh+vXzQDz1ybTYKmQ+Zh9kOgafzV9ziYUv8
buA7vsC2HpCA1dvz/pvIWYZ7oq+dCPIDIo+I+OoWE9Na1bLDDjDqX7uuaj/GMeQTX3laSSlLEmW+
zSNgEFEGUXAKDoFOE0pJ7NiJqzeHkaJ6s6TBEDb5S+grGFwM/b+rr8jghthsdQzZRKLjeJ3Ivs/G
HvKalF+xp09I7ZPPFZ9mYd36BadOb4WgBsypFHQrW7I0FadDoe52Wbk/kGqoCsF46w3NhDmDZiPJ
Lc/Bz8f19rAODkDb90URDePljb1iVnUD4crCTj0RMSXaum2TxEQsjZNZm+BGGXF+mnG9/AR+7ckS
QaLzRhH61P6AQ6eXnnkj6XqnhKZmNHTBmRU91Zhl8SZazeKECzifShwWyfWxsl2w1TY1tS1xJ1er
P9E9E+8OKIRF38D9KNMsN0awdHmifvvmcx6NDR5//SsUVNQhsT6rO7fpZpAcg4pVlrvXsY1a+xxd
QkY6pMV1krIWGlWAwO918Qx8cRyquWjrO+BY4KIKE/daKamB+CwroklY7F50C+G3qfQS5zEyot3G
flJ5aCztAhafPWg+i6oQXEuKePmKhUhOYeUxmt/qT4rShH9CMQzE4uUja5IoUpHpv2swpv+1DC26
qg0=
`protect end_protected
