-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1wqrLqH/9iz/zNV7MC/nFZ9yaaTIbqz9tsMYgRJfY328+8uWhVGduLbk3KWAJLhMNsabseX42Bnw
ATXSO13OwxE3fBIO/moUiTLaxfKOsmryySmRmxypqMgfzmLYOigDncbyFl0V9cDBt2GuGMrojYr2
ffbstH6xUm9tF1wQxQJWJc2Iw3UjYJD8Sw0TdcVWyQ+BCNpP+GFI0JUswWGDYEEijfZxB57ZPh2i
ZboJWNVmFH83j9Ub5SOIQQw801qhL0q4HGF7G40tBdaP5KmNsymgsWUjXxEJMwOcQz26WbuuEFVk
7m1Zn+wH1inMdNMgi8lvlAReB0rshq/NhaLghQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
CydTXTyG1e5fmMaFlBu7RkUXjfKnhYZ3iKRFtaNedELzcUtPDn4AfAmy9vgPRQ2fwGMFrshrnjOn
B6iPMbub9e3xtu46MxyOR41CZ1ZUh9I8ntbmK4G+V1zWXfJAacCiUzrp72vtMhr2vlyCj/VKMcUu
BuYFXets6sbsBp1KIfs+EXunTEZIfEeHs8cTP1akfP33X+TK3t7//2J4Hsyp/GUbqDfDP4erzyID
5KfPWhZf+opExYlowUCFmnReIfHPr7lrauJs7AeFQ+HklyO+PoPeYWKvk8ARTyqMIlpWpRaDKfRe
QU0ynTs8ElPAXC4hf4at6FMIonk5XsP7SHLIzSGLipXgBVCnTAoqz5lwYDwO9Tv3Io4ndKGDE/ND
AD4O0vazux2cEcYcT7/H3YqHFW2BCLF3v5eNhwCKSG/PNgzm6EBojJM8lRCfO7RhSvZpv7LtWkhu
oifpx4L0/hOLm/sG2uo+uEhLzpRlE9G1qBBvLsOsVNPSCpb4SoYVgyAzceOUV3VJlUacy+JiXx+o
CUBufz5OtWRqHwN9dwYgMVq+E3IBjb0KAGI6vRxAjUvEM+MMZOStn2tJp7WUYsgoDSdymCnnmcmG
+VS2HKkKb9FWMJH4CSB13AEPGVZb4LWXEXM6kvWFixAzJUjzg2F8Lb4iVMFQZhu1mutiD2pvApbw
uyrjhiqFMM7smFnj7pdbOECzVbOqUFZNpO8ExUmbpkX4+aHX2KzjJIRBv1JXenVZrUX0g3n/gv4D
Kom6TDDLHKOGtSYmL51kR+T7+oFKC0cUJxce92mGT8DWZjtYwZKWnVWUOKvCv5j6dLgPuNX9/5Vr
dr4Axxmk/zPqNme5wddE5/+I2Kk5GnDOdilgc3PS4zTPAWAvzNcWqAWaCJ4egkdI6LD/0qM8oO04
jrKyDMZC5pBTEEAQBsHGm5AzSV2S8ELW1GXqFu1vqieWET4nMLFf6RKt4DzzLuWgoc95Qt1vd2Tr
/pP7UCzshNpvdYwlFmbV/eiwe6NF1qQL2ZehmS3LZfDUjZKQuh8vWDOSy+lgllFBGhHxEMbMY4WN
WVkpHEs8wcHhgHIF14IADmZ1PX2OSgxaI/lHiNczMhGxmNXNDrDBIO7L+IkHaoqLPWxlXCNs3cii
5LZ9XoBPGJCpYhP/kU3pUARds/3dIeGBE72vg7n/ce3lqn2n5DY+mhhmFdsd2czDnSZ2qRdIFsFK
oc+QG6PdzOsg/TDAC79q7/fFxrLkStAMZMVogVwQ5IqNtyCQuAJ2RuOMJzqyzLS237N3mJetv0C3
StNN6sR+6fOZJfmsfrzzRGrqGOP96aYT6nAtmLwJ6xsPMgQsadVrxoO2tJ9Yki4nf28aDvahmDu1
YVgVEjToXCYl4bUKZ07qsR8qfbX690Ra2ICnr9ghx/amlmES/A7oCK9/b6IYGJPnkOpThZAvbQ7w
2U0ZTYN1y8yibCjA6Sf4YyZECv9BC3OcVOFIVlGXlgpHT21ZbF4oKpHWw40rLYeVsdVwADrLy6+m
rW1IlnHnZu/LW2JCa3jB+B4/u4ROdUmYTJCnoxJdv5hNGyeu61CpIgafhb0dlcQEkCbxxRQWRudj
KL4X47RuDWph6p6BB6+egXpL2Nb5KT91UCpeC6BhWXyYTZk3MMuanz/4yslQkf0gH3riAcrld9za
i15hBJTL10bgt9gGyQLOrCL3VU+LaYgFLE3tXbvjhPrQZKr9acoNIhe741H/8NVhLAMY5fGUmMTd
R7L5hecblZOnsrfXh4RFej2F+ZAzWr9pICqBXkL0n0shNWrO0NbZee9cdGitRKbPMT3KJ1ceSsOf
g9MrxcrZCylxulcD0bOPi0+DPOJ0O/55pr0hE4NuNC0hOTgCSEBOo3oBxmOSRncy5xSZOgmnhlfH
gP5s+SbsY1P7ymjUPkH0UH2Hj/o8AHjfrsjt7ndPdSLQJ1vXWWO2fE+J/WbEnd7akwujSX67d1cc
WGdFYFyoyKy5KRfvKFArUAd0a8EppyICNUEXOeCyoYdAcLGdcPZ4Lzpl1d6tPGpjY4FNS3n68Fcl
1FGjJp+pkky0uDoEI8wNYFIcNXBiyLj5oZflno2u9cc/z3voDPuft5dIq3UZg/fuGaNSAHyv+ifk
Fb0PTSqR5a1f30PrUhzrRVlKImCBBphOE42f7V2kkjESuSJj2bYCrlHtqc5dlbY3DnM85HB5xxdf
BmVsVlmukov4j0nPstHDepZF8rgRMKQPRi59ZAhCkcEfEeEvN+XWV3sWCMK6rT7XdJjX2xE4Sg0y
Uc0kB+SOzckwEQ/oIHQFzVYDjDm/CD0kjJ94D7/llDuKmQUnzJ4m7OSLc5j1Sk3i6e98U4KPLsob
l753FsgOIPZxXEd8Mi6yJUVP0jdVqyjykFh3wtZAMjQWWSeiF+MidL1NRVZregMTs66B/cQ/iGsw
bFJrXhJG+GWJ7oWMKYY4ZygR699M2Yhl+V23pYFjxsbtjrltysMY795AeaTmShXmwlirzoDXDmRm
SS+kSZWT67h18H2O7TmIZqy4ZKnmK3g8E9rEzhmLmySL2ciVP1mPVnfN3/EeYzPANUvbfLiCNOGX
SRLLtv2rWf9KsrNsFPb/HjEfBra2016MqWW6baXWL+LKOqTh2BN5CbsFZoULZb2+l67x5wC1vYKj
93kpEI1VY6bAFc6MgNHB/g+RmIresOFaKnuxt3iWAQf2DrCWC5O08FP3pYVR1WpYB7sLh12BbZ2E
u9c6MZ/QkzNkaSHZXwxAQpp8Hz2+mT7WLPtbprxVcKJv0pRyfKT8IbXTOH/wBMvMSU6l8nuVIEVh
FDYnqzTF4359zUtPLY5yBvCEypFw0K0ixXTKT25LySXHQl1HhgEfkVin0xHq1gNVc9rL7ajNqECh
ivJkveWrHN+h5X5ha34QeXop3e82+AonQ7JYE/ac4tGEAVw73f7X6aHaJOcg1gRxQ/HATMHl1wgA
TAIHlOqTbk3KW4CrQEYtd7JTsI/KmIdysrJINI6jPA706GfL/2WCBRteVGWp4cW8nq8JPzXnP1X1
7aOef4d+0CWOeIaVMTmkGThrfARDblpEOwEWIl6XfqHoAmRn60KCYlDs33T8/8OMqmDDNdB74YBx
b6wg6r6DvN9IM4ODCpSpLYdIFxCepA0xHXeLiQ0b3eT+d+Y7nxJ3CdoLOzk79QP2QAW0VkFiRz5R
JvyiTkeI9k5nLT+ZJW66ZiPcWz+EBJ+2saVj0hO5aS0czP1rT9ABr2lbYTp+F9xCJkBKpzeQV4iS
41tYmZAZRWbEjj3s/afywIfcHOveF8DzGp2ePqNYqJ4frnwkjwJyQcg5EJKXYC1RR6LI0h8jHlZw
jOuVcs5xNa+jfhyuuraD+YTD7Rb0U31MO3ERTBkXZwSOmI+0I928PvnmVKGyg8GN8XmqWbR2oFQq
5QXf659aHN0D1V4hVt386m0hoybRxQc/38VRKlVMNiQrZUVlquqTvZtmnnfx2y6+eR/CmcOkptvE
SjbrEpGJ8zN0BN3eRO9Gyh+pQgIgJCJFPWnGtSDIuuYpJlsMTvXC2jufCrfD+KdOor2vMjuwgNHI
cdkE7DWbm4jfE8vzvhOKBl/W0uL8SjM0QK3zfb3Yw511N3IWIJkWiwoD7k/UlDnZ1XmVr7spTx2C
eBA8Lzvdyns0OvCMG1SvOUE8Rl15Qd1HHkca/4hPq9r8zseN8wnWqguTtdSqKu640+gMPOiswF8f
YwfG0PnYqWtfWlE97RSZ+3PBsigdowvdzHBPGhZ2c5Q6UIyN3wx8uPCeo+73bJl2mzHAZi3HVMTY
pjQYe6BGhUomxKtLV6i3gk99J+9PWLa/VaBcvVKi2oSbkQQs6aoo7ZtJzdIWzTLfR9OfPaHPGdpS
+LVJJKJY9bRzofazHMj/0xBJal+jbuoVXmln9Wu/9xOObesBqd8RLh4ggRGK9Z4cd4L3v9e243Sa
0Ey57mU2Yuwf1zARwvEu1fCwH2z72SvXyWvrIQhqCh+mSKwbsgUfNSizw6JietMKAt0q6IeKf5va
f+aoGqpnbzKjhPuWRKz6UemFzlErn/RddBjCntMM72+DCPAiuDhL7jEnK+L9Hh8b7GGW+Y5tBMov
/73MCTuxoOg1elT028DZ3Ql1Sv6N7Nzbnh2LC/X5XbeIaSvgczRdkb5dmpFysn8WuKNY0rXXMmSQ
pABxltAyPPRfnHv0k79R3fSexBVcq3xPEXiZvU9nCFAZdvpKOAZ6Fn7X3PRCPpHGm0anP9SfG9xC
c4AshXTzAxqGxhuSQ96DDzxcvH8gi9UlrXXM9mH54wzQc8ut/vHtOGVu2AKgjrG5uO6s9iCiJsU9
8OPqOril6DwrdKujpO/fzqmvT7FiLRpWALuaKczxBqEjCC23qvfsBUdAWHJjaq51rylBhCk/2DOQ
eMd8Rjgxe8RY7vkwkzpLJfosEeoJ3jVZWt8qg7hBYII2hX4vD6SZcI8ExzNs2OayHVfRPLiJQ/h5
vXFrEzc/Al4XK2OgIehGuypCpc4so93iB8KWjraulLTh1ylApdwVPW4pOSfSH784zq7fP26azj7E
EZz14D4yis7qqzh0gXnLMSkpRzp9FdYbyeOK8jjJ9fxFibJSru4oYGTn+yZcoLxyRNVLrZ8GYN2t
vYiaJNEupNXNPwC+zqx9WV1iIC5mExBDx1bunCcYMVkAByl0Mp6eafej4hUI25rV0g8Cc43Pe0t1
NbWeSnz0O9MjY07wmuZLddiMcbhj3bId0HmojJrYNIOq2HLHLoYGH0t+6bEkIcq6uMLbSFn89YqG
oFu2yQ/RdjOkivYgkwn8tpSiQvDkL69KPYoawUxUk9iimk69dbPvSqL6jRsNLbdIOh59X1ERSkIi
TzWZ0x3zDDmmlCKi4dN+z1k0TN6k4gONPyGqky1IKa5jRdaNH7ZK4kT1EX7EFi4P04Qr5dFzxlXf
lYM6XjtqbsgJZaJRw13wyzMBKPQhdHSEvgTtZ9xcds/CWWgByPMEIYHrVoCRg0OG5tw2rXNkgZ6F
GwSfZ+zeK4bMhnKYaJYOuLdA+slbZQ9Uem8IE6/sShQarR8iFXEMhd9jnzs7q+kNR04gjr7tTuxa
GLI6aaCkgGVut3Zryq3sdSgZ7YlrRAh6vZoFoWYEoEaKZ6o3cFcUGdFBTnor4enTD4aDpByhzMYg
u8t5ef7HH6240sHHZESz/++jugwb9nA5aWuoxkZy4Bdx5LxvX4A5DGb8cOWEnYNPSE8VhNbPunAk
VcVsryJYSVc5aUpnMwQp+yjfIRMOz42bZMqR8tyq+v+4fvrvlFyWrglAtGfi40TITvMDI3DT/Yz6
qnTXysV3P9TwNa2QtGlMV6Bfi+ch2IwyxzFlKFqbZ5tR7u5C2lZpea2byA4cg2Bn0Ns3AEmtf8b4
WolIIj6K4vcRwPTkqOGRXFMuIFSbLTXPaRhx2b8ysXiZe3uR75s4VMX5NP3BvaWwCn2Yuxs+UXj9
P/npyic7lnP+0IPboO9f1NhyfOYW/EOqWuLkE5iSDS2Kne1In1Kd2DR8ylX0yFt4XYtk9hK0UJwI
N7QHNlImbSy9E/d69tcGN8jeVJwW0ATdsg9sII2j28lR+O+A9z7udx5Fuyde5ph1KEyeRw2phjfI
6h3bkUHPplNFp+Xgpi6NgP/wU/+xeS8BqdD2SLNvyQjDHtGwZ8H2uZ/EhIfb/yfCuN0wG+Hf+8sO
/R+4KMipaFd73ftDqYXAwjb5/nb+wG8DVGuHEApcJfTVaqa73K2aEMUP1eILP87CDKSa4z6oTVRt
2mH5do5vwKMhHVjEf/tf6qc0us1cHTP/T2C7XwlzrO1UGd7u3RyrAn4NCCe1LWBIi1HD4VYsOAuY
7GOk7tY4KHDjqmXrvhPv8yuX0EKQOxZfdqu5XklV0beoZPM3oS1oKkIXQyuXUfDDoitBLVLBfPav
Qvq7OVnBoXR5mxv18FWy1GRDpCYriKA7DhKbbR9uihFSjiXFxqEJ3LQ2SXDxNHWtLBcQkko5WJ1f
l4gDz5vMD8KfhV9tYiAgFKShyyFEXIjOyEEdJFjkirH5GLqh2qRoOXKMepJB91QMtnNwL40pZ/V7
xMqiWIVd222EvxnZ22cO0P1Gyjg4L0yhxnehHwR2cUNvLzYD2HRWcQ/XAJGep/j8oV8KJe/TY/8d
oZcNDtl5gS4D9wZfCUFnqYG+8esBadIZUWgT8mWjwyK+2QVXO15MLQk6HhQg+1AXSl3vOMa6Lw==
`protect end_protected
