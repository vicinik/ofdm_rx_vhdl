��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*~�)���>w�f�Su����cϑt�ڪ�,t4�EЖ�u�Sߒ�ޖ����,�ĩ�M$0"�R�~0�!,k���<�]H.I���"w�Ȳ�(�f	:&Ca� ct`�Qi��v�*�By���Y�9��c@&-�GQؠ����SA[��(k>��ǐ�w��\����i3[Nv��@^�}8#���IR����W�l�K��3��W�P�9e8� 
�)@���t���3`�~�Q9��T-J��;E����
/�esT*HU���d�	��K�@�ie�{ΐ��m&d�j����G�J�Pk��w��#|T΃�8�ѨCq��ʃ� T�ü(/��P�bf9
�Og�!p?b��^L��ʋ��bd?'��]U��<Sm���#�&Җ~z����ʨ5�Lz���g3l�?��9�-6���W<���R(����ގ�$��T�[�_"W�����fآe��B��V�N~qE"�'7��F�&R_��e~���J}n˲9JG	���8\�5tN¤2�|�t��n�2���?�
���ђ��/~G��Ց{4�g��`6:Ui�v#8Ӕ���lS�X��c���V�?緜���?��)��lBW0�U�?2:��o׼���i.a��^�Ɖ�g�!ć������
!�=?s�!qG�l����W�cL��n����e�#h,�;�M5+(h��BƑ|J�5�QK(-�q�k�p�\B*�D|������M�'US銜�äp�%�)����8f���5Ot�#3����V�T) �,I����V@;�u<j.��ʱ��P������uʙj�r+T���6}�6��S ��Cy�tN��mȉ6R�3����9�m�]@`�;pp c���[�@؁*#�p'â��DZ�S�.XN4B�)�G΄oE������x���>{_��$?�z�3��z�Ŏ��T��,�o��e��2�d�E2>�frN�4t;��]�rh��6[����(؆a۽�XnA��0H�������[���cA����<��:U���S�p���)�9x
Λ#l*m�}�z����@v��E%��۬���:����R�J:W7|2��<����Y��*9�V_��T�?�.X_��E���N<�?��1k�Iݿ�>i�2D��\�`��_aG�����G�DVrK/�I��]����n/PA��NI{�,���!硫r�pmB���w�_,�ɭ�Xyv��Rq ���i���44�Q$jݴ�%�it�Ԡ%|����gn�v��sG/�qM�u�6Z��c�$��$����;0B��2�e��:�v� �a�����\��B�N��.�"��x�� �m#\��V�Y{]n}Z7�QTu��~������hZ�h�􊣛���NbU����$	q�Cΰ���*'Veb��)F`R��篌�OY;�D�	�娰���mV���䀉��W� �X��rh��%]��J�c���G����qH��nz���1����|�,��zo|VT��ɞx�Z���p�Q��y, έ7�.�å3�W�gD�4�X��|\*Anٮ(Mzp~��a�Uw�^����De��Ð��-���v��02TM�ʞ�t8h�,���b Pg-#cJ\�0)�v��XQ��k���To�u���,�����'!3FS��IBh#p�SM߾\6��h�\�ݎ˘O����[�jW�n<m���ݟ��<�+�(ګ�3�Z8�gmd�2�s�����v�/����ǮM
���?-�`}������|�a�H3v/�f�V��@g�S¨��6�,�e�����s�3L�X�%�g��HG�f�o��y��!��Μh�J���ǘ�7R4Щ�Ħեa�v���I�����Fb�Qrg�A�yk½{E��w�Y�ִ�#([+�k����y-��FqDO�D����N�7�}L�-�jo�B�mr�Fl��9'5fG����Ј��?��.j[�^;sO̪�S	�3�G-#�o���لA�T���u~谙��w1��2� �3}�<�X���wp�����=|�W�Y��V��|Zɛ�%ſ/���Q4�5�z[Z*�Rm�l��A���L�j^v��%��{�:�SЕђ�Z�d�E`qn�v���cM6>*��:��C�<=F���K���94���t�	�9lY�Zz��I���h��cf:��+����՛ѯ^mȍX,@ّ�#ZFЩ>�IGc��[��쫖o�m��;�bf�����?�>�4{TOú�����Q� c��m��?Lfn���3�Qu�Cr���?=�H��6�fA���7��G�4D�j���N��S�f�"|�l�\�?)��T��)���.Wa��N�wd�<��啿���������_l����"u�şЌv�n��`M�7���ꝑ��{�Z����E;����)E�6X��-%�Ŝ�T���@wg)���a9��>X��V/�t���U�-���6E���J�I�`�O�!;'}m��?�Iwʨ�G��b�,a'U�s$��4�#�^���F�ȆQ��Ai�ֺY!:p9+}��Ⱦ�m�������uOb�9��ك�����zhM�&�W:ТC��~����rq�vP���X1��k�>Vx���
oO9���� T�Vn/�n�Ow���&�,���: ���n�o���k��� j�ݮӦD��'	�u�
��$�d�W�$佨��M�4� Ǆn�*feoCś��VH���~��fG��Z�0(�:.���N0��T�}^> ���'��y�"��s��*����>�ۄ#�?`�&�٪>�'e�B3��?үO�k�OV��N7�����RK���a���Zg��~�5��r�}�eb0k�yD8����m�H� A���	,FN�����lK�	y��)~��s�k��h��dA����D��I�g�UM�Ar���
��K�S�DQtF�K�*��^��~��
n�;?�A:�t2c���pg�Z��wS�r��<r��0��B��l�o��e��!^ TiJ��C��!B����h��89�m| 2Y�I<�m��ry�|�(y��
t��g����#��ba(��%1���2n�/��)F#�:������lz??�(�!v���,�'�=gmG3�lFw����p-�h#<�G���O��i���7wv)���Cj�?L��'洍�U��鉻�U�0Լ�C&/��v"�ѵ��,7��a�<E��O��"�G��|Ɠݸ�v�M.<3��Jü��-�ǭg�ʀ��?�qJعZdD�	��m3�oʳ߯f�90,/�D-��̬>��u����5�U{%S��gg|�%� ��������oR��cxص+I}�q%� v[�O��]֥���q�|`k.�AvA�L�Lme���L��_�y
��l*L�k��Uպ��g���t.�3ĴQ��wN��b�E���K*o9�p��`����H�I�bKq�k�:��<]���F�0i�;^6|O�&#8v�H�
Ei�u�j�Jw����W���=M �9��m����)��:»�u��ͪ����=��A'��o�������_F��fQ���Q��5��ɚ9	�b~�:y�U��	��}m�7��<SKMO�:+�(��^��M�����Q���R�X�n�w�X�����*�K��e��L�G�8���E'v�9i.�$�/�ߺ�[2h������V.� J��u�NF��Go��D���瑝�׹�k�r�<S`]>k[�Zen ݋�7⍑ð�u�Z	�!��ă�I(	�j�=p�"��e7��+���~(Fҵ7��Lh�Rg�8`�I����#���]H�a���B6�q(�{�w�k��y��!�� �M0�F*[�R��-p���@��1�� +6'W9yUY�]��j>K��+�4�HӤ�4�F�D�pj�ء�2tC��վ��LR��\�߷�!}
؆pݣ�5C�
�Z!2 "�Nʣ��t��m3@�h�x����L��_|Lx�����V��@��&��ϜA�{��� �J�a�u��������r�z>*���ܛ�t�<�6P\`|�p%_m%�Kڠ��$������ٳ�% F�.}� �n��[�I�e��Giԕ�f��1�OB����/RQ�z��w6~8f�Aɰ[ǌ��{��1SV4��:d�W���=����0�g��Y�����4ȩ�bdV�2�0�;��J/�40O����0�/Lۀ}�F~�߅۪֠�Ύ��٣�8f������
˔S��sL���.w~
�M�u��4@8}ס;�^T&���.cɥq]J��%`C�tӽ�g�9�h�������������|��k>��r0�S��M�l�5j�7��{W�*�B��2i��-��|��M� (�j���2�����y�Pl��7����}��t倁j��fY��~�|:.cFN�A��)�Z����`�({�ɼ�-eM������� 	o����\��of��PQ���E�n�3��C%E�<��o�0j/,,!�
��G�r���	�h�����5�]/J������n*� X�,ĆE4��j��"�0e��=M�����ϊ����"5��A��O�6��km_�/j!�d(�#�hN��|�μ�F'�dn@v�4N����b��bG��?��:�e�.�4�U8aBhյ�� B\���OX˂_Z/�t}�8��I�3�����<ƑU�ј���(i"����\VM!k���>�.�g��#k�_O�l?��׉�0� ���W�ʿ������'\&�2_��f����9!
���6|w�������Olqn�v��<[^*�����s������z۷E춒�W��t,vL���*�V	1�n��_���������-����چMW�ε��$چ�i�F!�n6��H���`�׶�{�C�D�w�[���g�0��Z�^�n������e��\k�ěȠ�1��w��DI�9�8e��-dj$�0�̅���lr�8��GU�$���
ywN1e'�Ҳm!�	0�\�W?��11�-�_oD�f*����aX|���M[@|�%zk��c�EDf�M�� ���@��S�ES���A�Q�х$�^2d>`y,1��<9?��ا'ݢ8הL��������W2���N��m��%O5�0���/����
8�`s�m=;�wEߖ����;m�p�R~No��j։9T��D�@FYA =>(܎�؎�VV@��L�4���Fgd�1�#i��a!��!wFX��D�7�Vy�5T_�/K6�,�,�	)�s>w�t��S����F�
@ёd���d�s�
5���	��M�3p���w��o@�� ���!�O'Y�76���m��'��LI��%_b+��7F)<_vKʭ�!>��2bOzzS�,��۩�X�y6�c���M�0)�w���O�1b��<h�[�>�%[|�j������f����]�C>J��|�cn����Iml�o���ÉP��=�R��͂mU�;�#鲽��؅.S�Q��}q���d���gW\rq'���K���N���m��e��4b��ae`�R8��I����*I�i��k���8p2a}�����޾6Z��� ��\]�@��ٮC�g���sۖR�Y5��&$�^������r{ЦWa3��a��i$����eӜ�:�9K���Q��6!��0_�]�=XW�祖B� ?�2f~��n�w�n�vqs)�w[�a%�8�U�	ڂ5��n$RS>�ʿ칑_m��Յ�j�����t�[%{�]au���̑i{���P�,���L^P�T^$v^��&^���B�s�<�Ƅ�7��]'�s��7=��;��	i��/��"�L���n�٩�W�CG��g1�.֟��͞�d��w��	x��Ν^�1�{D ���9�.F�13��{K��>�����:��a���`G���E�����6b��EsX���.�p�[�T�T!8{�=�G���M���G����Z��ދ��S��� �kЕ6 �`R�B>_�R��aC�j��D�3K����ZnP��	��úo\�R��\�B�d�{>��D]<8�B��E_~�Lkj���Q o���5��R�cv��;G��6�K��Fw74�b�'/�w;��мF��fx?���0�� �٦��| P�:��$1����?�v��%]�������Yʆ��G=�:�K���C���Q��[�������z��"u������Ж��Gg?���B��v������<�B�*��T�#�f���`�HZ�K4!A/���Q�7@�3P��޷�&��Z(������jm��)���W7Y�����'�DVBU��j�`�v�,'���m����ޥل?��X��a���Λ��Z�g�^,�'����G�,>��;ѭ3'�4����O��a��B�N>�CНC�[4T�¶�~�`!!�ab��K���':g���Y�lܛ���1�3� �s�*j��˄|��V�?fX��=vZjZ��+�,�ds	y�C��;��C��#��A/R#ʝTP)DZ�s�
����,�˓�'>i�
�?hgd��Qqg�_��K����,��Z�N:����-?��7_�o�P���b>�f��q��r�YA`�1{ľZiP����G"h ����n��1���?F��Y��0׺b��������g3�n������t����֨Ӂz"�m�0��µ��k���@�ܝ������\���q5�>,�L >���