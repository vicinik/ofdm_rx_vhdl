��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�g�ezA__J�o�W�FM�u��6�GA�f��;]fM�|.�Khƀ!�2�c�5U|���k�X�5�����?���o��|�JĪ��¥qe��܉U�\a|+���#���/<��^����fMn�6�ӷ�Q>� ߆�Ѫ�ޡ�0X~PіܿƬ���+c#�d���cu��m�����}j��~�X��Up�
�����"݌+�΁6F�e�8͚a��T Z�Qج%�w�&Nėo�h{��8���2E�J�������p�E����}��늘�.�%z��;���L閺��z���IM1��y�7���> �o|V�|�#��]��I�P��z��Q<�u�������ݸ0�k�9�P*��z`�O(��%�jQ�g�� �Dt����➤dФ��RuAuݿ`Lf��f�vQ龈?�k��\�$�yN���^?�U�R꼓<�q&�v�d���.@̷	-b@>4**83# G�����+��`�6Y����R�u]%�#J���R� �7�Y�fIm؉4�7>ó�/􂱤�Wţ�W�F\bz$�x�FK�b���c����D��q����cC��HJ^�����
���"*-nJ��5a���T�t�9(v_�"�#X�~��G��O��c��ff�p�(\� ��R�㱹�}���Ao��a��gq	�v{���Ȯ�@�f 80ZK%����FgX�+ؖ(d�����4��e�>�O)%�o�Y�l�.�S��T��J���)����M�A�"Bgȅ�EU�$�!����j|v�Ϛ �Wv�۪�z��ԏigXV>l����J�x�V��EH˪%}1d��O��M�c��f����C���Yj�/j2�?�]@K��ѐ��oXH^�W���7���OA��L�-n�W3�5L@�aHx��s��H�鿙�2dk�L��;|�����y��*���3�k���!����ێF��`��͹�t����/N�at!
�[�]���v��̲/���w?�{|�b���ϵ9(�47�Nnֵ��n�TX��@1$P��L�N-9����l�F����!�)Y'7�]��qD��V���Cl�D��t��dE6�� N�e�v�h;�V�kY�<T�'�r��J�T8/�e`5k��6	�osi�"�E*"R��W�4!Ϣ��B�����^���E�=~s]Nkt�Qi�y��jm�*������;{N��%���u�)M�I�z��ajIͨ �['�JH�Ⲣ@��/���h({X&7P�Y�<?}�J��o��E�ŗ���g���w����ă�f���]2�6�z�E{	}M�m���dջq�Tم��v�1^".�L	�T��U���R�(��Ø&����"��Ґkd��G7��	�+�7��̸5A�Y����y/|�{����U�T�Q��>3�Z\'mdN7�Z���4��RF��gw:h�E�ze��3uҍ|tVY��+��wl���R3O�	,s�5��J/�<a�Ν�k�ɏ,E>�������~�V\�-Z|I�Y�N�7�����V�	87�����#�6����j%U`�b���V{E,�Fɽ��i}Ql7mۤ�x�}� H*�xcW"}��l�]��W���jCẄ́(v��`�*��0��E$�Iz�`�8pjPk���Њ��k�a{7�:�[�k8z���s38�Sv���)]�q��9�+��Qǲ�w�`�=���Fj���*p�.<���ø!�+,ҡ!i��:<�'(�C����'�R�ؾ�r����>�)=YY�X���tp�I�;U�l�s�E�v��,�T'3{�޳	v���a��mES����]0����zS�EQ��O�u�?曪G\���ȏe$�[�ߪp��<����q��B̰į��ÿ��^s�Ϻe�ƈVn��l��M8�n0�0aM�ʲ�B�f�5U���c�3��u��I�r�~>��&�(��K�-M�f��c��t**�0V����;E�c"c���9U��%�����E������M�n3�ܮ"� ������f@�]�~[���`�3�爊�Ӌ(�����* ?X�U�,7kʖ���a�1w@���[Kw3~����tA5�7�N���`Ƥ��s���D�ۿ�c�(4���Ugq��^��{�
�p(]r�p9�T\�-�}�q�~�u��0&�_1;�j�ä!uRU�f_�_X��Ek��b?��.��77#9���/|p��%"9��M�g��]�ٛV����<����B[ǵ���G���u�\�s�VMg�`�vX~���:9?c�Z���=ZQ�W�G�/���#r5R31���%�-d�j�}1���(ӽ(Ng!7�U-}�6*]b�E�[�^��~���ØV��`�Bh�]�V������9�3��StP��V�����^�^�F_͖S�	%<��A��/CZ=���b`�W�5�.�ro���g��`(Ue,�a�I��X78/�S05�`�X�)����� 䜍�g�et<N�r�u��.���٬�h`B�%������xS��0z���V�/KA=�Z�1E�{�#���D����c�k��gD���w �٣�D&�A]��T`'��E�.�'��?�V[�̥���%q{l<Z}�B,N�����2c�Q���R�^�A�g���C��YoY��HAg2�I��à��q�93��ǌ7M58)k�z�){�Z�6�����B^�i?��E��4�f�Ĺ���=��2�F� ���D�<UM�֧������ƞ�b�)���(ꬪ�3;�Q1�f���>�2�@�k�e�I㧛�pD!��L��g�Pv�a�L��.N�:�/4�u�Mn.���2o3��
����1���,!C��mAxջ_�Vi��G�m��*5�_�^�p�m����{��j��ϐ���k����kK7
d"��y�8x��3��x*F�8w�G�?������*�+`��JG�$w�qv��D�� +Ix����㡻Әr����1H 2��Wى(K�D7עN�#Ib|�#!��B���H�j�vvpi,�轸�TP$�
���9>����y�A�o�q.�_�q�����8�F�3�Cթ����Y&>T�����2�w:��!�c��EJ��mxG�c���D+5x�}]{�֥���V�zJGl� ��I���3�����'�����pRe2�q!J[8�S�Q�W��*��_���0�7o@L�GK�AƔ�c�&Ԓ���ɕ�z=�| j�u��VG�]50����O�p;�²�߿��_66�9���|T �ʫ��K�~��*K_[����ü�;�)/��	O�&:��N��Ms"�4'��X�����;��_�G0��k^J�����$Б�Ȟ��{�6�N ����+��H���وT�T�i�*k"�>��o�3Ϛΐ%�yE��i,x�,tLN�`�\n*�u�e��m�hg'��K��:�\d ��Arg"���?�sm�6�uy%S���X<e�������]��{Z���P#N�Y�Q*x���$���<��4��.�3.i41���+�j�!Q�`ٙ��{�5Ct'�Y��?��o0!�E�=E,6~�`d�'ڕ���qmn�n<Ir�����b���cP�&�0bȼ�&MS�%k���L*H�-�կ����v���ѫ������*�;x���eSl=!��<.8,�)m�N�Se���?�w-V����	�0l�iQ��)OT�7*e����ɼ���"�iE��D+޺�Y�J =��툶��-U���!)+J��t����w	1-����� �v�Uł	�g�xx���tBF�|H�&����t��_oJ�ڲT5��������)t�N6��=$�+�,j��I�3���V�b��=ɡ�������9��s��w����h;I���v�X@P�g��v�c�j�/H��T��������]�{�G�+�M���	x�;�n��A����O� �h��ohl���n�v���l(ώ"��G �9�Kуv�Y���=��g�|�-"�@"�͆�=n�Gd��s��y��#<)�������YL��r^�� �b����v㌜]"2�c�6�\P*��G�g-8qc�7E���s}HyF���e}ۀSϖ�(��M��	���;J6e���k���H��2�q�n��B�]|�i�rL�������B�{�U;6��z)�KՁu�)1��r���ch!�����PB�M�(?��4���9��}�⭌-[҉{��Llu���SD� ~���=o�JooJZ9���n�ux�����.�������&����Щ�2&�W����N�TtߴQ�{M��"��فkj�d<�Bn��,��:1v͖蒟�ԑ�(���oL\J��MT�6R Q(����RO� i` �⢌����{�-f�{u�ͽh�{�V��úts��F&uj�UY��)|pȍs&'��U���")H�+ak����Q	�*�ჵ���?��>���`M"���Sme���	�W�R��f�^١��@�������0}r�S䭀�h���EE_��1q��V~���;>���(ߗmһ�V~].B��e�W{-Z���P��m-��"�W��H��ϴx���D=�MG��%+mZ���^�1l��W˜�NI'���]�3�N��C*�,wJ�3�`ie"�CX���[1��i��`z㼋�ZH��$	T/���c�#1�H���G�J�D�x�{�v���6e�C~n�o�(̵֋���O�M��}�v �&�F|_`&������^�*x�W�S"�����n	���>pލEt(�ʨ�����X��ey9L����먳�C�kw)�d%4{C3��wZ�@�n�9D��Z�N��Yݚ���e)�n�}�
^6C��G����C;*��ՙ�q��0�G�Q��SN��P�z�uշ7iÁ��4v=^A�����py�RێN�0��?�9G��7��gHv$�����(=���W���ف���Wg��5h�I��@ٻA�� H���k�S6�x�_%��h��l.�&��� ߉�4�ŗ􂤬o(d��C�P�)�iP��
�L�Q��&<���X�L�-�g޺��U��Zb2����*Z��F�mp(9�Sw��jdJ��<7x���,���YMc4m��u}��I���E�Emg'��~b4�l}�Kr�u҄y�#L�����
��g̱��C�j%MbAg��(��B;���}�+��["!V1m�a��3�O�P�n��q5(:
��ƣ�Ư��l���V�N{h�GYv�0z��9�K[���W���W�}�=�dqg��4�$��U�	]�nC))i�+xd1���ʘm>�T8>2z��f�3k�����h�=l����_T�)js��8J�KRd`J��b:�n���p�L�_�;� #��z�K2_�D��G&���@��߂�{֦-���g�䁬8��QD�g��|;���gU�&�o��jx��rx���"4[#d��M����8,j��A3�m�'Xs��d��/��+�����&��r0��3!�EX��+N���uS}1̃�Zٌ��O�6 �A#-�Q�%HR����Q��5Yl�0sW<�ۙ�����l�O
���ҩ�ݒ.^��R�WļL7���zˤ����&�#��
I����������&GFLv�Z��l��Ce�z�8Y˹���]N���F�2��Y)�d����y\
�*HtG���s\�k��9�9==���Z�'u�7�J=�ډ����c	 z���|�!�W+]�q��I��@&�����O�f6-U�4F��@|K�ޠS��w�{Z�L	p�c�0����~b�TY�h*�ܝ8y�N�I��uI�V��TD��k�]q��@�=�o����!��R���N���yɢ!6tZP�m}��/cTE��W�i2-��+��/s�@v� ���$�@�ߘ@�	_� a��,wC����	X��c�Sr�©G,���x�[;u*��X�ji���нl_��V:�z��Kj��8����v�;�<���R���u��<��m���ݴG�ؚ�L"�\��R�&�x�m�c$�≯��	~��s�+��T�/:1����F����Y����0lxƹ����6Ӎ4������yA[P�h��m~$i��"��<I���)�xi�ˢ�5��naEHjL��C��S�g��2A��6Cy�͡r�o;��_LDybB�x���wLbз� 0��-\��&{%��NGF�|��5�k@�P*��G2�Dwɲ�d�\˙D�@�P�Qo�.p��Y�|BvD�JŻO�ȕ ��U��:hg��>ZW��uJm&���Ւ7[�c	ҋf�����[
������5����o��s�������ʌqٳ9�qq��P-:FV��.cB ���/���G	��o��f�"�pW��w��c,�i9��|��!�� ��7���)_�m(��F�����k8���N5l�C]��J�7E=N��~}D����5��GR����� G%�E�a'��3��Z'��d�sS��i{s�Y&Ci��}�hr�'�ш]t�p-����Ғt���I�����8�<�wG@Ж���zgǮ����	�Kw}򥜶0۱\vd_|���؊4U���Okz�/O��Q���Ǿb���@TW�9�(���� �8;�P���.'�j~JAI7R�U3�Wī����/=+�)Us�?߳�ǔn��f��9��Μ�|���w�"��p��H4�Lz��ݾ�}޻�ҙ�08�U�h��lk�U|KE[e�Z�d�"d�G&<~O`e|�@��.�s���t#B�w��]>�M������Xo������{�������駵N�I�*��r����'˥=�f91v"����f"nu��"�a����ZD5/9' q{��E3n0l!?h8�T�IM�I�4�F�ƾ*�t���ӏ��ƩYc��Ok�}����9����7o��j�z�����vH匹��$���t�tp/6l@�T���^Y"���Q�� �3Ǒ�?������C�%� Mn�_���O�2������jg��0��X�SPTfKq����Q.��D G�V��CS��#�T�9ʍ���*�;z�3e�N�!u��X�Y+A�y���'�D� �����gݡ�B)H?�Z*���T#�Td�O��I9?�M�'p&�|ܞ�e[��?,��]��h#^�Ne	�O-Ʊ�>
O������ܚ2=@�~����j�2(m�0�1[��3��Ճ�N-��W��բ}��g���$�h&lJ�d��`.�;D�#�)?0A�iA/��Xv'+:�#����]ho�۪˷Y�Q��:϶YC��]�R�0��,���A��.�W��f��8����,�j䫹K�Βf^�otjm�vy������Y���:ٲh����J`���E�Ń?����1y�d5ܰ�=;��~]/�����>���#aVH6���'úī���P�)�OYl�F>D"0��uDG☧�9��u����Xw�r��}{eD����5����Tk����c7�nV7� �qt�J��A� �kFN@�U�4�9��9��Jgx����sÖ��O�����1#�G��s���D�)~
���֡��Avp�}�t}:��g]33��#\Z���.
8��8�vff(�W�ػ "��侸��e��@o�sq������E�����"޸�Z��,����&�(����`���8�|�:1�}����@'�~;�k+����*�Pȭ<����:j���
=�4=0�Q��]�D���d[��oQ�e1��o)}8diV���c�ʁ������|��r�sA9��v@�V�9��k�TI���?:�C�u�V?7��z%�b6e��O����$K3���v`bj�L��H/�F1�/wq��k=�Y�~z�IC����c�u[��x?Z�:��Qb�`��d�ʄ�&Y�Vd������j&1JI��Ȭ�RMJ��y8ǵ/7����f��� sB��{�����^�lM(�`n�ę�i��-��)F��>�� ǂ�����ێ���>Z��	�+0D ���֋����w�t�f�W�l������� �,���b��Ş�L��n&K��!�H%��ދ$x������o/ux�`���	�N=+�`Բ�`���Q�>�����ʳ4vS�ﭦ�5c�75��S�RP�l�p�c�����ٚԸ'Q�P=ć���=-�:���>ec��HUA@0�y�{Z _��Â�0x��#'ˇ)#���dv�O���夁AhxZ����7�vc����,�@M���N�E�3�$�'�<�֗���KX�f��hbk��O�
��%>�L���3gl>T3d8T
���	��|ږ˭Q�����upI�j��ꕗ���w2�^|��<Vl�0���!5)�߿�Ð��
LP{)�+/��>�����>�1yˡ�j��KYI���66�;z��T%�Mx�׫1�TT��a�B�N�{�
�^���� p�9Ǵ�ˢr�'�n�ܵ?�E��D�J�,~ke�� X����� �3�
��X �>9<N������osy�
r��{���_�����uC
�lBHOyTJ�I#=�w~w*Q![�ö��@�TIo�)��'^��]|�_�%�J��YL��P�qi��bcw�d��[i� ���D~Q�VIj7Q��^���#�LI��J��NX�rþÐ:iq�H���S�(�g�DG�L��:�O�#�$l��}y҄Y��ͳ�(K�lL�D��u�B�����;u��l����V裘P�03$�ѫ��D�Ӹf�����EnV+y�Y!�84�	�"���p�t�	�h\|�3�6���|���=MF��` ����
¹~�L�w�W��.��5��(i�k��^�������q$��!!gB�K�X��;^p|��I?�U;=�D��m����%!_z�ТAіDny+�R:�Z�P�n��CGis�e�-y������;Ҁ�R��BY�o� �T�����<�eTn2uD��bn��l��i�4�E-o�'�ʰM9�����tYj8MAK�= �ڀl�4�q�Vo<T��`�aiN���sK�����<nT�$��� +��t�XÓvǙ%�!8��!���´rY mB�&�t�L|��M
4�=�Ȧ[�r�
:�ϋ�Y�D��7`m>�(�4Ќ�	σ�^�����bq��a��Ǽ���q��ʙ���53g�lv;3}\�?8�@�nN6�Ȇ�"%�=Bw��b�K~*ľg��>Po!Mx�����I�I«�75~���O�=ݟ�
b�mtly�>��x��)�f��Ύ�����_\[������m��*�gi c��n��Ҷ�k�}(�I@�v#9��V�w�qXk����6�T0���"z��
�:����K���GL��(h�O}A!��S�k{��p�Ld>�6]�1��Ü2��@�r/rl�����ұ����|�=�2���T6��(q�颗L�:��#��)���Z�ۦ&}� j�Be��RW�<��.�S",DȆ�#�d�+xύ��"���TFr�%&R2D\�V�ɝ�k� .f�E�I��ђ�fv�&�:k���G��8���9?����ݽ�|R���{�e R�t�H:R�to�����7����j�Fٜ�� �S�O}���
��h��E� =
R�ŵ��[SVV6p��'�H㓶1B�{hy3���1�oYo�ZIp��G�^<Hz�eI�v��E�H��do���e���؆H���r
,3�JB͹O,���M9k�m�)�з�����[ ����s;����e!#���O�~7��(!�ޝfT�1<Jb誩���$�\+���/���غ/�C��"�b���t�t=��AN4��C[�E����xy#���q(�7WV/��'�N#U1�9�����ؐ����N����;d�YԊ~�+�>�p�j�5�"�a�����dܡ�z�ȝw�S���mS�ڠ?�Z� '*�v��>	4��l~8_P��ysͥ�[�Z�*�F7���=���MժK(�kGϽdY������O��^K�=z9P�6�=Bo��~K�
!��:��;��m+�G����[��2��ں��9���:�����N�`b�t��w�����ͦ�E�ze���?|˟�ůc@'���6Ԁ-�3" ,�*m�����x��ߐ_ًeV���B�UDN�P���l->���7����˦v���l�.z�%ܺcML)�l�g�b�����)����@p�&�*>
�L����U�Џ�˷���>�A��%����X3��^��ѹ�iR֋���
��1�5ɢ���H���e�F���H��~���O��T�Ƞ���:�Ui�w6�g�;������Hd
� �O�2�ȅ�S+|�; �ލUi���B�����W�@��Y[��wI�`���	��+�eA�sV�?u�,�.?z�LߥW����ѥ�;��歃_4d��mwL�	�j�3���8�x72GJƝ���)̽c4<��~G��Ǵ0ӺI(��+q'5�<�``�_㣨��ǯ������A�fI�x$��m[����ڀVs��y<K�UO�P��e3@�n�A��Q���� ���� I��\8x'�(�kӆi��7�/�3Ȃ3�&{�T$�.i#���8E+(æ+2�bT���&���C߾F�+tC)����t�G�d{K��:).��zד��XLz������2�h�I%��$���5:����F�aXNGoA+�s�Dn^��J��H(%�o� Y�ik�����>�c�s����"�?>��S����ֵ#���e?��];��r��Rc�݄��ݎ��W~4���,��u�Z8�;��)�ؑ�6�=�S�57u�PM}7,�l_��a�c�/��~+�g٠u��qu�]XFĹ�-O��M[��l}P���$����##H�)��D��*]������uD�߼]k��AP�Y�lc��_k�'��h0t��
@��k����m7D�Q�X>�6,IK�����>�g��0U���6 z�F�aA|�����W�t�cL��s>;W
<����g��#>�4Y��b�t��cä��i��E���;�|zIӫV��U�
~KݩBUz� 13�������Yߚuz�nGD� ��XR�vM)���!��8�Z���VgB}Ӱ8p�?FY^���e<\�ι���Y0���������d����1�9���t��3;z��4$�^nn���s�Ad���֊�n`f+�A�PA�YD��,�Q�5��a�w}���x6���%��7^a:oQ�ŚL�o� #.`ؗ�:4��%�v��7�mh�a�آ�L��(?@ �O¬��S'�z[��P���'@�.}�Cu����5�����X&�dC$���˒��FZ�-�ANzػ�^� q!��QD0�j�1z�0X٘�((�o�Qb��̈́�?ks��{2�n�p�M