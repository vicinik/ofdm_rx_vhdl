-- FftWrapper-a.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

architecture rtl of FftWrapper is
	

		-- Components FFT


		component fft is
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			reset_n      : in  std_logic                     := 'X';             -- reset_n
			sink_valid   : in  std_logic                     := 'X';             -- valid
			sink_ready   : out std_logic;                                        -- ready
			sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			sink_sop     : in  std_logic                     := 'X';             -- startofpacket
			sink_eop     : in  std_logic                     := 'X';             -- endofpacket
			inverse      : in  std_logic                     := 'X';             -- data
			sink_imag    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			sink_real    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			source_valid : out std_logic;                                        -- valid
			source_ready : in  std_logic                     := 'X';             -- ready
			source_error : out std_logic_vector(1 downto 0);                     -- error
			source_sop   : out std_logic;                                        -- startofpacket
			source_eop   : out std_logic;                                        -- endofpacket
			source_exp   : out std_logic_vector(5 downto 0);                     -- data
			source_imag  : out std_logic_vector(11 downto 0);                    -- data
			source_real  : out std_logic_vector(11 downto 0)                     -- data
		);
		end component fft;

		
		--SIGNALS
		signal sink_ready : std_logic;
		signal sink_valid : std_logic;
		signal sink_error : std_logic_vector(1 downto 0);
		signal sink_sop : std_logic;
		signal sink_eop  : std_logic;                          -- endofpacket
		signal inverse   : std_logic;                             -- data
		signal sink_imag   :  std_logic_vector(11 downto 0);  -- data
		signal sink_real    : std_logic_vector(11 downto 0);  -- data
		signal source_valid : std_logic;                                        -- valid
		signal source_ready : std_logic;                     -- ready
		signal source_error : std_logic_vector(1 downto 0);                     -- error
		signal source_sop   : std_logic;                                        -- startofpacket
		signal source_eop   : std_logic;                                        -- endofpacket
		signal source_exp   : std_logic_vector(5 downto 0);                     -- data
		signal source_imag  : std_logic_vector(11 downto 0);                    -- data
		signal source_real  : std_logic_vector(11 downto 0);                     -- data
		
			


begin


		FFTInstance : component fft
		port map (
			clk          => sys_clk_i,
			reset_n      => sys_rstn_i,
			sink_valid   => sink_valid,
			sink_ready   => sink_ready,
			sink_error   => sink_error,
			sink_sop     => sink_sop,
			sink_eop     =>sink_eop,
			inverse      =>inverse,
			sink_imag    =>sink_imag,
			sink_real    =>sink_real,
			source_valid =>source_valid,
			source_ready =>source_ready,
			source_error =>source_error,
			source_sop   =>source_sop,
			source_eop   =>source_eop,
			source_exp   =>source_exp,
			source_imag  =>source_imag,
			source_real  =>source_real
		);




end architecture rtl; -- of FftWrapper
