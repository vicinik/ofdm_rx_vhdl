-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
W4ItM7NzejAxzrl5z5K23PUKb5l9UyU2nS5abVNPZbKnvZOtpoblUNRu8d8FWb1VSuAHRedMZQSp
OC3DzAIjtW4aPpe8ljH1gT2B5hgYdp4mbZ4A/OIiwdhlMqVuSpCM5T9HtxwFPmaI2i9Mx8wvLpGa
0XDzv8XDZGZbfxNnXdytt7nfLJy522/Xl72QkgVLkKcTQFXuxkTcYoYXbSvKwvyUyPnxiTP5i80X
ySfvPuazQFA3yaW52MVG53ryt9h0nwzrbneXe6IPQh4SVzppU0nwkcV0arTI5jze2joUg70rGV1Y
CTHxx9lTdntTL3xiNVdmRc1MbRZFVspsxkg2KA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91552)
`protect data_block
chqj6+CKR4TUwavSGx6230fiE/dDMK4GCau+K+CDWbzkZRPv+EgI3W6SXxxnNiaaumkmtNm6ilAx
SoJ2orrBKV8nfHOvAlx/8HsEFVyK0vpEjxqazueprA259L10qp9/8OcbghqGlYHi9GDyQYXz0w1s
orNN55qS0r0gWkshwcPBdcNITcCoL+kBZyICSHOlq16lO208Eov5/H0OA8cLmSMhgM+K0CxawZrh
8mQCMexsL6Es5csFZ2xR9khk9XpTMd74Nh5jfgGcrl82ApkXX2paUZ68QnJm7v+kCKA2hdDSM80q
8YFNA2rfXaKeThoMXqcfpM6jHA9RO93MOacLKWAWGPwliDNa1kQcAbLGetnazH6hPZIZyNEFYjJS
8kZTDT41pdzOFJU2j6qp86QeGPwzkJ6cWDD46hcEyiHykkuE6kPAeOGECQPaX3bnRfQ1GO5QBKL6
GVgVJJSIA55gBvKZwN9rcr35V8MaCV7eaZJ+peBD7KdgVKkyNwQiArXXp5BLMtulskc/sW6aurQq
6p1Q0WHbt+1I3REdMCgWADiuAc5jsxuuUZyaBgVKBwtsg5iCgTnSEY6Lap9jLlIvHavJUy2T9l0j
jrVka23Uc6arlQQjn1vUhlHoAFERnR+BdU69SlaRY8dVDi1ghLI9sortx73dNakFDGCxwZFsSkUB
g6384EyLKW+QJJrB0YFi+cZjFQKUbfzTn3F9Yu0gjJ9fDUM7Mlwj2sURmLy5aCDaHaCFVSolO0mP
iJubsRhCno6Yj/NWVllS+P1pQ3lp/x7LPPqPbo0Xzoj4MmNYqBj1wA4wE7vEKSz+zMVvl+TSgI4H
iFhB53JtN1mSoLHGxHyb31J6yOK7b1NgcGsy1dXDyuhMKJADCM6OmoD7jqA7j9F3svvOuVQ/B9V5
y1YPaLd2sUWc7Q9+jQ9JX+DvC4F9dkgKYd3CKPsOTbbExYULs3dQwBF0HgNVO40cxKQJEcHAr/p2
l9fr1RHZSvK9R4Nk4TB0NkTRnYd9/Tm/EgMvJu/W07phRfLshZKfsi2HqC5hzpNMSCooEgV8YkuD
ZElcTpim9TqXip0NvE0A37f9KyVEVLmAvQVBAIgHybiGIIIEM5X3Bwaz3OQ1aihby35E5nV1+0gh
BrpGQbX5IMrUO/Xtvi/vvFULrj9Dxlb1VBx5AgpIchQhwueRW3ON5OQH1JVuPWERY7C2EgotF0yY
oI32NxMkdfUJM+vI6dpslmuqXC8NyjGY+WJXFgd9HHoGFHQJniKk2rCk4KxorkMNjZA5afOHWjUe
J2f0F+k8Sro0FIDtvhvgQnJOC6+mkU6vwj6mDGBx9gQ7eVYeoF/gfuX8kQsMgBWMJ4Ua5LaEkzsj
7QwnIHi/U3DmZhyUw4bszy9TBSBd3wsJQj1AtcnXOPn0izyTAr7s+DBIaQsSPmWuPeequ5MX6Bva
RNKYELcnGnCwDwJaeHhB0pPn/xmvp/SreOPAT1xsCtF8fw8qTb1j+cjumVJAK4SVbdPE9faDncgy
GFLTu/QYXSeDzeFutIJ+HfHVuEYmV3BoZnhr81krD2ffpl5GfXrPxL6MqN+U//SwuEskzHA7+A3l
hMmqhFEC+tCqjGVwsjo8r64J18RHPwpDj8jNaaOpjMmqiYG2VEfQl/LG5d0qWZ0/Va99vlNnGgYb
ogQGi6LUHG7pt0JLp42GnS69EaYvWU3+vu8zt3NP2Ch0a4/QYnpvfIumXl+G9Of/WpPQOdnN8oyF
V/TciMKdCuD72gRfNQEB3ebQHHyU3rl7A7VCmPZA3PFTxndmOywEUwDGI/m2AkzzQnEGM3D7Ycrz
yD0yhxprJdFVabZemk0Vtmtc/hoMDcrtbFAUBvLc2hrOvXRJLIsy8h7BVYZIOeCOrX7lNvbpIXOT
E2qABjUQjQgL6SXd1dosKszq7n52VOvT49EBvZdJPeU5/Br+8pl6fZAMz8iMF+DeEwb4MC++rWNo
agvlGvaUnccLbFJ1h4zxu2no9QUJ+qZHvHpJRnZC2Yxt0Vb4aqqSTfwt1NXmUchWTqSWBJ95s9Ze
FA3iahaECJqqo9rJzcWqis4ionO9e25Jh163mluDPvaBGAMiVCAKQA2l42hLXRjMoRQdkJHXmUU3
iJmVogE2hAWblRT+5sdDm9rulxQ8Dl6bSpXXz9V192+mzhNDRbN+XCZFTo8ZTW3hHJhbVjnSsdKb
pTkxIcKGGCQKJRcu7tqZ539u3h+3l9Ef0OapP3io0bsd/GeJmrePkzBuT32nnLU3XAqzzqMrBEe/
J5t17KTpc3mTdm95zC1GC5UzYK64aX/z8oSabj7/HLcbXENkrIZpxN5QL0jdW5FwVnCC+2OLmrV4
lKXXZ0EJ7Pm4yDfvlS0CVhu6mlI4jQrkTlJlMgbdhvv+THYVQP4Rv8d4TJ7EnffV0bB8CjJJW6w9
/EZjzP+wd5+a4ftmDtc+PHpjAfXzdfZehU0EJhDWqz+sC+S9TJ4syNhPImzp7Pbra+tBsS1cp3AU
Nk0qTKie1zjA9CHYfNs368OYh9XXmfg5PVbXK/zTg11a+ZO16j14Z5bVns58PHCTKC4te6hKZD+Y
0rkw8RsXrYLBdWZQfbdi8EutYVuvssBRjcsEpaAEyyA3GrSNDbnh9Z2lleIWZKi+MC/UWtjnHTwR
dhfDHQL56Z47I8+tJibKdbiVqOIwI7rXuT4eROIGYWLn38n7noQfaRMAkUlQbRJH3dXn7cskKtC+
UUJ0m0BuKQ7tXKDE0ngxlrDbp1PcuS6V5IyW8VrQZJz7npONRw3cTlixNu2kztDPjKVOanfjGC9P
/TNJotKMVr3If0i6cpret63a494BGfzpZ8Uo1DhhDOmbTs0+QbDHRb9BSRKOuO4chEZRNGe8a8IY
ziENUjBuEJSMokt49+Ppaf6tZjoV2eQtlKueHdZN9vCnsdfn+YDcRR/cltwyiZeFqveG6BdTtmjk
+HQ+1OMfRvjdR8NQqYzsI0fN1WkYQWJd77vkWn8Af6rrkhuLXT+g0CmmJhHxPrclrGDPsL3Kfofe
jIdKZz7T4fwyZzXb7BxB8dqPsLeBBg0IW9IlT7qgSwe9RA//WLkAuL3NLlLsLodmDqnFE/nTk88M
YzQtiwjud+8INNuJPvk4wJeQW4lMKqgasvl9s3X3iZiKYLNNqwg3JND1O3hMIKGw0BGq+lFW0oHA
APpKZxK0I6+zIAMNSUAZkr4xkxBNRGVC2T27PPrJbdn2+VFVBrI3GkAMKH/RQteE7pqImssdjf5A
uKoyU6YMmFIvp2T9zRiLK7Ys7A5VLWoN5JSCu+HST//H4akNg3hTZWyVp6t6HBaOr82KtyKKf4SA
scjoW5oS0yDw7aZ802aoIuZykDwCsITwJjocNzuH2gyv5VTBmxTDKv3+Xiu7Z6/i4onVlH1PMUZI
+BHsR+qoF+JRigjQrui92GCFj88nUbM5A2T4F2KmlYuMFXb2J4WQyTgMom7No1bJ0LU3R8jFGiYz
KO5yCfIQJQiRv/Poam15DaflKgu7Q5n76ZL9X4Xbs9enxXRrMfgMp9UVngoUYIr+5AzrtjfwdcXq
hv1qhLQ2FJ2xMnAoGzagjKubcGrs/tDOidTu5mBlJt3aG0uZxEmwvXNZ5VbH8Ez7yosUYLWbXDOi
Y8PB8poRNWPdzxvpgA8PIAdrCMBhcrEyvfDRfd+SxSHKJisqMyBTvcxNY/l4oKVYtDjk3wrdGjPh
CMxNtnbKAsuIA1TyV45d+VN1mXDDFRX0faYcQObv6dIbahpZh7ueKTNKiXDYeOI5rrUyFNttFCXc
E5Mo+gdHuhqhMDR4cjbNEPQUyvi65qVO3EdO/ZLD6QDBB4YaFoij+eg5NJrJouoBGOOX9TZ4e6KW
hJMtbehSZHnVLmDlsDVcXBi1UPHJuWORLXB9D/bC6YFdhUuKOgPGBl+zJfgd1Nx5mIDIa0zGDe/3
PecSe2vNFHNcSljMZ8PndXLfGCU5eqIV85AbA3FdSVuvtWZxRh7FiJXoqxT4A2EAFEfAnv76sZvC
74q4Hsx4Ujr9qnlN4PY21n5X8tRF4O2jOhi95XlgDRm7xxt+0Bh/m54X1R5ZYsqmCyzsDseBt6/E
NT1WnELfdrR4MHysU3soLvQj/dpvf05sSFF3wzWrdw6hGdesG5TZyNh4MTcRked7DUNn39If4qFV
Gl52RrFp7FyIQWg18Rt16ZUtAaeXz9M5bBp9GWXoOfpio49IwfUBIvEt3TUjUjWVdRw46q+ItQgW
Gip9EzVH27L2CRLOWXi/aVwQr6y1vrf/Uvw9AgSUK8Qu3lnn7GuLfWge8ZJtD8lnjzurSi0vTvbt
EmmgXhxfgKdO+PaQOXDxv9zIF/gMNCYo5CzAbMw2IE/0+v0svVM6KOOE6vboCGD5Y0uBCqyL39rJ
SN+K6i9u80dMUjPKg7hvIfpgy5W1H4k58m93OwkAbrGlOeE4M6S5ojNKZ3CaAo4WIDHUanoNKkfc
qCiXZl+gXACm8BlLQDT1VRoBF2O0FvkzeF5OE8qTLVIP8VG3K6iobIm5a+5Kyo0HloM48wCHIq7a
nTKZh5ZI7rdAHCHkRGx0vjrjKLccJSdcVMb5o+ZEE1iyL6rbE/jwwxFyjjjrMrdSkUOkD5QGIdXM
p9HoCF1qyL/rBQRMJKEL8JhxWP29mhin3sb3fHckqpwcks0WfE8wWl46hcNUq9S2/KmWBfM6UaXZ
Aw8wObstfGLTmo2S4BAlIAXUHggdtbhj0gxX2dnh8FWGc+Pngy+mFw4WdD/DkzJHE4q59JABljsO
fSLjfLCLUfkvuVzAkSgsM44pus95MA2+RiZJfyekXwbCamx95SqlXS85hLrmePIJsDok9CQkJm/+
Ck70Yf4LHVifoT0Cj45scW1prXzYplGVCY349RMggp/dFo2JnUDrQXctDPG5cHzDjlUmGn6Vvsbz
jiHgZBJeXnBMZoOCB81oBz1Jm7ayc5dlOg6hVRlDXv39QRuDwboi5dTRnxzRaK4VWyav7gLOFSob
bxOZ6W7S2k5MPa4tjP27qBf7ozBh1mDlbRYtMtqRyFrwzdvpzBNnFti5Ju1o/KQ/iN1RqgaFpFCd
/OFJZFAuq8oS7TQURO6nVQmJb/RgocowixscxsHuzfqLm/6Sh9Ukmq70wbpBaJLlqf+QGsoJW8MF
j09wzEvFrZIZO+vVgWEOd+SUMs/V8pXWQ/NG59CQcbRXQ3uu8qYQ0JGDKc/6I7n6BLldxAzyieHN
0qCWlXDRwdyyUgmJcXK/b5NovWX3N5vcUYHQAp0Xsburn9LuQd1RkiCk4UX4F4wXkuTHAuamucSo
OAfq1UJk1mCbb520f6X0p/6SWd2AVVmzkE7tEKJ7UlW5P4xj5KtmF5noqy9zvyKE5ybXMm8AV3II
PwHqDPXshUraH887Mh9z1+16Dvh0C8tGZeiEdhlFJmrpgS0YLh4yBiJ+XkWMbCvagtsyMHqm3RYP
eA1CFLPNz4Ksvb1qLBI9nX59ZvLu7U7wSrqqOCHbaUvoHl9+kJT+V0InfhpOzMn2UXozcQpo/TxL
i27kDqn7BoYHVySj8HrIrHbnOWU2zMYspi19C/rvnUsCSX2GhR8jsJWcHesmJk1qEeh9OO5FT9ge
MZ1MQbE47kRVUu8yXlMmNpWEeCBCYhU8UF0+29tx/7/c0h5n/ijGuBhgUgVjiOXkjTvBTmfvKtWs
IIVphCnvmH6GpeT3d1K78GhkLm3yQtRnCJdSu2abY1c4IZVxDLO0JvCAK2K8StVaC+A/4GymvsJV
Fw8hKhKUukH1t+BlNmW3UQrBE3LgZVdPMlEh5sKkO1OqHUBuEmoiTkfUV7wZZ1Sr76jTUn0z33ph
KS8jK7vOI/ayZ0LzoV4m30s7VK1aJXMggRXqxN2rvc4vcOar1RnoIz9ODxV0sc98ei21PNKNjyom
jQYmywaVsO+eC+khwTHesuas5lN/pJwW8v9vF0QVnauR07zbVwQdiJv3ci86YicjcuqpVF7LJDvr
5giXJ5hRFXt+0aEyR/pnL8kZcf8vaPj6fdz5rdKtwXY4Hw5OdL3FFQd3NJCr8ogGn5wQgVhmnMwD
99nsy5MJRjVV2SmTZTQ56kPn/eT5IScyRUrVVqb9acFhj4PFMsCiu8ksUyMrO01jWjjSONQhWtZb
yeBkRPvg50Ls1kQ255+aniSDlvhecb1pLRTul+dooqAiwfmEjqMoIrxejT1ue4xzVbRNqlFaXj4K
uLtSE9iUIizH0+6FpWt2W2Pjiaf9BRwcqht+/XGsRHFhayy7N4qfJulD9Ld+7bQsjhZUTgZS666l
damJrB+mU6PMu97vt+t2mQtFsap06mepqv1/CnslEqCG+QEsgSp5FZrmHodyHqXCGGELORrrV1Wd
SxNkuNGX8AE7aU5cLUDx20Vr6hy4aqaXWCuvwXYPrYyjZFqVo3pWXZIeaj7GFt7GEOOaVkosYCqK
zQ/0KpmXhvonHEOWpBbKUOwkJKpHtl428o1WEk3z2ojNygW9C5jmGBNv36AGT3PX5pLiRwoZmSzi
xidCPhv2gti64eUwcaYwj5BzF068AkFZ4DYuEzDn8QAlsEsdLTMNDFxwE94Nh0YU2izTR07G60aD
vOpG/ko00UxkHUIyVSGnnlbZ1pj8E7ad/yEMkmBsuhi3sx9Uye629YRqTZQviN2KZWpKFz4fcVQV
v8oYhPOzE0flQXr73RuK9/0kTzPX/lhx8Q60dvrBdEi3erwYtE0dEKSr0ZUmVrzCc2QpCs8Ce/YM
tNR6OuwRviFmn52Gpi8rCTgz6cod3Lmjh2HExcF8AQneA1+lNwTOhDWGQXs+S74iXZKUlFqyGZQv
kFIkF7wF+6XrRMUbLGQWe2x+RnVB8JtmO71g/8xL904hayK1nemtdkavWOcncAspMdN0OSSUm8W0
5GumqiKqNAtBax3CgnKOs0wMj1HKdbqwR1bbWMN60wTB6xuY9HccSQVJIxlAT7NvDZavaak9jQYC
w3S6qI6c9YnLoW0KS1ZvzGlvHrRqJo23zuSc88L13xRmq0bQ3laRbf5qeg6j0EZ+UhGFmlES66dt
cGnxOjR5gJ5ZIx328f4Kp1jesQhPhwivLaxAJYhKxBUrJccacrEehCXmQ/+ab4U7IgB6bIulZSrg
d9O1IAxtLRWUQh/Sz9hJ3+eOd8oJqV1L6LHYoyO/IT9uHZ3vVqI3hrVAwjgDlWzagCGVofkjb/A5
knVRITynOwAIBVyvkEZqNE3G8B+34hOHitX5riau3uqkRegvyiQvm/M5ttP+ENSlMWmCUfdIzyXy
/xma/WtvtbryOcYvjUKa3GFN1rvY4umTlmntOahYuUmCjHIa9aplj4+gY5PuDKwYrbeaAWXnmbeg
P7qe1cIDycg4Pp8/J7KjLMYvjhpQ5/bswR2B+Di+9RmzH55jDRc77c7K9gMlteV1+/b/1urKBFG5
fWpFOygQ8ua/d1Lq8wFrGYzdyOQdDZoGAUaxRrmVZsyDi9TIXL6qHQl8j+Kd0aphQ7Fh3BdxBxfS
YN9Nvf8WcsMDoc/jECNAU5ySFc04GllleiDfHvrwFvV+7oJAPq7TTwSHsZllhtypGeJmk9avou6l
IG2YWILwLAdShYHN+NOBQr/Gg3HVRrLl9u6aMfmx0lYtuoAgawedxEZt2L0WXYkhEoLobhqKkHLp
CbVY6PGzyLXGuTA0FguYiATqibcHcIlPXgAN5jlgokYVAB/mF7X37vseYiVTPcmFfhiDJLK1rLLL
xWxhSaJaHvlue2LlVkL1rq/Y9jEkSe55QkbF12U6HGcap+4VqcCjfSv/95iluG8HOgjQC8NHSeA+
CxtZAKrJKY6N/2kfnEhDTsR6wFIXx4mscx4uEYUBF5n/oU9E+95WiYbqII7eBn/mvb4Gl1pQgJtG
vy/S0C0aWJPSVPuIGmdTc5iIIQEnd1nxV4BPMOOagL0NftEzyBQ/nov8Eu22UJXGl3DRufqLjE2A
74/4T9fZ4wHoZRKFgD0hRE+dQ4Qepy+cUN35yzgSqDE4Q5jO+zYUthXTLNDIY3BU3nNSwaQPefNM
zsn8Nr9+a/gyQCv2gziaO+PtDGnf2juQ9mTKDz7ucWbm1RfBGekD61JusT5SH2A1OHdr45ZGiOcU
6BtBI1i2fxFTj+vhzjkzL2zuQo3f53hoVVZ3395/3YB5m9Sb3iGwuBfYUt9fTeIMFPQIyvylkbOp
FcQHXlXQBOQw6t/B2rYJtIfvD+OQEWRvM6hqcZMt5bsblVAiH60F3KlrJIMw7SJFz5wyR0Z2XSAJ
rAqYX+2CpuWJgSL0KOtN4tAtKaFKFBExABLax66n5Le3ui8qyCJbXB4/WyGguzmXMO+3s9TLQuUE
hREOOixFMFva4o0SsLGv70dcw0fyxyv4c8QndM3eZX7nEHOZCOy2yC+VKNdgdYof8qhePFiYTGoT
ZXCbSfoPwBsb7F8XWNqjlwAWDo8F1y3VXFAs/aQUl0q+4KG0giW6Hv2v/0jAcyBf64d+dDkGh8SK
SXeUpl9yhpeLzqjV8xiOV+ab/46XSnOI5ZFxa+nq1DTWlgfQ9n5u/wfh5LG8l0FxL7Pg/lPV8nLB
AIrneRan/FIPR0NgrE2WhrN/1JfS+6Cm9cQMmdZwZJSRAIcnj4WezkpX3JhRzfK2yXqiFc/Yvb/q
bSo4vE7259y9x3ooiZsyGnYP9OF9NS5KL4UWFd0Cd/DcFjNCuME24a3iiRcrO+HBWQZOKAqLQvuV
7+0Ssk7WbOXxHc/oL91dGqLRyatdZY5Z5tAjB2kwQHRwhYeW6QcAac56lrEQTokmJ2siApnzXuqE
J9TFXTvrkRYfSZVZNXbB7fXaDe8uWERI6bvjcykAEf/Etbs1bTaYDTYrs5f9+RLXW5Uskod4SaQl
RJxzZ7NbbVwGlUJ9Qe9qRlTVjx26Ymlj5lW1CRCUivAB3FRO1kyvSYse+Xw7xjMj4+yo05tjYsiC
yxQlpn93+FcRWM+p5RXMfMJsFokJCUL+b36UDPsV0b+GyAIUwzbCzytSrZ9hgi/ev9paIknCEXnh
CF5GaTq6RyGGF6YUDkJWSUA5O5knx8ImOjYjqZqtRRc2S0Mp01WsGXf4LZXThah5GWA7b0WqzDK0
XvR7xbdThkWVvrF5+2n2l7xsIDKoGSzHA8+xTq+g5XDMrggzc0r6crWdrCKi69UBb9xnYw1VNHse
1bPCXjUWnW20aNDeWyMP1H+Ejvn45x3pHKlTBeRZki10IPFxBoGqAjAOBZO0Byi54xFAOxt7YbsW
vRxnA1NjSEI0a3pzEgG3e7pnCZIsCExryDurAAr108iwc4zPFHsSmNOIR7ejjS8HbWGlTghGqkUP
NHzI9kTzTHsmBxPRd24RFJTfoS0LH4bYV+pkRbRoDJ5yG7aPF/mz6xTKY8WOeJ5iZIcdYiv9Y+Ns
9ihHZC91DdSx0Z2cVxkqvGQkcoLYEHB6tERCSLuaZAeA2M3jxX0q0BM5W+n5A+W8SI4qVMGXJiD0
5eHn0H85yWNMutMDBmvRPPJPXlmT1Cup+odN8Ckp+3FqRj5kCp/ZQH93LbST7qg5RAqO//pFxLX0
PdAfLR4wcw9MOrPBnCkDcYnb0EQOtg8Ilnc7BpmZ7phyhfQ3HtfwCfK6aXlqgde7S26iNRrcZoju
Gynxy67LQZ26pHnnt9x/Aj0wtnHiSDJNxrg5kval0ZFBfFfjkeZ2B/Q66AB2xJ1+s1TTExbdQA6q
wl9GrnVWwC6h8rdOE5KMrB1+BBvwmkd81SKMu49kl69KNdNOaJ/n34rYA8RT5mYgZ0MzlmrJTAZY
DkGCAd984zvFYpUtTvy/Isc4o7vPOts73VWQlVlmZKj1WLg4EfTbuv+G/A9S8qCgQ1Y6nObXQ+sD
ZX/6d2snPF3pKYf8XYjQJ2iMxuZu14w9FbLv0Hx9N1TkXxkt2Ea06iJvmbWSJRh/PkB/esD2vqMC
j9jro2+bEZWekM7RTWl+qIHqs6prd0QyTUVxpRg99OijJ0zwNm5Rm/FDByrsq7S6iJR+4yIxA/JA
9i4hzXZJ7NQx+paG7VBkjLVTQ7ieoEkKXPEbWY8hVmARuO3ZpXQBW6o8t13BykVByVskVsDzyDhH
rk2jFKa9KCSfNZtgs2D4IcaiG/iZcR5kcJKqjt8Ehrs1o5JaKYwb43SKo0UX1SaVt8LocMk7pHj7
UvO+edyn8bpS6cGedBbPVb+7Kqgw9RM0qTOTmaOQ80tpwuT8nk+N+jCteWo8Dfjj3dznbxwmAC7M
eWVu/l6Z+mWew2eLpRKoisGyaAKKlXugTh8mEqNONoMmCtLWvC+XiEOfTApGgggZZQa6Z3tKc/QM
ZZpoIXXfpuVA8tWDqgB90KuhmHCB2pH9u8OMufY4BQCKjOjJsU22atYipHjK7779+FpEmzJwfyKh
BuDGyoesNht9pRGyBqu9xzN5nf3Ehz41wIINZMkcBowzg/CGipiVfV1QnLgeiak6yTzTD+4E/YUi
RvKvduEjYkDpX8poiIdWOLA3u3xM5rq2GF4x4dcgp7Wn+DFjrQjBV/jb2TIpOP1ecW1xcLCTNOL+
q0BOeLJujyZ6F51S93eVeQ5PX2c1nV+LrCYwfm4EaFLliHzdtcY3n30E+erPagmfFSsyLtbn1rWD
sBwTojNvUGe2LNK8TI/Iu1/uCT3lXaRiYxqMTRTRsDyS/FYxNOwvAzUQcrW1rf6T/9IRLZX+jY2P
LyH5emdFUTNvn5MnXRR5g8tR8fKTs6e5JWkJf+PvJxEkB/EzhRhzHYEqazWQXxlemKKuNJHjQ7kP
0uRPJ3cVNbfC9tWDT62+soXBCv/4FIU0MGG70UgXhgcxxtQNM1uYHKQbccGlc6MIxcEaKUcC57fP
uxwc+Pz/ZlmIi8s2ILHBY/BKIytMyFV360mD58BPNXO3wor0Yw82i4PJ3zDFegyWj0sT+k/u/yyI
bEMp+wT1/uwS5GVY+Q3465V27K6QyhSTHa4FPM7RQjOrWwCjqvKViiT8x33ZGy3Kchue+EbvExCd
dt/iuI4Fr/hlG6bLH03mVUFmlp5qltD7apY3V69HIDzbzR00tDppq4i3TmAGMlZJZe3nI/Py5XK4
yeJwNDDrbThbvGJ/0QxAealJ5Muekkr2q7+YbZqGc5SagmcvdW6eWN4BpmvW7Sgbdq1NRjnAIIN3
uI1A8kIA9D1wfWBrOIaF5BPIzs0JT2oWuqg4LZnm8TzbYrbJS7kmlfKzaQKj4CYXhpZz08swG89v
6EJI3/324o7npe8UHlc8eVQVGodVzOb5xqD4h0Wcx41hf0sD5rGds+5TW7+7HC3TwPHgZTdt8V4K
NcJWwFwW26QIlEov27rlFJ3Pp9pQJ4gPCcVjrROWHouY67S6Mcc7O5PBnTds4i616ZuNZ0ENJitd
iWsqmoNV9nt1ElCO5k5+9nrVwaeJg2fZ5intoy+TA+zGIhW3b1VuOlmHdGQeHxeNQY/7xjJYfXjP
1+6KlgvTPJBlsGKIoQlOU0PmkTTNdjSIFTDAYA0UPeoDVQlp/nRvjh6NaCb8iyZGFjW2lOgPfrvA
Pzhjpc341UywBsfcQooeGhiJJS0Z507BZmaN4KoCBrexrOrBTLUb83xLpQaOTyw/JU2tTFFIKZjq
p0UmhytJWmpuo1REQEXQjkQRz1x5PtD2vpQAEtdqwaZpwQQZHkAVXkuH24p8q6HhkaI+twHNSsj6
sL40JJigoQxvFVlNsuJNFKU5GNj2nyzPimO7Mo/9JgS/oz6FVjZ5KrTB+tD0mGKhr3e19m/TyIkH
jXOsiTWDtdIu3rfxv1syHXQ31+su9IZANiuAFGsWiRI0FaGpzzcN8ymd9FnhjKf4i0h81mWxKqng
6NV+XxPHfrQ7zijzhlQuYNwvs4iGA+wob5eYw4/HMKboQoHbPUoBn2W5/45V0ZatP6byLneSW0T0
p0Ev1gJ+j7ri1H0PobAQW3R9YdTiLS/A19kI4YXebTS5Tstk2+tHg06Nlp+nYEDTfzuFMYmkNnLz
K7/ZFsk7Fk7iczoAkAn6WEUJNvmMjx/7bPGIBWc0+W31dLIm811oH4VSUUUazuZIiBMICwK97vkj
mtjpGAVz/PFyWFQ3oDBO+AaVw8JYVNzoUQqDdGym1zEx+H1fjMjp33R5K0rmME4nEVzuxjqrX8ki
972OcqRnPNaEYp4tl8UtE69KYi5N+xfcV/qDEhiMuv5uSSK2eTMi5Gp5fGZc9R8/db8/E6Q2Fguv
xQqLewKz6f4lUa94g77ChEwNzPDO6a1Peqp2D5ZXrUfr53u7JSF5BbjWHcnwPNfsH1NDjS9mfrcI
2EOiSda+dshDt5/ERwyAv1HPQd9aupIp/7+k5DLFXHtH5dxDwFZ0ulZo5pAmz6OjHIgyR8JR/hLt
o9nM9lD3Rmj9stHZ54qTMfksmi167b00xnF5BkztPay5Ai+VmsmDUTuncqhpNg4peTliM5nKlrPv
pH8l1f3CVz9j9F2FFsRFD/y/QSM6yZxoH0/dOhm4t1zPsYktdZjn/qIDF/HKz/prIp8Dn9Mu7Jpy
s8IETq2FcI3RKjXfan8xYhbQe90kofND8HWro12wM96/dtOfa4s+axeClXRkP1EooDrMPI/pUQjv
t//fGCuEAXZMuFn9HMPaNp1iSjHFbNm/MQ5Uud3XVM+ob6vYECJ4GRM4drttPhD85KqlHDGUrHGl
8BfvwbtWrnk8If6J6tTGw5wzyAKMKD/Uo9AvN0Qc+p9D8YAlr70r0lJRyGWBK1BO7w2mntqoAnjg
qy+UkEK+xtDZlFvvLpOVOHV0KerAckCMSVDM0LWwoL4VG4HZEnniSuNnThEIHZb7C1BJMjxw9tB8
Ih1X3QcsigWDJDElPPcuHNMzlAYAOP9dTeNQZDGEAuOntUbkCsHYtlZyyDjN+tjtE4GwlApTavRX
iBA5GLJP9N1QVrJc6QjPHCWuY968vtXTz4Mu3V77xr0Zr45gIXs7qTmR2oMcISegMWOjTLqC46oX
AGSTzvTn4e/mYMp5hRAAJGC4ONqgwnyUvrbU95/7Ps3fB8XkNuxKM/R+jBkgQHsgRW0FqD83HG39
tv2suRBFdsPsYajdh+66FmREQAykXHSoWvx2TWIDxGJXo/FiG/YNljWbM9Dmk1vYi4lGT2bu/B1o
zWxeaD3l6lH3RTm8Rmp64Wc1G4hvvcdU9bllDDUEP5enY5OqYrnVqOwfYvK1pnYAY4nb2p5unln/
/cWpXpLgNfekeJ9EucAV008dIegUteih8Xlvtr5DLXO0OoXqdX+mvTrAcuXgzGIDz2KhHQZ5nHMJ
I/AOTiAScx725/o8PAoxwY0qKMQs63c7Al2Q6HubvfqVGfNEtSaQ3f/3MVErqPVx2E+zvxDK4j2d
yYbuXbx2/cbVSuNkhpp2eSTKfKBc9jRA3Lm9nO9wHFY/2PU8P8GiOzq0O+cCV/vu7KtennqTwo2g
nhdbya+IINvFaJgbK1B0xlF5ZO5Ktq81xekPx7uc6f0AHMa2LHzkUgL+YMSCOF76JFQCC2huQree
HEO4p8BSe6+22RgmzYJWFcYZVECKMc9uBKC3/6TWSV9NQ1z0C9X8dCmsPp215S3z+q9HMBJz5MAf
9Exf6L7n6xF487buSwG+Zv7JnMGKHQVIABt2oVS9RWi2rGuhM2YyFCZiXUPQ6bUaGbfvbsBsJZ9X
0QkuZNMdXxkUF4fes+WsFCzRhb4k6zTQTn10Yki9rR/TURis008frRWtcBBEZPF+eS/Df2fyNXFs
/qteedQel6ZTzhUdzkNpobqvy59FGXhf4XDxNSoKxBEubAYgcxkRAiVbqwFwvk0JW3QKNZ7lDUXt
0dCldRz6CU9nI+7zOxQPB/Lutkd9K7eOAcCQQEClTeDzZo3fCDkJOk5VXkhJWkppBnXaL6oNCujL
Z1dNzM6+j1Mfm/V5neHjO5ZGEd0wrTUVvBP/eY4wCU9g5ODof7NIV8dIsoIkXKlweQo4I0TftNHw
i8Il2xJ+kmyAzLO+NJ40+Un8Haye9dFWjcxnUG1ywZcMQVgtl93NEOAjSPTw5RzplVxPC4svyFH+
QbrQNEzSDT2AppMKr3ClhzX0qF4bFMhiIOowslmdFiFJNK+wF+i0L7uR0RlGtQcRAWOBZe8vMAVV
f9tUWANgydekQ9FhXkYpI8pd5hui0xAZqxALG/R3JUhoDq7M1L5PoLawLEi8tuqRy8RDcIXY8eai
WCd5QWsZwmbMvFGPvwrhUez+E2n6KItnJBIPU7vrJ3CNp+eHMRaqpUzwK8PGAe3mmFn5vx1R9crh
unCSoYY0Yb9raAIRYp0RslhxdyR9V6HjPY627jZnwgw5zv0JpfOsHWYgZ0Oi8pj8/zaD2pZSIddr
vB9rN9T3hQjxT3htD+xvDZzoOB4SAxkR6s4rvs4TF/e7AjJo4AuzMo355BFpLBnApBtd1T5BbFZd
2hLPe0kZxJtzf+ofRUovduB/ha5XcJkNbmP74lVJqz++r0k3rVlCegnqyxXt+aw5T/IsArWuhGwD
Ry61IMpCPQyY4QKlvPjPtMSsMXZ+O8BUUzYuy/lBObKnmSIEgBsdc77vQky14NIYQigaEwKhQmLK
I/VwJam99jFZfxmuSzTCW1Z6HBHkRVe6DnJUw/eOPGePTfZbZFCt6yb/KW4DJ1n1aIPsRIKAJXy5
m2j8O5rhT951AO210pxINCtFvFoqqV13bafPuZsXWCwxTyJdz0c6D7T859ZSMWzqBlHC7JFBM5Uk
6WYOoszwfCOm5c2DMJAg2+lm1GuYQ5bes4JPmKW7L6AbTOAczoZKQK9wSwzsXHCF3JAsS5nyd52e
rnBgzoxSvEew/ctxeZgSprDAXAmMiwJaXil//GvZDpG8FnTuTr4ErPLBBWPZT1JWR+1PyeVfrGwT
67Kopg8XFkWDQX+MkGTpd6Sn8ao4gbCGpU2XAw+s3GhpJeU8HsWgiXtZVpG4yn5mF5hIEpPmofuC
NSLLnIAv49QwEk2lmlV/25jPxm2iWsGLsS974uByKsGRKMxhi23uOe01Q/1SzWZGTaQu8uJP3FKM
mesH+N29rRMmC4N9AXN4rdiD7HXI/Q5cDzaEjL//bOU7yimyGjvpEA1NYm4RbaaS6m/pTz7cu7WD
iRLl/pIKU/qfDMZlrT4pkUwDBxCVZ/sRQGpgn9IrlTqa/5+Ek8xhoVZtMptEANGqDcF+8wDXPsho
XO9xGlBdOBxkf6sCcN+1Xk5wrEoo9TQAcp/2kXtcKHrvn7FYX5UvRSQzoDgC+WmCeZ0cfcc6oKnq
NCPBPQbhX3VueNvVuNqB5JjR8kpwv1R1bQ3u4gVSt//LA8lxC+zcxjFuLl4i5D1Tkb2zyRORNwQv
szYVP9Lb1y9RKp45TEM6ON435YwwI6sthNrhT7AnOgiBfQuCDrMjkkRCOiunRelAbHAQXrFnkpEH
qmMmM1XzvXyfagY6cMgKbO44f/XI8l3+838TjjHM61emSCfujaoilYSuXNU1OWVrTVSnbxXT5sZh
w5b5npePDsr1lxkW0jh+FKLXlqFboSjbYFxR83BMQelWaS7Cgmhb44IF1ClGX1R0wh/8G0ooGEWr
wK7HyPJX6CmdFzlybZBkjptjJ6wuqfRi5ihjPqLypkVhvubug7QPsyngsAwDtSQmo5twRgKaX5xm
j/tIwqmdkTzaOZyLbGq/euu+yLKGLI/JZ6dvimhny2q2vQXILklcXCKxU2GXfvClYH5CjV7x9eYR
9T7MuqiMnx6WnOM6xkZAy/WijQhm+3AwDg63wv2D3KQ1M6TGbTdGYB478HJ+m4jlmz2ltzmZhOs4
l0XAm/WtsBlLeEDn8XE8njhwluonJ/yBkxUno6C3TjSXlDVEeCXaHvEBTGx9vhQeiDtt2pjyQ8gH
JS8cGnmmcjhV+VA6ADjOFrw24ky/kI5Aoc0P46kVMFmt7ayLCHFo2MDzP3xn8do3nureAs5q6PfV
BpfqCdnoa8JSq15k9TtDJT7vGM7DxdD83FD8jYNsv93o06ZioXSEBSX8/PgQ8vOimQMsqpK6UjgT
B/HqSy2JyPZByLfIp1hcB0djoeibbpEB1oVaDsGp3TRQ3AsYTpHeFchUbUZ/P6oYM2L5I1RcNN/i
5dO6K7vNWG4uSorM6WR0cz2xLtmxlEq/znq5f96FzIUVNjvr/ezCaJctv4ZyXEBweltIa1jhGsxS
XM0PjKqKtWSShC7PwEQAZOFhIOiKm86ZHqrilVJLAO1QB5HPetOTEKFrBJYYddclikk/f4eCjnVZ
85oZInJCw2ozoYoVjd7J8mgWLy/oU8ufHOzj8fQknr+P0X1zr8f+7Stdkt+pwul4nzYjg93F2Jmy
nW2DcJvIA6l6nPNs7ggilmZBBXO/flwEwnsFBT9d6PymKxoLwW9umASGZvRJ0ilGtUTM4liWHkGX
0YqRrdsgjbQkPvW10WqnYThoxqoEbxin/6ekqSzvbg0R3huDDy0m8AjZQDu7FMvPoAfd7oXrIUoA
bLwuwVHPNUxL8pGh37CdZSmr2pws89oQUh3zrWb6FiPHU2FoCkpdJKXKMj+ZabQRXBFhflismHP2
cukn347BEhCs2xncgl/s/50bW66ycm2lI7ZIYCRvx9bc4vRGnbTWn7CvYYIzETh6LYxIrx0zZr2c
BcrJthu4sIa4zTz1teMolXWPsGUpWwGqlVRb4sf8B2Otanu1xkNWDRVxo8g90J1Cm+nAVyxYcLHW
0ResAEaXSj0yQPpid55OBt0+fHO6yqQJwKJrgEGZBJJ3tI6QdnE8xjvhfggsWG8PkViXItUcmSM5
u7jEB02FomXRXpb8thnzHFL/DJ4/fIxMZnM4byMTBsYKhAlW3hxvA1bbM79IqoKPRo4K10L+ctUF
1jX+kTazTbMQCMnb4HrC5bpMjZYbpwc9UA1hno7UCwDrvOlaigz1+oit+qORhMWPBNuydQqS16o6
l/tUd59rMYDtAJ24fNaWUaFjxMiPlKemrn0Aot/RkS1uMQeLt69T6wNsePXfKajtKwxahzF8FhHL
b3aSHxUlgLvW1wKE+4Qw68s/IcjcmQYIKRm38CS87uHJpaOVWWw/kCGJht+AwAzX+z+uxusj/VkS
H6AiTJedyNbqA1Mr3L+7ZOaWxuSBmfYucXxs2d9spazDzgrHJ8I4yr6B9z7nDhRPHUM0rtrow3Pu
W5eYL/fWWNUB+4NtGJhpdABxsbytDbMhlYnvXEWzPY1DpGzefpMQ2VSkoLFcUpnnJtlsU+VdVGEw
7hxlqw6VFkjySH1t0rLfURSOD0lFxxRXeNcUjRP3Eje4tisU/84SyaW7nQ0Qy5VM0RFimtFZn8zM
zosH+YrZPJgmq0oNkQVuD2OkeNWJdr6VPHBRxQXSJSKkpT6PJhKKDy6l637tg7P0jowRtiyC+Qgf
jQ3O344FJ2lsz5JhgKEp+Vub08CN8yOHbzuNJ7P8Pey7ATkGSzmFnl0XcDKXVNGUVSWChGyXYaUo
pd7bcEmKVKXzHlKTuL+zrKI49GM2udVAJ/BVgPVpRA3Sftb0g9ieIOCsd7fx4af6Ftp8wOD8frpP
USEH2dlOIhLse5WgBsdIZvUw08g9NMa1OMVg/OT9v8Oj1euHnlrmk6uSczicpNS1rz4STDqpSklI
/2U3z/VfEHZsiDAKeIpcM26cw6qCXHJYiJJ+uDsbsuk9jhpp/0rXB3X0V7mt92LY3Y8Us2nKcDqx
ntnYMpCXQF1FF4w08kzuKXZeh3Un4j7GLVQdWNTLPeilLEI+JMpG8RCvCS/tJAO/ouAj+MKyd+dH
G2PPDniJlX/64WERK6mUXtZDQIdDfqaJT2IMa15K3EW5CD2BsieOEXp/AtUyWobd1yA1RQhfXYm6
GiYrlCA5fqYbQ1htLATZW1ow9oRQGQM3DXw9ciIpMmPSmWiZNoKHS/FV32C99HJIMvD9LjHa7yHk
MJaQw/wGmFtXPJ8IiNw3E2MvkIncf9YHH6LKeEcmukakvuHO2e4YKCxDDe6bC5MfsNcl1b4NePk1
JszKsipKdoGJUyg21ByL/tSboPWLdzy/kptOvDmE8jW/48I4dyL/kqZCwL+qCU0R8XLM69jrCBj3
vY7159A3FtxhTtkSywjfttdKzKzu7hm62Q/glWpM3OP/0BqSlDX75dZaDChLIH4FgWO7D0uZNahT
wY/42JXyntNYceIcYhSlsoFY+mOvuuQZ5Ravr3yE0wEYH4isRAXdgDUjnwlibioeBNaFjDLILdPN
bj/zufTkaznxRSgvDaJlIK4sYlZtXQCop9X8LkL9Ky77UK7vcgozlL8LjvsFZmMH3kVWanqnxsjW
KCQ0YuBqCg8IDyKPlJcIs+WXElgiNcNFnd7JjUkBZwHDOlDqKgnBicqJIGj0b6627aAOjcERi9zG
GMYLr8v21sbKnClnkPQCx2iBOpLecbH4uXdyPAe/4V0nNg1mOlq/VCED0xvH/+8qugPA8bvFP1ml
mgArOZKO6IeKEViBTUCGqeLpRbQiM0bovNuNoxnKaZVzcAHdEa6I9QrIv+Ck7y87QfQLsJOUKgbB
JoJeT3RsU6+m8dbmFlzQf3vDhY0tms+1xgt887W1cjptDAMbWH/f9pVuMKJ34s5n8OoBS/KuXUl8
UQqwdiBwixkkI9rLGuYjS6ZQnhjaxfT8EDHWuTMo1w6+tkbTd2AV7sFCaX25sMwxn9VK2wpivhsE
Liep0XB8ZdyOtu77FIewmEVofIlSggZKYKkmuJNh871PFfzatkFL6PwG1fKOKoBag86ri/y5g3Hc
4uPpI/vrgcmvWjNqjISzgEVWI2OEcj5efAuc0w82hIqv4X4EAtkQum+4nxArQ9X4HFEE53M/s+IK
eaSlSj6xYlruYx+xRQxOR+cJor7A4DP71Ha3MEWbxILRhvd9ht9zJSLmWfJKbMobMpM7DYeA6YnA
2KmRQGKvKZWHDTbpkDuknYI+WuPaANIOysRpE3+bY3tCcWqpumupeoTTDhxdeFlPPu5B8YSR0paP
fU55kxg1aKdWCHP/rAb6hS/QlBQ0MTuJFfLxqKVSxms0/q1hQ7YpgpMNah7FDPjWqIQhQGgUAdVF
SW/raG66H0+7iJVJn0GfgW5i//FOJjS3miKQgp8oQ4ysiPFhMdi6TSDY+0HRTOyiLu8+Ol6ks7q5
zdq17VNp62woTUVnA9/E1zaxpbi8OLAX1kqe+bst1C6I/5IXyXkehLjwhB0q/IsjPWBBrQUMHxOw
FT2Rogh1mqPPTdIlK/nTyjd1hO+h7ss1iL+rNMsDMNrnwnL/LASlvK9LjO+fx45BtSH2y2yivoub
sikLutHPfEUKHhcpbuBA6qjaoGEIDmvlpxW0XP0igv5Tfx2exz2hQ7XSrBfoHs+AIyv02jmartBJ
hoV4wXNICWMlGlvbC0fBA0bDF/Bsq5ph1x/qxMF9u5DMt777SlPtQUMqoZ4mogtKwg9w7vAPcJR1
F6fnNgDC5O0TnSJ9um0I3ZHFp4yNDcc0xSxvohcYqxgzHr2g5qn9PKhAY9EA+3JyMpzShHeGqdKf
xpLvHl+pYVUgLAJ4Qzodua6yMbPA354IjeC11QyKfMCOxDB5EEYK1s3ns9WgL4ikPZyNERcyw+bH
D+yyQHqcIFc/zEE0WleCc39u9EIUk3xFeNAb9nh1tYeHRp2OExk736RmJ7sQy49mfpbC9j/H+7Jw
QxTY/vGACan+UzKGnTR5VqRBoxZipfrdTtOig/2PGU2zkhASbW0qoNKw1DrcwVYkZ/xK8b2ZAIg/
Hd+ITZpo7vqCaV/3hzFseQt/XjE0OZEvCP7yDsEo9GqEeiJYQoTAYbL5bZTwD2QcgJN1wJb43em8
epke6O/hzhs/oRsqq6U+Y/dOhwUfe6z4Xs54Wbxa5DLtxTrLNcNWaUE2acC5aU5EBLk554mAFVx1
YsVVlrQQ0Zb+xRTCdyJIGt9IsrVeXexx8i3/DruxFP1GSz62oPgO10bQzSwqfllkw4x8Dm2TRwPS
5CePBQeUq4dv4mbkNLV61xurMshzo1qxVfLx7YCaqX0P5TcYp9KD5RwvAVUVN69tz4uri1M8eLUL
ttRgVVaimhhEOfpqkGS9wEF6cBaVJ0bnAN93N0ndQQP2TSiWaMjL2jotd0auPs7L3uAW3uaKnl7j
9aOuhOHoeH2X3b6UL14gnx8MJf7++NqhHeCadD/etDb9XMISEBIWjp9D4KmsPXRPrLqAczVHbj44
kEDuuuOAlRosRSALW2nO34S5QLhXqkIYEfBYGz9PFPF46PcebiIC2EVGdK4EEK8xU32vnvKZPexg
xdvV+IZNJKfmpQqbcYhYnu1j1lufn8Bm6p+nF8AJBj6msKWvrr28zCoGdciWlMdEER8qManDAB0Q
2mpw3kb4yFkR99x5/Pj6OPpe6aAO5D2Vhrh1Zsu6bJbRQcCPkBZnvVEins4Ayaqx91NK6a/Glp75
Y403/vn3Vfj0yOE1sjdFd0WnpEeU/GHDqvSRmk+YW79nQrDDBRykeQ/Orct/6Wb+nKi/zpabX/IM
D3LxCbvimpjWQG93QUsAJb63vCc63uHv0TCKo+q4dbMR3Q/Upk5BNAmecgAN/nFT/mIZF0myGx+j
YANYcP4EP7AobaK7LjFr6Xl8x1aCK0vf+tdZVWoRQqYBWvsfCMA0hN4KWG0TK2d3iyo/CDRjHq9W
8KtvRz4GtEep95xdOWHWfiZTsmH4vt4jqDjeZh/AsiyXaxtw5WSEnJwewokCh0J+9zS3NGKEvwF4
Tves1I1GwX69OOjVTgl3uAa35vAZ2GwhTc6r1kDM4WWBdEyVuomsjGRG9/eGEQ6MRcXrJl8M5hI1
zIp/Y85ANdY65bB2iR6DuEKWRPTEGNXyWL5dLUAIUX8/RreLj2Xh1mj6ISYZvPE0o3MWDhTkaxjj
c1EUnR8OrH3dvGKywBMc3arh8O2GZqcFVrHPoxkd3qyz+EloWFB6ICC0q0Ga94GPZu9eROm4i7Bs
bGDDj78S7CTtDWEYf9e358frpU7+XPMoXXS9eL3ZMHauY7ymPgTOV+znM5K9pCJpHg/ypnktrpkU
ZKjmtswchmbSaPsXCpDxadz9ftfn2Vnl+6hmBuNTVyIc/38HKqU9hqCV0Ab0VDXxdiEt10h7gBM3
0MakxyxlIJXpsNAQx87SQPtcpKBNrVrE5JBvIAQQpNt1UTdmQ/sNwwK78DC878LUqAlI5/YT3sYH
wlTmQin6d/pBmU5OiaOZ4DPHMRXykeaBA4W2PnCFds9ZFJ5u3ky/aEcxVRKnFvLKhfeSeRrdOgIf
I6/9FQh8x0lbQEMyJ6WauPHNNca6TpYyKZrjd46ZYDUzHx8FJxacwaD0g/4bWAGFEL7M/gQsxSdh
guGCIbGuMSsYn6CkOXrNXc4NYnW5Q0QVsWpA4IxJAq15VbfP+9sDEH8ECuGNHQpQFmmM0luTRZfk
1nE9OyMtQec0XspnBLVeAPB9MYWMSmRYrXE2hbPat+Mpgef1qeJf7ZxId8ueFjyrBrMCaMskEJyb
8QL4t5Zs58Gln80NHg0fIZ1cSPW1sG3hEIp5LVEncTbLMhpsz56YvFh+sNH2LhFVsNpQat3BH7IL
YQzMa2vUEyZewt/lR11NL00d01qOjDk4d5V8Qw0pvooIZPEYDGsk/eCZRVQKyO2ghnj3d8+MAVgu
wQnO/CG+KTPB/clLK+H4xIw0NOH8WdQz/lA9AqSQJe0qF7QCnDrJtRQXtH4WcVzzWf1l9Mr60uLY
0MVHhvBBoPcBlFuYe37z1N7To6dLwsf8KfK1S/PKjU69DoF+Kt0zl8+jsLgdhtmHHWZOIXDd4Ra6
YrBxdl5/fLCZ8+P9jNII+Dv64XwXJMu0FQQA4G+wIxNmwljNQ5CQMEoIKMic3SVhEQcLPT7dvuxa
zfitGTP4ohyAy0Kn2t8IIsidbzHQ9OvYC+aUIr9J/uL9hQCx68NGwnirpQO+h/4eXD9ElcdtATKY
Qge6Uc8b/4anByG7XFg7gvFcLc5rKU34uB0bwhAMjadkJa1p9uDPx3NPdeQ1F36QKxuZLKLJY+pZ
UOmrqERs8ewDjzyothEU67usu07LOI7zybsLlVIKMUFdQTYH/4PkD8OaYhlrpmiLEDC0PiTj2aUR
FAJ7tp0kIsD+nFrg/M8iGRn2q18vItFa2zeXE0vg28+werkZJ1yZEbcbQ5n7ji/WMwJEsxRHDYiJ
on/gGGljNDEMZxvE701PfB8MWiRE/yCkHq/A7eY3PTPxHIcSmKtaLk+ARXViyHVKsuJllB6I9tku
Hp8nioyIrrrfjUL7DEu2/y6CtTgpkZ1SF0b+U31zA4g9nFWjJtStQxIgRm5281xyaPjo4b14nVag
3wnftBXHY0HlQ6uVcd6P3p2ZMVhn44vLxn5jlTgTVuIdRtzaIFpOvy6uNFJ/HEnn2EQePAqD5ATF
DjxbkF28QEMCAPjwEi1H7boDt3t6CHYeWVc8sLyfbCeY1IRSFs1o2jGAr0twRRa9NeCIEii0NwSm
CzT4Y8ojqa8hylgxyy4DCSyOeKQKFcxT5PJkfpQYtFNQJV6R+kKwdVHslAZ+xwJmgVA6I3O+4j1n
68M1lVll/6fZWIMwtK2z/k4HMZJSmvhxmTf2+xLcEMN1BduWwO8leBcqgJ38IMvl46W/xFVP23wO
6AvnUgGkeAZKBB56WhmY2ZVKMy/XUV3BcljB8+d8aAgfOLvl5b/gh7WyZewUnv4oVcOUuHdNlQii
E82LMu5bUfYFGhdHAf81rwZG9ekKzI437g3oPICV4rzd1442jbtbv9J0NMJ2R5Ijzqm13izjZOjR
2bYfBH9+IuYtgAYF7WgzNOuOXPRuvrxqrpIrf8wIWSmGqVmruKuu4M3qDn9vHynrN82TAzvXNtMY
3PxhItfMFrX73XKakjlCGZUPwrhrYwU5f69iuDs22qHwL8i54TN2Y5B0imfDwBxJ/TX7m25VWGeN
rK4TY43wRAVodE32YEuIn/s262e6+Vk3AaUwiRsw8I7Dv4Vtrips8ayK/KKkwqiNjanQ1SPINzG8
3i2lxxfbJkgIPmR0OQdTTSlOCPcW0zC2HCG62Y8FG5+a7zrp9KgjP2QICq3ZTetdF8R/2kOS0ev4
heSWvNozSY3jIt6e6fW0V8WHBLQTGymGiJ7WLR+RnfOAThE8/3FChmC4zSHnW4atshBLF2l8iC5y
iGIi+RyERYx1qCf7wXDIxaF1x5HkcDbzR20DKivuCFnUXwunVzIlqMJDmOl/rbiSU+HeICFEMTRa
qQ7Ds0UHQV4Ir5kHHNRoCbVQG1pEUdRQezyZgkGLa+mwrpwE5EMkc7oPwNKcj9xwh9T9W/wqRa85
pse/zX8NIUYTJg7KYOolRMInVedYhOlDvsi5YyB5Lo1jb7sTH8rYIPC/hXtedqNdz1xdsirRvbnN
opmqZqGZI89DKqywcRXgVMcKVo+fKWYy5455KRFYab6ry0zrTPyoh9cDJBlOPAYndmR1fYhGCKwA
tWH8bxPbS4lwW/jLv8P7zG4yxn3wvPtVTRNjVlx8sbgblSgyrSbRKTPT2FzcQt8MAR/yh+17isfZ
JU/1DOT+Rxv+560LBOwHFO2k3HzjtNrVvOQT+h2JthpBgoYKVh9+M14hG1mMbaq195eneViHIRu1
JAn2qzlq2Ic+jg4TSb8TApIr8gVXW60ZE5buQcW5rNyojM/wI5lqNkNyswTMDQBk4vf1ZfXY53me
sGNM9OyyuBgh5DVyAU+Sf1JVRBqTkp0j41VPM8JcSSolRVTLRG0enefpM6VTGkeS2SDLC/r6rwIo
quxcqeVo6CHXFIEnX/54ZBkExoVd9/iN6ibtYFH4fYfo+QvM2GU3H4BR5Qjg6WtPg0xXLJfpF2fn
1527PFXd3M5TU5i26wZ2H4Xn5cyg1LZygd7lFf3eOTvboRQfSqw2znpXwJUByX06Lmhok/GK8C8t
QgOI4PDe0QlSzuuvKFxr5VHtVAB9n+JMsRH+wvUQvudWO8oGW5QgMOiSVDvzzhRtZYgqEpB9P7nh
qmqIJcCbYWdarV/KLaRC1wDBk0e07hNtgJWXMgtGfyvuUtWe7o6BMtkikABhbrhXOuncsWN2nnzs
72Uy9bOVLrRTMmVPEIVrI3Li8HnfogGYHEcXcnFuHiwqMB0tbL7Ydh0S8hwJsxmdS+pI8d9AEdlG
JvwG7XnJIPjTYiiMDjPBTCgWYvvsyl6jpTE1u7snHRmPCiATsRbcRpxzE8QiXx4on8zdE/zbL6ZZ
2KUhWig94uHl3ohTr+V5EbXmXTZTAE6Lqc2KZCdJrZdxc44JwWReKxLzozpfQ2pVv9e5+N5MQ4h3
jl/ao6w8ggnVVZiKTuTV4EwMGrYoE2UP1Pytd/XHgQ21o97h8YVAU0LQGdWr6O0XcfcWWIqSq3pq
VWzsGDgjD9mj1VZ5nhJy2QTwrSBnpksNZSeCrXU9aHvQPP1LUpqPc3WpgRGWIs37z8sMzEVSCoX3
cpiZfHyiEK+HL+JZTCOqUy4vmq1tPjBnaADT4eV1NKkKyp2xXiSDcz8lhCWoKur8EfUTuSsUEdhO
rSmSC/l12pzemOOFNyHJlPM4EY2tpYT5UM5CnfVQxOhYLN+ljZxFESkfQxNTjRTfiDsTBjvOxLw3
CKmHs4QndifR82jOV2sk4JSCVKXrvdaye+aCjtK0lfj0ISA7IMQFO0ZqF8YWF5Fh7bbmZgTKnUNB
xdvuDaM2vXd3RcHFX5idJRIuQ/IEvgtDiKQNS/pgLYCFUQhv1l7OZPJczMFFUfLwTkmw33SSdxBw
dkSs6PYV8W2Tiadrm1UvVCvsZlBsOcET6OBuIZRLpi32VuA7/JCbe6mLuGX/4d+eBfd7HZVeMkPe
0ngzvQo+8sOZD7RvTSq+jHlvzXnjgyQ6dcS9mFIC71Ow7fHBRwmA5ADgKYEsdDRnqfKYdQmp62TS
CQrdifAIGd4I0FUq6g8se4N6bGqgJEYDZ+Xa6hbyUT6kiHpuovEkg5y4xQnSX6JUwD7Uzhk3AUcB
0wWhNuIlUihu7lplTD8mkfnc9lw0U2ZaCb0Offo8l2mfyxZwt1D+KTWj0N3ddfdHpUxT4X+smK8p
DyG8q3927Gy7FMeR7DybKd7+TPFYWlI94z4xIzN5hFmkWTHPX2n4sNIQ61GxA5bhioiJ/uKxFIMk
d3Pl7fykZxDUqZIShzjwu3/D4zHG8zV4FQ/5txXzdNLTOdLouWi0eDtgGk3hSdOiYtxok8llhzVf
7eKra2+0aBJi/kmBY9oC1ZImiGaEKQwWQjYJv1hwi8952rd+w0kbSPBDKY14pJ2rLyu5GWPukY9z
n7KzOJ5Qq+ok8pWY146+pJPFMqMqMDgk/XKO1ZuMz+tuZLP3CPqlz2z2C3GU5Lrhe7O/V+Zvcx3l
YM52hI1XIfKYqgnTciTlLLBRNTuqO28lPTuob85kLNRCP8v+JbBRl8rsY0ucdnY9kIwSPXCIJuJ0
kOyf5nlH5+oYcgbmsMeGD8RvD/hvODERS070oenNM9kFCrYd/RzDLlbOiXzoFqzP1PblMjN/9elJ
kOBUobByO6+3PYe7KnYwitqyljZtHzGRpMpWCAl1tLfjWUMJEwacqIJSPQfhmIl+DLbpfDkYZYxp
WuNCePUSZh/qPJUHZiUB/ppL7tHlwDBeY0GNd2A7cHammyxfSJQ3PwGJ/gZQu33U25PWYWZ58ZmE
Vvy98bMWRJXB6pc2XYhDYXV63jK+vZqouSfaRZ4uPKYQmmRha11dWmIqoMP8KuPoH/YnGdESAese
zy8SYs1aphlfXAlN+kRZwzXVdUD5X3ocZ5oVAsBt7U2CiHkZiJolZxOUmm5WnO3eLq4oOr+fDVHL
5uMYbOQJmxlpYnZlTUa5M6N+hOsk1ItqYJ+5/4WK2+8sEdfpjOTvM5mRnk5ssbBcf8A301f7gvdo
GFm/wP+6ctmWNRXvJ+C1UzHQaM3Db/7iu1FD+PpYKaLKX+/NQVwNAe4EtCiDj/pLCOylqWZWBsNU
pV/8qQq2eAE5hmV+b4o7+bckDydl0SGyInyvy9QNvc9jCrS/opRExGGXqMDa0DkMki16mrRGzAyz
ABS6KandkW2/cMPQWKyyCfulPwWsKthUedZHLCcQ2a/Sa9IHJVv9jwwEEMaTwHYFaU9wB+QJaIKG
EexNm8GTMGQHo2jdPYFtnc2yhkOcfXmOx6DnHCWbs2Gndmf7WnMj9dfC1smcEsnSF16TS03ACpar
F254KUWzshPcKIHdZKTTDlaV9vNmu2mBQOzyLniQ8fewefg7QQlrFBG2XwZ9HQyyINvgdqPa0kuN
pskHlreRYc2bwGT6peDpEwPxTfVhwZE/Z/mjIg8pgp/Bk01Vy5Z7t+G3S795ixxPQ5xAZUSBrLvZ
t2IWSzKTK9E8FaQyU3Fu6bfT68JFA/mmLhwDHwsUgdAALg1seFvbjKNWusXBGqOwUc3+XDeo1j7p
XVR94499ZUT7TKt1JGgb3+SYR8R867U3En/RX4Yo3TFx5Ki56mfEToXAEQLS8r259lqCwZfBcGNQ
OgmfPrh/TTn23Pb3CqZT7raC/21mDaOm8Gjrm+XHDu3ssbBJV8y85bOK5d1FBb5zd5JMVS3xOJVH
tfi4vsr56wFBPp/4XlaPauEMiv6wJFiqT7VjvVml+8L6yH1NvaCu/syMOk/rJFk0/cvDq5/QRzzv
s7o0HEenXe28TkK+zDMYr9lN/graubQRKt43PvX+H7Cd6xl5c7L8ROyDuLY7k4yLXAWZObz1xsw8
jeVs+KWTsYOMzr2RoLcuGO/ySEe523g72JPvPnjUXtRcNKTuoH0qKnRaIX/g0k6IEc7f2gAHYFKe
vrfXt0G511A+cqxLcasPHbfPwUF4pMf/oncMLeLH9ORMqsfIXmAL1BMNQ43Py+IHTjBh+gWD0Mar
TxVa65f2Vz6HwvzjBWF6XutANbLBL9OdqGdL1WERUg2OQqvlziFZOmgoe2gPApRaqgRA5Rkd2Ag6
4elm2wX1VQ+5xl+ui5sZCLI/dcVmgHUBwy5hQdO4pIYdbQIP623MwMXjQJRtWEyMQcsey4ZXc/0Q
24x6CKzn7YUI8Lap6CwesXlKMxPv4n+Vkgc8fl6d6kNvfA20l4/3mp550Fw+nSuCYWguVMDDYZof
GcY3VqF2OjZmnHoKXgfZkhxNR0nd0aCVOgeNiZHrX8vjA+AOLFAoFob0uGhIi/AfGGmT2P3G+aG0
1OD9tHI8KgpOE9JKOM3kz5e8zHG01uGrcjPsI06nvYDoCI5XPsLr7wmjus6OlSL5ltS+12gjomg9
+GIMiulzwqd5ajU5Ox/FxiAL2ineAPizrxzgAk0lgQA8WzrxbvCJcjuV13V6Wd5D5b21ldiF1/nc
jUG6mD8SeIcFBcsHoFFivQJHyHNoid3bRxHQrHaf06bf5S1+1sJ7JFX/6QqieLN05x5qDvovZb2d
trBwUmG8r1f0aiRqDkE5xzRSZ0Jjw04CLtddhXgMofpP2y7xZIGBQY90FYXfD3dbuhnLzRRj6Tm6
/M055iIQ5C/FZ6y3Fhy8DCCRSHeY2CUNSYc0qfRP/VGltItaVdsLAHsD1o9C9RSY/9fOzrG5Etaf
F1MGAprGdkDbq30/O1fJolZwc1C0UO5gBhZkbldTW4gZqewnGUuK572E3hQkAkMcxDKy7NE1SOxO
rPcUNK+34BwqRq0SL9/xvGCxTVF2uFCL5MtJXHvKe8Ml8MoFvvp6XIvXKplJ0O+HC4MCIO2vVZWQ
ytF2i7GIvhS9WBYtLXM91pPbGjIpgNgon6op8CDLlX40rMCOFLrFiPdoFVZldXhcYgbFuJXf5YCs
2NDOVkEc6Bgb3P9GF2OB2yVvHI2VUku77Wzi5FHE89riWLRShXBryztw5wV/mbsCOQ9PtIr8qZa/
Zv4j3DgCwuLgZQRoodE0jVcxcOwZTS75f6P+o8scrbBzbfipIUJ5l6AHOUQ3TPAhNJTyLcmvLt9c
asRkZOXqbuS29wUCoFmq0cf4bsipkfWFY2IVdb/jRv32AF6d61tNeDfvpWsOHtHUSby4nCZP8wwy
nCzdyWV30aB72AcR+wxNukXlkgqVPYqRM9xc+ORnq+eiNNJdMHM0eMLY9N8WR9tiNoZupn3DafRX
QXMrp42PRSbAP9d1RoAgr6od0vubOTAfJQwGbBkHwMWoYFPgUrLemJfWfFBUGKZtvncbi/1zh6Cz
wE5ProKlNbkpkd4O2mUehwf+GU7RMqAThi7Bz2/0wTKgYFBMk5ZoN//Twf6KQvdioB7j1l0JIFeF
rpYM+LnaFKveyuV2bfkAPjsVl8KYj0f5VpBn/JTZrfl+smlO6EoPczb1SFwrGaZ1nkE3K3PZVCQO
17osBIfdDW0nrYJ77XLHAnLTSBOm/J9IQ/K6tUb25wXGI8VFo3OUDZx0ixqxrXWbAMg7SX8T3+Id
XWEkOfTmDHjAvDhHoP1mSHD7SVHwnJV4Rk+Xp/lL7aVuIbJEHWtShaxkpRwHWdhQrLz5I1ljerD5
DsuDjduLLclLojEUui0+rJDKcAq0JKgV+hI/mNoEhf4/16iq+8n7CngiLKXtAKaW8NZmad8Y/jnL
xSDKv5OK+HFewVgwperrwA70rVdpU8DsQbIV+PC/AZibut+GcFKTqRf3GaQDMFV678URJZdlFnQi
gjI0KU6v73gDnwAG3N+Ah4nxREfRjC/yGZGqm6yo+bboXQt0Mkj3JM4oGLKbT/u1PAzZ4p6Ib60o
xg7HS8+CR1T36vL7FLo6tHpFrdYj/dV6OH715anxe25E6jf3eg7hcNkn8vrByjzmVbix9og3kitD
P1T9kzpkc4To0wxgm/raHRplgJQTgSGYSu1MIXTAwz0qtmOtP41McqskhhjhL5eFH+p7onvqazbz
BHwc3FB0rDmJKhY/yCTvr1BYgIko+pnAWPUTRkSLulFExpcysKH0tMWM+ZkuNWglw7FP5AneqRp/
zLLqKcao5Eh2igJ8GjcX7HQZKqroMB79s/lXPvIVIZ3tn4pnStEV108ur7FK5TotCV+MIs6hxU+W
xIr/quS74X4i7HLUWI1bGRGkUq2XD9Bm3CueRZdpBugNi1VujM2RUSd8WYJq0PeYPHgArYnZ5gtY
iWu+0YZOz7B2MrHG0b/1ZeT2qAnj5XlcMuhEXIwVNeWivjl5TjyrYQ/AQ/dJXl5XC5z/WJQo5DAk
7g+U2p/uckC4Oy2nI3/48KsqwxP13kepPJfGoanhJVRpUOGvqbQxq3KtmPDlwuCT34WGXqcgFztM
olaxPoIzYThvnzJ9QWqwiyIQLT8V42GdaIROMZR88CJBcMlkHKfSfic3j2uj86gCyN2Yxz20Sr/o
7g/LnyHnoIqkCUWEdLAWD82Mru3bpnxH8uw7UQ5sd8RmcT0P+nAv6s3iCKldWLWUHN9fqTNm5cSm
RQz75xVIF9vxjU6UumNkxboyyHmaUX1K8kfIb5maN6vPqcwpeVUUqLUoo2eW/TCuCFRUEESUxSDD
IGecSaW9mCP6fieuSY1gSpdKTPXrpY+mBs065L9jhCmwy3rTbQerVGrS2JA/dEKZS7NKx0jkD63N
MW7+bLNCbNLy4wqyO+mjrTq9KOHi4eqwJ1/UunXcznFb29JN9X3nJNkghCAFteppM3aZJUJjcRAP
Pb22x+Sovckfxp/BYopkGlL5VUKwLRLiMnhGVEZ/4jWe65/5fh4QRRzVJ0eSybA/RR197pKb0Me4
7bHTisGNIFaY0paB47JAO/vZfTz+0ZWdENY0oAjSe2i9LevhLxj8cudLSwxqFMEzfAoUyNqI1psm
YQPiJm0Bb/+ZoyS2nuVlEpJOwoyJBiDtzZ+u6nfoD/yJg8cO5c59gC6YgNlBjYPwLdKaW8HqDwT7
HNjZL+P+rKxQ69bmM6muguw3FyRXS1RvnCLww9c2RjZ8bos6nP/p5GO5W7tTG+z82it6qCWXZvjF
B/dXaQtXXHI3urczbyUrqaN55N62z7qlaM49r2UDbGSvzR4T/aM/ZvlLceVG/X9sx8Te99UWjfbv
oN/glik1u6STsAgenm07W2n6AF2vxqH4YTsc+rUnkI/Yn+rgkBV2DIq+gPxEL0qr883mVvRs7ccD
clwwM08JMFYQdAme9fns/NfqA3ySLdOAqhMGhZ2N5MbJDokuWfUVD8xRwj7w7FvJT25tIROHNosZ
ssbGaMrtUiea4mtn07S+b8I0ocRhTrzHC5XHjtuAgdOFrpD09/mv0oRBewus5+Q88feAB07MP3st
5yx3wyUv1KT9KOyUTUX3z+2zwd/TtUYb38O+I3pGNYZMg3ZdP+oQJ04OtU0hkLw9RuRHXr7fn9Pf
at2O1FYjv9HMv7RG47HJ7qva2O62so3w1vLTD8L9l7qCUEamtUkMVxMlm4n+HohPBAHTvR4lKFBc
cqEOBzG4S7cjgqQ6Ib5krasTOLmx1HmPWIhnQvKU4ERqgL8jnaMMo4/WvUshiIhZ9Dm+J+Q4zpJo
QRx0rqRWWH71zINKT1ZLcDTPH/h3Vip88nzfU+am0IbiEmXMHQzsdZKmPJFuAn2hc/UaggBRxD5H
1h2H07m99mn+pkuLVcdjIzP9RruR6kjAdcZUtXeqt0HthqucacpdAPGKKRnLgSCpcaqJ/PGzvoaS
8PdZawGlEkkagPjesMNIK4PJ0KsiQBDCb1c+FYEBjloxKXe5bzGuT98Ow4xLT0jWgRNYimkipEt9
AxIHyZPp+BF60s0V/DkVrUNzZIRLYc/70cZN8lSQPuLau2C/mHkWOM2b+xLuw7Rw1v7UQQD30yYk
SXxLRrT/PF8vfWm4vgS7zomznNELzOcz7d3Pux8Zm8SnvFpoIHV1g2x4Bd+cHeIwAXZHBrP2qVx5
UnUDAGTVtOHwsrh5uXkDrAcIpYICHiL9T5GLz9hGfCQRaRivqeE48u00/n2WbY9hzR02VHcW3wJ3
RNrgzNlMFWGtSSzgRBWQ97rHnOua8uGtGlTfuCZAIDzxoRQzY8smnoktrjW+RKiYZ8au2elaoW87
v+v1nMSfXqKKKjlXEkmzs03uZIRCleRKoPnzjjOGhVpI2Xzujwg1HOz0VFadWahveyibYdupu63C
v01rIDAH/04VnzMaYFK5V5d/jKqIzBmfzA7GnGVRwbIpxkyVssfYevIF3zj4y9hqOn/HE4L7KeRk
5Z1w9sSf6x0c97E70UHEXYNaCV+NmhpAjkDMT9SbPUPlbHyl/u92ct5/dBinG7QBXK4Q7TpRpZ8Y
HEL27GDgDjAHFABmX8f9xjNIGaToT6fB5d64yBtf+luvp2wK8Ttl1bcy0IlaTEQUCIAI8NC2RaZA
+9m2S+DUeMHdqhw00mYZI3j9k2VCjRTxAjXAOw0slqRe+xkwrjHL4xuBdWFa5Dyzvi/yC5xILnEy
BLtRKgBByotgcobv4HbK8g2YE6gmjz0Amss5olXHoIvI6PV4vmaves6K+nWuMw6EMVbXhDtApqmd
Kem5fSn+sMaXJTT7xNMx9VIeT2to3iuLbvTiqTGXWWdascY0vZW4fupPJhBKZtuffSvMfIlwOSFl
AJE8T+36b0co3mV+4xu3sQi5RTT8Bf37OXxyelTmx7UTJ4DJgmk0aYvWKRf0DEeyOueaImK27SxN
qslO1GjXHiicdlgmjgziTwqZZsKbnX2e1hnRLGb9r3Q0LsIJJA5LOyZONXdNcW1Zr+kU4fxD2nMq
1NQWx7NQ/MagdWfsuj4fDDuUlmF/eDdtirZWPG7kGTO+Glc19+0g6V3et3/wqH9LaubKU0wHc4P0
qsidsQSV5Jo+7H6wi+rEebpLZrx5h0UjI96cUYe3mCogsJcXWtw59qAHp5sF6oWYnuun8jVX07Rd
tPVuR6DyuUegA8S6uR09K+QoTumgSgEZO1bjaTynT1Vc+hCVLbRpHtlU+KIl2MtF6cBxqj9NalvU
OOeyHLmtrQoZ1uk5UECSsrc8iXUUDkNe0GmFW1ES4h/ocUx2tAOeEoz99yW7Hr/1MDkWLf4JhHpP
GmH0iTxeJTv2gHxem1D4bkAQmdsZaaTY/JDxsmXcNe2zFPq2456QMIlLnNQZgoBBWABRnDXXNzvo
ihL+PcYkbgtmBv+Jt5C64r4+2bGv2B1L8+h9rK0hiicLVjyLr54stTSNmqWFicoGSlwWtC8nl4+H
agJ3rwdp1r1lDY54Rln4VbmyLJCDUtJhTeNWPXTh2Z1U96k3BTeKIEA5zE2Q4Bzpy5/yOLHn6yUw
fPvJJ+Hwyh/FB17D9jYpBUs5+jwuGFMFfUZVS4lf72FXwjW9R/h678D132W0HMYAlPfocz2K7vOm
wGVBrTuxeA/jnKFsRvFst7SW3UJYNOOkbnhyrJ2r8+VldzkTbOxnGMOmpt5ufpcDNAugVA5/PwOT
3BwEG1NdNQvgCgrb6a43vcMOyVmB4Qab0ibml/cuVfotPunnOxkLyqs6052SUG/8Wj9NSGZd+RQW
nqMOWevksei/rDgXFRz1Csx8jZpyZ7RTwJbeYCM/R7aHoEe/iYDoyKPAyGbTJkeLLPm8j+eKg0C1
aMsjxIIE+ukF6DGH2Umr6Vo4nhjTcFsp/yVc5MKz+JtTCBLxQOMecHvnURlj6qdD3nfMBK746Lxw
cHJ4lMLcHFavLYl/NZoTPWQ0tObrqMyRZoCA8oW3EkwpUh/3u2OqGHkuSF3h9Kl8na0z0bApaArX
dgYpmAGqbcR0AWdA+bauncfrGwODnj0+7P1ZS2FRnjXYjBnDN8vXsWOuw5++9L3AY8etA7HftuGP
mN6tMUZtFMesRmmgfYlggownIPXg9FZHND1AqcY6Co7ghlqyJQP6qNj98eeInriSuQ+3OC9eJkVa
PVhaCefb1HCS24CYmNZf1WLF1+rjurNrCKSHxHR4/uDCHq9SOY56s6/tIED0O4eTL0ZWHkfw9ZKi
CKYSgzROK8FD4XKTxW0BuCm35699WbCv78VWNUveDXvk8f6Pvr4sVW2fQr0BqUmrzvlU1jypFj70
+4p3yWntHPaAd5/YjmEG/1ve8RCSnSC0hDodJEh1dYSJ0W5zJua/mLhQeFRrvCywr5eAo4hHexc9
nvLga+9hBg66OPPVgIZDtu/fi+r0jMxS3F0nLhJalvbkIDLb1smdZMs0ijQUfhAE9ZQ0UJr4Ea7e
U+aESJDQ4mwdntBiZrjDa+EmnyML1GtUdwOG5SdSC092f2n054SUoPu92q6E/5VDYIXEdsl3DBIy
VVtdUV3mQSal2GIHXGeKSDWRBBkRZIxuw4F7Upg30a6P6Ex5jt6Deh7gz2eNnjoMKcef10dN1owR
Mx45o6N+lgYI8Rjc4uaM6QiS45wbn6EVWKVSRV6FVccEI5jgsg5xUuWkq4FculxidyF11HBDMoEW
tI0cEd3HZ+AmJ7ywJL2GPywt/rDcDlTy2RyPT5rlWUv8xrmoensYl+wQbSygwVt156JpAf59EHCb
e3qtE1Bn/4ZnD4SCArrfSOcQQr90WV+aOhETa96GyxQzzQpkMvHZ4/xa30mHEBBwhAzALKGD1O2P
XooKyRnErj9ipdc1LaJHo3qjspty7+dBDEQVFSfkkRxdo03vM8nZCTdPDEy2nyobCAIzysPQzvSx
zwToyFfajAVwjfEWNu902xeXrTr3Sesg66M5i7OVNlB/9B2J9O6ryvt5pf9fIBfKVTea7tHn+sWS
RJ4un8Aywa8DXIt45SI6TMhQEwlG6EFNwNnm7ASOohbiTcObAYtqNLc7Q/IeY8ge65BcNFIIpquW
ETKMbZWUCN6lDWgzgp07A0rXQ/kCNgxSA3ZDsV68Hjphov2bFtQGS5V4wIIZPhbGyYq7JuWILF7O
aseRbgTv9aLAV7MeZaVja1q+CtQoWi+BfXv6vqBnJOML8gIV8mP9rlXEE9N2rkur2JO/XOZWnAOP
am99yL6TuuxxAsSEtrOqAKoGUoRXQC646Gbx7Eozcd3NHBW9KFR+JTeLrZWsrRwUwfXF+xQzAm1g
IvoUNAKbkkeDzFii5/pA+F+1Fh1FQbGT/rp1XzyHdMB3Og3FD1ve+Wab/UhUiCo3XVUomGPk3lus
rbXsZUIb9LJ1YfrAYu2nB91r1ba/jbkKmvsYHMYwZbSi6hWiFgHltDE6X2HrUKQgdCKMePF4fglM
ZoD/1Wu4mvL0LbG1tYp6ORZluvHfFvnIYd0CuFbYYiAhs8GL0Pbvz6sULkccc7pRYneTqIo3yIgP
sBDaKApLDw/QdtDFQV+qFGf+TrXpmh2Qm4niQ2u/2OyfSTb6wa/ELvRQfoa4KbpxxxIJuPmYDjzR
2F4nqMXcYJqlOeDvx4/LAWkbpD6lNmYmrhLqgQLPqlDLrmBeCrOXeNv38o9EcsIFil+LcJrukwtE
fnk0q4O4ID2GrkEbuawRwnToCU0t+WLs3KiaR8zY5MFglHNJCrOtwolCvxkSUcNEp180lqH678Uu
2Vbge1p3M4DxK0ZTbOkUWOAxXLg7PN93Q3Hp0r/he5+CA310w44ZqB8PSYI0lW+G7E+ydgnCkggp
dDjjKAS0DTljvh7GNa231oquySouI6vYToIENOftc5Y3lKSxzUAuOWQCC3BqOzXrge/ufOyKqdhX
e28otwUK8f9PdAqGN16+0I/Wu0O06V7wuliNMfus3kklGzfz9apullBsxPOAwrI07jm1F4LJQ2RN
XTy8lL7/IKrNS8o0jN24gbnC9VbEWlGV7xWkRJDPOONIDUCwLOzO5VlxqL1hsaFSGAC+E8q6rqph
wTTzBGMHC4qVjWoMwqOwQpkBcmvjQuNmgerteBwbfK32NF2j0Uxgh0aBvsTQ9G6bR48o9zVDoVty
NBUa4QXNLiI9D8AJIYpNFNcURlPpBoSzXzIoOaFpYaivuU6lRgl5TZfTPm+Ph8k3RyGFgAF/Ge4n
ZgRWc3w14NkUCjSPlMY3qKbax8lWA7w5wygwigV/jezt+0yfzwQK5QRJDJNsEv1Pw7JQ6yIPyQ2f
mc5ag1pFRLh+f++GpwYRh6WI7RVrS+aJ3kCEaWfBzCPuupp310jlHcKM5vKijzInhK7yHjGXItsm
TGTviQzCCNKCkpzFyRnPhgRcZ14J7ew2car8vyFDeKqNagSsdzVOL7uo6sysw+YxM/w8tGHQmAEC
VBNILlkWbOfEwgHpcc6OLqENTT392DS0V9Id5nFKkRuOmohDhBqCrWilIpfDM1eBqOPtX0sJTz3u
mKMdkuZUasZJK/AMuMcoUB+RugSE3iBkWPs4n0yKvERxSUh3HTXVpYmiPavDoVIDpAqjYiMReN+4
5FNL42tIdsRUkP4lZ6OroWjDFrB/vwnVZjsm/WXUCABUXYiGAkhCaCyrnMYsypSAHXIAdehSW4G1
TnDpxExwbQ3jHd60kfodwOYejNCmdnxaBX/KNr0gX2mnTZ9SOyYXy+YfZaMwx9Fr44cDs/E/xcxA
MiErE/9L2vn8wGLtpC+Mb2fsQCY/FcKYHyqZKNgVFu3OCu4AhBsNuEXzbJ15KPgFizFw3VA3RYzG
LL1Hsi8GSVddEDyQ1hCaTgQOG/5d2NePLyqGcWu3utP4L3akbUR06kcXyNgM23HvXE588MgVPF++
GrxTU7+Uve6T7lH3RzhAPyHYJwGaMRjXmovt31kqBaxhlw2ivfk6rcFslfNeuyzC1ueYCN619RZl
bXzM2BHv1axixg5xhCUlDSbqbeNznkTfgyJQ5t9amMdPJvgC6UHfxONB9smkGYcwprs+YsmcYgTD
1/jXypZuFqK0E4WWmbucRPv51hdpM85IXyjosQO3iFNP/11sEWiG8I4AGG8iTeS55sBPLrgodhCA
Lb+eG81jjoCISSNaco4DKkam4puCWcKPCYTUKYaGJS1lFbxQIK+nI6s/vL5VpBV83ZLVgsMup2ee
+83eqFUuO6cOo+iff0QpI9IIBCd1hJh5hDgquDABHmPakB87s7/8kWQnHwa5FDg8Hgn4tlCDlaEu
O8Z4GeroPt/XWm2Xy6UsI2EJu/pwUu6rt6hDa4wfiFI4z4siyESXVACA02tz+0InAN1ytAIxBdcd
RT+BFbB2iGC9oXU0HUJVa1X/BOXTKB2VJ5KI9mqOS8g/BZJQ7eyfdFHuw2yqDq+PfWcOySYfcBQ/
iwmX/NW+CrrPdp3+/WSl445vvnL0wVztGjOwKxrrt41ViasC0V2lH9tcqLKCaWdxN/k8CrdqyX8j
K3dhY/6Mg65DzCTjX3PcP7qE9NR/jkNMTShnkcoHavk6nEgSmz8B7KEhRgcKiiXqQMrz9rrPes7f
y0+Ncug/yHIxSnwOdEOT08rzO4MBghsgWieRlMkM4bnZbswvYMR/Z025WN89IUBMoV5aljV+pydH
86shvX0OYyXsZcShfFQNQHoI4zlIH/+258igcqz4Bxm0rwAqyKokpXNpkELpUcn3wzVJKHZGk6Ui
49cUo3zURuH0THRYizJPser39z0kfzjc7mM+2GLB4ffCEHgIcU0ymVU6fqIluPuMJNbNvbCyfzOZ
c8oxJkmGxrImJV0eMFUu2N5IfZ+c2DaR04u1Ay55kPBM5NwzDldwxJes6Hprd1Y8qVz0UxwH/Bds
Nqh6ZtX9hRWCRXM6H8LleVXCaNV7wEjOgFmbUc2aYerz9908bbC8ywQde+N3HCSKs02trnlyP1UD
Qx5xem47FLhgMSBbE4i4QQqrSViG8ZPEMCcxy3j3NGT2p1FFTCf4Nlf8Njt8sb6w4we6YCntDLj8
wJfgpU/IK/QK8++BHOYgOoN5QXBPK5FY7SmX7L/lGmasMNVYcOSFK+lPWslat/XpHw6GdXC5WuKJ
usdKUZYr63u9pQMJoyMt2YEJjxc0s+/XAEa0TEZjKQe87nn13hpaLrbSjL5h7JNNHxhFyg7Hi2xN
tNDLDsOwMp84lHZipnDHcKgIDDsT5ZMpus1jQFfJGeanj7f9hngdjYbKHrUw7Z1QF2DEf7pELCPW
6HAwcmEfASVEHI+ab30DS1fRZSY9JAp8ynqT17hK3zZcVLFFgyHzgZe7Zgpgymubw8/Z/7Bw1PLa
Ph6tCyorbYNdPVPHGTY+phiPs1isOriKcGPeCWmCHJEqIcBgK3YXhXTdvI6GADr+zwZT8UEsQG9C
FyMj9dXd4RiJbALGAy8zrakBP5d7RBGcVQkPVqZ8IOeGR58hMMlaeglRvMttUbNM1M3UI5PnlFc1
uNEn+hQXM7qVy1Nx+0P4szCg6zkjJF1cHeB31E8BW0aPhpBfa+LfAedWYmB5bnKmbjQpO1s4fg6k
UABaeDsIyzmv8eAccCSy+AHI0uIGhtMuorHXNyOwuFOB1fYG2ImdLuB/XSl7CK+QWQiJtAnaeN9h
qn0+eMpWw36QorfPVmAI6WKWfsKkCtuoqo7YA7bEFApkBd3cFROLHMp+6n7M/4cXQzKsOhkO8n/L
oNBmJXUqvyzUKtJ5P4dr5QULYQT2d7TzaLNu3EuLmRMUSCW6+N5KXHmQ2efI14yJsuI3b7Ui+ju9
fxl3qkZR968ZO7qIp01B6SAIVNpftWrGCfqpWKYDAPv589P8iImuy/3DbsDUGIyF/pt9pcYJXjz7
ilHsezXiPrNzgTi4uhkUrQ3ZiO9C9e+SeHfTovai+s5yV94TkY2X/jh3yXhmOlMS6YPVuB0IWoJf
2eDczRG750SQ3qKfEYjRKdOgKJGariLo8gfi1uxqcZgQckmUQO5zctdeBhdPKikiIdE2ypCwzhZX
zkW19AbRThzyxKUKtFKMCfD8Lwbc2huI2UtRx1m3ijOTsAXQNrT9WxIRR7wcvtpN7ZyCbFdVG9CR
h8UhQ+Hrh/16j6wOwLtRV0ubHDLgD9dc8n0mz3wUc21rZ8M7ZRZ36ZjDO3vx4OvuoRFc/OTWIkUB
9H4BohKxjJQ3IWhk8whF41HK6s2B3GtlvOTqBpYpz6s06V9JsGv14BlOL92Uo5iCSnB7nx1TW1Lj
BbETsO5x8pK7a3zKEWE+xIv+OwpbKEBDRJAIZo1Y1Sjk8t03BYkydnXIKGXpPH9+mAk+DF5teiCT
MDiyDFQ2YAWKlRL0jTaMnifjgHzs6sjwFokYIoeA+K37Bth+LaYV4mx4y+gOonUiLXA+7axrjxtK
0qxxMpyx1UF50cAL0LwXPubw/3gM1y863bLAx27u3z4Rxvimp0N3qIhHsG5f+2t1wJAvI8rBDhfD
BkJq0OvJNedIms/gAA4YNmwzamVU9xIAwkl2UZD55ylr79PitwCcIoXEWxyfeF3mjMpXdlILYGJf
qTxh7akxdMVrUGWNNj973hL158X/7dWonXpbanJdt90Pn69LCFbY+8WUcue8x05+rDRaWm7G5Ojk
O9xsDU1uGXr8+YVmcaGVZzzPoXQxyxy2l3gAl66m0KeiS21DPjRuZqrn9HHZ/wRgzzO5tGxph/7o
9xXcYtYuDb2W6XYwfgLA10jmESuXBOMXVS5B3EmUZKMjDcTbHgMWIgjNxcuZmhgzcmmNbrlMxuAo
ET2m+uXtI6/l27HDoESmhpAgroRR+ABkaDA/rmhq3jH9F877omBB40J+SboxjIeHQX7T4pjWX6v6
aPeMEnIvkQo2m10ACDPavxfG0W7PWjsDkJKucXXqil8FuugCbGLjzI1HW0W51XIvGe9LXcPdACIG
lEJEKNm+Bs35Rkq76UU4ksZfRFnxNeo/dgEe3bflgCv6IihSnv+zElA+jMPG9zm0zZ1atwfQAMFI
8ok+meqmImPdv8xAVRCuM2QYbjT75+WtedyclBHWqgeb9MXc6Js8fd68mJsLGAQ/kE1XARgg80Ku
B872BltrU7rec2L4ItPcAnfWLrqMw6lI7i7KALYG5XSBLc86ePUD494qDxfZZb9+WLgHEv8Qqv7J
cc3+oy/YOg8oKF7RMF5tdoUeLk5xp8fZ4Me1ZT/6EiBchhD3HVVPuK2+c+Fsx1URLxttqFJ4w64k
H/L5bNfW6AB9JtsADL77Cm1GPbSDp4jmaZcChQYxvR2H20j0wuw1J4kTDw/2eDsXd1qYar5GuPWh
lo0SuQzwfs50caT+DVh4QbU5cPtu6ppGb4lqMr4zbN7CEb//1Pzuy17QTpwWl/aNkxUY4nbKMHUs
YhMKur2wULb9hvKZ7RIMyC281RuLy+pDr9v+OHvlYaB37pXSRhkMVJyV64MzqLrr/l0c6NF881EE
vCOvehoJuzGNPQZUibGcodGxFMCLHG8l2LTSCAfZfHsfzbY9j7LPNutare0kq3dN98aToofMatS6
GKis8ZmRirIYRWsiADnXkAHEYFjgpvKZw+4DNq6dO0MuzOI8l08nIZkK1g8bYVgAVQT9R5QeLMSr
wt7bIpImCK1ZBmZKijwj4vigAgOFl84bcTpyP9dvK2gym6h2qHysByu1FNBstK1lKMg9M7da9hA7
svwozYwOBDAtTIvg95hsot0/Vo2DCIIO75lHkwh/sy5XHph7fItkkIKmKwYb7hbcQPqN9Zxpv0cc
495zHQkQ5gPI8EwGp66sex9nLfM6Uxz6oY3/pm8BQldVMu9/X9+3O3TaaKF4htuoXET2irHvSrfR
cxpK31H9aqkYKq+Rvx9+Yg+vrmkxcBqVWtZ2quwHKe04EMeNdiz8p9PEXl2JUW7g4GAJTIMkApBx
Kf1xrrCSa9gFL3wJriJUZulkZ4JwJe6n+zoN19VJaWE/3oZuZ09Zqzu22a8AMc9w+0qVjxoikhEd
HHZXitAny+MuxUuMSwf0Pm103k5mZmNgszWdG6LdWKrs0llelNm6UDzC+hSzj9OgzegzGP3OET2h
NwUcAmfXFUreoO2wBJGfk4MtYw7WUPVYAyA/oLgjna32eng7+mV29tA74vKp5zwTL5I2UcoMD9Fa
sMMnfc5F2OmjNjnlpSFImYHggQLDuX4vSWpO6Fjzclg93HE28ff+F25xDy4YmsBwYvrvLe8ljUL1
vbAz9p/I0TYLrml2BuvZaOa5QXrWRfhrQ4ZcetvWcPXqppmrBcKGiW9YUR/ZfZlbFmFukN9o/QlK
M60da0OBWB0LKCWg5QAwQ+xUgfKWNnIXTwF1rNIQRiqLDnuTRJavyKIV0JezhG7G/juM9+5Bs4xF
w3OdKD0nVP3CKuMIBt6zIG05afNn1uU/b60/YqJS39PCoBgtYDd46d9WCTGyr0TNPMA07353e1KV
3iqRIzodhepkp/08WM9WzA0Svs3HeceysKwTkhaMGtkhtwYkrf+WEKoj+hA9cS8qHv7Z/Li+CWr7
ECAL2Lgry1iz0oLjEAwGY1gCdXzGCpTA7KHJxzNY5WzO1Qd8wBkznT2s8Rx09oKASgACwr1xeZrc
F4sKDcGP0LPJ//Cvi3AwJEMXIY2sewnlIOKT9ldJ85BBXd9lh2X52iN9jxggIvBB3E7PvnY0zLDT
GCHk03W5TEcDhAb8QkgXmVxjDeB+q/33J/l7s+Y787x4wQsNJlcL3/AMCQk1VAr7G+ZxoEuVWrwe
52fZ1O1SWifrT9XQR6QDY+9lW1J6iVoVQXDjzzxvyi65hTIReW80xycgLCQkd3B+89sySZEPN/0o
sDMJXPIiOe6WsK7cIMlRP119l1o3BSJErf873V3F5hdjztI02nXjYnhMQ+oeys+EnCila2w6HOOp
h4F51R5Uh9IkK+78dTwf1/KmahPARdAScAWXY3ebbyVq07zt0qfGsznM5hR21DUt4BZwf8xsRfZ5
qyTFUP3Cgh4xjRTS4u9Pfd7FKePO9xB1zjCdF/0GerQeWeF4V8hMDmCXzCxzMwT3suV9MzhyKIDz
sXQKnLVdJfzYUZG2GXqxozLAuRFBuhFaHvlo+rp3ClMTUo+xgla+Mr6AvDDp008cLyn9szO/7ptO
euv41W1hDcw/d4/NkmG11aN1lmFNgM2DXZSdU4n1CFwnX/w1I65BkBz5WTXK7HbOsjMygAJ9Of8f
VaJRtY/5q274dcxB+zTA0/BVJYrC4ZuksIZ9wC7Z04BsOWMFpqkC5aIz66cw6PjqTPhP1KQqdlhd
o18jN9M5Z3V6YOlTuZSBNLXSN6R2B74+zlKiY08j+Y57LqaQPF8RRxOw0VKMim2IigpAiHXRIjih
WUvjTMr/2N/uecXaxcNeWLhSHajonuxSr3o1HFFs5Cke6WCS24Uzd9shat4/b8/RnDTBlhdYpMCy
DnARQ7fLb3TUd2AV/ePMDj7wuoINYxtExicNVPBvHkTQzveppBMVWzbnPeZsIPzfhwkDdoZrJtDY
8eqdJJJeSo6CUlh+8NEVC7+50ZSFnVK2yZMqAkB+o308+nY7mJz9htJxXX7NtuwgqiD+hsgGMGsE
NWGch4cxRUDgXcJT+XWL5f6E6wrEIOuQMjhYywg0xgWhVj0QobSY4+WpETSj7Osel53h2jW3mgEb
r219eRaY3Y3CvhaSHciODV5EmYiPkLkvBDMxVNwE31ga+dJvvjHBcmknwtMCEThqVkcdzfAUWFg6
x/SUExnVoxMA2F51LMWY7GafqfZSFEoFlObMEBA9Ej0XUfp5EFeIypal6wV5vlvFj7KU/JjPaQ0o
+EDqEnqcegbQckaIVunedt/8o4uu/PdTIkmkOjUy78ARasyiMCq/rNdPkbblFEShAoFbXHSkyHSG
GvFAW00cFQoAuB3Je7fg5m6VrNAmm632XLs23brkJ4Ja6XHdR4XRsIPzFXiQechuGiLi4z6Cg7Q1
wHGezGIspJiIzS+FuH8rNDYmJ7fEUBPPiKb0ArabyD62Yd5mOcaI98HdC19K8cGL90ajkw7zDA+Q
IHc8LRMAHYJGi+QrdwkLjb6v6WiBDqZ5mt/rFKR3HIVkTF69degSDtmhnGSnsUdCisMZkemUVffK
sKuRSh0q+LOJSYP/6IqJGmxpemtFoptWok1wybwRGo/dPN5sprzWoShECfK7ClmIrx1ecMENHBL/
+5oVJkOOhHTshWwKx5tnnGM53wD88sY1T4iQg5qdSEYmTxOvvZeys3gZ8IpxiDHxBKu3/xgOt5q0
vbCKnGwwu72efgX98fXY/pdoziVvU78YmjjhESSmkdCufjgj4wd1qXWnE8AGjXzVWHysAL9jYV9w
GWfYiuGGTUaLZrevcWfR7/lzMoE/WlmB9qwq4myDDJLWbm1TwCAGov/0pVdImTdSq0ExgmQ6LcYO
Dr+M/r1soC3U4G/GLGItvnPPaYf2zYsq6hQwAl+7Dn+Xto0k3TcOurlMr7//8ns/JavRvZc568wK
U3kT5CReRptHZrUDCkqmPy02qUrrBkgSUciDP9iabBmClb4Y8/EPEm0PfAM2MzyluHR+3Y5DBgya
TcG0Co48EW6KnsA+08TBauF9lgFVnq0PdzVPfosr6YEMPw9U9Msr5cjg3tXT0UmY5VN0lrLiuSSI
Na9LVYHwBhwIMXzmPhkHNdj88ZZbSCfZyPeBftagcIZljM/wdeuUA9cShb8PbdWlBvMNuzkb87Zs
pCL28OUofrfimpNeIyNpzGrgRqOItMTxaY4nNKu7OTBw29xLjaV9NsprNOrsiym/AyIMVRFDBccy
SquZGLkU+fiMT/iS+3/dI5gmST3PWRCEzshivLT9Zh4b59zlPxwgp7uy2NVjZK6hG7MPMZ9aRgUo
EGugqpsFTVK5SRqbnfuOP3neb4Nvi64B8zMarQ1pGgI05K2ecW08Jq8o67A1Zv56MTxUTOq92IbQ
vypMQVhIlDkNS8fjOmu6C2iHdarit3uI+KvYYy14mqg9IfTnhoLketMYv64mIEm/5o/geXrX1Lvm
JEoygAm1ioIqV987Mc5xYHLbSH+loYs2V0jrDUvTDxF2MP7V4aA/zqB3iSnVa27nUG7e2u1ockON
TeIEw8wW8tTPxulCDNGZFpMp0TLVztB7bGrGP9dVY5JwGv/IvaughFVVovzbivldT+h0r9fipOL0
uHxAOXEzdjepEElpFCbfgiXiGdBov3S4WZgM2sRVdPnV++7Wp4k3q1C5snxzm3zApUKUKcX3tzqm
QHKoRZE8flMvWHJ+1qKMUUi3QJvvky3e6A5UfnPCP6uNZ2N4tGVfg20iwzaPr2eFbcGbiknZGXg+
cGiEMq9DKqRVsibxwHFAp4JGPJbkg0IvnWgOo+G1As/QchlHmW0zLve5YsSvgfb5rfpaRo+xyzJ0
enBXWY4EbqzhYMBsZWP6xsI2uMNdzMqs6M7wujD32C3anJu7rKK3rRGsVI2e+Lhmd8pG+hXA6gSb
nfIPNPw7fIR3iOOijKYua6HlJaGR0mcIfEfvkNHXEg4Yr/9LCDvDQyMNFywl+L60mCVDpSCtnrUl
S+UQKuT39l9u+MmIZDFFWgyIZBYoGh6GLFi0T6zr5pex874MvZxS+PyPSPtXXn5xxXubMLrqk6Ri
7H0PLQu4ivhwhomQnAVN6OPE3/F3IWxWT6M7/oWt9uajte/bBZVV4G8aHEkwZbp1HF4+pzClLd2F
68LwEDwd9w1LlHlOeUq8h1QzZ2oh7A56f4pQ7ZqA8IymnMTgpG4A/1VYMPSUWSxMJ4xQ3/dByQzP
JoZfkopuKwenF8JEREqjuIngKeh/lsH+C4f+kC+te1dIBUKFSt0AP4aLJsg9s6qGgW7eKfKXNMLI
ExJ9wt7oa4SNMrtlpm3IycmTD1jnB4hwLSPzSKGkSX42jxdCOwBQGIhgcErvqna/SepLe4GMNdJJ
iG62SPsR+alfLd3t0wmf5Wqoej0Bae1/SNZ8v2eDQ1d16hwPLAH0KYUgooydbC7S2sIrumTi4yNY
F7e15qdj8ge5EB4LEVCczoQax0shFG7XA8eAYtMrW40XfqEr0niHXSAIRnbSaJqthHkzDrKNsTCS
llSNVFGmNpNKGyhzRXEApKNBFDq8XtDQUeMtTjRZFgLi0kNYZPQB790HDmLOCAAg/8IGh4nqlS5Z
nQ2/Xbmybmiz4+lXfFS+YJfJMVwWbvqkH87w9Xo8RrSvhA5zTN1HEeXQtewAUX4xgx9EAN2nieit
EUgAc7XRfcINVAxTFQe9e+Gv9/qdOAVIct2ZUhNKbKJkh1ic8NrpJobvHuw51wknHtFG7mOg+8/a
FRZ0HHn0IG7tO8CsYAs8bBhib0r1E9QMmw1tnz+ODMKThd6hy27VrCEDD6s7fBQogLxpJ2spkagZ
PQjdnBCX3BQiS0IuaGP5odIhpDJeCsuI4S93YAx8jvkOEFmoj8YAuupfOzlBQRfNwKuu9EaS7+yB
9YFWUYcDTXOWo33bo13JFSEnwqx2t1gR83Wy7qL5ZdYCi3fgzvOeUVn9RsMGgDpSKKMFsb/olbRL
QyUiXBTNJSiUzsvA14rH7+5H+M7S4jaS6rL8WnztJqT3lO+aZJ0yDtWJ5pgLnk1XhNCtJyVVjf8s
AOIZrr7hY4R8Fufx3VkfoGZIZRXA/1mRC8U17eTivARpyPKxoCXoGAZ40ka5V7Zs4qC8I9psS6rM
aU1K6Go8V9Tt9ApyAyLkU4JcsFOvQ40nX+Hl3Mn0YQ7AeqITCmf+3qZsf/VG0QsuQEt0noWosoOF
6jQ/CHBmeHWuue66zISpBox/32gOx04WCVCK0rkmw1HZN127COMFztRYbk3RbfcCRLDxsSfAZhuk
czBI6MWIEAAuafNbxyNVJXq5jyMxwo7a6yUNkOfg8Sflsp4RUQmbCiT46DVIu63O0svWD6aY52kO
8fljqJeq8l/pF1pqXyagJJhHsIrveRR4zAhG7DkLEQyB7awRzNZxcC4yHNe8fIeJhPmZUDm3lHWC
SAgEahKA0gayZdK+0Qc7Ivxo4rqtQb5/oyNkkZJ7n4jNeqfmkuHQw4wXCr/zXJT53ggnob2mt6SN
zZVgYxy9zNy2t9UmNL+sr91EU9vfBOgMFsFAa6bGVCkC4UVF3E8Mm1FG6ww3Yg4dCbwb/Z20lfpE
e2I6a0dNB6BDc2C3AQYIqWW/8HnwjXAcoE+bRpTWNECfoWLeYDENIOiV+IsAQO1fZkyBsn54zkVR
1IIYaKj8eMewIlj8n80z2f3kXc7LOLvMAWtrYAe26a3y3qPzu69h6omdtAixB0ptuTBrvLFtBl3Z
niTn4TfjAKwD//UPKdH+bD+JvfvfnZcykpf00S0YtjwM1pfHw/2mkZiQoc49EVqC3TS999yQgzcd
qtWHfB294xBNE6IsnFasRsRlDh4foovvKIC9bm4ucZSr7+4zcocZZ35xt4uySaXVNJP8t3P5ZnsI
ORtnwcaG3563Sz4xVKlaTQkePZT/xmKEtzuGxmhk/LGCgaFYtEXRkJ/TJv6jPDAhNq8TbaaTk8qV
uCOIuOeOR1I8WFc3b0h8ybgkpG6aT2YVLAj1p505uTiB7bw4DkOQAsMfeUjK3NME3B5HoLS2P5sb
7yxmv0OV7NlGlhgOK/ufDaB6kwJEpAT5j6LwrYbqYvv6BjF6ZtUpkMBTAxyB+3bkFWIM6tpO7Y8Y
TY6B0KtOEGU9ObWp0nvn7z7IPpowD8clmCb+NQo6t53UrUNw/bOZBcv+ZG60MnDSF479RdWgy+UD
oH05pDZOsSVTP9wuWCc9FNhJkBVp+iD4Yr7x5kzxhuwzOoZgrswqva1x9ZVUhZDOGqc2YUX6FFls
3qX0gRvSUsjJT/w1WOA+5ApzxrrRKqTUsCmRSn28z8YyOmfdzpKEqRfJfduNLeB3UuO/epg1PJB3
2EHYjuYRYQMF9HdalCmrFWnrxNfTYUrlzsFBM/aZEbQZigViOG2yHWsKve+75umRRE1+8Tv90G5L
u/mhPWaKmtzkXJeGFIdNIRgOtjQQjEeAxnAKKEfqzEWxDEGPcRVSrhKXl1xTwn5B722S0NAY2Li1
iy5aTYGm/opUU8+xSVfyad42ucEqLx1LzEG+VU0Lm98b5LMNEldkiNmh94WN/FlLQRROAhMQYCdU
xiVuHOD23ovOk6yIFNb5vUGXwYJYsRSkDwbsd5ROm0zqADGZqTFsncHQxEKck1l59pGcKOV9RLiZ
W7vikKy565mT9vzW30uBeuFDMRqx5L5nPEsgb2kPa1BnxfbMeQGPUIvaSsjh0CSzpknhgxzkoa0b
K71Fk8Qam9LqylAWVT9tao/tBjC4zRsVKHuzWnoSRpyNOE7k6t79atBD9cgOL6gNpvR9RY4zuj+l
KovSNO/zXWOx+fjfV9lLRD/6POQNB/A1RUsXuDhwYCvBeRAFQagUqp9zBN4dQWg/1vQoE0DucpP3
PL40R8dUFDHOyxaAu5728deQ+ZuR0CwqLr90mGkDFL/Ru/lzV9pzjov15jX1ZG1LIGrUfxZnSn7/
bgTNUeI5NCH8UjDXm5fYHlhupL7+5aO9CkOZVC+/XWwFJm0BAHorLJ+uFFBQxb6i5o9tZXeSKHhp
oFOh013n1efyYH6GX6QgDPJdIJrWj1DrsluUs6NP6vrWYSigt3ifDrAe/9SY9awJSDC3wP8NUNcx
ZlFgyiWE7iecn5LMIvejZrmFbvMP9P1dSF66uyZmM2DWhsKgwe+wYN8v4lIXHNz/aTKQDyukCKrz
joW3UUyF3NGeZ6EaAW1z7PF3+HQGtqaStwLWWOXEIu1vTkwL8suZ4pNSW4DrJU/2ajCLbAfJwdOO
6L2CwyjnBekETAGyT9+HQ5S5IqGoLysJUIY6fTenxOhhaDs2VG/yqb0Tf0h1JI1aiShAHew9saXs
mmp5t2ujv2V+vD37foORS90FKRQvTbqgbP45Cj5phf2KbOrCrmQfdmXsE15JF2uNJnQ3EFcqeZ2t
tI3JoRwa+Fgz7Xfi/u5lXYT9I2QD2WNRe4Hxs8yEJGZQDG7anZGX9QJ/wWwPbeb+8smaJ50QuKGt
tPBzwvBgdIKyRQ82Guex0WQnThmRDJ3AQygvpw0Evcqt3CnV4GYuSqzWby39qL6YLkV4JjaY3wtV
LE7UQvLrEj/FG10oFgzJbPjhm/9KuVAbD5FUwnNTFi2940c7X+btUtXUOcfsaoIJLxpHFu8/PEeu
j5P73+ZCxB4dNEFMCxHzne3hFx8c10ypT3H48fdNzT+pXEGpQ1gkY4U53uOLPzRKZCjU0HFVyEoi
qR5XFMlWcVOj1tjhoLlIRIKFpQjz8cqHNI6nJ1rY6hY4xkxcxSOBUJ4hMtiDxJZCj9B0Ha3Azwbr
QCZ7ohd7Uls5+KEcKP9c/ZBbM+PkVNLdgilEePCSqxLIeEC/IIhA+j6RXgS/a7lA+bUSBZzAACeT
hkoSO4saJ4nf4CFCMgR34HuGbE9XkV4A6OdFCuzO59zT0SsFCWSnNRqqm4T75Le48AVErgD4YZth
+mtzXft9NeUwPlBPgtLvCkgzt0z2cMHHeaxJYxfhJNu19cP8OkWZEDtM6sgT3qe+sGIR2oipp/OK
vFf6Q2yGppAJPyw1XzPwJsbp823ZB//08olCQr1PX4gl9GFguEv/qmfK1yI58/v4kRxuC4WoOSH8
Cy2a5xiC/N+yeaxyyS5USJJitd+HQHi6sbxJwEhUEDYadXXYgvAdwTbioijUeMharGa8VfKeQo98
cJ+w8n4GMOBRg5T5JwQeuUexF8Er0n34/kneB7QqnHIqdWJ0HJOCbzIsqdN1eLXp375xrTL37phX
dt04aeB1Qa9aMPNE/1zhXkttaWD9tyhGGEGYbUtQ+1i7Dl1zRlPBGEyz621osdf+Zm4gXiErQElU
lncdqj0ZdxH80wJBSgJRkObVWa1c0cXri6bmMoUaasnRIAPckht96VEMpffrC5djzP1ujEBU3//6
q5RGh96oiz01IrDxJ6bgkwR0rUQD6LD5fvVNGgSwoeV9W+ePqMt0f3V7RgMsNUewzjRAapJO0rfP
k0UTwHh5GqtLBUquP87MCeCOwt4WeMOkj/mu8TIIq1kVUjwfryxehxiSohvCbq7p4mvRQsaEbpKL
nfdg0RfoSMC0ZQmCeOczmhC9PFbmLudnpBPxqyfjwg7V9ZUPiihW7OiGzvIrCJGP/zqi3phT/mMf
jvPJeng1PEomzF/RPrHtCSSzww7MzDEEXdF1pikDIUx7srbfcoi8XMyjt/tMAkHU0oVuChrxs48Q
/vYjOnIxUZN6At/MmGbJJvWAjCfGYLSLhE0/E8r8/B4tn9dXMYgXKhw2lBlBYVqHxjRsEcvcAkQP
EGiSuah58Hkl9dIVE59KXsooi5KWd51bEj9wmOoLiqW6w0U8Qu9p47AVmcp4EitzFhzH9P/eWjq8
H28UPFIQh+UGMv58wZUfpaXeZ1rmyBS6hD246yX0+8Zc6m8187o+fXvT+j5GGcUgOAn0z/aL50ry
lwb+1q9u9fO5C56hugGgzFwuiGtW38VQFsdFg6VtcD02qMyj5sg1ap6w8NrWHgbiiCE/L9XEsNvA
RlVQqYPKCGinzZW3iyBxyQ/3DR+2+4bw7PTEXP4uyIW/553o655usfSF4RWv2Zhl50d+6Y86DAba
KGaQjmck3hNNUV3ONoYzvCWmcxjEhAPPQD27DWALd4GWkItkTUG024j0dX07Mjyf/DL2i1tI0YRu
zHyosc7P8ockHvZEPV+4my+VOdIJv98K2AXxr3L67SIPe4AtHVsh3C514YLQ55HfmWRdqO1rBjqT
XNBd7pYbmkqBms9OVPTM1uHzzWOrihcaeRHE9uB+4+aUtI6SdusZFBAlaGkfNe9sfDEUKpouzFlD
773efCVan3LWCBBorqmeFUyAUfBgrmALhIsrMDDel8qEohjh2WwtNIQCYyfrjUQHfRhrxlCbi9PT
611rxja3Z3wM3Dw5PF8kXlOCPwKBxoLgGOCgjhHIkCuBRd5ZUXmwrk+1RRoVy9Mt5KiBSLoYoy0H
jALnOVo8bpRYzImQRUMJF2OMdg3aXx7i2lLUifnvTzhOk6rNMgzC1bmOfkkrI5pQI6adK0mQxFgR
qoo6FIvLVpURmpC2RRxKvB4HcTs3ycgqe6EqIAFoOPBAhAoqI2m78eeZvBkS1ZabgvqLZ+1yUtGm
lmtbS2JvvZi4UbiFNDN/br4TuMSK3ATqg4XPinEh3hpe5ilza4qdPWdYGoeTcBkQqr6rsU6uClCq
tF5Lxz/5gwz3ljsccPvEdA8SRwTS2NfoqtfQvPE7NU5x4YiCsneB6/OZ8uAa7bEvnpLm/ppH8/03
tSY1mvGF0d5B5W0HrtKbXir1NJTvl1qcUnUSpAzxW55b+cvA6hmK/2OD+JOtjHO5tlwbmU78ixhZ
VDJf++O3Ew3HPpzJAcNYCOUp/Raf3CB1WQ/zjaNKhdaRZMOAcUjtKFJdaVN/u2+YtgvEcgpsWLj+
v+RPQ1L4e2SFlyqVNbUIKrzGF+PlYyxLkoQDHllmHifU+wYUvVHUx/vgvupCsI/s3f9njwlyoxdr
Vllev9qjAWezF03iCqBcfWLkh8yDf5QgGWgwrf0K2Q5/PPm2bpZQlueg32hqrZd5QYF+KpJXBsrg
D+cTKmhzlQFyYBXB4Gq53VLnMx+8ROTY8mphQaUCOgusGvDZy1hMwCTJgtNCBGgmQQ+J/RQ2m3hF
T//8fEYDzwJKHFNEIWqQTtI+ScJNIE1iGZTSthzFdhhr7Aw39QiccXSxPiNkMiSoUGuD6Ff6hTkZ
yFMSEB4jh0mMg9Xtx8Hq8KO8NZMq7y5YbE8lw5k+RUQOMlDaqzSRceC6NblyTg/oO7qKq6saiuWr
TCBGp718Xy7Ez2IKjheVnIX2BZulOIuShNpVJ5VmclEmhK2U+kjxwfFYIpeMB5C12DFSyVILOM/b
rUNIfxZnT+D2DaecO7dxlOZMvJbeC6KeUWw/HA71n96EkXxx4g8L+zUrK0tHAM9wW9s59XCdiTQy
vYOidvlf+GnNOpualAHV/nMHqBGAeWIF5NRRE/DnrZDZLMR5LhdHYaaLuR//q1Th2tk+3EI9LiZW
iLNxxlLGtLqpvqd2vquIpBOcBQDcXig8x2v44EGAHLMVq4yLYYfHSlmk6gpdQMLK3hMRxIOiJBk6
7r7mjOVdIM6lz1BlJGN6JrkII62NPuA/In8hmd8TZnpcM8mQft5AiWQEL3on5mmyFHKvM8OF8hQ2
d7pb0fuzP74y4MUf2fytAb1vOmVg8mu93EoHPkTm8+OTCP7Poi4g4Lnx1UK2VN1GEIhxT6nmK6pO
zPioMjlsUUBTc/WlUcQKiU3w3kEYZ7QK8OVuGN4P/UCSJKROdknGyd6aCxgy1pF6A0CF6mpuLRKk
NQazLENBnXfW6ToBzArxPsVFQTKL8bTGZZxNCw4+NEjA34lBk39zaT8CKes9+Jf1Qpq1G0OiCHJK
URMOntLXo3OTu7MAA5zfcvabt36giTQ7VryV2Mo08GoxQh1O0F01zIIlUnOsrQBse0cfEZfJDazy
4Ikd7FnFfhr/vZtchW6+KRrsEjGlmVGtazCJp2sbeZbDI/u//qys8EdPWTJGw1H6F0z21fvOu/7L
ujVlBho59RVoAXty1U+kXlqgPt4scfgJEoYGPE4wnzC7PM7AaW4mZa8s1WK/r+Ok3qi5mgBCkIuI
567i311XYCI38rQrlOZdRZBzUbYXAH18zo9gLnfR4bZdT+oItuyVzERED92dsUJ8TiK5BTVqY+LG
eUhrAREvApMt3IBeopsldEKxNTrCk3JiJbeNxvTQfeIAmkuvRlnOn2p817fYqgIm7pk6DromdJkd
m2DeQ2m4rE/yHNsMHa4ljbPEyhK70/kYaHhJViH4MxT74jilyHCKaibVGaG0T/MhIZC+4t9lfVqN
rS+UblwU07M9m+FID3AEtqUpFNriphVyIxGFhFQbNXD4tf5MX91No790j50O3GpAjjG5QUL6q+Nc
1lAEhSitsrZWTuWFox/vkZTv9V0qL1blVIJ4T5xNoagNDUBtbT2RcKiMitb7j0PVAT4wcY4PTw3c
AyUlpGJthhLd4YIy8siN/CHp3rLeKvY5ETcqA9c9YJxGtJRjU02SM2wDM3RJTVWY9quN2sjIhFN1
xvNPYTkx/2Kge1DYOY0Bf9cSp1IymM2+fu1yEa/fdcg6JMzcIHAY1nv5Dolp/GC069S10evGy97D
0+kYPNBi3cZwEG+QBNfdKoiR5/uuFJd9pJJdLFb3xgKozBcCXF9tYhPZwZX6zyqgzqrbaQcjRqJd
G+2U5APeK+A82Xa7D0DZQwgbCJ1p3ylb5Y8ij2re6Wpc8sjeC66eZiRH5HkgmO0Wheb67j9kfNW6
pj8l0wyW7lzIduvIb7BEBMAZL46YvNVP2Qerp0KXv1sBqfs9DiQPt4bFn1TIpcPq7FZI3KxKGVX8
fldseZQm9j4Yl9NqsorUxB0nxsqWvXdPApjLLccfoYCZCwAJC0UMj62hlDENshfwkCkakhL5ZB+B
XXg//owlOvg3P0sX8nVIpKJmopsjfZ+pePln3mNLNtIL0K1wULazuADkaG/TON3lIEdqAQGNfsTr
D2EcP1SAj/RCf8d2/YLmrQc8gM3/OV/sfXxG9uvLvLPfZHQQ2WM+SvqK5VnI8PsWwDJdGaKb/11U
HDRYOTifUqa3L1368AUfGfyYWQhA7WNen46UzRMzE+GCI0Jvx4M7tlV6Eg6wqpQJumfuVHKb395T
xwQmq5EjjQXo78AF+Zb3tsAezDBLC8A0i7cdcHvFHYE3GfIxq8yOfG9fP6P+7bLIR995eyoB3mmy
n6P7jEYnw8+AQjspOgncDwEmmE5ONPp+15OLBYaL2N+1OA/rm9JhvXdlVotlpJVhCgLZkxzseEms
rM9MIO4mPkmpJ2E74WCvZvYele5xB2G+m91tpRA6zuG1vDdVnUxMSr6J49c003/awGpbA4eTYmh1
8ZUCOrjwM5mhdx6GE2CFg2FMvAwU0IyewTdwsZ/nbvmAIFSHGykatGIqq51KLLkE8liMNdcZBoGG
2JM/GQxAkT2mWuyPTOmAPFf5544TLnD1s2tQHdMxOOghqxIIcn00N1f/Vc8D7drl5VSNkEB5bdZG
DkhD4wKIGAjByau3O59H2OWI+j7PZb62JkhplW8PLcgkGW3pP7NS0PKWJUYvorwI8zYVNrojEMGv
qEj6hLrEC6vy18gXPTCTEbZiBoX0YJROuYLA7L2iTiOnheqFt2zpGkJKQ8JYx+88EnDGfBDkPQG6
JUvVcxDY4w/W2yjekEquUioxM+BIbHKfh2WmcUyhuFzzvn0hXv/NygV3L73RsLzfS7JZGF61D7Ui
txPrHLUhSiOMa/Ur/ynM8CHYmRBCzZm0UEV/eosBnbB5p15WmKsYPE+n8smd1mNUtzWxBHe3UYBv
Lj2Drz0kPln+M4BYEvAr6y7PyYkKx1jcMDTN6m1AGHoJfMRa82XwAG2Z3NNQPs5lzCTFEsy+hDBS
8Lcbdm6+1whHy0q/NkzmHnCQgTY4szGkqHZcfVamTsYF3EloQrth7Hz/vHFHA1Tg6UlXvTHmcl56
QU7bsykbWkRl9MgVCcn1hjVrsQqFGhVhIHHic4FNHYZiZcPRJFPDJlhsztDlF86Mg8x/Q8/xuJaZ
Xe3ix0SfEQlybbjLnbZm3s5Qv0mVGPysfdWRXQMWragOX18vrsJNqFY6bwe7kK2c891OAQEZfdSB
P53Y2MrjPv47YM9QV9DgPfnAuDQipt1hQ6TuxukKcMKHEFi596HKoPEjqiiWdlLHl0qfHL43spBi
Es85kRwbyb5psCWeqcQ3EZ4YWAIskxHAw9+8zmuWy2WKIuya6EGhRED6tt3iACf56ZvRl8ZZkLi8
F1PD0cEdM0eBdD/2gAzPcI7UHME2yIQYIYsnJ47XOwE5TvtvGuUjDvXhqefc0U7ypfx4XXpN4KU9
PzFZZlT/vT+TODIGUAowQOH0448ygHyYljr46pOrApwg74tEJIlMiukKNdcDybHQ+XksXjMH0EBM
vwsCnH1OMm+ZJHUlzZWx52HGJXm82SDCbd93Z5ajUdV3G3w9fV4cRQdP7ozs+Wmq0qQ9MciBWSED
7dQ1LVsR/dUvRI2y/3UprUgIzKblat4qrlpUdOE1/mSytKVuqITG1K0Vh5VkBQGxzKS+H5c/OHwn
pzCvIl9bgBHnm9aJPZ9rRWVMV2HAkRXHaLIXpSsgd0gj5AYmpP1d+QMnijURkh0g8nTmKn414Cne
+t/bCQFltuZMVVZKWnIMYK11JXBqsgfB5Sou226xyuN8b6liNbU0jX65Q2g+JOT7q2Kyg0dm5DzC
xMz3lKnYXvUPH4HaQHuXPlh0sq+gtSpk0Gc46YN1gcfRBA+Wc+5jYhApukdN3WIq3tFvR1d52kQi
MnnaNOTbs+1xnxp8Ck8lTdGpD6+GlitPDnjISWQz5x4yOm0P6stYtXouUnOpqDUGH0O2ML6hr3ew
poei++MHN4PCWceZ13LRgw2dH295/KdPKSSqsQ0pex5Db+LNd0/RDwGK4PdNW1j+GHVpSOhfgamp
GD9ftFbf550n4SnKi+uIxS8Ga9467hzKPqujUCp/C7A8Na4gWaGb09RP9dWeO15ZnYCQonKzg1cL
01RQ2Jl0MtnRHsgHvN+awCZmqOTyr7zyhgfkkl1ljHbJf2D882AFsMw4Uw2cd8KV0fyC3N879dPW
yXBKej5DjUo0IIF97s7cxfXHh6EINh/1HRtIKibbAAmnvZrdQZtMxSHvur1HNln5twcZ56LFbp/2
CbXjMNS4QACGLtrxaIlklVpADrJLryRrzik5ZZNewNgADpNPJ/X9sz6/t352xTTv4v5fRw7nSn3q
AFItmeEm5BLPta39tG1bnSAMlCQjJLo6PPEO7XnfEpfrrba8iOo0D3mM5iNm6oNI5S53/oVb7C8U
0pVm4ye8ZMg3WS5fcKOVJjBcdigLfJARuWD82LP9IOIKLaEJKmGVXJT56W2zWRaHT0wIDlypSbx8
d5h9P3HkvRLH53ApG/CPzr5eKpdK0TT9sHFpZgRKSh8ZIekGXrWF5Zk3WWDMn03Dpy1h5Xz8Q35v
djqSvkxtpPO5wDnJoUR4900EuK4jzw6Q5TerRG6Tlwb3vKI8J+brJNYGhYhnro3+aK4Vc/ZGeHVe
26VTU3NyHKdzRVib2e96Nzob3OZGDWsO0iJniyY3CN+JeW5797pXMR6rNChTVxx6gb6UUUXlq2mw
mdJHE4Yx9W3qrbGGgtCSYJmy7SRGny3SSYaaxvpTBMad0A8vLVX0oD4f4q4cy/fD4TCHw4WLM3WE
j+sW34S119809w/zf3S3+UzmlIgQo0tlgck7VbTGnaAiOR4Zc0CylXlEEHN9VIpZhnKXrqg+5C5Y
oIsFs4j4hVnXiDKNmojBlEvt/Zj/buFXMtywfBKdVTfO9s+FsA0jmpWg1CmVLY5WCptxaXrvIaoY
yaxkuoUMLrM0tM/+pErHaF+JhNHOp8WiSuySu2SzEX2S6rauV87VygWOWLwmjVyuKl5JIKa1qHRg
eXF0zexcZr3SvCoWl32/JmWMOBdMkSpyjqMiThxdSKENz5bAsbmD/OwkFmEz3aluV1NoeUISNv7L
0/dToSbSCW64xkjy5ffeKnl0N3Qgwb+HaO+BrWOxJ4ITKmV+NeKv6SNuzYn6SiH3THPu3bNzXzOQ
vzQpnzhx9DOzDN0ln4J0QkwP1eFk7hWDkjo6Ms13VYhPdn49pgArduJrVbtUcUDyiWs+09dI8D4K
IccuD0rCYcUE7up1tMyxONrd9YiawaIVc8S+9ejcMllJaSoOhHxjO7mrkpxHSqfqT5HzOlYrCVww
7/C+JT9f+xNe6K6zUp5XdVQ9QYpMBWyURwCGEhS15Dq7OkrkuWs/mLcAgEu+mHZ8+QWeZ94W1ZOY
Xg6g5xKvcJW/jBCbhRLnwA8HdYwd8nMhVWxkDTSK/xVvkqzrjR2XycEZbAjuiFHHbOVja4VbD/7e
YgERg36x/cF/46sqzZ3APM74zASq4CkPytPanHv9GPx3vOE+MY/yvl15dZNkS5Nwe+MUtJoWfcy9
j2zYSvNP9OvTONmCccU6rUV8YpubyceTUCeGPmkmxjNVMRnpZZABGY+8pIwwr/XD2lNimE/G8IG1
Xmuh3H+fzzvF3Nq9Ovu2o9QZZufH3vqVLs8KBVVayr1HDf9Y1xAufbV3O2o2hGeK80Uu/erUTVuU
zd418kGhlFLhY4kyEvgJM5g4tSspfdHRJ5BNxJkim029kKa3ZuxA0SByfN0fRiOmxroIndtHs3TE
WvL45azwVNUsWmuLXk9J9wq74K2fxUdaVHkq02OhgAl0YHmQQtUN2oXbgNiPHIq1VVWvlBioTVWI
KZ4wamsRTKRwyrdH4HxgnU663QiTSiHKzIz3uOzXq8qVDIAvwmlWSKL4jsEPrEWHl3lSsk8eAuXn
erVCx4oD7mF7q1JMcHOPiEPi8APGjWJ3jCaRhKwROdxJBBLyUarcINrWqlFOqFHAtgZDNxI9jVsS
k85RlGVPczZaipJeRs1UkUolrc2PtvsGFxJgVK44c+LBU0HFkb7n2nFy/dfFFbuI6g93MIHEO6e7
zKL4nppPGgH8+lP7puPu516qglhcyDppqlRHjUP24WobWeZfjlEmNww01q4z4ce0MOb8XhJpx5fS
Y5LZ5YKTt+Wvkwnq9crQX7BjPyKStCuKqMzYX5miJdLnb/rrSSb1p6qUFRGhHMT1R0gPnIB6v43S
OkkDg1ouFgbz7gCiWGYRAWDEcFKpD6sPSh++Jbv8QpDqRF9y200KfoYQ8wiwhhEENBdP9JtGOVaf
3UlB5+LrD3y32XHk8ojUDI0g2kfmKE5GDQRRt3Mop28fAusr2UwBtqXd29bI0+gzO/ZHclS4QPjl
f2J3Tom3UD1GETjjJxSw37mljI3ODoSbiTB72Mim9aiObVheeGXcSqHPyrWuNHajD9S0CkeDe5DV
ai1FCY7jFolNQ61Tf0XuAiN+oQYkNWv8wmpPzXf/XuMh0Hh9msCIzFSLtS/291UPgPptICkR+35V
HeOvu+/Im/pxDfB4FJdk5zJgNPQD6y+tG8TFoLPxYc5WonhvgVEv/6004sCvbC+ccNtltOLFl+C1
h4/seOqiA0xPCb10YnFzC46a6vNbTojr5gFIWpZp8GlpwB0iBHZDUSPbb1LgJV24O56nZu5iG3JV
U/WQGrZLo3zmyn2c+ZvX8yWGaMan44f5zQqmHhNTp7fFCtXczdBJ6dEkZRx6wDRCibLkEt6/a9eH
/aCKlZmNM7e0tPjyEHBJSMIGqu8cyZKzPHwrG/LyZcljDCRZ1ewJLtzjhY4OV/znCIgIprVyC7rJ
UtafCxcZg9swcrSjEb592FRdmduiY9a6Zh8V2Q8dFHMD+TeblhxG2JU0p0ReXPxJJd2FtVXcK58h
pftOd8HlFmlXnc7fN+0PaAb9kI6+6Z3kaS9V56iQ2kFw5RCOURGVgBbalSeAcSRk7bymsPTEd7EW
YjIJuBMyiizMedahTTVYDxjJv3gH7oZ9XWraqPiq/Bm8ooaIsKbqG3bjqGtKxHEAU5Xz7pTZavL3
fEZLiYjSDn+7WB//Cjc9bRlhvKJGtUz3SfZz3OQxBMG7H+Ob7dIuVeDPMMx+Es4U0n7YIICcwX5u
tVFCoiT3tblrKBVroNMZRCwE5a9CLmQ1uFHQWiYu+Xy0V7c6v+FmWNHjOl+WQxfEeElnC6k+44er
QdW+Dx1bruvinQYZ2lR3baBCGjhsaWJqvYeUIXmhnt9hCcjiKec8ApqZKDHF/9jbsZWxVoUPB/dS
jkeHxfko1N9KJ6vauOpvmo8rlWt2EO8uZO/UHMltd5q1QPLDLeoNSHXA70W8a5jrZ9LAL9t2nTpU
v2EOdM7gEI4wVxKG1lHs6RDsbK/XkKKdu5ugSz/KP9qecaPoK8JTg9q3UyMVKEh09pPiEKHDjiB/
d7VoV0RF67APUFbgoldmKADhTehNzC2r6mEIhkVDO697b9tuRxgnyiPLmwCr/WnSwBGtErk17/ni
gXUWFc+7QTwDNdx9OK0JQopHKl1dccqeA36qbDzvDJLQqF0VOPgBmKY2RrtHqeosVHSiW+rzvn3G
UWW6qYCv7l1vRbZmw8FpTK2CkXeAm2t9MIYQhu7TtW/DPfPxvsZsop66rj2mTOZXgxJ9iKMKE8Iy
qoPUbpSHST/CX5LRlyMFbIliW2kGZ9hygGcNZCsZFaZd121ByCoAKNBXb4D1M0Es+gk2pcgI/x/i
yfPucTONHxOD8/vz6Swqy4RyzFqVXseSX3SMauePkR5Dsfzm8jTC2MwwBhwNKHK3KGvpwjQV0mgm
bZP99l/WMVSygQUWNOsbaCk4bBceQIAqBisE76/iOlkuWfZCbtukCoGB1KtEas0ONeXd9Nk2bvlr
f5kvgmE4HK/8TGWYvDNlupXoNUTlgW9cTdbaohlnepZzVgwgdiSS0D2Wq6THg1VfBtjZG9lOKdQp
nWf02fmg58ZnEy2A7wWqPt3o6zWjja5E0L2W3nbjXZ0/qZOxWjt/ULXX8NTYhdFz0WdT5XwHLjy8
KX5/WLlOaeZe0f68iLB2TThfBj2IBBRTT9lvwDAqHG6Bj6E+KavsYkgwCo8Qp0v3Lj4RoL10CkqT
2wGTNtHtWmm8Y1012yvCe4n1tTQuVMj0kRUh4ieGcj39kCyO4XjUwNia+iLFW1Pc2GyGPQdLva6I
jqrFoQJC/dkxX0CBAFbbG0E+iiLXgMfHedjyIRs6YFQYlPDouSGZ/A7lV+8eZCLOmD0uCK4cIVT0
zttTu37Xz1QDSVKt1p1MAYJL4L0YmZmgi1DO5JNeTBvtiF2mC7E49OGFOJwYqyUyuN1wdPM8A+i4
mGK3AjgqoAl9GyToUGh75mV/Jtg9vk4bAvW67Q5WIsRIfpg/qhUeEk9SUPwS4AAIT8R4Mur1pEqv
ELPH6ZnhClhbSNW8bslZW8sq4P3UfH8woinay8B19auNZJaLWinksC0J7biQ2TiZhqjufEZ7o9pZ
T2PayHvTXXZrxVImIVgjbHX/hLU7ciEemK6sPP7vfw+a7MnGiYKUQU8sti3eR5vOUzOzZ7trqeBH
T1F8Q8coSjehzITej2PoOI1FS1CSAFdPL+wn8hrrfu14WJAOwzJqhLzDoodKi2DvynsCHi4iinF3
55zJXWOvHSCQm5xPt+fkSUW3DC1uGuLIHdWwTS3dykealijaUGQG4OcsOMArLNW6U5JzM28aj6hZ
Jo75OLZi1Ailz/OuhNh4gG5Y5Bx9CGhU+VTBZ46SsFADbvW0fO4/AdmRf5WofJF13cZhYQHrGuBf
p2+kYMXAxc/Tw5PNMpOjkWmCqPA6pPGfqWItB4sxSirDcFX/swype4Kzve3b6wYsB1EoH/kd2Lue
MkYSRiPZfVygYrRlMhGJF/c1dc1YdqRITcvRZ3aFH6q929XPJdswxy4uR3p/hA88PA3bWEFn7Me3
ZI/4w4r3PQhQSUn4bLD5RXK0G+S/Q4St+BPOrNIBJe9qF29UZbtLDw+G6ygSax+HZn1O3vDD2M9U
y7vRkgVyvRsKOJdrXqfGmQTZvHT4o8b8gnImGJ9wvGCkFFL9hJP/M/NaFl1T/IpAm3Uu5cOjmQ24
lO/lJpyF0QRk/B/qvfkcot4lsuAiU57XPXNFsF9yOeJgWv7Gob8aeXE9tDdcR787ARghUYdir+ed
7scGQ6isIEZOOKvIpPqp9hPkOwHhjd28ZtYaXPxsAkS0h+8WjCszHcVcRCsf4Y7NdsJa4WiWdh7R
0ESSVZ88MQ3nShPRSZMWSnGofFA/H2atlPHAqTvhXjLi6wQK6aSUVM9XQZKfX+R7bWXOz2LVUVmL
TaZspHl3fqw+ecT/QHDEeZFqmiPwEn8s9086icmZ5MHb+norwzgEcdMzF+jvrhz2pERx+WgZZrFR
ThIpa1RjVCFUy7yKHwzjDd79mE+X0HLoAw5mfyryGFfr/oapvhbtPfnZ690TLw6/JXOL//6hZOSD
FswX1b1ivzRpcu4SjVmOa6NNhmcbPAuDa2Jz/VBpZKRmPjotKqoOxIxvfEYZTmjJx8XiFR06LplS
VsyRhj/GA9Bm2gMoahQ1YPiEvyQPq/I1bJoOZ2FL+kNkPz0zFTfZ7TgBbCpdkD4DVJ/qVjSkmmq5
MU7s9ca6nycYllQFQCmcN6AxxkAWtlZ+W3kR9sSsYs8iipJvcY6TEhC1yBKWqVabtleVsP2/szgI
9B7VSeMg0x8bWf6QQdi/BLTZ/UMOLCjfr8G9wfjyRcK7Jm3/QaCnglB8K/WjcAEOgDpQPVAgizkA
fc2jIwC6iF9om9fg/tnGhtkyY5mA5ajHoaPnMA4xxXYlGktYIXRwr4vApTqu3yfeEbOIZ7yuCGKr
QcuReFMb18AQOHFT/teDqUGJaOP5+8f/IlJHPPcJq7DHhNDn9y4V1DSj07QeTXkRNvsTLVEewx3w
9A0vFhVqO2dpEEFarZhF/tDnZjCB0pVBBnr7Y0OoxNKIoO7CB7r8mb+eLHJyrp8p3Lyxe1puhP4w
QL4CylQCxprqzma0BVP2KdkEXPUWH2EOhKOr+m+i5GuqJaJWrwJW+6LtAltm80iuHTYqGgRz6zZz
zIPw9wWcN/eCGEr/q2q0QjZ0JmB8KjiGDEKrBYIX4WzFLBv2K0cLkFwsMBNRTWpnrENvGNWPWy8V
I1lY4iwZC4RM7NxmEoe8hbtlvWa1g3YtxBzmFpQH7fZEREWFys2/N9x6nL6lej4VX7VQl2CGpLYX
tKjM19dfJDOARa33sOn16NQ5WY0O5d8Um0aPzpa82K2MnY4SvkRrWk4PncHCwW4Y1ZxAgt48Ld7M
zy9rA01i35Egj2I9ptsQxBFYQW4akDqLHxVLXxNOrGI6GezjBix/hWLJy69U4hS1J1ab80dJnxRM
/BlNfSjVBfnNLZYkTMjIh2hW9odp5j8Fd2ITy+Tb2hZQpdw3oI/JpQqOIdHgaYmibIJpflZzFVx4
qExUp9onsXxl989AcCY4htsbZIlmuD28U9tneCr4ST/WuGcNc2UIhTMTu4PyM6ElkjrzII4X/8Fi
LiHlRPUQZzRjq8c4U8+Ep6gK+bVnv6+ozv5erBBM1K3cQAf21Q8lvW7Vu83CsGvso4TDk3GYtPk/
gx7BW+yIkJW7ZHK3kckpgNy2ey+7Fv2H90aD/TNP0vQ7IqmMchwbxG4pKzphsx0MrOWleKElFheP
R7b6MHm0ye4Pcui2vkvJbr1CeczZ/wY3ecxCx3z+FmoSSwBNHH0RlQDISJPTJX2+3eQ1cj6t/l5o
zqjwj4+4WA2KXdk7bPXyPVLETrnCk9shkGmQiCuzHpc71+mHQs5jKtLaObwyzIvdeKnc1rjG4nFj
pEbWQdvcen6++eiSNNYm683zPo70Ipqc0Zmr5AoJq9XgNAHOhP2Kg2jbtkMaNTS1365otzvap3Ft
8PauOHhgULjoSNVbk7O01T97jecK7yYjK77caXXeEAY5Dn5z9pP/+iruE8gBK5qEXRN/vmlvuEbO
+CBRKd3owgFfM+fOFuTKq3aaps28AoAI0OjWgOgXUosUhyPLJ8wO8iVZ/vdT29TQCxXsLwCpJ6mx
3KdIu5L9Z68xrTBG9zyksfgoEmLM2L07cdIpXqs6DhT3RgOVEtAIe4U5QTOucPkif3Z2j7eH3DhS
iCFx88uCaGz+BHJrpR2veLmu1AQrTeLUcDBScZ46xR+XSkAda/3RkzSQKyJWznW3P+lJYg4q1h3l
XoKvlZzulS3G4lvqQ+tczq/MTQy6Oen4vsySCAhILHtA0+Ak1o/BwFytdTCJxG9IZYAHi4yAvi4a
O5sgGLmLntwyWDhtajpGjWqOQJudWf5gvcZTlpta34tFmKvzTxlEdOaUY7WdOoIh0PTZSwTWX7j/
8btFKvh0/bEEkhjmFbmbp2wIhTLZGuWR9smhq2lviyk1LExeypXZIMnMBVMa6Lor82+OWGrGY7ag
WnXDAGJZSqhvI7O4c9/8GY3+wCf0IfQNTrddgzBRz+IBOODt34SZlohcp5h6xHZ9ZWj3rWVfLP6k
rHUUNa3Q6038j0ZOV/tc+pXwMu8kjnaikbg2o+YpyXXfT4a7SP3m8lqUahfHtNGJ3gnxL92w9m/b
siUpDLukzT1odUauo88DjKghTS+vR7DxoiiEWBKDcpT86QfxPBhKGk4KeKOU/T069ZAmYmRCWfch
K1DcZ8qcqtmd6NHrhkR+xTY4tJZwWVRjAQrEFeViLEvFhqI+AbBsT6ZaGd3/u6n/3qWIxz4+ZmxO
4HWHsOIUuw6jGxVJEpqzEbd9tosh7imuQkVbGAJLZD0/H5WfQpNaSE2oZUiMgm164iRHXxjq96Gx
5OMCtPzfJQmvvxzCROfw/25WEnlAIr0nSydenEFoUBjqSrB325VPkpWFF18CvBV8RxztSrECCbM3
zMdRjP3l59aYgpnErQlQ8Y3oxuVdhHELEnE/sjF7WaEfcMrW8tLbg3S8a8kJ7veLUA87Hmk9EW4b
/RyZSGjqp8kW4P2Wyqq2yJgmcB5r/NRFgfIRT+0YhlHrgyP6fnCgsG1fToZVlPIBq7Hi4eCk8Np+
XnJPEmsXIszWFR1YWY9Cadht3UCcYRuf3tFokkGbpEmjssw2Qzt0VUMMvIWARYuXS2zTxXAo2qXn
a9ORwX/A3MtAxGFiIG7Y2nNomqJue8l/KDDypqakpmT5YY1wcApgXsCB168gpqJY1HGyifY9AP98
wNyDbLOsXmVnaOzgWnImAj+UKvtrWT2FeRVe9iJ55C6RX2eP6BqaUdvub7X8eoTsLNm/NxNVUzSD
R3kF7Tzu5LxZi0HASyHBc5cApxIRQPqHKNoUcUps4lYJ9xEy9LkZCKbE9HTKKWFOPjNp9C/nBz4K
HR9z3JrvX3HduYlvwZ8BUsc2koBuQ+NRrYpKcuvG2Xr+KiIbYqhqbDpYdBTOi76DAWdrASg1wTIT
2agz1+oDiK6SdzcjRYuUtSX03k72yCYrS0GTEVzmKbyuT8jYvYgzqpN6mVWuksqFIZNEjsG7NTvK
JDdQlis7k2djCa3JozYiixvUnbM9tpfKrAJT5TJG2za9e60nIEEPTSeQ8BMisoOKU29MsucFHr1H
c/5+1D5sUxB0MDpLGaZFDbUzm1iVnCDqsRWcTX92/hJK+hj2YImrZPzi8v8LpU2Ud+2eu72N6R7Q
9rb/7WOgLrbxuQQG5bXugGix3HvxIMYQKIwGRZ0x3oEAO5FUYt7oiX1saBKKtseEcmmde/VKiC6u
lht1sDcCOdyCTYSKPKyOf2qtcf/ngqzYZGLV4QMaTjfUc7qNzRSBsLcCMU5N1vrvlTWCI+X6MxUy
JVZL0oAycx9l8PoEitkA9DLfA1cPj6IPmDm+9wIQ64iEvPalKWLxqZzNoiQJzvPpfCCmFWPRnR7w
io1yjyWwio8idsX/Hb1/IrwllA7fyufWfULk35gx+N0OeCeoDHbFzpniVuWIHC3IZnKFbnvvtM57
KIMWODDL7JeZzglbP4sCiF41VDGwuWiR44P5p1NSn+23e8p9Kc3OVM2t47dpDvskp9Y+gBzpD5X+
0b2dxAxbkVuzXQqGGYKSeh1VJknjxuwJSMtRDS6CCrvCONyT3lVkQqGe/yEDBjTwwFP9yOSlha9p
qb1OxTlWqTDm0lvK6588UU75UT5KRChQU42G39iF2qTUiKUPZeVV9bRsSX0c89Sfta55Kea6H1FU
X2FmFlp8Y1ku79Ihc0WHE0kGNPdP5+TeKojS5jcHgw0K9F6Cxfo2UgMzBgte1AuE2BOxuG/L0RMG
NxhL6GKGT5O+TEd6F83Ekr3jtu06u6+/ttLdWaqwVFWPXdmRr6ONPbNFSv+I4LkjWrQtlIreK86u
LYw75/DeWHqWl5ZykorN3SMsFeulrddM2ouvN5CVNSRkkPTdMj2cOJc0Hyej/vI0V5blNDZNNCln
9bFIP3zdRy9XK/nV2+pqRPtUe1+PZg+erbEd3kAQWiBb/FoU1mtNJFQM6+4g0CnxOho/JaEF7N1y
HIUGb7Tj33hwMbD5MDLdBQ/Yku1aggY52dGzoy4CrzFoB4aTcBwkwD3S2hzR7RcoD2ZCDmDqa1ju
3IQvOICUIzb9a/Mqyz/T+bSy2TKR8Kijqp55G9LBTB+VPlcvfPTa2n7h/H2faek9qJh8Zy4k3/Eb
N6Dr+lMN5/HZJ2IZsuh18/iv6eiko+846IZm0LtJAaadquJCrMCCYWh/ID9hanvjChEYIlFf/9ri
yKy3d+NlpTlp5LZI07mNkWtc4GqPS0dgwbNuao6cWO/VZOkmYETrdRQCgwtPrLTXhDvr/H+nwf6m
i67F19i0IimwQ6fYTGDnGcupfZPov0twtYyKbUZTOQSURqy+qN6d0ibpqsFlnO+b8emeRC3k3Vk+
lrQelCuwYtxqAnG7y0Cgf0n6CgUV/bXdEH+yBWhPVfyR6TD+MhL3UhJEqxJJgQQy/Ez+SUoZbasL
+Eyl8hL/3m6fHXSH4dePUkSt2oLaUKELhOyYrhmTTG+5z1F+By8XqvoKlx6Hctli9OtqZpT0TFvm
8Qs9O6e7oyA5/twbgxD1ISi61otNCwfu/165zC0H9gt/Mk3/NpdVsiAL6hMIXtFvbhJZUMPYdI6J
uLNoq4NW96/8/nyNobNNAedDDb87VZeE6C7Q6ymwAHFnJB1Dqkqv9oJdeYPZsWNX6DVzl5lOuB9z
0IXIXZFS+JWuZdKCO4Pbi7egYAq/qbnRCt51Gd9C4xXaJm7YSaeBbLjaRFlX0vTHGo/T48hiOpIf
ticsBfo9MBaXyGguhbIWNZ13bcuNCK/ecTt1wccvnYvaAFowrJkaNVZd1NC/nTK3Uyb71g4vP5KG
alTOGv+B3o6jhE5zETbRJqxk2Ou31Gwv3qG5iXOX5JAP9PuGGA1j04P8ZOGHnsblhqG53kf6TT4n
xzTSUuVwP1fW5yMJqQOXqTc1s5c9fuZOqRam2yKjU6VpPSGFgDxN9wSg2qcSzr6P4TfwzjVvFqsc
edEHet+jKJE1knMN4LlY3f8gUG8MG1xOW0LWry+ISO0C2RfgYCLO2dsKu1yrxpgh5p7CPPvy6hBA
xzeKRu9nTcegac2/FG2HKqD/0Qz8jslLDzGli9kh2FcJTV8riU09ivlkdzRWFBOQRXMn0QfP4A90
Oo5yukHnUkqygbjoh3ncPfle6zOGKL2zfLmtT1WY/c4+PoegeQv1fB0HS+SGeTaRLuySeDln9cVY
Yqnu8Dx2eaUn2MuX4cadJMRzOYEwrqvsgtQIDxpb5GlhYqhh/JG5bu2iehAOtrbgSb6IcTN4JsU1
smQ2yhYfzoDhwSuxCTN6y1nQpXPzVAnEPQxFEFX2skGmFH5ay+tUvGMEYGDE8QQ6EkYLvILNcEL1
c1dWC8payBJlOserv/J4ahVQcRkpvcbQN2qbO6HI2kDxUejpchKTLeobfYKf03PDqPNLSqdc6Bmi
FKJASoLPJ5UOWnSWYJq0uxoOYA8B4FALLKIDu6TsVxD3BqHgKlW5HQjRfuWd28hCkqaF0BRQy8Xe
vYaGeINI/XgTnHigr8HjAvAEB9q1O0QcacijbwNNPcHK5E66bNO5YQj573Dx/XgAPs26KOAPUx8Z
w0xasUj1JZAJdqM5yQB5p/cpwT+TdMPWqZbAV3kb/5haxK7Iyoi+2ZsGlbZcCmwxQHb7MnYMfFn1
qVtWVWFcCwOcZOiQ858aDMyAs+bHVUcXVFBwMoAyltLG24OnogVFigQN162Afw+y0KRR204jxJZZ
ocf3c5BYCEHZ/9PECed3WD7Vaq61AJu/2bLjvNLnYY1eMmPRo7C6Zv8BxepfuwuT07fpIK0lB+qZ
SBbHAFBWSaNAUyRtNHo8jd1GsvqxjXF0Kvc1wRYxN5NXcQR3yNS29yo80ri5cNFZvh+VeJuod1vG
p7sPot/42rC0ISw07P07/tx+ZIq2MPmzWIt6X4bFnfZQOucZBimHsDnOwE8AFo77Iouby58Lw6l5
iUjbH6TKRhgGSrR2b4PiqIPNAx9YAk5vucjUD7aJS99ibrdJgnb9htrutwargLTEViEbDXaVYSip
tF8qi15rxONQkhnlF6nrk0SbzbbCDYfRt54P1asshPHdmFE49Dtm6gVNjz+aepEL9fG8mcDKVod0
UFMkyfxv/gTSpFEUQGfjs1/k+Ey7E6/LBuyqaImD9/YWU3gkPSHojTgnaMMr2/oEoahRkhqJLxaU
luw3xsgaWkml139FXV52OhtGi7fBQcs7xUr5W5bgR6t/3gJMdLhNX6pGXQxvHbjBckrjLNhSEbqi
cIPOSYCQ4vWHaC51ixLV6X6N3aWvcN/gpJ40c8A2eouMbSIs39v9WKu89nUVHI5vumPllkjnJ2PV
9yKOylEEMiAYO4z4CFgf3mp0ld4zuth2n6RNSisoNl70OUIez1tnDP3Gjugcg5qmCw2/ZJItUDgC
eld9iq64ITs6HGHJ02BGKL4CItyJO6EIUGP8L3wTeBPYv5H6M/K7LJrtY5ebUN29B/ki8WATWHo9
aJCB0/ldDecC+kP47H1FnbEXqMUN3EUwD88lUfjezQ3RuKn8fsANpzA/VmLhnkad74/oe3AwBJoD
RL2CKNa32cCqjovI5GIQ0R1KVPrCT21/vkBxK7ryU5FhJbdiZLa3cTtKKkRAYonF9uG8XbfiiIXX
Qi+T/G4KyruhuE4C6g2X6aAvudxp0fAk08PI1QSplJ3UGPGBZZDhYd5W5b9V0PVJ5OcEwuoH71aO
ELJWQqxz9YpwqFdwnRykMojYiFWnpwemEThwtOQ+FmiCSrJJ4lk9wl0Kb4CokcQYBDU35awJvcAV
kXjKu+ZEfwcS1xXhV7YU2p3kBwMqJqpYGomSW/Ag+8qhSLXPAaqDJyabtonM8TpAXb0WlUhkrigh
4eB050/t7DlaH+ZiQIRLQe399ZAy/uLc13M7bmhLOQ5S5wQE1hVgwIK6zW2es1nDA5PbFJgSS3YR
/JnjDuuBwUyck0fPqzXCVXXoa/kfgjf+WSJrFivLeV9MVo6gEAWQVscCJWeettUBf7Wp5cGAuW02
n/+W7BYznZIVss1NNh0m/wm2twWEbY5uesg753rYbGE9NWMIrZ5SAxyxFot3R8rXd1f15M2X7xOF
pApdQctk8fVoF7C4FcAybN8N8PyUjk+lZ2sOVTSmTQeAzWMEpq1g8pfuEb7c+mJKX6cwzmbyyJ4e
ADOfjNcrH0Sd0j1ZtcpDR0VTMy8Hyu7ZYBEUIalO5mdDdWMRNeYOTJYsb5HO2jxLsOWReRhmJcwL
Kjv5yxvje15TJjHqnopWnHXwIlb1hKPbU/Sz6OFQYisLiU1wAGfSXhqnK/DhnP1Awh0/IaElQt0G
kxS6TzDtJoO6yHHG1RdXN8jBR42Uykb6PSc8Rd5lWqNt+9gn886RZYjP0uCsbrYE+BRdRkoHZHA0
vA6GUEXsFI9NM9lcezjYSBtAPWhE4K6WFKOaAMagxf0ZgbAAE+WqTJC2THITacRw791b6jGApg3c
nkoXl4bDCr2DVS02wYUSz5uHxJu21NYvxxbxC4WrnjCbbHc/MTD41hdA+oX8vzb1bmjdhNHrUvel
pxhxnORDz7lXlGtOEFw7B8GgVRaMBtSCnoMsrI+dMvtTpBTGjldEPbdwN0jvMbBU3fFYBTsgfFX2
It8U99JS3H/3iE9ptJ3OBGqrcUUQkBEjqcrXRtAAiAoIqPpGgjWcmaXyPCemk32L+PWXSE8sgqQF
x0Pr1v8RlSae80MTDlRwKFy4G6RJOBB8hfBXp0a7ZI/Z/jIdfTKIe0MINRu7yVmWyYvWV/noT/09
WFEce3Aw+uXIzYHLM7dEXpaW4CBkGZP/kZGcB3+ZmyV360h9ZbumoSiKsyIyXn6GdrWQvho3MMoi
wzY4LYnLcGOJfnpCSiuCYDwK9tKwYDXipB5RXX/3KrdQvahlFLPJL/zjTQUD0UF6QV1OQOhsO06Q
QJXdFfZCITTI2RitaZjO6YJqmhKqbZQvx7mjWmsw41Qamh5DvoQN18F/4Bf2toPI7Uti2/ahnwAR
+Eg+g75Y0FDSd/ZM43968+YUbRg/xD4VutmO5Q/oFDTJAk8vVlvlxsRj14Rn2QY4CAtWhpRhs62D
fybDq5xpfT2CdsOVzcUJPcP3wK787LMXWb5DrFi3oyDhSC+bRJGc0TfEkj5Y3kMS17sw/2sAAKTb
6bNOXNuOsN6tMQxXDrhahmNJKq4QSV2iM2TR5bnhUOtLOJl8MlrHGfsx6qqAMuAzGKbFdv5h9pyP
isVXTsU6ebO9BGaBPv9jWjMUnTe3PmTc7CREbp4c5wMGR7xNLfQMtNXqwWRsO+Ak19S4Y5bixc7q
ez28QeODk2zip/eesAbTdJ4wp2gS8dIfo9hAdh8psgcIeatAwGlLT9fm7b2D7eK38fqOhoOE6CnQ
z7oZLCE4xyiZoRnP/GX4F9xnQD6mcDpH+O+Twe9Z4jcxkdFiBYq2lDdDL0x1CYhL5/jbMxUxykUJ
mZl8Cb6kLkSIU3cHojxqEre2UwAPl5jDlAZQ1JT9aE8d7mWqeBwCXEp7ro3t7gRBVoJNKXs554PF
GwzpYh1oVBS7Q59XGZIZ3/THrmgVxw+ABKCjdHeVlFtayzKKyjbxZGXl3i53FD70sHH8elYZrcxV
Halc3CGJri+whhloJxTgzFz/kZbS2KwamhN27qTQ+xYDXiPVkx8doCWRNRXohPm9P1aQoEaLDWDT
uTBAxQzWy41mUlllBqXn/3Ylua/7H544JM+K5klR8Ok4j4+CCoPrPNOam8cYqgmndMUD4kXsbtZ7
HzgUCp41isFGkEdkYJ7XgoPYr0HGfcNcfgR71mJBsbVGaZAXl8YtaVRgW7NKV2w8KDGqq/omsuPG
Et+n4Mt0Eqkk2I7utiew2qr8j0N0KFYDipj1UJ0OoULwOVGJa+L3zsj2S/VBWunzFQaPc+/eVgyD
Nvr7+0cWe4XXgNMXdJsl4po187An8FQIv5GWluZQ5ArRyke01iPH4T07V2jc+EEXv5Cvs5iPZVvB
PBsXv+fZ94sAsNB2CyubxvViGOrFIsFDF8LHHm7ClkrQD70Ldn3efgRkucDdTMlGmexIogh7yPme
uASc87Kdl6BGHDigFBjHZfI6BLJz/ySepXzXXqM/1nRf8NcsuoJ0MHCrw5s1TpjYS2eS5f3oNN/N
jKrEYAqNwsuLsoAsiSYX6TA+mv6cti9EJS/FdLEL93cVev1pHLhfnN/5dmR2Osi8CIZLRC/DPN4v
AccgXoanuYptwp+fPxH4iy1agJFjlMWTVCZjvzXDUS0vpUzZbBSykeq5OG8+P32bggx23o1uV8+N
JMMO9jJNYMuiQ+Fc1e8TV/Pp6ai6PN3WNqftv6o3Kp3UbmhQUyJ/bgTIhMXukyXGpvpN3anatw22
K5ob7814ysgl0Fw6+J1sp4RLQIc3UzTsqfkvf68RXEcRKD1fMit9/COuZVBxxRGNp8IadhOyrvsa
9FLfObMH9OHPYW13+l/Au1anfG+U2/jtlaDhl1wanmOaAoyGv3hZYbnF5E/o9bqIC5Jv3w+vJOgd
mjGlb5RA/9MW0434NwC9K/UsCBevGD2Ncpqtspt6PrKCuRUXvzZq5v2aB4T7jXjisnfwwabxan1g
RVIoKWfr64ugcdjr2wiGwaETibf7Q0FRUMKAvKP6DAAX3RhB1BePL7aNQkQqKjUeOe6NzWzDlxjF
s2Tk1LhC1mMupGuYJJrslRa7+oYn2AJjO/L1GTju8JDhxTUq4Qw8Rve0PRYdi0TSseERTGgi1bZJ
BTGVbrGLmOPWrUAh1PXvRn2wqrbrUAyIDq9zB2JPkgw6uFvMph2sJRIk3emHWVvLS+wbSyhdaND8
sACu16G7CN3tMlWLYQxvxJI/4O7rQFJhvlKjtbfSeKmSlS8Y39Q59IPLaH7kMrQIgHXFNVo+UKnP
FVWKyosnHnZZaGITYjKwKnZO+1w+DGC3IYLKA9GKK+oZlsMhGloL67WcAv0nSOJWBUMcK7bvKIr5
ReiiubQuzFFslxRMkElaUmvpN6jBhpu7an31MUS8SaM67PtfsLak73aF6Mfh74rb9NvH3wOaoNOp
+uRi97lUoypZxEG07tjoIg/OXZYR4muAaLQ6McTiPEYgqDUF2ETvY4wlwL0WeEkb/PlXib2D/Fub
BkZyOPI+svcs9UvdX9LrUM0jhnWoI/+sAi5P76lj0+ZRhsrQd7Js+zhokd5+PXZuu3DxQSyWt5dv
0dGoM2RRaw0JAF211DMvLcHJN07mT27JaiR8mMUwWPvrWyLOSLbZRTWgd8veBjv4nOJUZ+aV/CN/
ZdbGsavWU04u435/CSX0+whgTHLzVU664Spt6YX9xt3MHkJVI5jrkfli+sgJ8AM3xnMRCwYvXiOD
wUFalLQtSieCM/ic4cmKK4A73mrYbNvuYetYa5wbIUFckMedZ86MAlKLSh5lVDwXD3ZghPRqMYng
Hxnf1Wri5bW8ZnDcuPcX+MWpLrCHZKI01D7HHn8+RAEkF1I4/05/q8IIR/BMQ84g4MMmhqQTGO0w
p2kTqtcMpZbnilWJS1yofMChN2VqLGjaUggf3cntKz7Y2gshC2e5H/qN5PI0QiDs/bQsAJQ6ovbi
K/tDDKzhcXhiqzcTuMEPajmw7K0fJ/LvDnycJnrJz5CEYcKad2ND4F10me7nZJ3H2PlE2O4rj8P7
9WEJBlzAWZWn15HhOfHtw9sl8vVTkzhH2dvGFvmc1f0Oja7rW5+dvym6xFvlRqZqOE/9vH7DUrJA
nQZ1p5IaN/HMNhm7+itAKVS1KrqmaBhNrfxolsVCnLCL4ICmz77KeCKvnSQewbD2Wt5AoZADm1ch
PfKZSfh18crxYYWkOukQnw/EUH1SBmxUNHRTrSLAjQWljldR65bPwitNtkylnH8uTDuCNXPYY6u4
WqcNy5Xfe/FEtKnDbWuiJbSDHK1/OgOSQb3K0bQL30nwmUkxH8qnbz95BVzVGGAM3l2tD+MxRQ8M
BuKyQMz/jgDNBfxBqtWKazDHp5Hk4H3Sufi+gyaODFGsmQZuDffi3IonkmYIMn/WsrPJWuSlVWWC
SRWegCBXlnQCyEKB5yE8QWJ+mUZc+YAaWprzWcDzMNh0V5aF2UykZRXnYCRhoxhNklfHGIpcq+tH
aaxHZ85cXQPJeMXiP1VFAvIdg2eOoLyGwwRhJ/Q4mgyhvvo4++OvaFG6UrCky64KN3Y2NFDXr3kO
w30FIJkvGz7DBc7f4Xa5eiOFMjhrqh6A/J84A/aZIg6oals1jftu2qPEcz2zTGMoU7XkIeKCtLKL
wxbLK23Yzl/3SzpTmsq0DLR++d4b2e9j4e6JNN+OyLWR/4TeouCMfbaMFVHGbZZafRExpw/z3aWR
mxalHgD02Oa9vCsFo8+ShlKgpMzJCATM/jnffaEOJzc8RDxMcrkvO6GEn7RMpoGQ8poB1+rbTqsd
6VJolqZn8+OcsiYeZ/WFY2aRATwPL6PXyOxJovBo4U1jarzZWfxzCUGdhTFp/ptEKu8ZgzvkudDU
AL6MZ0JEUNRpwU57hIWnucwOdQWfnttY3Kbvew5Jc9BS8gBR84jI2lf2E7Y7F5EhgLEhOJ3PIGyx
WQA2xj3SkvAXw/wHPi+N/1Y+1fO/hptPSC2iuViTLmqSV8evQW2w4vewl20nZiDUZJzJyM04JOiP
eLwBr1sSDICbTxoJOYeRaGQZi23KvSwfALdXpxiKE4dJTmvz40ma/kxHYgjxSCf06+nbOgvIlEfT
2HBQ3qCKFyZyOPwGNumzRwwjbUZ0n9jOrvksbjIlEXBC5j5K3kwo++Jeda/XGsD3YragJX1etPeP
+KYk4ezBJBz6S1Jq2CuLcdj5aZwceWVF8zwkCZ8LY816TiNAOUVC77FOJ/56dW3EOGUqxw7Vl6Xp
f8oOvEQyCj4OMlLfpxk9Xie4STsYnsjDb6mf2Z7oOcO7oKiZzMVvwUzAz+MAWIJ7uV+YfKpZpifc
6BxheIjBvvEQzV4hINfDlvdQmeElwSJbXN5bClAeMhCGuJZb2AoaIzM6DFzQ0vFDO9vP2tRxCTgG
bo3cml1Uz7GXjmZaJ42BGssxHSTCDaXudTe/pFftJFcniLZ7qy34Aih8fXde2blqj32S4TCjAkvI
hgV31xWIj/nwsQ5M9UOsIv9Mu7ZTVz2fNr4i4jdKSE3EQ9R8pJ2bQCcaY0lgb7wpS9qLdPjbkfVa
jPBzCFJGSC4/dophRwlvOJpQ4+jSVwdeE035yF3+xm0ES0xJ6rIK3yzIRy2nQ2p7XjhVipC9QuiX
Baq8Algu3rmmw2xmCieQ+3Lbr5L182z+Cas1L/uTonF/zGPrTWn7q0+iLBOw6gnZ6GKAjqTHIeTa
WIxVBugc+rK25SS+LUPsaAG1GFapCXXUlkycaLH1tO1woxGKu9pJmtmhNcNMBcnUMHe+gUeeMevr
Tuj2mOPJh5qi4OqISr6Cxam338oG3ccwkDvqFnqh/l9p24E9L5vaJQHenYQYwfgmEWkymRHtAQaM
vGgvwTG0Aczu0l8RMzTQoX9ShUdFcYiPSw4Wdq+LLEnDgva1JyTEnoS83jR5MCp3YSHCKlbYuvRK
ZgKvqjlMt0y9TIVomgS8aSDEem09GZIYnWLmgA0URDte6jodAGtlYKqmK2BnWyg17LII5kFIHhnA
fBFx6qyKVToM1ta90v7sOnajOszR1IMl2AChV/L8DUtndH/BAg8THEo/HZs77B6wvgKHwPXcvk9S
AtKb0DF7PMsCdszIbefVUCpIe5jSbBR2nufs/qDH+JrVlrre9KafGfNg8D2QyoEW0hP4ZnfiMMsH
iN36taqysTR9RYOjJuadC5Uj6H5XxHa/HSllOxOUHjT+oZAWoGU8yR/NvxuCpkUhEDOenudrmwpb
NJ2oEI60oOPuPVgVci0VaFM4UZ3FojJDCg8g2gOePWMOBEbZ+ak9wwzlfnUpIlzb9i602jjP8RCd
3WE8LtLwIpPMbW4nJkC3IWs6hNTC9Pf9Jblfbf1WFFOG7huwdWY/sF32NNDtxcK+jlTZJXpTfx1/
hDJvLEIO8NZ6gwv4qaE1D2CPXeDYpZOIJzSJgcBz6ROUre7CfQz1i/gArdRRoyEXs9XZpXIqD8Zm
avgp9NndjJM62e6IddqELoGKytS0ePzwBtmjVQbWr3Hbv9od4I9UZf4T5QCBlJqrqcu+mozno7sb
CAxfq+HtXhgnPioi8+hl7UOOnSPsEQcUr4k+QJ+Y2BdKIRuzmeStZmnuKFu15qAkYTNl+hjWGXiM
1Q5wxH1mO6VGQ3pnbuW6UICEmaqMByTSeKlONsQzi0Qe0RJKrgvnajuk8+7jsjBZ7atxBUFSTVfE
PbF+pbNbnVrMXRlDK2TRl3WvEMnGGl6qf/g3U5Ei2WXz09BdsJ6i+h27wVUVR8SRXQKebM6vDE+W
RC4fUZ9eHMU38g2sJj3+GYA72SqzsdNLzbuRFMKftU04D7WPKDrtxjpM07Iizmp2G1XN5tBpB4JR
jJc6/GPLril47SvBpLmjiPLhhyHw8Y+lf93Dlg+l/H+tX59V6XU/MZ9MsAfMqVFSUjtgcUFGbwgA
gg615ucFlBtMi4E2NlxuaGjE0FZrE37ihKdESBQceUtf1El05yjB/SlHP3E/a0V4WYb5ukJfOPqV
jOeTbnaRdgFGVVKjNkJ6Lw2ghMG2TgePa8YUzOhB4lgwVnUoxlfkxnx7ql91/dzHyqzJ5LPtUbLQ
QTzDuIL2bdjVYe7LreFXeF2EPv7PSjR3iBwnMABINbmy/3/tNjDBTG+dmLxZx6fD7r13Me808R7g
rgqbPRxPY//AbsTFPIpe1q4FKUhtw77ncd+P85XI++lLpJX8jZuM8yO3mIosJJ+TYnSesVZde9xf
ziHFtUboZ0/FPwlUaoSgiU3t8V1CSFiGSucYfppjnUpQBAEqTugj2FSvYWsH2mzD/wbNUhaI/uK6
ApliKiftboS32lkkK0297mJTW+HtFY0tjRLjqO6CHlnpdnT7GZo4IWZ58ugz5auZz1SEORZieUD5
Al8Vu/Tyb3fZ6D3ADHD6mWjNR8DODmgqGzi4uv5ZSPaP0Lq+b7vncAiH1cK9g5qk0hI6eo4v4rRa
iglylLF66lBLl7iF1yBW/S7jiPV05HNgD2vw8xiKyj9bpMYs2EgYxRW2Mko8L9AJS4lAgNJq+kxY
AqE+ik75sIfFujcSlJgEnWJ3bgOFGK3aD7zLeOWCCEZ5zXtbA4pL+rcG6d+FEPtDkXUYsBr7ofjz
57s3e8QCbMLwwWWotVxUykRk8A/7yLDvTH1BNruWf8hs1FZz89PGRROWlbeL4nEnUKA1VDWOENom
YHrsRlxebr2vX9uSyoItvrtokx5moLWQ97zKY8s9EXeaGrRVQL+gJlN6+Mup+CBSF7mZ1+ZRpxmR
ZyrWrqn6M6yrQauNK0DtctUDEDRXXk2X7qfbf3lfD+KT7AFJvImFamnR2xBpPXcOakW28cEbiQQ8
EsKl7ClkHi4eDSTnNIB8bBSNFtiKb2dhcmJ9//LGUP4IlyPgdvzPsCQzO+V9TFCl6g1x9vrb7hMN
49/+FcPLl4I4dfh4vj2Owr+8D7rxiMyKGAwsXFYErlZF1+pRQswlSVSx27qwSB34msS84a0XKNJK
+JKwZFp9++jhIW/sxI7oSN0Umpr84qhgdVHv27rq6FFZ+vlvy5aLPDa2gdhfxOflmrVgnJtL+mGR
vByH9vFcLZetDUN13SDDFyCA4ogVvwBWWTcRkwK2GO29HUKIsmbupoJA9sf2GwcI0iBppaltL75m
tF5Ke3vtbWVFIgcjbQXEpLJkZBgJ2rHeckXjzQWvqiwus7KKDQcRp9qRQ7UpZ5W8JjU1UZhe1MSY
kVR/tLhm/e+hFzWKDgDtlOI93pubWqLTAHvZFpvteDewDcGOm7vrCwm7sIfznKBh4BFonoxp39vS
an5LjroUF1rnRPuMpgkuTJplGYOM1Il/7FnV0ydSrokhffapg4wICKjRdxcMl7yDmLFnSx57crf9
pA9hmP2j4OLu5k3FdSbXMfbfrr9v9iS1r8e9Ll97FqsaeMyzIvlBCTGMvM6SqZcNC/WIyr3wIfE2
O3vW8DQDZ1LitSqN33QPusDU9R7ur4Zq8iUFvCJQFIvMWVMjxlzglbdklPrzFYXgTFVcEIK+wu5i
h5gcRq91QEjcWXP5mvdlDl08NvxnIJCDGSr3WDkRrR+beUvXiglkm6SdpK1XL2psjlXxTT6kpLqw
l8S3Qo1cUTFwQQXS0TeNipsJQGYXJ3aLZfn7yKv1t06TJbD+XDIchu+FtgAdN9sDqeEcz+4tOLIC
fHBS7wKdDBulqsfRFZLm1iTfMhnl9ZQPxPDwSqy//QvTFAPmAa0CqpMXgx+de6ieRpudF9itmv8Q
VurICNmhAuRg36u2CZHBNjGs6783qqECy8yY2aijsC3MYbV4Fuh1FVvwff5HnI/Sr6Kdk4kIkSl0
vjqSTzvUCsuwUtidXrYtU0vDWX7EJcEl3jly8J8liq46sRz6JsJsqRSBwh9JgCkGjkCQ8kMXL83n
KGklaGQ0l1RsJXIrGkElamfl11dDpdxCgpBGKjOb1FO7oB8dfVPQZJUe5ZsvGSLCKvbLrFS2bl4e
mcQYaQXA42F9i+4GpKOc+iqDPbTFbEPKy5aG/jAyle1fE4/mVeNC5exN4N9epyuFjoaBII3irbnq
1Z4K6/wbsSVTssccPPYTm71KzLu5cA5M4yw1+MJDQ6F9pjaKhW9bBKnmBSstkXL2TebJKZ6YDKaM
28RzStQKh5slzXiuY4TC54sqPUehwOGknoIcZ4gCoZ2ODi8AFegfYX4OMlM/JlMy0PyEyClx5y2W
uEJjybenMpH7iMvQ/LhIEgSsdfZZFuHPT8e19tOKvfD13YCT0ahEsq6zWr0A94qc/cW/9NBQCFxa
tag3D0CnI4OezgJc18kvhk1qzS7o9wsca63jtQJz+jTODrXMuamJuSbTNOrjoRSsT5xv+U4kXS5C
QkGe4zHOc14LWNGGvNDBSuYdD5h5cvXeiA9CbU2kvB1psTw+OFUxDjlz3viKoR1nqaQd0la1/eAx
CQR652XlXtf0mBjZtaiBl6nUj7rhjMcxSfLa5aGC07g5YSnedgLB7b2xWWSJKJMws5VhCR6SoD8J
0OgWjLYccubR+Ux7X1HT/OedXJ0oAu0e80rFX1Qp2mJEGWR7Ztp1TZN5PHCrK1fxYRmx/v+kS0FW
G4hN+RNT18o27vDpOtO/pg/P0A74HW5gTLza3cY4N6h+izNHkfXQbuRpyO518eFkhRJUrQa3BJif
ve1GYWGt46jV3jy2oMxRybkQZQa6PGoPfHinZsWes6N7EOGpR5cf3ink8k8xS0WolGL1gRBHsQci
fyCyO1GN8c/50OPTlU9mUKbXBg9fPuRcnyNxSBTaBHQDncneDIV7G7+EtOrLUiPqRYRx6l37ohEY
U7/s5zAd53j+qYJriHY5mSq2hTwh/dC3NyWRv/lVUyM5C32MK90WdK/DgdlmKcZ9MgzHXJbsP3xA
5arLyaAKfCFdwtZtfMRTJoTg5RVy9h73lQ8qqbb5UQ+QpEzapsB+Njep17ITAPnpjJKipaEKPedY
25nkkKPDowGTI1K9wxC9TPF/HUsnS5wDnpP5w11Rot+Q5kWMrvQIjmCjraoQ2orcbIZFWS4R0Kuc
rXMN+GelOoUvj+/JiInHAUE4E50Io6sPNO9M2uWLm9qrpriCSLT9MOQVd6/aTX5bPIm538JPAlW3
h+4Cxn1o2c14+WnhEvUFqWtypLOg/FnIVD7C5MKqwZWUr+mNqdLOfcF/NEcYnKNrqO5IFZjF6eZM
Esnfl97r0nc7uFY3LiLYrOb8lMXiQYGlkIdHjZ+1zO4GQem1x0ESOMKPQL9w2KpdxrBprYftUJWv
oqX2Pn84yXyzLYSiXXOekO3qu08PF4VauwPqPNEjiTNjLbX9dtc3PttEMHKqaQF/+/GI5I1KjQjp
8yeg1GlCsMpy+MwCWQKxH27jo6z4DEpg22YFlaHWdtBMYjfBRbN8BkUFm89zlRgldxM6DGEG+LuT
QMtl6c//feFF586BgWiKNg5mkGojiJOsaLkl2wdTh7pqY/1xBh0rIjjR+KkM6xTNpLnS7Y7sRnXn
Bz3yWKp44IiKhkqdMzKp9XwcdInr0CJrjgc+U5SyHjfaCMXfj6yEQfLvjBjwW6jvE8j5+fjL5cFY
pW6/PeTBbMbBRzLj6myqFP9F11jSpcAJxXny/kW3/UQyeGLwnKGmdtdzz4slxVfhURqTLbIZR/cb
6gvU1xgSnaT58DTxBXHC0GGGKAD3EP6EWlQ8WTWX4uG3Jd9kSokOSm1MIZx8xVHEv6xPN+g79NDN
GpJABPjN3F8N8Ka4KEMKcS3n67npH9rkUVuYmLl1/v10Lv0Sn2htw5PEd1SGJk8uvI5R78SkfTRT
PNCrYRqeOdiz6hVPGmfK6hAowVhAOz9Wbvk/M7O3aD87145pASPt4VSsn0QGLoqS+V4Z+gRNFaZd
PFu5rWu4IUN+wk4+SLCCQhxRQYmjxSsk6jvGCB3Rp5CkADthHlM9107UJtsKU57v+9Xj9v3SJgXp
Y5Uy8q4qTpPyyPyNTqHb8axaMGoMRrcyiZyqOUsM79nKgtIIVQiuAr4HpfAYm4B3DFGdpo/WkmV7
RAiFYmomuZGnwWIq60HqEpPXLXRvjEi1zzsg16ow3uCR2c6H8b6LWhIAT0eN4ShHILUwlP3Imxzg
Cu5G8urSf1w1/lVhgLtBFQO9zrf4HbS/mLMnmNZQC8mOCfmV8qzWmUz28NJ/i3PU2h0oRbk76vAM
Ps5Ms6pO0yCpVMFsBh08AxlYjcFFWN5pDx/nqG2aoYwaRD8cQFJSJ6LM2sDpeQ0HgnHblWOUROd+
JON9nIAxeAudf/6Y+/GHgWWb4KM3zyjDDWBnRxG7X8RydN2H1Cl0SkIs6/3NPF85xAcEM14Z8S3W
8VjThU7aH2zXnT7P3RdwsYLXr+VomdKCndvBBl4Q69+0Ju4RL0A+GcLF48RIQO2rFa968dP2UUfz
1oovyQTaY7gkS1KJVLGPk71vnfpUY+oxAGv0QyCfzCe4HN0NUF8prYUUsIHr71yTROIoAIE/Ncwy
wmqxVP7M1Za6K+pbyJsdxCtas65XoboWmo3mWzPmnEHxsij57xjE3tqIxMHNZ3yRxlPoPaW/Awe5
7SycWSG5IUXKSCNaSwPvx1QTVDbFTgFz2uo5PMyJPpkyeFca7/obsed4HWkft9v0tuolRBbghDEJ
DKm3n97Rmm+bGIb4V/195CzQHmRZDmfouVZ9bq58SwW9uFT4Rg6xGw9xOMXK3SlobL+DG4W0T1uo
ywvmfOz195AEbxCcPIgXtV900zDeiZMwRWchzuwr9+i9TYlNKWifJ04GGv1R48K0+mOQ6OfQbnj4
w8CoMHlkNZ+wcUjyLc0vIULFlnWYaTMQ1U+Mnt3etTcLKcnmWDwn03cp4Rpool3IcOgk7YUfsKqF
FmDlm3d1xtL/7b69ZGB0DXQPtW0xfQwBdHcvmhjWMh0ZanrzNGvcDkC63V9Z/hkPq6IKuHUZIBDg
D+5giayibY6/Z56QwwmmeSEjGDJsbLPmGjqtrobiKzDWCQt5UGc7LkkrHsHR7Sz3iB9RRUu9Aoz8
pClxkknfNV8nmXBP+bRP1gNcQ/wTceg4zWHfvW5rKQ7wbvx5Jv7JOaBHuZWHmG681A2ryzjoKtAE
5rmNbU5V2bVt3J93HT16dvLMO0j9xwzOwAdfksLRWn+5zKSYARVC12UaTkMr23BK6/RR+7sruDAw
+KRAJa0LdvXJgpPR7IWAu1kzl/UEOGxoS9UVy643hHuVO+c++ZwMj615EthOPIe/05tsEOA1Jzca
Rd2o2ChByTqQjtaolba6JsL0I6AOZme275ppX7Ne0em1nWuTGxQ7Jcgy+mEBdNv6vYBRRBjUi8s5
TxvAg06pOJEOdp8kQu6yc7anpwJJBKI17S/zEQXunMljuT18Z9QPnJTPFygz7WYCSWBjcsRUISb9
mrqGmAtwiYR2QvsZ/7ATF97kLXvm938JM3IkvRiQ9e6p4Tsce0PdbjgPair/0itq5d+s/eWwmKhA
M6LaoztYbn3kdDfkiEQpHG9g5PczfqYiotZCoNgBfRwSqkoH5/e+kU3aBaDwXu4qRrOlDKyBYWuZ
wshxn5asukIO/BbcddKZlnre5z7ccamLloXuvZEY+02tUTVQYFiaQy6WFKf8BrOiuJckJxnpGbQn
tLqI+7YbsDIZ2BENp4b2EpjsIZhdsCj6P4NLuppcuSE85UV87wARjGa8tbAQ97wW4F2lgzqGn6UG
/LCGjpst9ynQd73jr7dofKfgfVpQmWYd38peLzGJDihkx3Jum0AiZ5u/M679Ier7B6Bl37hC+fZg
IofGuiSDcXSFxTl2XnIerRv0DTsk93kd6r9s9LOTmOCI+GfPNjYN+4/Z3gAgaPtv6cyntNyJwVgu
ueIN1uMly5vjBL0BI7QPyMcfrxj8ecwfjrvQTU0RZp7o9SO29mVrtLH2QKliNXbKNYS9PZbolmsH
2CTc6sMRXpFs1YyXple8N0HN88FDnAjFP95/GpbX8uinvM77SLOhUHVPdI5yVjEw8Quhm8Txqmlv
i39UoC6UYZN6dBjBmnKoE1JICT5XGFULbQAEiyL6w1yNyKTflMUX56iKn1U+V35JCb3FqF6AY1a7
7J3qv9kvvPxy5HfW5wJ8xGmKokWD8N0ikyW+oBtpD6JGx9WgYodz+NFgUWGICzOSUoQHz6zJLGbR
WfcoSRAatSjjzIA1rirObwdtcRjThviCfSkcV0x1iyFe30lvN1YZrKlrGnBwpW6/X89wEBrxY4j8
ZcCRTQzD1NlXnP2TCNek3MCCm/hesRgsE6HJUOV0Xvv5CZAUrh2wqzS6YmEbIb+LCzvLMbM1MDyL
UX91p3yaKDwCZIqMVK2pDWHS3SlHFof0ul2kNM+nWLNDL5g0VkkyWtNudhmWRHFeaFGo6xVZdUKQ
jarGC7f95ON9oEaAQMEjgMOvXAreNadwkxRopIV/kHJHxOvz8rqTgnM8xhVoLNETU4i4GpbqyVKr
NbFtawNQPzYA1uaYQrzw7QzKoK6wubii8LOJyZ7bfbOFnHkbpHO/Q8nWxom7lE+7suND9pCTyBJC
/MWIj8n/CI1zgky/jYP1UppJvo21oNzJgppP4K/vRyyUqVjTK5UlAx+7bPhxToxddnIPn7sD1m+Z
9Uy+dLNkA3X8Mz11M8Bv552698TVryMqwPNJQ4ib7SRNCSu5Gf07mPyXVoWxs3/iqB3cDd5NTcx/
Rj3BfVw9Cs9bN6X/0ISW7F3eLn7xh+cxWV8wMzXifuYqv3xgRaJp4sawycXJZapb1m+x3wIQbioJ
rH7lyABTiD7cT4aZdpgGT6MUh5q9LDticG763f3pOTdhjuv+7GWDsFwd6j6QPuhLMBxV9+p6/Acs
w3RU3sIJD3Q2dQhcb217dgSWqnA3kr+TQGcpnoVvYoOChC5eMg2J5pXpAybXBKLPqnNe4EAqggbx
hPf5QbOD7JJnfbjYkfKgGj5s9H1u8y4b95TnrQ67TcfRxXnGKXkD2S6VhBoOGhxhXPPbC+0rZDRg
wA4EsnB30cdhXRvlaQbY9gnSbL3BRHa4Rl8VZdHqzdrEB9/S2L40+SmzE/2mstiEojWK7CKZKNA5
0RcmkXYiw0xRkMQGEKRK8PYPPWJwTWPbRdqBhnMGg1U7JaVIiejh/NeHz11DmS05i/4I9NOsd1wi
44I9kqKA/iMc22L7mV6dJGKL2idwgQ9lMOcQte8VJ34xup0e+7uiCda2AOZy8cMxjU+i/5ZRaK2f
vj6E3Cz19ogcWYMW5Mucyb4LwetTYu1U9bT9/KrNfRcjBrHJNK6/eaMNKwefIne+ID+NYD4N4vEB
s3x4b8dcN7vg2aQ49Wn/4R5b2Hnk0hPM3opwO0G0GfKlDdkUxEMY2YvT8472U3m0Ft7tuMyt2ljj
s4sJE/44V0cA7RV5UmQ9sISBN0VpOMwAtehZttWV08TAmIIJDxOx4oMGTEGtl+4OMTr2hmH3OBDo
OC6wE5TkU6rPZQkn4NhXb9gdLIPZeOIx20kCOOs1yw3nZ81vU9H2uv8a3j11syGQtGTPea7mH16n
IGW6n8HniExnkJbWC/95wsb4rjPH0bJvnPfOmma1X8B7ih6dsBfY3asjWK/rphnrb/bHMyy+xi3L
TD3HjJbfR7Gpa5DGM9Ixef8KISzgsvGU4/z5C++95l8XuFwNexmHiUkG6J+yoSyuC6Jzo0tPFCr6
RCw1DX00w4Uzs5zMGqhsj2g5ZQlmbvZX+0Iczi5ju/8PI3o+EXmQb5wOG9cA5sZh8rLo65I8YZWQ
U3iUPOFt2JU8wnSrhP/ja8zYQO+2sIiXuPCB6AVtyxUBYBtSn3ye0wpquXIX0PxHBQzI7pPyHzUT
3q1dFT6f3erofE1g+e2YBn8O9vWk4ZX/vJxRQaZ+GLGuSwV3KimJYCwFhWUQzSFCSmhxr7yZy2iw
BwrfzLOymUiigCRmZNWi7kU2m0NuWZXQlCBW3zNKV1vUWpbfoqXXPn9yHCZwhiu3cX92Yhowuo0K
qWufC41mDmW8MFtMckU318BxWCsF+xxaiuZhLSbdXQNQyOlEuhGyeE/xWndh7jffaOI0o00tbm9E
nHbq23RVrSWV5j7hq7K10SngVBhKiHNA35Izq61d+meDTgJOqq7m8d4TYB0JrsUxVDVKKnPW6ZYN
sP20a/hhhPmjkLSjaW2jSBqqKlGt9Bl0Ff9+K+RngEED16reRIwryQ/owcLXDWGsydyHlU8A7Ykz
Rad45IoSC0EZnM/uP3zs40tMoNZIWPA7FLGekpw5Z0xGrmFroq399En4JRVWWIwTKk8ZdltH2W4U
NMVAvcn1h2AWGXrrlXG96zthjx1HkNFhkncCxUNO6kELn7jw8DCZoz5hbMiCX10XW4zYIyblKtjN
y6pHgYH5uzl+pukUpVSnRLlurG0A0gaxt1P9edYIm3pXqI4Av9X7liFAz6rESFI/Yp/EKvVBAO2v
epvnnTkx1+7TxKu7cxTgAeqB6nFDqlGcoMNVX8gapKBbShdoyex6i9//GE/lsQEleyMZLXwkN0Ju
tUIjFzxd+otiVFEtlOd0JNYgKoCMISUeS9LOe9wd5O+PhDQ/qLGlo/9l+186cs0dnlQoPSZP03h4
I/wb9hswAHNKsBw8HaTfwOylgi+EwuxeJPhynRl2qWqpCagSiYjTA656o8oOlx0nMI1bblTIk4t/
MV6EvRiWVupiv8T2Nj+oMn5Fx6aQVDcp2+3gTfT9WDEx4cNy7TVR5Pv6p9qMJ8A0j5dFMEOJJNDU
6NaNKsYb9xIsdBbI0KqHyZ+tujyj9KVNP8D9LRaewb+sdxcxdaGD/fsodrI9Z5Z+o+RAeyc3oPuE
WO/ccyFFdpHey+Lvj59nVZcTxg8HiWZLmsB2cw7G8DYLcz2srMCCyYMVyUeVNpOmk2ysy/1B78Wk
nn19ukFNp/aJIP/b8F40CjV1OfDM0rNZhsRVWowYeOJY980a0aRm6/PoLnAlY4fy6K2e+sOZi85j
qFl3XAahfviMvXlSdgcFvx2gX5DfXB8P5sSJYB9LpIwwFyJMIFo0+4W88eYjVI++T8BjVgZ59Qqz
SgKOED5f6IDpk+BJ6uv3edRr3EQkTdUnDUzN/Bya8+BiY8CuczVJJv8L/Gm7r+HOlp6M0TVVbND4
3BJnltovEIRgbR96pSdrj2E9cKN395hPEEQkziJb//B16P+dMLcTH5qJl2DLZL0uGFq79a/dsgav
tVXh48biuK7J+/jKaf69ir5uXg1LGaGcxHXhVo7USiguTP/XD7qtOHb2nkEEFLF0T7TctcU2afl7
Q3tgiwLDoQKOXvqd6J5VzWshtHITngGVTBMB5+fssdmBdYDh4DEARmJ1hQjJL8B53heC31iB/+OY
G32MN4kMDgNgZCcFUk2vxQEu8Y/WbrRb1goSWX/jDkJsxmutndJmw6LqBzyfPHDTdxjCmPE31voY
uvTJs/NGuoMvQz3I+s0TmTPiokZ11NlJHOghCK8953MHIFSgJgR7nb2uM4+xwZ4OdvqZ2FdePDeT
RVxG2eWOhtsshF5uNksHrDW2ERMyDStRxeSxuP/rWNRNnpAa1FJwVj3etQ9I1R2FphbPEY/wqFhX
JugP2tFEipctdx9w4mqckV2LM7XdOA/v7vDuJexZM1WmQbBn2aGR5+m6SzO0b0FeOqQk7ng/qjUw
DJ/n+3+CA1JoDJL555omZLwKK/rn2sqQnzHE6EdHw67bqfx6R34lHvZa6OuEyWdX9z7miN5WADug
Olsuasto8ef0AuNYaSmUoeh5nfO3rA4RXVJdzSuZiRI6Tnc7GmZbp1UB4OIJm3PojtzLIuuoRkAG
1OB1WpXaIh5VzzzF+sfY75QmRlWFjqMHez93rhzmey8SGQ4XFaYMebfq6vyQR6zwVI6EhN0+uRbH
unD6nXb4Hu2p4dAo5ZIurzBSvBBSg4YMUxXHJlj0e+Kw08L9DLjAQvjwq0aHAZjjt6WHVDghcIq+
akAhaWEsjLXrN2LvYmkDJQrR9d/n67Nj0HXlL7RQfeos+ROnhNFW++1nnk26kPmyNPHPJFSJuLrQ
B6JboqiKJvIdmQd8b2bApU/tD/3h8eHglJLrpd1vuDxvlvhZDfoIzFOaPvFCXggLO0rsXFg+Ze4j
0Qm6hFv/yAdLXHhykZrqbBDJItOAwSI1E0De/glXQocmSFiUYUL49dzDpDenLUc/p+MQyQvEsHyv
Yk+iY98r/7RYdhDJXvy0jgS0KrT+MPndBB2KmtVPGHxmVjMTQudZoFL6yV5tLCTM55Tnjcg8UFL3
6djLtScujO1nH6xr6V3aIPOs7TDh4LhHPmlFbo/d2BHvk+zy4ykAf1oqWWKqrJdFiBplhSqbj45P
9QEK/8gLL8zfcoDRYSVP9a7eg1UqQUR+9C6w+U44ehbDaucwDi1P+MFGfsqnpaqfDPeBCyMY0gs1
tBoiz0bSc8/SEZm+Y6TjN7PiYemuryB7JDXQfhftOQYMz/4cQc+MizAQYRF2jW6ZdceQL3wxgRXb
Nt1+OCi85xaJGH9DbguwgsC7PRSidrX0FaFyH3uXWN5nheHH0JCBNuvu3NaTCWs9R0fWKH7ttJD5
mm9ACQ9frW9SuTSkst1zrI7H9zIca41WAaiUl9chs0yQ34V78efUk4lKZSpEDCrhpbno4RSooUVr
d+kSzfYWJdfWGrhuLPhLQ7CXPf6+zIyF0YUOx/HsAE2XyIHKODO4wwntmWtyT2y2G/NB8Nzfckhu
sdBD/1Y1ro1dHiF6pnDDqEPQV0blio0opO6pv4aW8w3tWZ+q/IU7R3dcf5j0u1ahgRNFQxRhxoPn
C3CF1QhFpdF9tblJwtdOG5WYgYsnrycgFep0/nWOF8sO01eGYeg4dfN3LT3wOEi7kn78mmD0VpmI
6PxOz9qcDP+7Q+q0hH1GbP6n5udnRz9Tk/VLfkLnXWGsz0+XeflYFLZZAnY+tZKHpxmqDRjMyvK0
hZ2AJA5++9HSF+xzYwzs0YAMR/mBLDu6zD922+cPv2zuLYtBwXlyNsPjke+3/mr5/oKhy+5K2Mep
cYkn5iH4+M2u0uhjvi1Z0uBwRuKb+tkeyomkUjDP7LUndaon+9sY7UZu4o7Z1Lr4eSVacHNQaQk4
9RHlxTCZAgoijS9omjQtTZzMLZz/n4Qd94sheDLBm8DdDemuB+iiOWiU8e4+qU8Sacyfv8bMXzcw
0Z3kK5O8v6TRQ9tfIrSa3OCVGRcNTuSNHizaSNE39Mkc80kZ7lzbTAIa7CKrva1tjAUIJ1JbOPBu
/pDIhxoAduVclrYMa/5IKnjefFXn6DjkJJ2Jxq3mD0RbiX9nbV0tvl6TI5j1vewT3pFhctrVjFpd
3IrVUxppb/mCUrLDvBo+RKwdwdjcPNRhhvVm/ZuSDc/YBXzKAcrLtLQlHMnZ1pNIVZbKcvnxmi1h
6SLZND2hLe1533RjWOUIG0nUwkDDln2NW4xfKBcHIJl+2IKY9GWrbkk7tWdXMrFpOZUuEq3eM2yO
OS/lvFLbcicp6KZ5zncIhXSMmi9PnPUPrbXRNVZ9/IqmuvfHjmdz0/11gOyUPSEp2HwkOi4DWUNC
5Al7vklGPCsyFf0B8L300aXu8PyTYjjRUJanzl5Ym+682L/rJGKS/j9rLXXSo+kX15BRb/yjcAl+
ir2XsJ929CyGt9RVeb29GEXncGTVrNi61Bb6gzAP5G4Od5PH4fbI6uJyayVgyrbkQw01umE0nUbL
tUWet/fvL85fyku902TnY71vPyxjCPcn1doQW7CkM+gpBOE1X8U7PDK24MRdCf5wl+VmdW66ypKS
Q5rizUWTxdo3zsz0DzM62wnTsDz89FYj7vmfrI4pLkioDf4exlku1po/JWPhekGzXbL1x1XMDfII
m/O68pNVhGGDjA5yDGITF/GvB33RdCfRsYEbnQ5JwQoiq3SzUYrtHPEWD8hLBpB3YKx8wCDp7f5m
AvG5aGh9FKom0UawZ+MoQPfdro/fBg4k4n63CF4kQwDQ7FTSH8Up/RVfMpIC1CaccgyCBp5AV7XR
6JF21eD6a42EVt8kuUzfqKtlTVpuOprFooHZ+glocWIRqB/VORvnQi+b85oaPuURFq5gOZYP7VBa
3V2JRu7iEZ+Suo7NqMljMzCHhrDNfCewOzJTjv3eQfUqS1y111b4TZUEAN6yCHOCRVFu/OLqixI8
eFhTzW5dYihNoQZyKjTIH5XTeYSvYgISNy8q+3vqTLkJOFxjyL0JLphf93VI6eX0G9OmC0a1f6wB
E5q14Zj5wTC4igJ/B9i/hVNf5dPSPr7WfeB+K6T8FkEGYXnSSk5ofEAUoVtQjhcRKBgH69HcLuuA
Lb89++ossSD2U9lb1qxZ64VxsXIaR5uTksHASCE76kxT6AZOfbRRAE6bseaE7dW2hZyO9gnGcHg1
6pxHghM9gib1TcrnYbfQzoAhQ0eTlp06UgRZ6JpXyPxtN09eJCMMM6npLjCUsQ4BzALxm+Es+zvS
KpqRIlMxclTKNhbcuYL/gPvw/LPyvWD3w/LQz+mitaH8YxjOUzgjd8WSotPHXv4rvQnqZs4gErFB
xn3doMZruhri7GIvQGO5L/gZq+kwmyV28pMvXHNFGVnR1Z0RS/4CCEDBFOXJIewk1Lttas3uJEwZ
qJXAVFajQeWNKCerwc0k3R0hUudkv3y9tgx0UflrtH4ugocgVoU9qbZ9qwpwBdTN311ifS7u7IQK
mBZk/kxKLnp0Xew81pc4F94yxMo2mQIBFn2pGfat9JtybGjqdVh22FzkjSBZiJRODzVH1Bx0AWPs
+mJY9D0Tib+9GCGseHKVb0iNa0aYU3/wJUakMEmnasBtvDRNP6/6P12GModpF48nV7D+NyM4+Uih
ljE0oMQY8zRGYCC8MvFq4DUb8Pm3IJWULsBhKEYc3B+i9W19LRghSTxmdd5S+B1n9f8xzhqL1Nyb
dSSlutWcaIwM3k8VH1UbWL9ph/9CJsjmvWvXBQn2NRyZrjuMifNqBUwP+WGnl4D4DC52zgg2Hvtz
J+RLU2j90IT3ayqHHnw+AaNaVCWg48I3jnVMD9h8QLNtKhyj1IODTcqHiHrF3qrKZPyt/EzAKdkR
9iOB5yEqtMPRW/PqCeeWr3/W93IEAp5/stnrGA9dIfOhxu5uJu4XAScPH6cUFlOD4Dxwi/H3fYUg
8E4YuAnCvVKBormxwJpc3GZQbJKbSHQpAAwr0+Kwq2FUEg4hx68Iy1waZTZoJ9MxyRyzO/mqT8le
E3Vx4nYl3p/4yypOi/bBEe1+HA88DVp17aZj+7f/Bks4HcAkmlL1Mz/vk1Q3rdnkPAGMxoVD9/nr
eGD1gaVBXBkC4bMOXYbxkuSXV8E3nMQAk6GpyPbZNUqa8K/EBAt6GowWABPausiIeIzvcKXJexeT
CONK8+KG/OxG+un+bzQh/wmUnGYCBYKUgPzwf9fBgZIr0oX0xocG0a/ZFk4h2mMVBhoFWIFKxaOO
Ag9DhK5jSHh+Fgv2FSAULDkeObKvDB+H96ivdr8VVHqqrTmuIrGFJr1GW4JVfqAewXjpJ0QA15sS
TQ0kK6k9k6o5PtzJwAMe2EafbQA49iT7f3Wup5XE8gAFtKheYsxFMqXY+0odk5buEOIvrudqjbSG
H/4zDGKY3upY3hatwfBI2cnjkxm3dImtrNj9pP19yX2xO6wTXDJxXVycmckGvVtVwE65/xSZripZ
777dlgdkXR+Q5u/M8fTIgcEl5YjjZ2ZzP71ojMAK/9ZUAcwWIpHnrLhWueMdNfFTm6WuTr2zogCk
No6JRrDxlvm8wgtzlorzTU71viiPan9U4K5ieflp4yZaGgvxgStKIpPtRpCnRnqelBDS+CQ5pfv3
RRa1ijLsy+9oRyAmry1Ja87rtKTvubv//N+8ByqYmCzOa56CmUj9kTSkTfmbIoKj7t1AykgN09w5
ZPj5wBdBqCjZtm4O7tgNaAkQ8Vj/chzILFdVVwgChItD3LaSs0n8eyW1byNCCcaxK1JgahxUTBjc
WgPcnsgaVFbwYzybmvrgswUiVlx4fNDjlHdTzkR2i7uAgS5xx7ZEKAbyT+sDohaZ+28l9LHsQwzH
ovGxY6uwTPc7aok4givQKcAdF7/P8kZu8saPLcuiyG3QhG69AVYBqRnBFkPZnBL9AialWSKttMRn
FfAo4xUob2XKRNZKNYdBotQaydazckW/v4huUhi+t28eYzk1luiCjqZ3m0dRRAEu9v8yUbUvuMnk
OQGhXEugA0UZLBkwiZ62McHktindfo76qtxfPKk+pJYzvMC3yL0Gm/YAG3mxxLXCEgHB8pDSK0Vb
llTge5Cjy1h3qMmPLHAYBE5dpjA2EkTzOKiI+qnIlUvzpoAwnqD/Iq+9qXRcv4Ax/rzLQn7cNFHU
2/gygFfKG1OuRCWi6z8l9Ob2+2FZyjks+8r7emeuPhEP1UdPEttqur8D2TmQiD0jAUqDxVEfA3YL
ubUTJkHjAzXq5V8VUKZ9K4xhbyO75vnwCegDEWo4mJMeMLgggE8UOk7fsI6i11iyF3ivvY8BpXZf
JDSRoZ6hTptqberTtJVaOZ8oMGdDvETIN1LYhjiLvcstPPgpzfx2qgypc88dbQAt+DcBuy5FMBeA
inJVQebicaQVUf3t5mV2HTLCPDWKPP8Twl6UpT5mBfRwfPhscssssVNlMqdmYQMz4+93Tabsyi/2
Y50UKPGaw7pkG70FYdSdSWe9ZNCZkxhDWKX3jLY8x4tM7uOjA9rusVQqzqDCIog7ZyNvUzd50aNp
ATUkwWbFsrJyYRz4lUa/5qMZlfeYEF2FKpVEkw4Cv74ApY4It5jDZrNfcWuUuxuSeiRo24POgzy+
VAxW7YULquhvbZztpTPY4c0FKa/4+9lwVZyG/ASX2jpD2RpVtWk1v/vBGxqD2K9yDdZdoSbhADT2
J2KpOxG4o3xo9+TAkx9mtOwYm1ZuXtOf2rqRby23x2EMYtSVPp8q+4VKSankE1v+ZORgS/3xdcpu
YV8UWpjSDqp3luxU+v+fqGyXeTQkBvYjl4P57b5TdtBW6lc8v1mHjDnslxY5oeYk6BeCEFWacFBv
2KvVZ/omJDXygpFQyPMojNKX4iImC3nLlrb10prNZLcn3pxzjawyHpadBUYr9B2mGW0oVZs4/enH
syhTCeDQG9SU+Et1Yhpz7BuTGA4PvD0VfdzFm/vssCxz3CRusHmaekei2AUi5YZlU1hfdO7fXsRV
RFolX5rCnew6Rlly/9QfrQnnuwZsYMFH2AMuYasleCtGcRJ2pYXGpZs7VoEvKqZYeKyIayoJw1Vw
nWJRrX87i1AV4GAbMOAqusN+B5ginvhUM97exIJZSsDWn83RUYngINiKFFfyX/ayz9Ng8Cz58KHW
0HRsfW95TRIkzVupIOtDgeSAdwk8hjmehnsx7eTe6dj/hqDPX3MSHfDSyajLpSoflmjjfYDeOZDF
JrV+nvLHiMOXfS22Eu883qVmfxEnQpI1LIAKrkUl8F4/F+UmIfKHEpZEtFQAfrxMJridGD+3Xixl
5+vUGiW5dB6zCcoIM5AvmPGufu+etCf1E05j8+TuiBvkI4ih6Nm7eA2tOsvo2Vlmrl7QJX2/4xmf
api4/0mdMGmAFt0LBOY34tuqw7mEQ7hT8SitNKpIzxH7CSI3Xg4CxSGIVCaYOaiS9bu7naVABk9D
kJJGM703PxMuILYw856bhswapGMpAXluWQOtNPbxVQ+kLvrC683aIkm9reTDKYmLsavAKGvwpIkx
akxd9iK5JYwioOnykfRozXwpvRFAalSrg3JrLyMJrvNb5iFN0GGTFjlkPl1cFo9kGO7c4WlKMj8m
6fPXHnZVlPmZeLGvTn4SsEa+0GUVU6YQwh8vJVEuWMUglU2T/JlzehNybLcEs2+JrWoBnHx0+7y6
fegY/qDpTNbW/WwgAXEajPoJSxMrD8lDO3KBvbgJelLccxifECp0y6Sl/uvgAlxr/ojkkGO1R4PZ
8wrRrMp9SM0/pi2gJva4KaggJx0GXlHdMoEyBCpy0QGlClA4hyLAO+7OHwJ8926eGABU3i0HsSNC
pREUfdSU5TplDHopkVFL4DecBIXv12WV8s5uxk+KLJubryfrnsW744BQ3yz1qizBjjcOfBdc2naR
WSX7BPuGlassBohhNlpGvoNTOeTCkSYudLkn/pHYJLzJ4PmeTGG5vMur1vhCyoblAcESXTPhlW8y
tyFmZ0GBIDx57v7g7YZjSsX4KovitckuTUkFi0HRObKLQKNjJk7X75nYYuOvCWNyYNkXv9Ngpgmo
8YNWH/tXwKMqdBCP/hxi3eeaHTbBNW0M1ApwME0x8XCfuiTvkXvmxtZbykebiAnm6TA8rOsZR2r0
oRregJmDsyyti8fW2laRG3OpqYO+BVc7M5wUmSxklst/QyZ/Rmizy2xOWV5A7V+9O2xKGffJDImd
7tsM0fNjLcWNBb9vHnyADlZoa82YJjrthOUE+o7rzzHKvnm+aeGIr9qv0A8nucC2duXrmrp8NtE7
5P6MbRHh4yVohYIGp48/ztBkDRtLu+5i2nmFPd97xpdl+wH4VyUBxiXh7Lik0Ef0FDpVrWg+WzyN
QK9ZHasPFzJLazMmD02Xuue/vPcbe/OFIUeYUJ1MrJGVy6k7BcABMGQddTCz7KDg1kCiQygDkbD3
SP3DXp9EM43lwtLYbfUlHOtJnKGgug/7PW7GeDuj6qJWw7YxMHfCOaYdlIHsXlyZJ6vKQnzbH6TD
BEuTrb57eRCf1cZ0Cwj9LfBwjYD2z1QMBz8mYJT9gQ/eumV6E8rxZnoSuQIrnhSKXpJQSOLddIzs
/s+oNA13nGUWCVVT14+IVLAHWzBHrUq5vDtPU82Y/1VYRB2Slb8W2jVgCIuP+/DGses0ajS2VOZ1
dxzD+OBeMTjwXUFKn/eYR4kZsHaae+dV5UbGQ6Jc8G9lN6IyC7cbF3fw/uftkXFwbp7m1y5hlpEt
uLf8rzYn8IRePkmmfGq4S7nyEryjp5hGyEAMfOwdRr2Xai36R0K4d+tNYCq5rQsQWPH+5bzKfTun
+u4fc4crhpFaikuNrPWjlDsU4zC25mYVUvTF8jmb7corn0SB6UwKbZk/Etzfss+qZHn9eFUOQvNm
1WewBRorA2UU7bSrA1Z7p9DORDIhaeC9tZKEvhgXUOs/E0Iu/2+FC+Hvs3AaQC5+xsyAzGfclLQ8
r1VyQIo6eDE97v6L8Z/haxYZKWo33PqMrd13SpvR4jucPD956pGBOYA3w04cJGj2WOBP3gXGtkSj
tx36c+xXZyXnqsff1kiQ9ErdbJ2j8FyHZ1dCdIRH/e7yi+ZCMlJ+UxVfdVRqFBE2CcP83pwl4kLS
X1Dxlh5zf/tYTJNXpVwHOIzOgdHBpSet04gsdEFIBOvmf6s+ZDOvlFhCK4Eol22GtJCuLn1HvEWa
cBgEgQ8qW5qOSG9ZW9oyq5LLylzikCYcgJeJlJZiU9YcUs6LJgD+zf6kPDruR+1TXlHEwYWc9Qfj
80NR2rhdWWOcc59dpUZtd1Q+T4W9ic/CI9yCErz8oxOigKlG50QnjB4PNuCxIgSxZvdrLnklwgKE
mqsn8X7uHNDpffKBjv52txk7Ww4knWcR6FdxOvGWfQEbMCvuc6hKVHeO5GW3iqNNBMliCZQ3ZKlO
ecbkIild2fNbpBkNUjh4gtLTuQZgBldDUK362wWK2rqZo3fbrslWTKvMhRoMoibrbEPyQNvOcAZB
CReV+IYZgKNi21tg35NLlUW7oPFEyEzW3V6yR5vnEcAp26vzNHIr+ZsnybOBuNYcu1BX8JgiwmF7
RY8LQSTpHoRvO1hl4fkwePMqX0xij9uThiV2z7cvbb68T0GsMHrx3hDWH71nkh22ddNpaAv7GAVL
KNvZvNr7ToaBdx+6VnjBydkmISmJdj5fxG57AJTVda7shNMNXkJW+mt8hC8ySQVN91jvQAb5uFip
FMT3z9x6YwgCMNVlD5zpnonws4nNvcC6viXGHrUUdNNguxoQ78EJ3YNhtj7RD56zvZw3OBxvmIEC
B+nzaBY1gBouu+llpRLSOUgFbF8BQLpEli9oxDsOy7MupFO6XzvyaBcQRZULZA/vzUTlvcSZ5ham
WcS+r4ncSVoAR40ipO8B6r5GMb5R3vI6pbY9hYkArO5MOCJ/qk+mnqnilNL6Sqgqs4zCwlLbD+uP
1FdUd5hpdVAq+YykCRIZp0MyKs/pQzaZ9l9Nar3YF9ooMn5ldau8+4yPl6sN//AD7lynzDq5RrW+
ZIblKeGzV12UhGD70wyJ0G29UB/XPkGj2qnv2Nex8MSqSMFKdI4sjQcZ8R/YOMJwjYk9DzGJf0B7
49lF/VTOspE5itGhTQsKB1lTddr+B1MpmsnsACkCzWFmEUu3aeCoh9Rx/i+PBlbL5GApVLIP3uC3
4Bcou/YfE8fEtQGqsOif3B2NxjIMyQ/aqRCbRE39YyWnVVOsRypuwa/1nMN2zDdZq7Oe32QsJSBG
nNaJv9GeUQYcmYJMoL5RTZFcC5DOd9zDH3QpMpv//E6t77MW+stlS32bRPtcceT8zu9wHOHvdrKc
ILKuMRIf1CXln2BJkkLyd9w0uDlbi+yhBuNrtmU+rLqgUXsErC1qqm2vXSmU1JEYP6Ey3oynh5UR
ab9T7wtsWaYpXpUrcG7ui/087VwD1ejx0Tg77RM6NfiIryBn0+Wg3Xq+XWC315dQE27m7h89zS6A
0l4PCmhJz+RRFKgt6W7We4myRLrMS05KCvd/oLHbKdz26IMh1igIS3MIVQxwn2uEOdaZeIKjxBxR
Pn8Vbzm+LcNxqFJXRerOOf3WQbVWmFVxGOk23cpgWchmH685o9TlxeZ/qL4JvEa7K4SIRDIehs4l
5k6c9/RBZugX/ruP+dgvgfzVg71Zzcj57CPkmkHsX6seFXvprssS3JOS+ebLRnmaeHCZMrWjqf/0
Mv3WGPzeMYeHF3ixNbdc+QTjxsK+9y7UWCRw1aPx63+77McCDmrcHiwWjU62WiR740DZED+g+aL+
Zrr4FXd6i+fMNy392XEzkfI7cplicPC9/uPsHzxUMMVE1z+lmsl3sQSYdhtlAGiQRvlDGX7JKP+9
Cp4Z+uii797QC0tupsqluUykJIpt52ZEcu+V4jtQC5vHoqPNPnzhceQ2gBAvH3R0i6UcnSWmUD3B
VxgBqltTiDPdcJUTfiFtNVwbuv+xJK/KosR5xD26BXF3w5TILVqMfT3TZcg6rdGfhtaEz4B9ig8r
VElRur63Vwx9F8uAeiyFqz7SgLR2K3jXDa2UeaJmWHH6KaXsXer9VLBWQ+tJzgV3In0jP0cgfxGl
QJXJsUck9NuQHyNiX8XBqDHQNxin/AhaGLkL2Y3ycCSvlGcFT7N2eBjeknpzJyhkKiY8qxJSNK3q
0JbD3pdzuNjZFFlWe8TJNbwQgOifweYOrkrJ/5p14M4l1ZxKMRfcZnB05REsSktmnlS+301Lu6kZ
1aFZJmKrHLUeOE149GcQ6HN0QcKHTcNDSKMbPYJPqTFjzTiB6l3siae9YebfOq0hTVWDowE1YTqx
zX08LkRW8XVxtM4T99NkQyPCeVmRwweX9qQqR6c6QOUWcPr5VrR6I0QZJw7g/7esTlyUPo8K9/IE
k1FCgYR2Y/G7zlFcic06Re6dZzDdgUw9ThhLfYyneysnbC2lWIte6nign2Dg/QOKgIbRK/2M+jRj
qFuxKWEij8Mi0ti3V1klRi4slTGP+QNx1TMK1Stda3mej9Ion5GoNidWF8Hf9sPrnj4yPpHQW1gI
2YXjIG7S98kx9xkQ0u5dTs6pVl+Ovq7gF/21xu3kkVjmkhosiznPEuxn1zkwnBGjgS3krh5izqg0
A43E7FqU4F01bvgB1Vu56oTwruJCDuS6LHCAjT4p/eP/t70zfSTOQiyCj5pmeSEJsWObOc+LbDA7
dGtZF3DnWmcNu82QjUOINfqAmeTez7psrc8No42SoObwb9mwmglWpS2av2oerrsx5kDGg6HjVMnw
+Z6HUllmsM3VhbrSyCQURUljNp8RgHiXf/AssRlSIv/wFDgnotVl4wN6N7h8kayLkew9O96qCVpP
PpFDZxAAAuAOjPWrAwF6H71xdmWX3fM2P80J3kgj/rfTNzMvhTNCT84Sn2Z/j6Pvv49xGNdBOzjy
Rc8248WMYoz81Y3Ld/WiGxlS7Ua/9h36b4VhZxw3VwS2p58/3GqarIQWNnGQHyN/pAFkyqWflKc+
p0Yu2ygaqJGkB52ABJSzzSCqojdPPWRkInOWqIPWS1SrWCJ3p/C6taYvoNOPD14BGEvZNFnio+wG
/CxkLtwRSIR1ahHyQEvTEuQ58yvAWPCsZY6XuQ1fU4o5FXzAgkoCcxGWS7vq8lzVIdAyogAjGI5b
y9G4KMUpHc8an8cJJGXgVMpX3DBwc+7IF1kQIIsWTW9xo6gchQ9ZgtiToJUHt27EH6se1WWYKGli
S2SfVGehZ0ZIsqTHozgA/UZoUKGK99UoM33SxhwVOfuQ8THHFwcxud9wj8bkOMeoXoDj0rQKYelu
Bi7iepoX7ZRwOLCf1YF0kvebEehx7BU1HodxwgTbNBWnLMkE6NR3U/jiwADRdxRjt7JBrpE2g77c
rBI6d56A7ffFsVSPWd2Z7Q79zZ5lxoOoiyOihWqQLdxV0PyxNQ8Ub1t/0E+cQxge9OcXTjUcFxVz
9uVK8X6EJNsDcdRhyj69sjkjIwBczRouH7Xi/9sk1Z+Pq690guUsCJUm5exWUWU1H5MrbvNbT/i1
fNOyOFQTehTs6pMZSnHcqbPli0T+NI2nEBxaVOQnIbkErpcbQF/B2pluCx3VOYSe2OJ59jHv78JG
ptFVaFT/WdJZYCWFWNEcpjW4vz0cU+KdIgzEpqK0kPSGPByWsTz4H81cnOBPVyGGL6RBbKJZOFSu
yR1HNVlMoPvMz0b0WGBGbv1R5ZS00BIiplhNrELhlP7i84KaN6ncgMdkOugEp9cZcEjnt1D06L34
1DMeWPojECwhvEnbWgxrPTmYkdyPw7fRC9aeIIW2ztuUyxXbfRI752sWHulgK5rNbEke/nFO/md+
Es7QKi9LnFp1+5HzYJCPFCNW59Socikqi1c83TxAcAXZtuna9gMWrxTfsG7XBLpJdy7MG49CfRnh
EVZuXVvdfZ8vXkrHPhEV6n/q/eIZVaQ5LLvbWAYXjh0jr6IlQXxwQTnInOCaAjqy6fJUcn/b3Ig7
bBj8ziq8+nbDOIDNRXnUSZwi4A5jwohjDciSZP1MLXEhrdep25+kAyG5a3qlhQH1KR/ur208YKkj
hhl733Kc09dv8KalObYjETljX9PxEGnTmp0uoBo7k/TEmui5/uNJUYzOdAkmXB+f1FEBvYvlUiBk
9FimGsS86gmglQslXwTdVWBKWX8uh8HEcWk7RPC8MkRE7hofgctIv71Se5yef6E4Ii61/zeOylPK
yX5qhnNezDiGbYZF+XNQse8r2FWT4uCOtoYqQZZS9KSKlP3Ko+Z4dzLbHPrg/NcN03QG+atspPUk
M2CXXzt+YEISiZVEIGmJN+P4fstEK4Do8RW3dgSEkWl0eya6fi1sxOEnnSS5n1qxK1dcoCXJHAXk
A9CBHlD3MZP6rgRqxB4YK/xjRUd+WU/BL7selyyt9tjA8knxsiSu5fENkzJaIFTcJQT3aEKzKT6B
1mVIlnn5DDpF326iBCeOj0ew4iJ5Os0yHE9HIAA1mSnFApdBmVDXRuO2ZA7S+ET8/TJPJtJ4ulDf
ckJ8YFOxPTVUgujWN+Iph/SGM9g9MIr3U2hYebCAzYhlXIL2UIDQDNAeXh3JJq8gwHzQa7xQBV4j
xYp6bRuq5k8KEDLOBEqZ26fi4zSXxJ2OLZtzgkJLTbhbjgLy3bv7g5V5invKzVM7Ir/rBIeefGZN
rd9gmUpInkJTEHVejXYlVTg9SYOClGoqfDECn36/Bbp1wXOTuLJn2xko6y1hdagV4TBTPRkoBdGk
mDDks8K93U9EGK1ovxYUtidYz8CnYNfNEbyDvNZO1f/OmgyFmC1Epa6rVRBmh4c2QZkjFoHVi8YY
ZFxDzzyg5U58OuaiCWL+JpdDDMDqqkvOAGS/h76Hjwr1oYZgtsV0BiXaxjjv68y1FQKkndt0B5HJ
0a9N92b855eCE2rB0DYkt5bPOP1yoPCQJGydyusuTbk2nAXmp3J+E8TeAF2s6QKyob56o0mrAK3o
bRX33lAczAz5oiPx+lFbv8qGyoBsjYnCsoO4n88EJ3GouxXMnztXjQGeB5e60knuF/QTvQSr5h00
gATaz9LazEvBcaQ4urhq7hUGZwiNeaHu/NxPQVUYgINB1MrjPrBiXnA8JqOko+Eiya6HIgaACyyv
UP3lpRTHJOugx2r3n02zqWp4FJRP7quDHgV5lvEAT/pi6WlsLaX+r6KbFSmAZ36+Fp4Uv0Mrwr07
bvEAkGlAJ5x7cRFLRMWknsw8R1MqwMguoaqyxwhNnf0Y/hhXpqukNTjEH3J/iid+99RQhkdKV0xw
PhYQeDGYIqDt8ru0mhKhlAaSOapR6g8glkkXYJd2oHOX6hHBwNJulfFj1RA1GFdhZDV8nZp3PNaR
lHoZ3vwjstBCO3zG746K1XuQvCdQiBHZ0qcMpvYhxZrchcpSsrmyjboAhn6wZKHKMSGp8O2+YMOZ
eoJZjUd6zZaFYL/L6hVWjCOhKFim6t28WNKlQsxmCniS1S5jSHDN1fXErm6qZtlZZS/UIdzfh73r
BbEpWry7arpfONTZ2B8rl347xrOytjhyQcycJwE512Akc2cj2poagaxh2MI6fPPVyKE3jGELnkYX
WfyTi9g7/BkBmnWER0ABw2ersl2ldIK/yGQ59o48aYYQ5sfSSfmaOqZD1lliEK+aqdNefaQtbsGy
4qztN5AjqsZyMelXh6I4CgLhsq1GPjvVSn2zBkdt8PY77xWQ0t6G30t34QXE2vuzDhqR/hA56QL7
wsB/xGutD/6Fh1UBDvqfghPvWvk4gyyDatDHMHW4o2tgQCHJPuS0wUZnn5ruCZYIKu/rKi9ZINBl
E3lX9mvC8n6UnQEy8tQtxUHLpHkHQa/lI4gGI2PH2EyZ4GdEG2mfL3KQIsGDryaAQ3kOQnK6OISH
s0yJcPzy6pGS3ai17vpuNyxG9TtSvSylpCg9FK4QA6gnmhLsb4/SrzDt4fXpF1hmX/uc1bvqdWMu
totGP+Skds38QRiODofUi9TCEHfndA0SZpldrDE+JAoSnMFAkEbLfGMpGjFnQGzRW3BnHJc8gMdv
eggX9Ync7AR75Z/HmfuRtkNQRUyvOQUThfMRp1HMwuEF0eTyetDi082hsrLK9oUDleTqw0myBP5Z
unosRzk5sXXmPhDWuzuPUWRuLhFDOrFTrO3bKGnu8bG/yR1Z1eXbjxwox6AbJNXwOLN8ff5Clb2K
afUs9ucYct5rd/wyMGv5TmonlDSoC7TPEh016F3MV8fOty8SEuorL/JntcJ6tuLSZ6yUH7kcwzAv
tMGjEXrZwguCFCRVn8V2QvYrzjPeLfRODveFLLDjy/YsZU9OU8BVsXjp/pus3jFzX1xLaF0sVQJx
WkN4zaDWkSpAUbLYVkkJePbZO6rcI3yOmklhSfhROaW+eTKFegHgqhLtP0PprwO7QyLPTD/kr3T4
cXvLElRK65SJW/b55MJOKnsckgfbxDTiGMhLD6Xg6gHwc51KCf2+Lya8RHvtk83xrjPz5N4gVief
FyLCMVvkUhS0juudia5NVZLb7HEDoE1GF4dqt+kGiH3FubvT1r9TXICWpN2DgXV8uu7CoG85/5cp
94JtNY78J+vl3sikY9loNgBy1I2qEyYq73HhxdXWsgGm7SycaUQeHpNE6ta+E0MpT3JAo2ZaB4Pp
IKkvWmkmA1A7aXAXAynEuayxRfdgcGLjWb+tnUbHtGXtjRrLNlIquj8AtOMnEUbkCYLpJ2tpuwV4
aY0SYEVTy0i/rQyK06kI1FYyyushWHGuG1PIEJJhx00Vv9KZyFMNmJOpCLjgGtXC3NOX3Lo/6K31
mi2aCmWgJyfpx1ADMkhw62YmZxQFoF182Bi/WaJw2Z9e+NE/s17HGGCIaGJAzbSFVcrRLCDbRZmc
ve+xaPk4n7WgyF+TeYpmDnsqfEo+Fu4UZMLL4aAZIadajmljvO8PmnQHL/Z5ScmEPkp1qxBkB7+9
VZJ1O5XFeWC+62i1V1eWpsZIKQKneltQRf4By4r9Mkp1UEpdKbAaOcU9S7YKGnl9PnpzOHKdn6nF
wtVjYEhuCgDzny16+tE+pvTAoxZmLbcECA8spttD4TS3lDnjj8inXS5NZWQb7PurzM+SW7Hjx4fV
aOvIok1KE/qXrw3inJsdH7haPPmGhPNW/dwqDHwKn2G6aXXCMYKZaKrjMu/xHMp6l+Z2JZmNcDWQ
Qgrt/N8/dwCzgpyx7VVZ8vV5+CxaoBnHfNwmhhWX2PgelDElzywIRLR+r54/R2Bs2cflRPNIYNQM
oH1dUZQGcHrU/FVxy1zFiA1RhKhiv2g3rsW2mzODVhh+RAnD8pQzvbH+1jytTcQfPCX1y2yoqSEu
Gpk9qJ09aOp8sh9/xJ64zILWJmvHoPINyw8J5zCnOD932mXybdho06mP129KMZQXqg6fQFxTN3Wq
LArtCZIEp7zh2mfpgx2mZsm66VQ0f90WY1cTztY3T5vhz23LqR6wVSfrplMhD9ijLFw2n/molhVw
tgwLUgg1lGRAZD+NYl1FyvETGtS3HHz2DVtEOES85gZ4PCL7C0TsdsjIpB/9w3nExDNm5rkYVviY
R7HZxXsie1MVAjKscXYMrgMjTok3rwJbQqLp+C2ib/MzW9IDUABe6xIb4BFO6ReP7eTpQr+cpvQR
0KKOQzWTt4O3N+BO6gYbo8xhMsdkQHMg91Cic5olN+5SZGm0kLiyJNtzGzr5hl/Y2KRlOP1f6avf
qt2pkPNxjpd1Kxjxqmv5cvORgDnrHWrcvb9hZImJ/yUz6rSX8f6SV/OPZS3EqIBHClNouzi+F3cj
rw1xZSZULvRgz/X/ompWM78t20gOstrkiG9IMXUPCp/ECuEz7Dxb76/HU6oC0yTa6gBZDeWV/YLA
ks4GBFDysp0pVUf+y/Ynno7rOzQHEyjkYKwGE6oQtsyPobhzjaGrwhO8ZJRUESWKZlyijEuT3l8O
v7owosVSGOHki+sz59dG+aRMGnsYSXsRt91FKLvRsDNEoqbTzVtbR7PBrxOpbLBseX14tFdUWvt1
i33oHWkdK269fdM2Gqp9hQiMUvCpY0yclgdf/AunbymtO70zQO+MhO0SynAtSmyiDl6dfRt4j8Sp
qmqGMhXDIlaaiYTkPnR5QniSgXEieaRetMuIAQFEHZtH96/XpmYSDbf9Z3kCRrGj/XORaR4q7j6y
9zTiQ2YwqJRSHU37hmLrI2/SV9wOwFApRENdu2MOizGhYmWxHTFBfb+qhgAi0o+bbCwWy/77MSzl
vgMqkI8SIjbX2ycwzw48phFp+dzCjH1uAFpzr1fReq1NBz4DJrzfIAXHHvqaMfVzhvblaC23BJ/E
7lwz2xsPi13Pl4UOkCzslqIeGOjSWhEurYQojJK7+BXYAHRPCyHSLe6cW45k50FBh4d3EkoDMN4t
NMWVEweishOo+QDOzjhbKys/chFYYtIdpnZY1R7J2vV4wAVLGWU/Gc3xoPaZ7BL5ic/AuU42rEu+
5/u7VlH+DcCt9xbhiEgsgsipdxzPrUAG2yiIdZtrdvy9Sw3ee3logQYL/byPtcqS48HtPeGMEYey
THAkmSDogy9Fokz0qRQW6vZ4Rrwy6Ru9NC8Bou0+Bb9AON4lStlM1onZZyrB0H3+9lZrId2zMoMh
MLWxjgxGtOP7iTanZp60OAbSxn+NemlbSUR96F1RbLeZhxnbJ3+cCkg8gl0bb+YLcFU8v8OHp0m5
wyM8R+tVcDtNtySFWms1xNZGswBxOs2roD7xPgsT6JQgoHdVZWOx7swSbcyW8fm0ksmlVVIHs2MG
JnaS+wVTiBWDspcc4F+lVjz7M8E+OSoAvYeh+GmKyqGMfbRYA4Th0zbT8WjVy8+aNqEr9gITMv14
SgkPPsYlTuKYW3IeYgvcgcxbqfuqBIkgXjLXj7xCZFEi9Bt+7fRmoJBWBYmhO0l8PfqBvkfF9WzN
OdnvlNlahGg/rGiK/GCjsr1Z/0AHvTOeorsZZbeh0WeFq3IFKL4l6lcqxzljB52qbLj99BVuLHvF
spVmCXEqT1cv7gf00uqAofWoJfhiAVbGFlSgypl4C8JX+UlQGjo6dOWd03VYPfvw+TpXrRbURT+a
80OOtUVVPuAknvuAaswqEevpUjHIegDljDO1nfrZuv/1JqdkH3G4j6ORE25wt04oHHypBMbDT8OQ
RgblhlWBJsAE3mU5jLB+j0FXrGQgn+eDN5D1/fxp9kgsRRn4jC7rFS+um5N9CePnDA1VFlCDvbAb
KL5jWbZVb4vFeDTzZF1ox1Cwy3hRjkB/FQDzjCSBcmS3X64tZJCxZFJlnKNLQHPDxQ2e+STbZRkD
xq/0LpxR+ACFjvJWZUb1ds5di6lZkjAyZvzy0qmhWBGSA0AcksGi9fzUY52OEbIP6f04odZqRUek
FM+LJT5Q43xJ9uxXuqtJ7LqEENcxisjG1A9pD9hQv70VhCugfjF3756et1H5ntahXh+jhI8vpUIv
crHTVogAljKjbMQDW8jKjm0HXlPSF2dbC/p+rThdyLJr3H4DkUVCXUZ8mvcq3PVwoG8tgS4b53kt
6BP+0vlwrNn+h0HDW35tFPhctcuC4M9Gow2m5u9Qu+pbktg3lczneAPxqrO0/YyaHi+UMg/X0t3i
KdSpc1qOwPb0wuPJWrt8rRd91Zk3fVIvwFc2WJyuCvzKvONs+jvhBSHtEiZC+PZhAWuTLEnGBuWX
xQU2LVzphS/0Mnov/Lhe8vxXEsJAi+dWd6SNo08PvMQJ+8n0yhflBqs3ZjN+cajJJ62leBJ/WtJC
wVfZmPTPC8wc9laMbUjeTz8wQDM1Q7ZVVYcov0y/BIG/y3f5eaJsLBuwTZIHF75ssMZvdz4UIIAI
V3G2pmOeywq4JsvIwfB0Wrz0KZ6iG7QozNnLwl0E1W1ou1RyHatEajyQv9cMX2IKay4WwyQO5kDJ
3n4ZPpKHHFpFFdMqlObujwRq1hbLR4wpET+GlcRuOXuWc2gpW5eS+n4K1UgYwP2PbUcCsXc+CJMe
eW0mJaf4Bo/FO7Uo1N6dkcI4ZRLtq1Oyiv2HnJ11ub/xQC5A2XuHzUlJ+MViiNEkJQGdLvK+cCun
s2PeAqkMhWbKQ27wmURdxCuuZ1ZLEijJ7ubhr8JiXbV4YuekKzgihxnsEZUWN6tIGhmm0kL7P9lN
DGcq9VUQE3joqtio0s/JxncbpOWsoMk0O88cNVCsZHmf24iuaoLmHF8LsVabtYQsPYb/te6di8nk
9HT6xR1HcJa/FNI/sSGkMV0xV6bm4Blm/59Fm6ebiCsgb37Gy08mQPaUH1UuGf3MdbjWIpagjWnv
lI3EnhwZl78QAspf884CihLSlKaNufzMJ1RMKW4r4neJfbgCXMwp7d9gKKKZS4aXZB9S9ZJtKhME
XuUhBVxBhVI+oFOKKZYVus8Q/v1Z9UTS9S7ES5RGzIvykqceFkl04RlSNyYLygmOOK69eXO2+Ies
LmND3ztB5UMRtmvYBJRBw/VtFpw13UGDHw+E0LgFYh37IQqi3qQRVCKZNz2fza/if2h7OYleGQo0
AenXCiNp3Y4SSm/ycHEuOp/L9WjsqtyF898DmCzJHbWIUMgMDbCkSQsRBF+0Ykuc83t2L/ZhbM7y
/TzBt+A82/B5fU8M9HRpQKD3hCLe6YHU6jlwrcg2Uf14i6aNOjnHhng9AXIXR1t8uQA8JCvCv2L/
q25E3vxMAhmzaDaU2VHR0H9Kwhz1FVKQOY4wrmarE0s4f+3kr59WSxocgJD8swCN50DkEVT0kbCb
M8hutiboVJ4rp4NrHiSRGGTtN8dxlcxBLwXrjY0FEcz2rqJnY6B5ambjPEII9UyUPfKSjE6+c600
yDZPpSj3wgAL2cvjROAazlwfNOrnUyoHU6Q1d2UBioEzHQpA/igBXKQt2qc1iPu6JByI6qNTDjjS
G47QOiCf3KadCzOmJZ9V0ay91jY8v5qh9LLHAsjInBgMho8LgEEjrV65tFwvM5CFOLd8TpdsB95o
6rL/Vjxj9ERjXv0g6QHc9bdsQGszp7aywkZgU133rkZafi2PHjnzT+zYZQ3suDok6S2hLwYg0Uy7
b2y0dAPB6bJv1Rx1hr1ygrnpMAu877C+rIVNz+LAFW7RMtUgvkRIxGakZx4xy5Yo/dNsarfTtM6G
9MmXW7IRWBG64N1QeBkRy+w8DYW1Y0aRXWUrJj0Q1/m2VESuov9NKE/nhIZ6ZjkfeQy1guRsOxtR
fcf/lIJTjTTHmy7a2d3dffQfT8/uv9jVhUb1I+vVjDyXblKJI9min2njP0d0zw/8J+dalPEI9KuZ
ga+gD4Ts/k6T2V3RKWR+ggDww/MjgPmMj9NyAunX+6JuaY4lNXyguEJlTYSbYqoSv1lXfsqH2VmV
G2yq7lUazKZn8IN8zPo5yZIWbfolITVAAxaYJEiZYWddgfTDG98WaoO98HqjK/f4DGW3rZr8B+WE
lO1yxhEV8kZ9hqomLMIkbex3PNpE3bXAVJ1NMc+6IbBl7g3o2tghhvXIi8sJGDF9zqL/vhk4BPVo
LOOF+6rDJc+0pzmZsjTESxZZOgOcGRAPXl66TC8rzVHsDJ5+ZTMKgSNSAEiYnU9Yc7PUSd8uKufM
rHOljhrE8p8yRd2eMWyHIMBUjNiABjbH9V9QAzgao1Zixd+lTH8LPS7r6qvtl1ch7rnHxQPn4jqI
DEN3YTCTOm5nJYWTLku/DSmB6pTCRIGKPUfV3dpAkmTLO4glblgQQM55FY8OXqleBmPEXSXtbm4Y
BLYq6VWpUH5dMucClq+ukDNMitrj0U17ghXAsyFaGceP4phtEaAr/2tR+eZOY9ycA0/I8g+9wc8Q
Gu2z3CptTtyK3U+PHtpJC1AoabimmqNjdK3CMSRlVZPXNW87VbZ+kp4XxVBNt8dfiPu/gWjHZ/AV
YsFujXPX+VpU5d2DD5vHUfBI8L1ar1DrKcfJAA+SFYp4pAs20dxvOFJISP8s40Vxyg2NPtNLXQ0U
dlLvuHq0AuhWzfajgEesIXfHag0gKzvhDx1DJpHpkv4uaPZs7j+n1g3KGYebb6RfDNxP4OTQhygJ
CsihDZioY+8t8gK3uw3yoFYOI9F2av6VEhuYjC/W7Aa8cRCxvC526udPhHc7EFLQ/lr1KW8rKYZl
mpJWiG4Q6suExPi/+ACCR95Wro6Y+aRz8u+3K8zR+l9oKT98nSZ43jGQd3MffRVSvLG0SpYx+QuB
h8GZgGl6i0CvwgX0YdNduQKy9NaLGZZr8lK1coEm3Dp76zv8XurZG0J+Z05Pu+ZQs5cywu584QvJ
MM14GwJRGKltUGaToDPCME91oygDkU7fXj4PsYZt+/o2JoW+xFlrd4FH0I+bcg68wKZRClbevMfH
UXBHD8qFU/O+TUV3LvpOHUAJzZRH7QKGNAdwHdT8eLYOQJsgC4JjZ8WRT2RdLKarQL/dErMheVdC
E0Y+6ZucX8xOoMAyvusMc65BEkEFF/VEuQ/0wLvXESxIWcDWeOS3JIdt5GQ4oEIwnVIuDvam/hu1
2KsjRY8zjQNO22c49qJhQ8fcIwOhV7bAYy5K2AGMxDz7x51L2JsEsuwvXujeQdX4UwgnZCKd0CFu
9WJWO16qKTbWblLjjq9nsIvC5vTYLyqaCQBRnPdmTDgrcKFUHc9x+UFh/81/iM1R7SFxnm+6ueTs
EePIjSOjV6d12hBnNxRLNj4e0z7gBsTliPFK0uOrYEFt/6WtnmDdMeV1oMhLsJ6MXG79GGpguRbY
C6s/ImwiOaTFuQ9W4Z+wenu81kkFlv4r7EdA4f/BkHcUxQmKaHlJArpix9GnypdFTP5m1hRfAWt3
Qy6B6mHX81PBDb3MFg+ddZ0XOmtsxwbGx4GFoAu5ACjJ1qgjMHwwRW1e/uqlHFc6SDpHU6668vAf
V2yC0FsDQvDvgs5W29w8hXYrjk2DVPH0jIx8IbDb9fAdByxxfpWLih0L0xf83hOpOoL489zBKwHu
s9Opf5XCWnJa9J/WQep0NcVzCy5lcmXMx6eMuy5+h9/AL1ZYC72Bm+ODIc3+sa6cpvtxPmcLYNlH
8xdJuEsEH1g2xzpYCklgpXumcAuArm26lQhug5GL8ab2iXYVpij6ONBbuXVcYhRhyZwwAY4df70d
OhOc9KFTgQPHmrjmlfLNGhERnOUP7H0RaRNaemY3F6JKN/bIiUuFXZ3jKof/+hx95PUa0x4JvMyL
188ZDInkvHb/rL4ZzFQEhIvtadp9AteC7R7JNo6C7qB485raSFEaLWRmkG1TBTuBCvxdZruJ34mv
n4o7rXn4OrvW/uTK6xouKO5m8OBUPbmOF1c/gmVEpexQUpoP4CPvXmkKH4aTommQkRXPhwn9ojq/
JTmamT5taOrw7ZDtKHwV6u5gxWUfFYzWaXUGEFmtaUvv7cSdXOaDUB0TVlxYCi0QJK7ZssNta0ME
lM+M6mxTNzzjRDkWpZOP9HsqClTAAFC4H3vAgW+Nk9ai9hpv6PlLYeNSz7bVnh60tPEZzZ34G8wX
E1UJPuVhTEdoT32+VU4A1Ba+LHYWwg6spLYS77o8uxSWJC4qysP1yRB5sSbKqEop9I2FXKDSYAzz
NKK+kb+1eC0y71Ewbiezz5Y7TrNuzsPfbEH0MSmwJ7n/dCecihU7FUonGs7SPUhasl/FfQRz2+/h
ckPPIJMoSM2QubRkCpZSU7tnYfQX+vjuLCR2cvoez3xBKHQDfj2ueytvOc51adfgMhd+nYVy3ieH
TNwRk88kc6QAsT1vpPrhkfsmO3lvB3Dl7r3CfNriWQ5l+44yMLZS7iDrc6aHq4ZAnX2oEfBerUJR
dgI8gxx+BHah3ftxyMsob2rtRlRXcLeHBdRHuX7QMB2yu6Vz7oiJMxiozFfwf/CytIUsOBlvdvPM
xdaO4KaaLbGiGIAqxxLsrwvzyChZlQxmEtW8iIdmXxKScTkNPKhsgPgCCY8AUTvyKvgKy/LWnveE
GclT0wpnMSkblcj1wTaXKZPIVE31hUfQRLKsScXl7zjnkuqWasudGNrOHKb8PPt0PFixMeNJ8QmK
LDtQ48SlwqeU0u3oL2m9BFE2/sWnLhSpdeRhzwXu7mMgxsuYpjmogZtvKFogZeLnWDRzsWmF9u3G
ekiWsTlroIyLk9jpnIu0uwOcIrUUe2I5HQRNxXulT704HRyVnBnDfGNgZwzyQiMAlOuqfcIaFY61
SjL2tl+SP+PKQTBjtddRG9l7TYk3SHqaLqLhVA4JXMajMTqZgMmJrFr9YNmu1KuXtu66CQujpTBi
PuXXNmb/YHVi5f4LsFwIuV33svhkzhrVJjKtG6SOoJfpJXco1deJCNReQjxtIxGEvh0ubIEek9Dq
7Djtx8TLtrvXG5m7dAlCTlso9sckJii6afXXpWLIkNS6tVB/5jlOccJue4X3sx+gwquVnmjPzZhc
bqbRCdTJFI8iVN/EKLM1ETfAeujzVGN7DKEYrTSgI6oIiFMCnhvhGF+VV+AIpNEAs6RIlvrMVSud
WqCLPUQJElqGzmULcMKQQdD+Pcv3nmOTLSFcQMmYc5Xem+IVpTgKFzWJ37pJDpjjDApq/6AwfY1X
RFkvOD1ez/eT69N8OH8rE0pAs8B1YrC5z0CSv5M/DgPlYVcy14WYpqM4UyWF71Yap/0YPQxQ33xL
sG3h+pEoBhJpeDRhwGiKsKHWuuAxQD60eHFvexLqxU6X+caynCxU5NjL54sM7OqASIz+wZUx3xqz
36fxcXYTiQ4cgpeRUL5GkHfGejHPMptAE3xKCZuB4/JYKJAQoa7QSzeZBQpOBDeJTjMDB5d6Uk/m
tND4vqcv3zLWTzgjj/bEXnhQBGHoJ73lSUAn9IHz7tytKGLaQjrMuAnW1z8Qef23ymqhUWZtGzWm
YCcFahwf4ILNx+5f1TGl8b2x86ILD7YfGY/fy4GGwPwU99zwsJfdae0eFDE4jJ/J/DaNQTPwLr//
pfj4eHrl4cwv0yCFLQeRE0Z6HF56uXAk7sqBQTXntJQeNdLh0Pav/XOHuz/FD2k4YR1hjsxN08VU
bWZm7g1DuQpb1fkVK+HuLlL65IxdI86PUllcvi/kJ4ivhWS80sCAdYYnViH27/N8IZK2CcNrqRPp
8NxsP4f2OSAS+ZSqcdWP1mTJtKuaclg0gbLyqUEPV1UeuimJ1Twq2Q0a+voGYwtEaQT5kbghw7GB
PvmqYk+VgliJm0dnwzJ8t9YvBpWHwbYb8XSzMCrXcBc/fZx1EDOx5QK8CbDlpea8/rpu/3238BG2
mQDMtjhsrWQNj5/2+QqASGIkl9pyi92RhG1SHG4AvwRdLUq8uwsVsM+X3IVRLw6ZOkIKkeUYPk5f
TSZG0M8Q0YgMm5DAvjo7FiERC62mgc4HCwo0kT+tiS3qkBjWcPbmYgxvoPIixtrj9nQVu/bC9hlb
YnrpcE5aGlY9tnIHgqfnJyV8Hn2ZnbdQSqHvqFinqLcc+3kW0hyBM5y+Bfpx5eQ1RlVmbIjldHzP
48fD0NAm0x39/aJn6TPHJLjV/jV7pTF6IikGPBGpFGJop5trJvA2Lo/66nq2sKccqSBZSDtELIeE
DnjS+SeVJP/N0vafmqtfoGdT87N65tIRjfEwhsa5CsEEAbg8ZFty2Z25Ay9ms6O1jzXKCy/xC7Wv
mToa+XTGmtE+ELmB+qUaKkD3m0zfn2B+a/sOCrZosaOKIt3TWLZqJS/Menq1eg5ZXmDlJ1r3NK2W
s7LAjlvlV+lxTjuYWhZKZ6j83iSDLjkdNZCPmGKy4hU5zlT1NQXxL3dSqDHpON9KYVnGYBuyY3S7
X9UZkwkiBZA5HUviShODk4iq6Lxz9BVGHsyw/muDqbcMRK7ejaMvyPwqxsa7DGtNbEFNkAnWdTt9
deouqGzXrmHcfxMyqGTQIR0Mhl6CQ+/JNdnpTYsJULDQQzPy6JmZQ+ATlgMCRk31loo0TrR1qDFu
qL7RF4r9CPuTWK1Ah2uQJzR3+Czu2xiy/EwJAGFlIwr0SG8lnnOh9QTG1JXlGfnfRmVhrOtiA+bD
KhjBq8Y3y9k9aSnF+SJhhgq7KviU2EX998GjheElIDtWpbZBQD7AoORqs5O7VDTJ/JUQWYD9K4Fu
unV/KA3R9HQbcQX0BFGNaORbeYoJZn/8g66b5aGtvWYdz4c/v0ztHcTqTbc8Sh3yXOtJc8XgFSgm
xdoUbmfPpvPmhxkpsK2ydER08TOVXeiz2R6hTA+PYHXokDkybfXw0wddgm+l/qGw6bpmCj0C9ZRu
iT0UWZek/rhByFCFfghWzzYkOAmC/I/fkz2tuETYo8SVPwOEGfA62u+7+ZDkLpZ5v8k+vfos1OTx
DsRluOOZqQjGAilFGhcep7DyYD56kG2F3itYJYA23LN/l4fdOf1OXV9y/YZIFmgFLjdpVRLVzQvj
O0tTzGHxA/Ermaqoky6PJ/AzBudxaLJwN48wf6pEEEjRFwa48ivFkQ3+zuQ2uUUik1yvmz5Ud+Yd
+UXKF7XmUjKbfuWPT8HRP8UUw4pfoHkOGSsQp7P4AnBTFgcvPuXKoFkJu57PUAP6i2aINpGvSdQL
uy+AE3pg/kRh/epUc2WFpcx1Lg1QXHTGFCLivONaSUm+Uo7ErKLHec03LaD3KJ/Gm8mkeiUrBQbA
QQ53KXaN9ax/sgewt4tdGIZCBFyKEvyCq0eGLBSDA9rBMevd7KUsJAiwgpDHI68C+Zho7EdNQ304
fQmt3Nw8OzuzIp6sPDfv8vF8+eY1YL0OAcTfjhduOKUBnCeMfTMbOSO3zT+XbqbL/3zqJiRut3kW
DRCxZZvn9clEtN1lW38T6bw/6xqHCBZGiLXkZ+LCoGOw1ZbZxX7rTp7DMdnm0R092WKczC7Pj0fO
6iX614O/KWR4hVldZw29zPdKdkDFXaOVI3Vf5jK1dbE/G4nRhnd/f3RtQqLCyoFokIAnbhtEIDV3
xtQ9412AYRCfLh48ZN3geFo44o+txSIAuEDWjpPranZNGGfO+zgPal7o0s4tb93R1BMofPJSnUdT
tp/M1UfimGhgG/Puye5UqeNT3MZgzAtfuiwwnAtYWqvAMLzx7npEiifZV0xJRFA6TVtJsOXOhvs5
y8TQdOSdLMf5FqmNa7KhMBNcrauOQH2KTIA+qm2nyVkSJI4U5vyIbyGu9DwaDhuFzVucDPQpzlZP
6BO/OhawQ5aPYLcXx4A2lZrUQAtURQINljfOezLKpgWAh7yF1VEfP/umkTUHlnire3u1uCCWFoRl
1V/MYPDCGx6z5jnx0e5Hof2yrEq6WKvhYcINtiFny3s51KovdRoto2ZhiHgAx2Ny0R47TkBIFr9g
N8TWN1TPj14I/lN/LngzLbfRUjSZVSeIAeXy2af9J1mpaA8sdYSyCYkU/hiPmZ4o6ovPUL4YrIr/
LeJMSZv334sKxmThYpWNyFPVTl/KufOlIlzlycvSLHLeJli5J/491p55SrrgOFu1veA0ZbF6bAYA
5TdWI3INe+/+71Qc0Ym1bkSEZPvanjDCVHulZjabx/PzF4lLEr5M3LhLtpH6/U6pSRY5S1lDLUjE
8oabWasspWm4e6hEtiKZ+Kw7vuWYYMEeFDcNfzW74Ih5oWiql2G8F8/vzVyULA8RXpbu0+v0UuY1
QxP/VDIg/RGlSpfgExuuraHrCwa+aXlQA0Qt81othdDtMEq3HsxdWn5WlMt8Z2228jDNWBltpZbd
JyifYm24ZiqmNdnPfDzOPdgUEPdVACLZWCyrJus6WIJIY0G78Zl2NlZkQ3OPPtNVHkwN0oP3LiHh
zxlu6ZEYapkIY31367UvvusZuZfosUJzhAhMlszRBbUQ9JrBWmFuWV3dlU6Pi0o5CzDDxfElDSK+
70kufx1dZnODgFXNyqs1GBNkKEg/Lgvcbfws+1nzG/pIsc8xtX6kqKzWyJP3u0MDtFtDBRthKG1T
c1kzLG14A/uxZAdzUtBNzQJimLXac5LTqUH3Mz+y0dOrwHNz+X1wMLLSdFFJZ7oFj4RV8rVCwXEy
NnO1cHCR1hTLlGmPHZtP/CDfdvyUp4JIYyUZTCZXt2zT3G7uajQskYIWU7xKvyWpslVEs2Sx5NPd
L2RnkCrp3WHT7Ie6DnL+1GbwVq6bH4AM9uAzoUdbJ2MeR7bRAVAi8KyNkf1rLHfj8Fy6BHA14Az1
uzSdZsynpyGxciS41yQVatMkL+S5/Js1V9BvMoXnjQ83M+7IwFuM5E2+CGdbur4I0iW+PYU69di+
nTpZnb3t2q+4CTJgKCPubLl6f87IHI4z/2zKu6gO92FaC2rBD4hAeS33KJom8MAX7tHgrdSpPFnS
XqSuzgJ7XKY/m0gZRe2QYuaqYQamvU1Z6xIToPsUfcUTFiVwl7Xay+4SdRoauGZDme3TTVHTjNx2
QuHCSi7VEfcz4/3zCsmbs9PbxlJEDpJ6QP5aLK6cW/nimImyFtjwhwx77e9Xk32NjcfU24rWlWS3
RytHiUz3+Cku2gtiqPixK2rglstC6M1kzzgcjk49SQySKRZFX6AIcdwVFQA1SzfEwbJj507Ah8ZX
HDzDnOKehax6hOjAu1u5o5BqIrz1lUVdESB7UEmM1IvC0YsxtCrYRYBzHik7iC3xRh/g8iVv4rGj
3nbT0xvZi7BXoM5MBt+kzQ6mESKCp1fpUc5O0+dORzBaKR7kLu+fTLwkM/5GEfbiU9rQW6RatyCL
y/eEm+eyIDyvi2a9FP25kuXxYzdvrKRVx8OnUHXHQpQu6uVMAA0UQ1wJWLnCVM66zkJhG/yfnx2C
obuROn2IbnDZ0pHmdbOchr/mvN1prhb2tAyaN/A2dbJXEjZ/JKxJxIrpKwB3ZNZjaR0uwVNl7tTz
idmqbLb6VhtLPU43aRfouryK6NHlEb0gkI1dp9OKGmXnzjj3RY1Gl4HAiLv1Us3g1sYdqntf/qVU
GOT2fcjn644OWR0UPpRFCNUJ6wXozIcHdxFPZ+krTsyBoIwL//xXIYjEWL8WPELlZJOfou8nH0YQ
0IM9R7ElwUH7NovEH5amVn+sNlQpCxylG6xWzb//cO+BP78srQvSLw5p1CU/qe7Ac2c4H/Tipsjz
MUF//vkejkBDAMoghZfe5IaPP7pt+HAydEqoeaGETALtyl0akEfq1cN5yixCN9apFYNdD2BP9Gtn
YxkzgM+CH3uib7fk4ux19iWDzY6ANR/0j9Gg1VYX82aerjGXUV6nMSvNwJy7xjDEqXYkZWEN5l2v
1BCDn/Wu4APQhCBvfnm9IEavzbslBrGb4afc7/hpszDSFCkpyFzuqa0DME6saLPUIPx1vAvrYMu3
sX27268NRNynp0Zwog38uG/KHDGnY84ANaRI02NAqRsHmVH6Tyv3gPwfk2/0GpFftjgTxpoChE0n
/POzGQlhgbn9T6dl8girDf1ZnJjaIg/F7fRtMfByYxx6m+gp9zX+JBE5B7bZj1h3G/QwxYLoPprk
ZT66jm7VL733A4ykF3NssDbCQZ3c/5BvlkiDuBWolGJU9WGrJmlG/WoRaQXp0B6b8v6xKYo93Vv2
O2ZCwo+6hCDy2FIRhfkUcVPMUNUEwzTCp+Yylu4Iqbvw/XANAq2HCfqjTtkfRI41m3DIDMGww0sr
OmUK+ZepXcg7yMOZHhy/+HgVE/DPcgcGcYauccohDLU9cmUEj2Eo5VKzGLedE3n/T12U6ko4P5n7
DJfEOJqDuUaAT5zK8H9tnuujnY/NA2RtSE59YrlodPuKaG4FH/TBANIpQge509TZ9Uke8EoQfxgq
gReNT4rjSyVYPx6o4hoD4nHOM3zwUdyI7aGZiTlwojA0HTgRrLh0NHUtMWTBTPPU1l+xuww3doQR
QaejGZACR1SBhxh1ScVlEeZ1TPgaCPdGz6OjvxHUQLgyF1OHTRs29/38R9ezx9Wsjk8JaDtogTOg
GSlJBYcj81q1Gafcad5PNEWpv24F+RXXXk76Hx6NvEZ2tBquL9fDlNF0z1VvZJVoSf1ZyEc1EBq4
Gu+XAZLxPFa+Z79ske+WM9oPIOW3PleEWmtiS1AEyBK+h81I3viDo/6frfsjllhcx7zVP1fev9pB
DP+ugLwJSLcEikH1FPyU+BSDCuGPosWdzt1KEmzXqSChyCMWvmfNBTFr7H4xQmO1s8piH4gekqku
SeDRadNE9ylxZOQ1hyQTIrUrx1EnHdsm2RLqdruVepug/ZS9BwuT+4Y0NCti5kyaWhJsVJkifu3I
eogxC0i5xXIqDNpJtVdaqi5U8NBx3/Ww4rMnP2yq4Ewx/KeCKiHEXzPmNPl/GVgapg4ZYleN2ysT
rLis3TI6oxa2uz+b4AYM9VRVlTp0/Eya1lNE3QV53seLBRt3gFJj0GCTzfw5NnbovrqroBn41Zqy
Vmafh661An5zML6IFbkKhQVrjrGcOdui3fHRwqZe3NPOz91yiad0xBHtUrHWPSb+kUE4o5wYXyQm
VqaOQgdnV3pX4qqvoCza3vLVqqY9UzlOY1b34a8VLbfh9+IuPMmXXWprwByZv7YanEjsypDGo8e1
jpIriJEL+qbr97dBzXsMYHntL0xe884M57REGLcchlTFQBADDUpFaaqwOvo0JaQxp9GdJzsAeMVi
O02SvCcNo24RfSUnkujYkvR0epZpV7RtS+/6rGtFCRXc6lBv16x/kV8bmby9bUSD92hkyd1Is0A0
/K3KRbhEEsvcCW+ZG6H+OgmzsnzDI/w7cGVubaXWsFo8TOnr5uvuVajNKfWM3LZKjdr+bhAA558O
cUiXExPuG5Oc8CqVi1o48zp+TClcDxQJORXthbS/IWdAZkoE4Bs+JvyD1BV2Zi9pfwDu2Tw3VnSZ
usq2MVOneIe1WMCI5JuyVV2OPRRCGRijoEiMUnAJ4UXt5KuNct8XkNckleUHYK7t6OOdT/KbsW1r
bujdFOURPCkYgo0vkFkdUmGutIjr2pLhkMpVkLKnEpLRMwz1TN8mJYpxgi33PKQsuO/TaXpGB2Oa
iHjoP3Ex7JOqvbeTUfQqir7Z+h0CozDzkLg60/81So/RX2380/hNQf2FuDnGsLFPppxRuB1QKUBn
1f+RCa+Cf+S3yjU8AOv4Grm0I5HVe/o0UvSPsKksuSLtEhqOCsB4vpcknikHrXa9UPy16oOQiCTC
ndMPvuKUntsln8CEWUKETh0JhZXavf3WqdW57BeN4FOSRgYSFhXgjdRp2Jhac8DusI3tVbyC/Ryj
U/E/567e2l3wznUnZDXrTKMzr0A0u9xCfscYuI34/W03OHj8EucxR3jIIV1E9HYfArKUEckXZYBb
jZzXuQdZ9DcuqsPAHbOtvU3stmkI5ISGu9R/P4VkV8Vfp+s4tMzIx1HcPigjnVCdPxc5s5KFf7CM
brMG9We+bOacpdWcKkAPQ6ZiIWrzaR9ViRLW/uT+wEHfIiFlRrra2Ox54LJeE5TVxINOkmA0W+Wb
YO3NaqhAP4PM6WjRr36lmbREo5UvuYqLiqG9bfmDQRaxwFRgnnHi/yGN67TjwDYEKapBperYCWSF
7lQx19bjNhDxece8RntkavOBdDSilpV4dcTKAxJQcRC/u68HdFM/LUG+Pd+TohO1qcZZFBn7Hsfo
uFsuvsjbODYe9+G76BE7gNUZ4F3HK09334Bn+6eSn2apG0Ultofi1TkMyEI2g+W410MxZeLoDvPA
Ujda3yU/F9HjDJ3xQgJcGgixjDmNa1+54LlSybAs2ZZN0INceVLJZdYiWhQS8opXFFCyFYUj+NyC
urSz//D78DyUQnEXaMAO9hvae+3NIxnAP1cU579ZT5d28j9Xbn721/ByHjgBySdrI5IIlQyj3zFy
iCdIMtlidlwG1x5uDzouPWsfNcXGhxI2eNRlbFqLhiNw4+rmQcnwD6oNUSSmfqFWPmAO3SqkwU3O
Du6S66Ko9bbQJt/oNSXGOpMsY0gfgWGT3iEfYzPzYYYaSX95mvXrLHBAn0OBVt30cy+k9NBtIkoi
otjXQCPZKkzoFs7LLWXqzKbQEuLSbRZAiN3cBSqB2Eij0OCXL/sR/Yf0AM+WkXPh/D69FErs/TR5
UcwFEMbhkTh795261CQfZhCFJUh/YkPMLvKnnN5bOM6v0VS7nglbefKv4hVgZ4hvqEtHHjWhLK12
FETb0gpx/xqds1wIOCGnrDQ3PWSKSsHzzuOzeftjss50U71SZUifPLinN6alZaB1A5LCuB5Q0aNN
paGOl5Zx6EYIu8QVX0pTSL5SdeHru9JV/ay+2VXtuexdgeWEW7zsfNWO3/IPSTIWGuYyTvxDsIUg
qbCSUolP16HIgfVa9c8kwNfeM+uHzaHT/aOpQ94bEHVnB8jKumHbGQ2aDo0mj1kfKlNntRUBkY4k
EJ80k/GYfhpTNVbCV8DY9pt2z/B0sJCdE3dH5PnZKBHdVjvs5hFLlZB17fxRcyVbnbv5Qqj0CZZf
bFzlTokvk+QDUOzCwTmUsQVoyUUx3pVC0O/P6g96dK3jujOA2A4EWtt4YGQFI7R24EETd5Lcf9eU
CPC3dbqpgafmLced3PyXqb83z+8tiVc6W81gm+gyV+/V3F+kzkc+YwUvfwxgEpWWskMV8VbrPyKG
4ReZwqRD42UNQFV4bgGJ0wMnVBw01K6xa6ThS/5YCx8w/TzSYk9jYR6ZYhW2w+He/DqAJvY+eu0X
QVg1X44O4qRjJI/JC/3BsfHT8A0AmsZZM8FTRu28J0VwtmXpMkcDpnq+sUsO5qiT//sPsOAIr3o9
nMuSIuU7RLKeDR7mktGunoFMp5vz6ApCz/fAE/8jx74XHT/EQ9zt7+3CIgH7VgnjMmnJQtK/yk05
2LSD2S40q4WbqLIMh0Eipo6vDutBjF/3MxUy4raWWzAYlRMo+7ZHhj54pEJTVirSAttcnvju8e+F
P0oPf8ZihYf7GFuevinDKAI/Sr+RNc4rVYv9PhKfPLab6dyJh1gToJn6ZHSsA0y756aO4JrrtS/X
j683aHKk+j1jgNa8XWY8DIj9T36Mlt0LLqH3HZ54ExJwD4x3NwhpEsvEO9t+B/P3WesIBlBUw8/7
opmls4VSJwkWtdtrKgCWh1jliNUc8pPypfK6FfvDTDJ7GOWiDoUitqKHJ5WDRjYCyhZhxqHHQc4Y
xxBJ9trV6Bhxg0YZ9Mbby5jB9FRIWxXoIM5t22rli9GeYr2JiigyaLNf0GdZBpPi2r25yKZX5XgX
bPPhwNgUVsc02X3/JBkImcv7wQdXCN1hWu/QILJnhLHdiqcHlZVGb6SOcEZD3TN2xgPR5UN66sKq
5h1r/TPcve1ukaMMNBw7sys+BTZKboKo7HyY3ta6t92uJhZ5z5SAjAC1pOfF/pK11+wjiRvYbX4H
pEy7JqMZjzF08PECGIpSNg4vaHDeRGNuZrs4iJBuK2+2nwqjJ46O5vQJHdthWVHXNX561ZH48aAc
tWQWuW2UatYPYnDj+rolK7Y/BHo63dODsi/HoCaEna8F9gT+zgSuSxlPaMzxPaVIyv3UP7mKMazz
EX0DSJpG4TUzVDpzzkK6uNCAGf376SdJpsb7Hm4vXHHncgQWmCcLtQ4eeSSht61BnWZlHlh4W1B7
3D3ncy5643dU07h2xsI2r7DyKKyEs82gB3c3AGsrfGKCTfuHxKBaBywyvxhduz3EZ3WRkbmAsTWd
SUjwYFrPMj3KtQEUmUGszsy9KItHN9jZiGGxClJk7aLpmC3QbAO5Bp17f5WFn77KSP1bwUp7uNan
xFOw8uBy3l4DsEx2Lk+je3t3wruLSECuN+z/b7xllJ6pRr2XX97dCJqgv5Ut1wuyk1h36zyBktVD
FFrDe6VB49265+unEek3wfvvVfaX1qrhHWUCjULO1gJQTDM6rKeoM2pkIuWq65RVvTgVDELp0ZsG
5h9KpEmUt2gYIH7m0lo4k9VyYBc+fp8+gxRmft54Yy9nzXhleeXon+XO3pEsMrRodwrO17V7CIpt
OsV7cJcXfsXr92ez5zlGZlFjJGuWH3rP+qyAWmQPz7EM5d0EYO4O7ACgGRDUasuWVoLuKM8ectLo
u8ZURD4y9TlTDDY0awhZ8mlZQufxEZa8qpogvpGgMZpGKRXDGbMWCEMe7B3o5Fh0Ncl9Edhy3B56
Xif4YAZTZsnJHkxu5X9cgiA8sfJOCPcgGyxcEAHh/45rl3rOXbGz8iI/pCHuP5zcMbAxreOWcAll
eXBTCOP/OzSOPgrlyphjAs42S8wF8UI8+lhtK6uIZA+wYJHz4Qp2gNHsXUyMv6mFdU1gzbie6Dtg
ysUzU1u2b6rR8DJmHh5hd2erErHtthrQ4H+Rq/mXaAJKFNgF85CmRt7pWNkQ/EmYreZ4+EBPy2UF
ib0V4pUCrRXKZq/CdpcFBkekVcvNaGV1dDTgLO/aZ8dIpa6i9kLqFWLmMG/1qiNzlo1De+X2ixSP
G+LcDrkc2dhhSicNE4fp74xieGuczfzeNE5lShmgmtubSzRDJZfxkvSvpltLnVL5S++t+NVJSdPe
ZPmM6xQr8d7aDkU8Wo8S7/t26X/iYujtrB7G3Otsv+flR2vlTAPR/RE6DJN72fD34Jl5c64y12z0
ATOoslzw8AX8g3XMs/klO57A5oUNtzf7tKAogX+PSiK3smNCOEvdvNJQ6PTfBT4ga2BT2K/LIrtV
s6EzFKMmh506QZCB2L02+sqHecoBRiGImtyzQjQXgDwaDuWGdLKNEkKYAVuWLjErNbD5jH+pIffM
w4GxASc2wQUzb8Ll6C1May3VunZS+vudqSTCf7CZMb2e7bcWRuBVwi5IQZsofOeBbiEcA6CPO6oY
QDWgEDqUaVqXA01eHH0gthhrUc1trIZd+21tB/h3tCo2oJ0Q4V4fddxGtcQi1bFLA+A27wz4Zw6M
1t4LnZFjHOK4/QsqVLOlOrI5r6JaenkZHUSbZwrbU49DemX/Ls/7mYDz9Eo4M+IOiNGR6UWu0NOv
okQeG50MkxVCiIrNSxEEE6ChuiJTQ6ii1dao0Vr5f/HXeuQ7tAoOa1WFCUuwmSBZrxR2i3cu4HXT
iClGWbLIA1xKmOd2L/sdvKvI5JF+hL4mIxHDw9gSmvDrUWwPtX2R5d3p2/hdY0eJUIoc8CSzUxWg
XhnC2KGMCxxu5+8fxZtwEADP+kKfkNCV15npZghQtLs6OCgvX8liWP64EMcYYFfa9/qKz1+1uRum
VZf+bKFDrPHegjmvKFx7QmT+xHlSHRsoHZOjSBLGV5DRXIDU9W4uyHkrUFnQg7i/v1XVO/t8vrxa
+JelMdp02KfhntQ5wr86f+SEWdlJ0JX7IR1mT/4lYkCXHnMP5+QD9b9l3XE/bv6HNirjDcY/yYud
oKYZaDzABKzvfwr7e3BtD3j/F++OxLw8Z4YPm8EhD71l+nKm3Piebceq9cdZVxxAHm7i4M04P3AR
oF2yKmY7WbrKYboDfSVO6863jEond9nl8fJ5gIg1h6YAduSFMVhmKs8U4YR6JUq9u9+Ka1dEsOBs
vJ+3BBem57OLjSzEsMFcTCukV9cQeFRstngu9cjKm0QKTxzUfXMhCuaEyaqx1dXXfrnnJgWqpFRT
5sjclpwVVfoRDBzXwnb2IywflZORnrz9hRhqXsB08H2JqMG2o75Ovx3r2v2xSYlE9oOzhfsnBHrP
LVY5g7A4ViEQO92tfPDdz79kw2alo+LPmhSjLaBcl6foUI5b6Su77KLTxmJjPZ6JS/GJUum0pTDG
O3OsHm/8wxHB4ULY68vp/2nFbgYBXsUavrcMx1Z3W0f75Cw1mw+BWWANEkk4Ugc10k4Spv1eRjR3
rTWTH1/6JvgSTPdv7CWJPUjilxNbWEWTBGEa8aSShy8DL0Opkxj0NGs4fmayDk6/JNKSQ3iT+s56
WAwjxE2IeoFwpABx6K94j+P5P0rEo5prAiykJdwVzH72NlvWiO5VgfUmHw44S7b/d4QzUgq0NG20
ow/18TMXqDjM4KM10D5q7S4nqoAboew9q8a6resTxqMvp6Eqfum/8ucbrk4aJNPAOi8vatgTKw/6
1u8DofGteKjpPH+hNVuoi1Gc+c35lnJsOoFWNLtpRcXuZAi8b3Fpw5WgT5z1e67j4rd0WvWAFkq2
x7IWOP+9v8FFEMyYZltpLUSxIcgcnmN8jtbrtrHSaGx0ShjgyQv2f/ckbiVV0ya0FiuZpKHydzMN
1OS4KsTyyGj2AWNu7S/PT+M7corbqlViIlyW3FM2tXm3okn6e+Ls7OGfQLQ6a6Gj6yR6/fxH2D9o
bWHdbnCAHYwejDvwF+R3mNDK6N80+Wny6pcOa5py+6NiVB+FkSwPJnNpWxjjcF23hQhgT4IwGF9Z
vFeKTpfycGCe2bmwD3/6tzFxMllCgBEjQ1fF59n3exKkjXtMl9YpbCSnNWQoTCDCbyp/Q0UsjHOp
BuXEFU4U3LNYtluzySwIbi13gOrsP5wQ23Fu+O6nMW7Kw7I/LtuQ0AMBPbnOe+Q/JezdJLz0JGME
OZX5IxTEPvY58PRPAQ3k3YOuQdlV5igLTQUNFjN84E4Y78BC5oG8Tmn3oQ9zZLINoke3uxgJAxWd
kM98Vkl5G12RX2W0mRjM4uBJioDRNnjItlMb45YCXn1NoFT7jzBMwWSIVwadk44EfLJR2NPdpjtb
95UCX07/y+3tYCsqtjhUrfYbGairRp8jaF6J9yos/yWJQ7Y2MuegF8WKAYvURLM8pgttWVKkmXOx
Wi/qqEspAVWRjhAZmHXg/DMhEx3mVz0zh7STiXiAuO66887sTWf+LWkyB2yxy+6JZyrbuvOn8SZl
oCzXr+SBLFaxkpWNZ6reyr/6vIAHUsYtMfpaL/5PaJbfWQt48I7cF5CSJ9xjyUvt9s/5zjD4049t
qMpSbis/Xuio2Sa0uAJ56n4/vcDJJIvwmvmtdAeRhBsBEXVVWU4uxQPIYn3EGFLrL8K0SNSo66k8
SBgNpXwcNN3Bri+m8ZmeZkZ/FE9pd46RWrCGmJ0fr4UsxdpFDo+DkyHzurn+EBu+HXL7f2A85C72
s31ChwjnprWeg3oeNKAOUgLJoIsvDo1M+E4EuCSQKu1G13dr4mHnNSfDovhcGqeuelJp8tTaa0n3
95O8vJCNL7pBS6GfN/jymP0URuV4hHrPTCgM8E1OBxmkoSuugB/ZGvO5eLXWkr+MN2ZydwQmn4gO
giIgkrf19p8584Gk3kHW/0kLnnAsigWYZHdfbloO/6BQ4J/oQsTxki7kJgtPjWyOrAtR91iDCuVC
7d03wcgTkkJMIiBIrnLJ3uJ/hs/YPZGz4UGToaF3dFS8kSguKrTp5xjZ4NwtWIgiilhLAGplArS+
oqmADU+Kg3L41AGxUIdrSpxJqU5CeFFlGqJAUDXdppTq7nlaZfSZVNrejsD2poihTkER1S9YTkXB
GxB8tnJJs+mjkCeAaqWKRqKL8LQevAGHqjzjeBk6PGY1PKfNI+qC1XnUYEgfk1b4qhTD5ieTBnjY
zQRDauHa+lxqZgffGZLt6eQn3Zg5kQ/xTneBf+8qC2hiSqzXfFr5b7KAmX1lR8im78g0tsXB1JLY
Yr49D7q803pHPdnIy8Ca1tTsJf571Ei2c+8mQeDMNTaDm+nGNF1vCpr08FHvbllry9u0kZu5Ykuh
hnIQMI6DmHZ/mJ8q5wHZ24pD74gq4zb72WyFKcV4HP5T1BwGUvG5TjU6RjwetGzmKgSs46ja4fou
d1v+uj3KGWWEKdbIpgOlX0lrZ+fuUCewdTgWn0cWnvYRhDNUYRpGsl5n8HjAAmgl2Wi+Wyqwa3Vh
InpV44Cx78VPMxgbCCd/0M/3k5x0KbdcfTSROYi7arpe6Sz49fxxZM+9RGRBO7YJ/xsfCF1de1TC
VGMAZk435JcfcUQaXXgpGaQAAJjvWIscaJMkRHt0Z249OiyeeKXWlH61VUw6v7QCK95zi58yXUkm
ZhZ953mCzjobdYx704QVtA1Ya4XKl7dzAzjcr21GJ9hgEuqMykWqZzPEIUGDECItPWPRCZ8m5FMZ
9m0/onu12NBRiT6tksMO7+VXHJDcni5uy0ly7ZE6uMqlIgacv/ZShRa/NjqPeEUzCUyRGvaBj/SI
6/F3Y85ZsrlwX2V9UD6MTUt17o6CgG6w+v+18TV5tY+f7tYYImk7p7ZWitNIJSV/HivLRBK64U0H
ZK4ef6ww0k5BgPMCJgAo4c933EHkokpkfz/a/78ucM6yLFe+sUao9QnpvxW8O7AL52ziJjTzVr9J
Yye/mtpZtlCckpXpRSfbPLdtrmdzpx0/JYk307I/sSQCm3bBjqogpx9ORgKWoLAh/5mOhuPjl+pT
bJ3U7MIPDphbGmRsyAds6HLoi5Ar401+ZU9Ixj9ei/Apx14g2Fgzdvkzdn3XyTNl8V7qpf+sBiKO
Jqm5X+BchBHVh9F+9RKj8nb60yh/Xt4/rXJkfRA1V1warvg/YELMFHDku1rq5e0eErRR5c9RCt0T
DPo2YGqHXxa9NNMjbZzdvFT+T1ZvKZxEIMw60wGWUceyhj2iurmTiJEdPSYDY2DYJi5tyhLErLyG
1ZMcDpEJ9Cp7u74m83HIlIh9L3AOfWGHaTuf5TvK625lEHPOtRlf2o7O1xiujFiUNC1/smjbVCd8
tfCSKQxGzzizqkfZ8VZZPkS2l9Vwh9nzGgbyxGuswM0soMx0RZhujB1XW9dNkJkS5plVMwGtWWb9
tG8gEcWFdkVGWSZQhwtoT7n68qrvZcAUt0SbIJc5XzZVUlSuXuWXGlMq/KxX+I/t58zaQASPepwE
YaAkLuGN8i+4/jFvHc47q0C752EhTz6lvNG8MC0AJkvsaCrsaeBqIqdnrMwj2KHNualwyUD6DRQP
HnN8URYiSpvueNhxXTosFixox+31KlxGSAKudm7tIcXMncTngsmVx4kXErssUYXM9AQKHcglmP7u
lD+oP21tehSocqIT4YMGaQAcon5ySgtuANcS39MNaJkhXmVmJrbI+C5Fr9WZ3naMiy4Sus+9IW0J
wWpEtt9PBpEK/KRK/DOikQDYODPJLhT/Fnmif5I83TGt6O5tZg2+T3ODg2kluEZbgMv6cWd9sl8M
Fyn1gMGEV7Q8yMnVlXOJgJaNuBzhLyEbkidzHF0/IE0kzfpX2IRHNfXQt0lxE+pL3wU9iM8X5Yv0
D/qvEZBE5nzI91P44Rb5wC0fzxXZAsyp5c2SxVfGmf3E8QJI8ouFp4DzVDqEkB7Qx4wqwOpgkRtW
FU99X1r69pSY/2zsZPvc5Xtx1OHqPRzAAO4ST+9IPPMYfO6lvDZDiuWahl+QxhPrw0BSYkxG/Dtf
e24mkoUqyxuHmKgRTGxq5h1rW/R2N5s8Lu3MYs/Jmleop+jypGFaQn+S0U1mI0FbhgCW7dH9RfP8
QU5kfWTOG8ta5C+pKUVzQOpnPlYQhW3h9Id51OszP5Yck2EyZx38f0QnkKuorMpVLWmgeor3KNQ6
oI/XQAi18x/B4PLwma3ErPHd+3dQm/CQNSxLyhvDaBM3V8z+PIcxugE7b7qvfLla3FsawMPdaGz5
sMn60xe+fiAsdHbL3efzK0DMaFw93QttTz0k+XM4Krg4K0a4KrhOiLWXPm4MuMyzR201R9IkwUuR
JiB5zj3UCy0JZj7zDAF0lg4FDUCCyPdrLmo1VPJhXJ8bfmkJAfVYZu7I8dB4EBQYZcAcEfB2THFB
UQPV5FZtncHbrxVWFvqmxmpSCPozqm4L3tqzGfbSB98imeKVaBe5CuTL/p6/C1bFCugMpPypk8xA
pEhNmKQp2Pj2bfLO2YxVcOkYbVCuuM989eXT/d4joCC887g5il2WbIdnjYWBJKmw4NJQNXYVhX8x
Xl5/ByamZPyB4e8ap8Jhhn3j4BtthmKa8apZpYS4fg2hXY8F3VwW9cQV1KvvZVs2fCjOR5kyV774
nOrYpehU9btjAGS7heLCwDaM5u4h2560u+qdu8Webw4Dzpm6O+TjUDJk9PYFFDmh+fgPBBgn1VSG
pSw1zI9nfYXvWGyr7Zhe2vLtVbH+WyBGNmCjKKKJrienBEvCEaWniv6SUn8kd53K3MI3Bk+0wWIf
c67CW3ZYRo/hARyer53E12lerByZgD1punPuVbic5qpT6Whrpzy9Wuic5KGAK7dm1yocf5tbRuFQ
n974ByNtnRkVawh5r5X1Rr0G6SOh4Xd/78jevmAgKPGJwqz2pDpUMzFKRNi4q1qXxXc7WgYJKm4k
v9304+N73+J/vrwctBTszO76bqT12lgkEmFFY4Ika0Fud4m5LTiyZkn+xJ1ZnXSG/kBGm+BPXWZg
Rm580/t1ORQ5Wnoe2W1TN6JRwCdKt4vz3V7ynrovpQRj4w2tn23TbmPNDmPl8iCh8kuTOxEX4tRs
2Jaow8jgJlGaX0ja6ThlHebg+L0Y5EgsHDaRAKvm0pUlB3SWOudcrMDMgT8DVHiWtdx8O/oqXR+H
WT8GuBDbAZdnz9iHCDEt1h4+L1lUrwiAFOczOrCFYAj1BIykLoREWXL9Ga9CG9OTsOHlMdZ1oT7K
2nLITZTI7fvQEUqdpfFQ5ZlQys3oaBj22lVnfIZL72lvddifOzVvvr5QP9tFFbTZ/2h8Vgswgg2v
VGBXfwl9T+EbqUx7hVXO7UTFcdUX6BYWV7OYfFES3CotvJw2y7I7V2vojshdRrXA6sFCE2tRdY3H
2qDjF3KTGxabIKId4PmyIaIjZwhiJn0SkPPxA5xygh9ObwfoTcTWr69/+OBn097upv6jr9KMoj8B
jMfpJE48rlU2ipseSyhKE/Z7zlD4qdaV4nfrB5JqaPjYFnT7YWvXFWgifHZ0Hn0w274b96DixQ5s
pnVzfstj8FNiBoyiZbiWlXt+HQWxWlmPNS55IqRmokvpuKE9iSzYcdqsJTKoNkJFp3Tf3/xY1JWA
LKhI8J76xx8im/92vBGKcVWFbTlQA9hj0poS3JzmL7qImM8Ue1EzgqbgJGEpfNEUFOKIbREFMUlQ
J8whWCLwDYCS80GyXVjUfHAOHOKmFhu9GXvJSEyDPJl8Sn5OhcPfqdqV/ffydANTnFbb29B0hgF3
m0BPHlf9VAmDiJSvcgZIdWPES2gzjUBbr2VamakHccv7J+T8CM1H9iYyqrJ1Oe21DupXEln7mb65
8thb0fqtZ4+EK7sDjQfTeDgnPzUbg/Gv0/deUYo/ZidbNJDBsWO5KUwHRwMeTfO415P4RYHaITCZ
MmCzM8iDkP/KCbWlwtPi03etWtXqyMISUSjCObl19DKGFsH38CuvxEFkkSLBe/GLiY9TwYLxEiAz
2GmxKmuMBmV5VLNKfCrbCZ99P7z8W3GO6LV+BqEatwKayQYUtoxEDmjTU9Q9gtID2YWhhvHvkXhL
UwFDoU4nMItObFnVs1Xb2TtUSp8sht1ofsizyH6ivVHA0XjPQs1Ra0wZ4QyXThyZRhjEu491x7ii
A/qcze6GdV+8rBs9Qo/UUpkX31dg6QXzCM3GYZLrp81jyphKymC2QbPgk5vmuoqwsbgkRd1YhK4W
9gZ+M6V4dviWHLtxhcuLrFdC2HQZdg3wjErrJEHe1KvWcqXpV/+axjeCGJ6yuOQxrvfvA1PerBDS
6La8FWeXeyK/FPiIGgYVYRw/8UB/koUfiHjgwq+fJ2gBDd7s7xcj2+divNUsqD9EhJlKSLCPEu7g
Alf9WUZ7DqyZ2L6YTOL92LLU4DoNevKD2g+o0tnCO80wrI0ZPpU08eBz6yX6Ej7bQLYZ5zkDvikd
3U+WQ/Pp8qBxdghbGLqXvCaUJnm+5MvzXqV5WjWZhTHSZ14YtgMko0HYIUeRed4QFio4EBpmPTWc
sAo94crwnXQtoQErs2FI1f2r6rmmcuxhaDPT5o0DntyY1UEEPVucqGX8w/2U8UFHCN2+JqOR8/FT
J0RYAY/K+tzYZ29DwnATjWhaiQoSQhM7LFj8afiHRnJ8PzRj5sFHjXLU72cIUQ4Skml/DFLcdal/
xPNnMaAV/UR4CV5me55k4f4tLjeD05Totcbj0jdTgpo0SIAPCRuWp8Sqkr5cEbFBWTBjLo1JlO18
9MMAKW+xwqdeDeM9KRliulMsgugQnjiuVO/4jvSt4qzns/fuKggT6eYH3XbO0xKZXS2X7txbzHpV
zT6gHuidn4/z1qMuDDARVkY0pZuduxxW8oGu9/FU6xQLux38iII1lDzixcowWZEmID4D7wqfqU8H
v494oTTCKsUSaqRJulOaNdInARRsoArYaOvvbn5Gyi7K/CgPKzfCM9/yfIiaKCS8chttyrSVchG7
YNvewOEnP9QvqyXZTqV6UQ8nPbNkYFzzHaHo0Nxujmm1ooWz9R9JraotcsYvPVG/41exYKZndCfh
A6ym6SyIM8eJwUykh4Gwxp8XbS+mIL8/W4+Wxok/3sOzpCBohPK6a9YeupET8kr74B52OfaPIWCD
81qScKF6zhmzo+Niin19goLTBW0sOgae5jIQWqK655vUcmFvPRwe+L5MeDtoeaDTiLSrOBPJRzYw
je5dHorKmJG1wg==
`protect end_protected
