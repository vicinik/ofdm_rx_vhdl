��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��Pޕi���>da�wz�D����0�֘�n�M�zD���RB��0�'��Znp����A�$��e���n��ϡ/[��2�z¡��g�65�?���\:Ձj�z�ܺ�(󲁍-ι����9ٟ�`��� �PFy��/_���*�ܚpٳt6��ˆ��ѡ����[�I�.n�ϔ^�'��Q4*���k^�N����M���&s��?c��uod��57��f���s���A3�|���y����@��-1���4�~�x�#��@��V�N;pP����c��riS.���ܶR$������S��c�����,�ؑ�`�k>�{���1��Qz�.]L�=�|�K���W��*�I�t�̳�S�s5���p?�L�$��aH̝r���|A3��Cx�8Ir`n�WU�hlw�/$��F�?R�L�v�e�	I��ɗNP�RƓU�p8�geJ ���#�$2��m�-J<0��@nE{�X�ܔ�p��;�*���uR�����H<���\X�T!�gkZj'1~0ʥ�3�j�UcO!�Bu�U�XM����Sp��3쯿��tm�4�NlM/���"��h���|�#�v�W�i9�Z�׌;�(Ӄ�Im#���qU��y�	�������߻�	̦&�`��
�d����xr���a���F���@��icA�����eG<7%):Q��SI�iD��A�@/`�!z�[���M� �e`�ǃ�X�ݚW���� _$�!]��~��U��)�����qۣf��)W�4坔*D�΀�9L�ѻ�}��F�?/�4F���z�7H�b+4�\7
k0e8M�fj��6Oʟ�·6��b�b�A����Eo�R�	��/~ 異.�"ѻ�X�]���z��b�(�2��Ʒj|��u�ț�tv��
��[�:ܚ�w�h`�.���j������Վ-���������wr�����k�(�
j˞J�'y�s����iդL�6���$C�Ӧ�[��c��V`�����'Ӡ�I�|����z�&b��}k-~&�O��G~i��[���0/4�M�-�O?��Բ4c���FSx��*^���TZ%Z<?h���(��f5AM��r.YʩV�,��ow���XkXݏ���,��Qc�(T���5��Ĕ=w�����O�w��:V�d�h?���g
6�(̅�*��i�4<�Hő���9��	�\W�g1�Nu�F_�>���.	 zD�ݙ�޵ l�a�mm'� �Q~;�+��AyV�C�vIԇ(濅5>��W��ج*�wj�[֕/��C��f������4���J7�)�Y�2e�Fx	/�����9d;N��<�5�����|В��l��L����7K�$O�,0�O<i�M��H�q�l��O��O	·��kn�Mv0�%il�_#|v�6Q�qa82� �&�)�L�9�ث��VU��1ȉ >u�̬6�qe}�	N�=�u5<���堷��q�Xf��A8X LQ�wH��e��>���Y����C;fsÕ6H��B$A��S|��4����-i�'*���U�ngI4 v�k�&�Sx]�M�h�s^2g���7)D�H3>��{�(�ĺ71ʩ+$1�m!����? �S�)K��xW@>�):ѕS��G�_Йb �&�0E$��w{��D2rsI�4��?��Q�Uj�������L���loY>ߗB������=�%l��C'���S@�5?q���Z���������s�<tȮN!	�����[陶��ڲ ��n��~�{�t�)�������)��Tv9�[R5��T�~�_�p�I~������O㻑OJ�fx/�����S$ba�_\w�� �+Q0N6K|nZ$�ڲ3�d�##�x���X��"\���e�. g+/i�v���8w��s�w�C=�ƿAk]�A1�1n�l欔�qw�����_�w�wv��8`ӦjETۀ$�@�!p{�nC�(�R����p+J�ɽ�]��3�q��q�	b~��xf�29�I�F�j^N! �7�Hŷ��7�XrO�>�!�P�����f,�D���)��$,���������b�&�{\Jp�����D'�µ�Lp�a�^�i���ל��㛊�0Lm���[���ݽ�.�1V�2��:%�\�/�z����>�����U��f ��Ɇ\�:�g�~�]Z�@=�^H'��=�}W�1B����M;.�)��i��T�t�8�/�-�.V����qo#��[>����)����NQ����� ����� R�܊�Q��P���,'$�
�Oh�b��?Xy[����՟1 ����Z$iߟ���K�֓�r+P����e)/��	���ZER�S��iV?U�RC�0CI_���9`�s�a���[Pk&�@��x@e���Ι�}��t�$���U���r�e��T;�U&..D7�8E`�%V�J�?:E	�K��*����h�=������הq��:��Q���](���?���d����'��������D������$0�~xg����Y��#�J�g���`����*��[-s��|a�~��e�lA�7�V)ƽ��2<�e(&v�d����>��]g�9��e�����Ji�i�{��[������Q;ܱ�Uԩj[g՜:B���mc��������k%��N(%�I���w;o�7潞�J�gpK��f�Ft��K��G���uM�^I,�Bg5��h%����;�V��&�{Z�D{�����=5N�^u�����}Qy��"%F�WC[�1,L�&�Nd�P��J���Z[@%�s(g9d�4�{��p��}���m��R�-������qi�$���͕�y;z[vӴ+�V���epm��
��N��1n�����)��ZFz�ƴє�4��]"���k(\�΋/I\[ BK		�������e���:S��Ǟ�����5��o�ab�fzB�9ضRA����X���بS)yz��;m���:7����g�yK�b�k:���6ӯ��|QP���]�h}�c醔���2��'YfJ2�W�1m�k��-�ƙ�]\�%���y��䆚��ם�����U:��ݏ�����ˇVUz�Wޖ�~��T�X_��kW�~,y��j��U_���Ii��t�LœZ�A �&('fé���w�>�ci`�����0�/lA�ͣ�2U#D���V˜��>&b
Y�h��M<����Qz<^���'Iд����% p���?����B�m�	�v��9��D�̊���]�X�$�&��|��ѣ:
k����IJ�̠�m��n�U%���d]	9Y@�i���T��R�������	q�Ó�]���܁���?}���f�>x�<z+U����?f^�mb�.S�n:��3���թ��[�^㷤�B�'�1�O��R�>}����`�8���}���6�˺A����3e���'!����5�+���c��̹"d�U�.M�b��y%N�LV9%�z=���f���z-�O�V������3e���J��G�ܹf��$4831���Er���w����mʔ�}`�#��Er
G���X�Ljæ��D��91L���k�N�!�}xPg9ً6Q�y�]g� �o�M�'��Ud��a*�����#'�U'u���g@�K�@�qP��y\�c`I-�����D��:.�xI���K ��EĹ>�XuwP���7�b�v�m��GD�S?�Z����|�}��-�G�qrK���pK�)���Ay��O��i����]�@��i�d���~�A�+�Z*�Wk�ci�|�5�&��1"�ds��� m3Ι�g ����9+�Ugkr�/o<��ذ/>E�D2rW�#�zM����P΁\�q�%r�D���<C��8c�C����#Q�݅D�g�зC�{e��>��ߩjrc͂��!Rm�]�e��X�����ك-��-$[��:�u����n����a{0s����[\���\O��͞:�'oؚ�������e,��Wh����2v�gg�<� %o�}A�[�Z�ʼ���C��MV4���<�J���=�mZ���s���6�N�����ø�v( �7�#b�%�瑕�*p��jF�n"�Z��n/�-6Uׂ��/O��0n�� ��2��>�,��`�:�����=X�$��b��кGF]l�2+}�zTIFY��<�6�2iQ �#�^�+qd$����S9�+C^>ވM�D,dwz��(3ZY��Vm@}���	�����׵�+�.'8����BS��E��mn!.U"rC1�Ol5�f�[�ȭz'���$�%��O������\�I�`,��0`Y�LL�O����/�����[Q��f ;��3 C������-Q����1����vn����j�������+C���U���˭���9�G���m.�x���ͅl��q�MZ2�q/��i��p��`b������Q~�?Q�彗�u�Pc�P|D�� �&8��0�d�����:RH����!�s����z�FX�'�u���Xd1�݇G���~g��牋W��^���4�eS�nun����쎱@�&�o��&˺�V6�5����>|� ˊ_?H�Ic��hQ��D��&������|���|����?�[Lζ��tV\N�.�]&��s' �U�*}��Q겍���8�%�l=r:�^S&�O�I1��<�}��֋��M�$�ڠe�W�z��o{�5J�2	��,���'��K��Aw<�9*~�~*��-W���k�L ĸ�яnf+�&��(�� ������Z9�A��n�(_�kD&���"�l[*�W3"U����S��)���unX���b7�
aj.-�T� 0�x	Ⱦ{=7�^���}(
u�.nG�����M��]��bq��4^�8��vy����NMҷ��ь���-t�V/�yԓ�?8/Ul���g?G��s\��<��$�6���GB�c�s��7�@/A��3Lʩu�ؽ�ᅋ(50h�w#R!VX���H&�U4��`$y�� -ٻƩ�R$�DM�6�6�����M��r[ä�Q�[L�!�v�1��/�߶��M�a���?m�O]��wiY�3��U�˺,�C��ĕ���8�fr��� ΀���&�n���0=��^W�Լ'���!Iԏ�����<��Т�f'�DHm ����ޟ�N�<��xz~��E3^�WÖ��)�f���o�r�Nۂc���,�-K�&�uv����Vq����T���`�;cZ����~�T'����_Zy:�F�Ý���w޽�݊M�#}� oK�[���mM�\h)�Dh��'i|4���8�K}X_�̽g:���_ٌ�^�T�_��i	�"`�ѥZeJU^��K-�,sTRr��몦���y$p�l�.���nE��5 �;��/�&��L��E��3̠�������2ȝ%i�I��d��� L �(o�t��'���pup��W1�q7H�&ίm��;1շaW�I���?\ֽtOG=�|z������\D�I=�.)���oΛ?M	6m� �G]l�M�@)O2�Y���7����
f,�y����Z����)���ǖ��z�P䃖�TR�s�!E��PW*+�-��e*Ѧ*��}g�8a���;���H6c�Q���D���G�-~@�]�H!ɬT�6`{���x���]�;�7���g��^vZ �|������C�,�ԝ��5�hmu���.��t��*c�!��fb�T[`���/�7�_�b�D�&�����]_]��2��V4ooUC���P�%D1g�C��������KA����qݦF_��w�v |���N) L!M$D��b/U���[P4(#�r��u�/7�G@B�M�V���� ��iu"p�����n�㗈�of��I'�,d٧;�/%ҋ6B@A6�JBI�rh\3��@�~�{~'D?0��_������壛
s����^޻=��_�&���#���H�i�:��o�	�1jYl�����j�o�*=����2�Egj���TK�e�1�GzW+�T�W6�Ϝ���L
�?}O��� VڜR��}F��ճ�:4Y���}��Xo�Ϣ�o;��G� |��u��PǊ�|b+����|����۝,��O�+E=�S�XM�J�S���i~������N�8����bG*Ԯ���B��p�x;n)�3^G��G�e!B �yʵ[K6�S�lf-{e���Gq���/�!��+X�Q���+7�S��N���"�D��2�B5*�o��g����8����0�\�Y&��sk/�ӑ���#�t�M�G�@ЩQ1Ue�4�"��:T�g��!:
]>Cy\D�wO�s���!�0#�
��	���"������8�y
Z����(e��=�i���Ms� �A��� QG7ћ+g��ƾ�����|���Om[�!zZ��ϩ'	f�1�m�P�A�K�/�@i?�Z�˃�^c��!h�|m.�C�˰�u����+��N�Y�Hm&�8�{h�㶖d
��1��:^�U��&�)�S�o8cvβ�x����%1��?ʑ�b�����Q���2�P+b����ȝ��[:}����m5�D�r4�D�]@�� �\��O�5n �,�8�>�'����������M|�4f�q�!��#���ÌO� ��d����6Q��
���1��Z�����"��="A�eZ����Ӿ��EY �F`�􆐧^K����$��V��-��_�z�.��5��v�R(�U�Lcx��9l���z��u�F�*�e;DG�9�=o$�b�Y>	5��$N�ºΝ���i��}���2
qa,�¼w�N�fH/#���xaoܨ����M�3�3=�
�R~B��]箑���el'5G��~������ʗ��h��p