-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gU8Qg/UK9yXAPqw4hadT+99w0z8jC+mzX+mXp2jtqvvLILTeUVUnRO+PEW4pQ6Cw0y4sbB3L4YpA
vPVBZ0abraXTVl3j656AYcxzr81evmp2sQHjYZFGttIS/BPFMytnV3O9J3vuyRZFSVtmUrSl39zb
0lAL5u/6d/4iRDpEpKd7vJRNE3dG2lMR/WoVMIQQT33263jVJdIHfEkveHa0jnJnrd8Fqykkqs8o
JdAlawpWiVxxaHY8kYYO9pqb1pA+wXz0GaU8UcaHs26jSkbjNvoXXq6eJ6x0xyTer+QRVmBXN8A6
yTVymep22aRj7CplW7wDzW1ZHMmv/8kstweVsA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9920)
`protect data_block
Yho4HSn8SIjh6gZXD0vl7F2YNVREC9V9Lm1UyEodQnn9GOrGByaGV11n4VSg48PBQZzO9TpmcKBs
tPi958+xHPUwIpEoeYy54Y0IahxaQInzavU/rFi//blGiBccTTNARpE0yUaGdAjGBifJ74qLdLwR
eJJ8B+31VngL9cYBEYX++KSSzcHeow8iicUZXB2Us+I4g6Z9zX9RZNAKjmQO5nFI+sbMDVKH0SbB
p6p4abWpGlqrfSb7Q/fPmkoo/4R3H9NMqOoaxARzaDaXp9l/IMUONBVDHGDt0RsVgLvOkbYJFtKY
C643+QU8hbhQWFCvmolYVEys9qAQlKup7BwU8JAc/gibaf8U/EMKL7Uvk+IwJ0nRjuF2S9Q2USk4
/phxRJUobkZQVwSMZDTkT9kdvyycVtsrX61F5CQai0NyPMMo38VAVcDNKOh+EyMc1GQ3tqsKJzqq
TmIcVjT5LghQ2WBLGq4p04nBe65c77JNU9UU5RLS/Mw2d00rze+60Ym52ebORn3iF05AxUo7G6XS
LbUsw0ulUNqR1PC9n8kDTmuLP2SQkknLYhdiAStvt/rBsb9a4anslHSEnfg0LXEVaoVr4sq61El1
lpMOEsCZ4fbgYilSIPSsDthJ5Yice+qslx9m5Du98gkdc9RNvqQULmmEgsqz3C/YlW9VhBpqHxN6
PR/uJ+Fbt4/tOJAxmrGrzZWsemEHt+Lf+AC/WRSfItzlmA74h9w7ouAcpNhql0uOG3JymyqyT+wD
LmnZznwI0fprjNE/90oOIpAzWyUDSMJOW2R13YhyA3dT9zTMA1fiXXt7SQuRvrZO5bvsmCknfkU6
eooSxQfd4AXTYwlypmg3PJBIeespFcHl49PPaFDJ7HDxvhoV2xSbWBNLChoXcmOEwxuE1tI5rPQU
tnbvp1BTUOwueAr8F9BKGjo9ixFbB3pDxcOxXHDOqCkWeFhaKlGKRTuo1ZiX0dAzs3EqH09JYgzO
/9ORL8bh2HJi0mOT7guL9u+GDim0hroGrIgk02lzGsSn+Tg8us+fZMTSD3m2pxBl83Uj0lbVe7fK
MoXf0tIIDlVBe+BZwuP2PpZ26HrhHgjS7cIXOw2GDFM0dF9pK0o33z+YofLSjIL5dFroOm7Qps0L
y6STIuVlZ9vWzyTgCQS7JlewBWXKe4X2TXM7igRhW9eJDCERt/r971O84jLUBIMVc8AoiyarPPe1
ADUs7Z6BkS6DDzmOU9wJ8kGwFZpviPOVztYGL4jnEtnOnDiMhW3/3c4MZvuu4XriDHR09XmeTN4t
Icxf0cEw9042c1KNPD28jUVHs+aNJ5VmwBmb6TiUX0ozHXo7y+fg+aRssKjHvptjmnRxHHGg8aC/
2gnMMOxk1TXddk0ecWbDl9SYF++O//SrSdoKisd54WisEahxOnKVGdTda102PxShg4VGWWfpzGU6
k6Kj2eDTGSXGJxLMZBjl7ioLf1f+GiQK2OCLHwC3LXc8w5p275/6uPGbi3Xxf+PBn+UQyFIuSPWH
9qssA3vO8ykXkRtOtLQIMOkFHs5wF26fFdmOoqGdQJe58upZYeDKFG3T1lwYTSNYnU3FFC/Eq/PF
ofxHGzLE5elzfq5mz8pfzzY2sdS3EmIFIJEzgE9hyiyIvDfXlhikMDxzqu19r7TJgQ1a1usU2FNU
YGRT4wGZNSwk3g/yfHScgpwGkjEPOopn4vBKY0LDc8aKhBQH4YPOhk5Dp7c38wp7Wz0HVs+Q/L+i
Vyi2qTnbiF861ln1qeC56Uh1JH2xWXElb/HilRjhBf65uuCX2Xc7GAVCI/5pqGOyQMWPAlGzwFcS
P/eX4P0Lguar8WeW10Jxpb6goYuzCRxOw6G8aiXToYibfceFXS1bTAALDOrq7pdMcgnWxz/Ss6vO
PPN5sC7S0wpLGTm1CQen3hINW0MpYZFm5QxNNz7KewBa4X/0IXCo50jaeSYCPf3b6VTm1w/yLVaT
oDPixSlIVjDUw5n0SRQEOo8CRD/6aaaNnp8V/unCLh+uzKGi4ggV0P0+DysESAVtxcbEi6yZ7a9X
rOgTrQ1bck1JoH9S0Xc7VofuZs0p1YuVHD33kKLPZ4IGS/9N7v19f8uW9iYsB6DuPmJ8g92pyqST
bezKKbvWr4SVzuL4mVE0X86DhRHT4GBBYeT+CJAACG1g0uCPgLVnqMtL9E2Jqjjml/ZGdvyu/EGb
dbfiLFfwKA56Xw/V9IWaR0qrCUTpWjtDazL8Os6tO3SesJd4l7RlC0AZ431/RBNBlw7tQRWZRu0P
dXxMNfrrrDegcBbAAycu3oyo1gNt2ekanXgLr65/sTtYCoL7Qtb2k0iQlLnCDEnZQ3Q6rrmvZ9Nt
FQSnjLwVNFgx/X8xowcdi+0z2k3naSQI0yUt74wmHMAZ4QaN7WaLlQopJSlVbCZlBjcxuV3pDNu0
LCrBdRkkeT1IM/hBv61w6bELaWSx4/z1eJCIvjaYi6BEglp/w9G+6p2XKLSMS+NiazPDGdZsCJ3g
/KImAfa8ItBj6kb0syi7dJqWi2Wg2xZnCVYyLlvvyNHi2BBv0VfR6ShVqT9YtTf6O1dPuTVCZip1
njKv1URY+aBDROpCxEOp+EGp0Il7/A4oemj8rguB9ictxU97yd3Srdlkm2B15RAaJoDtRDJrcKGp
E8nJkIsCtnzUGndyZMX/EddyAEp9bfR6CSJE4h+JF3ICCnQRmnaHKHN5ONHtmz6VJju4rLINTe06
L6gGQhW0X1tTwgJ5Eb0n1pOOQTRJ/pMWZGHVqYQnA5YwdMmzKMSfudHF9AXSoulv1SNl4A6XmOt2
S6xAQWofADVKQvvnBTdrH2m2Jst28f9m9D2Nc4VZpiz9dYCJG8Rfrzxsf72nFJS8t5nReVGZc9Zw
HVu/DgSLQYDUQtugsf3unk4ToBF3RFNigkftnGCR6zeSRamBaf8UJn6zE19zVWdeBFBHVi9v88Pw
pWf8no5dzBy6yDxuGqVLsQtUyQoIznhTzOAK2GAYVnwB0BfFMf9lIDk5vWFq54qT4kcdbEUfyTjB
PQKSGcg7dhy8tSfvx2ncMXwHDeNDTkI+YRAirU1wdex9Cpw+k2RDe3XmPfxhqNfwDeoOu0vWz8VG
JT0RyC2xVGBzQnXrZFJyAaTOKr/gb3MgNQVfhgGQP1xI41tyfvDjdWElAdLDfvPXcHv7CMbpxCO2
pf24DFbXyWGN8WnK/ilahAfv7rMxUTbD/aSmojMVnCLMOrfmFUWSqAlUvDTtrPXmKnnwRJPzd5Av
3Z/3531yTRzonhb498gF+ab2oPdcuYBkCncHyzbnPqA4WN9+o+GTUPDrlm2EiinNAqHTyY4YrByW
iHT8QY9BKihQ+AinYAUdxTdTR5foBRl8klOH84tQ7i0tDPU2Pg2FZsbPgRWu9+XJh/G2SSK94eys
iTK9wY4Pdp1WjbwcjmejO0AaIwQLjDsne1LkGivmUa1jUdxP/dzh8HsRauQfG7eucLK9dIf3Hjxc
m5pMq47MBDGjwns8kfm/NPzwnic98IZmhrmRTVhfaBK+9VXNg3WUFCpWRkrVy4eXisGaoW7seurL
nw37c1nyrk/V2ME4KS2xbSi8wsbXKMaAfBfwJTn8OLW1do7jXNXpmIeuHQQnAnV0xK6/Ifrc6UPg
vGZSJtCRkVsIMQz3/NGmt143LRh0lYgYBywFMxjij0ucwSdFoafx6SnwGckVgrnJsCLaTe347C/f
CZRn6DwJiX08kFGf3V6YNrX/oPq5xOCCGE+bmufN1Ip/8whZFDLYymkOIKnDZ9/YF17AofEngHQS
ncIByaywYNQ2VQVMwaCFxk3CL1w+v8Dw2IkdYW+zQE80H2lM7bpq2ed3OjxH3wTI3pWp6pU4sKur
OKZLbSq/b6HjNa6YkB1ZivZ1fkfw9n4z1zbyW8OVHytGJvRJw8vzL930PG/8wENxsZFpl1f/glci
QRaLpQ1naq0MC8jKL9tJXW60N0dEMYthpAqQEKc7L4QN2SnwaL1un9RhQJEn8WLoopY6ewgO1SM4
sglldB3Z0tuN7xmGPKnwgq11b7n/khZuZC6l/OgffbTa0L3feZtwsnuMyn15h+kaJFDMjC8670P2
7bIP3roQzFP/3v1BXrWJRbNIrz+TW4Ye8HoQ3zRUTqkFY+04LZkEVTmf0Z9rt9/IEoSDmZfYeKW+
T4NVCXOMonnV20KfxNl+2IVtWfPorC20ux6rvCr+moS/FWm26/OR4fFYQAK8yxPxth1T5gvwPIFt
6MmbH+ER2UsaJYYv4uQopo5/P1JhPK3/Ed/ADBS0le3e6vT9f1CMF9ECNX9o1ZwHvL5WDAeGFYo2
CPKYCDN6NZyhmEeARoAlNGzih5MdEk99ZZPOhLOP/LmRRuIV0OPPU4iXQjDCkECh0lCXySIgH63C
oiKhcHLbEaleeYEtR6lziTqCnlpS3kHuSlogJ2O/ILjWK5GdfHzv5Z7saCSJenXcYPgGJvD7xxp+
NM7UstNfjJnK+PxCtCt6pXG7HBjA2h9uTPXXNi1mcM0456sRgAybbLIlklJ23GgQ+CMwPrrxOa96
TOXLwv9iHypiRTefmx3Q9P1ksqb3V/UFMN9H8aEbcX50XA3zClJXS0JR78HP1kHQxY+vViONr9fv
0UzgzPFfDd2M2BSshtjcJGKxh3azUjHjLwBk22/7VOf+hapQNlgbXlfX11CZwN8Zi2ahkKYSeSTc
js9SxI1k+dW/XHW9QsSbwXBYrLHEcvIWhtj6cVt6W2xH0oSk9aWY+PCGALuDm1k43wkZtCsWQlns
KFLHNIdI5loUQK/WAzp90UpwDtGps5+B2xnUOqWxV7KQfuoep11SYJayC0GYGHf7yOnXQNwr/Mf3
ZxX4jep27c53O2Cl/se9UlvktOVumgOUe5slaOzNfSMEUai6OPEPsHdtQnc9rg3sPZmESg+u2iv+
WmutFtCIryGHLmBS5H++50XE5GB6InVfyi/Gnz5yOoeUjC/WQ4kJ1qFErQnoLGLEMWyP8N//l202
nNP+jIfViQ7Hpwj1kTOOdRmJYTjT2SsLrzHoWSXqwp6gWaVy6hWTYiSFG9fJQfGc7kWeK/KCJh/Z
sO+CGZvkxVHm1pfoPkA7n9IldH8MGaj3K9tYIjVrW/TmoxcP0iBcP9QBZHmXyASMJc/+hdkRo8+T
AQQjCnbmgAJEESaHDu/ThD9XG/hxm0SlxbG5/kvQJZDWgnQGwysglPV2nc8/yVVOwq0VSeI8SdeW
eV+2hNX+lWvA52oBqQWB4PpVDa0DDY/wJ17BThGId3tDhrhgyfCoX3FOb27xEjbllEg9krDINHsq
iMuf2Ro9z8GOLu5U4sygnvO+r8iQvp0XQQSkesprfjYnSlFSLUWgkvFJL3Lyss539Zup0AoilI0O
n7bevZvVFHEtBEQVRo4sIMouwqJRapi/obEiv+2M5zn4XScOgsKm2ilyWjYwSYxYDgVug/FICZiu
6hAjakSBnwAhck1u38zUqLlvSvxVoSPxvbRty9rZWzXwm6aLVPjR2qA7cMWm2719+lcF8SbxRuJL
05V0EQLDjih8Nfe4Zp7aS6nCLZP9sMKYFv7pndHMOaGfTxxGoieeD+mQlNxNlY/98gCuZKFrNm0d
8QdHmfuBv65UTN2E/K1aAt81JmKUpoU/aC4ZvJGHVgGcJ5HuxXRakINfssuZEmtTZncZFQUtS8YY
Nje0icW8e1wigZXRGGpweVHIPzu30Fg1hvrEm6x9KDwAtZLRH99hMXKajP93qoX47ZwmVLVtl5Xd
pzDYpLIWy+goHmXEZQKArwgrLCSDZxUT8D6TtiOMTu+eqvCqKxpIeVuT7StxSptKV3KkahYExX9i
CL6HKHqQFFIuAxj8D/bxWa/o8IvaI8m7zGF1PhdEGwbdDy0rJ+f7hJawfhrxkvofaqzjaj3mcvsU
a6DYvlNGAm5UnkDEIzsUSGWb/Af9KCPxGC/SwapzXvddl8yIX0NqPTTig0XRMY9wStYd9f5CjjQT
eqM18KyiwtS+NNZ93FoqsCsTyhrtY8MZRZIXQ4NR+gFW96IT5fu+gBpT5mkhF7wYFsM+BtZWA/ig
+kGZ8EeDSkWh0IIa4hrTS8CWYZCFc6V76mEQBPZL14SrgyW8+2/Bo1d4VibQWi7LsOfVu3zKYKdK
csOPdX5luVoTU+Zz9VSSl0/C9RYZydoExwQJiT3KQ9sL1DLWwytNz+v9p4C3wNw2gJD+9p8qlSue
gg+sFT/ah9BGCmnuPU8E8vfFTyJe4tldCxZ16TtNxzXOHG2u6nfZxwpS5keRbrW8iVVc3dfbrOGP
fvrOjrK0eG7huobcS/Lpt3ja0I+hbEjWdh9K95g+v6jpQa4pW+6BpBmzGOJimtq+/Nbt9lVfLJZE
wVmG2bfY8WgiFwiPzc2Uj3P3z2SXiOAhrb3h/VTcf2BK8B06Tf7QVAn2bhgVk3Y4JWG/VkHiz4An
BMqt71iNZY/C84rppkNat3oLGpAbWXFsL060/30v59y6uIqq6/DVwIsf7sx8tgAPwYskw7TdKyzy
y8abauPb7gkfYOxH1zGSHy5TCH8PUCHThYQNbrIf3wtnE/a1uyBQgSt7LzThvKQ39wV2X+cFNWQ9
1DMSzulSxSuj6eU8EqOa3b+ll7QbLFPVb2n/8p55IsfzPEbL4a/LUQlQBt/2BDJwUIhqDWpDx4Xl
CvyQyvto+I3idvlRz70da3u42ARlPTbqJlUDt5plL3fNR/O+fbbdtoHN4jZIm5VEI++UYLAff1KG
diLy86AIaxJh3e0AGKzkwB241gT2WfnQUzFiM8FphcwqdaQhltXbikIxUnH9A/Wppsdm2+ub9G/+
fi8hriaE8m/liLUi94Ht8+fe8WOQUrMEhLOYbvU3jJutt4cn4APcW0rDkaFiFC9nAjRHOYsGtpyJ
lau/pRN5isiAAUMIniqHuEbD4Y4avdb0+tWKUE/miw7qCO4bohuolR9TEIkQYDZt+OXaCcJq+pmN
edfBtdLMS6txHGOYiOPPQoXIc8jQ0/KMTznUPE72QD4vFYSmOPdy5GOToEf+J1lUOJ5brUE/aHrf
1ZYJpGGH/wj+0f1iRvQyb6v8droHf76o49DUZwT0wMC0mPu0nGSbcY9tFdM8wAmDJQOoDNWSIebC
HYeDO/vg794VBYInb772QpGSiMG1q7sM8i0AW/4WJxMk04zvZvWt8ivWsKm/23GCJIEHfyAndhV2
6gKZS9brQ5MlgSaEk5Bx4qSQ8Qs/NqWdaYixNZfYo0sGf5ss2O2wq63gu1+j/W+RxBgwKWzXoYiu
GqhIHCP8CWFFm/JMUjE3dssROR0D0quN9rahs6DOYTGr4b02kzxPmvN+2a9Xsvm3QlbijbTeVunA
7nVmP9DTpu6pk9ZKy6BDVA/ddgLMKfU9P17H7/N31m0ZRWILH49vhOWH/4khVw0bGtNqDjvtLDff
8cISeRxbzLXoF3j8/v1Rg6IIln9AmQhZtlgWx8amz1sBhw8DO94/1O5jwsoTXGIQJnbnYWLkn4Ak
kDEucKOj2R99adyobK2i6EaccKPeJCRJdCwnXjFlNoOM4M0TEymo7YXRrNBw3gOzp1o7UvSI1TQZ
6I8Le6vJr4VgqD1it5rW/TKTQuNV4yu85+RsYDngEvH/1ndCC8iJ1F8EdOuDxKXLQYNqgyssaAJl
2G8gphRc+5JzPhG+zuCcCnm70XkFh6AzJ561InIwWns++mbAQUkvMq5hw3rPin/4gOOXQRdfvTur
8U4P1M35/uQoyXJc6HZCpqiQhQtPrbeVB0BgRxeNGwhOsf5HrqXEvXDr3gbSUGa2wQWtrF91GLeA
DKMgow8WK6uJ8arm9M2aKbGbTnOz9w4jjhT+aXiHaRXpEYrVXhRI1+IJ7CMwxw9T5qvFRPzgAmaZ
mbPb0G4+nZi+ZHCwM3mMfB0z9x8TyOQhcPs1/bN1H8aT9YKDHdrfRev++UI3uLTsUR9w04mU6GTP
54luaEOwM3jgl0uBtaGc5OJAznLflk2BQdEeWco14OiRxlx2plfY1IiuLey2Qhe2gcR+kfz3sCt+
RhhMiGyWAg5BO8JvYlYf7V/atPhy2UW6WUGTe4ApOBAWKgw2DJXEczaJO6kY/9ClC5MXBUxv4HEM
PPWAebvah6qv3TDBdCP6si0S5cAQ6jsRV+EJB//Zm4S3FcZQ/8U0nLQDKTF0kukQhJuFf/qcjBo9
AFh/FyBd7GjvVjj7yGSSoaw+a01scjgOFpLrJXVhxQlWcvpYEO170UN9A0B44SPp8PLGHX+/NRDa
3esH4HbsUPLAE1Bqccn7h1ERlPYxTpBEug//tbd3Ih7I2zfYhOe5i6x/iR+lubNJUljDh6cT4JM9
BUGbs4nkXBLaYVLhCJttJgADqiZB/YzWM8MK04jPjSW4iATHZWFQFZQvSHtutCVHwW2QBunQBhnC
1oOS5hNynkemHTZmD/acM8hvBvdY9CkdVA2Rij2aqYhhcNtY2hr6OvUVxd1txrvb6wEePAV+72au
gugmWm9EfkYytHlk2HJupHXAy2Old0SjWwJVzo14hW0HuFGqhbYvCSNBpOypoMv4POJfthrs1i4m
QlMvnayW6J1Wk+lwTnnZY9Fal54fz4t0xjvh5aunhjJ7r1DpAtX1QccTpIN/SO/YC3zCcEOWnfwm
tzvgHY7BLSpxeKIKNr7qaIPhpIt1Pzs1dH928xnpYrOEVzgdzXQk5qOqn/uva/qvgpYfKJ3ozMbI
zlyGwVW4B3ZIq52TsseEmxlxC7thGpgLEH3dZN9KzXsyfFxhInK6jCTl3+W7miK9QhHtwr0lZsQu
qWEZl+uDGRtn0PkBY0oeNMaZ5ztm1kAUDVIIGCTWEvu+jbcKbWnLx6kisCSNA3SQAh7RKJJ1WMdq
UKWpLzHNsWUnnFLAvF3JIHXPHdU6jnf7aOftkL/V5lm5SFJPZhDLDC8zhy24ywDZgHhKjgFSW9tx
jmLAfurW1zU5TE4habTjICCsFraDPieYse4RDkxQm+opZn2lzNvJoxPO1wOuJVPeFSYmkSQKQOY1
V49KCjBXLgOdnBFQRrjePdrkOLzwXB9srp/Toh8LCgiRqQdTqYUuVXEFSgJWJoGVT5cL5jPzceS1
lIes7B0VsR274t5steaBWt++3cuNZQqce9zLbdOQhK1ZBHrlAwlXB4bDOfDjUPVlsCMQ7oFK+2T2
GE1CZFu7pwR1HV46j4hWcBRM3oMmEpXz+jCZiLw39iefzNPoN04fe/uwZAMlYUT1rwFOqLd4nzRM
2bISUqMqYi0lQZiw2YQMk5qfFsel08brqbV/t8bZhVHgg61Km3q3pFlpC2wGWZAxBVLKU/ugwcDF
Vp73mbTGBQzgIAikKvzFXdQOumRXwevAYYbdOXv6RnMMtaCHGo+WpvILuzbz0kZTel6K7H8Wt03t
TcFDOuPcf8/fvQF5sktLnW0rXJ9CBNeOg2JEbCSQZDIy6zoRPfi9DJTuNfBeZ7OvnhML3uZPvu6O
YePj0rJHgSs9vif/MoVpeIAaWxU+AiMn90Hc/HpWTCXSuK9cVdwTWh4yq1QY+GlWZi1naPj/ZEA5
44bq1Z3nDH/xVcAFef8PgcN7qTBl6MHcPYhyN9KMIjFOVEZtsp9N1mSjJK482fx+Jc+9bYA6fhP0
bXvWSbg+Gu0qGmACk2phpbffVUBzdgIrVNcyhLqTr3MbNL1MYU/78dsQ739WGW9yUtuRMF616keP
Cr/JDgOoOhxs+QOZG7vB1yruixREfoebUC09g6EmvlJLwYvqS+RxqSr7iRTqFAJILfLhB/fYfb55
K0eynU5LImfjHNX4EOFRcun/FYssxZC0sYXQB+xO2bUOu20soaCATXptvz79QYwJqjgVKHxMZz60
sgbTT3xqIVQ2X5XXG9F0ofzZq6Or6+6SExfdsr10QRhD/UTNc1H2Azfdza52km8gZberCB7IxZaH
uSl10dVrEU3Xyp5S22QwE5TAqNlYlRl+g2HHLmC6moPzf1zA8CNoPbR7GawB1GmTcWbf6fb9XTY4
/JQb8yoAGoRBBgs1LYrpqoVVGrEeXoG+RgOhUrgoMkmwlRbixfg5Fl0YU7+gDInMqKrDeis/AdoK
xNjylGrEpOamHCkiyLu8LG7znBM0R+IVB5Cmgf49Ahq7+HID17VXvfIzE7h6poXtiDLMfHT9AZGf
7/sidfJ7Psuzn5l2K3Lqw1Yn9pL574njPGJbRH8q+HAc3c6M1bx+RU3F/dtYAb6oxOzltNXVgHeP
FA/U6axKO5u6Vogj3THK3vbsAL9W4KIO4g/cEuwDOorIZ2Yi11jB3veuqKsXAr5Ckx47TW+RGZxA
aj4+BwXwswwRnSARxBxYl9mML5SURO96mjkBtRSktcmGTHBnpLnFaPMqW0eNB+PthT4D7V1KvCee
jzMu50himrERZGdVPnndeXlpr+WHQxyWbTnQ8L2EOdeJfr6l+f+Zcvk1jnOKRq+egDKfilVtuOxF
/maaKpjHL0LWCyFg2/aZUrZIt1SrrCmgQ+ANk3st31CjMEwBc7rGJ4hvY/cpboN1pcrlX/5wr2de
+k6yjekzrRPpoEhj9gNiWvBrqcP/UjAcgy8GgtIndVKk2xvLcr6dOhHKDeXAzbcqtLLnpfwDii/H
qPMXNNNe0DX0pJCS70W5q5Kgk2dsxsnuyd/A3b34jC/VuaSvplKDSgBLzNsvF8rspEJqPvVMW1Qj
xOdNQVSgK+bkswekyuzOt83WpW9EmrG3+I3qWRKhcHOb+RzozWt9oB+Bw9dtYJssUcCMdhd/5mFJ
oFtypjeqSHpBC7UDaiz5YbuexxLmitGTcLyVDOFbit1tL/S6ZLZi/FDpT4RqcTHu01AOd5lGSUmt
3H16WL7Ay9o7ZBjdbRiSrFLrI+IYh5nzOA+gz3r3NjCxsAmAbk09CRmQwq3XcUpLkaWIJ2bdzMSD
it4gEtD/Q/ZOeiDJBJioi8C7LHDejRD+zo/CxoTi1Rx0vh5eBFthssUIPRoE4LDbhOwRkHAx372i
8Gt2edx/50kFUfkjIWrnZABoPjBfZ79M+vyrm1pZi7Sl4q1jfSjJrdJqIXfnUX3WR4nhsr/z2dZz
url8J/F4PKkJPCmLypgFZLPRQvrQ1E8rnSeo86D7zPI4KpFgcckUMUOZIKlTv2UJ+zUKPdD9q2jR
w3N5H5D0dpukFwowIQtkXblXOGu32aAG1E4ATkb4GULOW2EC6y0cbT1peZ5VXKIQ9L3k1aW+0lmg
b4MlXU772m/aCghWWtpAwBRR9qzjrAMdRv0MMhO6fRZWxmjd7+nc0kjoT9wM4nzOBNQtPQ47IvZC
rV8plRyMLEfZHcwCBNQ0LHJ4WsswxEyDAgSTW4IS4qKOBE2DmBEPBX1BhtkqowBTvNjH799NQE0+
2L0qjsuWMsjS5ZVop9Z0oEZZXFzDIp0waM6r5bT80/HdZxV+eqQC7z51mgx4nBjxwADCExxKV9wE
equWNT/QL42AEAt4RW3IDQwJVhYuXVkESORdonllURP3mvD5DwWgtdtk4+O4CQoEhA0dGMNrypTJ
OLbGciqSci1AfxNtFR5EaT1TXlIie5uoUdIF0rgtvzvl21YIdIGNOFjSsngLqklT+QCqJFFhibgu
fPc1t/dAkb8qxk+wresWxPdI2ON+IXGOMq8M507usNZIDj1LkeG3yUmpZXonp6hwN9ktImrCx5QE
FqvcRPoVP2XpgiFbtNs8tHugHz4EFYnlXdio40b36hAnUL2fZDypSydW+LdwNeIAwTxh+FaBc1D4
lelLARpTkGgaFPY6PN/GSn1bzPpiU/GpRurjnN+J33kgLuknnXRvuojHCxlZK94ZGXB3T8bbFoSt
kIwURogx/D1NlQvTf1tOudR/2WYArMPjq6A9xrX4pP9/9CTkPIJ+UZLPB0Mj50HiLwSIomt8s7r3
+4qrWGdII7r9/8wPYv30V+wfwFKEA9UjIs2mjn5AeQHlJcJai15ycaNsxzatUX3pNel3zOIVlrVo
v7+iXh+9NMxN9OVL3xB02jVdxE6txdcpAfx67BYjUFZ7YF7H4jNWzUeQxykCYaahJyOIlFAp+PXN
cWyg0qP3BfI4aFECP9dzcgfOZtAXVujKnhMyCyy4w/akmcIsHj2+L2BE4wAUnp07XhUENR4FDgXf
cvDFFoR5lWQl0XDJ74+RvFPZuU6XjQaX1FX1BvzrxhLtttdbwdLS7aTxblLCNvsNdRc+VxeRvXd5
k+QosvSJ0bKU/BweJkDErvgqjSvbXxjVSA2OLiyVOlTM5A7gZYszosB2Tw/hL4/hyT/EcHlxJLm8
gKRn3tXrd5ysy7D1vcPpRBmLpeZRgyIPnAKspzBdLcZfQD4zns4pw8NrzetRRCjMmf0BDvcbCE/H
B5AbPHYeI81QSL/kx9eY5U9a6ixdj/CnQAqtmo7FdXjZLcZwSiUO444FafMUhWIFA8Vqia7mMWBP
GSLnjx0aCc1d2arsXLI4mAf1Rihbu14Y6jDWDiiI9D6ROwZRFTRScuf/Ez6YTKc333NU8SKWF4lF
Djgt/75wl+37GWrwl+JuDbwf2iBuiJRzZk0Sp+KteuQz2QpmZZGvClIRzZSIba04Q1q7EdJQMfjt
EX/ykwTz1fOQ/v56KOSjt13XfmFmLZnHqE/dhIVGnKXr/OsUZcmRL21xIolgMRUh8NnIi/3KfyBy
zCYVQQtNfzPKgYLsN6ZR/yRbEnWaEjCgIssWUeHx3M9vDYXuBynsJVd+EfgxU7mRLn6yMOpV15uu
KepurpiIzfNthSWh8VMuJOTVNk606eOQv2ePzEGjSd6hYNYavdt741o3O8OQpSL3a7AfmYICVQMM
gCPOPDNT0q9XtahNji+enhWM45vSB73S9P6qzSYuMBTeLSUAfo/oqb3i3B8MzQ/wIV9udf75gn4z
xNTOMx3dgeecAbBmw1xwj4PZc0ryi9yoafpOTXLf1ngW3yCnVoZgleh5+sCM3naz/srvGQg+nK3f
EZh5X2Un4cQV1grSzkuXotbw4pyM89IIZe9Ty9aYiTFSn1oRoi5qJovJZHq6+p5GQR23BWgcRxXQ
+M3xsxiyNV4Ljmkwl6edQDoxNgKFU0T76618L47WgdLN8FlJftDiou+IL3v+gTq4zR+MH46Csgrn
eQDA3PrrdvslJovPVzQvxCz0nSrKfruqRmWkxZXYNGSH2/VX4AbAbctEqahV+k4Jr4Gzkj5ZVNFN
QCQ=
`protect end_protected
