-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FOw0Pxh1/V1s9WWunweVY0n0BruT24jo+P4KYHt4I3CGbZYazIp4cENhhsrrrIrUbHZzhr6EWF7C
AhZdjmUrU1QWdCnEizfVLIIMlKG4RkMaJS5fF/KezX0Tn0TCovxZ1f+pnwEg07vjLuqCoCy9PwKj
8pM/nOqM3gUU5iYf7jDikr/7B2qEHyYrlyW7bZt/Tpo6qvjySRi/oEXIzNYRvGksxDNsW6FigFsB
q1XXVJiWBkzSk2Ztbzc9sjJgyDfhiwOzi8sKmm/TS4rIHDPQmD/dzFEqSVXGVwRiwIUkONc9C7+3
XuQiE8gAd/rSXBnAhn0envpna9nTmr4YgWnFFA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2960)
`protect data_block
XxQMxom6ZikSus3x1ZXl1Js5A2CdfRWSgodWFOISgZG1JqEVpAY57yX3sEzsuYveamoxGTQND26E
5LML3rWpTvr8JO2/JAJi4+0EL+s0zw6w+rwGdenLwlsjXU8jkHx/dUcAGkTGpZjZQs4Zb7N60AW1
4KO9CEA1YQQ1q17Vbqet0kZ1xtAlE2CWZzo6/4y/WZNDb7h+/tnGWxz2r1asQXS8dX59ft2YUuMM
SP/cgmb5PYOriYR74MSApdNihHCcWA52BjrftP703SGPVthUmYzgefSaagOv4L0VuxPmK5sf963S
UarUI+6DzV4N9qChz87FrMbBc2glRpqeJW+tBihuB92qcNpHmyq3VQXbCed5u0RFSbT54vPy9gys
Sw3ZVWTWXNZ3abSpCLNxSkweyPyjS/yOhQJwCQ9PfT4Iyh2x1S/kI8ACPietANxUY++kzGxAfAuu
OGECo3n//+vuqhtziApd+Ft5Mh3kliKFaKpV7a4zVhu8H3eD3YNGqs2/u/FrSGpG6bziu7/q6wXn
MAcOngubsj68n2VslyjXQa25TSA4jtj92iof8fWzvoxq4WoRu8IomaoFblBXZV4hkOpcmdPFvP2G
LpdkcZR1ok/66+rjqiMe5lXAkmEdMku2s73TU/VQTfZl91pbk3UXThTNGztfhCdOwqD16PeY5BFT
rWniIPZ8JsDhxm64kGieCVqZ3dD8zWSG2VAeZaglI9AN4MGfGr2gtNLb2XpEXW2bh9oj45Dnkh+u
31qD9zy6Vmpw+hjVDyIUxsxBmmM/vzeBZHPiUzUAngThT1nH2kNOjQM/uxWwU89kGel8c1cIYE04
reBNuuCUjo1MyhTOqbtfTT2nUNfFfy18IMQW9gpt4W4bQ8qt0iT1c1BMEV2OI5AShqXplc+MPBGP
A2LL/Z7fVdiOivq13qLeHBKQVdGlO50plmwncx2BS1F0c7dyKz5MAL+CpPZKqAOMx30vidvegVX5
W61pfPCPpllwD5mY61C3R4V7uYCG4DFWV5+rL7zqIMBztmG8f7yMNVoXXOvMtrEGVFyqpBW1FICh
bvtRFArsf0thsMPJUlo+tHfa8AwlkXilL+VquQ4ViFB3LTAqaJQj2zmMJLdPw1Of85Sz2ckxy/xc
QalVvv9Rh/DrP8LoNDr0tLUvFlBHucuszpW38N2TGNKsg+Qu9Nvgg44HVam26waoCwmquXFZfB+s
Un++NaLHQc59DS8AwzTJxFX07IAOpdGrOh4F2qryvAcApT+ZT2XRbpeoXDYZw6+rjXlGrlhQVh+M
nZokHwS9eyaZwWZh0QcIJIU6Rv/msJZrV0HhPerI55TaraFsiidn0WNrHm7ArOLepwEbR4dMXYtp
lJzZKlTt+Ib5H0ijGVLxttYt+yMPL/Uymd+qv6U1sRbCYKrIkXGVHi9CdIuPziSDKU298eCmU9Cu
oIJU5Xo2BI19JcPdtmrIRPkSWXcweXVbZJgLGLnOZz8G+ju5rf66nDxKMDUq8isnkQHqMkxTQAFy
YrsxorCpPF+GjPh6Uw0LOON4Gm645/LGEIaTNbLJz9jVS2AvpLOOdWZnvcjw3ap8PEOVM6+SP16k
RY2ymAjlJQAfmh99NKNqCh3fWB55Mp43VDM8r4Z6IX5uDZT6SXSqSGHBYL3LzJZzDp7XG8pK+e3X
1qJoPwmJ6+xhKnM2QUlYgZ8zrEAKAHgCzC+4nMpzd6CQm16ZKlaNE/uG2IPwYJ+8hX/YqshF4nQ3
J1vyyp+0h/uSKy7x2Vozw24BimYgdHC0rnc/Z+NFN6VSzqHwv50BOmD/htjK5t4ZnecmEzdZ9ymQ
Ax5/ycrqLUyPSOP2sMdTlgXXjrRozrwgSc2bJR7zw8QlZNUGC1p2C9b7gnDk/zqpJP2a3SBTw61w
DWaTsLvbIdGx32uRZqQGCp/BKuIXy52ciofsWTdAzBssaEpSzzLVrtz9n0h8mGAAuZUfceCQK7ah
g+XaOBMlXpoZV/EHvSlppzm4h3iuNchC1JtxWDBcyawPJiVZBpY01ZCWHkjd8geyG0qPVjR1y6cL
QFNtrFC/0kATckiEVh2DUoQEQnIaC2Im/sI4JfdY7XPgWTic3n9Lk0JlKXDJgW8/D71Jl/VlFHdV
s09Cwr3eJfnmCyuCR1GkbTYdzNeEBx6aC21avgqzn2U+YNVE8P6VqTyD7B49JMbxitqnmannG0Lq
Trbs3JGosSOGIhLd6Gld4c1t/KPWsVS4ZSNFS8iMid9wq5J/KMwX7smDU2Kfjg7TzvDSE1+PHror
k+q3ZN8ubzYR59oTk/Ov1pOwA+RxTqKZ8PAguuTxB3VnSOKSFnxdnfGItxrmwym0vT6MsNWgOTFv
lUAgxIN0BHmt8iqKkS/uGbVp6ewX/ycngNlMFSidcLqcithTPR7cUUGn2BMDRGj0xW1fAWG6beGw
xzEyf6s8DzGC5dY1xeJwOEBlBbZ2pNx2ks94yi5Qdfxrz3/0ucHEdD+X0a0grdgrcGOdp6lwkWXt
b8g/rEhkY2wZRoMrLnn7WfY+wilQik/hp7wuYacPmVButj/rqMxloUAabD5oVD5LrrboWQqaN0d/
0EgG5gI5ESYvN5lZ08LTKIP8CNzGRINGftzdCSuX3uMNoqZbheXOyArqRsd+HeGUOcMp187WoDEq
yne4A386wVlJxxZo78rbWNgAnXp4YiPijcrfSLrRDSwhBTbcyUB8rnwn66IzsPHl1Z+67HDe+yUC
z0VvOGpMGvFKc7xAIAtzS0s5XQXJ2s37WkHZyaWgbj9BwBiaFAvARD27jU6KUzduZz2IP8XDUcGu
ecD+xag7Wo93EAaBOKIE9owaHdkv3QnNni0qVcaqq2VBdRgDU3fLqTw9+gfgLXiXX8LqQQF2oTqm
F0WGgK9OnijrYO0nHbxnhbr12elymNxtjX9KYQnLAHbL9xVdHYPnT2bXmNZfh70AoYpF9Iv1JPvv
XHrsdxHzIe57LBvUZmGJTuXP2NmOBcbRuZIDa/lxzA+4mUzIQ1tvEEzy/YDi2cKhp5pBeNiFToFa
1SFxq0JUo9jKkbMlyQVQZ5p2r7siM9mlyv0FgeOBe5LslyObMcK0QFtS42TOgBay3zW7ObHZwZaF
t/GQpEILoDaeMV/hiRk/68tJY3UioMUaRD3crYZuSsvbh1O2hUOpLZyB3HAy8rbc67qc6Ij69Vli
7rhktKd0VkKMvpDG5eMCfMIFE1X5wwYccpt2s0ZuiELWlOz/7soHKBF7W8jotlDwPc/9txGa99GZ
C81R3BGS8OZWC7xHnFqxWSSj4IhHP+TPTZxtw2p48AQ2YGQUYF7zORpQLVEzb1egFM0eeE33diUZ
6IRUQ60PvG6YF9Wg4s89FrEdxp4kTMAFX43iamFeBokxJkNqM62/IwmKYT3aIt9dLrJGoukje3E0
Q1xbEkUSnge/hn0ZFQxBc1V+RzYoMdVY61xQO8HyGar7YU0eIES9MB37IJEMCcvSYYLtBCo73Gxr
P1P+rUs100ZcNWlCjF+WevYsu/5Q3K7kAHYy9dHjy11dL5cd0jT6G1+N7OGeTSaWYnZS3Vrayk+N
rhgXaL+VaK6Q2Q9VVvSHYg6H3fJNcvfdQ1qdp6I1slZ6mYccOqtIUDwXOl/nI9cKUEtTq47tIqQ7
Wp95UOsJMq2Q4L9mPCg1cknsn+IJsle5Fr86HLvhgcQzLIeFB9+3kLSAkM4pkPTjSQCQIhBnTpMM
BsfmaQ4eWWS2hel4nHeYHnGJGBLtprwQaBsjYUfg6W6otQsQtJUkv6dKlDqJOssUdP3R56F/wzmV
XtSpHZQymIKUQGuqaflQvowoAQ2Yp04GrdszFYlBcIjDQznZ7wO4arStNwbS45hoXPQz6Kb3Q59W
M0YaVMgpDUoPQT5SJVziobxstSSbk6xDc6bc7IuYIgOBnEwJ9NuzKqv1Lz2FpiM6ignP8Uw=
`protect end_protected
