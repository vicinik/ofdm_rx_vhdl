��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P���S�+�Gy�*��HB���l�W��y얷U˯��E����ٝT��]��b�S��0��~�&�� Lg�.Y�??���Os�����KQ�)
�ZP����Jt"6)�ổ,s�#)�x:m�K.kt;��¹�����<k:o���J��!1�a��w�]�	�ZfŬw�w�<�T��6F��SL`zj���]�Aug=];.��?<�����UjxAY375�IQ]^[y ���_��K�s,f���Be�l���3I�G7���pP+~�P��!�g>/�U`1�%�FfT�Nx+��V��f]
�Y�B�lD�#��ፈ�޷��3C��� P��c��%����N�6&��V��\p�qB�������5���A��TrWzO�;���B,ʦ�F*zS�gdP8�	y<i�c�M82�f����e+�`�moAC5��~K����|�0q�^������Q���r��J,9:u�[�p���ʥ^��8j�[�enيsn���zs+�J7":fǮ�ufa���ݵ�(��$1��.�
�d����2�2��ӫnw#jK�=��%2|��wh���_�fBW���� ҄�<����v��܀0���bP��U����k�[y2�����:sl��o-VX��=%�)7����{#�VBFJ�
�(�~ܯ�h�1�i	��LsCSe�d��0a���U��6��ì�C������IL�	X��*2E��>e�"�Z:5���Z���Q������n��������-2e)�\5�m���p<gv���#���,���m��Q��ʍ�Zͽ���FţÄln⠎t�UnoF~�P��C<����n�Ѝ�K����v�,����wQ�fI4��h�����t�V
�]�xA1��R3�d9#m���^�X,���z\�u�Y�t�'q<��=�jv]��-	�p��"�������[n:%- ��RCP�&��<���&��s'/M�_��c_�랩c8�:�����yIei���~���RY�N�ôe���NR�qo(��s����	�k�8�5_�Q��|�u��S+�}Cg)�t�L����J�	�F�Ġo}���gv�&�~��k��O��Ѱ)�l��%��ҝ��[�:�q�׉���N?�� ���]��1iɾD��j��)O�����W��jJ;F�$�[�c	���ܮ4��/b��U6�/m(�����i��{�˩�fr¬pC.lV�an���`��(S�/�,�ݤ�u[A��j��.�59o�P���D���0YYIL[G7������C����H"���-%ʐIT�lf�yp/O�Y%mG�8��2/��s�$����e<��+�ڰ���&��Z�,P�Q�S�+/��!eo%��Ü��V�f�o�'W�Z�	�q�<"!u��M\�=� `x� �}�c�f�n��bF�L\jU� 
��֤'��9[��:H~X�� �31�e����