��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��ĕ�Q�i��hb{êX�cFk��]v��z0� Oh��l����[%��O������K�n"Ɲ륔�[_vp	K�c�A���x�E��^8;P��I�[H��L��v�Ix:�ie^W��a�R"�=N�\�-i�	A���c<��\�W���tJ~Z�G��~7����|�Ie �^���}�И�s���=ɑ�r�~�D�ʆ�Bkr��
mWZ�|T��;v�H��p���剿>��7��tE�eE�=~� ְ�1�I@��� ȇ���*>_����bê�����娵�$�M���.�S�z�����Q�=o3]�D���uR�r�@n�Z���KP��ښ�F�PWe�b�x ��SE�;�l�s4������o��uv�g:i��[�+��gȇD��]�W�o�t��∯��$��lv�K��jSőY��f�@���ee�Yb�q��p$��!�'Q�ƻ~����}�s�(���h�?��,�N�5��Z�K[@���9�W���N��3���!�4\�\��o���(�y��(`�ச79��(��Oq~�qD��S���-�ݲ��Й�{}�hJwQ��ue���(:��O�:d����[�
����u�ƙ��q��~��C%��yր7R˰��{��ܠ-��]	���&\vE�UE����/'�w)uAp�P*m�!V�:� �f�b����ʡc�X��(����>�l��
u[�kn�,��[��렝YA�:�gCpV�F�z>��EUv�������
d���B;NŔ`���#gU�3Gϛ[�6�����(#hO9?rm��"�v2j�O@)sY�D�Tw��>��߼�%Or�-x:�H�}��Y��x j�J�S n')R/:�{f �Cu�6�:����Fa+B���<���ǹ��A��mf�?q.5���\�S�P�M�����t?v�K��h�DU�qk5�����%����Tq>i����|�4�4S�a��{y^xɓ=&5�:�%�� $������*��G8�c2��_�.��\�_m�|�^�����@��O�,�xE�WU[NT9�("�S�m/)ȩh��W!\�MF���JL��:��Hgr̹�o[K㒣�Nm��{��=��+CK��P���Υ�Ƞ.��j�ks�@|Q�������"����b�+��gm�����B�m�7�h��2��&����߼���J�S�V���ԡ�m;��^8hG����.�P�M��<�>��d!��i�aKV}봭zs�w�mæS�XV��0i5сۡUx$�d�m5�,�Fi��vvl�(���ϣ6�>� ���/��EO�]�Q-s4e�1���&��H��.&4���k�Ld�r�%>�PM�c���C�ލ��:��/�|��Q(��-����gH��(�P��eIlN�:��|��{x�j����b4�j���)����| �`§�2�?hX4Q��a��t�`"wG�!�
'<�9���XAuOo�:轜5���d�LO�ƒ(̿-X�,_7W�%�;�~ۭY���׺ ==���؊�R<" Z��u��Av���&��g��`�Wr���k�]%�{��W������+u��^?�#��O��My�� �ң����>D3�i.��dL?�������bS�,���:h(����!r(e?V-P�u�_m�=��(����sk�u����+��0O����KW���wBs�͚��G�lu�{��s�H0E��~O��r�L��B*u���R�.���{oG�����,��}�_*�q��d�9<bSuA5�R�!�E���E>�i��U�[�
?E�?����ZZ�s���YQT$f��CS�H�-�3�	���|gi�����p'�9+3�(�4�4Ұ��;#���x��+6m_gޑբ��T/K=uD_8\��u�&e!��s,�����TF1��܎v�/0�s�4joWT���ʬ|u��E�fWT��=��m�ad�&�ؠ�����T���zg�+%o�ڠx�4��df��t�6��b(^�-.�,ld"����y�S��M�:��(6��@���������X>\��R��
�������!r�z?QL�j�wD㙤{>V]���|�){� ����������������S}[2%zlqYTV���;_B�J���j,��f�0�h�8ڴ*_"�f,��XBJR_��>�������X�|��^P�����`��iG}�]z!.�����b���Lqu���>�5}�ٰ�T��"؄J��=E�4B[Q�D`)��c	��?磺[筼uT��WH6�A�J� f��w�5L�}�	���Ҽ��Q���bQ07�!�zMk{<�=���3��y*4��rX���9��泭%� �3���(���T��UCd�'q�, ׊���� �X~�����b�u	�ڳ͢�4��d��Iz]t�i��sit�S����N�73���$��o'~c����,:@�Z�t�: 8?o�T�U��v����1��X꠰�����%�����"�e���c.�0*�������
�pA3����h[�1�F���$֓w��H�K���Z�8�i%Ȁ�i�C�S��9��W��؞��r>��'x<�kf �N��sD���&�̿�2b�频2Aj��\t�b;qI��)_i���R@4>�U�o������ґѶu�)��Y�Z;�0��c�v�� ����gl��x���T'�Nnkx?�W�q�� �G$U�Gϵ�nK�p��@4ߡ_q�\��
S�u�6����A�����	����e�->����(�̞E�!�c�K��c�Y�}2$������w3����=խI�!O�m��,giH&I��,�7��μ9�����_��؛�lt��Hz�qjg�r��V���1�h��j�L��r��em%u� �ɀp�y��0�f���;�Z)hF�}9%�c�vC�'k)����V��}���&���%6��M��YS���K�0� �K�,��FrX@�@>�MӞ?�!q�ݾ����0Q�i��2�]~&��-�kd�+�|SW{�à��X��{̣�J�٩<���s8�X���:���+d�ŲB�6�(�ʆ��08íu��P��.���]克�7�G�Po`�Rd��CY"x^;�G��MCP:��7h�"��G𭳎�~.��[��r��5�Sp�AW����SE
oT͕<�;�eL��P8�;��ַ��~�ւ���@р��Z�V�f��h
� ���iZa��D��,�LY��	-Gs!��Sn�RJX?����^B�P^��.�>��C���Ӫ/v7�4�Ka���nR��E�6됥/�U����G��/��	�C�C %|����.c�K���1������ Ɲ��a������a�HYXY���x0�������S	񽛑��D9���q�D�`ߘFG�
dC�f�"O���6LM�mm:.��w��&�&�H��H.=�.!�K��F�`��%��=��?�w�x��l��C�z���=ʽ�hJ�����_k����i<!��c����ZÛ�l��ov/}���W!���-fگ"�_��mt�z�(fP �yEW������ȖFFWl�c<_K��J�K����#=�?ԕ�u�ž��#U�p���ҁ�j��$d"��
,I��vLQ�n����98W��N4zu�a5�(�(%��6@�~��� H����������j���QxG��Z5�<���|w��������T� -[��A3a��b�1Na�@4�w�K򚫪Ɵ�u/,�5ձ�P��x[yu������t�5���$�Fi0~:�vn�A:��%�7L4��*���|�I�]�;*�Y��'%��8���� D��9�r�� b�
�!]6��M�+��UKM��{��X�#݉�4>lo�j�Y4I�M�u���-��� ��'�#�4K��6��o����7�^1m�k(v>4�g���F�
-$���y��R�ǵ�'+�غKہ�<���ЏǬf�u�9u��|��D[Q�~���늼MY�F�[x��{ٯŠ�{���B$f��	�5z��h����q̯�L/�e����!�P8��!pN"T��fz�VAa�LFDi��B1/�y�K����b��B�`DL�u`���n*�礳�d�L�۾�P�`�8�xѢ���������=�	��+�6m�-lP�4�%��������CM>�m���M1}l�"l�x�6��(����� �������* H
���.@����Q��(�E�3����W��,��Tqi��ε'�,�%&�Mo=�m�y�O7ԍ���C�N��K��^�U��{�Fwn�1|8^0^\���R�5A%�r���&�҂%�SR�N�7m��3C$PW.A� .{7��x��F�� �b�\�V�]��[1��Ҝ|��߃{`:�]��v���$� f5Bi���g���h+�~�}�ʮ��,R%����tKT���ɒ1T��;��Xo);Z?�����,E�rI��L���ŕ<���];dIg����祂�*)�B\r�(�j��S �������āCIB�i�9  �ixi ���M9���R������CK*�l��}oEH�Sۜl�ۂȠ�_$$�93��{��{�����j7�1!N���c1��Y��'�:P�����V�.�5g^ْ�>�;e��f�R�Q�6�f�ġy���'q}c�2�5��;+�����l
�͠�t"�>#�,���	� S\&!�$jq�c[��.[��'G�}-U�|�Ĉ�
ke���� #0/�\L,Sp�����||a$м�m�� \d����	��'�=�e`N��qz�ʴ����`!mԍ�����Z��Ϊެ�	���Ae#Q������A�Yw�9Cr��}G���M*"ɂ$��
���-�Vy��p�:��5�]1�@�E�
hs�t�A���������i6�C����K�p�K�	������B�{:�ϑ�9=?��U����-��$s�K�}W��!���S�����tM��**'�Uck�1!lU9�,d�-�37���'妘C$]�;���	�\��?;�ŗm�#�b�'O��cH)���pɸ��$N����	F���ѷ�zK�pK`x�^<�I�&HrL��X3��L�m"��{*:�Ooi��i�� hĉ����zE�ٷ���-�Y��U�L�Ǳ�L �w"I�Y����?�'Q��\Hd��H얯�]U퇮G��D�bV� |xf�\��H�G�E���=c��������v����<����m��<�@��5QFD��$*����K#>=�\70m��3�'o+��}���s�7�1��(�Tg<����1��Ι�R�X��C�� d�t���u��AWW=�P�C0G�!)�H�J�՞Ad�yf��|�_x�]f�9�*E�/��75�1��s1L����uV��Y��{5����G�b~�C�*x�ߋ���e���=\ȟ��5�����i�~ݙ*��vP����5��E�ks펧}��]��dȍ�l��Ꭿ�*ӦHԾD�h�Ӥ�%8VH�B�D/���~T��q��̿�����U�R�-Ea.�*��
;�ݘ�0�;JZeqF[�Ԯ���\֖F�4�+_�rA��N�q,}�w�oY�L+U,��Y �
�V۝���K!J���1�1Nj�Oj�ol��f�a���]啐��#���� �O>ɗ�:����q7����#��Y:[Lo��^>x�Y2�@(��]��֌�<�g$I������a�d� �@,e7Xg�8̠���?\ۓČ��ƌO!/�*�.��p=Ƭ����ƈ���|��m\�e<~�4��^oh8�Y�l���6 �(��ą��t7���!��?����1��m��)�/�h���U�S�a*��j�5���qft����*(H��R����,�a��˛���G��3l�R4^��t;K��
P1p���Z�*��ʗz�H?eF�vo�����H���g�(~��	����*S~d -��a�l|�G������<�_�/�t�3�X���^#���#�t���1S�.�@�EddM����;�t��}z]W���>N�O�]���q������Z�A}K�^�G��w�j7h�9��:MѦo�q�K1�;]����E��G��H����H�ιJ/���������,��NH��]�դ��o��M!@`�6ߐ�CD��Q`˽�3�B^6�π�̄��'(�ͅ���239�0�-/r~C�"���٫T�x����l���A�����'�?���>����2�ص���:�zBn1l��ê��H[��Ь��E#��u�5�BaN*�R_4��W��zl�����ܵ�C���H�og�+:뭑x��$=�\�I��C8l�˨�6�?�;K6��G�`��" �,u�ŀ�x?h&qqB y�8u��L�����X)!����&�&\��q▲�{�6�Z�'PqzUzԮ�~%բ/L�nY�i:��+�X윽K��d�Z�bI8�	����Q`�~���E�!�ME�ޜ#��m��WȖ^���t���j��<4fu.��dz�e�7)�H����]��Fv�ecѝT�GE�,�Ed��ZX=+�r�X7su�j@f��g�&��Yi�=5ԟ��I���/W��
*�7	��X�ҢZ5o��9\W�Mڱ348�ly~--�j3R?>4V.�W�����1r'=��Z��yF2�8eX�i�{����n���-�D�<�+B|IO>_@[���1nh�Ag�
V<���uy��ap:ȵ12:Ѭ�o=��yW�L���0�':�L%q�ÕA�c^�������ݹ���� ��Bz �E\�6=�c�	������}�R=W�2�S�^н��[QpIJ�]R-��v��ۄ�>.7TqN۬NS4f��E�A��P�� +�����1w+��}�w��e!���%n��1��s?��c�4P�B�p�wNJ��5Y��b�u�fr&Z$y��k�ژ[w�+�����C��j�%��U�����������*�૱7�G��D*��R��leuXsdZ�-BD'��c=ȝ�Qٚ>XR�C-� �&σ�]�c@�������7�t��l����!5�%e�P���R?C��HP��[ �0� %��p/�����Loml���u�j�f(�hIi���7���v��S�?_�G�������HÍ�S��(�͕�HE�{��=u��d�b0�4�	{�5!��츒�w��K�U���S]�)�2�j�M:��+�Y�Sc;�O�`���Lϳ:.�02��-p�P�V0
d�f%�x)+(~�Z("���v����*X9犗���0Ip�����['�s���1#<�����#u�����R_s��Ln19�weXkK�ٙ��-�\�s�]��wV>�B�<��)jurBy�~���ϵ���_5�juy.BHW*?Î�?��fھ�[�3iccp�w`o��P�� /�>�Ι��c��=f�7/ �r��Sq��sA��W����A���{)0��,p>�,��<;�6p���s3ND�%yb�.%���nYhS'~<۔f˨YC�u��g�xp�Riý��	��?Nmw��;C̅%Fi�V?~�ԍ�.;Ӑ1�?��#� n��ɥ�߱U���=�H��z�P��;�^����0�����\��-+6 o6u\�?�{�߬����ц�V��`�8�=|њ�R ?�ɂ
t_x_l��}���zi�_�!����|�JǴ��z`��(�eL��S���^࿭W~�[Ey���Q��2�l��&�a���c�H��ßG��)n����^g��sO�=�2��^ւ��̧
ɏo�s����<��֞��[���?D�)��(�Э!��F�ə|ܰ���Ȣ*Q�&�J9>	4�͎ ���wk����6&�6s��t���,���_E�|���`���E�t�]�g�o�+�-�����dC3hG��Q���eK�9��"�t�ku��*�����7A	oT�k��9R��#��R�P�zF�d����]�h�nz�����#~N�	_1FX�dr�����a$Riǧ�����dA�P��|�N��B�:��@.�N�l��x�<ß��@���b;/K���I
����!-N_]��3%mi�.�C�pǨ������Un��)�N^`�|~�XV��95�����J?�}:�)9$h�B���N�HK��BU��tfp�)c,���˥�r��`s�Ber.E��^h�@�f�1�T����l���l9M��dq�ַ���PiE�P�zRl+l[��b¯��D7'�i@�q[�@W����e5T�V>[��e�/-������^_��Vf����dA�<�Җ�W޶!þ0W_&AA�?
8�g�j��c�hp׆��`M��s��FdL�Z�x%&���l�~(�UOg�ھ:,u0T^Ѣ���=~Z�Ŏ�Ck�LH�a���d�5��U��@���uGUX�G��]�
��kzެ�ԏ]+�`��6�����"&��I��?���p=&o����=��k��ƾ����=3ХML��܍�TDx?�d�\a���V_}N����n#���2��I�Nw0Vbz�r�c�Q�]�VB�嬗�5�ix�K����ٹȂ	�fi|.n[��U��=��_֟�0V9*LyF �?�2�����O�)u�������O\�:�f�sp�(���`��������T`5h��fˢ��>�������*���Ġ	\Oܶ.�G��ܪ��
~W�,��;���㰹r�L�d�����8�"K�L`�0���=��Irv�g2�C�'6���ً��Vs p�	d���n�6e�˚wd.us�h�jy�壜Ɗ�='ƷC��7 ��x�:�Q��H� MǏx�U%4��)M�-5�9�E�u�f��y��>m%�
���R���t������F��5j ��Ȉ-a7��;b�2�0���n�������������%�wH6�SW�!0J��'״���"�C���&
t?�Y��2.�/-��m������>>�4���+�G�	v�ض��$��ǖ����A�m����J/��>��O2�0�i�i�z���z	\�u��kos�-�F�wxn΍Q|t	�bV�u���}�۸�J�5�a�Ϗ.6�܏��j~m��/���$ؽ� �]Z����O!�Mc�W�3s]c��m�_��*_�关إ�;�DǄ�𰒤C�ԫ���dQ��#�,	ڨ:2����_�m\<���n��+Z�ۚ+�ɡ%��������B�k�4Bu��goB��CPсU�s�I�D�k����'[4c�����PpA4��,��&K̕��v�K�F̖aQ*�]
��:[���">�m������fDCF�qqZBvo_�k���[��Ҡ�pS��pU`�,��X�r�5�i�&	��P���Z���HDȷI���d�]���A��a� ���Ӊ��[�/�ѐ�q��R^A��H�=��z�A�m��)�>��s �������0Dd�l���O���Vt�FM�O���M�����H\R�a��m�G����&ߔ�w?��w[�Kq�;N���@,�>�B��BM=�ݫ���q6X�rv)ęh}���y V�t�ya[��P_�t#mo�^b�$�G(��|��c*�:�=�W�;[��^��P�Vz��C��(�Jvg��L07T"��{|6"`��
�W�vK�Ĝ?�>�չAm�i��%:&!�Ր��<�@ �tBfWbm��"��g]��3O��?��x	9f;O���'7zM�>��a��Ǥo|�`�5Rw��x��0�:���5�w��<�1�Eܾ��Jq�r	�����~Ս%�A���,9y�,�ƫl/����M��� L��I��`�X��k�D�m�<I�rm.�h�6�u�"�|@ːq��;�c�?<�p^����e�N�7\	�h����FY�X�&~���	Nԉ�tx�  n�ߒS�e�#;�g+��*Qb��zm�{h�L�u�"'U�a�i:Uz~�����mb�g����$tD���fv�D�u$�+(�.Z�L�T�5.�s�O����7!��JlXg�R��a�9��S��X P�mbԷ9���J�[��I���b�T�Jco��t.�R�ZJݝnn��[�>lw8wN��~}>�%�&��g��I�b��n%�z��G'�v��wN�p4og��9��ԓa�	��_g����:�cK'n��>㛨�_�.������}��3��"H�?����+xNM^�íx�,��y����c�P� iDWk4`����S)�+c�%sA�2豽��e�_�C��ʆ!cY��%�?^+-Wj�{l]@���+(J��Gv�2o"�iϜrR��^T�ץu���������	�!��~�_��f>9Xɱ����\K^Q܍�>pˇ�
u��h��)Q���bp�i*0�=����"��5���ѡH�:�e읋zJ��}W�}ge uTGF��>2u��y����*�%:�w���a��7V����Y?�k��p%��-(Q�}�ڕ�4�sN��rf��laVH� �1�rL��G�����ж��v�+����T���uG������V�ľ +�J:V������vi������q_��c�W�E��$g�}��ŏs�=y�3wc���nvI(�~ ]_�F�R�Ͻ�K�m��������a˫�-U1Y�X\�q|�"g�����C@8�/ɽ\��Yx��E����x�\�%�7�pI>o�A?�M!J��p|D)L����W�E2:�k	�����D�a�h{<�m(1����h�(i�U�Y�OS��-dO[礒,�
odr��P�,Tp������(W��C���/��y;?���&9�Q
y��g��|
�E[;�v`i-��h=��x3�$\4v#��!D'�1��n)��	������i��B�+r��c]e�#�>c>�B(�o���Z�_�x<*B ��bA�G	�b���O�h�0V�+XǪ��õ�m����A|R�p��W|k����_ٖ�o��[0�̭�kz����X���U�h��;Ŭ`��1Y<��k<mXA���ɅU�����k^wo�5���:�_%^���Si�� �S^��S�i<r
I����B�,n���|���v��*�Ti�i!��\��l�}�6m�(��$��΂����p�`A֭ੳDGX�4�7����f��Y�h�93� ��q[�$X��!7�J0�Zwzl������'Pb�I,F[�џ�CH��h���(kO�Ykt1���9��3C,H/��!�PFZ�ujv���M� ��V�&Kk/����ǚRJ�(�&\���$�ք�޼N�Qbڅ`ihMԈ��r����^�j�,��wH�>R<Č�X��QC�?<c�o$��Å鵷Ų؅�b���p����n���Rn�	?�pb�v�ka��ݎ���(��?� Z��]�y�N�}�A���x"u�;�(��c�U�8�q�&A�+�T#�+!�RO[H�T��My��Uɚ)�*�8��eV�b]�&*���\:���F�����J��F��k,��ՋKj$L�%���<P�YK�� ��|�����fL�oA�y�gT��!}�B��ni5�@�{$��L��M���鬋���_���S��
�˗c��I�$��q8���6�Գ�4XHg��WZG�(fy��E����i�n/����-���qH8���4��\�1��e�O�#FW}�E���4��~?�ET��x5�R,�3YMK^��5�N8�(q�0��a	��N�\��~(����3s��Y����#5F��������9�.�Ml$R� M��4v��t�|����w�|���Բ���[A˥���@h�l�v�:x��5���}v��3oT��S,�1.�/�L2�e.�r��A��] '�L�:�.v��/YDl̷�ū0�>�����E̤Ɯ.��SfS���� �Re�"�T��uH ��������rC���i���hR���a~��?�]��geV02�sT���F�Y��}]�g5c�6rG�0N�)E��pq�&��7xE�c��_�Y�x8�X�髏1ku�S��{�pX�NM���Z�f�����|�v!.��'��7YT4�������iI�g�SMMA��k�7@��6�2ݭ_�E���Ӆ�)S�'���U���n�hUkV�<�'���.�w�4�-t�8½m��y����o$ow���Ux���sY��E���1yu�_*�0��8ULT[�~|������0*6�k@���CBκ=�	m�܏]�*l��;��mPV�q_������_s����<�QYZ�;�x�>�M�$���}��+s�&>�B$ޙp�P�9'G���z�]�c��,E��9 3����8I�d�W�t�iqa´)c.;�j����M*ӏ�M�߇�ƽ ��yR[�B�IZM��xJ}�.!`�?i�.���6Jso���v�(���hW�>!�/3��o?r�2+���欪uPtV�̛�2��ק�O{
�d��[Y�+�������('k�w�ն�vC���~�+a� +R��.�� s�l\��ı��=5��]A���_���zC$��V4�؇̮��W<��X��8�v������*�aK��HVۂ3D=Z{�95� ������v��B��F1�רb��Hܜ��p�aw
Hbp8'O7Z�'P7P���`��(�F��v*�Ә�TL�#�+2�q��+F�
WK�����o�;r��䇉��G4��?�u�4�+��ӹՍ.��P�Q()}V+d��@U`a�S)�$U�
���t��(:*�x{X�����=���3i-p�z�z��4��z����D�6h�d�>�������loZ��T�;���'�XR����`WƓ�{�����x��]5'`����^v�tW����N1���L�.��گ�V��.)�~�)F iï�N5	��I�����EZ���߱w�f�͞}9�Ls�_����p�gu:�T��1�
[@��}�42��Ơ�z�����ݘڑ�{��U �U�{O	��r+�1���
�c�ߴk����u��n��4�y��pcAL�{�����O�F�D����H��-s��H��!�O�y�G�:�ћ�1:�GQ�p���mGeX0���~��}'[�R.�i��#
���1x������"f �0Xu���$�i��k�#ڬOˮ��>�4����aaf�4� ��A������z���hJ��G�q����&�5-7Eލ���V8�_D�+Ux���@*z�ՋG4=k;&B@#��l����z�����	@�
T��5o��@���.�����xX4-�������W^�PGHA��T��q�I{��^$�A�Z&;g=�%�͋.`��u���I;�_U⥲���*��T��6��F���k�Y��{��x�)V]6m��C�0��_�N�Fz!�A�'ZE��'�`�����~����L{�SU��J��P|zۛ�{v3��±��_�|��?���=�|2/hC1-*84M�YV�.9ӕ�/Xy��Hf@&�>�0Yr�UjΑ�Q#���uG� �eB�iP۾/J����D�V1�Z�Gq�К� �)�������f�?�;���A}	h�a�S�w������9�z�-��/��=|l�f��������|$㨟�����7�eBc͓�����ӎ��~����� $c�x�Z��"2����R��'�9��X�c����\r��,�t7��4^�ûu�|\������6�\��01Gy�/�G�:��	�d&�"��+�5�ue/L���)��Nku�!ɞ��X��]>��B'_j��Y��X<����Jn�ÁB3f�e�4߭Ѣ�8��8�):<5-�<�բ�m��x��l[��:�N�����gU�f��0K �#�ǎ�M����`��zJ��q��IX��$4lPQz�"�qBO���kگ�	�U9���0Ӎ�*r�Kզ�$V�tGJ:N����曊$���S�k�:�,j��`�/�n?p���U>�ҙak��=�4�YB���nv��w� �@���F$]���!uo�,�Z�
2�IQ�)!C�<�!��֜J�Yde�dyn�"ɔ�V?�vq6��`ЄQ������� �HK��7g�=8�6����v1o�b��B�hym��P�ڐ9]�u��s.%�/��ѭi-�JK������2�|���וC����b�j%ν.H\R������~�H��3�[N��0FPM��z���}�  4���uh��ҶӍ5lb]��w^�G�(����4kTX�R��Zziod�q���Q ��Duh�~_�ɉ�`X��sp۴����5�[�7㶀]��i���)�܅ZNK�r/�RP���H�[��^�pؚ-�rd������
*
Lk�ԃ��=g����С~�VL	��v��* VYq�LL�Q�M�`Y���ԥ&M��H�3+�أ~�V,�ms���{$!h�73��e�B�3����9IKL	(s�'xq���=���Xά�{^�t .R��0>�'w��; �����I��QV���v8zz%
�=۷��u|�hw.�t�[�X�5������ѐ�J���S�Koo�(3R	��KF�TI�4���l��;��d�j��͈=��4T�&�!M��_?��I��f>r�wh��^	3�F�{�ν�y���@ΐp �CM�������`*�t��:{py��	�KK�^�j���˙&�.��Q���ܤ��8����r�i��Q�Pr�M���i�~�e��|���W,�a,$�ٙ�u�R�T�j��U�Q^�-p����6���9�3�g�E�𘫨��ewTo�g9:�v$�81��a��2��i#'��o߻��y򹭔��W�7��W�����)�*�G:�7�1�]�B�R��L8#S�~aT@��:�_.(`I\�+wC����R�Ө�ʒ�+��P.�����݌e��Gcj�d6zN�\S�S�I��lu��� I�duҪ�[�D���s��e@ΓJ���F��̯�a���?�'G.��F1xoQ�}�gܓd������ ����'�ˣN�c9�$ԭ�(�J��=_��1�&g�}o6�z��?N�^���i�軹��;/v�m�,���6���������Yr���a�Т�C�-ǻ��;y�L�a-(ɪ��Cc~z�E�(�i���\Üahd8J�%�W�Q��Cp�Z3�K+�$9a1��s�W1dJ�f�j}�v ~�[�kzl�0���C%��5l+9�����}�I���)��"M�ɴX�kA^��B\��Ss� f�5'�P�d^=����Ko?
��+�M�Ƶ�UW�ˠ7,
lƅ�#��H:�c�0g9.ƽ�Z��-��Q.N ezG��R8{q�v���8(��&�P,��B�{�x���}cf������hhi�-�x��`<c7�8��hԆ��L����X�f��6�nɟ��s0)���m��)���_v�U@����2�M��n�����R,�j�c}�b�e���R��J_������D�}0���Bp��p�ނ&;԰%�'3@�m9�zCa�:�I����!ʥ5��o-ef,�A1��7��� �gdR�����	��b�N�UXj�|�܏+1��VK��v�h[-������"�J(ֲw
�J���+�-$U%5&*����r>;���������}�>y�=k�
>����Z�e�K�l��������x��բ�x�tQ�������W�ݳ�4��$��"*���U��}s)�~J"�iz~�����b�8�}�C�ߕyi���l'�~p7�(ݥ����JQ�mρ=�)�T��y��'rwI��L�S���hZqN�����*9?�!e�5�C�7�R�(/v��h֝�4�B���&�q��Ǔ���;=w�o���ߩC��X�Py��N�D�Z�}EA��a���^ח>���R�*��h�G�F2	�e�q>)�`Z�5+�p,\�w�dʤ�kj���>���:�G[#���ղ=Һ+:��m�S�%Y���u4���͋����y)�6R[h���X�J5��� 0L4d�p%6��ї^
�L�T����Q#O
��7	v���W�0�d
ǫJ��T5�ZG6.;������<�L�;Thҡr��?
?�o�ZȜp�9B��HN�&�,_�m(b�i<<mI�@ �`���٣!��o�R���(+�Y���eb6�z���&P���bK�!�Y�Sn���K���Dc�=m|���0{��VR۝�J=��m���H�O=�ױ�	|�n)��n8���$�d4�B������ P��9U�N��ς��&f
��sXw�?�B��&��S
�'}��.�H$�܇b[���+ol�K$�@�k#�"�yf�3�=��j3n�Б�7��1��m�䝩R�~|�W��������	�4�����ֶ�����9�<H%���E���`� �ӏ���1ZӁ�K�@H'�.�kN�om`��_�@9�{�UH�ɝ�bB�=�U�NI`�S�]��n���|yy����L����Q��o�gH�63��os��;	�hy�0!�\���l~`y�?]���NZ�!����xq��G�$h�ܢ�q���ptн?�ۆ ���"S�a���`mt��\�N%�Jѳ7y�׵�V��������eT�C3\|ရ�]�Mf����u$��E��UZm�qi��o�V&4ɜ��'����b>�!��vG̙�A+��(�0����:����Zh��<���*0)ѝ��I�en���YjO0�<R_n��;��&:J�|��ϮW�M����?���3ݜ,��J��"+Q�9�y�Z]A���#�pz
R�4>�Z� tC�ʰ�L�p�zD��֒�=4���_��ƗѺj{!Ȑ�YY��V_Qh�����=+?���n�)J��Rw]/���uk��^�x[�ƚ�b�HY����7�s��3@+�
��é�����/$#�n_��$����̺�Ѝy�p�����"�~�s�U���7=c��|�V�g��ˏ[���tΨ�\��&���ː�x���)���r0�5����; '�Y;)^2�����=oB,BGI���眄�*�)'9؈�h�ѿ��&v�����vL"��:����I�c��B���4)�I�2��<fݴn� a��~���ҵ{G�E�vr�F�^NQ�mUh|�^�q��eeao��̻��?}�k���g���{4����'O�y?he�7ی���UUɞ�~��bF2Z^t�t
�"�h�J����K� η��5�7�N)���CR�.9�f���<�^?�";�7^Z\�����1���M!�8q����3�O�>vL����K�����i�rJ;�5���IC�<aZ*�X�&6;���5����J�V�I�~ZK�� \�0��ؑ�qG�MVbO�j{[p�X��˃��L��H�'�_�Y�y|���sv�ԟk��b���{�����n<�yٺ W=��/��3�uB�Џ����u�E|m��wP߃M�V�iJ�]z7��,��>O��r��gR�l-8���${���?�+�j'o�z3?��1����J*=���I�������]��L�;�u�f�}aĭ��ce_��#�Ó�xx�2��I���}8h�U<p>�B0[�k^��u@��g�K:�%�M��Tb�V��`y˜dɹ$��R!\��"[$a�A��WM�\��Q�|�~N��h`2SoIm&Ӣ6=�?[6W�e��14#G��/�^T���H�!~�_!���f�
��7��yQ�H�iW�5't���	�@�g���A/�d�,܇�|'�� �"��w����˻��Vdy��~�ג�5�D��.�E��@W�S��?;�XF��u�mT7û�4�/������K2�]�X���!�>d�p�$ѳ"9L1�ӂ�Ӵ&�����f��Mj�P��`�L�[�s��-TrQ!��Ok�
�3�6^Z�#.X���>J$�DױgbOV�y�����˨ND?�h{��:�
�"��2^���ʆ64O[�uĸC�	��)��,�x�!fDT�YFB�m��t������J����d'�څU�=._0���I�꽧�s�b���Ă�L�����xj�+�ud�'2kt��K���E	�n��6�_�?��;,v.3��,ff�g��+_�x9P{t��}&ؚ&B�ֽ�Sż^���:
�W�i�#���[���L
R~>�\?�9��Z��dU&>-`�����;&�8w;^�&Ue[��|�g3����?��kk/�
��i�h�6 �k����<�B��A�*�($�����TY����jH1�#L�ǹ/>���S����?߯#�SZ�v��LL/�J3J(��
�O�;Ùk����J�V!s^�����k#-$6���5�y�����9��Rx��q��tG��βZg�W�Kv��cѹ�Ǯb�CA;�xH��V�~����I�������ṏ[ �����BjQ�3iN�2��DDmc� U
{+���p�j����HWF��������V����{��O�m�ގ���I��h��䠎d�~�'���~���4�e��FJR��p1+����|i������ v�l�<|�����̽�qU������΄��KѼ���Sl���睘���Ԉ��i����	iKK�YT<����ҕ�[49p�cm;l�(��sdV
Kd����KqB�u9�����'�{ei�Mc���E�t��rtA�o���b�	�=�_/-����0'ղD3hH�x{e�t�Xl�R9<l����16���&�ͼF`w�b"�|��v���O��j�ey���S�}����O�`�,��g�Т����!�u� �����`6��;8Ķ�խ�6�4��	������{�Q��5��0ު�E_T�g|�E5V��n��_!:a"�.�jSt�b�Lwm�m=7�;�oE�몫[�Ay��6G���F"� ?#Z�(�� �}��q�l#
����&���c���fPJ����Yy{�O���T�?�7���d=����b�iB|�!6��oN<<�l)���ƈ��J��nj���]5��3��է߄!�� ׮�u9��Ο�Im�}��F��VN!^(����bM!����������Ig%�s�v��;Ӵ^#�[���S�]�r\��������zt�b�l�7d�b����I1��.(�p�]QE?9>��&���uP���پ��׍��Ϲ�7{z|�p�8�&I���w�,�g�?��O����fN����t�ք��a�_j�s<Z��b�[XBy:-��L���Kc��wJJ�%��Uts��[N�F�7�>׹����WP��)T�s���)�9n�ڶ<K�>|��q|��Mv2F0� �+"IM�,��ɲ2��VBX"1+�̷c����j�OL���:a�����7>�gs����x��`�ҳi�V��Pךڂ ��Cs2�Zs�4�ࢺ� }K���Hbm�(Li�g��E�-EgL_��qJH�WTbh�k��o���5{!�#5>�Ԉ>��Q���tsj��tw�	e��R&ȇ<'�7�+�h}��p�-ȟ������x���] Jt�������|,�i%1`�&���c�k�H�1,��0�.��~֢�N!��BmA)AA�����u�s��"���Ȝ���{����bsD�G�Ӗ����&��ST�f.:�dO���������@�q1�lx���+�?ϐ;�2o�H�1@���d=*�V�-���n��{��L0II؟)r3�@Yi%pQ��>m��c	�8�ݐ�nC�'��8�"�����+�	l<z��x���;�y�	�����#���'�0��;����a�%[�� [Q�Dp:7Μr�����\8���+�S#˄ �:�&���\�#jr��%���_�"w�Z�-��Y��������"�sH�!���$d�i��0��h��8y4c��x$��us/�M�K��kӭ啘{��0�r�[?��V�C�Ƨ��*�OVJ�Ŀȋd���.�3���_�W��z��
.���k�I��~x��R�q2��V�F�nsF5/;S~��Q���H@\�F�g����
�fD&\���j0��Z54��|��ε>��9=ppl�����H!!|{����v��Kw{�'�]X�;�kr��?���Z(؊����-�q�f�̣V���ȵ�b�6�$)A��"�1��}�J�\���8����7�=WKo��@)���9�p��W��
G�?~٤f���;���|,����s�O�:44�T7�C���]@Ƃ߉��f~�2�t1�4��!���!�Q=ɎE{p�ĭ�y�N�����`�� �f��_f{�yT���M}Ї��"	�L&lü!o�j]�r�Nq��Z��R��`�7��� .�2l{�|��f�MmbkC��C�"E�~J��0��-�G���\�i�_��d�{��ܣ�+b�T��6�O(�'5h��(��q;+-��e��~�\r}�h¼r�%B��bq�ʻO��$/Y�+F����4�cŴɣbZ��	�Ge��i����_��%߻�tP�χ�������qJ��N���S��V�]���?$��"��{߆$C|$�ъ��f��mO G)Yw0y���R�l�tH�p���[��\�D�YS���*>��N_�J�$u1<y)���i
�&j������0}��f�؝��#�W�Ȩ]��d��/?��%��9�O��蟛�}�9�~!�r.$W �ѩ;����/��q�5Q��m�_a߬��9w)I�<�Ձ��~�.*ޗ;��f�I91�A�O����l �&͝6Y����(��p���(s��
����t��Y��>�]�N�f�ty� ��U�%˃�L���*ʬ�DPj�Dj;>5}��WN�9"Rv�p$0S�vE�2�cs}o�3$�Α�����e�U�a|͂���
�)�I��M�����3̈́n�[U4����;���,c Ir=~�{�B��:'�el��at��Eq���9�`M�mwM}'�7Q4$306�a}DH��P����O�<As���>	��l(УQ�����G㜐��oV��r�]K^��1�<�r?���m���(�~��,C�7��8}�<{6��%�d���e������)ƒ��9�B�T�_�2�4�Y~U����/��t_J#׹=��y��4���l���������vn_��T�V�?Dz�tT�6��������5p���˷��A��`X���LLh��}��S�iҍ4E%s>R�b�I;����ס�T�[�M�G	
�lL�s�Ȝ���� ��5�_��z�3x�����W�?�+�6�|e4*�p������T����²�T��]�QҔ���@��s�bcV#:Yx!#�=��N"=�.�-{�E�Il!J���x�{yݶi�s���ی���]+-�'a�A�1L�g���$-��Hʇ�Y
��@�9�
�P��|cR���.$ lһȹ'��N�<Ճmo�n��Z4w��Ö�2��Ϳ7"�!��rd��v� �9_�_os�s�1=;��A7 �.��⿾��6gb�G@�<]?�o/��d��O��|��
B���`�iG�6Z�rʻ�~&-)����F41K?��
�4�*"���6�w����Jl�7l�����iG��5H�q�� �Yx��w�c�؆�h�!mhdB �Go5�A���j�����G�1/ۆ�pvHFW a3��:1�!��E��vD�=ڟ\,5OF�'4E�1��h�X��6N<X��֪S ���}H{O>���j�<'�DwH�e�e��O��#4� ���k�[$�����V�$ѝ�7�-6Ph[s��t�a^��q�Z*+Mo�#�b3�?��֒����K���z�<�����g�~_�."����?�@�S%�-��Y0���v�f��}ޙgul��/R��B�t����o�nP�����spF�?��ʠ��	X�^r�J#��f�6ߊ�l�߂�I~�O���k��<O��Ѯ<�ӈm)�پ�v��<��
����-ֶ�:�r_�����v6�U�v0?8$��^��iһ�m
ۢ����=���L����?���uW� V��{+��SW������ �(p*�q�&*zU�2���n���"�k�)�}Si�pC�Fh���N�Hu|L���}PC�2o�6����w�qbq��lҪv7��}E��<;���x�,+�	C�Y.V�tsJ+�Q�5]�~�p^�������IE(Pq�����ts|P\�o d���j5A��!C[ѻ/��"ZIU�M�9�0X5����v������_�[q��w4A\��f���=����XՂ��3j�D�#E�����'��]������>`������=�d�<�J��0�&Oy�m�{2 �X�.EJ3j#_��>@s���H{S�ď�ɉ�����=N���Q�R5Ё�U������kv�=3�c�F�z�bv/U)����`_ʗ�g�i�%n��+���r.��S�&V���`{����B	oEWO���� �;��E9���Ux��`��8TH� �V�$�U�����a�v;���M���D�[:����C����6 ��}���"�W9�ߝ�kpC+kfj����,��$�/3���I	�󥅵���t��>�1D�ŷr�ݧ`�����/�[����u�?��)��z`M�ÉA�c6��>`h1����W���.!]�b��>z݀{��D_�RQ�ݰ)
�W�������8�5�6��@��s�|y�3)܌yy�X������鱅�5�y�;�&��"�ҘX\� {�/�ccY������_��E���)�88L���;S����E����CV��ȒL��뺉HJI����	�ִ�zhtl���?Q�%[�'l�2�	knT���?��%����k��ǝ��2vO�b�Oޜ5s�X���v�S���,�"���+p��X���?6��8=2�'�qc|l�-bU����U������k�>��Ik��\nK7�F�+畫
������?�q�7ú;���1L ��;�/%ϊ'{)�eYH̽:P�Gv_#��1��g��_�'v���t4b���X�c�&:Gl%Hߴ��E6>�dv%F
�#���q��;M����XAvh�L�T������~��.��b)�v�����ZԲA���I�fV^�R��҉C����<1L�6S����G4�b��)x������H0��l���|v:��)I6�&� _���I�e��/�7�@L]�������������	<���������a^��?�Ah2_p@�������9�B>��*FL��CCU$��B�+mSR|4�!��LU%.����<H�����N��2� i�'JTѯ�χV��U�� ;�矀{M�e��uτ�i!c~p�UIe(G��� � y�;��ʨ<Tꝭ-ͭٟf A�C�����Q��~��۪��+��_H�+0{Gt�c<��N��o�!��"FH"Q:�)�Z\�5��%8�~l/�O�u���]/�3c����K��g�P�w���ɻ8��Ɨ��5���N���szݖ�����B��A�!b/����v[�u}�Q��ز�!���T�VRR��>�{e2�!�@�&\e� ��z����^ɜ���Z,�5bY�Vf7?��6nU����,S�\��b�.X�=)9�t�7�R<��7��C<b��"c!ҳ�3�=�_E�S����t��Ԭ,���g�t��\L|�KS�|ҵ�wN8E�����[���������i�0o��p����'�(�Ͷ����Y>�U_���9����RGܧ�Xeէ)����>/�Y�*皣4��C�\�)�"�&��8� ʅ�=鍽�$>���w�4'
�H�>���ә�$��gG�Ir��
�H��vվ��$U�ɗ�B��Pʟ?�)�*�R�a�X3&f���f��2�4o��	VVN��TϮ�����g�i��9� �h:�{����}�fA��4	?[�G�H=�Qr���)��Ө�������+M�M��ZBpQl��&Tu-�4�B�Cde8�;���T���ƟU �!r���:�_)��?&��t��j��
Q:�T�� ���8/�ΘG��jr�ǚ�u
�}C�jj����.{����b��m3Q���o7�Y�Q�G��- �����9cq>����D��;+'���]-��`H%g�h�{�K��D蟳87�����ț�f?mX(F�5�V��0���u$+��q�"���e��E�є�Z8g������Y��D AuF>��-�;l���(~q0�TQ�ƌ��=94ơ"������E��	&q�I�L`_�zbqެV�X���ak�/�4�܏,^�h3*��L���G�6@	�x[w;�p��r��׮�;��o����c�('dh��8}�ӿ�"vɦ�9�vr��>��
��cg���� �zf��1�޷_>7���'wZ��j�*򙗽8�h�+o/�M����V׷v�TԫP��-@��@w���~1����)&H!y�>�*羊ל��ċ�I�&����r�n�������AC-�h�U�)S [dV3t�3a��k������~Du]� bT,�[�跅j8�x�<D��l5��;�T*�A�M��bS�.vt�7�Yyt�c��Ox�Wayġ��,I�ECT{�+(3���elCmyF�u�PƄK��Դ��+s@q��������r1��$9-�����/Nh]��h��˵^�l�L@F�����9�QB>�X%;U9M`a���f�C�v��@��^�Z��!�N#d�Tɏ����>Lw=ݔ)w�E����zaUw?<g��B6cr����K�'@���PK��[�g���eo������c����|�&�����j��5��-�ոQa�c�~��R�H����j1Y#$�����/ʴG�����vO(�s|���;�cܣ��IN<{+���L,CO��/E���N�g�N�П�w^�;��J������yQ�OM����T��A[��]��'sX��R���E�^}���Wx�T��:�Ln�!�\��4jf�##��^OD��O:n���w�r�mz��E~ZJ�?X�w��F���%II�_��'b{��|������NLvHDa��mǩr��B$b|�O��p=s��O8��2���u�H�d��g�n��%���p����D����l��$�Щ8���}�Dl�!�N�ɑJ;�V���ƨD/7�UZ�A�U��/�����-'!��1�Kl�X�\��):݈�ȒdP5�k^S��:)/��{�X�۩��+T{�l�#�|YB��=���m�!��/�S'?�V":2ɏ���2	J����L��J:9�ƃ;���ͧtPu�ް�w�0a8�Q���92�*3��HC�.v޴	�]�{�D�&61F�fa:D��2-
XRD!7��7BqX� �|x�h���̹<����7�`�4ЏHq�R�"-�E5G��O�L0����>y�P�GA�;Ռ�=���-���G5mq��"wK��ދ��I��r���P��H�?�S%)�nz�����aS��GIPP�+�[�u��; SЋ47�l3;�k���������q�נ*N�3X��Dl�:� `]���+����o)���r������;APy��V$L?��KC�g�۽:�7��'��7H�{e���o���i`ԉ�����������s����8C�Y�L�-',:	M���I�-��-��e)f����4ܜ�s��Ǿ�:x}��Q���9}qLp�|�2r��Y~1��d�
��ʑ(hZ٧�{	ͪ~�-�`#M��%����/ԑ��q8 w~"^�.��/�\,�  H���ˮ��g-���u�V>Kl��`�Vg	�_Oz�l.�i��cH���)bԖ�O0���.���PA�r��qȊ[��#N�9�QJ��N��0��UW�,��u�6te�6+�L\P�(S���`�f��ȶ�k�~Z�������~y@�\ Ċ(K����M�?V�[�C��Ӝ�BG����aN���e+���E�@� �lB�C "P~���z�M�`��E͉T�:�J��Zx%�>�ǥ�H6y\�ƣ�z�s ꛌ�9<�Y��� �"c�'-8o�8�΋�������Q�7�����PUO-�	x�a͍4������2�B�x6Uz��u$/������"A��J:ݰs��Oʡ�3�J	����z`��KyP�]���+���sG�G��_�@��L���6������(���RU�
i���ȝ	z:���"��Q��.[+�Y{��8M��^��l8E�h3��<ȶ7͐�X�k�E�;�]3y�&����Hlq���H��;���=:t|���:c�H#�)8m�,��?r|a`�QaŽ���1��?��nu�9@Hn�)Br�O=��b�$� &��h�o��.z��˒���9�~C�s^,󇀐���Xv�R��gKm1S&�^��0�c�ʻ>��U��7h~Ɲ�I��5q�賋<W	Y�}�1�ɩ�aM؛��N����q����t9����%����ɰ_k�"|X�UQ���1|Y��[�⦭�Vh�4�a.�2^ns�_4�TS"���	qf!VC��l���K��-���}��թC�"=���i@Z����$m�ui%�m�j�yF��r,��1����=`sY�M.S:O@��B[�X�ڰ��pF�l̘rh�W��P���m%����G$�p�췄�}������:��5�����9�I�dE�^!Y�`>�[)�͇j���b����z[��>��r�Mm6#"/���a0R\�*��{m	��eS�LO8sS�nU�u_�$9�M��a^��e�K>oK_������+��L,���\��[�ԍ̨�� V�#j�zͫQ��on��A�J�;?.tt�I$��ːp��I,�����i�/.X���(��x���nL}_=Z<ܪ���8(Xc���J͇�I}6U`��&�CɟP�/*����D
���SP�k���j������j_Ï�L�Q��4����x]�i\}�&6�	W���a���ҥ5�o!���ۀ��PU"�O�,�Zׂ�w���� �h��j�3m�B��Zde��wbi����.��G|x�2�̼-p���9�(J�9�D<����M� 02Sgֲ=����
C�l����VLd�i��30�D!�i�0�O��I.e���U��ఫ��F���B�ud!�A��Vd�l�9�_���p]�h>A�G�g������w�e~\�&� �igvN=%���G�c>�5�;�����W�L�{GOC��q-� u����)�z1��駳9z^L�ggp?^�c�Φ�;�a:7Hs�.a��>�Po�5�/�mh��`U@Up�7���n&��`뭰D~�q?k��cpZc*ኴh�1ױ�e�
@][�:����6���Jz�`%6�u}�����}������G3�k/w�q/2 =N@ �-S��	6r�����o=�md���Y����VwI�Q�i ���I��%�Z4?�H����#��iK5"B'�����r�m��k�f����pݍ�7kD����+��UhHkr���g��pk<��9��CI��Ra�c���3�{/����"ās�����~�ǣ����mj4��|����{���R���J�����~�ڐJX�@��',A݄���X;�j�3fS�qH@��^g.�����0(�4ܓ�U�p$��?P��:�)|� �3Lz��
�af���"����:��I7J�|�;�>a�{����,��� 5O�ZKm��פrɂ)?Ĕ�17/�))�,��ct�s�N�q�(mZ���ѫ*�O�\���i�##4B����_(���Fd��ܟ�C;�i])4�Șs�(�Jχ��}��Irp���w?��$��d��q'����]�����&(��ev�pKpJ>���(�C~`.�� ��C*m���������J����'�|B�Q�)�i1Z�����Oj3i[���cƹ�����
���C�ȳ�^~2���^1n��&�y��p ��7��ǉ�'�_+���jH��A�z�`j�URH�NV����$��'��/C����@���u��G��y��o)	aSU�811���=�S_�>�PzX"�ax�K�-i-5[{|	��R��_:���:�i�����1:nR���<�7�r�oP�ZnW� ʩ}>u���ǀ�)�����G^+�?������������𹿗zx]��:/��q�, �}�ۜגTD��H�Vٯ���p]1H����5>�˛�A�h��*����Z���S}==h� 9�jB��K-� X�oO)���Y�B� �w���3��L\���ذP{��<,��ɦ:� �w	Eޠ@0�jXAS���������$�.��0��Ak�v"8D���y�,�~�⿦�4�X����ǳ�3��#�� q7��ʓ#\�����_�3g���\��LI��ssԘ�(?�#@߁�7J�x�����c�8�&x�?����%Mv����h�3'XBp �H�~�!k	�u���*X�|^�u�����v�ᠮ#��_ӥ����	���*P��A7����p�DE��I�6��A)���gM�533N���_t��q)>
�% �	�3q3��_c��ԭ*vV�� ������"�r~R4��YrZ���s�	�%qDm�*&��߅,� �Q %��
=��~�4�$ғ��?�ȸ�����u֑�#��'��N�F����Iv�����D����'�SD�+�*�.��U�C��$�k����&��v;� ���\v(��|("�87�/U�_�*��;@�BqO!�����e�$�+���+1���}�+�QO����XUL6}]׼n���[���O�����:t�GB6zA[���1�ny|��O�-����܉<���!��DM21y�ԉ���#�L�7��~ϝ
�BG�Z(��>�.��ɢ8y�ER��x���i����v0�w������1�ŧd7�i���z�фd��EL/���$1��Y����%�k�V-=�h�B��U��gє�#X{��.����� .f��b�eU�E�;�o��?q��9���Y�������c��*�te�m��{��a�GeP�Xt$M���*��mli��Z7i�	q4Fs��Y����a����q�L����-���ف�
v���gt�(��m� ,[�☿�\_;2�{R�ي9FfW�MM���jO��15T�'��w�):��BkL�=3$ݏ��ű�5�O�&"V*�$��xYD�u�)�iMgO�"��`)>I�v6P^�5|YJ]���e�?%S�Vz��nQ��_p�FiL�M����в�}�se��oٱ�k��\�!�F5Vy<�:�C��י��*P�M����u
��taQ{�V+A��l�|�R�]Z1Z@�=�+���= T.�bN
)��zd���*z�%��"��fI򥯪��4��ċ�?�_W��+������bf�&�A�e��:�˳���,��?�)-o�Ȧ
HƁX����r�ֽ�)�暺LN�1ll��o 2^e[�u�����;��x������qL!l�b<��J��n�©C]���A{%n��te��h�`#�P�H!��O����z�̣����/yc��	�������i�Kѿu�-�B�����"�����~(f�/�^�ۄ`�P�)��}��]t�p��-����y�.%���>3%�b��$Q
�_������j5���G?�U����Ư�|?��q}[��{I���R�x���8�xs��]��Q�Y-XRM��&��y�����f�[�&���gf��r�2���B}hG\R{By談�MT��y� ���ͱ]��+#��dݯ9��4ܾ未j��أ�,M����ۻw��؟�0�GΤ��eE��o��6sȀ���ɲ�*M�P8�*͕uY���j��=�V�j�p���M��[��]�=�Ekז\��4�h�3����	�EG�r���;.��*KS'G՞�|Z�o-�,�����>Fmv<�Op��`,�X �1���S�^�xf��2�h��U۽�q�F���f�������T{b�#�vU�
O}��[X�*�U[�x�6��p��[z#��g&�Q �6Y	����c[o���E��?�9X$�:�P@�^�:����[��躬H�CF�&�����E(+k*+�4�4G��s-���	�%�c��{���@�g�y�E�V{ݧ]�W���bVb��P<�UD`�qexqRM��
[5�ݔ�Ӳ�����~�e�ۤ? ���2��)6_6*'	���ڬ*��T+e; �	r�l�=�mb��K����9 N��8��_�t�F %�QS�Su��^Pq=;���Pܨ���toe[r?J�[o��A+IzY~�x�I���L~���v�
���^L�MY*
x)l�gą��#hUd�܉/�g�ۤ["���:Eo�P[1�HM�C�D���p��`E�~�MG(�I�~	�Rм��;g���i;���/ؔ2���,5�a(��qY�_n�G�3'��Wo|�E�K�-�TX	���e'���)+��o6��CK��g|	�SG�I����B���Ao'B�:뉘�-���~%���"�>'j7��C��*]k�؊ �����~?E4�`�&Q��[*,w���@�����m�:�m_�z'L� �sm��7C83"k
#���#cwu<E�p?�;0��G����@h(�5ߐ���Z���ބ�v�����G����'�a	,� RC��Ic����i�v�О������J�� g�"�1�ˇ�x����Lq&UP�Ň'+��^��T�eb�uCܼ�����E�i W4֭W}�y�ǐ~��S��6�&�6�I���T?��R�dH���>S���J��yF��o�g{�L���N2��������Bu��V2��|܃�0ՠr�4�)$쒚0����MAW
� �4�)�:�z�ó�XWF��D�O��]i!j,!OD����	X��,��Dz8#�����͉C��;1<v���^7�i&�W��6Ke�G䍹D������"b�÷7Ǝ8�������]�4��F�I��	��i|͸��:�s���4����kP��:�e��΃�E?�]5��$S��L�	D��<����0ۡ�qj�l�4'1\kU=Ud}g�In������G�R��^����^)��n�7)�s�B����9\&	U����}��V��}ٽ�2CC�Y5.h�i�-W�����9��(�͡JsH�o�de':
�#�.~f���v�
�c�s�ù�W��
����bSiO��5�u�lH�5�,W��L���h�QA����)�+j�1�f����D�1P���=
G��~��SV���`�dVKOE�����;'�h�\�Y�"Y��]���pRf��VL+����j0n�ƹ�DQ[I$�WQ��`�����utV�G�{���K�zCj�nX+���A�K�mE�j�n�X��%�-\���d�������E��f�Bw�%~`~�V|�w_�^%�_���t���l0ǔ*��R���#L�U�q1�oNR������'��=��U$~�Y�5�~'�ʫ��dx��<�����#�������s�vӖ%�;>��T#��{�D��ߖQ�Ot ����||	�T�S��g�#e�_����V���z�m��ޕ5C���\�{KU)%��H3��J4*}��ٴ���,���pU�e�CP�H�Y��6��q����|Ȋ�ᱍ[���Z/]�)�����j�۶{�ό
sT���m�������W��i(L�%kn�:�.���D��dA-y{ܔo�X����=��Q�*��$�����,4^�Za�d��8Xb}�m+|Bt�O[��!@d����8����V�v(Dٶ����]}�%�X\*]���A6JhL��)�;+rf/v�C���lD�ɕ�����_�n��Y�۾���&.����y��u�Ե�1B�#Z���P�s�D���VU4m݉t���0:��Pb�,�}Ҁ�ku<�JJ�[������0I���}��N�Lp���-ɱC�]K5�?f�6��­}�q�9��,7mN��!�6%���$~�?��1�#�)�S4wڅgܳ�h�Z����Ʋ�j��(l[������wfB�7��:��x	v��S��L�b�ce".���G���+��`|_��@�y��������#��g��uB�Jm�u��H׿�c�z����!Ci���-�c��_������֡�^�n�2� �4��S*�Q`�s�'� ��������n�+�Ih������#K��W�����5x�FY�INXڂ���lIg�������%�����������i��Ï���"�aJQ4���������q�c���7P�A~�ur��3SH���8V*)���'H�r9�L���ٰ�Ӫ��xf��j�����~Di�1s�取��������=^O,֔^� �2h�"�d�`�p�륗�A�&����bYQ�C��� �&�d�I��r�͖'Q���I�ѱ���U�'����#�_��9-!(&��Ak��[�e+� d�^,�O�e��sv�pԫ�2�,���S���d'�R��r���\�~�:wo5��^w���j�tZ*�b�h@��o��u+docO >�~�.��/-W32�6��E��TM�ۿ#P��g<�'�8�b�� ��v쬹.(�����&��ƵV��:2��5{�6�f���I����$����$jXO_ew 8=�
%���w =�Zȥ�*#� �z��M�,�d��I�$K֡X�\Ju�۽v��A0ch��&��֔/��Jpd�4t�y�R%�R~#��Q�u��w���n�h��Ǚ�y�1Ǻ�v�m�>�.���	4��hG�3+�E��uT^�!{Ѭ�P1ft�ivڡP�пn���̗�R�X~��#^G�Д�.��?��c�ԅ?t�f�
[G�snW8���������!�;���\���0chĖe
r:�m����G�3P�L��ޢ�8�n��bio�qE=3�5��z�.�i�\�Nqş¤�L\O����]Şp}\NA`Yª���[V��?�o�?.�. ��0�"��� ��꟩q�
�H�h1�E�S��2�}<�|y�*���m�r�� �ݥ6/�RG�&*�XqK�֕�9��C@s����k��n���J��!�VY��\�ò�X�I�f�T��4��ҷ1T��3X[KCR`kNc�.��k\ϩ�xS�'�>����IF�'	��B�l7wLqx댕&�ZmvJ=g �@o\0ȝq4��c�8B�ƕ?P��P�fV�U��pLD"��Tf̫z�SbETN�Pz �� ���5\ޟtԸո��;xA�����
_�Z��=+]��o?��{�C���xY���kC4��j��q�б/{��ſ��!�?	��5A���fJ��ƨ �j�S|	�ǭ<�-j�~��`���!u�V8i�Z��5�,-����<M`tR!��v�L���͈�	��=)X̦�k{s��B�.i;G��H�sSn%G����I��'�!ǣlʩ52�T������Z� 7:g�J�(z�ˬ�h4�;�N�x�%Qy=�W����+��2�̊K���}��h��K&)8�L�x�hCdl`Ĺ�q��Ym�A�f���5J��9�? �/�N(�M=����$n J)Lfޝzt
�����.`Z�M��i��[-�J6��;P=�����wB8Xi���'�ZF�+��6a%����Q'��M�����M,E��0܏�����-��-+a:��<��X*�|Yq*åB����X���V��^�rc��X�lTɄ�`Os/� ��҄Q(�������<�1>8�n�Ѝ���7���o.PT�7&��萏��ɋ�{�g]�t���Q��Q����H�ejض�;ц�S����>9���;�w��(�|�Ը`|[8l�K�>�JS�b	'���уF�ħ*��5q�ep���7�h4׼�4[?�R��ls2�!�#�.8.b��10�wl��:���Bd������͞ѐƸs�o-�h���P����L�ɂ��lW�/����|	�F7������p�Y�J��/�T�����2�d�1��OO �w���0�������lV߯��~IgB���O�ߧ�@��A�����p1ym~�*Ԭ��AD;Y���;E��D�r ��P3�z��ҏ��{ۗ�T�*5t�௿m�/*�+!t�L�^��3��������0�"y�&�b�M�Q:?�ۛ�����h�J�Nv�6\1�y���� �� [���9�H����-6�Q�5U
jIOd��>�i^HI�;g*�ZH��9Kĥ�ޓΚ��-<v�m��?�L�,Rr���x���õ��z�|��~鷘��mYn���=/�QUr|�N���zl.!�4�������RH�7�w���]��o�	]b0f.պ3�����\��s�-Y��NB��l��?��ɺ!�ϋ<��5�SR��<��K�1�dGx�qf��-ՠ�a�ݿ��sҙ�Fa��3D	KA����%�E;�r(2�sm	Q���:W��O&X7��W2�.H�m�Cv[?�e�ră��:ck��т��&�G�FY�eS>5���U��?w@w,�v��6L��u�Xfv>��K�������Pe����ԹX����L�A�O3�̐�Gu�ЎX�Яm �`l��]��붅 �E�.��J0��fU'��q�J\���������w�)�����z����̶	�go�7��:"��:��7��Jr�b"�$��E�آ	r��Q�U�,�औ��:㤾�v-[�a�m/�[�+]����t}�E��:�v�R���V����X��|��%4C ꅭ&!�B�
'�Z#	!�7D����ds�f���8�J� F��vKg�����g�f9�RR�l�>��ggU�j���D%h�
���0P�o��U:�yx]6��Qf`nl��[�#�%�I�Ӑ����RN���C�ǒt*�?��ߚ6{0Vʾ�
�^<�"����a����(�A]屵2�.;�3���3�[���O�^��3���RtR���u�b"g����i�����-	�AO�x��[�?�� U��*z���C�9�R����<&T^/mӾ�.��N�|hՀ��siM,�Q��ߺ�gz��������*�+��X-����ʊ�T�^�P�I�I���:pe8'p�	��gB��T�YS)��3K��T��3󷲪o;��ݍ�#%jt�_ilOg+G�X�1ן�L��*�Ƣx4{=���d���|\��b7������^����=�E o-�U�B�HM�c �o<����p��7�_ݧa|��W���g�6���C�"w�%4�ۃ�1��]�؋["����0w=����A�n(.���_1�u�S�f��Ɯ� 2�W��bR�����E���������e7�����)�:_�m�E��9�vc��X�d:�WM��Z�Ey(��fxMR�O�k����fL#��vu�Gh?["�O�@��Ԩ����/�#��S��|}8�i�B�*�p|���E�[@�G(��E�mЄ���&�c�:��!�/T����6�8�J1\��8�b�܁���poQ��������	���`@�pH���Zig�2s҂m �C��;�`i�G��qD4���)O��rn^3�㪣�޼�Z/���ea�lW>��/*qo����\�L
��#��.䗀�Q/
�1�"�@B�*T$zf�)1�u��c�|�q��tg�*Ϩr^�����ْ5�!��^�b<��j�)�����iM^�l�o�sR� ����E����v�hN�|d&Ŗ`�orh���>�7R�����>v��(�%"X�q�h������b��kz�!j���j��~_������22�7EZ��A�)ϫ�^���q�9/��emN��o�vZ8�s���u��!U`����7^b�:nTV`\�t(pӱ��ĳ�M��	I��������n;�����,c%zRFq�ѳ���� �J�ςg��(��<�t��`�A� �C,a����hm�"#�3�y��A�b)�8Q�o��l�:u=�X�M��_7R��94�<��u�VD2r";���r��%��ZX�*����\�!�,#�y��I=�1.j�~�c�6�{���ƒmwÿى�z.�bV���
"�T�1���'	
���L��K��?IK��DdgLs�ߊ�<��?�5jZ:-"���r��
MYK�9"k�׉g|kl�4����L�2�^��֫�D=�8�N��U����Y�������h���.]4��8Le���O�4T�1�� TZn�:a:�zC�"�[��A�Nh�� �K�	hƸYZ4}�B�2� ���L*<Io|o	�2GM����nS3R9��X�ŉkLR�aq�����t����se�4�p+q2��w^Au�M�����ㄙBr>�?�2����fwv�	B��\C�m��b�j/�����^�k�ga5��\E�ð�l�<���Cg�C�������=Pi֤������[�{��w�?���7y5�)֪
W���0	:L&�ƅh�Ev��EJ<����Ci�z$��c��� ��X��Z ��\�p�)T����uk�����+�."|JX���ŏ��W�}4�V5�����dg�ë��w`G�@h6� ��>�czGi�OҲdNvqҠ�	0�qZ$�:[�����xut�7U�M�������!�zN�M\���-j�_G��+��0�5i7s֛�fb#�1%&G�k�;CT&��MƓ�����b��1��f1�9��%ٕ�o�+>v����C��k��N��5\J���f�Fk�-�kK�*i��mlw2�Le��X�46&%޷�#B(G���4�S�lE;�YON��Ý�{%�����f;�o���\R�Ĭv	"ہ&f$�s{X|̈́D<g�����Lh"ᢻ�s�m�<Ǌ�x�90�`�ڲ�̕>����=L'�P��ْV���((|�K�iw�E�WC=��]꾨�'&�s�+��L�QF�$gj*��;��̩�UOؗ"m|��|c#�W|	v�P�;+��
o����ʧ�����ZS��-![uR����݃C}�f���)����l`-�F�ͪq�i�ֈيo��ˮ�����a����
^	=����I�u�o]��'����K���c���ׯ�g�jỤW�ey;�D���	�"����!����[����j\����\�'���X���Jv�q:�m~�����)��K��f"pҸ�����A@�/$N�&�u1=�h�<{㘆7UMl���Ս��g�i�>�_�/<��zē�Ca��"ݮ_>��C5�!|^��o�!�!6j��~Z����b���'�Z�%8+a�C�0�3��(P'g�(eE���S�&���f�4��O$�u�ǿ��U�	��.��A|���I�V�`k2.ڟ�.�%8s����6[�V��S�݊2��Hkw����^}��.31���{�!�ǂ�B���� C�!�_4��`T���pS8�H�b�x��qf�N&a��c5ܕ�sPeUR�v�����Est[�X�C���y�^�
a/p�Ts9fTkf�]R�Y2�_���S�ʍ�w�QX��g�	���9�C����i݋��N/���*�xQ.�l2
�LPt^��q1����M�����m/&��s_nL-��7;J��p���'���y���M�d�3�D%I�����7�U�}�6�2��P�,��ʋ
.]8|����[���,P���25�Sz���e�.�����5�﷾I�z�X&���e5/�K��u�]�P�ѥ��
��x�F�R�6 ����D�Xm*��B��M+��%��DÏl��}Md�Cp�#
�^M�K�,h1\<r�t#F˃4�l��m�Z|��SǴpx���R�n����0ѷ��܄?ȐE:�e8����x�]p|�c��ƛ�o��qBHl!�7��H�B�д��5v�JY�������э�� *����t��+O�a��n�	��so0�m�I���:F��鵥��x��1;8ߕk�*�wYo�͌4���^�!3����[��-׀��"��Uz��z��.�?��Ò~�KZ�!��Y	��ER3=����i!��~4���|�����6_}퇩*��Y�g
a��O�Q��j7���IA�Nռ�P ��	C2�w����2k({փ�c*���g/���C��oTw�O���nT����f3�\�>K�������0t ��l�s�7�hL��L��/��zzM���y~��������ꡨEѡ�o��ET+�W2�c�<Es���f'!�~:~�&�3��Ļ�tgL�	9z�{���[a�%"�/�*`�R=b�{ʄM{���DNm�j���ug;�gJ�*_��>C&��sn�L>��w��X�������1-�E��"�d����vO;p�L'
�9g�n�`���E��1*2�ths�珿�Kh��Ȁ!� :jw,���(\Nꣻ�2R9�����nSuR��p
?�x�n28X��f�z�`&Jr�aR|��KE�:�x?M����=�4|pՂa���f
��K�<�=�P �L�y
�"����q��fkF�́��I��Lݘ	dd#@rٷHho4����$; ��'�q�Ɨ�V���8����Z�8N�p4�4Sخӟ�$	3��U��>����"u,މ���s��شR��]���/
бbw�ܧ�x�Z��㎢=����=��
�iA�Xy_P?�a��C�����M �U��p�dn ����� �j��C��('-��z,x��a2�!���������(L8�t��k�dDb�Ql�)�RVy@M�y�������]�AF���c�b�	�-�Q'69c<�;�&�a�[\�T���sE���&��x���Z����T�;��#��"�IeH9v�I0>*���.�{f�_
-e��I�ه���W�ۥcƒ�S�����*��Oc��T@7�pJa�;�v�`海��5���pi3���b����f;�|��g�$�����`��N�xH�!�m��Q��O�
�a�&Z�*_l6<h�1�u�Sڷǚܒ�g
Ȣ�$��Y����f�C��X��Ի&K����61&�8ld�T�����:?&�b҇��ha��iD �WӋ�9O?�i��+m
/h�������RjY��x�c檯�捀�܏i1�{w�&	�aJL.���j����(��(?���+ۯn��� ��H�[���#i-�^���_�'=ͪ�JvqO�蘻JP�߯MY��iiDQk%+��=ck忢�׭ހ��Q�w^%������k�"E�};l �d4��	;�sAj)��M拰*�@#m�GR�Ԡ�p�2L���[�n� YS��H��t]���XQ�h�6��x�m�&Ù|v�Ae�3����6��M�Ӊ7^��P��/Yd��S��1�f)DD'���>u'�T���:���t���#��Y�<�S�5�j�$�!�Y�yF�O1K�;��Q8�*�c�L�ȯ��Տ�J�G��Ɛ����ӂ���1Q0�]�����D�R�i���j'�������b��l��ь���s�6�f.�R�]�`B]��/��C�tEW���{���<�ՠ00F�ncov�tQ=���g�A'�'��ѝ:�����_b��[�>����򯏒/����%�
`��q���9kc��&��6�����k+m¡	���o�NM��w�[�w���.j����ۿ��_kPmd�@6��
Y-��4� �+��p��=��/o7�s����L������Sg������B�m�JM�89���/�˜��#gi��U8 {׎��sܦ�����K�5�;�>��.�؀băa��=?�(�A��/ C���fo���3�T��oO��ŷ�Q���rDE!|�Xs �_�{��%O����4��o�1�5����9�
�SĀ���a���J�QhÍ |���k1�44��',j%�;U[W*M�wn���*t��Һ�꺚�?Me�;}�ü��D �}$�p5��U�gr���ٰ�bZ�϶�(NWy�w�f<�ĭf#3mJLt�L��H�?-V��.q.�䷍|7���C�F@�U
����Z�]�]rHh@9pj�~��YD�����<={�&&�RD�:�k7nt[t��l�G�Uo�0N�%�%���J��$��t�j��hM.-yY�q�&7�l�YYt�>%'�R�D�e��-��t����~��|/��=�Q��A�Y����P�1ަMmC+�*���,{9;¦�b�x�!�U�JO�����N���NJ�:�SV��ɕO���4�" dH�`.)HUZp��cc�D��X/r��O��L���)��h_��:	�j�gyW��H�LxU��Z�����6<�C!������YK�����Z!)-0s}���(0e5�SD���c�^[����:?MiA 7Zz�����vt�=�g#Q��0�6(hTV���x��b�ޱ7̼f��N��s?��B����g�����6�6��[[{����h��V�����*0���Vj��_%��}�$b�
�ƜG��~�����Vf>)��#��u�⻭UL��̂<Yz:��εMz	��*�,�y�Q�_��GEns6i&m��HW��JZ��V�X[�;��-���먔.�ނ�A)^��粯����,�[u�٨��.��`�eV��&�m]��d��/UJ�X
��y�-~�|ܝ!Ԓ�te�
�^�_I��|�'W�w�~ieS����Xpi�21	)��r����i�,�.?��^Rr~_��>��}��	�BYc~M�O^\ 7��Yp�7�ܽ���%�tAZh�fPy0(�#�4uyq
}<�&7��^�SZ��C���M[��N�4%�!fP�W��U���d %���'�H�ki��jQ�993I�^��2�*u��Y�9�;�Q\��k0k�xc�fVDc�DS��^�5=0��C84Ҋ�0���k�����ɜ������9Zv�{WkD=��	C���<���}]j���)bm�A��d&���S5=yW��e-�v(&����
:-[:�0�Q����w*%}�[��N
5˂}l`�Q<\��_��v�M�5�Rt�S�d�gH	E~܃��W�RJ-o�9��]~�7z!?�+��z��Yz#�#�o�h�6)(��uK�%��à;9����{�tB4��XP��V]�l��LC�z�@���^�>ډ�6�� <���;�Ū�5(˕����Vm�U� rܠ@r����U~��hI�̑,���f����xr�>�]A�v\�
S�]��v]?��)�w�ո�V��rm������`UC��ׇ��͑��N�i��#X-��^c�j�r�	dy��9e.j�����jg���a@<}����HC^�c�1a7���S��;K��rl~1��$/��G��̊��G��~zzg~�����~maF���<,���ɥd=����7�~3jF+��q���	&�É�����\1Y�����@X�`��l;�d��}S`u��o4�d�I��z�.JLs�bfExg�]�`7+:�F�`+u��6�����F���
�W�������IL�_�a���,���[����[i�� ���x1g��a�m<��79�ݵ8s��h�"0g2� ���yσ��t��2
^�x���"��M;$�X�����}����H��JzгP�%��U���ދދ�X�CF��?�ѻ)"�����=��A՛M*%Ϻ��	u�V|>R������a����&� "���
|r��Y�Z���Y����V[)&���Ee�S�5��6�tul�X�R��|��V�N�`&c���*�
u1�$�WH%�*�&�~����r�HF$�۴��8J|�f��	b�Wcr<�
�s�4� *��t(�l���q�����?����zz��Ke�����(�0�9�ɵ!������\e�w�2����˹�:ԝy@�%��Q��&��,�?WB�}'�д���Б��(U+!P�@]����yi""��˽w$��:���.V��Q��*�����z/>w�Ё4� jt��s��GrH��)����!ט\8rRs��=���V�l��J���.�?M�ˣN��_+A@f���0�o���jΞ��]0���RC�A�9)Aٻ���^Xv�BW՟T��d������7H�o��>Y�S��U�@�PL����´E������D�@3=a�:�b���/֖mP�O��!J�?K��b=~��`�q�sY��|=������5cK\�ϙ'M;���Q�gdy�>O��O�<_�ѥ�G��D�~�ړ9tbar�j����#�p-}��:U�k�e�\����n��0���H��WbJ!������jf�/��#�[H�����Q��e\��{
`k��$i�;�F��b�������5�/���1�G����O�2����6L�Xg�疝�����JU�N�j/h9>�܇-ķ,�z E�+�R[3g�OC	zE�HĚ5�������^���|6��o3lQ��=GngY&���#{`K����v�&U���fj/����*鲦�Z�~�O���m���x*T�Z��4����Y�HW���ۦ����P �2l�ab�$�>�=A[xs$ ���Yex���$Jz�O��lp��T��	�[JYZ�fY���<�:X���B^�b$�VG0$�>�$�ٗ]�0d��eg}�ֵ�b	Pa�*�����w�<�n�g7$]��4[!P3��0:��� ��GtU���?+a�d�ʤ�Ã�G�Lw�z����1��� �/︬�WG_�U��G��ғY���_�1 ���Da��uq�`���l��68�#�L[��̀����E?��z�(
BV���H�`�y���� ��Y�c|SѾ�m�!O���C��ېs�+a|W	~]ٸ5ʑ��/D�ɍ��	��m��E\��oq�n;���x��0����SgQJ�3�����M�����P��:�w�eE��6}Ĕ������
�q�A�����'�����G/G�\!�#��m����T�cE�|q�IB(2�َ��k�=2� *&Ot_L����?}K�4��-����Gː�%��L��[�B"5�-�P��3W`7Y�I"q�Oq�g/�e�L�"J�Pz����\��L+�jJq��3c]��i�Z�ۼwBqp�^����^��f�G[(��t�l�X�HT��F��&;���h�RMIll�7M��H��;FU�x��E�,=u����i�H�����pH�����=��cH4h�����ȴKys�R�ZEK@��n�i0�rj� E�>+�4��Iʪ�.|1O+>N��ў)����]�z�+u͒T��B��?���(��g�@�NU�߽�q�ģ+f���_gŹKH�c(��t���.�����%4�̽�*������ıYn5Q��N�@&�&�t�#���޻���{��)�aXܪ4�+��'��ce�qh�*q,W%2��D{�V������&>@��4_L �2�Z�u�c\P�!�^i�ǀ/���O�f|00������D�;���X؞/�H	�t�q���~\�' |�}$��`�C�wA=�&��oJC��Oʬ�,��=�{c!����<|�t�f��3��q�gW6/x�Vt&�!�Q�
@�T_��!�����H}Ҭ��T*�	���T�O�GR��ٜ*�#�`z���Sd�H8a��y��Hd��X����r�����P�T�@�]}t���M>�o��󖷛9��X�������#ƙ�Ai��A b�V�sͱ���
pyCF����\Z�a��X(d-��˜Wz}[��$hܨ5%��#����FU��ܨEe8���9>�#���,�gwLS*�q���ތ�1j��M��4*w�&XYS+X'T!ư��"5�p2/�8h8�b;��G{�v�1dBՃ��A��N��W�o]����Up�����Ap���Zx9�m���S|�2�Ǟ9�JԪ#8�t�'�u�,��`��gI�J�٨���޶H�.{�a8�E����^ep�כ�㕷��~�r���mD�>t�y4��<�;Ǭ���zА8��1�r�����v��� ���k������� �|��U\'+�"^��-����ya����W;{x��e�2���j#�7!:AI��%�N7E�St�M�¥5�K�������쒮G�hq�8%A���FO���#�/M���)66x�b��J1�X��I�GE���D"Zq��0snK�Xc��B�ղ��5�����DXF�痣w
?B��g�>t'�5Ϯe�8w�ਸ�y��z]�� e��#�F��`z�\U��ʸd�����x�p�j�"Bt���s3v{:-�>/*�M�K���:5�e���z���V����=C�Hi� ִU<T�"=(�V��1�C'����L��V�D�r|�ֻ	謉�?�-w?��3���U���.U���� �9�,�棽�����r?�$�8@j�U2,�属�Z׮�:>מ?��J�ģKH5i�Xҹw���W�og*�����ޏdoZŉ�e�꣔J�F��=+.�u�jo�=n�~P(�C7�� ��#a�T�0HAS2���6�%���WM(�M!��8A�yG�ᕴ��a��8��R�g�(R��oa:(^��B|[
e̅� >s壐D���I�HY&0�d�G�����o�����j���m�}	|:��hю�ݙy�6�J�n|��4#��.[W�����F�E����c��R3ߓ�)�4���b49#?9A��Ssq��@��P{�H3V
�^���0�>��Wީi��z��
��ǅ�e��S�'1�b�����2\P	��B�c��o.";0{��t���ܫewc��)H����x*6≃��W��t�j�8�c�gF��}{��b��'Jmj���>1`M�$�J�>�������<�A�t�@,/L�
�V��y�qH�Y��Eo�10�2�@����㻄�xR+�8�����9�p��bʘ�J�Q4cE�������G���֘���Ž�x������bԇ΢1��|�U�����U�d���ٰO�̘x���ma��3$&ķ7	L	ؚ�u�߫g��}�ѥ�a�H����cŞ��m3:&�kX���\���
�#�۸{q�d�ȍ�Jҏ"��k-�V�9�n5{B�LT�7.U�k�A���3#��qtg�|�ێR�(J�W�T�o�w)�(�!��O�|�\Ƽ���Gk���|�5Z�GĮ���^���P�=;Kw����	���E�U2~�N
}�t�^�R����].t�M���{��f�Aֿj���k�,+�0��0��[�Nr5��FkM~��)�FQ�\�g�бrܱYV���u(T;A
�6=Ya[S�'h;�C�CI�}��)��
7i��wU��{��4;T�����3dM����!�w��`��p��㓜���i�}���&�L�������"�\��:Ob����O�>|1�)��*v���q��R����gWh��1�t_L´Y�OĹ1'g��}Yrn�c�����N
�	 ��7��-�}R�_�-��OY�<���c��E�\�	���퀪�wz���K�{.�a����C���(��k௖GׄIr{@�;]�-f`�N$�YP�oK���䝿�Y���6lF��\Q��K���&jؼ��:��C�:��eטj�#���q�@@�5��
k|f�_>�̿]S#J��A�O��� ��_;�12�w4�0���F0�/�����\'���;|��af0�8���nd�9p�y�,��9U+�k���Y���t8�mӷq�{=iA4}���GvI
����������;��Ȇ_��d�x O|��.o�<l��<{�\��bl�u��)��2�_�
�~�Si⒢�g��K�s��N��U� �\$B�Mu���|8�}]QL�%˩�j����T��K.����l�V�`9�*��Fk��4���~R1�*�4�ա�-�%��#��P�H��bD�h}��FZ[�{��ԋ�A��$U������5����Ҫx�+VF�_�\�D|r�
���jRX���+�Ė�^bӂ�
�HJr����}I�c͟��S]���z�n��.��.6�	�ृ���A���p�7�A��U���h��������2*m��A�U��a7� \��72�|�t�׌Q��mb(1��%�
b�e�G�sm�5�J�*�ʐ��w�����#�0���ya�a�JK�)�*�l!B���9�q�&���ߤ)�-`:IK$�(w�1�G�1�Cw���[
���l]���ħ[�Sm�yj�XS	'��#F�Z�B�{݅�)J��c%(���>��ufI$�H-5��e}����?����A�/WV�����_z%��i�N�5ޠ�,�V��g�q���e�<2�1�(�2?6�!J�T��	��n����w�5N4{z�HקVpxȼ:�z��劜�r��R^#�:}(N;�ɜɄ����]n� ��nx�� -{�"rн��,��ɍ�Y�C�C|f��MSџd���W�}��<�����ز��
T��`�]��wr'L�"�(��Έm)�Q��D�����e��� �d�Q,ӭ5xn�KC��]�u'�vLo[��`�Z��^$2c��M�n{Vb�!����1(p�ߙ�7�����f�-H��<����ۻ�OB-�(n��2JF���>��o��b$�����K�`E���Φ�(�p=umL ��w��$"�tX�7�r����ے'
�I��8VI���������N7�=Zppx?O����W�fm�g����zLF�n�k��=
�A��2J��}�}uq�@K�
ԫQ%V(R���,�2��X|J����O,��뚶�N�5���,�s�8�{�[α�ǒ���Ú��*�����?o�}d�M����ek4![����(E�Xۊ 8�9s��C(mpʒ�S�o�{��0TڌIS���^���N�T�W�Π�j���FD7�	<�������&��=�Z���m���n��B��FD�_��,b�j!gAN�#&��]�,��N��E�Y{u�|�c��*K��W�N��Ʉ���M���C	9ɢO�
���ʤ ��)
��k�}��U�u�A�
V2�!=ܹlMt��w8b�����c%��hn�zfe�[������_��%����E-�sllkS��d�����T�FѢ��x7;�$V�S�<>�]^���׹f�wiu�G��b�~?��� �g/MlZ�u�,�
L��tlʔ�D����t)]�FV���V��������NМ�!6נ�7�z��pw�8^#A��DN��U�h.S�S�W���^�S�L*ٺ�`_�%��]o6���9��br7L̒�~T�7�QS;�ټ%5���\[O=�+�����6!�Q�,uƪ]>�Q��o�Wf?@p?�v�-��mק���(���9!�q It����e�Ol��ٿ��@Զ�1fN�h��ϟ��l+G�G�8UH��Vs��F�,�6E��(կt��;T=�T�ڟxr�: A�'����ϑ
F(d��>F~�o��oc<�]�g/�G�����s#5Y����Š�I��D>��w����er�S�%,J���E����|�s{�'����}$�EW���՞�z]��v��\��g��� 2�V6�H�M���zP4`kYE-v ZCj�������(jBH�ED�����3kبbL^��V@6e���0�;V��֡U1��m��Ղ��_�4�a�}��e��#D��\�eJ:��IP���%��t�y��в�����֩S",&�|���R2T!.�:�~v�n٨-	|Y�t���)��;��-���'�� ����k`��5p�w;" ���q�-3�fe��>�9�si����ݥy*��cM���`�괅������5b�d줐�E���p�#m��S�T����YN��Rƚ��<�@�l��4��8��OMӨ�Z.mY�G�v�����<�H�M�[�<�tq]���5���? ]
����F<>r�UBs��۽�r7���!_����t]���O��h&�q":���r;�n���S��8U�%NP�i�����p�k`b&��?��I�E����C��9� =Y��+��8u�:}��.��"����)1��_���-4"ӻh����xU��i�ɾ�g<tQ�!>J�P�=�/!���N_��8��Ozj��*���Q�F!˦������ _"��R��N9.���˻�E��֔��ro���N~�~`�0 M�ԣ�Eo �������JN
�<�-�"{9�;�nG���\�uj�	퇈q$�,)��~s�평�e*j��=��kwR�!��ug<ݺ�����/~e�@ֳ�G�P���QTs0'w�r����'�+�~m�-�jk��]U��A���~k/�Y/���J�[�\~��J��������V�G#�dq T�ɚ:^w�hE��KT���5Wk'�@�#L
�n��ᣆD\Gb�J$���9��i�����Aχ��%a9����)l���X�0�Q�q�ѺZ�ā9�nE�+���Y)Z�.�kL,M�Q^���D�O��|�V��^�!TN��� �*]n,�8[�`T
dR0JTP�V�?플1�ى�ݛ^�XB�|+�at������i�[DA��U��\rY�z�`&�#�u�{G��)���yI�cܴ�.�o�(1�����y.����JH�@��-��`N�I������F��C�6�XiJ�xE��UF~a���r#(�Zم���uj�ٕ�'T5�.�݊�@s�}/w�긍���	B�.<TTd����Zp\񩚊F� �b�	Y-i� �����Sn��(n�Q�Y]�{8��H�x�K/�k�J�C��S�q��%�]�Y���g���9�G�_��#�h��
��� ��bti�Z�_ۨ�1q~%i�."�,�@WM�����\�Z�kΫ��d��j�����L�o�^c�gu�y�+e=�@mQ��#V�ZU��$cuM4Utԃow`�~�i����%�؜�:���}�MR.���Yb3쯯C��zŀ���@7B��2C>�`�T��-��@�B��8�c��ט�a����r@wXS�2蛡�9~"}YN��{�+�{FcR���ꮑ#�� Ћ喿4�LL��D�,�Q~��]x�����0�j4��*���>c��#+3�hp1�"���U8RHI�4t�������O�B?���y$'c(ľ�ձ�FdU�.'3�\��3W>,��B���eV�LtREe�5+hM^�wM��q�l�Q��G��3��ާ[�PܰG2�J6w����ƣ�ԃսi��vGa��)�8#O��g4�$]����L��p��e��_�4�½?J8
��ΨSy��un?c/,��s9����'�4�I/]�Zm9�s�K���P��,�pƑ[��NЀ���;��㭫hD��E��&�!����B���+L�ƓC@���ŋun���5��:�����{�*��}���~��>�2��2A���j����3~e0��2W�'���֍�q��k��Gªh�z����*ப���K�`����C{7�L�fd�����oє��r���'*��a����e�Ѐ�e�t沙���8MTt�0x�tt���S	����kv�L-ֶ�m&�0�z�m���o"mM�̌6��E/���So�tJ��C'�<��L�}rp �8���>V�m1�0J�rs��.��G������k��V}BxQ�,ȁ�Ҋ��:��V$=i��saku�Z,�1�F+�y�3�W��L�j��?܋�uv>�mud��67����bS��Do��#��OW��'P}FqIY2����\Ц��8���)�P��6w�������7Z�Ȍ��Q��'��_�
�7��Wu+�o�[�NM�)7k}����$���\���*�;�;\�W�+�~��
3ώ)���S�L1r���v�_2^�XMíu%O{��O��g��9y�X�7oM��u�ɍt���m�y����Na�&r�/�}6\����:R�$t�b׬�������1W��d  �9}T
�1F]���������)E����,$��剒���4�T���"�$��ߦ��t�G|��=(/2})v ���(�*�Jd��Q̠�=��ŨO�r�}�����] B^N����5�ͫO���h����bY���(V�[�I���h��1��PN����݇Hq���C-1y��D#;���	�|8ʫ�q�`���Ʌ��K����h����J:I�﹘�U�'�<��(�W�5�b�|UW]�X�_`*4R�Ȥ��t�_̃u�	6Z1��hφB}�;�W	$c)�.�������1�!�,�@MIr\Zs`*�{�QGS�@�a#��E*�ʑ~y ����k4	z�**�9���;@�A��%5�Sp��D�^�«���$1i�7d`@���x��UD�܋B�{������>�ǳ������F���B'X�!�re�Wf�x�vug�R7����Z���⥸���Y���)�љDx�����/[��*bTI�T5C<뼗���`�2�?��*�쟌��7�Pn�RD%�X�dq����%�H��t�Α����	 �y���$��Z,��t 3�"� k۶�I���1�9}rZ�%|��	wWmN��H��w{���9��P\l�tF/I=#<(D�E8.��a�3�����D�ݝ�Z~���E�0���Z"¢Fc
f��aR����[�+/!�r��?�����oƫ�����Q��!����@V,��_FL�&��J
A7�����B��b ��f�;V����أCZ�O�F�d�e���pT/U�5C���s���I0�-����ُ`�����ehTAuw^Q�^��r20���hLP�b�6��_�\d:h6�'lYV=V��9��2۴�g��ցYgс�h�U��X���g::�z�ݏ��Z<��r?C�]�$�E�� �xZq�*�1%�]��M��Or���G:Ԟ���a��D6YP&���ּ	��r8L��kf�,8�(�%��*�f� W��֪����ڧ�]W[�L�T�^p�<i�!��Uo���B|���9���1�Y��{ ����܀�߸Z�}���d�_x��щ,����-� Ԧ��|x9j!����.��+��ï��
%X���
�0k�`0�����=H�I�NM����u�R�v�������i0n]�#�u��R��1օx`�G���H�af�7}��+UP�"޽�����Ui����un�ۀ�3m����B�%B|!y�xr��t�k����P�%��Ų�u�;�v����O�����)��8�)��\���Pm���C\ѻ,n��EDV$�J��L�%O �� _�*�!�jjb^�%���uLD�n?{��S�v�B:����#��Z��H29���}��c��a8d2�ӈ�����jHi�B'�8��Iߪ�����L9��W	�0m��耹e(�#0adĘ�n��^��ֶ�7�{�QC]&v�}MnY�L �+���Ə��I�0^,��ox�&�JT������B�zt������. eg��Œ�/�|�_�l�����V�|���Ъ��7"���굒b/<G�AuK������W��N9!���a]��ǜ^�Px1I(�m_��'4_�Q����0���b�X��I���;�YwIn��I�;�_�oJ�P��	������zKO'H/���
&�|�D�bi0ͦ4b�+�ӛ��!x?~�	kg8v'��sx��L;��
��Y2D�ji��n���OQ��F0��l�7�� ��͛�wj=�a_ƺ`�
�l�MtE�����FG�tʾ����!3�gѵ�Th�� �;'c��0:�1�C{j~��7h��S�@���
P��q({H��SBB�����ܪg��<J6����`�n���Jߟ�T��
C�F'�>�4�L�����b�Xk���$K^�����̧[���AviW��� �>��y@\l�U e��I���6@9 ��� ��QK)���F.E蔥�8�\�Iope�\���!^l}
����䑭��n�C1��r>��_b=��[d:$�(� "�	.�hP�P�8�	b�|J?.���=�-]������$.�DG�GV��~���yc9ADh��� �r�fnD��O=c�M�1�ٵ��-5��|
ٕ��O�v�5��I|� 3��n+�}.j*���]�N�?��PjE<9m��Ӌվ��|u���ѧ��ݺG9`œ1�r�G��F ���%��dE��$ICaɈP�����0���x7���ޭQ��wت/���4�]�'T�_K(C&5���%[5��J�@f���L���xf�c�R|3��T2`I��躌�T�
y=ٟ��b0f�.���	Eo�Z|����`P��Fɷ��c��}Ŧ{�]AR����c���]���D�����{,�.��*3��ً�[�Z�����\ ���É��?"����q�Gz�Nu~�S����(�u/�I,%��s:�wl�0O�14H���DK8���X�ԑ�'V�P�$GC;�bj���ѩ�	-�v�85#����SXd����0t���y3���)+�F��`�k���D����f�Lz�
.��$	���_r���>tIT\�`8|9�U<��n����u����~x�����q�x ��*G��q��Q¿*�PJD�x�1���s �Gl�!�������T�+Z�C�h��1��?٦���PA(���Pm�r&�-V�z=�ѸNkx�?"�]\
��9v�\�sRq��.���1�ؿb�g� \tÏq����y0�9�N�Y;��g-aHh�?.�Y�hbE��2͵���y����/�_l���w���$�����!�ɐk���� �2��.ኟ��l	lO�ZO���cY��lsw���f�q7���T���z��*8�\�_J=zv���'�F���;_��#- R�	�4��S�	�Dǰ=S���1Ɏk�3?hl24�v��vO�� :7\���Y�z$�z�e КR_jq����#�7$�~�e~����h�5M7"7��u���x|����9��5;҃��^N&P>sKu�,�ʛNjG��<��u�����m�YȋX�M�#�6���"'�H1V��cQM��5����z&@6���[����Eԓ�k*Iq9G](��J��l�)������WU����UM֠@u�#�Z������3��4<S�M�[
͓�����P^�"'Ƌ���f4M�©�\}Sﳝ(Gk���@Z�َj+��֯#�S���|�凅����E����ˤGSR�/U��d� $��>2#�t�W�����LN�A�ɐiR��H�%v%��/-+鍽���=�ǫKgNUCaL�.Ɣo�SZ�p�Z6o����2I��1� ��8ď5�P�g=���͢���gZ["����E`b:��W>?�y��)�+�+��y�r�8����*��8ZU�>M���{�MO��W�A+�Գ&��bS�~����{n�.����	�9�H��Sc]+B��p������Gy�3`V���1)d7��\�Һ\S�zd�Ye_Щ�k��^(�N�1���0��Q���\��`!���ὼr���i�N��hպ��;�i�� q��c����ޕhwڨ#�5��zƝ��l�v��r�b'E���^ҵ�G�<��X:�ݸ�	4�Q����3�00G��!=X��������K�'՟�r)�Ɣ6��$����[��f��Z %�uR��lۓm?���CI�p����خE�D�n��>�L���7��-ڗ{�T*:�)$�Z�T���lA�
�}o|�ߔ���m��,d|�7p�ק����_Z�<qc�֬�i���<A��ЪF<�8
���p������4�A�rV+0̓����A�Z&p��~v=N�/�����I8z��PfJ�^�~��咵B_Y�r_���#���[;1[w�A$�+�LI��7m��A��X��V�\��g��R�>I�xS[�t�>j6�v5X����Y{LT#��n�Ӗ0��7�O������6v�;���d�җ��4�w�8Z��yI0�*Dv)�Ļ�'g��Pf�T�o����/��9�a0��C*����E�O�,���`;�8I�m���ٖ��T�c�	)iB�/A�ms �#�3SA�Wô�A��]'���[,����9��M�d���}:#�{���f��W�_�Y�#]�E'5�Mv��B%\�t���s�yg�^"Ξ�<�$���9q���l�R�q}�ֶ?k��~���5 �,�a��KIw����0N9��͆�U�=Q�v/D��ɾ�2 
�3�'��z��S(��H����]��3�{�](�I\[o��x�A&D�5�'@P�ܰvK��@%��Gד���g�kGM��eɶ�X9uw��{,�I!.���ݼ�a�a����L��X��v_�Xy+��P[��D���k��U&���B�=�a4l�(�U
r�iJ���V��wq�v<n6�.����#�z�vkd ����-������)���R���a@�9���>�8�`�5�>	��YR�NI����~��<�m��j�.sw*����Ob<�J��j�ct��NWI�Z����%.��SG�`|j�~m)�.j�	)J��������K��L�C����G)��$�
�s�L�U�I�(dL�#9E	��>��Su��~~g�bh��'�nN�N�F�d�0)&�XW��$Ly�-1��nYW���Z֗��J�Ul_��~�>�ZZﯨ��}g���?��$p5}`r4��&�T����0���+j� *�϶�����~��PKѦhX���m��Okǵ�^f�!C�"m�PW����jT���y��e��qX��L�t�*��q�1ۓuݮR���g3Jo���gt
P�sI=�]b��{y�3�{Q��"��d���ۄh��݇������*�|�Whxj�p�s���a�c9�0y�G\&�Y�c1*f���d�(�=4��t�`�K�RB���JÓPc��Z���X�^8H�P�ez��j��tӹ���4�S����Q��Z��P$����1�Ƶo%�V����f'�ωc8�Z�}�>e�~*b���:Ģ�#��ZSvH܊�(��?S�B5���G)A&����U�Ua;��Y]3�����	�q|P��;�+���9̉6S�?;�n2b���Ĉ��.�����H�q�c9R3!�Q5�?�7$5�a��-�ʖ��	r���=��`�/m1�nם<Z�ك�6m��!��(��H�?x��n T�z�(!��M����oM�����+�v�1����F��i�z��T�k�C���6�`�GWlqEwsV�߿	A��~Ɨ�
RG$���%���9E�����a�;�����e�Q^RS�}�����7K�nB��؞J�7?$�&'�Ű����>�謪�����O��d�<�K&l9)Fy:Aʡ~��o��O�'��W��͢���{^ky����$Y��.��e�|���w�f��g\�[����R�Lq��Lp��B��g)�q7ܪGf~���b�B՟R��e\{�ٜ�0�T�����8��ߜ�%+��I&`��㹔�~���@��$���GQ�Dן�F9w��c�3Em���3F?QL��s\����F��Ǆ�fV�]
 "K�K�~9hrqV>ћ�-SP��E�$����<Qo�wϜ�Z�h��S	��#�?��(��/5�wi��ɘ���?�q'Ʌ�w�;C�"�RU��*��z���7x�utq��=��/�K�Eo�%�����'�g �����`�K��	]cd^o&��|��w�H�J3��cU����T;��X�T��P�9�<4�����sWl�@М�������8m/�Mu��c�8=��]&�ϸ͛b�WU����@� �`��ϵS��P�!<�W�|E ���k:,3��A���+�ו��G�U#w��P�';�1�RD�r">����p�.�ym��hp���x�SK�Y࠳���C�N�0o���{���)< ≴��jh�G{���#fqXu<ݠQ��ө�%ϻd&�n.�}d�6��@��Юպ��M�>�~G2E���y9ًE�|��DȐs�C;���K���)�{�&kw��Z0Z�"�}KDI'l΍�'�Q$wZYk����M�������h娐夨$�^�6JL�j��!���\S�f`�1��_�(�|���_����t<w����eq��9��Χ�tbq��Ր��n?���n����ė��A��Q��}Q;�{ro�}�xkyfo9���|�Q�\N6,ڊ�6�j�d���W)�����+�e�Qŉ_�9C`&�YWIK�T������xp�1�C����\7���M��u�@�nq��T����m��Xe!0�5�vtx)���}�c����O�j�U���B�.4L]��^h|�c�G���q����$ M��4Mu,�����U}�)��b�w��<c����AJrU�������^$�z�վ���a-f[;�K�������v����ag�^�����*�R�_f��[��p�%�l*�E�@��S������u�-~O��uɩoy�J�9@��Mo��Ȋ�-��Ol�FT,o;����F)p0F/�Yܒ@I�1�ǯ:��X��V�{�U�(-��> >��Q5)� ��ì��%�Ũ�Y̐�^�"��db�SX����'��{ٽGid|>c��bG\�}���L����s��[� ?6{���),��%s�0��E/�S�U��ӆ��Hڼc0���*X?rl�w,�&�Hb��`,��m���'��҇u$�%�U��>�`�2C��F]i|`ޅ%��4������Q��P'�M�5f�����@P�4'��SMs�`v�(~�y�J��^���z+j�v	d`+ۏ�����q�cڕ�4)hѸ4!�3�ZXh>s�,���Ӻ�l�Ru�ρ�w��>Ϥ����Z۱r�ڋݰ*�)l�3�r�RX�z�*h!!�z��d<e@�J��gӹ���R4�)�(ȩ������T�c��е��Ѧ���u1';V���]6��;t��F���,��pi�M����ס�~z��o����".D�JP�e1}�ߛ�_Ļϣ��+Չ5�f��p�g��ɇ��`���!����5��ѓp�WM*y�&7����"׺vj!��[-b=���XR�����QE@�h-�,��T*�2гu���$I.	�~�%�_x��ĉm�ٖ ��RS�9�����˪����F-�EP�ۇ�܏/	��l+�Z��}�g�obmܷ�:L�[U�����V���G���r��d�'��`�Z�
��m�QF��Bbפ����y��,

��0���Xw������ǌ���-��M����@.����~�2E�i�n��A?��{e:zl:��D�Q�A��'[����{&�8��+|��,���G�˘�_<\��%���Fp�8��_v�T�$r���rN�� �B$T�?�>u]v�^6��5sK�;�X��-̋�AZB����26'��K��E~D�z�v0����`A��+O����X�s]�t�\��׏�?�F���u~mʍQ�Y�z�<r�� �+o����/�����/N�7�eOґ2�y���c
.ل|�����{�֛]ʨxŅ�]b)X��%W�6E�_'_��r&��z����nOK�>` -T��@�y��pTàX��Q1��]÷���Fy�&�r:r�K%���Ќ8����l� ����붺)�2�_%�8��M9:U�?g�.��tʌ\�@İ�K]Y��[&��>�p�$��L�����r�ylsw-bm������>�-��Ĭ=�ҟ��5QvR�x�G���r�>�U�##����R���UA�j��ZփI4D;�"���e����/�-�e2���ޫ�t��!�!~��fVvMjW�b�pD�
�{Lnn��l��Qfl]d��8��Ⱥ\�C�Kj��L߭���p�Ӧ��#����(Q�rJfd#0��(����&������~�B���ތ�zWS.S&��m7T��r ��2�����m����v�lg�ɇ���Ô�٤!�ƒ��@��
Ͻ^���cA��P�MA�>:�4㔺��d)��p��PDbE�8��=М]�oԎW%϶b2x$���0�6�wSi��q΃trz����uY�@*��O��j�}/8j�,�d<��J�4�Gn5�	�G_.��[e����<X�}���K�~�rR�i��)�"�;5g��1XI��33�%`�̩�K�wp/3��W�A�_COa�dl�~�G��9g|:OŠQ6�����<�I�_;7�#^7��#L6$���:#4�C���C�D�*�*ˉ�OzBSP�i���)M��,�ک"K���i����Y�?�˲ĺ�O�]7F�T����AwBIZ�罓�Z��o�m������{�+���9B��J�&��;<E.����c[s��jiL�%���'!�J��lzԞ9zPg'�"��͒?:On���R	}�\Ro�)y�uP��`Z;Y�T}��s#�U%�P:"�/Ǣ{0WC��g0W�[藜�`��'y����C� ��O'R׍�n��o��q�R0,$T.7�<��-b�H-��R 5�e�Y��m��3K�&�2��!���^��S�\b⊸h4�m:Xއ����ͽ����_h�u�f.7
�0�?+�t>����$Aˢ�fy!~S-�l;�?7ҍ^;,��=��2Z��R�w��5a����M,�E�k�ռ>豆o�T�V�C����r>F��e���ӛ �0���S����y�q�M'��ǵ0@+DTE	�� �a̝k#zqօ�P}�-�5���C?ޝ���ss�[2x.�\�$|��~�35�����i�9\;��� ��U]���Ss�HBepmA}������?�����>O��}q0.'�F_�v8�'�����{Ft/í&�vJ>{@\���� ds��@_%R7����\�Ts͊6	����=׉0��1$���`��K�̮��L����aҩhY�	{�����q��ۮ�e�K�mF��̐p#lcXM��M�mՕ���f���]i%zUU�}�m#�������a͟��q*���'��n��E��YE�I�tH��!.\<aKLȾ�R��Y�7��
�3ߞ�Gi�̉M�3u��y���S�0�/(y����_�gg�հcV���}�Rl`12�R�"�}��+���ms��bJԗ��^�ie�um��;�U+"Uj;k�Wn�3w6���,B�
p$A�I��;p�IB�F&����ɺ1�K� ���$OD�Ǥ`����-��K�
�'�ѶLN�T]��|�ER+��)°D�DX��~�(��8������*HY7�ئ)8 V��ӽ���U$��L��a��M���;� �z ٰƯʪ����n���v��5NЋ��Yf�18�|.�ۀ=I䕼.[���^rm��wᰶ���1n���0CCj�F�	�g��S����~��n�)(,�y�N(�>DG������0f/�s���ϸy�����X�P��L]~�j�)���V�?�	���Ǽc������2鵺_�A� l�}�\Vu�=5��BY>���K�g����h���tr�Σ�>�<Jw��zM�g�H-���RT_as��q`T3��~��O���_�n8���V���}�x��J��]���j�|��X���~g�n8��˨{��p3jR��`Ǟ�e��ۙ5�jK�����f?���q�p�G�'�X�-�� �co�-�=>��=���Ao�h�g,7���"��E�i WY>�6A���)����A7�:1_iw�+�O�*��%���ET�?E��}%X~�1��d�z�k�GT�������:uݫ�|v&�bCghv�o�k�����o1�G ת/Pl�ʅbA���|?���C�DpA�B���6���8�m(lI�>����c�L�|�́� ��L�\�������2���N\6�\{��B��@mPӐ<���iB�:9(f�a-ٹo���tV�摪�<��q�6?;���f�!a��;���0( F�׫�\c(Vdg��V�mث)�rq�	@��l9tj���_I�t�%�Ƕ�p���?"����N�C)���KwE�D!k��
�L��4^׃����V�w�]��d���&�@/�(�?g�
|lզ�Wq���G4c��Zp~����S���W��cR�P�<ѹ���q���O�`|�i��c "��P�@k?3O.�%!/Œ�i*^���:ie�;xdz#8�AY��7��Y�-��(�k��]�i��+�D��c��L|��V۫�+�dt%�P8��9J�Xs��F�����S���)t!�%��r��w�hH��J�-��t/t�S����@\�g8mŲ���*�dU�e~�f���'P��TB�_���nA��aq-t�e�YM�V}G����9�:�#`��H���T�+�Ee�¢���6��|
����G�q>�Qk���7Y����4FݬHX*FZ�m>TZ��	8'�~���2���Z���W|��GD���H�XE*�^M��cU���e�#��h��?�� Tթ}�<��,�v5S���lw]ķ2��a;-���uKzv�*�~����|���`D� ��-��;7n��H���Д�&�H��)"�JM7v����s�˾��˕e����fPl��$��XF��i�yL��ma�D�ڟp��]!��:ͅ�R�+.��`#X}�؟L�w�'��	���V�r�;�������#�Ccs�"�ɝ:�S��RjU5�QL\o3؊<8;t����Z$,�ڨ�*>�dT�_ۙi�����5M�A��ZS�Z�/���E��,)F�]s�@�1�(����y~��������tă0#4B�@�k���*>:.�k��E�=t����/c$'� n���NS��lc�M�ZE9h��-�cen���T(oEi҄�G���bsJT!pU̹	޼������m7��s�DK��$��krs>��'���F�
u�y�5QK�������a�+Coa���yW��o;�vJ�R$}�X*�H*�R������1������`��8)�4���,<P�Rpc`S�uA��D�Ӏ�w2s!�~�"	Q7�1�6���-9fn��ۮxh�����������oZ��q��D�e�tݬ6�I��~T�'fa��.#�� Q�����0��)_BuƟ�ɹ(}7y��c�����K]R�j��w)����t���sOMmC��i$�%IEP����#�4��^᭗�	���B�Gg�����M�P����h�jw�<��5#�{��"��d���V�.��+,JY
�.眛��3+̏Փ!x�jС��3do��kV�^��|�1~�<�񨞨�.썓��4~�o�}d@��@�c����Id�[˞��	� �Λ��{�B���_�v �TE!T�m�}��?��'���'�2��m�\_��7ν�'��$��}���-Mѭ�ZO�cuQ�o�,ıZ�T���\Q�B�J��P� �*�GQ7��01�_�G9�:�r��,2�g�k o�~G��� �X�=7���׀^�de Z>���BN
�[TK&�R�j�\I ��1����^FJU�_��O"�X�)����	�!X�U���L���Q3��V�}| �g����'�3��68�]�6z��5$sƳ NKw��^]� �N�ڍ�FV8��`��J��aFX�2"�����{Dj;��f%��m�HL�����*�q���y��̖J� ^s����k\�Q{�m��R =slU�:C���v�ְ�c�	�_�4�������=��	6�hV���x�2	=r��Q
�֢�(�\�*�3W;� �5�lXJ�a��q!��2
_	��H���Ȁ���e��PI��1%�E@����
E��1��vۋ�/�����5�]S~״��w3�K��"��}goE�����-�I��_<�]܄�i���j�&+�w���m��;�"н3�R@�wqO�kVٱ�FZ���(���jM7��R��{uu�
3��ܤM���(���/ ߝ���V��u��B�ꐉ�<aQv�þ��c�Gk��� -��\�7�t���jZ'2�7^}>D�;�5�7n��iTѠ5�0r>7qG`����(h=6�J*F��O�l����r����=i�pL�"� z]�%=����|�z�;+�I�?�NQ��=5J7��)o�E^�����4����I*�nǘ��) �n��^����\�<-�ASc��m��Q̳e
0�yx? "�'\X8Fho��S��b�v�K3f鼽�I����HG@���Z�����A��Ed��rk7���wo��0jn�����]������^0�3C����O,f�Mx�����J�Q����*mX��F�M���v��ϜE�(+�n������O]�d�>�/�l�����$�(�R��`7E��$���0������@u�0����<��~Ǻ`V�;�
!�EX��a���M��+���q�r<�0�h���̞(�-Cj�ET��������@�q6�8`�^y�q�ɚ�Uf�
s	Ta�.��@j��o�J@�(7��6� �x^��eb_�"��G�Q�?��ж�#�����:����!gj��96��o9���`xI�0�V���u#�X���d�d}Zh��Rs�o~>БǦ9��T����=q��]ޖ�4y��-0����%�p�͡}Ȧu�#(��ٱ�}�:�*��x��X\ =ϗ�U�?��"T�`�������W� Zc7 �:�å�E����1�=���G�[KGk�7���5`/�����g�m�
��b6��E6̈��.�#��x��K'�3����4_}�"�#�m+&ޱhGoHmc�K�[�h�{�A�Z�u��D�֫E+)��I�v�K��@F�V�6��)��/�����K^<�x��,�}�H�pK��]K�����N�rI��D�������Hw�a�o�O\E9ެ�˓���xz��3D��46_��!�2S��jR�Z�x�|�⧩o�+�]8�����`�ԡO3��E�=��X8m?w4�x�h갎we�����j��6tRo1���I܄��P�Mq���J0�9`�b�K�ALc#9~N�hӝ���W�`���6�v�-)"��" �$���G��ewǍ){*�7^��C�4[��2ح�t�tm]0}�-9
m~C�ǡьwc�,k2����aU�.���>��p��ԝʡ�HM����?��$Q��ħ�xR�ve��Q�NI����8ۼ�����޶��x���6�<�9��k���㷀$|�5�޺Y�n�%�j�.�*=&",���Y��L�ԟ	���CH�xèr�m�H*5�v���y�b2`'-�J(�^��"Q�����'��xu�?��R>����K|�G�=��R��a�~^�)��x�y <1�zRF>	Z����y��R��<Q����d�P$���E���p��F�2�N)/����0�WNCb�s�Q�[�O����P}����[)�[��:���;V��Z=����6�0���4<���	t�n JwZ�<����엸�m�����c����D$�-��$`�N�5�ѵ|��~!S����1%պ�[��r Ɨf��g$s=�R,G;����<1����ʔ���V��F�B���'�:\׫����\c�M_��@GO�-��wh�z�W�U�L:bgns{4��'�diO-�r$��&��ǲȦ�r�z�s���Ց=�@����p��4�7$D�6�\ˊ:�>�ԅ;ɬ �z�t�!=�:�6{���-'�b����o�u���T�
�����PO�-g<��署�{�C����
��B���WO�}�����ђq��nc_��?/K��Y.H�z��N���,��ꈭ=����K�s&Wg�^U�W�I�`z!�Y0Z��;�R����F�RH���?��Q���e4n��[�|\��Ny[��|xt�6L�"k�lʴ��#M�%4�A���w��y���,#U���@���
$���� �~�,��6�h&��
�o�_�h�����6f�8����HU��Θ
��wCp�"�;��T1���l�o �aP�&H�G�5�uP6F!�on*\��ԫFQ���;W�J� +NA�_]��{���Ǐ�K5b�~8;��e�
jU�6�נ���Jb-*_T�~9�������{�R�=1�1�6<�u�f��!w��I�I(�B�d�� ��w d��ij6�~��h��b���ݠ-w�m�e�9k�����=����G�����|�)Z�| \�傇�<���d�?�f���|�2�EO?K�c2�t��O0϶%E
2˹�pqX��3�h�D��+M�ZS�la�98�9��<a��9��:a�8��;���/�O�Qv��R̿��҆ܛ;c����6B7{F:"5�o�C�浀�Z �'k���-���sh�r<eȷ�N�A$�!]yf�2�����d ��Z��i�r����A�<�B(�ᮗ��P�i�Y8�Q�b����e��]�#�!�&���2��Mc+���@e_��;��[qǶ����7�C�y��)Q#2�[���"�� qT�0A��=��_���ɇ���7��̝���s�����J��)��Y#��8�"o8�u4B���&��Q}��&��8@F�"�����[����C+��
5���4���.�ɐ�1�C[=���l��וn��p�.^��}�R��п������ϙG^���J}�<�@�,��,���h��������o���ur q�v�jJ��E
��&����$�@yKp�����i���QM�5�߸���6&ϋ�����5�� �����R<<�.ڈ
9t�"I�\J8QC~rnH��ȎCZH��YH��w/�'{�^6VΗ|��k[0��gE�!����
�`��2���!�[#�z�_�[H����9+��t$���?X��m,��bp㶹�����*B���F�m�E��o�d���-���<��A9��rˀ7y_q�k��K�p�S���L�ۮ�I��p�\�@n+���>i��Ԇ~��
�c�uBQ��3��J�ݥ�s��Ȧ���م�������+xu��8�׌��$FE)�X�	�+QT���d��
��azغ ��R��W��3���
7�k6��Q�]�5OQ��^�P�c2���²`�J�s_1_���^�qxHCIX��� ��f�OQ��?5�8Us|��"V�����KM�e)�o|;��F}(�V��E˶�8f�q{�a���b�C��0'�1��)ꀓk�.U�.���6��d�&�o�Z50� X�����ӈ��]i�/ar[Q �c���?���Ud%P�A�d`�t���$H�B����C�;�x������'[�yc;hQ���r����̢���)�޺H�u��ǟ�.��mZ��X��B�׫�oTȼ��e]��|jn�;������Ƥ�Y����z^ �o��H�i�H6EB#RT�$�3Z@���xA���D;�Þ��HG�*�H���B�ƺ�:�Cʸ5�}U�������@����K���(� ~}�'�5w\��n��Z�΀Q���l:�^��4�))FP�3�n��M*��;�o�ut�l�V���H�0	�C�G�����َ ���P<�;iۖ���!{3�O1����,�,���>S���FO�}\=�����H�����ʄ��nq�_
��V��U�E��W��Gڥؘ�O'������;�zv� ӰT,G�@��?!�iH�,�����Ռ&�5	��*DX�2�V�hg�]m�|R�Z �|/�++�w3��(5|zR6s�*��h��4ڪ ���&�Li�;7y�b���Vo
��"ͭv����>�=�%���W�����-"�v�6<���F��}����RM����*���U��,���^RPL�{�q$� �jv�K��|$��C��4���xz4b(T�P����H�����nfW��䣲��u�p�)�D�=��-Rt%�IVK�j�^xl�7$�P��	e����*9�v��,�-}��ͦ��}�Gm���o������plz�{��Y���lvk�S�=���,q�Q�h%��2f��.z}h�B��r�m���u��̕w5��Yz��ƕA���ZJ=��q�b�����bz��!t�8�,��!�u��Kb��;5YX,z�O�<__a�-��3
�[?)��p]���b0v���e�,`rC9��	�$nC��F��H�z�d����:YI�d%:�A�q�Ԁݬ�u2����}+�w���r�ǰ
I�gGǑ
�Ŧ&Ws�O*��,����T_��\Jwu��^CZg��5�680x���C�<��MY�.�a�O,:��+�)y
E_�a�e��el;�� ���5��i`0�T�~�A# �Ȉ�Xt
Kfn��f.}Y����ޡm@o	�7�%G3�e	�K1�ͨǲ��_�+b��8m&d�+=��8�sa��Pm��S/��(��j��q?�¨3�ś1��{�:���%T��wĄH[�*�d�lg�=�q���X������EǚWD����%�3�5�?D(�����Bz���h+Fe�n��6!������ݾ��֦�:���H���{*mm�B��h��M �lu����%���YQ�Q܆;<l��$�&��D�>X�>R�/P�zް�P>�k��v�� ��q�~<��S���.�����$�+���#J�.�;����n�h��W���u��ǚBk=|KMب<�v�,��iȁ����x��!D4	�R<��l�y�J��@25���K��LFaTx�*e�ߢ�"�K�r	�58 .`98'��Bq�;�H]�L��f�仞Y����
I��R�=�Y�@
�`��1�����cJ�6V��l����2�$͝?(_��m/]�m�]$���ɠ���aݐ����q��5��-ɯC��ME�(G�QY�b�W��p���,G{5��k͵B� ��L�����ġ�@r�2�dM{�=r�Z��+k�gzH�W�jLu4FNYΙ��	\<����w���>ɒ1���,1�6�i��3������nh]8�,c�V���F^�J�=��Q�w��&�g=�Qaw yU�6]��Iu�Vغ!b����Hku}�����n��}?�dՇ����
xɧ��G�G����,ͬ��g���ڲ�9�}��`6��*�0�,�������%�}]M+�_>O���1A��,GE����l�~���^�n`B�G��·���q11[XC�,E֯i��	'��5���+8>��Z�0�h�*��}|S���;���+|��Ե+�a:?6֫�z ���i����X���`���1�(�����)�rY�4���
�a[������Z� �[{ރ\�y�VA��.-���ilT��W��:d�;):8�1��s$�+���E��j%�{F,!�f9��nf������:�cL���஍3��t� ܐj�(�Y-k�Iz��^�W��)�?��̤Դ���������:0�,8�'kzӿ�L�PQ���F�����`OP��6n��ɍ�t�'�H�,��+���� ��'_d��&Ց��$�ܬ����S
<D쌨,�Y�����?�x;S���8��t������D`!"�}�1\���:�P�ta,�PWB�Q���&�x���VNaè�N�����qG���$�c��.��t+c'a:��}؜�o�r�?Ռ��	�����r*խ��o(O�����G�M3V���2Q��PP��F$�LⱿ%7:u��;�9��,$������9%�v��<ީ�J��q>�os��rrp���CT�Ad�-:
�&�+a@�R����//ּ��=s�����ʗ��i�mm��R�<T}w��+���z���x��T���>	���z�q+{ w)���=H���td���]�H������*tϹ�5�D��j�8�N��F{��W���o�&��d�K߿\��e�wŶ��#^�݊�kw�j�%�唛2�H�sIPW�����$�tD�i��Y�+�"�����j�y�`Ȼ^1���A�H�u�w4]̣̿mĔl����ۭ>/�����_����oՒ��G��Э�Q�أ��&q4ٲ�O��d(gD��x5&@]&�j$tS2ç�e��m��\�*Ŏ�J�%��Z]o�_~���[C\o$
��P�o�%T�`Hu��
e$�]2TO��1��Ǹ�Ҷ����Z�'�I��B�k�uDT�9��Z����kȔ�1��_�|}�H���X!_�U�h)��1z��yH8q�������A�tv�> J�n�F�I�̒3+ٙ;��}����K{�Û�*�qg� b]����:TMO���-Ej�U�~������p0�c���T�V\��fM��v!,\��>E��|���W����E���Vb�䟐��W�b˪iA�������>�j������whyVRm*XX����


/�2� �oQRô��	}Z^8K;�׾���a?��r�� �l�8o�	 ����XbQ �77���wq&�����ȩ���L8���6I"�����<ث�����%���Y��2J�|�D$�F>�
[�k��=��(F�<z��q�d����	l���h2aI�n�f�Xp�Hm�,�q	O��1����3���qA77o�%�y�[�0P�zx���~���A�	�Rw�L׭��N���\�vX_!�/0/3@��;�!�<	7����[���������[q�NЅ�I�<K衾����3q�ҍ0W�QS���؁����,q��P�>*�^���6"d��>=[�S����j�uP����i=�8k"R����v�4���<^����E���<4a#յ�ȄpD��WYT�a,�db�=���s/��^��hh��l����+�6`�@���)v�tl�(���4�|t��+�dSO4����=yA�Խ߄(���>6��6�!m&B�(ߍ�mY �(��ǽ�)�s��Ǩ�X�g�#�eX�=l�� 3�P��]E�<�9���ץ�K.%��VE��D�c-���Wz���<[�ُ I���r�$��(x��L7�J�ux�!���&]j�La����Bҥ���e�et��s����ת��űM!&�ܺ��͓c�4�z�v��*]���א�m��K��R�ߘ|0�Vޢ�a:m�#�Kԫz��gm�����*|�������}��y����hW��	�����y��6
��t'����<�i������xW&0KɁ�D#���-�M[~�����'<KZ����48��Y��g�A>��N/c� N�L�r��N�<GVt�����n��N5&�}��S �PB�-��_�/�7���e�7���yd�����ZA��h��N�~�Kmՠ�l�8L���7�h� �����P��8dccg8e���|Hܿ�ĒU�N{%�Xq� �wz��N��;\�	n�|����ii�qRE��RSѧ8�����}�d��s'f�{�v^���osVv�T�c�]ߞ�;U�YnJ�3�gt)VC�HxF/:Zu��˒iv`�B�H{�B���͝��8D<�@���+9݁�2��U|-	EJ2L��Ak����g>�qM�2b�`	^���ѝZ�̃�6:��T�@���4w#_a���P@/���P�З���Y�W̪7Cn>%��uQuu���*Y��1*����v-�b��}5���w�M�ud�Fh<	��w������W���A�3*�b�;�C��jF�Rr�wӒ�
��Nnb���O�.s������sz�4�p(%n&Ł��i�V�Y��od�A~:mՍɺ��_Gs���Vl� �dL&�~5z�@ܜ�M����.���A��/����������QD�v_� �`�>v��aa�e:o��-ڙ��d�ι��l���0e5���惣To��qJ�*(�L+�J��[����}H61�Nܷ���D��83?�:�1�]d����)��}r��zo
k�5S��.J����eT)f�P�N$���ޠ�~��s���võ9��Ʀ���68|˘�Q7���.���Rڡ6����ml�U|�v#H�|aJH�U�D�*6�j.�(��d*V`e$��;^vCj�\���a�rE����|D�h�����\��7O����0��;kT�Q%'	�Q��$��غR��Z�������K�j�鋉6�˭%�S�+����$\\�%9�Y7J�C�	5��$�+}����&1���]J� ��S9�ִ��~L��k;��R\/n�Oɱ�ˀ���c��M�v�~���~K$ѱfب܀1`{4����s��V?|���h�	H�����FO�	��4�!Zڇ)���僘�$�5G0T��rBx4�HT�xGi��l=-W#���l���� ��/=��ԍ�w^���n��,)�w:�?�ldo�Ԓ��4'�xs�`����kQ{�V�Yg|�>�H�x2e?��0ztV�0�Y
D�h{�]��j��Q�ċ�c9w�P��u�O�Lb8���,�@'��u�Y�t
"G�ʷ�"=
!e�
|��򷡽�����֢ڻ�� �k�@|���`8�©�M����>��IAٻ�!����;�M�h�P���Կ��{��}KEvH�d+�c�[r����$7���N�76̜!ƶ]��/�P%�:zK���޺؜kgg�0,�P����9 3��� 7G���|&$��h���ͥ��{��@Zr��i�,��j���(Ts�C5�ײG��7��ϗ���0�~���I���ʏe�[[+���<��C�d�}CʱX.r�&�p˦�֗��I	�I���l�A���mE�m�_��nI�]h�G��J���ͤ�0�{���ւ�4",5��
>]���j���߅m����)��5;���:umߎ��ދ��jhP����w��6�S?�c1��>J�hVō���0�f��n�����Wܪ_�_��r�������̩s�ʝ"�o��D���Fc�پ{��TB;r��XP�Q.`�⃣	�����36�:ܥc�#�v�A��+_Z��,��ށe�"�bޤ������$y�Kl��.$U�F�����?@:n�xg���@!.uH\`���
� ������D�M쇖��1H���a�q�͎KU�0!�;4�+����_dт~<x^X���y>�;d�2h�]��
}�bV?�~�|bi��$��0�)�"∍�r��N�(T�)؉:\9U(�qa��
,
����W�(�����J>��z֩��fa�BAH(�~����t��g)J�P�9]7Fb��o��5k��A
g�]i��5��+Ȼ�*`����F8������.��U�04��4��>	�����1�"��0�ڬh�
tڇ�� ���qw���|g6s�����z�ƻ�뷳q���אR�'쒧)�d���&?�;#���Iq��M�!""�JEHǀ�����a񲢬�R�~q�:��:�O�Ѻ� Y��o�}�z���-'��4��r.C��[�Y�->P����m��oF6g2r�e���Y3eQ��27y;#��ޱ_ �A|w���N&�(r�"��}��Z;۱�P`�[��Y����*��GE�oh���7h���:<n�L��n�Ԫ][m+��Nb���7E�>ء��x�@����ݵ�vҽv�[�G<��h��ʵ
|< �Nଊ~�����˒&r	�e�Jk���n���
#�+�sZ�S��wy3Xgv��f�����+3HC�����m�%C�̮��j]rMwKy��`���¦CqZ��θ -.�� S�w`ü
�eep�:��ѷޯ���
�{��
߭�00�=��e�Z��h|m�r?+5��J�ҙK]�>@J�嗩E�q�M3o~+D��"��(�H	x�O`��#s�yP�M���2��9��s�ۈ�dM-��w ��"^v2� �7�p�A��%�EI!&Y�m�)ybi�z��נ�W���}T?��G���|"�I��|���u�ڪeľ��ǔz��f��y�?`.�.FVN��!?��V�Tk;V�!�*-P�7a�Q.��8Ԟ8T�w
�P�����v<����u��I
Cc�R�� k��qf���M����)¸{zI���5t8���N��N�A�i�|���wcw��
��>������w��XjY,x�Z�  ����K�P6A�ϙe��@ /�ΞX �<�M'��H�1�Vv�q%�v\1�C)���4#�40�շ��V�G';C`ML�+K���L��Z�0�Y}�Op[��(���I_�D=.���𮗖dv���7�"`�Ĭy;�����a,f�2w���Y��(�=�&&��U��S(���	�+���l�Ĉ������h���̂F2'3?�U�W����"���/�^�C��_X���W��N��!@ȳ�X�C�㦍[va-$3-ok�֙3�,��,�C�ێ {)�t���6��/�H=�}Q�S�{�B%	�g�١JL�o�>�;�ɖ ;������|ꌅ6i��?m�D����J� Ԩ
��_a���}m"Ŗ0�E�n�4��UB��UB?��G�Bs<��0E��b���2e𔮱h��AԘ�5� F1����)\h�'�6�;߳_�Y6 �	_��g�nv��>A��rȘN ���V�e��?o��N&8Bژɓ�n�w&�Q+Ԩ����D�_�ӿқKɣ�+_����y��{z=#𯲶��m�1����x@K�)��Y�UdX4ۢ�xi��[�N�z�/Q�\�A��>��AJ�p�F[�,�P��~K8k���~td6����ޜT����}��-l~S���j�q�Έ�鏠r�㭓di�����̕�B.^�ȮZ��%�S5Qm��
h7u��վ�;8�Mxm��/��w�DL��l�mt����j�߿'�WE���F�����b�""Ҭ������6Ʈ�y>%���G��$�[0��Qń�\KH�9�^�Uv|��|r�Wt���I����>��;��i�5�� �� ��-�v.>Q�p�J�B=.������Ux�-������|�lA�;��ٚ'l�T��Sj��p��w�)���~W�ܢb��V _Cs&h�}�4�=�{�=n|m^b��c���g��o�8Xf��N:�
͢��\)U�8�srr�;� ��� �1A~
�_ُ=I�M<z=�Z2�fQw��|t�gHK�����7�~"���I�)�݌`�*3��I"�ʇ9���d�o)���"�hJP[�9�y��X��SCK��XRBh��s��R~0z4��G�k�-�M31�$?�Ǚ�Gx���2�� �G��VYs�ն�#�����#8�՗��#�����	����MG<��m	$�[�#�+G��.��73WF�$�8�kJ-MY>Q�ҏ%vF[<tu��GyM� *F�V:]�oV�����ބ�GlMbA��ׄW`�г��wH�F5�H/}�l�<w+Z�j�t��V�G��[�v�]�Fi<�+��K��Ĵ`�K漳U�o�0\�ȟ�Zs�J��iT�bU�T6ү�RE�1��LIy҆,�D��PV���qIޞ�(�@����u��E8r���������z���g�*u��k�kV�>��x��>l�5^�*/1=|�+�p�Ai.n��*�u�S�r�G%�j��@D�ֈ0$��N̆��+����`���O��z1=i&��(Kgd���r�hHξ��uh���ѯ���. ec`[�%nJw&ȍ뫵�����h�/&l���k�$��y������p6� 3�WҰIA��Zi�QOV����������b�<�>�ǖ�v�./SeA:���z�Q���y׫�ܔQph�GX_��l#v���uZ�<q�(Ʊ��z�bb
���#��R�6�[���)��ԣSр	��mտ��_�̞б�kC�8V^#yv<��C�ȝ�Zu���ɷ��L��^
V?[���p요��J@�/t��=������X;--�z����W_�,�=j
�J��/e�{�~��8ڧ���Ϻ8d�V-�a�ܞ���á��0˙o����_��
�]���-�5�A}7�}Z��������8��d��̺撢*A`e'+���ia�68.�;K0��&���׋aź/׻|�0� J=y$i�6RaSm]����yL��(���v���r�1��e�5�k�qɫɣ�L8�����S
c�w% �P7u	iM0��E�S�XM �� L���gi�����8	�����5PlVP��3dq��9��CmH��@q��F�xb����o��1|�?'���uͮ�I|��r�6�-L5�ъ����G)��V�#mUru��,ѡ(:�:����2�w9(�I��S��ٰIe��h��#��� 2�w΍*��d״{I �/-�Ԑ����>��B��J��)09p����x�j`�ݶ��c~Ç3t`�څ͵��������ւ��( �}_'��K�r8X�r���I�0�N�2�8No�3�}e�A�z*��<ͺ�Y��cCbU�WK��a��]kY��,G�Ce� ���C-�R����{��[�ވ|3���	G���n��!��\!��@E�t� 5�2��=�{D.����_���AX�5�P��.d8���,�yߐ�KZg	!�$X?���f��ʦ|$��Q��f�*�����8;�_u��G�A/�$kh��Ͼ�P6�h
?ϢԪ��5>�-�^�u�h�o8fJg@- 1]�7u6����z��M��������h��m�!|Ui?��yU�H��6��@en�Uw�A1V3��.T�5�WB�~-��VFQ+R����!	�;ѵ����`���5ɀ��;'e�O��<��n�S��G\�1Z�	�]�_�f�P��t�y=H�!&I�6�e�+�e�I�[��� i��:�RX��x���[h%fv>7��t^4O���3��S�/��"����W�D�=.:�OXa�v�Q��l���� az�2Av�8��Vj��5���8�@�y�ͩA�W7r�G2$�zD��a@׆�G��|Rm�4L3��Np���:��#+7���fi�c2z�K�-E��U��E5�G
�	W��xR��g�<	�	3��]�|G�H�r��VL��uI@�qn���	�{�󅉾"� E7�Iq^�}o+�q=f�p��1s-b�]f�?ZD�u�]0s�S^I�a"�3�+��lw��7����sH���,c��䮇Ҁ`��1D .���9�$%�Ր�w�����S�����(��,<��9R9����>�O!H�+��*�q�Xx&4��K�u��2��Y�S��[���L=�J!�q��$?�E"��&&Yz�,�Z��A�4t�=K)���V������<>"�?x�/spƑ�~��;䑩vAwrES��bb<��M���}�k�AL�.?�@zs�(�t������Kl��C��<8:��om!�o�Y"7,t��:����|���x���Ưe�K��p�W��D1���y���s��(�0��0�;̀��/�C�A/w�ȵ�+`��7��{�a�^Ο��IFllo�FxZ�.���6�D9`d�}�
�r�!�!{*z��Y�U�Z{�G�qI�r�Zv�UIf/G�� ��Q۩���d�g4��M����C�_��e���D�+ו�2^�#�@`��}G9L�mb
A�9�#'�sj1xu��8;��9�Ү��D{�JO���y���R�&O���O�Sx����,��ITF�g�`i�p&�f�8��D��]�(=��qG�:|��3(�V��Y�[?�.K���\kG��cL����Q��Ƕ/���d��\�֠e��� �t.�� x޻���m���:T�E)E�3vKKvkz���zPT�.�w�4p�i���r��Ô�`'���ZT#K�'�3�x����޹i'��E¶�uO��<qNy�~�s� �r$dXw�+���e-TT��ӭ�/�R��3�:���pW��𕶉��+�5���gjR�y���L�!U�Z�����Tˊ�{J�S�DZVE?�NVK�*ֶ�P��isV��i7~�B����'0�Ã�!���)ἤ����^�@�3����bž���R�W;�B_Eɶ���-��ϾJ�n%7)� �[� p �)(�w'�>��W����0�O��rR�(t�P�ܟ!��ˍ�a4�C�N��h|�B> ^�ZJP�)�Q'��$E6�k�b�@��/��4�[O2[)�/+a]ޒ�tQ2�[3�u�6m_nS���3Y��> G՞I,�J�π˝��w�Õ0�a��R9w&_�OO��M������[��>{�rB�e�P�W�����@�yݯ`��Mɳ�0+�'���V�XD�-bS1�RyW�%3*�����6x^��� �/�pt*S(� .��4z������6H�*��������S��TU�����#k�Z$���Q�bU�YZ����x���'� Ea�Ei�vo7�򺴌�2(����'hZu$��l!"N���鄩�w3�����fu����~����e�/�/�GMs<�ҸE-<��d��撮�-��~� ��^;Q��2yBuG���Q1�Cnе�(��t��F��s����k��m�ɷ��l���n.ѳ��v�:x!'�Sxp0�K�f#�Ti=�v1�{G�&'s)��")@<�AR�g�HwX}ʹ��#ِ���-??�߱aA��_. Fy�T�Чʻ�%�&���*n��$�"Ў�N��')���-������"}58E����9=���� g\N���/�/)Y��1��\�w@�T���i^�����{ΠnU����L돊moH�Ѳy��R�3�Nrm"�7��<e8��b�ӂ#lPڰk'�K���7�7�J�B�����~8�>L�׭-�"�"6zU��S�0*�}Z�(�],睕fZ�]ܞ/����t 6��A�P$�JI/\K�T�&Ė�^�RLz�0�3ac��x������a�UK@�m�����@������W�|q���CM�{m���UO��m��۴� �Hq��u[pI3���)]�#�oT��,F>�b��:�PW�/��x��ʖ ��a]���;�0��;I��Q�Ô<<u�R����8�����R1�h�
@��ND=�na���G,[�#��7���ke.XHs�̿�6T�a%!����|����"L�I��1�H�c�����M�j�_�h����"}���6m~	�o�;�r�?��n��&��*��k>6
�n� �t.H�=��{�;��#<��֪�_@�?��Æ��(����C��;쥽jJ"q�^ϩ\�"np�wX}26�q|[�Z �"���B�a��r�2�, ~����;cd�v�Dt����~}-0��!~F�C�U��U�ʽ��D�ui�lK��U�2�>�r0�
_�Y��h� �;�x%DÜ����	���l�W�j��VZ��������sę�wEh���(�@}Wĭ�-ăc1��/��BM$)�ؑ�����q�E9%��xc��1R��`�)��S$y�>Y![�w��"?�{�;Sz���7(r�#��Zs6rO	9�J��i��5�KW1����P���0bV���y�I�+)����*i3�\m����X[�!��f�q��I)��T�E�f�����Mk�8٬\�:�x�D�R��^_��H�u(u7�Ndj�$��|0t�p��D�Iدϙ|��*2Yu/2���'͚���2��O�u�L���a	�6��
W�U%��5�� z ��o�� ��MC��a�ed㢃gE���DĜn*��`��|��8���ʘ�i�S��줆�&��Aa��Щ*T��N���2p'���ҿx�˲\��D���F%��R`�ި��Q�`[��`� �{�j�tYGJ�&}��A���,A�g맍�`M��#�P��m�J��S���x�Zh9�%��`����*�ݹ7ut�L� �8d[�2��]�������-��==��]g.���m�� r��%�M�Q��Jr"��(=��� �V,yl�$RE%ކx=<�Z�]\�����]���r�ST�E:�ᨴ��wm���h��0�O�rݏ��v�`=dbT�is���}�W�RJB]���SL�h�P�]�����&�i\����C�L�X#y,a}�+w��O�^/T�|�
�~o�}���pŖ]��	{;ٰ�	��YdS��_�V��0~X	���C>f�����M���S�H������<6���}*�uDQ���?��]:�s��� ��R��Լ������u�R�bPY�a?G�yF9���R?Q�g�7M���=(���$��v�a��C�-�H�O̚��h�e�&�_�D���|�8 ı��71Q��+��|��-X[��3�)ލ�L5���䒓�+y��A[�o������)�gpa�@u�($���d:�p���8�~e
�')�NU��߷g��V6�P5=�O-��� �@��n>�`^rQ�9��E[�qK(� b�'��� >|�#��G_~�H�>����J��/����kӥ.��h���!9%�(��	�#QU�<��{�Pq��t0q�U��eq���b;j��������t�P��e� ��5�ؐ�9���F0 �66��rDB�o�OG0���:���D�NQ�[��Ou&J ����íY��C)DM��QRs���gȜY;c��f�N(��=ap�`�q�:|%QN^/�n�@�:<�����2��=%�!8Uƫ������A�_+\V�E]R��t"���쫙^ߕ��5 ��Bu|x`�T���o�qd)�����y��i;;+s�[��Z�D�y�\�Un��6Ò[Y�Sx�B9U�d!H��q���ah��AgN��``���\p��J]��f��ϯ�l	̪��\�� o�%��h��HM�o���._�95L����0�0��ޟ����j���}�m��fzi��`�����`%.䦰�3?���wH]#�	;��w�Q�������+�j��8f.�h�,�]Z.�n^P=6KH@jG�����7�ov��5�;8 %�N��3`暹^=��(%�oG��d�>4�ؾF����hd6 ӹ��V�x~��4��0��
{�U�&�8��x���Sk\��SW&=;�w|l좊\�s�>�U�d���y�"��(�Ɋ��7;2�ƌ�")]:ji�P� ���i�ev�>��O����]�q���
H��v�_9S�@	�]Hn�w�;��n�mL�H����F)Y�\/��Qٴ�s��B�^�C�Uk����'*}���:�]�?,���Y��y�YgE/܂��_d��Y��0i?�5�\;z3�$�܈��be?�I�/
P�������Nt9>nl���&�s�S!��E��]?[O��
�����MN+(�g��
`�F'8^�_h;է×�q&�ؗ��QrZ�U��������C��(q�x�^Z�Ԣ{6��o�H'p����6IH��k7%�^���ɒ��.�����0�-�p�K��~*,r"�V��"���l�]�d��OV^J�.��U�r�m-@y�䗠����`��-L�N�Rw�<�_��؍�զ;���ZQ%�T�S�U��h4=�d��ke���s���� ��W�d6y��JU�?�u?=-�s8uS��;0���o/
qFZT��ᏟJ��?s\*?O�kw�J�0����S�%	��7�r/Jj��z�f�6b\���5�=�'	�]m�)h��?�y1\������X����w"7L&(�ǰ���Yb�Zt�o"G�����e1����F���7zP]hOk�&<��6J�HM2�����v��찑�RoΛ��?�J��Ȕw$b����0њ�I�f�z�W�xDn�ĉ����I<?r�3�g �̌I;�	�0b���@J4ku7j�Dl ^�>��J��P���i����K�޷j���FH�RRR�Ic����^��	�]\�	Bb�w1+ϸ���=O*^v)5��#5}yv�y]�2�W�˻����Bsũ�W"�>�?
��Zɽ��Uh��>�p�vWI��+�v�F;�Q7���/�H/��<pN�*ꋹb�'���
�]�gȺ��d��xpɪb� Y��g����3��⓼w�3�*�b���;Ŧ����G*�`�;M&9��V4�h/�r0,|�n� ��<kl!��ƨ���a��8��Y��;⓪�D5�X/�ir�	�
qP��^��ްOV~�c󻋽ʚ7��@��~�,g�*Ha\K��Mߺ`)t�4.2u���uI������� �*2�ā���S�E��7�Ӗ6z�_ķ�!.�k"��t+o�n��^cN'�u+��Y��X�N��jlXȘd ��xBʍ�S���&���։)ow��x�6/e�z���tL��w�$C�5,
���ʀ1�{K�0����-����5"�����y�>3� 64����iL7�/;e�����v�pq|h��l�P���|�+o.�Н��^7hi K��U�"��v=Q�RO�z��:b��~�����Ps3Ţ�P�1A8��Gk��P��iӦ�����c׵H$q���ã.�{�	 -W}aѐ�(��7��[��<��uU8���mR���[ƞc/����̇���ۻW�����Q�W`�Y���O|�������k����+U���J�6�GS���()e'��[EFhhH>��P�Q�ݪ��D���߽b>�/�����Ta73o:L�pv����@Z:揟�S�5�ʏA���76�_�b�O��J�'�җ����#4�1�8"ps]Op)�>792�h���i��3��K"l��^O��"��E��n����oH�Z�ip��[�5��+���T���2�1��a�G+�嗱v�+7��"�Xpx��U��1'�t91� r׭�����T%貲H����G���]�D�>��8�ds;�"<i�4��#��h g���'u��3�����h���/,�k�~ b%,�X)�x����Y@�Y8>�T�L�P�^DZ�XӃZ���w���;��������uBH�y����H�d���� �hs���+M����	���JPz�t�ez�C4�@��u����T�~ڊ��{-��F��M�)2b�8��EQh,��,+�]��y�N�\�ר~F�3��+@0�c��L��i�{�~UhO�X8ePa�Ŀ
��C�:��ea�	%�aY���Xs_� �Zx��͡��D��NV<�C�}tsY�C�^n��u�V�n���Wux�@��2�[ww�|
�`bK�����K�Dp������Bݱ<E�\-G�nό>v�WMA�En�1�%B6i��,�m�Y�i�8��ZN�/B���*�a����&~���&-Q^<;�h���i��5��j� ����I�{��U��IS�N�Ɓ�����>�R�y���m���L�ZV+��k��h���m
�7V|tQ^"���"�0�M4M�#X|�7����Z�b쩯�*2�f��r�G�Bh0<��^��u�ɲ6<����p`X�l�)�" U�gB&�5+BV��]/���L�c�1�=�����Ѓ�!�Mׅ^���V�;#�:Fw�Ude5K��"3S� �p�oV�M���o,s�Ӯ�w�k�?|8J��3Q��-{P�L}.�.ޘ�,pG��ܡ�Yh6�6��A����AEKݓ��TC�;*�~�!SLw������E���0��n	E��U��}���S_&N�����O uR?�q��~�K<-��J4 ��F7N Q0̳�w�m�76|�$�;8zZ3]I�ɞ��ȝ4]�P>�M��Zɀ]�aP����wej�2'�@!����nz��Ȭ����G3��^�16c���d�Y�yES����Q�&� ؕm�y��J�9�k��7i����i����/c[Z�Kp�Xq$qM���5�-�/�%�9����g'NX0��0AU:��~;�����ZH����g�{YċK��mӂ/�R�s�����
n�M��8d�;�/����!���ic?��S[�O6��R�"�J Ͳ���e�K�Β������ ��I��-�U�q� ����HOږ�#��k_UT�9�����.6M�ڇ�۩=��1~�nu��"QoHŠU���v�w�tM\��א^��zؿ��h�����#��	þv�c�I��#��傠�b����Y`�B�G!0�3w�n$��?���7�>��+j�{��:`�q��dA���j\e�1��(��g��iL����Ȓ��H�о=6���6���Tڈ*���3���cEz������]�&3��ട�
�S�Gp��S������k"#�kښ�u�:r;Y�i�j;�nVM��fKr	�VCYy_"(R#�ŒP�qA�if�&˞+D��z�a�!��ה�O�g�yE� ��q�#s>CY�6q�d$���`8͡��aз)�R�ݕ�Qe�C+6Vi���T�Z ���R��W��N0[���z�,�u��BȠ��;�87�ϭyL���H����"ucuX��U,�7��I��Q)��w�X�f&2[�DM���.����*�g�=!���w�./��U��Q���yH� �,4"��X��Z寫��;�\����iq����U�\����B��d�8��ϧ�d<N�o�E���[Q�.*��W��]β3H��X*&C��SZ�-�v����p�p�k�B��N���en�)r6�����{d��Z
���y���r�䶇o��%uT���#�&qHk���{�`zTL�O2z/�ۀ?��j>�oko
3�� 5�+#��$Χ���0@ �(�X�	Ƞ�I�VH,>��cte|Fիb/�2�n5��#.V����_�`��ɜ���b�D �M�+�=D[n6���d�cw���Y�%��:(&��؇�Ό��e1M��+��<��;�mr�����9]�\�=��.�5�����!��L�v�z�x�\�	SK�j��ʧ�M��R��O���*��fQ`�Lߵ�3��C,9��׸�c"˃�E`u�8�wA�=6�K`Fk8n�p�v���.[R��J�XX6�,9����kǘ����3/��X���d@Zh�a�a��X5���R�� ��G'd����PEe�/[J�#�R�-U�@3�a�/Oxa��.���<(�Dǟ��[��~�P���>a���u����Fc/!:�,:BZ"������cg2���i��:#G}sH��c��m:	��V��㮗��]�B�ғ>��������a�����Ua�E�kl2�ܫ�< 6�$�#��Y4ȑ���g)UbP96��TR �a` ��	պ��,$��=��P�q�˥�'�='%��?I������F����TOY�qN���ѓ�這��l]E�:�\���[٤�j(�p�[�M5y�P�<A/x�?d����0]
�����vM}�����7\��d��k��4ʄx���19����l� �v>Ҕףk�W���<��::��G��<�g"��z������E�*��Џ��\�KM^�"UE����1qM�['�#�|aj��gS�Qt*�y:�� V�J�fQ��*,�<����r]I�ʮŔq�ԙX����݌W��fCcA+����2�L��}Rl��u�n+ ����R��v�R�NIp�sV���u����#S�X��|�4��\.��`�Aw17M6<m�e�+e�z\+����j��Ϻ9�Q"��bM6D?�*��K�%����j.�P^⅀�h�PZR���ć }�*@Pg.�?!<Հ ��M'U!B��<P�{�[�U�0F+���{�AwR�\Eaؠ���V��GN�LS+���Xdgߗx>�}��^����D���[�����,ה_\�J�H�%]0xxuȪNF/�o�M��X�ut�R>�=�I���YK��A]�_�=��ٗ��aiI��x�ĮY��+!3'�,��+��'l���\���N��=W.���S!5�r��K%�߹�5���p5i��$�b,�Թ����DC���!�U땂�i}�g!�n.N&f w�Z1�"�wJ����� ��քJ�H,��n#k����6��3H�4�Ӆ�����?u<lX�U����Ӏ��e.9d��#��0wqzW��ctQ��,[�0oC8*']��zۏT�U;�_�< ��M^��7�Y#<Ȫ75�?x���`f5qp���.ts��X�Y��F�;�s�a)���ꄘ�w}/j
+#�a�_	����a�ރ�����9Qh�ޒ�:E;��^ht2c�ra����֒AQYN!�H,=Y΀��"�WZ��)Ĉ>�j\>���y���˹�ikl����f��3��x��;�ɯ�I�ť�;4��MPs(�N �O-�����S��Q�-z��"r �n8x�r��7��ǩ��}���B�{u��tE	 p��r- ��ߓ31\[ ģ\�g=����C���cRâ���c��@��ǕI8k�1_��͋�s�R6��Ӂ���4o�>�=!��)�՗�/���w#�ń#
���9\�4��ᒞ�<z~8��� 	�dD�G�����Q=TG8�w:Mz�	8��1�_���/iof�X91"��Pp��{mch^e"���h�\���9����K ]���7�ŐPl��=j��ϋj�5n��x$�Z
�B�|�i��7����G��Tg�x��K�i�W�IVT�E�zk4@$q�͆h����*����Z�����I��^����������]��?n�of��!����ZR8�a�o��{kO�M�6�a�6��V�w�V+��B*/mKE��W]���M��6t�P|�X��Z����!۹�0���c'#n�%'(��[�3�N����!��y�IS����ߨ���pA�A��X*ˣf���1χ.�{��ΫY�L"�jV�T�����N&���϶���o�Eu�n�E��/�;9�T�R6[L<jI)���l�:8�6���\[�k�)��6[2���0<���x���d@���m��9YC����B��3D�R���@���cy��	1���ny��'�4/B\i�(�.	UPP�Y�~e�kk�h���U3��o���?�9Z(/�wȅ��(қ����c�Wc}� �z������G�$�$�y�&��.灖�1E��"�P��"�&LC8��6e%��Ju�w���8!�����!�|YV�\����9����P�;Y�f˾z
/z68W���[��I�����}'I�������Oy�F^	]�)Ak�b�u�����X[��/o�Sʥ��ܱn�z�xgB�x)[�a^��B���/�o/���,��M�~�U@��0qDv�˫�Do�P�Ào6^� �$�*\i��8�
lK5܃��Ř�R7
;x���[��t��
3�
D����PY�Xd�+,�u�^��j�@zP&]���H|�+���&���f9�^&$؆����w;���F�0��B�𩴴p�_��B΅���"�Zȧl���΍zPcP��Z��j�t��{�w����vu�z���d�G�z|���];�����5C����d\A{�:]�͟7�##�TO����3���?���c_.�Q���52�f|���q�P����X��+go�'r���)��������s2dZ���Sbh@���zR�ؠ��]��v�ȍp��V�[;�ǖ�ݴ���FVR��*{�����!���	FjH���ʇg�%����'�0y���˫`9�kA?�I1��&����aSSSQ��C���y����,̗�1��&������<$�35A,Y�2�ˢ�(#^���ː���o'Z:$�o�Cu�k;��P�K�Y)�raE���?�+�&�` u�y�x�/�<�)�݅�_��#�ж��vNw��	��s�3�8ߋ-������~c�w�X�4����L�2�e���j#I���Jn+ڼbo���C��l9�50eV���vۏn��/�3y;" ��Ζ
��F:�������-nE2b�s��=Q3�`sM�l��)~����m8!�^� :�Z��i%i��!(�HѨ9}�릇��L_���?wP��))�s ��璜U�����������9K�������m®r�ְ�9�7G;�+������q�2\82�
Gx|�l��PL��L�)���J���zO���˫E�x�a��������#�v6��Qt�䞹"6���������2sv�?d���ҿ���z�UX��L=	!~K��dǳ�IX���w�2xc����5�:^ѢU��H��[�IK�a�������Q��)�"��B����&�ӵ�(o�1���x�_�&|�Ͳ�e���ӑħ��%���A��	�Wz:8\YW,"d�������� �3 +��E�{}
��/�g�5�d<�~w�~�<�܊�_k�i�jѰIZx�`-�w��_R�
�g:�f��{$�fS�� ��Pˁ���C[L[@\"�^UZ�}Y~�O%q���s���%�<�|�h�6vP����?��5[ف�"���ʟ��xL!7E�&C�64�1�|�嘯�ɮ���B@}O�d�X3��z�-:J��b���-��r�C@��jq������b�~P�( ���*{.�p��j>z�3�H{ۦ��ŕMԕ��_�񏄓��J�2���B,؉���L��$�?�',�^����L�R0Yv�1`�>�2 ��^�?Ul�"&?Wm�?F2`�t3%L(�S�a��b�i	���h���6Ĺy�w��VO���� �#�`Q���CjO�?�������iv����=a��65jr�^���B"��zT2�Y��>���Ûc��vD ϩiw�X�FۖY/*�%}�����'<�Q���eҘ��}d��\�@ʐ���,��m�LG�+��N�@r�T��Y%�/Вbޗ���͔b4�ƫ�mvXc���\e��ȅIT]"�H�Ϣ�U�$�)�x	��CL��B����d�7qe��G�]��]<2�W]-fD�U�xv}��[/\��r0��קJ��0`df�ë*��'t���/:�~}0�5N=	),�d�}ȅJ�U��/Ơ�R����'`�g���������6C�-��B��������R��s�Z�M�uD����ox�"�6/�+4��;q�|+�A���0]��[��(\ղu�p�%�<
�~e�%�غ�_Kn>4�)���I��4B>�w��,}��k� i�(���P[u��O�T�G�0�� �<|ZD0�����nkl�'�6�&���3/�?��J��1�RԸmgF��� ���yj_��{��zƿ�l�)9�\*MWF�u��!�0fh%�x&�_,�u�V���ԅ��~ߋ� �<�����7֡j�U������s�3�mGJ�Ǚ-�ao,��:���O)����vM���lBK�!���w���ߌI�>dǸ���ͶI��p4������Q�����c�*�S�mdQG�ld6H9U0�J-�X[~����S��0J��`_0�&_`���B��e �W]�I�o�\ "�]�~K���gh���Jg��B���th^Ve<U*���Jznw��ȣ�BaX@���N���(�[�k��ʒ[:���J���q^+`+�`|3z��?�W�����O��Q��sE�T�X�����@�Xb;�V�R�����n(��*�yƽ]sU�0�D;�_�
��s�6p�%����R��J��U�"�1�u�;^����s^R��G��m^����%��Q� ��}�/ Ҽ�!�H�C���;[�`8�ژ��X�X�d�f�En	����6�p��!�[0�=1��,|A x{]!��N�]/4�_sQ*�_=hhJ;����_�[�T��SJ��8����$@���-D�g���fː�T�Kې�s�U7��Xɹy�zw����煤���7]�#�8�M6ߗ�yV�C� A����Z�U;�pn��~nf�*ͤ�����{�_T�q%��1J����"�9i��mv�ɛ�wF��:�W���^)������b�Mm�����6�ݺ]����䓭���("�f��Sf�[`V�n�����J�y`I�XN4��f!9��|vf!K�E��=���?�g�Ʋ ����d� �G!�s�ڝ����
�Ar��"S����W�I{[7�S�-L��9"�.£�-��Kq����ٲ\oȒf��Ie�Nr/5=y���Ia�FI�R���Aw�eh�U�ܘK�o|TF�!|�7Į��<�2:�E���L�VIl�E������)@42���}��v	x�.�$8����� K��A�z�.O���+���;���A��E9'Z�m�>�ih0kr�wge���d������x7�ć�xBƇq�-P����F:�����ָ���c��f�*s��L�w��R
"�j�c��%80�xe0�$a��.C*���u��xZ�\�*����Ȭ{�}��N��&���� CW��'�)�Չ�f�7��9���������j��^ਝ{�䏮�<G3]�i��~�5;@_x���>�1༐�0(�K��aBfݯ[&tB �v�l�S7pZ�R6N}q�;'X��Y��
^?�ܫba_V�]��`囶���
ڢ�b�J��T�f���edY�v��N����p#'�?�o�0�^�p��i����IBe�D+��Z��i��(��΅AԠ��`�F�wnQ�����q��������F�c�K�]8�".[f��E����-����R�lt��vj��fG\?�.�cȹ�M.�x|�����-t�1W[L��	):E��Iv�nL���MR�N��#�X�jQ\�&��g_�B��#;����U�:�f�"�{�2{��@Ɉ
��7��Ε�Aq�(�F<�-�������qd|��
�Jɱ���l�P�Ú#�;h����5��ْ�����x���3h}aNu=����d*lF�ԋ�V�Q_:\�[$@SȈ��2���{�Z.a�ߥ�
��vVN��J��@&�-0�_�S�6��3;���}����6ځ�u�X�XIt����Q$|{��FS8�|Up�$�?� ޻�}��="ε�|u��L�`0�:���I�s$>��䖝�W\6�M8�n؁�.����߼��	����ß��_��j�� �W�^�F�U���\��x�c�f�SIL�e�>s�|m�z>7B�y�������`�+��߈e"��P��)�`��e���zkߤ� ���^]�A��Dl@Ȫ��������w�.S��9��rw��$���wu�:�Q���&�l�/�lX�m���*U'�J&w����&�憅��\bU�L�<�W`I�-��"P�E�0`�6����?�0F��2I�� �S�V)�h�W*�y<���vbV���#P�*��Ɉ���g���~@R� �8������4%纈�����L�c핋������YK�R�9�}�h�0)�����a�M��1Z�3��imŮ�tus��	��̂z�LZЬ�5k�MM�U�ܟ���#��*Ѧ=��=�(� Z����h��b��RC<�<�Ǿn��M��kM��j�px�1y��
��9�!��$<�u�Z�]e�����TӪ��D1 \v�g���f��5Q�o�:�Sm:��y^bn�@ �o��/9�\���=��
�1}2������0�{a����K���-IT�C֪��q1�s��s	Ke�x'��B�VV�J�I�-���|���<�����R�[h����b� ��'��xO�&Ԗ���f�JM+9f��c��
�+�Ny���ݯ���z6�*C@� ���Hl[�������B>��H �08��l���)�E���{�U�^�6��	��t�M(���"�T����C�1��󵰟PY�@�U�
��H��g��"4G��F<g(��脱�1� ����� 9)`��!��T�s�I�/�	\��Kt���f����ȉ�nO�g!� W�*�az~���{�>�^de ����?��Ӿ�Gj�����n��7dM[��5�����%�WC֎��q�LE4�	͹ߞ��3x�]����+���7����S���4��u��\��!*_�;�6G����Dx?��S�x���>���,*�qCgq�rh��l���k
����������C��O�>-�\��\������޴A�;�C��(n�e���ɂ?�/�a&�)��+P�G�8AJ9^uf�BpNl8�t�V��9%��"�2���m�Ӏ�6ڑ�g7p`���!Y=��K�WF�XJ��I+��"=]!DZ�gz3�>�1���\�̍!�f%��V����!0�N�H��oڬ��3��jpG>#����8Hͯ��|��>�4�xsS�"6��&�e�e�x�����F���bwfg��w��:,�n�p*�#p��v�,���2�(�����1���J��s�ޤSD�L��!F%Y����J��|�����en��b��<y�^�S���)?����kl»�u��[-LU�i�/+4m�[-Lyu`��];�,&���bR�[�{⨼��G�Z�˫�`ٍ5�j��4Ƣ��iZ""�Q��;*���nu�jί�	hH<�(a �=�Ք���է&t߁!sF���W꭫6���N=���^��dCo͜��i\wsF#g�(���\�
G� ��]���ɻ��iƂ��T��Et��-�K-��Ľz-��U��ܟ�h:;���7�
@�b�:���^��]�~}~�M�1�8��<n�̩u�;����pAB����44��TayX_����>�;���X��;�6��ʒS��D݊p�5�+��j�]��{�f��Z
�W>ړ�M�d�j�gh��g)���o����Fm�3I�.Y�{��WfƎ�\fV��E�>x�s�\YTRV{ݢ�����C�,������fL�F��x;6%c�0xm��,y<x�D�+TzKq9Î?4��F��3���/ �u?H� K̂Lk����6��Ԉ��)QX�����)��q���kg��4�Yj!s��+��i�#�B���q	4�p��ҏ_�6ຌ�:�]���I��Ѧ�p|�����J�?��ʮB\���~�f3�xp%�׺_ߚ\�D�$F��+�����3�J�X�C�T��f��)�z�W��PjRAH�8���AJ/y��y[��z��������Ӭ�g����V�F�����s�˵���*4�wRD�]��v��'&���ϕ��xp���T^��$��)�hj4F�El%b]�^��Z�u ��E�/�(7�d'�7�$�~�(4���oM��x�.�𹌡�E"�����&�N���w��'��񹭃K?e�r��j��e�ab�eR}0�����6��zDyA\�`�[�+�E₻K	�z�����y�I���:����z�?�o,>߇x0#i"e� 
�z���aY������n���C����z<H֙L���c����i-�X$cݺ&�>��w���C��P�g�
=�kՏT��CR�iD%��!_���Lʂ��kd�C�����p�D�C��1k�b�=7&03y���b�����ΰ�A�-�mE�������	�AT���9r���2�Q��;cT�~��ji��H�s	cK̟�Q�#՝�� sr�C�Yh��Y�q̚Z8�l���O�q��T�U�s��T�F�MR�xۻ-��H�p��$	�$�?��VN��M���pO�g�w�x��%M�/��D!�4��`Z��ȍnK�t���9�sc�	���T<t����!�;�/���U�t:����`��D���u8{+[�(r��*(�@zn��$@w�Vf�	�;`ņ�F䇾���9VV[Z7,,�:�����P������}���뭓K$�h����,U�R`|R��������+d�L+�F[B
�ڷ�3u^.Cf�&9�1��߱DP�����w+��9
IY��x�}����&�B@�_�Y�;��J���}�/o|\��Au{����2���Y�=����w�{7��dJ�X%#�R���h��~n;�ϣ�KA�]��vw.�� J�!�f�Z��g�:��	{Z���#C��n�G%:���<p�{����V���Y�úa���Cpk�"?���7�"�ҙ<��$�o��/�L#��л�wcg�g�r���;���)��8,3E��%v�ߐ�߿\
Ƈ��7��𨮋A=d��iuM����l1�;�i����G�o�t �V�2��ER��Ql���� �[��^�ݟݻL��@pcv?����<ؼ��Do�c4�F�/�kz���)F����5ul��Q)��$�n��KҦsl�+��׌(�-����S=.Y�TȨ�b�� <Y�$Q�0�t���л�x�:z�	��MA�K��=7�E6i!_
�Vn��?٫-6P���S�FN~��xVT)l�b��k����kF�G�h�$|�ޢ����yh�X����K@]�/�Y��N�C�����񸓼G(��5�5ʭ7��?����*�RL�ԝ��jO��?��,�G����0Ʃ�z����qAO4h�z�"^��(�Ҹ|��n7C3�������kw�����'��$��;�D���#�$�Z�o譴������e����S�����Y:��40$�З@�;�5#oV�`�%F	��#�VWK �B�`����G�i��.�� '�0��J��4�}$���yM���d�>/�_fu )�GP���d�������zQ�+͕w�P'�qi�ZS���p^�/}'��s����� �<(v� ���q�&N8&Ri�]�3�i�h?E�1|�P�1�,����)|v�h��`�Rb���&�����Yե/5��cS���U1�@���2J�k�5�X��Cb��1�J��F5���E��R�ky��-���� ��2��2�Ox݀V5�A�y~ETѹ��wÔ�
<2�ž�����%�_��RǣB����n@F~:g��+�Q��?w̯�����#5��,���QE%� mop�Ŏ$4�}�3?�v�	���x1�{b)P6���p�g[w��]?������-qz�-�
_I�%>'v2 b�X�)܇p�!��|L�YJ��%e!���@G�g��f�pU:����T����R�$��u?�r���\o����r��.�_U
]��CݱKG?%/����oF�R\l�3�#2���md/q	3j��屫�xX�x��m��k7��@j���A�%�#��#��u[�9�T�H���l��~�֠�q�Ⱦ���9��'-��X��-"W,����y�xY�� H-(�63>ҩ�Vg\��Hz��!]�b
��d��u�M��b4ȯT�e��|����ڎ%Y��e(���i�	�.NZ�Y�a��$�V���B��?����B)wi���]V�;�T����b)K��BG�+�ֻ����E)��$�іX�.����{@��_���/f�~nPXsu��������E�">ʅr�����07���qG��E��A�Ԩ�-���^���B=�L����mo�dw����.����F7��9��*�����e�G�}�7�Rxc�S�Gv����g��"��n�H;��S��Z�y䁩��C��Ks�K^�B_���4��U��zrQub��B�{����{t��;n4����n/�s#�*��{z����Pb�I�aL`���/D ��ɓr^'Je�pT�>?�3���m��bx�X�\�2��	ZZ����=J:4µ2�s�6�Y
\O��gW?���K�������ڌ̎�f���	�n�n��j��C�3�oJ�: �?9�z!�ec�7�y��`k�[�`{��C��)��D-L�=&P�.����s*6}�4�%cT.����$��d��v���l��.E���h,��4a;��;{�Xr��:@8�-����t��_��jQ��l���<B�]�J�<�
^ReD@;.J��A�D�R�W���]��I�����R!�������CR�����{2l�"� ���d��<*���̣Uhz3�bE��8`#�O��g����R����V]�_��� �jgB���$+�O�H�ǖS5��y��(�v9o1���b{���>��zH]t��Eՙ2�����4a�y���<yeX\^��"�v\��6����f� ��?�V��)�&]��h��������#���Y�~G~���S�l������YWt^��f��8��KD��e�uaZ��Lc��&��!����:��)��	-����$P1�+h ����Y2�i���߼(�}������ɽ}�m�3����G��
Y4p]^Mg���Z���ˣQD��o�A�c�7�r�1��6����#߿��)�uHX6��?�t����r$�U�/M�#e���f7��_OUg��ͷ�gPV�� b�Y���G���Y;�k�r�;t������6|�73?s:&K���o������M]G1�^���)�ʸ�)�4ـk3GMu�Z3`��ג_�)`�>O�'Y� w"�zGI�:�/+�yI��@��f��Bw�L���ՋK��$�D	mpaK��N ��e����)�����$�=qw���婙|r�y*� �[fWS-�+x��b�P2$���f����������UH�1x���������e8�|�DǞBE���<��"�h��p{;��jI�%�m$�9Zg7�P� ���B1"N�)���Z`���w}A�N��?W3��椨H����E�ݘ��<��7�ݽ��պw5s�{�i�n��E)�����X�:�vQp��]���]���8&Z�5��#��
Ѿ�ʍt��|uy��L߯�_T(������s�q���=��Ba�q��`$S"����1�`&خ�c����(VCE8�-~$������G`t�E�0 ��B�A(�V8{K�}[�����	AW�7b�w!��,�V���P�ɥ1���|�ȏbX�aw�`�N���B��e�0P3vV��A0-�Q�M�dƟN62�Nb��(c��?�N��iDEߞ��U�$1�4�o�x@�@�x��a�,(o�_ѿ)�ę��"[��~��������-��WO�t���N�.��d*|^�V����阾W,��FCtn�%�h�x|�Y�x'g�-���m�
��~|�L����+�$@eiz�/	�dr;�(L	���2M���ť�_\:N�9�]��۽͝+���̩�gղ��4���=�#T�q΢ ���E���Dy��@!�,�I�Y�Q;�o���+	�R���,�Xm"��X�pZ��~S��S������t��Ϊ�Z*���ֱ+_gg��[;^Dt�-[�L8����* ���V��^{�6���{��ڨxs��au��bJk�s�[9t��j]�\
��?��%+�ϯzK�L�9pB��C��;*Z��b�H6x�r��8�U�MMS���S����w�d������a��T*�~�E��~�L/t�B�p��BJ1�~Q��3B�<w�a�`;�z�0`J�P��N�V&���Z�7�+�"�K	����o����#���M��{6	�1;���@o�A�A�0g��4����\ᾣ!��C�ꖏH2Xi��E,�ze��N�0K�Y$MT_OhM�f@2�a��t�8�ᥴ�C\���f'�`�"��+��#C�*���>����u�A��_h���s޳�) �k��e��O�ohi�*Vi�	��`6Zem�I�o�L�¤K�Ӊ�� ���"b�7���ن��C���%��{���p/��=�FO�l��#��ҫˎ��H{�|]5��1p�)��G��8$AF6�tI���9yrP���'f[D���Փ�j*Hsu�T;�lpv�K�̴h�l_=!m�Ԡ�\���i����?z�$ۂ�|��a5���Ozw9�Ӹ�7n	"'�K�LX%�]��cM?�A鎌�r�	���Q,��2GG*P��&��.3 FbE���*N{�4T0�39����_=,^�����TY��~�0����a��c��_E_Gc�8/� HͰ�jǔ�ᢪW/=�2@�V@5�H#��ZQH�W��R��8It�%�y:x z�sW�����=�П[i�Z9	�.ai|s�g��q$6��t����C����%�����V8C.�>���a��׶ |�4r�7t ���~�ݞ#\a3��m�Y��?dA�je8c�1AG��^��F�g���bv�3����yU��@p�p�����7�fηa�%[M&sa���bx������O�L|�{��X|p�����<Ag@�g��w���C���9�����Jk�"�l.��ZF��N�mI��9���#�q)'\#q� v�g[_:UX҄�ߢ��R"¼�'�3B�[@u�S�q�_(�N��;���i�E¦��ӈ>i�ş�A�p��9HЅ�1��{_�@-����i���>��)��#z����7�2�J��_�$mΗt[4&k��<��[��]2+$94kT�������m����n%�`�_+��F� {:EEW.��5T�eA���[QO&��no���i�̕��-͞��ֻ�����}���3}O���Em4����4eR��9�'TUk�/iFJ�G�V�[&�(͔�a�'[�8��'%�Y�6����4ŔW�+G�k<�L�<���k���Rf1Kd5CE�ɩZ㐿�m�k:��5n�t^�m��Z���[	�ui�\�>ʐ�Yy�U�fz�QI,�z%}�_ �6�i���l���@R�G���G�Y?㍹�=��?�)?X�c9���[t�{��7ú4��ym+�@�q�;
x�un�%�_�� L@\���Ӏc�i�<En��7h�6F���b�ק�	��/�(��e0D����XJ�Ir�<{�6,�N��&�	S=�'O��"���Hyۦ��wx ��8/�	�ܯ����L��h5sNT��hH &���0	�A�P/�K ��\f��--~/ȵ^�z��<�q ��q��=<_!A�[ԁi#��=h|ߺ��L���SU�}1-y0�*�a!	����9tĐ@
��D�b��=L4�%\f�ӕ���$_�k�RI�O���16Yb'��,+H���M
��������q���C��h>������=���O���	F���XrEj��㧥l@8�{�L���$�������5��Cd�?���4a8c�ɔ���#��2D�$>�`��B* G����d�9<���O�x}o�tHK�_@k���r._����W(`�&k�oP}e`���@��7���^_�@���~�����Z6�?�vO�Y����oY5T��3n��?VU���)}`��|r ��p��f�M�=����%����´�u~&�/��#7��t/AR햦��t�8�2��|���G�A؆�f�Mη�p$�7����=��_t�=L�Z�Y#w"\��^[�]k|*ŝ2-�]����Z<{AZG>��K�)G@f#�Q=?S�:�m����꺫�1�$�SoT�6ܸ�i+�'�B$:����HO����
�C$w}:/W���	^�,̼�q�)Aq�����|H�����z�U�㊙7�_�S�)�5uQ��l�&~SoX4"�h`�i����Ooi�Lq��v��W�NU�[*W��L��2�,V)�����ki�⿔M�Z�w> �/ �[�
˙t<�<�'y�*L�[M��_ˏ,�1g��RW��|F�Φ� �({y��5<F�����Wb:�Οn��lb&��^?i������X��g>��Om��i�
�򂛟�-g�Ά�sJ;<6z��ؖo1�ڬ��x챐���H-FTQ[��w�[�3\���bϙ�l�;�P�ah���52�F7gs�M&�D�Jp16�	v�U�ކ�^�y��n������0{Cŕ��v�(��u2�"�4���}kY3����ͬ�����6��`�g'��Y�ɂ�ܭ��?�0��_���2,��{�n?1d"��<@���o��!'�ٹ6 ����j_K����~Y�r]_(��I���-,�.�|������5<d?J���3'8��g��x7�Y���=���v���Q�D2�ŝq��B �O9��������u6M��Y6U�Q/[G��v��jQ K�/����s:��ZJn?�u]���BG2�R��^�Jߙ�%9(���m�]�
�%�(�.i�ng\���7X>���a�y����`�p���)櫬�����O�z�?M)��Ks�l�uን�C�*��1��S���}1xYש�cH�)A^�Vna��$;�a��~%�E?YNc=��@z���qo%.�^����,��Z�$$T�Q ��K���b��>ke�O[q"�������J�}s1psu��K�ۀC��g�lQ����2iU���?�`4��N?l᳸(�6��d,:�T=����1wW�sX�c���3�
�/�f��ہ^�\�|�~�	h0(�'թ��[�#c����5��N-kP��b��=j�t�G�`o�W���O��\NW�E�XC{k�A�͙2�q���6AP�5�1.~zJ�Qy��W­��W���!,C�\Q��E��Q�C_��t��3��sF�D��jO�9�(��V3K��7������	\���X	�$;�'�L�f�����Ty��n�j�%�QW�ω��7�y��Mą�Z�W�;���v:6��y�����9��\����3dQ[oc>��0��A&ܥ����:G�#��G��ۣHr_r&������CO�z��p2��G��o/��|f꼱^Fd�E6����3��B�|��=h�
�*��aW�����j���'��s=�k�r�K�{����~�G�:�J�k[u@B.��nX2������FU9��5&��I�Vf���Y��%�#�����K}'4�]��eP�m��hlktO�$N���~��D�p�#+��~�����|G����ѝ&Ss+]ꄯ���V.���K/Y};n] U6�^x*	F�v8X(W�G�B_vJY]O<���s�zI��y�OH���A�*5V(�Z���z�^f4�o��Ǐg�9�d�~&_[�B�'�m�è�p]k��������g ��!Ry�X�\1����	�S
憶���x��^��a�� �s�Ow�~@f�EP��T��,4�g�٧Yv�����M )"��+G��[2ozЊ�b;�YC�`��ᒻ{����Q3�p�ѳ(]��?��ۼ��&�D�*0:96/�G�;V���vq|����Ҥ�:�!�6P��Y��C�}���{����<�g�4��s4�k�8��7I��JŷӸ]ވ?����jR�]�ðd`���3�gv�~�����t�Aj���^</�{���_� �o$�Ztt&c\Ў7�`���<���8��fDeT��Eb��4�q���/����=JŖQn�`�i�ם�M�'f+X~��'�f�J�J$'},�d�-�By��gUh���.)�
�����+�R�A�����)GYUw�L��.��3�]k߬H��e=�}�E��6F������A!N�BL4�o�Y����Y*���ʩ�%GT��-Vw�dp����@d�gm�k@FW�������/�.�)�8�=��-�i��- 6RdZ�3m�*2cD�2�&ޤ{��R�"�d�u����%I"��FA�B�Ŧ�#K��k
Ò��A6��p=�-��du��5(p�b��?�q��je�ۦ�a4wA��`�J4L4�*���;؝ D^{��*e^&0�T(7����3E���l��B���rV�B1�)��*�l���l�5V�Z��Dȴ�ŀ��ޓ[�79�Cb�m?�}T�6���(�L�ԕ6rI����+K���7J��+b��,غ10s5���GDĻ�F�\���ir���z)�FVc��ٳ��M�n��p�c���V�o��SaRx�>�Soc�����d�j����C���r���K��a:��=䧿�KF)�"db'��'��������oA~Lm����w�<�;NX@x����L-����nT�5-	(�p7��������[�P��ü��~2�S��ѭ8G�ݕA�ȡ¢W>�s����
����B��Aѫ�c�t+�o�U�R>?+�Ŕ��uk�m[�W�M�ݖ�y��G�j}�j�R���&�|�yI2�l˻M7����&oit�x�~*9�a,|�_��sW���pj,�M�ڈzdQ���I��)�-�(�6Zp���s��*6x���n���Z��ށ!0j\"އ=\�vD���t���p����_��jK,�(qg�Y����P>�w\�ُL�R���j�q�Ѿ�b+��%������.i5�u3	�B�!�@wEҨ;������@t��P� ��H�ş^+��T�>�us�W��!��<G����|	.��Rw��0R5g��WƇ��������njűPF��0�k�8" \z�*���a$��NӅp�H�y���4o�9U7�����5�N1��<9��"�:��E�Q���ٍ>\��p��p�\g��k���Q�EL��ʈ����Q
��x��ͬN�r��aY�R��oܘ�k䧞��[��iO����/��pޞ��BS�p��.:�Y� c#�����A4��Y�~)�aOof)��h��F�mC���˷���7Oϲ���c��W~?��_~�ʓ�<-p�bl�4�EVrI�������g��R�θY�	�-j��WT~0���<$�c��d�^,�g�iY֖ԭ鮁��|�o�O,X}��y5>����#ڭ����Ԭ���-����+8��(9��x*!˾�/B��y�[��[HLIɪ	��j��|-&�^�[q�qjU˰hu���󺙩v��ҍ��Aq�f��-�&�	�]�kZ?_U��>�{��;iQ�Lz�d�)v+\��0��Dy(r5Nc�lBJ'��Q2A�ܙU%��M��ֿ�b��I'?��v�#L!��B�(ţu��A3�^�\��Q5WF��Bap/9�E��Z�QKᅕ3¹��4g7�m���t
�d�����R��j�z<�W&�StT��]�`�}�"x��.�:�N���+���?�}^'��7ߗR���M���ض�}s��{��ϟ1�ce�K�}�.5Fu�E�|��a�LT��慹<�V��~;��oq�//��*� H�O�L��䔎���N��퐈��|���ت�JIj/���� ʛ�iC��ߜ��,sO�5l��4w�OZ���:�,2o�jO(!�qo\V�b�ڣ��Xa:n���̗u���fp۝6�>�r�'j��u3���:�I�->�y��VƠ�g�84��7޹)e0ϵ�ϯ$�51��S���KH���|��Vhd�5��l�U3�h$��c��� ���~�@�Y����;���37���]l�Ì���B�{�L/��7� �Q�,!�'^	��dgX��x}�;� �{�i�w,����~g;S���2����c��j�O�#�܂%M3"д��3���xeb�� ���w�9JW`H�	���"�q�<n#[�����WܔI��i���l�9kw�R��vWS����Yo=���`Э��Œ%���=��)�d]q��(�=���Ҿ?_HƮ��ѩ��يC!��F��iU*v�<��۶��6�-嵻�d�ap[ȏ�A�\�{����μ��^G��|t6���ks�Pk��[k]���p�T���h0ٰ��x(tp��B�j�8eR��V��⻰8O�
���y��X��]
�鰶6�Fu�Ɋ�7����Bǫ��eH�8��#˹$�6{�G��J��	ֱ�T4,�K��t�>
�姼��1kSyG׾B��1���b���M]=˄�q�[:��t�N�����D&S�ׇ%��{.�H��W��Qq�)1�gь�����/��.��y>:f��a�~�tz�#�zM����hD꤂	��
���`�����fh�f�L^�6(=ޤĢq4�]��H�D�?����ju��{���E�(��˔�/'k�ܕ; �&ҋ-�Qww�|�����	�5\9�651M�ѼC(�|\̟̈́i�Ye^�>��J��Z����0S�����]#?0��g�t�1�X�x,��~�uP�>���vԉ(8[�^���*�N^i��+��H#9ET0E���lZ	��ȡ����_��e��9��6�?�E�^ߪ1����Z�L.��:�l������t.�0�{�l�U��`�=>��0}\/�=��Q����dZ>�*�7��ހ��]�^h��i5��+=��{��2X)�����ܐ�g�&����8�-��@�s�"?�|�,�ҝf㰥�_��K�ѳ.e�Hwo:�dSp=${n���ƍ���b�װ�d�S(+�
�./?��3����E�=���ڔָO��fNltd�DI1Ϡ#�,�oW.A�|x�'9�q=�j�n����U���%J7ж8t������~�g:�}: �7!�raw�p�vA�;��4��6��;���9SE8QiZjK���뵳J
�62�[�2�tVp���n�J����5}��s�o��,E�5��-�u��k���v��u�?[_��k�Q�u�A}�=�C)y��q��)�=<��lP�眊۟u8�Un&��w�MpX�LB�����oKsB�0�9��� ��ڭ��$y��n�H�A7��C��K
�e,��_��-Rz[mւ�FCu�q���L����5o��u�3�8&��$�y����\��~��n{.��=��a���
����#Z�f��]�\s�y�t�d�o��w���n�Ȃ���y������u�*t��  ���n!��#���!PXK!|�ɪ��gh�>a#���� ��Lmn^�Y;d��e�f�'���S|=)y>~��>����/¤��ϵ�o�.Y�\*g�mQ+ו-U�n����'���Uc��sJ!d���`���XFv����;��-�O�#�	�t#���,��ahTaMՠ{k!!^�T-��6#e_��L��G�XlZl��q�������!�L?�"�ag
:�Z���t�\��x�	���}qw�:B#P����!D _T�.��S2^��k�$��)L�b9�AD�dQ��Gn,ޤ��
�=n�{D+`E�����j��^w�ɓOȎ�wb4���(,v��O"`&�2�9�a�da�c�Z!�3x���Þ��J"]����]JqQ��P�4�;�)HM۬sWj���ޕ���aǊ��g��%6����'�5�8���Q�*Jv� Қs�]?O�`���g$C�J�� W���F�_�ӣ���J��B�;8\������GaLF~�Ij17�r�����D:ݗ�)��7B~N��Wy 8� �R��6�����n���%F�1���#�y�������3l���	�m;4 �]h����P��.\%�t1�/�+ޠX��o�G~�@�н��b���S�@g!���Y��Q|�'��t�ejz�����E�n���j3�6�'�eS������)"3a�,i_5��W�i�vhi%����4���HB����3)W^T��NS�Ҁ��I��� =4����:=����%Zث�����t�$m�bɯ�&9Ņ��j���p�g;ҫ1�`�Sw	����+G�a���l�c�s3��w��Vf����
�������Nn79�s`5h�c[��Zps��1H��@N��V�~D�u��%#V�	�E�p+�D�љ#`�����6����������-@x1��������3(D!Xٯ��F���r����Ϗ���ͅ�5��1C�Eje�2>
d�������U��t3;�]�)i������i:�a�l~��I��g�i�m���,�-&yaGZ���q��];�{sMؐ���vu��[���3~�9�g荃:�]���C�MH�x�Ş��"���q@#قU��
X��~`<9MȖ���6>k�u]���������"�!p�Щ��4˽_�.��L筤EQ��^��b�����B�������*Q�d52�yQ�ɩ�-�M�������%��@����h?D�Z��_�TT����Xt��z#U����.X��®�e��жB���r�ǅ$f��IL�� =�D�?j(ڝ���Ai��Rܦ���}�f�F�)�*;Z��l�㰖��cv؆L����ڝ�	��d������m�c�Q]��c��;�;�n�p����gΙbq`�S��@�)��Zo���� )�3v� ��-,���鞲�?�4�{�5��Q<c几i�^�~/�,�ۧfy��	���v��⼻��������a�eu?7�X��!��[�q�]QPϘ��y�|�]r�?z� ���!}H)�7z�A��鬶�B��60%D�.�]�%���@\P���{�ujV�Tԛ^h�m�j6��3�M7���G�d�"�7�{vi�l�2U����
�݇��:�J���3l���^L{���6~��Y�g^�@��������"Ϙ�c*�~����c,D���II���eҐz�`XI�[��֧)�78>a����u{���x�����X#��G�)����.H�e���B�y�'dg'��W9@�G"Cc�C�����N޺�Ӥ���qF��n�^h�}VP�i��|��|J��4,6�_ߛq%�g�t�& ��ZA�A[+���䑘�E].����s/ZF���Z(�6?�{�%�;eG�'���j.e���d���X���$5yǏReB�k9y���������WI��~m���X_h��OIg�iT-����2�RwH��w�[�K��B����y��I��|��i��6J4]�;z��T��a�UQ�-������J�4�;��_κ1gFp���r:�a,�fH6���'�ux<)�b�=ZA����ߣF�C��uZ(�*�xe*�;2f�1!l�ᱤ,岢<�2(O�o*L�S3g��$�{4ؑB�[���`�_�N���.�2̭��a'��Wcp�2����,a�2xJ=S��m�y���V1o���Jm���"����#�+̍�0g��SO1;�nB�J��&��|,�2�\���`�2s �`�%`�W�*0vj��@|����o/���Z*$� G�P�m�-�2R��$�&�H:�F��%I1?� Tn����(�%yD4'X"�N �������`~�����vc]�}qT��/-�b#���}W�w7QORP>]u�Dv4�ij���[�y�k'�C{3Y�Gn|e�F[��n<[n�M�=�j�w���Siz�K�|����c����@D��>[�8������Le����c�T+C�h&;J�@_�m���p#k
����FҢ2�qAf��������	��u��j�$/��`c pLɂ �VG�B���~bq�����H�1�{{��:�yǦr��9������К��;$e��b�%��X�`��]�D3�Ǎ�V��?�������J=���LYP���PFV��df��T��Z�eϕ�)0�KG��+�$A�j+��Ү���٭�x���JwpK02i��AN�l��2e����w�y�9�`�!^Nk�)���I)��;x�MȲ3���4Q�#����z�p��h�T�@�E��]dh�Ǜ&L���(��~נ�"�V�+?{��X �>.*�T��֜���ѧ۷oN��B�ݻM��r��Dz�`#
S�>�B~/��G�_7y�Z��E��Ĕ�,�oQ^��J����d�kn�,��8�6�Qe+:'K���{��(3ӕjo�������թ�f�������(�
�����������<���·��7��ݻ���#RYH�X<�����;ݼ)dw�����d�p�<�U���J�/<|%P�.�C�_t87X�`�(zm��?O�����m�r=mV�u˷+���s�x
�Z�M���� �uG���8�șY%�_EG�	pt��iū!pV�V�=(]�� @T�B 'َ�x�W;�'?AH4eU�B�����4}Z����XE��b��2���ׄx�f���m��%�#��O�Է[�v�O��:ŷ_W��Y�_�^������0���:6���"0��xX�̤B��ҩ3�&K������m��/�u�4�u�]�OF-d)b����t��=l�r����#*MPN�Tnc-�+�[O	h�>�{3�'��bA�m�9�,�Gk��;tԤ�Mv==��ԅF+�f�F��#U](��+f#ph�>���K� {�p}yO���<`Ej���Ƣ��P�a���9`*f~�e�ERą	�SQ~�6�ʹ��E�" ��Ф�Wz� �����11���@�w���އ��YE�.�����;K�[��:"���������6��B�k�����_�?�����m~��Ͻ�9�r<��6�8� �ӱ��.�t
�Ew��Hm�^�5uce"ӑ\�<[�,�"g%�����㍼\���?(� W���l�Ҧg'G���ս���ţ�3B�.�RKθ{�o�zH�-��N�!����;�n�fE�(�V�K��D'��X[�k�F�}ަvhF$I��o�7�K�������&�J�����ݟH:��6v��]7���S�N�.e)�c����ݎ��z%tmc��/L��V�Y�6�1$����_Z�wS�k�3J�߲���k_28����6��.�H�>���'9/����{�[���/��=�:�̰֎�2����^�͗j�����u�[ v���u;���l����*r�������+�gC��B�[�K� �;�UJz����x�$Phh^r�Ԑ*B2v�ȼa��6�?��w���g���	���PVU3]�`��U�B�ʵP)Ӯ]ү}S��+���y-����NMbT���w��GV#�=���ç��8��,_iB��J)�A�FF��|���t�5�c��o9Q.���������b���d��B�����,�C+Q�:ɓ?����y�~�G1̂�Y�ьD��<���xSc�ܖ��0O-�|@�� o���X��^�E}U�eM5�f�\��Y�� ��0�
`�
���:x��B�W��g�y^� �b�vӱe+�#X��7=ښS��Z��Ə!y��_�"�n�0_%�̟�"���y�c�h�*��{S���1��u�'�q�H/�
%C���ɺ���ye����Qa���/1�}.����a�H�yk��d�'n�*�>^c�&�����!C�RVwG,�\0��n�a���㞔��\��5��1 �ׇ{����1��3�?v{E��"�P�St�o��G7���xx�)��e�10a�;�����v�"��4��Xa�ZR4w��cs�����I�ſ����[��,$�/wdߑ��T�3����t�M[�=F~�";����c����h`��S =���%r�[�VM���P��fx���W����t�I�Yz`���Yu��JƓ{&���_%�lYJ�3Wv��F�%�X�?�m߿�9��`�W��]�[��,�QμS���E%Ԟ!��Q��h������������o��\��J��Z�H�ɹ����a�?��(��q@�܎�w��"�;����X��/��<�_�� y��!K���%��" �bȕۺ��K�R���ϭ�� uS'�S-��x8��]~(���dY��b�0\%���ō��=\A�=�����5
e�`�۬)�	/�kh�AIHMv������M��^�7���� ��j�Sp���:9chV\���7@gU�l ���[�g]y�@ׇ\
���ߌ�
�dc0il-V0;��	IۦX���w�����ʍW(>����=���<�o���yr�ր�!�$+1ٯHΎ>�e�O�����/#��.�t��p!�_��cL�ف���A�TA�0���[����4���4��6��S�g�JU��� �P�Nt�Re�M�H���.ݵJi�K��e�4c�����ऴ�Bi������@��~'s��/]0��@yU3`+�ų9	'zD}�)��