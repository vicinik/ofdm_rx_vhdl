-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QkCSDgaI9qvexExIfBveoWgAMzn00P8smxy2kBz/Z2aJdU6cJ+GjhqPImu/svhYda6l4dcgyI4rA
jMgOi43T1h8TAYtmGuFOZ82glnfBRgluEB/GhFoGmzi9xEjKxX/HwUN3Q/qpvs+zlUyEaEKeLgF7
LPlYmU8EXyLcZwYmOvS34cNu0G4RS1bb4dueb1SlffQhk7jV+XkIXfR7lKdsi9R3os94+CcvgfDt
1dhUoEfpwIstI4utzCqWlc8RXXJmGIcOoEQeRoJ6iJlabwjNuwGzrg34mspzzfhaTZZEVA3IovHG
G5eL9djfB537set/m01pZrD9OX9wrA5jDaGkpA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13440)
`protect data_block
VnRf380t09G6Tl2xA/GJHpimBQqGANUbKCUbEBOZy8WQ/baAcdCjPt7S9uDc91aY0LcfVSdT5T0x
mV8wX5OXMvVQrbq3Lt8/7P0GSPGAhVO3wjPqEWx/FbvPswFOIruH0gU9waxaYMlTlEg989UzRl2m
nWmPEtFnbAtMtzw6x2nA1h1PM+ObFHBdXrh2/FalhKoHaWj1yB79Lt6UOJ4sbeX3CifPV4T6pgvW
/OYK6wWCNdxcNKpn4bKUQVeu6QONroVT0/nIBMveDToSExqMFJzzP0j/EFVodryVNPbFeLbzuoM5
sUSTITaapCXPVgrOfoC3CfIllYTcOXlZ5t37P9RUAqvYdmaqtY7uEC+3bWDjoIHEF34nHMW62+Zm
IuDvkgaF0Pha/tm3MmmV7P65IGSPQD7PsLOxPI7mK0ixiabgD8nYoAkWIT5M2zLJTzHYfLA11F+O
GMBkub2QzpSN04Gey+CVvYEOEQBR5QxEEeI4aHXS5Pb1QgLlt5yoBIaYe2I4jcoAFaXPBXWsaOyW
P4x5ymgsq7ZGAyqFYfvstJZXhVVPNnZTPV058KBN77P2ly2OjAl8hNZH2BFSNW7+xPdlgx5kpamM
Jmydpc34CJx4fADPJ05fjhiCRDrcxwKREn0vHDPI+n7F2pYv0kjTr8XPqolDw7Dm3dUBjX5Ls9zZ
1H6xPaWZqAqRA3fdZ08GdI1qwixc1/WNYcDiRRQoj7TwtSZehbY2SKjoptOG/NS0DK+cddsdbz9O
8bbGxm+C/kUqjBnYwn9GlCmZMnoNmyyNrBSGCXiqT2VlPiANTM1dZ9pW/GY70FiuUPhXdF5K9qVQ
Ibtjh3HgUctWAqmOFm2s1hTQ8Pm2pdzdldjEqwqPoYcwi1GlSM7fyPQnSPKcvSGLcpBZLpWX8vMO
yJnPt8/hgWwiEJTA44WbsS3lAS5va2Fl+vQPuQ4f+Jg9Jo8w2MMYn/tz1KNPBp3q2bd9ENyZCb+A
Tg5P7qbVNGeL8RrYfiU7MEhtJoBANA8r22gpyiYRQOAtLwiqDfp6qKu00oari5JCmpYp7NdAeHLX
iIO5Qw9jD3En9j6OCRa7SXfMGnhg+dTnuzAPT5EnwzYh352uSIDXrpN7qoOsB+IRIhmtdosp/8du
vb8eJQMYah0Ps0CTFDsCzfpdj3aG2Hm35smQUdH6gBZC2bjkDX0l98WomR4QzNEcmmp7PjM3upMA
X2WhRdNEo4jKAJB9tpWPYPUepa+kXv45Laawapy/v39ia6XhDzjoYeMxsJuRTE/ksM4BdClSfHOo
p712qRatait0B/wZmgDRMyWa4LjONaDssd51wkOmZg1psQUKSL3WIHw1GJW4VB+teGX3Qh/4jdTh
qVC1lSGiNO32om5pTbLntyqLr7PV4njtiVTYJv+JUk3349TRZlIwAwDum9RKElRGp53Hj3W2Ksay
U3eVQhObablBnKXVYjopYGbT9L4j9GtC29ecapemY4oNvyoUmF1MQNkJegr8bVrB30DAuQZkFLVG
tzvZo3A37StRMv0oenmVQuakB7Am4NY//5EcWeI5PQb/NIvBg9IR3KAMvtdwRreMXtGIpL4zcTRR
zjmuuT/54vUaeTpgAXyM7kylCvbsKMdcd9TYBrPFf4i7er7Ccf3HooBTEqc6pT11NM1Xny1wfr1i
0cr7Wc24cb0gr6cq3138OP6QWcYIRoWdVCtZmTKOQoTYhCC6MuBlAA4vPk8BkpNEdrDGYHCKRTRT
toiNpJMERg2jdxuSM5d0oZCbCkn9BBGT/l77L1H2HnzbRe97hs3gSv7QprC2ssQi2jds7vDTrX9K
y/QswJsfyUCTKO6sy99lHEMHCFkIEr6q/K9HCLGWTP+Cp2X7GSCmgOrErW2/IUHEz1RYrVH5fSlj
jz6I4cQy33VKh2K7bc0yjfv9gNajxNMEcsFk83tin2NzI/LryCXKBjAl4mZAvoZTidZTg4hsw3xc
7KQT69KdrJMrduszdIOvWvAnt0vSWrfz9du58D3b50U9/PKTU+diXVJsPwEfh1qlqBB58OhT8uYX
uhMla8nOJ6xFVnd9pO/iNnDDZ9cl4Bjj3de8GrTrGQrDK+R0NmkerptTDzIthYz+NcUzCrnqban2
lnBtec7Vnb+ZDa/j7pkykfkDVt0E9L190wVMM60CR+waLjUp5aZcd/ByS5AuBoMo4wQI+sIZxY9D
nN8I1waQ2pirch5dQsWonMfFVemaqral9Ml/sdL4fP25FHXk9YnH+7tIRvRpIQJ9l4ngcjDoC5bF
KqsaaD/kB1uqh+heqW8JcG3WMiIzmmJzPRXGjwECSXqAv2QzRnsl4wSt9/bF3GsvtPPI/5sev+OI
Zeo+gvR46621cH2NoIqs1YX5hLs7iugKl5gNlf+W/oW/JHJ8z3lt0nGNN2Xar6pedHErGoZhEl9X
h5gg2wL8DcZ7iCg98m0ElqqQzMRExNwSBtbFx6POi1QEBUPh0V488nzZxVamntKnuw4acrBhfOBZ
+B3rr2yTJNRkAd75JjkaV3hKl7wwQriyCXl4Owu1i6HSyDLoTKtrTAdAjHQCwOmH41kaukboFw7l
OclVXO9MstePBoJxozHtkHiJF/h4pVuLDpX8uxoWTUHwdDOjCxrKjCGKqJnAug/g3YvIyjcvkLRD
Re6ejCltjC3in4VGlr6e7Mf6Nju1pO9g/+ZRw5DmyAAgAMhJ77eWiiIv5PdWXYXAWq2HLpSWWXW3
I0xxbB/S9Sg+NMdYTBMtnkJE0kxo7kg7drB4dTW7D2mCG4/nO566wt9h3bJy4MB51E4StPUwVBRZ
6PtWqLHk8nArWduJSqW1kw7pnXXiwBYgKhIthzDCHXzOr1DbR1DX4cwj8tUtsbqY9CoduAZsTZz9
J7nW9ass1WClDYG6s3OdH4YeZKi/2L2K8oVWg87iSjfnB6n2da8xijhadOtOTeOLUu2cb8a+RFB4
tihFmOolm5EryxwWY4G5Syt0Dspq5ZBLwzeS1JUniZsG2fR1/I/bIAv+Qoa70sN6LcSYRiC9xY61
voMI1Cbv+M28x0jD2ztvr2cc8QE6Vf/0+sKnth+TSqExcpxmECWMVA/stn42pQCsSDt1KWSdH0fr
KnhXfy4wQJULH8qOjKlyd8CtDS+ZJWxeuYL9x4vlwR2QSfnVa7boQ4hA/lZQQZudFs2XE40yA2RZ
5/l45kn1wUyLYttGQqlKa5lpwtDQ+Oyy7HenAVI7obyDvwWlL/r6KZfoqYxSHzVHqjXQmPZFxBM+
q82gDiRa9DS1B6pxAO6KYctcxned3jgGKaHlLXWuZMs0G48NQmTf0tBSfmBbre33ML/lglMDuf0k
KAJ/YsJYtph8lVv3C8csG2zAIJm65VpJjpCjpuM48cBGMzF5KrDahHaezwRTrz/uK7s/o7yinRQc
4qCOHb2hPflfkcLcP/rVCpx3+LDzrwVzgXDLJ1Vus/lNJ2XIpqT4/WQadb+2E8R0IzVaWgtUCLOW
yvqQydIsex2QD9exWa4cbq6HaGI9lsQ2DGsXBg9pNIdD28ymrW38GU+YPFIndag7KaxYhsHhgrl8
Ar8rQcrXwGsE2SWzok+9w+Z80BtA+VvXrtFgrKZM8GRxvdxg1okrrcCUcwt63JbEMRl31iHvAc4P
DBER5jH8RHy0uIjTo4SGieF/YK/hmX8xMClE3z1JdkJuRE6KAluea3xauX8BdJcP5rexG2a8IOuR
nXL5CMKSKGc8cN9sDT6KFHI60rczRV21BAhlXG5uGrM4Oq/sfZj4vPuRHzc3BW67EwI9CJSxVr25
yyH6s4HWLRXvdUzRzmCaGL7GJDLLG0xBXii8seioVvHoZvfeprpykNk3YtrCNd+PuJhedlX1Xi/Q
fhoEm9BPFBe8zj1cEU+8SkuH8MpuN/dBIt4B8Vq8MWFWNUFaPLVxOQ/Vb0MHjO/7AOQDUMJPcogz
l6k7HEQtjO9LfYiqpqRooOOjNE/b/QoRwszdaH9CdKb5XDBE/9tqqvCRQhI8/RegnU4MErtkAlIo
lLzbZ9FOOcTRSm6SYT0v31ls+m2YPEHJD5qOzbbED8dOz8lvacgJqofpgSv/NVQ/wA7KBzhdEaMc
e+ZnDzrKvztetFBeNxMZzgIKmP0+VLMT/aBHVMcx7rk0z0+Be3FtviX5mKoy7S6KjhM9vApxoGx1
2B4vDBg92w38l4JqWPlQjGZc2jtXfg7HPBUP8RMdHVT0xhnDJnnXVYnhk272Q5pyuUzjk0OgtSt0
bkxsHJxw+6LNvRLvv0TpEFbgxeOxBY7UDR9Swx3Ks5NdVbuPmQhLrCEAnJCvPXrhpABZcXVgJX8a
+5x7jZMYxYtR8uiNbKz1xOSEPhpO0NANKJBl9nJtjlFGVxfsQlkXBDo4d+eg3IQ0XGbgV/XNpE4g
tH11qrxh3HU8bnSXF3YJ/ckJc/11YtIWuBN1oXZcpNkQkIf0BO2Lq4L7h6/k3t/7nH/UidSD7Po5
+l4M01Mffrxd5AECcyTu5+gqntdXrBX4S2mFX/zRU3NVtL9zBaFkZNXp67gip5yQZIeo94dXrMgt
QgXhj8JdT8vXSRKdgPVW6RkJHnSroaFZxQKw2Te9eO2Nyy1diR9om911kHIKEGqvPZeL1aySSah4
arfgUia4llFnxPTFjqGJxKiDh9MF45+3ERYmF5G3V95xs0RiMbalOsh3H/yhzTWI0T2YO5JSj//f
4FbGxKX1SxEClULDkHa/0W0VPQ1FzqmlAcob5iBd5bUMlRh4u0ije6hF4WRtFBBr6NfEhq8ZNUzb
e+Ot83X4N6FsDALaAoYCxthwv+JL+/dNF7KHnzyXHEhrBUktyaf9IfjwMXLlWxcqSWwxrQH9Oi0g
PzIFef8LkLoDvEvtKLRhpoIRQ65fIJpblyDmMKlG6oCV9qsZ505+goTTibEyO0iW1UCPElNSl2UA
zCMf7zeBYNpiPs97cDOWZ86IXmcBgWAgLl3MCDy27O+zUnPpYyCkVsVA+TO2amcu0HY0PKaSdZ2i
nU0F4UmYBB77IGUlDYlaszJ3XwKSnyeln734hYCwcEobaJFLlBOrsjHjuwUp1MHp26qZPCRiRMXz
grp/LNQoERs0/vJ5VT+3urCLN00jor/bFEGz7uOLHg1xLMOMcW4UwLPYqUtTfs228bIV3c9/4KB6
6wwk8KOg3btJNduA6Yn2C4QF8fRRgfdI+T1dCz+XgaQ5/kFXNf7YPzQtsWZVBvK32alxFxHJjcXB
j6SD28RXj9tzvXRpw6Cd0QOMKAzmqZ6OWbWclx0nSlOp/Xv+SkA+dwmcFc4x3epgdPu9xrHQcWwf
KsJ56J9PAYq4hp+1zHZeUkGyMfR2kFmqKPTBG8zso49S+cEoubpaAKzNv6VS9vKDXF2UZ2/ToydD
ec1K06JdkLdwoz9DFYfW8V/wiCOUxT9JLJTcTsDQvsO066ahjlPqZ+H7QjkWSI0Y30zqDClPLAOY
u1jmtTqqxtffKap7u/UHY3UpCsJmn9lQVNnsBqIRRDsPhDbXLMhRlsFFO9k6cJsh98L1nST06mMj
2S36i+a4vXjSWWyfjm3ej0+IIsjZ8Vj0PGQ/GL3+bQztXaUActVnYpApGr07hJ+60EoVY/zHM4zd
b5HFZjaUkoYxW4dUp2PKfA6Uurv++JORN1+Lzgf/+DUyumQFs8u8wOsQ3eshLwP3soE9MBPlxuJG
peNZYylGKbdBzOC49Ad8wwNGXwgbM6Yvt1kht+dVsxQSdLHIHrfMrWR+LjdFiOvrh4KjZyeR9ia0
ggXT0nTpdsJnctemcvkFwLrRpqY8hOaQD8hhMQguFg+Dz1uca6/50TCXrrR+lC/J2Ffql5cjNyLq
5xoT2+oF+zCe4Vdf+XFyWhvBfcgWFNqCvtDPfmykHBLlyGVtg8okZ1+OOp5HZdLOJbRypT33u926
EFh0iBsZ0BNTaKX0shkQe/8J/8DIVxJNkBs/WwG3URr0hswjNcxZZRZ619DgZkjhgE+VyP4pKEBm
HXazx2IMwOgQXebNzTGeXiP+SOVQ/28Px99XM/uoM39OEqVJn4SlteBHGhkgfb1+KqF1qidJZa5E
qcl5Et6ETAzZOaFEJZR9nfQVi2kJoYmYnng5Uh12PrEFq1XIVjp1rIvTR79ZTpUgBUGXhANLKv6K
G/RmsSVrVLF7+ym/3vE7nKGpQkL2i3FYba+XKH3xuA00zVGm7DFYA8N6ZMV/UjE2LYProixFhBYp
QPAWXacVOv6VVRioCSo9I6qxEyv8Ug+ENMrqsiJF3Z+WfzW078aPJGujzXsgtCbdoZlCst0511HX
Dkzf9VIhhkYAxwRJNYLXB6BKas5zbMw8JoN+suQnn0a2Q+cxuesiIQSi3anVNbLYaeJh4/DJkKMN
yACrpCMOx5JHl46T8SB3JaGM0u+zxjXiWg5rKAWYA95utHCZvYmr30BYSG33AASExiW9M+f/7r2Y
tQ3hqrlqMkVnDq+hDaelrOsWY1tT51kSK5N3t738W8tMWXpaFi8gk66zzr9xfW/iGPzRlCRbE3RU
VlqCEqcnbhoYTCUM43qwpK9rfndlYXm1Vh/5rdrCLpqX+//uL3m3Qg/XE4sXzNscw+5ByaiAIw2b
Jp6oIwV5EJ3pQtiXzWEmxjf9BkQBp1y1+eTPefGe37jFf9zBlIyf0mqGE+COwu5PZFwjcily0IIk
h04woLcRpwwX1v+xDberfDjwIyltQd/mkMoBr+f6H2KTaxiEyVppDTYkwpOIVij2mttDSP8EBowa
jl2KidbnqZWaK8Isy8ba2PI/pDlEsnqN4NiWRLK/5pgNCRwmMKqsVDsgrkhsuHj4iLWHRnko5Zl5
6x5KivoV3jieCgDETi0yRsYeomRem6C3kylC71+YGy3aeC0O62z8AC5U/XPHMuWOHlXYHg5I7Imb
gIQ/+tBp3bPZKbQ1q/FJ4rYGnVmg5Bm02r8uJusHnxX8/w5A/W1z5Ehmy7rhWEwznDF0sU2n86vi
b6QVirbmehIKpAYsX5HJIxXeUKyK016AVrOW9SIeYiSmq/XooBPmON6n2vcEU8LiRCF2UKW/M9R5
SiUJnX/i3Y1lmX98DrjgyTDEZ8KOlyJ3U960MEBc8jLQaazFd4UG1ycNWzBajqi9lBBCt41si/E/
aduN14CFWC6eSXwCuhsUZzBeqfY0tBCGK0NiS3jMqF3o7jIgRoBm8Vv6IXGC188h90UD4xOlXyXn
7JuII8cIQV8FHm29ZNIo6WkcFd7rza6q0zXQw8nBs3xBjx3qI6NYnhbVhpi6s6hc+R81bsV2Lym6
jWK94ZEo7jQGCoGFaubCviNwCanCu3507gVnH8tqpvN0ZTelY4zt5OYO445mDxUkIO06/VC6L0aK
koNjVfmqwgjyfmlPcq+KWZgj0+cizAsUV6+7W1eFFy34IQoXWTDy2FLSfUdIdamYUGOZiAFQ5nQD
4qcUme+r0TmHMss0u8axuQITxlXL4bg5C6W0xm5qZUceBqNPLEIWZN2n+bu2WWyMtBmmiq0ixwfq
3QzmV4NtMBEmWlMHeihX4YN4YVnGdQpMm0ZyHFBcRUT63/7vpcmBf8M779Ljqz9+JN6TsElp13G8
3qwguM/FUmRjvJYPGFMkwEEdVvkdCQCo2bOn5aKBrF8c2UPJ+3RPIJYlutnC5ziVu403E4OaAdCv
kBUMZlQa/15tthYsZ0VnRf+ChCs8qLfEy1vGfm7BwpopG0cwWHyDmmuHDnrB38da8bdW7UE4UwTZ
0GXixxoLF9F15VDZMH66RrSxoulSNvX4SVeL1h8Ti/PBUj+8mjjlkjVwOlwG0S6mNu6uj66jMeUY
ejccReZPpHeX5fkaJOyWH9QKvC5BOX94ZJHukDXRaxnFgiFaiKNf2pMJFfniOmzfL5B4Q+rJjLF+
dxSomAMakri+xdiTXy+Daj4fqf4V1ioO9BRf0SRnSVslVMRa03o3bO9JNGey5tgSrb3coWT/hjuS
r7jBZ1uIzs2uXDZq5wMlmU/tNUoQk/tA3OJeM3GQumPm/KWDcCxNqap3rlpAGZQL8gbWYG6cGugV
XeRxAKVugtoJ9I5cH7HPvrzrjYSF0DF+Ixwoa2/hcbi4YjvKjhaQD+a/N7Oql5dYvWarNZ7x8Tbb
R2PfN4o/JGVm4ddt8iD0dX/cY+8HWDL5AbsChzjE3ysJog/LVBjDTw+cOkuYhYO24l8vIieclomR
tgDj6IlMNiostisXYvEhJRbCEFPmM8i2ErxjKENfCsW/GFZ/rAX+YBlVIGId0b1y9X6/z6ASob6B
zIgtPPgzCbcl53enONuwXEmNQyCxoc1giPbQ3RbzcKWmQcAvoCklY3Zkg8I6QMVoS15yIMnA9yjZ
6hsH642LO/VWPLyLl/mGlvRm2RxqZkRTgIc+UoEuvIDMY+z9sl61hd2EUaPcNfNzPFDI9XoVrEWX
YYp+Yuwd7hVScxofqde0027MRPrrHJL3UrD1izMMCsx2mT6PHG+DBd4pcAYEdhy4Djm1zI8O9+Y2
AdQ0FVTOnBSAVQF+iRMJgbpB6VucNb7AcqX6JEE/KW7BTAXzUV0XymWT1/V2IYr3X78Zw2dRDyl0
3/RuA1Qs4RrJrl2eR9UD/eZ/uCmI2ycJdpxMsndSMxsNUzW57yKNfVflIgpOe0/krWnLktvR/Ehm
S40BtgDXN94F5ticwfPvVdyaTaN3rvF6/z4CejR3dylUszUUwhvl5BbmsL2BmO+b6B8x+PDWLenn
dpSpahW2JI2bQmkfBy8HEeVUQYfqG5/qMXg/X9Qq8Co0CyIht/7WHD98y9olTPzqp2C4T4usW3Rh
FWAGLAEJIs56e8sD4xt0+d9aqd39olraQeO/W/AbcaTA8ROgE/EF9JPTTmwWg38YmtY8amdSix92
sJUoWymnGHXafu4EcUTW0ey9pLUOVDrb+uFkN5PlRk008anrS1yObMIj88iUbDObDRUKZjmJMCt1
GUyAfxT9hrq4UwQD8UB1jXJXJi7UahiqyRCItO1xFCpM8tDAeopib2fcTace+n7nm0C6Xh49pQrv
PR70heMmdLBcF0GcQsJEo4uGEw4IN78WWnCv7yfScXM29KDIC+G7VxyDiWN3EYXmzexxblJbJrAS
M4QgnzlQj13QzbphJPXfc2onPhgKe+dIf9JtURpcb2N19TkPiq8n0hHsGkaIvqHFPPJqc/aYcRRa
M37zFlLbUxgu3z0Rh+BA5eUII46Phqxz4tzheeeG9EUmyYhiOPlQEQaNO+ml1J13I+jDlmr+SiKO
g5skSFA2J7IszKTbPpUeKzb2BwL4b6hIz6SSLsi+I9YYVkQ88kaPX3mOEAU8N6C2G67bbVYdTHZR
5hQpZTkGSsLPgKq4z9gWNPNrpEOkwW/dbSp08+a6i7TNXFzwR2hyqu6UbA5Unf1ApVp+vfbWA3Rx
V5WJv4eth0yXrGa6Yqwt8yY2z9nna/p3M64dqEnl+1gHP59mupsDq+1Cni3JTCeZE5UzHxGgexZ4
034/kTHWrCUSU39cwQ35EbhmtaMrP+vMu0nEszeF/Nct/903x3q5KY1PfoBazP+Cn7+/n3yV15Ef
FrXvDDKs//Q9LhLAasb8cKjpSF9MvCCPJiFGGybkLK3hh40MxFwRmoTkdbHZUWsKW5mK3MnzSy+c
AnatAf1exb1+PBa0FOqlFbq685+jK5HQlVWNSmdXtZvTGLDo4T+oIudAqsO5cHyGHSjyNPhocAug
6VeT7cyeST5LdwbhS9f8gNZ+6fp7QX92bDiF4HX3WI/2oqOuXC+yYE6QIaYN+lXH+LVEwFgSJy67
RNplpWvORit3qQrUPIvK+NWPH+KvJmw5EWP8iTTaOODA3gUTeH0Af0m1lfWeRlenII4lspqkDY+o
1yMRRIE/sTsUgO/ukCCZ5PenwmZIcezmq1BLL7Vk64XRRzGa0grrWtKYdnnLjWLrp1Q+dNo8WEFf
Hh1lqgy5dKLY2MFXQwN8FEcMuvNTJM6NfYyAPLujfPC+iM1ofqoGS71mI4TbK3XE+sYw41nkoSAr
HTslgMa6jxKnezQRjvQlMTZObF54AsmOxRT1+/pJihXg9qOwqe1UTUFAVqm04VmlycYA29Ncahzs
auT/5YmIJ2MgK7cdBqTzT2r/wr+aSs4KpWZFx9wU9L+kP8tvu44PGaSWuHKmoU8RjEhJU66T1eG+
sqct3AuDfG2C24ve/gbzloeTlksxl99j7JOMuEdOb0b+TOwYEfuvuRkhHSHXHD8SYXcvpHuaW6hb
f8xpkcpU4NWwaDSeZvfC82loCMN0EvvXSkbNS0cmraW3BdFHznxnXwpV2Q/Mnjr4f+M2ISRE2b9P
jGpkCZLwjBjB8iDJxDA0vF3TXy79PTFV3pa0fI67kVMWxQ6tn5cgP8SCF1Hfx3msxM6NPEEwJtKP
nU02zH3+UnCaFl16XtxTPNISGV9ZtlvPOWzOlUC9Fk/oPKF8+SjYrpM4B5U0ZbHTQKCJgjABUhic
AVh+mxDrCyFODk6yTgK5AC6XYaad0CTEsKPPTndKQMZRuwm32JV0N7nxide6qeGqQ/lZU1uyC3ki
dii+xfmF38ITqucLo20MLCW7/C4V2LjJ5xxEcjfF/4l0SJtb6cfKWBDhz6uUcioImrEPTV2bd3MW
XnBwl5v1PNemcTHvBUdcxrNAjxeaWDDIXi8Ubu1Yhg9Vfb8YNDNumb88aFa++Js60yFGn9yyESV9
7up0S3cB3xj1SCJimpOjOJzXVRHqMNixcIWqP447TGCDlnZv9CkWESjwfOAuwkDUXcrva/RXNdcr
SxsikIjzviv8TLFm6etWpgHJCmRAKsmEn1V1Kpga8qcKyU7Gjck/IHMgEsZAGPYNO1kKVHbiHB0A
I6j8q7En+tm4+8og+GBUt/Xhd4DVP4jKU6T1H3NSn8hMEQDyvdJfcHYjm8xa6PPTqW4kbUIzhnXD
4+L7Ydk2rpNp/ptewGxWxKa6u1lAdP8E5liTSybx86vJOAK8zJg1BonXzVQtby0SDLwBLRRACf2J
oLRh7TgTf3ZpYqqsNn0XNAiYJ6//ko/9nECWK4WSUgwxyPLGe+ZNOqpfJ6ZVikivRTdrepmiqp6N
dO8eoiLbbVYhjscvpvmMDt3JDUfUjPOeNpNGcNlUXbKai4SRJBEvrs/Iifm02BpT4EAzX1bsIr8B
ZnQHRtn2erICUTLoksKOe+iq1WDTzZK2LElUwTr/GOszIfxbX9OAEHK9o87666p83XYBFGz+mWfa
Obh21OfDBJU/b8Js9dNI5TAsT1fCbJPTEV5eLQUulql8YMMONyJZUHaUC2WEtPxDB0Wmi/Q+I9TI
EZGBnIvo21/omgAO9dA7hUaagZn9yISKxkam7PXlvAISYTGF1NZUDdbR5ZR18WZBatbg0stEMK7k
6biY9W7SpYOJPMZal5o4oqQU6f/wWg6tb6MlUXaR8fVU3Tw6u6TeyjCOTVmKvXSPLtCMZNFXcHbq
9jRh61R2fgGMALrMKlJ5ubPK5BFGSLh9Mab7NYs8ZypLbK3vzLE7tKsUp7/wBF6HFWaDhOo9JfEJ
mlEK6y2XxLm9kjuxa+jR04GcLQl5RKDGzK36UeZ1Nm/00rbB6TCwWjl/qLVPBZyECgIJFkmMbJTS
JnAAuG34ce8fsBdKYdLe0nH3ujfPkiaVZupJYqUBgzYYnxGQ2vXc4u+AL34DquDtoCAoZdC56IwB
2yIzrF/WdkIe95HfbrmfrF4j+0MH+Fv7xuVV7XVueewwVt5diruJkgKqRPJn4PqPKNLmZPNb/G3y
Oq44UpUTrwFNu5wr/O/Hcdlw5sVt+0typGvpOcJ13SGAiqXJjB5VMkwLtt4/4n1boaAxUKFONkOw
hqU4o2Br5YgD2DQC3oeiJE02PB3JQWJnL+Kl9EEuTzt4YDNKDCa791YjVCe8WktwCT5w/T+zmc+2
QYJcCSWEWNBaWa1MHxu1/uWT/hK3R3hOyZAqtvfSrWrOAeAa8AD9ug/hoZ6F41y8Z+YuLpgLkd4T
0QMZcG3BYGBPEUZw26sNtPoU4rFMB3Gd+6yo5jLVcTRTLXzPpnVUcWmS4wCPb9L1x1qgpLQcxezo
bDPxf91QU6URDEYW51tn5ZtJ8veVhWJDIAWQJ3OTn7XkkztY0WUMPgk+kK270G5IK0R6BWauYx4K
LcjcCL2O0Eb+GKIt+oAxbH281QlN6PpHYeskQztFxFbsbabwUdXaKNbFNUYVmu5TG2cTJC2ypehN
2cL5Yc0Huel8FW5sQXyErpo/6aLiCiBdylCDsKjxfoiVb3t8P2LgUyD/spiHzBp9mGXCjbsf5AIb
vtfBZviO4FaMSg/OzLhPWNncDCmYMBPK/DCqwC6DM9WH9pEP5p2FVr9d60pRwBWKSvkqEHrDM6B2
NpDKVyvg7zQ+KGyblLYuoOCD8XOlJRDWtpp4rYTYha7otRmDDuMOMKBvql8+haFBp1PO8YxhOCxY
USfW/XaZ3ObIxotLiD+6cHgTYkIaIhwrogquYTpv0Gc1W5AYlYBzL/asxZ+DZ3dJ6qcqCKiWkNEx
hyEbZHisMOezW4+/VY2dIIm0SmucoY0SoVXkK2Y6x44/SH5vqMqV7TfvnVXxJQ487P2nXtqwpPZU
rxDaMXol06AxSzOcLFRcPaNJ/whK1+BmJt76e1BnMbgou3c+zE7RgJzQtu0pBnbvLW1jZ3DVR3PH
pKU3UsRkOwjNjQE2Q9M87LgtnKbGk1s5kkf6w6M7VBOPxtt8K+fJuI8TlOB3Fu1ECFBJ/iErtL4b
PhKrACw4tAoLxN7zFXHgba+lqR/kw/XQQY8vkXDU5pMVY0qEUf2pmhgh/7VzF9V4pxYm/vHd4lqf
4cWg0aC67ShGciHA+73OWNBFuGqBxYPOTSa/hZKgW/tqSj+mru6tb9DtthxCCSXO7nJkjiTUPH5b
GP2jCh9MlrN7j2+vWNmerY2WQqk8Mu1PqcWUN0YoPBstRcAZBorAegBO5O1p5qkKQvHr7gO891Ph
JAK4hG6v9MyGcMdDSRw2YdBxA5TUNBkp41WVvAEdHBTUrX7qAb1fhUmtktsQfTw0vhwdw1eJo/ON
VSJfDzw5oVwZFHM37kE0hE2GGM2Yuf4INe3RK259xwhiLQ012lpxEp1mmFLkQRp3X5axD+fZT1Ll
DEl9+TVIPPRqu6Nn47f7eyUhW1ZnEdXF/SKaB0+FfmJDWjVtiD6hhb4IZ/3YUH/UENrBLBXY8aBl
lBreIx33IWORpZF8Hww8GoJblZFccwKGOl5yW0z9WV+YlgYfOI3Raj51+Q9qO8l3BkP466pquw8a
bzX09pCQ5JLK94XorQVANzfRi8TXvun/WPbUuShbbF4QRmRrX4u+HLnLKr5H2abotuNvRDgcrEhu
rADXCwM3MbeNi+x4FHAEK1BRgmKnBcXGFVo28iFo8yzCMUQzxNkb3R+ioqBhqkuGpEES78wPmW4E
AbOi6+2JpcYjrU9q/4yxgDtE/UC1mu/RVGoEAErvjtgRhvCYam2uClO6aIBTU51tGvHZrcqVwSeY
Zgp6enGV85G5VRbfuMO9AT7sBNbRBJV6FGsNdsZ4epTLmufwn4clpd/eknDhCqWqDPtYmUi5hMOw
uoXMqoUAAYa8eB/1n6pUvUP9Ho3zrfOGNkHyyC0Nfd7yvr3kJB8C+LJiCbWEsVT5z8cE/JTwu4bK
os+HctI0rfHNvsTfuIcPkvMHH6SnHE89/y33zU43Z6dyavk1nvRBu3FVCUmKqzREpRubSA5u21QW
hBywjINbqYZx5pacu1yqofRXpB50pXtgkFPWHncV/U7ut5J7QoLRSIlXvqaGSQFM/nb/VOcTsYqQ
h224v7pRhIY4Xk5Aug+Grgk+cDfuy/OHIBkmX8gSa4cTc4TCQbEJSR8i9pDn7dDczt5FpIMjuksW
MYo/IRvgMiHKOMUNSGEAj53AXk1repmo8g8xHthHa25AeHOyIVjW/5znrqDM7FmoRc2ZiRCp/YVV
VpPBMCowD/RVou9uhDjJJ/wWBFXKfH/e7DZKvLSWNMZFXxhgt7wv431yQ83m5VrgFSMY5CQKW7KL
t7c1qOKpIPC8nxCgr1ntNMMc/UOYGYjY96dldlQVbztAKOsiGj59XvNhqK4p4xFE5FhQdMSibSfM
Fq4I+MA5BVbYKsl0ihnqo+gCwqlZX+36uYgtvG6NC7Y4bYnPAzhrdqCSSpkNpXYH7bmO+Ot+XasT
E+yr6DNVri4XLwXSzQE86SIwyyP7DuFUdKjXtbBHLzv6KxD9+Mi4nVJxe11M5U72+OSjjYslTIVk
LwZwF48pQC9T9U5SAPmmPafnyPMwSCIBQE+RGvwwJq/rETdGqIT+LFsLFB2oDe/Ja1P0fbjjrLFC
pFTa22Bjb68/Hp9W+cDlhKl6nf4RARJD/hiZcp9vhiV8faqn5NX0HVQUw5ah3oPRuHRfqeNx/aXf
oHg3HpHXW+czyItUGkfH2zotShfHTOJuKtqyId+uubHalZ7WN0gYNtPBu/3YBnjolCkpFD2n/aBS
39oMlhNtUMGj3r+6/mJUgK7IKSIaW11CBULkk3fa6viVuXM2y/SkLzEqLIPYDMbSzJGNrDi7te8e
kRtPv3hzD2yZrPvVd0jSrmhvWNqUUpZ9POf4YF0BkhbxQH7Whq89rik6ouYrjNlYjKfmsdi2Upve
zIOoesCyCnvmMcD62j4p1wDCu9A49p2/RI0IhYQmRwnzyI7h2YLp95s5byp3RF4g6uJfMqcR6sv1
dcvLg1IJdluon2QaAQTwKerg9rzu33DN/m5eH3F29cj2UMGiILyAcKufaG5V02bTjS8+slHsaAGo
89tQPajjgJKTRVcav0Gb18gUgLjuU6bQkuAvbOgTIrY5y0eD64xVGq680cN+y9tKyaAxN+9D+j9b
EAENtFjzZDGvpxLvCy3T5SYRc0r5xBQc/G/nbpQLEndYdcIB36iTk6uWpOs6htz/0IJLkm2Lw0u0
vdp8Ssrd+i9P2uAD5P1rkBvMty8anCKfCh31InM1h1ZL46keZml/E/JkShLPClrX6VAF5ziW1vuF
idYiUAHBmNe4Xc2D+337WmBBE5Is9pEOOUlG1OihQDEzha22cfIgio9lNrnKcX0k7aQaGGkNVlCP
+WE+YdArrrOO85x2RGmSvRt40TNxXpaRMw3z2EhyluyjfiwY5OCJEP3uNOOx0VYkTyJjsWmi9Tot
JiwKYzQv30VT28XbbTXiYqR4oIO+nvwkAlx20QirxrjfvHJzd5yLj5Febaf6/jEb18L/unqAo4es
vxcN5lYGhVStJs5zbQDTNiA1oxKw7e8xRwGMr0jxulfhRhmQOXyw0Y2QxHCxjaXFpzjq8VXF5rxn
KqwKvR4hloqC0o8yElpJYLgJ1bKQQYrposcmsyRmO2GMECVtiPpOygMNRYEog4BI8Z5BtnB0mKDN
BW1Vm13UDOH2wKeNZCgyLft25lxjPJdKpcSHozmIZBGL5p2HXTC3En7m5s/Ibn7qQ2WiBDH2xgd+
Xh6wW4GeqKG0bvyFAKkCdMFYYGDC5ZmL3CmM6j5APH/BqNe6xyMAAxKTsiku+yBTpnaWN2tIbRW8
UqOzi6HraUiBMAkwdBIQAEEmeE2ZPlUMX5wKhIl1rBxYcshPJblkRCiSUtk/9a/WO2HykGkwDRId
27rSP4G/Dt7zmdB1F6Pls9Vgd8Fn209CjlIa+jQEA5yy5Yc5toXUCLB4NjuTAJxtL9g50qH1gzFZ
tBoSugNYKNYFF+TmdVVEI9tQZo5jZreTEJtBuxy6YhjEW2ZzlqL5V3HkiNAs3AwzISE8w8vLD978
6P9jpI5dEAfmlI4gAwU8G+19d2Y15hmVGCSf0cdYc3qUmwRXwJXVQdN02TZDFk2VJKz6h55iQmDu
45itEH1LN5YTTzoc37Hgrm+Rkh6C6jNEB4PRrCiUad2bICeEdGPAobehR4+gFE5YiVd9bi9cVk5W
wTXkKmmqKBrQpUtmdpSbTLVH/hrSxewUjJ/+1XAMj6h8vINqvmAOA61I0Q6gV72lMSiq+LC7nI56
3EXhSKRf2LwLEqHfNoqIw1Mj4V0Qfsnxl/ypkbPzq4Hdqqra+656T+PNLNuKRt7q+FaXNSEJaaLG
viiXMMOQD8GjsP7R/wQhmDz7Nc0Hq8HJDy9TDd1GVZQYCds0CEXMVkl5yD8H3bIbv/TRx4Fn6phn
2zdST4FccLV7Vr9qU6J4XSzbqYCVmQWDAOEPHTT6SozTYXSKGrGUnx9o+NtILtRItz0Y4fNp6P8l
NDBmCqlSiI4hypctuoGfobRtanYNwRWh2mmoZGNj6GnfWSr4UA8PQtweyNxamH9SvK09/rdM4lw+
GNkOc5cE8Kp6e1k6f6zpnjq7Ol9g1vEsUcle/gdWx4ZxDP7s9zb2hHLJUvKd0utmRfzU1fN1+Zns
4XYfMXC3apoLgws8t8j2gPk1FI/f9rWSN1j5uHxWDflMa8Y/oScQDf6JzEeWGE1jF97CA/bKSo/1
CSO/lqTSObzxo/TQ0rL5Iw68T5WDo5h1mzI8aFb7s0XaEcgc5y2BfLztfS2wZa+K2waKNYmACYPL
ftKsj/nLHd0Lzag2e0Ew+KeRTXKePCMCRadeRbz42y2Cqdk0yuCntgtIdyk9hd0b1VImWqBLZO3w
RtYxzTjfmAZbEVx5ru3QKC69m7+5Sa/eFF2ATh4f9Ex9GfLmlTe+l5PDNN6K6UMSZS65ErIJxoa6
JbLtD29uyJ/rZBrQwKFu4R8rbnz0N55YoTTV0R8CLC9s2pZ6RFVEQKO/RaUHcJKn3fC2w9+ZA2FH
NhKoPS/s6bKEun4vQVjJUl0L6Zo2wyvYOOBiNtROJmyVl1aafOhcokdud1gtJ0hFSZ5C3cVFeUJt
Kb4MP2JL+6xcPw5SbGHSECglCeAI1FnM6n3/ICAVYJDC4aczgZBVceaa1qpn/1+xmhbkkkUTarX9
+ERKbfTZ6x5FdMbGvqZ2mEHJXDFK5rD4vVrWw+Ha0GmwopE0fE6TQ3mqSIOgzVtbMJvO28/0RhXj
gAjNjtfAjjs5HTBRN18CPGzk+6W1BPiY5KwbPpO0pLkKj0UQ5/RfQ8D+G3Qzh3UaZNNKfXReKGPf
VCfoFIeW+HprKjfZO4yGKXQXSWKkxSZkRYM7NCVtn/MQjXK/W4jCKJXcqgOBZanrBgk8sRFaJmIE
AcJci66Gby4+GK0bVGOqXkH8Yn0bwVUMRYApCQXY0TSzkggM1msOidTyXXzAPqai6n4IN9GyJbOZ
wvwmOh1m2lWV/T16U4tt1aAnP7fiE7JSVmDTAxxZ0XZNS20x2jQKOhUIYpcB7mmac56882ujSjmO
icJYsZu7fKadNOESWpzIWcGgC6SXuv9WB+p+vu9fRiAPT3E+/ZrJiz7CprykS4+uewTcGCHjznZJ
y8o3CQ4plTXt58iNcuoyeWdyMWP0AeP/BOKFbD6CcWROPiW0ljWmglLrYNhYHu3/g0UYW5fR5BSE
e789Ty1VNt9zUAB+vSEYQ8wneugrYG7R4W1vio7n7CRQClngxrXCGSl7EpWHH0khm8BSGmlA/JGr
Gg/HpfhhY5LEqMhtgESy4CeulCu3FrlO0dnRQxQdCFhkakarr9tVOQfLeOvf3vqHpfr3m9Gk9YOC
mEV55Rkz9FlsVMfT1g5L5QPoEdfxVtISjTararQrgnZZnHCg56bqQLFLajQptEjTCjqKblkj/nnS
tbT6GU0Uwf6XqqWKxCIaklOKxoSzwO7JHrf6+ht7qk8IIm5yJn0jsM5B6f9OuQNTkJHYifpCbTr1
7966Z3kY6yOKHOw3vt93LG3+k41A3hUSGn/nPsqs3tqTUh2hQ+Psi4sM5F68bMgsGNvfbsTkmhRw
m1pKs8GJJAQ5/zsI4hp3RdNPduq04X/CfvBhFq8yv5n21ynzQV1DTyXxWT55
`protect end_protected
