��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒�0G �i�z�N�!�i��*
�tDt�y���_�3�vb�R��/��Ŷ�!��f��,y*�Ծ��?/��U��߹���Gn"�7=L��Y3��Ht�c=����T��V��t���X������ɪ.��ˡ�����It���B)	�+~������Z��zVfș��m�[�,4�0����@0�73�qN"����{���y�ϭ71 �8��1T�����3D�Pz���x�P�Ip�M���"6sд��ч����Å�u*���&��5��Eq�X����m�����:(��i��BΦ�jH�L���5B.�,���`=��c�i\����(�˾�Gv^��&SR7�,<�\��6�h"f��D_��B�� |8���h����:�pYE��C�r��9��r�;|�V���y��u���m'm�!0����"�l��
�|�/EDI�`bo��Fc.4��75n"�i�}�Φ�m8A.'��@�*G��Clq�u�XӚ/iD�c쩺:v�tΧ����/V4Cm2�6r�	�&
}��4�c`\��6]tv�e���T`�����!�e�)ɏ�8K`?/��dy�ٗܭZW��A�28��������.�SJ����9[|<�K�����Y�`o�m��`P�v�Wo�T�>j�Ў���>� �8򐇶���s]���~�����r�H�+�m�|���B9qH�ٿM?�#�����̔�C;���x�Qt�G
�;2��&:�}E�J���(�3[�<(߮\�����%H����/c�4�e9[v 1���p�:���o�P�x�ʙ��YL_`�%Q�[G;L�`{�)`�m�����|<�k�z_ޔ=���"{���y0��u= �>�c���N<�z)� �?a�||�9#�A`=��M&?j+�"+q��	�(�րP���{	L��Eq�C�n����+&���%o_@L:��`�s̆���6=]�PId���',��8�_��'���'��߽`ĺ��m.��/.Z/�X�z78� ����ܐf��oa���ψ�$q�̻R�`���,�_�R�%(x�a\�0�S��<��wW'��8w/��!� �	|��DTHy"�
K�m��M��];0)k���읭�]�?������i�Vs{'�=�Z��
2�/\��y����8��?~ص��H��E�+�rx̗��Z�����k�J���mP����j��1vM�f��|!��;.��������Ђ�s5⥿�0G�_p�1����N�-K������O
�����F�b�,ޱ[q@���Y��T��$?���~�6{�����e�mO��� a��6�f�W�"c�}����c�5P�GTdm��^�c�9��[!j����(`����b��
/�}�T"b�3�}�rl��]Q�[=�5SR%Z�g2�Z"�,�ve�hL�MVu�n6��6���9ݿ��^�P��b�{�4M	8^�m0KK�%������ɮ-�zμ���F�hg5�<.:�рZ�N(�plwa�"�hrk&t�ۮ������<�`���M"R��-q�Dc�Mc�{�}V�3ݧ���_��� ��0LDp@�"R�� ��T�zI�Pb���t�R
$dO�}-¶� l9��f��uUI�%[,:JU9���Y�rr<�spD�R1���C+U���.�j�hL�;��r=h��7.7���?����H/Є�pf\���8�'�3L�=�V��\�Dp�����$������v�� Mx�>�v��{S2v:c2��r�3�j�6L���oZ�Άó��w��d;�<�A(7✽<�g/[(�Z�9�c.J�k�T#����v#������ �j�0:�d�T��,�s6���Tئy{F2lpv������=�oĸ�ϲ��]� 5���xrO(N�=�%t��@�/pj�C�&rt�����r8!�s�Q7�x��,R51Z4/42�����	��ݸ�E$�RK��pM@�w�>z������Î�T����͋�._���
��^ ��X�����a���崞��j}%Y�g/~�oZ����ds�m����~!��|ZqW����^]����jY����4�[_�|+���D��Ն&�4�_��^�q��z<�a������yZX,v�ɗy_���Y8G<�l�{��S�F>ќ�y?r��w,g���Y��'�4׀Ԉ&��k���bvO0�W�Y�z�N�E��e:h�E�ACdL�g��g�5�U+�X+�n5Kf��|�"F�z�m��=����`cS�t�rk�ob\Q!iv���֫ZYr�h�5ٖ80�.u�	Q̱���?��I,}W�
���>|V���u�ܜ
^$���ŉ�L���D�r�ch龛�Ps�+��42Ӵcn�� �~�G��,����=Hn�"��'�1��@�1��з0'����a�i�EA%����@��s��DU#�7xpfnV�� _xX����RwW��A��D�;	yH�!��q�FD���P����؟���P�i����a޲��l�i��	�#�.�̠s�����l�n�[R���!����>!<���X��3W�ޕf�����79�F'l�3��-:�"������\��4g�9�A�~�3�f	����Vjs�������я� ^����9o�w�a[��	��H�yG��LGh>�&B�st��,A����Uo\�~3�pN��rD!���̰�:�_
b;��	�;k0�)/[Y��JPD�3����H��M�&�*V�4jG�La���Lk �4��j1jt�kWp�[4��OO	1ر]d�3{���D\s�;��^@��.�&��ڦ0�s��K�v��@�m�s.!�Y6���:jE;~�����x���S�P��g�''�e8�i�+�1oh�j0D�`�1��J���7���I�o"hw��n�ܴ��ƨ3뢔|���=�Y��	��:R��5� _���6�K�'Ο��Z"�'�\��CKW�"�+ ��%h�ĸK��3Me�B���<�c��`	�����\�.�J�.==���/�2H(j��˗��YC�ĳ:_'Z�}*��d�8}n�VƮ���H�}���*�t��N�f4%kH��f���C2�c�n�Ʌ2{�ђ\�ƞ����M:��s�f��[WC�����uݶ�E/N���p�u��t/a���Ș�Rl��'��	<ԉ������Ђ�)�f�{�
o�p�sX0X3��Q�X돪��C\গՈl��e�C�K~?؏�Z;��!�mⷞ�NjJ���M��	��G�̙O�,�T�r�kB9Ͳ�#|u/D�����9>*ݨ��g<�$5�pp�¦S-������*���A�����Hȅ�S���c6�l��iʂ�&{t�P��:�.�q��b"M�8�G�`�q�l�WL#q<���8�������G�4��Y�4�W|�:�p�YMY��M�cwz�oH_��e���Ƿ�
I5�yrwEo���x��dbu��ń����P�D;�z�S�b�iGObX���݆����`N�p�6镠=���V�&�R�(Q�`�
d;/�l��Σ��;bf@�Y1��s��`)��]/kf��U'Y0ja�C7�R�'�Q��M�%�N�����{�Ĥ�&J�+�<��1~�v���u��4#c@����ů+�A9�h�i�?�2�s������&��!�{GD�}��jr�=����ca/jB����2�ל���)�V�P����%*��{�-+�Q���S�Xʭ0���b;�����A� ���"=� ����Ź��E����XU�|a������J8B�IuÒ칱�5�p�ж��mX��� B��7N�KY�m�M^L�;���F��!�f��Q��c�HG�Q�!��յ;��tVw�����M
ت �����Pz��14�&V�t��f�> ?��52b���kW�Ϻ֯��`���".�� "���gTw�%���
' ��9��[] =�=S�����f��~0f����s�(��^ą�Oz�k��2)r�)Q��U�l1�����*��,��P��ϛA���0y�������YP��u:���W㞩�Q�=����l�Q�G6_�]��3!C^���X��ed��{�)���]���f��~X=�y2�U�TPog�� ���Y/��^��hR������
Vq���-�?�w���Fe�tyt�m�V_t��Q��ݣ
(����@a��!?Th�Ǝ�*�&�������[uȃ�X������~,�� k�:3�{�UL2�ʪRG�B���^?�S�^m���t��L�o��F�a���\h�A�%���1�ѣ��+�k��!	��O�K/�Z����AphP��,��G�kE� ��"+n8�ʰJUUxU4�ZS��!Ǧh^(.􅸯`������WPf����T�(��7T8�p��Pt5�c^0�a��\p2�~�Y���$n;���<��Q�ˍJL���/��ư訮q����u�Os;%&X���H��\k>��c��=waCx��1�-��������Jm����ح��W�1w3U��_ ��B��Y�>e�E��Ԩ����-��� �}�N�=qW=�)OOY�af���#�m�m7'OǮ�z�_��׋�8�kj��a]��T�#x��J���o:�DE�@h_����5m{�Q��w{7��X���Bj�z�6�?���N!�_յ]�/炋�� V���E���ol�o-��Z
����	L:����28�n�+X,�<>�{��!�X-��(���r����u�n�\�Z؁���]�:6���� L�9|1��a���U8��Z�;R����h�bYAT�'P>L[��I\�g"��Riɰ�8��zU�(Ӡ�6�ϳ��T���������,Q9��$�gP�SX�y�z�F�m� �0a<�+�%2JC��^@��U"2_zU4�b�:p�~�p���w��J�jCO��%��W^�߯E�>zeab��`��B
x6~�u�k�þ�������
�?���q��a��G��N�$a���I�3Fȏ�Kݭ�P6��{��S/.�?�RW++[/n�_弼��N�d#Ck<�G~	�"���$E+ǹ�ݧ� t�*����]߷w���"V�$/������~���Ғ��d������6N�Y��ښ�I�%�|���fsd�G��9��mD��l��|��I�c�qe�H�k���Ş��)(������G�#v<]��a�^@���&Glx�
��.��x�]�Kӗ�i/��!F�yȨ�����'���|��m	���~�1qi�b���kPh���dUz$a����<����b���<��ai<:Ѫ�Nt26����kkĺ��c;
��\=,��0i�$��L@$����w��R '��~�;�'Ih���fg0�"M�T�_=����J�{�j���颫9�Oؓ+c%}kc]��G��2�J���J����x�6��֐D�6��:�ىb�E���+���B�m���6�;��2���ik�A@�_���K�˅w5zN�zٜ��m�H\ؽ�_�lx����p�L��Z�/�R��:�J}M�_P������Ę�3�¹�c�]�o��ݹ���}���.��N3}k3�X�ȉA���d�,���v�3�y����!���>hEPS��}�b�s�(
�������{Ȼ&{8}�Y(kGVk�rȦ0-�k;C�fz�atr����:���f�*����$Fn���+N�}r�a4=$ߞ�[��zJ�c�L�;��[��	�9Tw^[�E ��$�������_Hht�dN͒�e�`zV*�2��d��`������˂�ΔJW���{�%Ù��_Ŝ�$Z�� ���;[�Y! ��U�U뤟�a�,C?��*n���|�|���Or�%~|���8O�8:CC�p5�}���^j9 cl��E�������	�G3��H9��o"�"�tş-s����6�-X�;e&�Xy����-�T�wN�wFLY��%���8��&��-W^���'/Z�����P/k �9W���ϰU���+�d�읫����1z�,�ǫ�~rZ����� �'���;�u8iV���T4������+�%qҭ����}>��*�{/����/�~U����^_��ߛ]� O����o���?6�8��h�J#Z5��:\�K�O�0D��
� L~�PH�Wl4"*��x�B*���쳓d�9�"��n��rp5�#Ǳ�!��xgssM*��'���%>�����$�j�Z�����ttzacȭ<.�"�v6� �E�t#
�%�i,�T�^��t��{Ty�Oу0���%��ʿ)8��x��i��Z�k쫭�>�N(O��M8޿�ǃ�H �^��\�p%[�x�i�Ҋ9��������-`����p{���nZ����Ry���d75�*GJ�Qf��[�ko��7�yw����Ɣ���'�D[86���E��C"���n�� �Z�Q.�iq�S�u��0c;�����Gt^�0_��]���&O�<�I����9<�ԩ�Wk��6�a
=������Ep8sMݛ���}�SVa��6��;���X����5�#��zt��"R_Q!��5]&��z��2�@Շy�[8y����7�m���RZ��~;�y�~)�����դ@����@��ݎJ�aso�����L|4qwH�Sm�����8��[��.��Hl��-������Is�Xs�y�t�/�3���wSY����U������&�{;�����[K�r)n�sj��-FH� �D�`����<^��C}�@��MO�~��	u3�
�՘��bh�PQ���/x������fU�SX,՛GA��t,�����O�כ��Y1Mq�^j��^�� � ��q�����C��z�;��!�Wex鱜ψ�D�#%I��ޣ���e�mâ���q��(��-���\��{k�,7"c��	"���F�ў4>=����������&UX���O���Z�ap,�����������:8y�`�ѻ� ]��cɯ�ZJ�`a=�U�ryx�Nz{��!s��kw�-�W�s)x ��0MH*�U0P��2-Ț1Ѭ�2�!1&���(��V|�>(�o&lT�>�*w*L���u�UC���Nُ����Ş~Zf���� �ƾPЃ�A�ȩ>�~KT���C�ϴ�ɥ�"y�)��ˣ�x�	\�s����C�_���o <2%O���� ~Hb;w"ED[������}�C�Q�u���y�?�B�=oy�<g�N^��Q��ϭ+O��d�:�J5r���;9ƺN-Ϝ�^G{l�۹K����~C-��j��`#�����SoI����<�q�w8Mr-~8����g�j�7��|�	�ifQ0�q�@�h���@a����)����DuK�g���#�B�jmJ9d��j7�z|u!�A�Rx (_�)(�mL��;�eai���w�d���s�F�0�9-j6�+�{b�p�������ڬp KC5�T	�0E�lv��O��"��|�ѯ�Ƣ�|=j�8v�O���W�x�Ʊ)�P4�o�"�5�ȶ��N���������9�O�m����!���_�=\"�0u�5 �"\�"B�N��b��d����?Y��/�̌6������ִ�^ʀ�AM�;�A�F����� �)� !�����h�"�~U��F�-ݫ���3��q+Q�&�ij�}Ɖ`�ۈ��&5ʝ<��r�ua�閼���⧷[�1O�N�rЮ��i~��82@����ʦ3�@a'&�
!�� y��-������s�H����h�N�pAH5��tUd� ��6��	?w�}?���-���r�e����yXE�9�5M*�-4/�MS3�P�2#��F��cw�u#.a��>��u�0e�lP�[Do|o�4
c3�7�ɘ�ի<*�Qdv ����K�5g*�^cׂ�S�<)��D�lɥ���%�5L���S��I4�-��i>����/�夞�X������@{��i�\��|��c�h�?y��Α�A�y��}|���G����f�[Na���������#��~"ҥ��-<�JT>S�n�t��%[�M��d�{L��u����?T�ף���\E��N:'����$s��w����b{PD����Z��ҮY���4�
�W�a���>$$Cy�#� �ʐ|I�z�J^��_�6%��5�%��#H�l����}#e�iMm[UW-�{��|�F�t��tJpio��l�=&S|�yp�,��0PY^ `0��6i�;�k��l�~6�-�Q��Q��=l��)�d��� �Lxf��X��� �׻T,r�jH�N����[��U��Z:vrS���4�g��N��r�r��P�Q5!G�n��h���,�Kz����Γ�GMs�&��(�$�nf�V1x4��5LE2F��]�w{���3�a�����UBN�7�E<��'�2�\�bm>�T'�ڸ�cT	rƛ�dH���ɖy��
^�U9�=7
� ���kaW������x�h�$�(l�xҤ�߄8m9�� <� �Ti�.���D��Ax�G%?��*{���S��/��=ĳ�"����LMN�0�=�:�����_=E/����	=�"߫w]�>�X�(��!X>@j}��Z$����^N���ae�0Mԁ�����Ú2}:a#wU�w��7A}^���?���m�ڤ{��3|76-k�gtɂ;Bڔ4��J���N��Qf��S5�D�1=l�ɮ�����&1��{��;�Q�w�3k=	LN�;8E̊'0d�����H�O;�6w�2��M��.����b��<e4\���ea�9�����~�I�f��������=�E-��s��S%�P��j3w�!;Y�,���)�G�wbj�IM���k�Ns�\�c�{�.�(mN՗�O�n�`���U<�n/�$g��@HG���}S�����/��:�k5�u\ 5���ѥ�Q�߇h� lZ}�،���.Y����1��ی4���z�S��,�����EВx��=�(��>E�C3������:����U��0��r����7�rqr�Yy��w�����+'ɴ Y���biHX�݋�^���:����<��w�cX�*ҭ�OkM8���3Q���iL_�z�Zn�(q5a1���g0�����4YO��^�!|�;�"p�  {Zя���RsC�l����+uB�tˇ��H7�,�t'�5bQ�}\~�D������ґ\0�8��-��I��{q	�6?�7�<�_��b�
|�+ʒ3dW��׸����������5ձ�h6��z�]5��d��d�;N��gvhY�X��;�[:�W���D�ƽ�� @��ѹa��a��-���;���E�h��IE�"�ٙ�!��ؘrbjV��(����F77���gJĎ�����,�t�.>�҉�L#N|�:�
�=�M57���
��w�J��o<||��k31��kJ�FS�ͽE�!��WN�����dfѧŞ�4蘡�y�3��c ���̇���A�
�k�4�c~�25TK�@�O�`��!�ha���s<�7ځ����@>�w�`u��!a<����wr)�8���8���a��Zam>���t��r #K�~wW���E�T���h���Oi�1vQ[����7u���TDP��Z<�����??"z�߼���\)�BBĀ S�nd��I�y��ybX������C����)��G�Gd�H�߅,M��]s��^)�u�j�����	*���-�U��/�ɨ>[���hQ/|T�&�b�N���dz�%�-E{o����af�3 �?�o����U��X}#�F����f(a��*b�p�i������P%�B@�����N.���]��^���F���$��[S���Abb�	M�<��z(��;~��<T�9U��еZ[��P����ۥ�X���URK U����D�q�H�@��R!����:���H[g�k{?�H"x\��'��D	��~b���BӦX��?�u����T4v�:@������	b\�i�J��S�跆�W� >��-��َ�i4]������Ǔy�8 ?J�B��`�J�(��s�+B=�Z�F��y�퇕�L{��☫������5ak6�Q��q�����Z�RG�0�����p��,o\��bV���8��2I�Ax�|`K��Wb(G�(h`(l�Ӝ� ʛ>�Ju��_z^���ĭ�l	����JR��*Y3���t�X�k{��~��R�3�Z���c�Z�Nd�XuJ��}�8��ѠM	��-���U�d�g�Ȟ%�2yV���4|�E$:K���`)��lQ	I��ו�*����x��/�H�)�I+�\�Ѵ<f���빧���U��"N8�A�����B���I�U��}�	%�%�D6�]�GIO�ar�R����~��J�&L#��y�
�6�*�ɣ�[���b��Cc�. ���'e��7ۉg @M�{5��e_����v
i�}���;�:��4�۞c���[����LDK���k`�� ��Hi����ܳg���|��E���Q���Z�1��t�2�!���↔��P��L/�;��jI��ר���hX�j���jw�ts��M#j��[������d6�<�0����O0����5���vPv&=�xڶ)�VM�X��R{�Hi�����R�m�_1���pJ��n[/�	��66��*dt�}�wK�{8g�X~M��6r��P��@��O���߆YÛ. ��]��o�ş�NM�)j�L�F4ßc��a��vU�qً���!`�t��Mo蛧 �*�%�7�Kg镅��!�@>��R�\O�j�}�^d�>�����>��I��@���Ƌz�i̓�C�D�0��N[�ի��r�%[)'k��hxMgT�#�\ohF�T�h��ܔ�V*3\���!�?�B-���W����Ȑ.���O(��x8���+�u}*0@�h���f�����En��d����nL�.��T�ja�������#R����s�6*ۇ�f@��>F��
������ҿ���F����ei#��WD�z��w�]�:��cUƳ)X����YL�l�x��M��VՌ����^�-Ƿϲ�)ޚ`���V���Oz��O��I����Q�j��£F�?I�S�8A�rh>���,�4;-]J
��V�t;��3aƝ췌�R��Fp����������W�V��[lA��.x�M#	���g��`R�_�4:��� ���@�|��KN*jߤ��7ʸ�1H�@S�{G>���� @�5����h>�r&|(�##����Q���ɧD}�[�!���o���;���4�v���|U�?��R�e-��O����f½j���|	 iu.�u��Ș�;��>�t��ڕ*J9R91��C�yM�j�h�Ӗ�ˈ�����L��l<�N3�Xa�d��������K��0�܂=�q�uUs�D.���_fE�ɉ$S�4Q��C!����E���p^�n�II_���69�.��
�٬ߡ)l�����iU��	µ!]�BlDA?\��AM��x,Nջ��}�5��`��]��bY�j�7�}�F�_��o�4�U��`��CR/'�
d���ݗ�g�������D�@ g�]q�HH[�"y�#C�{v�)s�6�}g�_��K֔d��F_��Og�ſ5q�x�>P�r�D�@.k�JFP�M��Ƹ�84q+r�'b�[���@�O����fM���Z�8(���t��W�I��w��9B��8]k�i����o�e��R�!A�m�;�a4̳؋�`0�)
S�ȴ>�����R�e݉)۸Ԙ�L��`��7���=�[�.	q���\��SX[��!x�f�P�q�m�f����o����&2蹲�"��/ K�,�GSRG�s�C(�Q�Wg�1�<�Y���t1]�s4$��1��#�ؙ��ۮ��|���z1�5����#n�+����E[�Aejv Sݙ��ZI���U N*�|��}�`i�7�~���b2�I}�d`�g.�����3FVv
�zL�y"�fE�K1t�Z�j��b��?��׋^�u�I"���r�گ!U�
�&�`�TWŧ.�r��_��X��K��`��ZB����~PxM	'��������ɮI *��f&ELeTٳN�����<x�i�q�Q��w�Q�(�E�k��7vT�BNj��B~�o�Ej�4�ɉ}|�T�$����`��k\�xv{T�a}�D�Õ��EY7B������Xp>.A8�{�hy�����#�v +�ZL���~��7�:�S�Kt~:�N�_B沝Z��ճ�47���e�� =�O :�_�X<H�?h�ԉؒiϣ�����[�����X���a��B�*���zl��3Eh|��tSЮ5.��fu�U�E`|�A/{�˵4�P�j�h>@��9�ӋX�Z�$l\�V����`�X<�L�B���E�&h�<G+���c�^���C�����L~9�]��{�zϦ0r�$���c-)8$_u���\Bn͊�$�% ��Ml=�W�Ǫ�ҫ����<y�'�X�j]�w�ۘRΖ 1,�*�~���ײ����u����8^tQ�k�3g������6JQi�1T���H۞�4�Ƭ�Ok�>�)�nψoDH�KD�?��4�C|j _�/�~ )�w����ZF�h����s+&�e*-���TR��/�^�7��Lƿ�vV�X���,~�N�E�R�D%�/�p�)��M��%�j����WRҧ'����k���S��gq��}��2��3RmG;�PKZ�w_��C_�H=u%RWtH5Ѽ�����ƪƽ� B쳚ڨ�?��H�?���N�W�aQC?AT�'1�iʷ��ֺ�u���孢��0%#�SE�sn��8�]�@[�8~inYv�Ȯ�H����ˋl4ݾ�9�A&��)R�������V=����~T����0��,'�#iJ7�&�oU�ir��=]���D�i�<񲧋D�c��^���jY�HS�Na|Mj���;�7�$�3�ç��fl?c?�+.�hs�c W� �|�T��cI����L2��������%��[k�S�Y�9��a6���ޫ h�2e��~2!L(�%|T���dl*���񵢝�vu��gt�!���I��@��Ȓ'u1�A����a^�u?d����o:��G[!����s��nB��LW�bF5�n�ky,�����</���#�w 낃�-��eq&��zT���E�b����k��p��{k�J� �Ӄ��j����`���zh��m1��B��q���o��I(,��|�WS%���?�!:yk$M�ξܱ�N��
\�����-��<N���:�Z�NA�Z��ef^�1�L+����plQ ���PlPY���T(a�=o�;j�D:�NR��+]:}q�4 � ���kmR�`O���t2c頩$Q�>�'ozi9e
^Rr�+<�I�bW����ؘk��|�l����i��u�?G�Qkc�/�g�V���.��:�bO�#
[L��Su:R��i-m� M=5D,�ٴ`�(lkm!Z7a*6#�7U���Y������V��))f�>D]��/6o���l=8V�����PJ�M�Az�
��a"kq�J��)i>����˽�%h
f9M�20�8Y���"}��Q3뇛�ky/i���-��`�'��>t
;�E�ٔ�$��2��B��A*��'�b����
z�B�%���ԹM�K����>2 _������>�!�L9��W����U���Q�]�e��!�����th$�U
.�I�zvMو����5��p8۴�U�J^9�|*�dE��1�r�P&�/��,�#��1kM��Ӆ��X��+}l��{���F��*�����$�@_�\�uKG�J� �"ӑ������#J��
��]s��}�G�|Q#��+�Y��D�;"�r��j����%i��������M�W��*��m'�SͷM����c�."�_R�n���|�)M=~�Q���h�Ob�,��s���3��?W���r�H�9���պ��\���li�a�2�Sk׆�d��Gsߐ�+��g8�aP����?i�$�A����Ro�5�A��2�,X��6X�4�H���T+���;�K,�-c��O�?P�T[����&ǐm�����P�sS�NF��N���{��ܣJ~bԧ��{�+�G�P��䈪�m7颵��T��N/u�%�[E�NMy��zQGW����ܩ��ߔ�\�/w.<Ŀ_�T�����O,7+�gr$>���7KW`Z	Ϥ�v;�KpA�� ˻J�֙��t��6�*O�]��#��;�t���R�h��i��:$�&�F�����ށ�c'2�$�Ҭx�i
��#t�A3	�B�?��M4M� �LH�8'�[���N[����2����1h<�����l	�t�/���|����L�]z��V��%��G��������N��d�򊦿�uM6Z�VV��u�>��% +�ےPnگ{�Cs�u8����4�\�.{�u��9Z͕�x�2~7NuN}j�̺ݽ�;)<i�~@��f���M�O�f}�S����\y~Uv%f��*�Y4k�ҕ�ܲ]Ҏ���t�_�\G5qx:͢���*��AW���J�I	~���{����@�0ݦ��je��KX*{q"ѻ���o�����D�d�η<}>�"�=:ky.�J���������*��A�|�TI����h��V6![�����]��j�'ҫa�<__
8ٝX�e�EZ+�#�>1I\���e'	���K��C��m�4LYL��m#ic�"��j& � �>�:���y�����|W0Z�rtu�
��<�F+g�^8~�����n��'��V�j��N77
���ݗ��[��u
�Ԉ�	�э*��rj���ɧ�mk'u'�Iu��}��ϊcIjt���k����/�o>�!z�Z�O�%��|�Kt)"y3��)������m������M �����[�Նה�����O'<�����փ�� 領������E���ty���F!�s[�)��^��5Ntޕ{��|Cɰ��g��b�&&���)-������a#Ht�/H^?U��፧��cο���<�iX[\�j_]�ǳF�%����n'FD]�c�9�o?�r:����R0�c��΂o0GS�����|�?hv�t��SK�G)��]�v���gс@��8��!��҈ldV��u)�O��QB�D#�� iؗjq���Bȉz���a왖���|$:�� �s���](�G�*�~+
Ř�/��nʃV�S��`k�q&s!j�����ɣA�A����"`�t��a�4y���q�uP�����J��#��*֩����Sc�v�S;$KZ1�����qFT��?���)QaNk�v��M��]9����'
��WĨ�sq�{�������!��[9���>�3�y���lxH��x�;�:��v��<{tb����v��6r�y�$x�K����xf�F����E�q����v���a�^L!�r�	�'�}1�{��%_p���A�4���̑�m�&V�#�=h��trr�W"�i��B�&�u5`p���Sw��=�E!.�dSM�B�9�ƩLfS��h��c>Qb2�2V�J�-% �<)�;�Ѓ�Z�W�ʸ{��v�U(�6K�JJA�~o�2�RSX�~�v�mp���a%:7�wJ�Zuv(���%�j� !�߿��R�$������0��6����X^�}N�@vyf�-���'��%XZ�A^�v��̝�u�4��do���m�M�'�9��l�~=<�e:�3w�M$���p`������~s]l������bݹ��v쟠��&�
LTw������ϭUr?Gv.C����p:N����sx���S�����ï�
��]�)�N#z�v*����I�Iz���|#ӗ�}�#�y{T�k�y0]��X�]Yd��eEiUE�U�q�S-�� �*��
�!�mpJ.�ȧsW+-���ܤ��~Cha�h�.?3��=���(��>C���L�eSE�P�L�m�D*f����ִԭ�����Q2��lŚI�x���U��ݱ�,S��^�l�����a�Mk��5�΋?Vό�ix�J�zwUD�{/�H�L)�@�un�胉����:�!&�X�v��Qy�8y��Ʊ'��j^�<p��W>�}eD���}�7�/f�8����k�NK�F$gG
���=3$�Y�v��\�$։�=�?9DS�\q��+��� g�%m��{Kf��G��k���-��g9&ㄢ1��X��;�4��m˃,���P�9R���rk
j�0��KW�*�0{'����6��p߇�~訕�e �Ԁ��������觀�q��m�?������ k�Z� BI`�E���؞>�l�2��V|Ls���6��	$ �|D �w�~�F��s����E�SZky�����Z�w�����>h�U;K\{��C�E@_���Tӳ@��B(A��76v�d	���?��>^�I��0���,��H�YLjow�A�)��a鴸���o����$���� RX�
ɐ�����7@4��@)��̓�ɾ1�2���B�{��nz=�L3���V��R]������(-�f�N�7�k�q".'���<��D�[$(���fQ����m��J�hƕ��A9U� 1�ݵ�<�F%��D� c�m��N;ӝT��\��G�~�Hn7w����6VKYa�,�ɢ.4ęN�`YYP�����%��%�2t�d0�O�||=(�@�I԰�j� ˘�?�1y�vDy��"�ܧ�?��FB�[b?����1ϪB� �L�m��\?c���3Ş� k�곇CV���ˤ��a�F�IS�$� M�4�B�?�Rc��x�d����m9�1<I),*a�/m�L@B˗�۽���H�vg��v��n�1JW���k��x�������Wp?�BX��Hᾉe�,�I�Prⓕ�/8XXʡZ�9<�U>�o?pv~��� ����MΖzwֶ�Րzwļ?��3bz9�m`P���H~�g���.�u.3o�t� ��,m+^�KU�X�ƂB#���*����7��0V
H��Qc�֋8�\P�3)m�k	�/�cq�o}���$x4M�x��d����A�*��a��9��L��������
��pS�wts��W�3ܤV)�I�Nrz\N�g�+Hd�4S!ZQ8�x
(%=�4"�w�Τ�q�ݫH�i"5�"�vO3�B&!B�rχsټ���\���l;������ ��D�&��w�B���j�:�#��E�qRFަX�o���2�\˾!SK�o�0>كgSC���-	��E0� �h����8x��~/�t�Hͅ$`�R���N��bT���"��(�Äh�l3L����񚁧Ѹ�A�ǟeƠl7 ܍�^��w���I������\"�8��9^{Tf�¤pȻR�+A�?�I��~���?N:A&2G��+��p,��[�xwm�g8���0��N��KZg��J�ա�S���_�V���W�mi��w��"��;g%��Dz��}R������ G2^8�L�]TI�-0;�� +�׫����q�q���-�gr�d��2�q�0��G�b0HH�"KIٕm��!V4��톤�PѓQi��P� �F`���u����(�ߏL����@"e�*�L�*�C��)��O��v!~=����r�Ӥ6h�a�����S��w�wrp%r�Yk��T�٠����/9�:߲��{W \�XԺ*�}Y�B���
�{1O}�:τ������Xi��؉��G����~$Ҭ:� 7���ρx^gax�36�sdg��-dM�us
/��',��������ǝ�tN��
��q^�CG��.-����Ҏ�x��:��#i�Ij���%SM?��[,�{~TS8��-�4��1d��6#���-F�c����_#9�e=Ռ��ܬ�En����0��C�x�M�ƢtL�w�dϫ*�u}${	@|�y���s�'wWY�H8E������м��Ɔ��EQ��I�[8�:�N�*<��9wtlE�jC}$H4�KYqY4F̴�K�m`ΞZ/����#0ź�2�=��.�� J�;����e�G�wO�1��{�s��>��k�zQ��m�[;`J`�UsB��%�v:PB'��J���jR%d4�o:>y8������G�>��0�Ge�QXӅr舏N�w�I�����D��a]r_|g����3��~�FP�T?�ޫ�1׸�s�dxs_a��S�x_���5����$
��?�/���H?�&I>�/�$��m������Ɛ�qPܓ���_�H8wX�#K��E����)2�Ig�:&���=�ꀺ�Q ���;p �,�.����%�8��[Y{L����g'�@��d%z�4
F����a+tP��ߞ���8p���Ռ�+��ݷ<z�i8yOF��pٲJ?rZ)}�+������ޗ�UCB-�F�C�x���bM5��K0u��Aa�)Â��p4�=u�sV��-��������lN�6` ?�k�
�7��x��;-������&�������c.�v�G�5�;"�o����z*�"���|��'F�>��;�"����+�P"y�i���d"��� 4�{�X�ʤ8ӥ�j\ͺ��W��Sa>8�_R�T3�pw���-x�M���f���g'�����;�;x������m�v�G%�v2:��Rc�BG"��"6P��X
���d�-�T�h�$ιJ�$�b�3:���x�y���S��Z[�mXm�9�I��)xm ��Y캁� ����+B�.��"�VJ��t{~��66��0m�fvXT1�s�������.D�p;h&exu�!��,�׏Z����i��=�(���������l�4����
�V��Qs��ǌm>��-_� 3�X�=L3���\ԅ��DD��օ$�Ųzc�,������blmFJo=��W|vͩ�� 	�"
0	�ܚg=.�ŕA3IO�G���(�{��S��:D�rqxK$�x3�)e�	f��/�␢��S�م��:�F����4�46�\�?U[آ�^u��Pv�ڮ�G_��a��Je*\LOEg�J��`�D�O�}
�<2���3�8��%����G�U�O�M���4�A�\�΍�C|ț�a�1���U1�~j�qZ�Hr���{q�݄?\��gƍ0�\(O�Ғ��4k3ß�:w`=Lla�}%f��J��N-Ҹ+,�X0)R׸Í�+�X��\W�&U-ؿ`��곛�0���UfFG�ǣ:͖D�Jb:?��s|�}��ܙΗ� ��u�WC����E�"H#�������~�\�T��`�O+dtRǲ�!�����Ml�+Ё��r�p:����?p��a�cao�J�!-y@	�?E�go��wS���%B�®pG����Ϙ���,�	/�4�/�6^��t���
d�c�wSl?��Oa��f��	��;.�v�&G�� `�����o-<Lo��g����_�GV�U���1�T;��7n������f�L�;[Mj������U��֚�'9����`^Vb��P<)S���~�,����)/�g��ʯ��%@@\k,Y�X��g���YC
�7�wh?E�e����
�a�����[S�)�Vi4���α�a��I�n��^<�˽�_�8�ť6|�;���d,�zG���K`��S�C}���C���7E�)���ѭ62z�>�M�@L��?��1�b0#��Q�\�W!m��1T�_���c|�ˇ��RJ�!����tx�0O��5u?��$낙�����>g�r�EQzJ�6:�f	�K�-Y��C���h� �8�	%�-��S��ڧ�1ږ�N����y;��9|QDӡ�ׅ@�/�s�3K⦘1�7 h)����s�	�Vzcf!���R�6��>g�b&2���-�m�']z�:듫��}u�O<ɝ6*�0uƘic?1���v�p�i�׾v��ulr��n!s"#di���"*�lɈDu��u�xۖ�o��Z-�rlȴ�<���'q�.)�d������@E���H��o��>�}�͆�Z�B�*4�AJ��߇�#�,a���Y3��qѫh�^]n��>TI{R�c�a����ZFyFک%V^O��Ve7n.���Jf�hO���K����Y�
����`���hyp�@8���5�Lq�m�)�Nr�^u��n��϶
�a��9L�UbƼ�HW�Hg�d&E����\P��Q��E���x]I�?%h���z) x �v��c̘{��30ҁ�ng�@��7FYjQ������|ìH��9@�O���1)���Mx��t0��V����z�" a�E����C�;�aߜ�=9�Zr��`O���v ����#4�[���bq�ʊ��9�FE�p1�����}X���(�����z[��NLÍ����',��ڤ��q⸶ܜDJzAe���[����C��<kZ��J���)�X$n�l�:0��w���FN=��>��g��	�tm����薧ݒ����x�"�c��������N��[�7<��:�K�J��Zb�/D��u��q1$��xd�xKǔʔ�]�T����aX�\t�xՒ��q�L/%�m��2�������)�-	� e�:���\xܽi��y�������HX.�� +�����[W].���^D�~��װ���[*�EU]@s.+��F����|����h��ײ��u���AQ��&z�<�����+��rʈ�D-믁k!�Dh��t;v!���7�u��i_Sq|�EǑ�x��S &t�1�BB�׍��,��G��iVp	�W&��J�r+�"F-��j>���-�w1�R�,�.��pT����	㢏���gx�q;K�G33�y�$�`p�	/v�ǣ�����ʠ�d�����f;Z��V�i��%0	��h���z���{�^_���N�
�uU
��q�.IZ	� Sh��Z��Y�����,+yH>�-�	�UYE��;����H�����9�HIԊ�K'T�0L��������2V�DEs7.��g�z_&�;��I#��[dnFk�S�m���K!�>���G�u;.�c���8�'2�Z������S{���9!Ҝġ$(^3&K�E�����<>W��w��S[%�*IA�N��z%r{��Bi3���7
.�w^�?n^ ��4�V�5r'?�B(-N,I�"��9������_��������
��`G��${���P�~���җD|�McU��L)3�(�R5�n���E��]m����߱z���V�e��-~��� +F��}�f$���W���r��#�D���������5VDz|��׻`�OcG�_��3�ք�Y�Wײ���[�Mm/��*�70y9������I­�,�c���niȮ���?�,��j��̹d�|%�WG���b)��?�+P��9��hfMO�/�ѹP���5���N��bs'��vR*�0�c�gz�t���7�&A�f����gl��Nſ�ϝ��pC��w�l�E/{)%�kp$�ƥY����!q'\�������DOW�7�vV���gl:�Ѯ���;�$z�s&5g���U�0_��FhYce��E�2�I�tx��"��A�b
v����[�b�����(�ϗ^�%(�7���\�Ɗ��+8+�l����F�,�^�SbqfґࣜnC2���n����'�u�9<fH���~�\iQ��d���_@�4_[Hv�)���>31p�'h�sj�4�S����9;��N��*��i�7� �_|�����b������h�c��ǘ���<-��ձ��T� [�ɹ�&oQ����
L��:�6����F�=��o���,�'���"�I�L;p�?m�o����c:5���է�8���[;��I���ι��̫��R��ޟ����\[�R߈����I�H�zQ��v~ � &;�W�r�����7+�\�YdJw}�0�Tu�Ѳ��*���H�8i���ʬe��]�s�V����Ix��GOĈ&�f93r�4�`Gh�C��=8�xyC�/
zZh��NV'�'qpėU��m[���&�*:2n��V�֡�@*�I����D�E�g.��YY�ݞH-�pH�*>��<���a��-��D�M�v�o��ʷ0a�$须�}����B<���Qu�>��'$��u������Ώ��Q�E"S�aI���)�%=t^b �ܶ���;�������+8IN���}�A�=Vٰ��L���Y�*�چ.+Hr%(���~A ۬��f�@r��Y�;58��.y|�� 3�X ��lϿ��yMM�����Y��?`Ѷ0���Q���3@��k��⊮������-�ϳ�L��g�뱏��@26t�� �Dsi�y��YNw	$?�d�ބ1��B.�~��zs�{?�o�R���{5T����Ai��|�k��B *�e�3�ѵ�/���'7��7g{ľ��=M��&t�p�$��1�nx����dy�愚���1��y�=�$�)�΄?�p�Z��-@���R�s�w����͐�<k�I�����"U�	ӈn�B��d��>�ui�]-9R4E	@���j�[�r�zGM��a*�$_�M���p��Մ�'�ᣞMc�,`� `�nʄoz+؁�{�_�<VA��Z����%]�u�XH���Oҍ `����{��P��(�$T�P����P��KC);��fd���(R3-�㫖Z^ecM�ҭ�L4 �يz��=�u��Hu�����5���{�,��t�r�},�]���4�M��p���R�ȧ�>�5�%P�;���7�p5tn7�����Yj���kЏ3"
�b�:�ɭa�@�$'��9��������C����������w�d�W����]��?��0;�l�/
�$����b��eec\����xp-r�Y5I�"��[
^?���I=���g���2����F�LxjA�# �����#�a�\��Y�ʎ@�[囩n����{N��b��P!Ai��9.K�A�@؝���çU@���sIS+`��﫨��N�%u�e��"Zl��mUi�������Ȃ2V�j��%ۗŦ�VbM�.# �����n��/1�?�q1B������2Ai+'��֮?�N���3T��Kd�y?��:�<݁JQ2զ*Cz�w�A\^3<��;g�=�[XU7Z�@��C��U*���
�W����%��9��޻���M����h���2�&�e���{�#rI�k�L��,����.��E;^��Gq�ح�k�8VT(���9������#�:}�}��l�����i��m=��s�i�2of�&v0���ړd*`����	�g讟�a��:0-4�Jwv����2L%�/A���<]Ϯv�͝Dۆ-݁�PB����2�-�c��~�tl���N��f�ŎWs5��/�CI�Bo��2}�c�.��`�*!�����5ru��^֊+���f=A}��i=Kl�_���l�M�\5����o�y���>O, ��7��!�$=��B\�k��2bS,� h�g��P�(�����	qw��?��=�j�<�-Î��)K�fO?L/F]�}tg�o�X+=3���%��D����E��5���0�!��s�։9+J�"��6Vr !�u�f���9ą=zg������/;R6���`��p���t$���Q��eW�<f̵ֺ<r>)�!e��MBo��d��9��_}�I͎Z�=\�vZz@���bP�PaP�ܚ�θ̿l��;����RG�~�� ����sB=-��Օ�\U�Q���ifk��z�^ 3�t��3�@�[�P@&�|S	���#��Cŝ��3��.��0R����+t^���T2o߼�����0.��v��ue��=��dmȃx[=�f�J�c��k㡦�,��]���|���h;45 ���]7��-����r�46˝�� Ҩ��1�f�s7��̈������NeM�>9��aW�Zx��s��H����h�q*�8�QlZ} ������j3MQF�ُ�]<�������hb��I�ݹ���pC���#�ڿ��	F=
QW�}|7:n�R=)ǭs��'�d�+_f�n��8�x${g��@G���*�g�M�"~xRS����A�?N�� C�s -����3L�k[�!�@f�ώ�����k~���u�����Y��6ͩ����AL��u*5�M� X��Nׄ�'�AQ}X@�c��Â���UK���!�������"�.���?���PqUI,��8�^��!�"]��x"�*X�ߥJ���RS��Y9��ķn��}����7����ؿ��P;u�N�4�o�fn:��	Y-�����zo[m��.B���,�	������^��v<0u"̦A���M���=U�R�W^���%�ёĐTH��M/���V}�`�E��L�-�?QM/h�l<�ߓtd�׷��¾���c�_G�������#7$�l�ĝ����Q\z��U�A�\�<8��-��c̱�J~i�fo<%D���<.��v�pq1q�S���K��jx6c�B�gq*��w_:����d��stC�Mg�X}�a�D6��$���0���8G�e��̺v[M�K��Ss8�]R��׳p-���׌P{�W�i�Y��U�rp��r>�`N���w:��g��)�y��1�W;����3�,�M�cr�$[(j$�AϹ�4p�
�!�K��,�ᚿ�?�^J������Z�Y�{[��Skg;���B��#+RA�JQ��w,ޙ��W�V*ᶝku������w~�Z���O���8���:S�Y�Q�#��)yҤ�t7��e^�ap�b�(2��:�C�.��	n'�E:Iu�G${,�HEܴ*S�H(�eŞ����*,�_�6n��F�'0�Ms�P$"�q��mS�39��GW(Q���D	}^�&Y�C�"�X�S��榄��g���=�����Db�PN@�&K���c$Bi�S���Y��WG�x����L�c��tس\�g� �Tm������g�
�LZ��{���t<�p��)b�q]��V�s7)�P,� �]���p��T����ʋ�?�FP�lqe��q�j�Uu"*Ť�,͖�.������|G�b��NSh��������Q�L��D���ަ�9��pr�'�C��.�#�Բ��W�(&���*@�d� �����o	I�
�W�o-�DI��#�*����aܛ�x����Kb�~��� ����Zȧ�h׃{l�0���d>����j�F�^�~��n�(뵿$�� ���3�wg4*J�3���Т{�E�gC�M_e��Q�Z�Jڃ��|�T�1]��G��N�%$Y�.Pw�Y��"O�C�Z�+� �R�K�/oV�8�L;a�L�*�{�$4�:z��1�f���(�3w��(�3y�M)k�Q��T�	���qb�N�������/\xV>���%�w�N��;�J��#Mӣ?ɠ����πH�̙�j�Jr���pX���J���t�uo����=�ETV�wmH�N�X�J|g+77�&۬���^b���5���^��j��]lc!]�Jo�S��FXP�2��^X�s[r;�Fx?���c�=�݌
e�wJ�L1ȯ�?�{m�k��ğ���A�T� ������:cb��g�N��c�IH}�_�.��>�:�w���\,T.�		`{�]#C�2�{k�y��5п���p���'��V*��Y#v��P� ;A�@��b.�u��CmQ���=��״)-v�4�D�Ml�V��%-�p M�vA(eh|��D��^������	5M�N�r>k�.��l7�?=��UHۉ�ݍ(���u�¬�d�n��)��CU�G@��]�Bp���2tr���X�GC�te����� {�H���#��=�#f\��M���-5��kEe�l�J�os[_�#��	�B"g��i�E �+fu�R.����\-|v���n"��>2G�f&���S0��R�=��۠�����}��D���2x�Z/bH*w�N�EB��(a5S�.h2IJ��ҥ�b�;��à�m$;�&�:�����~a=�ta��l�_a�@�2��5�S��k��<�"6���	ke_��r�o���4��̨
��
U*p\=�D��4���O3�����nN�m$�]oM*{62����=`�*!�.!�V�U��m�<(c�ӹs��|��5�{^Cj6�։��1����(�(צ�����ں~����A�c�����҅f�S�M ��N� ��ߦ�Do�sx?���Y�ӯ����8*�3Md�u�k�zH���#�FLȦ�CَZ ���ҫ��©�Dp1>�Ӊ���
����1}�&#3�4/wb���[�'��Q��6�>�V[+�sTjK�U#bp��F=��F|�ފ��?f��u�R���M^��@� l�L��:q�1��#T�,�y�f���_��B�(}Źi�k��>{AmN`�[��aw8߰G)$�Cm��q3���kb	˫4����O���Z�,0 fѢ�us��EowUps_d�	NOL����	E	�UcК��Lu\��)��qKl���x,	���еQ,�V�pg�C�|�����j1�!�*��aZ*�@CI֎�6���lb���:K��q'���=ƥ���|�!��WR �\���V�����+3��(��ZPǨT�WJj�I�n��i��ؚ�.��,��~k����e�"��mw��.h3�67���s�d�ٔ����Y�Ȍ#�0[�3��B��0m ߋ0fk]9m콎B�~�_U�mRv���9';�����'�FN�	|?�ۭ�U���L�]ᙱ�6ji�~ޖ�ͶjY)1�=�i�i�EV�fj��K!�ߩ�+�o�]�
�����g9�H�7� ��"9?���h7�6��+`iQ��0@��M�+K������[�L9Y&�;�w�
��F�$&���ܕEf��>�b�XE_`���CLi3���)�7�[����6��+����V����QK��J���@+8�������^�EOx��� FR3���zs�G���!S��.�)� �[Ҷ��j�\�t�[}ԽZ����BI(�;C�O��:�B�]�p�L�����e���((GqĆ��9�dؗot�:�􈨑#�9x?�A;�>.v;xς��9�KV[��M[:��lL�_�<#��2l�H.������5�	*Xb�RRb�"1*H�x&��mT#&��u�-n[
�{8����W62��ֲ�3������BL�%����������pN��jS�;�~�U�Hy.Գ]bo��H�i�M�##�	��q58<�'�Pa�Ώ�7#�Ԛ�k��t�(��-�Vo_K��5�vr�U_�5�����ӎ'{_��b��ð' �>gn/��b���~[�=��(�u����>=3������`�����������jL�D܉8o���T����*�M@iA��*���=��B����;GuJk�ɝ,���d�ݪ���<	��!��*^ȷ29���K�lR�d����rVuD$2gM|$� g9����fa��o� ��� _�L^EOg�h��F��>��:[��R�CPYQ����g5	fdmV��op*�Z9�N{F�'�8���)�VS����|^y%2���4`җCܖ��L�X
�s{qZ|o���`�Pf�w������HO�0�W�c�����bF�"����ο�|Jƙ��Q�L��Q�M�C%=�W5*��ŷ�f��N�u "�'���,jl}Z�~�i����,�hd2���D�F)�������n+���n�W�_fS�zX���w U3V�/�Ɏc�����[K��l Hcp�W��g��]'(��4N�RR�8�3iC�<���G�ȎoR�T&����|	?=�Z����DFRB�"x���[g"�a�>���M��\\&��p�����
=,�q�&�9fNK�>y��U@$�T�<E�A�.��*.s�ߚـK\*���t�Y&o��'nXSCTè�����ˡ"V*��tg�tUHeVQ��}��Ď�5��^�=u�+:�Lv�و�����9�d����M���ؘN��A�"��λ|Q���v���:���Aj43-�(u��4۹�=�
�����WJ����"�&���ْ�׻�V''y{t���
�U�� �F0�qh�� ���Z�ل&�f��lQ�q�P��F�A/nDXe��	�Ƞ֙�A��8�� /���k��u>ԧ���2z9�W�1�<EQ �cIG���'�Q�웉�c{�-�Imu�[�j����?���%o-���Ec[��v�L��[=|	��,��Y�Z;��j+��V��b�&F��F���_��LF?��S,:SI�fQ��>�â�,�tUk&��J<�{�Ԋ-�a��!r��HyE��N{.Ŗ*9�'�IF�v:#��Kc�@+TŨŏL8~�̓��at�AK�����M�P��q��_[��M��u��ĸA3z������ﶟ�(*�Y̎p���Ǯ�_q�ʽI���b2��Ov4��[)�1��p�*����Z������-��&B�|����\&�L����K��"M��Y���4�Roz���}�]�u�k"��bn�-���E�͵������9g̪��?Q�g0#�C�Ȩ<�ehB�LEOk�E�YFpe�l��d�KA~���N��EZ=��:�������O�<�h���b�ǲԴ~hq�q��{�LqP��O�3�Pm]��j � ��u�_\]�����l�ً��$K�w�ˇ	�DFp���HT��t8��K&��*������6�D7	��Op��H�h��趯վ�B%ӆ��uU�RSk���]�*�QX�bb���I
b
Bw��x �����4���w�W�Vh=l�H	�R���n��L����:$��ܣ鞛�/	��ڷ���̙EۑB�ڙ���ύ@����.^�}d�8f� �n�k�r���p�ֳ�z�_{��2{�qy�}�\+����q� |���8l	p�A�,��1�̦b��J1��D��L�6f�X���l n��񼰊�9��#Nic-�S;��"Z�y����"c��8ZIW�2��I,O��:�A���~)9��}�����
����o ��E��F����{BG��M��&�o3���/1�nB6��ֶ���0�\<������w%�O�9�2���蟹j��	���>K#zJV�)��|L��8a%R9_���FÆ�ƥ��\$w��d� ��3ynr��Vk���]��O��
��B�P`�k�e&u��N!��~���(��6�犯R�k��Q،�Hٹ⤈/h�r��-!���tarmj�R��5�.��������ť��:ۈ��Y�ͤt� �{)�F��<��,���3�b���X��f�iDao��Nx�k�9w��p�-(U�ܣ���2��x:��`��I�:\��_�1P��Jv=�=��e4e��P���l8D����D��h��2mۜ��q������p�����p�����tj^�]j䲰9dc��xLQ���\j�7�G;��M`<)X C�2���w���٬ʰ�s�G��/�Uq�R]������lɣU���s���c�"�(Mw�K��!���ꗜO�]�]� �=k�י��h2�eyL��X��/�%/0=t��h��	��ۡ#� QY�ӱ����֦�P8V��]��|6�<��j?���j�P��:X�h����8Ξ!���)�Bn����|6��
ѵ?���&aa����?(b�pnR��܆:8�>����RR���1��#^Da
��KS�����o��<�l�5wᒛ��~bSr���"���'b�h�շR�0j���[�櫋�Ϛ�
�jq	mc�
Ȇ���>8v!>0��K/ܓ$�:�_@�p�|9�|l�\ā���R~\��Ѐ��;|��K���J1K�#x5��i���7Nx�z:��hg�#EqfP��h�ϱ�8����P5��>?"��n���At�~���Q�9��[��.�ʭ��A�-'�05}3^��6��Ό�� }�ś���m�I����Sہ�Vzu�ѕ��8�@�"q($��9`�.��}�S���AGۼ���?�H2G.�_���b�U��Ɓ�_hgs��VPj��O��Qj��&�"%�)��ÁR]l���(G_� �b9�5��>!f*ެ�'�x/�UG(�x$��>Cgo�|ٶ/��7)'g��B�Y��yw ����]���ߦ\��:0����\�w<�Aΰߞ$��B
䗃`���v��(6���W@'"��_/[\�MNi4 "*֕[p�R "�C@�	"-�a#����$Ŭ�,2��h�e/v��m�󆺌��ZC\��s%s��l=#���E�F!H�r/_8���;^��=~���̀�
���c��a^��vԑ%��?왝l�{��_� �7�*�;� އ͢o�9.����=Ht���5�&ژ���Fo:Q�O[YU���	�;�����[�&��G��AY$�(��i~�%�$i��ዻ���Қy^FQqW����7�t�E�11&+rK���=���{$��D���kH�%AO�O�q��;۱ '?Gr��������\�'eD�aA��>��x!O�*��%ێ��k��ǥ|7]"��j2j�E۠�y(�Q�7���l
c<��߭Z8���l8��˝Ϧ�خ�}�� Zfe{>x���c@5�J�q@r�/�\g�j&F�����)|K��I���dʎa�˜±�ण�3Rئ���8R���s9��|b=\�7@����8�g�b!�:O�dM�g�@Ch68A5U�xP��$#�T��#Үg�|�l��r��9u����XS�9��X��U��l�1��B���n�H>���)T�j���P� �D�l��`Ό�Y�aGS���=���g=Oo����Q�N���	��~��k}�	ǎ�U���.��K��3�y~`�v&�����>�0M5�%-W�7�
���vQ]Cc>i�,F���2���A�S���.���j�d0wy�"a�j��_7�ox��Tw�ϙ�0�����|���fퟪ5����l����-�x�f���e���@�p���� :�&�Qx�Z�?�~l��q�UhYՌ�5�<I-���l����S�}�����Y3���)B[�� ��_:~=;[֑m�A1�A�1��򢙄İ���}�s�H{�5�P�+uԬF��mo]a����S��
	R�~ 4yRw�ɸ�Jez���Ӛ9��F�Z/{�&�,���*�nV���x�B-'P.���~D�v��2�b�k�w.��i��Bm�+߇2q�t�lx�}R���.�(~6Л�jХ����(.=hl�iN�H�EiIS%k˫v� b]ٜ���ee���'�Q:�C#J���q����j�8�;�ؖf-����%<[�x��W�@�ЋS�t��E�H��7q��eDe�≠.����x\��!�|�k�	e��Bf�f������^b�?Fc>��z�{ �����i�nzG���n4���h��I]Qڰ7+5�%�(�u���w�������Z��te���Fh�Z�z�+&����k	���#'�	4�s��$�q�o��5�ʢ��^ye��*�!Q��0�`$"�X=�6֤D3�4��Gx���Iho@�2���/�g7���HK�#ԝ�d�� ������YnDX7���e��-�e�5L��(Mt���u��B��~a;Ɠ9�ak�kH8%h�8 �t���mY��e*+�V��k�*��ȡGQBC��LAF���1�2�ae�0��{kw/Q��Xn�$~D|�1��H�)���D��V��>w�#�����T��P�]�����+��z6H��ʮ����*�H�+5Y����r�ǎa�G����O��v$^,L��.p�sH��@o$����d�����,�M*9EZ6CX�&v���! #z6b`T)�R�`>	m��	Ne�V�)z�,#՜51C��PV�}����:'t��^tD�)ug���=<��������.�zdO�����8���7��\�cX��!h�(Eh�!���\-�Kj^0�Z��R'{ub�zW��s�on���N�?r(��y��ډ"���_�k�K��H�;��4�=�ö����^6�/�8#pyI�&�=1�����C*��x\�^!}���z�r��`z`3��s�jc��X�Dd���/Z'����i=!}�3�nfdC�<��R~�$o��g��s�E�,m�jC?i�?�h�|����ӐX-��+i0��^�✿Q��7A(��X�o����xL4!C���b���OX5����o@��SB���{P�ko������gjN�O$"��<��:��g����@��Q�W���5<o�:ؼ�F�`��k��x":V]�Z���E�jA�f@!`t���2�0��訊HT�DԞk�J���?�d��]��C����j�������ƲmO���E�!���"Xs���)~t�� �b7 ��Evgj�
kIUدP+�!}�L�5��\�5�����,4���%�he58'�Q
W�1X{~>c�J�&�ݐ�V�C')![�w�}&&�3�
@�+"�� �fs�Al�|~��uI�b�>j_��`�q��ۙ�af���'�y#�vc)o}Bl�.,�����^˄��Xg�n��ӂva�[dt[��N��aP3����ڸ�_2㟚�رr����}����d�d��f��:3��|[���-gh�ʖ��ث��t.lhf���e�U5%n�L8��GBGsV !i�u�?=:��K��-(���L�)��@s�+MWswa$�z��!��	��Ac�y�ݷM�)&!�+��Y��x�%Tnl{':'�k�a�Z�8��
���v�lٕ,�v���(B�&:�ES���Ƹh�h����vz����9MԕXڐ��E��LD�D~i��s�<����/���%�j�5���wη����ժݣؙŢާ��}���T����%x���K�d�%BS��lIn��^���v�>����6n�a�\f�*��/;nJ�fm�ԗ@�i[\�K�Jo��`K��C-�x������E���>�M�~�p�P	,- s�>w�����UE���Q]7&,�p3=+-������	3�k-o2!GU��!��{}�~gѹ�S> �M
�A�psYa�7�Q�ckS��-j�$�Z�Q�挾���L�^�>��(��*�Ƌ�K��>�9JZ�Bh���H(��W�X���j�Ԟ��%���O UZ	�m�+�(C�S�X5ܖ!���	�E�'�}q�9O^��H~YP𥇈_`�?��D�1�٥�0��9�v�O���siW�{$�J����-<�u�e�e�ns���a�0M��u3M�\0��@� ��N�/��ߏ����j�@¥q���_��z�Ռ�T8l�)t�ɉ�g� 혋��T��9R9�g���QiAg�>�Yw�9�C�t�20�C�3,��G����I"3W���h�Z�tV�s3�%i�U��:�\�X�S�&��Y~���R�A�0_F�����/Zc���-E=]���sÔ۲e�4	�,OEw^yj^ ���NZX��O�lt�ς�Շ�*[:�Vs2N��.7�,��]�QP5��)U��5щ<���HI����čۦX���=#|w`,?��
xW�̏}��%�5�ݬq;ID�V̀~��J� �@������~[1�ۇ!D<UND\P��S�V��y��ï��K��&J�f`��̂:�v�o;��G&����w@yϴ=(Ԣ=A��CVGGy��G�%��e�b����WG>�!q]��h�Y���׹o]��m�\�im�9�����Yc���4uS#��@?)d����)B1�ޤ��BFB�:�e(ڕ!k�G��@�GoG~2	�� k�xsoB��Z˸n��K��8򥍔x���W��hª��b�����:�G�L%�ņ�1��+'�B7ѣ�����D=`��D=5&�C��e
����ni,V���������.r�\��L��鶍N<��y~D2K�n�FP�WV�9���+���D�s�4��(��|�M�5`.���]Dlo����>�ŭ��`�!�#I�G��1s��a������������/~��q��|���B�*��e����h��,�ب����8�%�[}L�al7���:��)��"lY�2�GO��w�W3�����2`� ��bp���?_��x��xgq��oCiNp@��<P�w�������[�ČzImR2�Z$�i������r���i�hny�rS�yC���	{tX!��
,��s����	Ogp"ln*��@h eq��77�}, ���3�Q5Z��VY&�t�/�����ٕ8Ҫ�1D�v���m�!���]Qb���J�skH�n����W]����x�9�m}"\N��_��w�vWxF����Y���ɿ!Z�7ê9O5K>�R|~�U{�慬-�ٙ,�q�2����	i{C�Y%�i�����ST�x@��^م�n�X(�庠J���ɝcum��OL����l�~���һY�&�7ab��$۬Wp���S�W�t�]V��'[,��p��í�nQ�k��4ɮԸ�X'2�	#_���-�!H.	#�劍s#���I�΅uþ�uЊ��{��o���`w���[����C�d�D[���q�7��(+�Nu ��Z�R��.����o�݅��S֪���Jv�����6fn�fzحJM�+�ewL	˥�u7�o�N+��﷾.i���A�"�#?r��e�"�_�.uw�`1 ��?���A�q�G��qfSi��G;���4���X�u����d��F�a��]@��ӖaZ�V�)��hm�y�ed��x��#U��caF-�j@
��n��R��)��@�>�6m�L A&H˖�1d���)��VB��u_�.��ʎ6�X �@3N��`*2�?D�#��>"�EA(��Kɇ�؛s�}�`.����ۀ�&��q�I@#�9?�ðSI��cҪ��V�jj�yv��=<c�y>;@�϶���;�S�ݏhH��PCI��q�f�5V�g_R�o}.��s�e�SU�XG�����[��y��7ㅴ:>;�X�SxU��3�GE�*�v6x�(dp���j.� �N�+��-��	� nI~���{.Q��Z�MU3&��3YUs��ט�IQ�g�O��]JѸ�!Ϭ���������6��s�	Bv�W�0>|�*��K.���w�q��u����%X���&V�"�0@��|��H)���&TrH�Z��ߞ�����J��{�U��?dO<������FeW�Q/-�F� I�I�X�M.�Ȍ#�4��k�E��IiOn6`of�&2igC���8=�j�)Ht�,����U�a*�m���}�aC�W�F���y�#~�xW|Y�����j�x|I�6g
7L)�4��v�xl���WVl������ ��c~ǲI���T8���C/%�.:��xw|�}�1eq��-�sb �m����β�`�2-EQ� �����zD���X��Ԋ��D������V5�T-nh���LFDA*�[B�&��;@�{���Oݝ�Wti���>��~��8�+���ƻ��Kh�8d����,H���Q|��|�tڈ�\�� L����fZΊ<�bb�T5��ai�pQ7�#��y��ũ�k�̳����bA�B�{D�G�Lo����^�e����k��Y*ֺ'G�f�Gl�mn����J�3�Q�E�۳��ni3��w�\��%�\jI���ߪAͩy6��_�G�罊wR1ik(8�2��p���0�y���Su_��R40�� V���)�3w;���a�z��@
p�Ch'#��6X�n�O�_��Uz!���ꌳ7c�]e6�q.��5�Z4�2y�%�4����Q���S� ̠Zɖ4�C��ۉA+J��~v}
W�%f�΃2
��`z*��<4�_�%��* q`^@Y���O��k��r5S]�S���v"�m��^)���QN��HЅ�RDP�5.���݆�P��˷~j%���l? ܲC�T�x�ݤ;XGR��&nThR��+�ayǗ��H*s� FW���@*[(d��q�E�j�Ӽ�>��O>i�0��)-����_h�J%\E�t./����o��.��JQ�λ�ɖ���$d��CȈ�6�e��ΰ`�vrr	C���쌮귱M(��U[���p-J���fp5�������5��W_�\�'����?գ�B��e�O��B_&!���OC��I��T%K'{�P E������n��������[��D�i�n�m���EV;�>��-��.��V�����>�F$h��%��)Pٽz/��6�Hj�s\���k��fmV"CPCD9�X
r>+�M@���9k:�Nߠ��1�170���ZA�����_�]�ߘ_��&g:�>���۝G����ɻ[�V�*��Q�O��А�Oa�~H�#]�Ũ��;�e.]��������C��wr��H<����o �J/�⡴�� k�d(�k�=�Sz ���Ȟ���><�*z��mߟ(�F5f�靔�	�;:��%�`W$dߤ���_�u/̭�o�9:���P��J�۵a8Z��0T����()���xh�����	�m0�?K2	s�1N��*����\'b:C!(�B�w��G��r���'�N��/'v���Ź(�Y贓�Ok���Ix�M.j�y�Sg�>=�|����1T��+ql�Q�r3��h1JT�r|�����:�o+�H�
����"�>q�s;�<2[�����~4�ٻ �ʪ'��$�[�+�7qC�Y+-�:�i��8,f���ƴ2��H����gk���N'��/�w| �z� ξ�c�;�-� �A��=��m�X^r��%���f�5���vV:�q2������������/n��B�H>���Y��7��&��g]I"�p�W��K6�پ�-��_F�k5&�7+ON����A�=�xgx���'�w'����6r�?���K~?�!
��.]q5O��ub(��f��38|��|$����SQ����0�.����Py0v��m%R�RH;o��k6߶b2���3xS��*$��F�̄@��o�OS"��`pnqg���`(H�>����.^��5r�h$H^���G�/�ߎA��4O�ڤq!%Ad2�B�G#�|�X�K��Q��Z
 ��X�nڣ��^�͗@Nr���A�VQ�V9�r�Ad�k�}0%[�a�ǜ	|����͒ui��7S �Y���O����]-ǳ��c�x)����O/�e�Q?������|<�Z�I;%;29-0��(jE���8y��Hz2(}6T6�*oD	���E�޷!�q�~�A+|a�BDùvY&� �W	[�8��t��Q'9��Pjoą`�rY2Hٔ@��PĕGF�^h{� ��=6x�[��w�p�'
�����%����#_b��{�RM6F�$od��@����oC�lyiE�7����6f[�<F�~v���tƠ�(/i4�$�%���%���Fto�:�����,n�PzmH�{�k�E��!�V���07%�O�@d vAס�O?IP��1���M���(���r	���ew�.�Oksx�B�Tܼ�3��셫��[Zu�M���.�
��-���>$3v>dDj�� 8�m��0��{T���2./	N ���(�Q�������qՅ2�Z�B��;�'�Mz?&�rl��!���sUo>�ʔ�L�}*��l!ՇB��΄���Ja4�G5]�G��[l�4צ�Ee_���_h�����8k�	�f��� [�$gɗ��Vʼ�ٕz��V�T��*��(*́�_�b����=�Ɉ_{D1 .�lS�ն�	*�+� ���.c͂����;��� bqz���^W�
��KL³ �Y�	�!5J��|�-;�c��n��r�&N$ᖋ��ߣ�
�J��2�J�'h����6�	����a�^C@�����s�+,@4�`>i6��q�5ўo4���t���Jܢ�|����Dwu~K�Z��Z��"�E	Z��� ��T5u~���¨L���Dh��������V ��S���^͜
�G�l&l�)��_[Bu��nd�������X��ٍ(RM��A7jΓ��8���m
�S/Au�_��-Dir�|�B��O�yU5��F�K6P- �B�Q
��0�ȭ��Ν���e�M�a81�2�^0۪ aҚf ;u~�5{pg�p����E�n6p��� kD��g��?��Hv4er&y��!���6��mn>��w�=j�A�x3����0���)|�#/�z6���&���ؚg��R�&�#��g��A4���F6䯢P`3��gs%W���.wG�H�	���7�T�)��K��
)�sK��qCS��c�lu�jĈr����]VG}�K^�l��+"6�p��
*�AE��ϲ�=T�Z�8�Ϲ��#ī/��^+5�~9��mm�gj�V�_܏��Z��ٍ�����j����~�����ʚ��.�w����\�;~�Ƭ6����� p��iNY<撔����JE�j!(VQ�Iz�@�G��TĈ`1N�8A�-��\sm��;������W��]�%l(��,I����B?��r``���G tT������Y揘��ME����zX	��9�>��љT���	�����&�����Z�B�R���0'T��9�8o7�,[@����F�>=���o�����$�U�TGi��uo�o����D\7��w��i���gG��G>X� 3���b�V�w�k���L�B����PZY�'�[�6=Z��ϢsG�v땲����j��F�@��YN0�M��
���?�/��GtO��9�F�����䂐e�	�Yr#�I2���@���|�X�/p�,W�.a8催���� L���%v�U�ﺔ�ho�E!�xSU|#r-�8��z߼* ���6�|>��U�r%Ja3�����6X���Tͩ�0Ѥ�Su�}�P��j`�p��lJ��Cާ<����V[F7唎��<l_P��H�������E���x3����%	 �^���ZF?�Kkiy��9JX	V�,婦
ȼB0�	K]���U�Mf����3�t�;����Ki�M��V,�}��%�'!���E^�"YҔ8�fTچ����)���� �3�L#^�
 �S���[�����$��9�I��n�6�	��CyʈfÖ��?������-R��퉊��j�}�&�:)7<�Z3oJp�t��X��dE�)���3 y��"��:����9�Ẵ�I�-��R���uܔ3�u��J#��
��x��x )�5��z�&��[4`u�Pv��x�#���ٶ�#���*�=��>FG��[����7YEI�������ۆ?"��ctu	��Zv9?��m�A��Quv�Q�<zp4�5<xb{��焱EB\!g�

��C2pLw���?�U��4i�R������Dj�	i����� pr��ty�'k��[�Q��oQ����"O��-[Dx������v҈�e=�x_߬�^sڑ|W��#:S�r�	R�X{�)U�\�  �MIPX�Tds��9�8�P��gG��k��to-�i)���6�d)q�N�+��b	�&g\<�2�Q���w9IAe�lC�e�~��$�(JO���e�-;	䲿��Fv)\�p*a�W[	D5܅p��[�������9�cjR#�v����a7��S0�=�΃�(�w�ά�?Q����&]{�Z	����T:ц3scߛ�AC��!�_�,�-���I�-?������+��[i���N�$��w�o�~�����|JY�s��x_qh����%�3��O� �ME% ~6ACՇ�ܝ�u5S5h��4�[�]B����\�z�R��3/���du��1���1:.� Xv�!"�ppY�p�j��9��M�"eӫ�{�����0�ˉlV���-�����}���<5>�k��d]���qa���WW.�R�*uh�<[����.��*�dHoWo�q�jլ�<[/��
���.
3�97�LQ�k�!�W��BE/�PFY�$�L��1��9�WMR�5�%�%��ᬽ�ֆ䭷�jt7�}=MQ� �#�"n�?�9��1)���I)e�w��]N�y���xe��"*Hk�U����:�F<���`�9r*\>,6A�&�l!HY��ԏc�/��mS��vG��Xz��3�b��?�����	����O�����ny��Ⱦ�W���hm�Q!��^�<��l�����`�<\\C�$֢t�V��_ņ�]�<J�@��!��_�%�7���l�NJ��ɏH�>���!��h%US�ZL���Y�� ������*%XP�AB��0�0���) j�RXwak]lC�>%��ɰM�ET6:h�	��gLu]�3e`�����Zod��Ë�lL��n�l�z�w2�?���v8�WTb_A<A^>�=�ݰ�g�x� נ��IHU��W�� ��F�c|
񮬆�,�T� B�=���G���-@�/E�����������)���E�`����{4mkР �#�W_u�]�'r�(�3~�bU�7�~�և:Q�VrB���b����,[�������X��^�7�����qlDM��")F�<�
�٫��<Q�j�|�CD㠦D���>����O�nW�H����������4[B�Rң��;��E��&v��'8�)�	r7�� �+Ϙsw���h�m��y�}�w��uE5�.���S���G�J�C�E���0���_��J�\�_[�\��6���>�3�U�����-}\H,	ö��c������ѓ��=�ײ	���T�_�Zʽ�@�0NMhHBG��%�I^]��nw����8�}�rA��e��K��sz����z2>X>%C�W��͢��%/Z�ӹf�J �.�����+�ņf�r��UB�mi�^�B�t����F����؃	�8+C�Apmz;\Jn�E�U�k��H?K����-LY��§2h�5R~��&ߨ���ObkH=j��t��Y$p_��i:Nq�������e�ă�V!�B�׊w��M�{��c�F~�:��OVT#~��l��R��s��i(ΘQ�������R瑀BEe�p��:?ɿ(v��@�`���(%���-<5�]�\�'������u崐Њ��?�i�U�v@���u_j&��+u��ݽP^2�5��,H�;L���ژ��K0���ay��VP���G�k�Wn`En��%��$�({YM�`�ೋ��o�U�@�,��I'��'���}7��.�����'\'����[%:��^���S��?��ī��%�sؓ�>�����E��[eW(�gG��7�el8���ta���Q�ۙ+J���q��D��^�1�.�U� n�g��3�&�&�
�	���pcz�"�$����MΕ��XeN�ն���w���������"#���?z�,3[��W5��m'��b0�A_B��)��DϬ�8Z'>yb� ��[ur	���	������sOV�Z�ڰt�`���X��Ϋ�F$e艂��F�	*K�sp�G&�^��'��$n�F�'��������{/a�D�|��so4sv��Z���W~�4�FC���@�����D��N`�M��̾��N>8����Z]��i|f=�"k-��O���ta���v�D�o���Fdu/c�t����ڜ�a\�s5:}˦�w� ��vZ�خw�12��A��B^F�P*��rn�Z�7��� 5�b��$�c7Hx��|U!����T�+V�״�+���YL�Pv�¯� Z���Б�K�������j%˶����hO �S'k�촤���2o�Q����2��B�w�q2�(�Bv��>'|�#*L���7o�����I�`3a��R���x��Jb�unL53K��Դ <5z������R[|4�+Y�T�(&>7�:�1^Xt�����q��7�״mD$ EI21��ތ�0��6ws\".��0y�K�D8/��ҥ!�'� ��[:��e�7wz~JM�i�P=&�s([�AVJK�)��V��`�q��A�{�o 8�I�uM�&���4�)k�4�(tf�d���f�@�7�z�Q,s�GQd�,��>˵� W���3=q�?zI	W1	3/�a�qfԝ�ݐY�y����\�-I ��+�rҨ���ږ�౺ܙ��"ך"�ٙ lx���agW@0y�7yNe��9 b6��j�m@��7W�l��A5Zy2�˼	a*|%��"Enm~�bI5���!�`{����S��z�Wȴ�]ѳ�7��Rфo�S�yZ�WU����jx Y*ZI
�|�Iz�(�N3��/�>C��j�H,��ޮ��wŀ�0�f|78���1�/� Vdm���Oⱖ���������y�ç@�(�GG$�0��kY�<�)u�J�>펿�!�)7���\��	{iNYЉ���#��&]���	,x	׷W��B����콴��>�����vӅ@:i�v�c8�g�� ��u��
S�M��|2��jd �$��"b;���>�f���;�XM,�>A�M�ͭ��fx�wOH�'DMd�������'+auDo�-��)&E�_���V�v��O��l��I���T�>�E��s�7��b(�s%+��c�r5�v��ʋ�+��ƞhf1�#����pТ�F�B�����lY��d�p�9`t;�;O-�[��Q��vF.U�<�}E�{��e��ܾ䚻���2.gZ �'FK��A{�^�W�#7�4r_�__TS���U���6��%����
g��$�%��i�&9y|ڹ�
�5���E3��_�5�E�%���b�%.@������L�/͠��0��7\��w-3��oO��C:]JI���|3L�/_��yr��g�A}> k':u���ϝ��41���4vQ���$�gܲL�R�d�ލ~�^XS�x�H�*Y�h�@����n�M�W�)����~�4*%�'�
��A��E5z����su/�*N���p936�[�5�fb��Q��'u�mr�޻Vs��%�����;���8��%��r>N �Jxuf��tpc>�駛�&\����YB�A��p�3�����m�T,�hb��8��.���x��[�e� .Y�s,��o�/�ñn��O+�|��9p�E� ��T:;�e�D+���Qi�4~㏀�x����vb�HkH������E�,����; >jM��b��@��t#�`=Cmɰ|U���'���?���]c�@ �=��Fk�)Lpͫ0U0M�]_;o*�J�_��&G��,���9Ǽ��;?�X���Q��2�����bׇ�kt(�R�xq���t������xp�
ш��9KjC(�IO
�a:J��t��*^R������Vvh蚌�"Fݵ�^�չrU��	$Ж�Fsf3�@b��!!�fB�D� Κ!g�Ѱ��{M�-�jW<m�E^a���f5tᅯbjJ��m6�+�b�)+��Z�`
')�c�T�y�+�����&�[g����a��F�O�"����G�8E� b�2.�!��(�O7۠3�n�u"�K&�#6�9ȃ�	�Oͷ8׶<���eľ�Doxq���_�kMc����u���?��WR�9���@Dpfǭ��e�+�g�<B�.ӭm%E����M�����U�_S+gOD52 =/���"D�	��nQ�2�lM�cu� �e�"Q�M^2�j��Eɻ�$5=e}^���޾�G'k~���7���(l&K�."4)΅y@�1x;+�[/�g{�x�$y�9C���)�Wt4oFxt@*�D���r߯y�"�i��Imo����F�>}�og����	j������0j#�驲�iw�Q�RKx+K��?E�Ux��<Ϲ��E���3���#W�n�܈�;B�*�9��#�t�.ux�d��u��be��E�)@����l�S]��I�E�J�/e�1�6w��Xjb�G?�TM;�`�tP�U�S��PXs���=d�=g�y��X
�����4���{#�4r�D@�A�,�߻�p�6� ݫ/�|]���У��;��R���l��Ucwp����~�N�ov�����(�@u��խq1�M�^�^���i��3u6١{|����h��36�6�_�V̖�V�Gnp��cXﾌ�D�=�*��Y�f�	-�*�l�������_}0��s'����و�T�������v�Υm�~�m"9��ݳ4r�:紤�#�r��JU�wdT�Y*���<%�� �c��@��ʰ�]���4b�/��|D��&P�I�{�*�'�O��b�5׺�</w��/���r󻕆Ý2�N#�l=7��?E�w�OT��%Xm5�u�Ns�e�t�����׵s6�Գ�,�3�A��&�[��5�]Q���dg���3����V��FH5�`�i��%� X�O���/:ol�'zI�#|An]������㯨�:�k �5��I���*��BU)9��F\�-��nإ��!�&��4�+0��3��7�?C�)X��*���4���z 7�B�`�9NP*DNf��ߛ"��:� x�I�e@�O�������	\;F�#/�P ߹�6l;Xe������,zD���]��,1����~���
IcL�/`lJ{�����0�]�XG�jeUf{gFh�ahD]"Q��6�٬�R�U�ڣ	w���yEŏ��]��Ӧ��D��"�E�x[�#@�����/gA/Q�W8��w������5t��g�(�%�%�dl�N=;)2�<nH�}N�����Qs@8��d��j�t�}|Q���j�^�s�gAV����cT�~hS�D|��hEe2�"!Z�~+0	���D ��]S-����3���Pv`��+��ZH�M�aML-	`Esew���f����
�.��~�c!]ٗ��-?WLv�GuN�q2���Y
u�)"f;�i�*8W�κ������ R-v�z\tOH���$KN�pT�섁g{�>5���a�uI)n	�-��6!��}�B�1��ú7x�W��Fa�8Z�?����j��݇�o �e�G����{��]Ud<�_���`Sq�k�o~p�]��#�cz/ۊȸ�u%�uyU�],q��+g<�姬%>0�'2�DF��,����/��y�\A$�q�������@��dQX=M$G�ٙ��[�ȡ�}$;�
/�\o����J�⤑���Z�mV����x�G;�S�����6q���u�in�ʙ�<}�*�^`x y?�R�l�탫x�Z�D2|�迺�C됇؟�E:��c�~gb�2@�p��H���X@(�9�G��7���e�AAa��=,Yؽ�b���k�*�RZcC��x��M/k��q�-��|�%B?L9��_9|��\�W�k>n�rg��b`oL�Z�L�S*XɎ����|�3���|@�l�����l���b�ƽgК�]����.�R�90!_��XE�a'ΟY����: ���.L��o6/@nr;��� ��ѪE�5����ۖ�������Gp�%�2%tt��H�1��mcU`��h��3������@�bh�������L"�D�
�y9Q�9�h��X�p��1�g�J2Ui�5�^Ġ��N����3���*�|O-�Z��b�#&�$qwo6�z�\?�r���(�;���D�wB[k�F5�\��H� ����X���B�9&>��=��=\\_$��&�G������E?�-�m�I���ڛ�TL�0�ع��5p���P��(�]f�����^QW#��|x1_%���s&b�bG�8�̙��v~邟=�� �um�m����xG�������T7���R̾'�q��4
��M����jq�DS�7�>ި#4K�2�Jw����)нnK~1z��^��_��Ћ�����T)E��t�һ$��OH����y$$c���R�C�v��s����р��nM4 V��÷2���g�m����"7�G�����]	�v��^
!/��:�춃\��TxVh�C�4���L4$A��qSu������+�@��_cj�	�Nz�jk' �F�!��ͷ�i�F�������~�$_�1�-M��P��TQ}���@�7v�s\Oќ*��I)�G�Cl�����2�=׀%��7ٽ�~9 Ô�<'�$$}WD�>v���-Yi�=Gi}�"����P��W
���k�Y��:�������H�p��ti9'kH�@Lr���`m�_���w0!�/�Z�y�;�|X��Z�P�_��UD8V-x]gL�@�A�t�ŬSFU�`(+=V��.``?��SX��������T3�@�Wl�Gmk�-�C����L�)��|=��yv��)}�,��	m�4T}v�V����hI��B����`��3�VO�iy
-7,����m�+-ze�)a�}a|�z��L�W��G���/��QA���~ =�3�8Cκ���.'/)lr�境N%���^5V��s}��~���Ur��K";\@P��1C(ZF�m���U�ڈC�@��VF{��]}�	�$Z��6�q	7<��2�1~~�X�_���=h*�4�_U�@�+ZW%��	8��ɮT��=Q������u��� ���=����
:#k�����t���^1"��)Ïd���[jCk��:��W�t�8��cx4��Ȗ�#t-��ϼVj��'nk 7a�"n�?%O`��eK��Q|�����W��� -�rF�ַ�
��5q;�TDbL���G^�nF�6Ů�Yh��S/N�E��wˣ������ijq�a��i��%��Q=��#�|%0�ۜE������!u��u7BE栓Uy�ظ�Qk�[��k�7��nl�KXF�4\
Uvc ����)��O�;�%\��ěX�����CZ��P�
7��V���?�2��_;�7�Ͷ���1�x�S��2�V{!��wڮam�d�
ݢ��3���z�RE&K,��O�$�=/��0o�π;=~k������L��Fr%�����fE)����Y��+z����S�4n�cD9 <��}�,��C�~��ל��VT7�Yˠ����X2�{g����Kq���@ƞ��]9 �:���L����[�Y�������Gd�]�1�P\,�����✘���ZW���(�W���7r/9+�['�r���qp������9�N=<h��m����2�pqQ���'�W���K�@���nF��j�n\i�
bV޺]oQ�1g�/�rT�C؃�MW�L��2_xnX��N�&t�nux�TC���� p	�T����rÌz�t�u:b��D��v��cH�w��V��,�.��p�1�W�Ґ����d�et6�Y�*\�Q�|��D�a�^ ��\7�D�
˹:b�6��uD!.9j�&y$)����)ICK���$��)���뢍�_�t�ƨ�\}pv�P�����B��TѦ%�s~/�.�&R� ���}��@�CbݚD����^'�SM`��uZ�6��+bU��O�J���.p����%� r������3����C�P��Zq2.xa��[��:L��q�X�(5� L�,.�v����)�9I����e�+ǟ#�)��$q]�Κ�R�qժ7Z����~�D�y��Q��E
��,k��n�m}�0����[AR����� ?��7�>�1-S��c�.e=<��h�CÖc���1��0��ڋ�c�O;�o��.
�hC];���ts%�/Y����Կ;�<�-��a`jw���+���DY+<7ٯa,����r
�������H���!��3k Ě�g(�D�����EM�H}�;5G��O<��$=��^]�[�r�ي=�N
9�r���WE����vD4 �;�������grn
?f0'^�O5���	I��8֡2��R�O��B����h�+*�������J%4�s�-q�YXR"�5�#�xzn��y��'����������@1lT:�����(ǘ�2��M��D�����͑��Ue���1���T�6��x�dF�<�H*H����{�9F�Χ��k�>	T`u��*j�>J	�$8IX�|�$p��a�t-��hbU>��� � b�"������W�`��J�;��#o�uCC���?ɵ�.�֠���q���~�p�����4=J��mw�c#e����#�����-#.�E��t�"�u��E�n�_��\pAC��^���f1n�gC�3w�)��(��'�)I�1+����\��.���_Ź6��0�t�x��7����MoGYp:���\8!��f���}�s����O�:��-���E�o�_�����#�º�>WI�9$��aezM߬��@X�.f�-��\_�힆0,^p����l����k2��ߓ�ZC�^��	5Mu��)4����"w�Պ�e�qj���PF��#]�,; ����1S���/(����-�!/żl�&��f�V�ot���ރul��xf��|u�We� �g�L�K��
�H@j�s��2L�q
b/�wc@�~T�j������\��h��r1ɢ{�^쫕4��R#���7�C�wI�ڻ9��r�����8;]�t�{P�$$���Lb�Ò.��ms� N�FfmΏ�g�K�X�~��=��A�g�-_���U4B�J��vJ�Y�-�<P/ gǁ\RcE��Aß���/�Ὤ��ǘ#�`� �gI'���(+���ߣa��84�|N<*��>.�^�j�R�j(L7f]R0��;��V ����$҇Z,=�q�`���
�o[��H9ӿX�܅�A2���<�[Rf�tmt���C25�%��w�
����	�w�
'��@�:�e�]���7�(�F�|��R����Ip����5�z�z�� 7�r"��X��w�⮈�oz��k�=�£��]�L��%����$;!u�8�mo�� mU��"軫Ҫ��v���7��N�����Gl&�� ب�RAŕB�d�����fa�$��?����-�h���?i�	�C���b!q�K�����I��]�P���A�ٶW�d0��IX��8w���/�X2��wpW���dy��?61b���!>R��LM�
�k+h�u�����O/�WWR�N�G��'C�#�7\x��xn�Ǘ"���K�:�����/�Β�
C<��l�z�c�,UU�����U$�A�W�;nZ��rꎽ�Q��(1��le-'A��3s٫J�,��Z�{�_W�!�˪��N�.�J���}Vwh��@��dr�Kpm����j$����� �KS��d70�����2��fnE�h���\��>�����g��i����]*z�.Ϙ�߽q�[�d���ar���W��tf���Ns���vTz�2���V�C���C��7y��-A�7$�����Fe����U:�r����j���]k�+�
xw���:��9F�L͉�W9��"Ü)�F��,� �njH�Y'0sP䭽�H�Z��M���"�F?5
P�&��G��Uw�$H�E��9?����d<-�N�P�N�ds������Q`��<lp�q��1-W�i��N��[�k�tǨcMG���9�����7O4�g�"Aj3O���W�z��N��b�k��kh~B��ů������2�Nl,�����D\	VDT�G��4��#�r�:��:>@��=��,�]>��+�y[����΋��~�
�-��UB#m��n���g���7w12��S�v~7�w5�
���`n:�#鶹g� 5�^Έ�g=E�yGO1h�ne��Hi���P��������F�g(��QG�8G�R$�:��MY�׃-^��^�!2Ŋ���i����?�0lt2ƞ#(�������r;��F����SDs���%#l�n�[��W-��������I�-�m9� �����a�l����n�������]p�c�v�P�H�ǼaXU�c�;l$������AU�'�/'���\	�A����$�*$����r|���NO��f���wJ���>�#Ǒ���*�m^�r���mK�{M�1��8��H�y�rdX�}�d.�-�e~]�K�/^����}Hc5�b�ǚWX��Gx���j�v"[���Ȗ,���_�Q:��)i^6Ը�a�^�Z[Пzլ��+�0m#<ҵ�#{+��=!H+Gy7�Y뿊��{��8|;�G	�S-�|e�>�)m�+}�'	a}	Z�$pU��1�X�mE--��Õ���1ۑ�kp�ͅ��E5OR�0[�H֒�Y�	V�/5�ʕ������A��r�0�.�	7c���he21EL�jiL-������c�[F{4�S�n�{?PΫ�����t����+D_�P˞5[�D�x�㶊��t���ȧ&hZ��Q��h����{gA.�Z,�聁8�&�
%���bi��C��R��]:�ٹ.��s`�QjtX��R�g�V�Az�JkMF�1����R%J���=�x������=E���Ę�򊻪�7�`5�=!Z̍Uk�>�����fT�@c�\St$��s�NV���礳�Q�5e1��ʪgE9$�x�������#_�'|�X�z��my�9���U�����5D�k��Q�T9$FZ�삇h�醤#�D��<m9%cX��ʖ�����|�{�!0�C$#� z��yO�=qxDe/r�����A�0|V�;v�(�HV�A�U%2�Y9��S�P`�wC�O��|�N�!x"�����<R��j�sJ)0�s��G���D��΂�3V�k��s��VP̦��U0����F��-%�m+���j/��m��5x�����#2��zn�V���53�B��J�&_�:;q9��/�b�-��Q���q1<P�Y��/�f��$/U�������|��d���u���P�[>(݅Jn-�h0g�U���ֿ���X�61��0�}��d.�sc��݂<N���c��B<	��tPG���)$��5%{{�e��dX��\�H��;$��A�PCF<by�,��=R�eŒ�;X$6����A3>?C��@ �in�]�ʋ|����ƛu%�a�N?s_M��P�qR�̈�l�z�ht>%^V�����̿2~�05��)�Ǣ&��L��E��k�It�4!+/)�}����.�:�-b �}~|�
!�1�ȱ���Y����=�r�y�;�'�-���O�RU�6�O�c�a�����A`Ģ���<�*斴�	�!=�~}�%��b�_�5U�??\�J0=;;��	�������qT��!�c�]'?�4*3�eU;M��!�%����W��A ;����&��AcT `�P|ƹ���)����L�n�.�>}'_���",#S|el���2n��	:N������ �{�|=N�u�)#��#�4�>D�D9�z�@&zW�	��Qw>״�e��5��dp����������jn�Ѝ:\�\MÇэ��Y�a&y�L��X'�F���ny���/<$}��$��E�ykw&,��v*LJ�R������X!��m�iT �Ƹ�9�%�J'�D4Q����EFG����m�hwL	R 3�-$���1�7�Oi~�3sI�c��'�ʀϤ��)���$�d�p>��!��~Ru�~ ��ͪO!}��p\�͢4EP�a�'��It4�����5���\]�k��c�sbrO��Sb�|��Lx�S}�XR\'��!�/�����wo�1�Ώ�򨀀S1uQ�����
����2��MLjf܇�yW�]R(�jY'�_�+��^�+��o�u�\d��<i�ID�������wH���Ñ�5?�����������p�
��fXG'Y@�S����#=
,c���r7�� P����|�)	�g6���4k������"�1�e�ƍ��t6w�bob+�v���Poy*X�*�| ̐9T��B�l��4����£�Y�0�&uE_�?d���[w��*�q/����5A�L߭��b�oQJ{�xV(4��
�2�C��vvJ+8!��]xm�e�f�A��\��ؾzD.cq���k,��ex���]u�%�ɞRQ��t��La��︝R�ȉ�T������ޮ�mD��'��T�.p;�uh��e�^_EW�xz�#o�pC;�)�T��AA�> (L/�#����$Zݷ� ������+�5�~�n\X'/�.[ 3���{�I��s?�ᕶ�[�!dh5��R2��PQ<A���
�0,��RR�������AC\�����K�����S̚�������o�j�j��b�&�'���P�;3<B9�_�$�����o��Ƣ
��oQ�YY{�ߔhaj�zRV�f$cͶ�/~�����h���FCg�?�LУ=��^d�Df�6!�T#"�/nl
�+=�<�ʵ���A@2�"�eHY^�)v{2.�׏UQ,f�-q&@����B�g
N��H�%�x뗞
V���uۉ���h�Kqk��C��]=�~���ԊW�[i�^�ZВ�ͭ�eS`B�h��8�]��敜�4�3UG�D����#P�&�E�vD����b�����=� 9+��˭���׶�4?~/pfU�E�n��ᵐ��D�q9E}V�S������$M;]8;��T�7��<~R�T(�E�j��~|� bzw� T��i� 5L�{�3�^���0��Em'���°�{ ȟӲ&�hsk�A'��̴�ڇ�ǐ�ً��ͤ��7��Gپ▷�jd8<�S�-����D8������C �M�ރw���x�N����a��V�t�Bփ�=g�8F8dFb���^���O�Lwb����сK�|�����Ô�"����M�\����|+y+ٲ�`I�!U!�C�/���cF3!�'fU�͉ݸ{ �&9M�*��u��54�`�Xle�.x�����zӥ�*ݴ���f]�zx{b�}��QsvĚ�b�B�s@��~	�ex�n�Q͋db�t���5캠��
sj�4v�8��O��S�����;��#o(k5E�#Mt�.8�%���#��9M��]"|R}[��,o�i���	��1��ܼ֒ƙ"˚�8���yCJ�vU�����'-:ZHolݗ@d�(�ӷ��4�}��Ց9�4����ʙ�R��%�a�0@����ui��b��K���Y���o���j����������u�ӿGU����]&�n������Q��Z��"kGݱ��LS�d�|#��5�|4�������V�a"��a�/��X�t��s+N�uNL��-cԃ?�I]�M.�ϯ-"��7�l�
f�e�
�چs���S�gT�d�,��9�Q���Ub�	٘BF��U���X_�h�j���P_�ķ2(ź�l�9��=�qB ��{.��D�1'}���N�p��ٔ-_pc2������$�I��|����1�&�J���%e����^����9Y-�z!��41��m�2����rO��+����'e��m5���Ď���N$�q�h�l��E��w��Ί�(�v:�Dl5�~��F>j�o��T<���ۨm����0��KmN hnO\65��b���|k0�C��2���_��F�����;����
�ݤ\l6�`w����X�g\�?��{�+Z�7
�L��M���ҿ*-��:Nҕ�4mP�gRl����+b��rP���vQ9�6�~����d�z�~��4�����~�1��BƱ�����8kf�˗H��Wf�q|_a͇25�[8F�ٜMi/��{Fy$��ƻZa�Xw9�%�:�8͇*��M�q5uE�B��8����Oa	^�T�${N=��Q���*H����2�L
4W�
�ˡ��J�qoM'�F�\���g�Mm�&��$�#IC�3��p�5G����?�l��4-��Ͼ�#6�����rc*��\������a�V�  t7&�f��ɉX픯ɢ&�9&a���}�#z P�	�}�j���s�R6D���ղ.�I�~�������MX<X��/��'��Eٔt�pL]���s�W�Zv���P�Y�2�ۘ�'�v=�䟺0�}���ȱ��X�H��aav��
@g�)x�6�2�O�Ƥ��H+h�6���Y!J�aPP�g�D�ￕE�T>�tsT5�mAU ���e!�y1��p!H�,�G ���59D��?��/�1�
?����"�F����}]����^¸�P�d@�n��%Z� �ɋtQ�09��5��Ws�'W7�S"ԋ�k
�!���!�ktG�	�䵑d+�&��.q�Q�f���H�J*�t���o<mRos�}B5۹�[��D`�c��<H�����?e��o�&a8	����J��a�2>I�6X:�i ���xzH�.Uy�@�a��Ut,�8!@�n��W�<]�ϫ[	�J�ٲO�۠v}m�ah�ѡ/��d��N2���l�+�iz���G� }��(�J��)��)2�
RWj�_��;;����<���H��gp��2,�{�mR-�Q�v�R�� �+�S3�{�2Χq?;�C�����Q�P.i7W�2��i�۵��_���x#A&�IR��1!�M]��>�,����QX�������)�:�=�ŝ{cO�\�	ѕDߍ�YM�)"�
�-]��Z�	�&?}G7���EG�[ڪ,Z�c�؎�}�����1h�φ��� �"�
��� ?���[�ꈻ��]��,sq#��ouQ����7&��[��WG���-醧޺��9Z�6˽3J�	<o�������F�P�#YJ% �W�g��2%�;A�8r��^��O|4w%��.R��_4I��3�b :�6\�o�$�.9��_��QC]跟� �J�}ˇ�p�q��@�M��XQ��w�;z��4֭T��3�W�2��!/��G�N4�Ԅ��t�z0c��}yw!�7Z|ބV�K��?e�,��P��,t@W���Kq�]�����8e�+� �n'�P�����m��*�v�}�M��,I��w�A�*��.����1��m$cri���W���,�	M�?�2�;����\�K�?_4��WwF��-�4l��	�_IgU�,/@������Y>;�+@���t��3Z5���*�?b5��Xrc�
�5�3;0�&�v��c�̩�������q��L�����~ӯ��8�>W}���
��É� ׷�p����&d�u_)�3����S��(�ݾ����	�������<���Sr��m6�d����j�e�b�3J�����&#}b�؜�G�K9������1*0�|,?��չ�8�.v�9�#�WE失Xe����3�Nvb!�)OғH
���G�4�s����V��zUܲn;\Ԝ��0�'!�����[R[�O
D>�n�&3�W0i! ׆ص��]6)�T��[~EU���ٶ�i0���%�4'(C�1X�Ru���e��ޙcy�%�t�=
��\��)*�=9v3���@������d�N������|��	�	-��;�zm�W~K�;�ߵQtI�m7�fz��GޘN��H�j��N����c
2�r�p-Q�+�#(���i�ؠ'.�Щe΀��bB�[��ц�7��(�S�Cb�%<x��47�L����eq�F���rg�E�
4Ϡ�-��1�Y��m�t����D�*��h��C�P��	��'�)d��]��rէQ�dkW�(�x�J.���(A�лj�3�on��Wa2�(pw�1�͎�Î���O����ߓ����U�y�*��ő�
��C�<ci�+�&�~+�ʙ���U��v��8�v̵眞*~7�d���3��ÑO��r�w�Ec�_ߑ~u�����Lv֞8�y��KK������y-���{�-q���a2*'�i|N�m�O8���&�tt�ks�\���GK^�`�셨�c�(Y���#����p��^L��`�VI���6��~x��<O[Q�I��ZN�v�.@��/������"��0B�'@9}���h��\%�U#�a9v�S��:��d�_���а<{����j���ُ'��<����=���eZ�^�á E��r�T�� M�V/8��	7g���.����y`�Y�$J��ixzO���f*�G��k􏠃�[e�K�)4����p�f���J��A�����#�A���v�4�z�!`t���j��
�_�1���!]ZU��R:���|�`X����Ӕ	�{�i5aqM�7���v�ȅ˪s��a�/���@���j������i���3�]�emQނN-zK}�
`u���q��5<;Ž����#t��n$GG��e/-���,���.���z??�1��Tv&�n������*�!"D�)5k}��&=��r.Z�<{_�?� b�AJA�����8�t���6���Ӟ�?�u�U�^�^i�ȶ���ѭqg�@`�{���i�y��5��1z�������V�i}}p0��0�o{|�C����z4����E�7�MO]yd�%�����ݰ�|���@.Ö�)c��<;��Ƞٌ�nX�
v�Bt���δ�ҋ���,Q��^7���8%��ܷ�{��T�B3��푞����
�����9牔���T�/��$�)�b�⏜���-��8ԏ�����K�g�8�_��a�F����������|��k�y@��+��n�<�hn�Q�_�7�Ҋ���4�sY����s"�0� Šs�2;�_����MI������t��L;cll���|C-�7i|����Z����p��"�,��?��s����J̕�޶:\4�X��>���A߁��p��$��	'v�
ap��Z��ľ���K��O����.��qJ[����vc�?���0`e/C�[���䲠�qR�;�~M(%�0�R�w4)�$#z�l���r-��O�XW�x��*���ɛ}�P�2�LhQ%�37�I+��`��2zĳeCX��4����&�3���+;�"ӓ�濠L�c��H���B�&B�� ��e�0N��huT� �i���챐��VL�K�Y�q����H$�O���*]�\D�]>�{e��T,\89�E���艮ՑD����d+�&ja���4u97�>�7��Y�j�ɶ8<�Y�K�O�+|�m�S���g��!�����2棤��>_-�m�I�UBL�FT�{�re����0]�/0�I�_!fzA��e^�Cz������l���ҫ(Ug:-%i�&N(��	���q�(X�?��<���E�O�e#�6�H�OQ���QB����3�� `
~��p��.Yg��CXH�9[�^G3<����d͓k���<����4��̖�сN�F]%j����tbXX�]񥝰P�a=�{�� h��J5���V]fZ��\�
SW�:��[+��2'sP�PZ��2��� �(qit�N;�; �Y�q�ԁ{ �;�xs�yv�'y�,�ze����DP��q<-���1�fe��v	�I'P��C=`��4Hh[D2hAA�(A2��Ǒf^P2:"��S�mi.\Ki�����ZH�
-鹪��G1Wa�"їM	�+����vh�d}����b��+��
SR!�����!�:9�xG�3�(QЌ�%?G4���x|b����h=kJUR��Q�K����
�
�@����y���������N��;ј�̌*a,w��Vŵ�!�[yp��c�n�Y�z�JQj |F�v��ӣRZ�=m��:�p�E����:�a����v�K�u��,aML9�����/!�kFu���X�$&Gs������l#D�:�]l�.��뺅�wnc;� 	x��:�O�����,��V�\�w���K?m�%D-�Q�
{�<`�t��g�����b�O�tq5�l���_!:�1T��:S���M�6��S-�3$�Z��]��Z����m�p��M���&-t*��Ǟ�x� �'\��ܯ��v(�Mp���l�\g��͋7�@�
~���|�
��F�+��5^��0o
m�C�pM筊��	�bB-(�X>���p���Ԣ���P�b����8͓	�[�~�Æ�����!��P�u9I)3�
���q�V;�O��~#�.��^@AᐣO�@J���2�G�.��d`U�t���Ǿ`�"jEO�Hp��h�K.Gj�G�R�R㭯���3����8&KlXݲ�U��1h' ���)��*�
eW'���c�[]�U�n���\JuŹ��E��n�i�ca��~0�	.�?�����5,&9��*�?�ے�bo�e&ɨ_��/�%L�C}.�/�� q��}��ˆ ���14�J�T�'�ؼ0y���?l9��~�:9�c���7�Me)Kخd���>�Ӷx؅�D�P�21�o�9�r:���?��^=&��7A�-�ǛR�
���mQÃ.g��§��_����).���HS�8֮�=��|`�,?%����ҳ�/��/��@�>���ѮI�ȥi��WCІ=����L O�ǆ�_�_<�у�n��c`C���(ڃ�\<�,�8��X��_
cM�ug��={�6�3O�lSb��X����Ј��z��V�e~��`9��9N��'��љ�V0㟮w���vCr��N��ӏ x�,!:/��[~����s������N�� JF]E�C�i��]��3Ae{y��	8�w��½�I����seOB��c=��O��L�X�-�1�F�u;>	�
��Y��]x\��3W���>������"R5lm즅.��){$RM��X�H�}3:��xs�wԘoc��1���U�n�B�;i>�
��O+�Zx��O$�P[�x���h�<������gF�^�jN�u��t���'�G�AF���D���a��nɻ@+2w&��~�/�����8򏙟�K��A���ѿ�1��ck�9X?���s��_�U�:����v��9�#�UQC'���F�_2im��R�Z&ߚ��73�X}Ke!��&P�B�����X,���Ř�`�8���*���|Nv���Ǽ��b�<�zҗz��!������c�X��5�wH�a�����r����K?�����Y�i��BЍ^+�^e�o��섴 Jb5�Ø��Ь�jWSz���b��^��^��a�z����Ǫ��7��L���*#��9�k��\�g[p'ޮ¾e�0���I]C��Jw�`2�ŃKvx�E{��q��Z��P	Pg��Ah���~&���:Њ�z|�Q^5��Ď�1����1��>f��3�
hץ:�z@����� }L��h���cXv��t�hV���١����+0�.��T�X�c-�w��&))���d���#����gs��\q�,ow*�u�Z-���KL��r2eh";<��\�D7쨫)TYwJ�۹2��6�����Pz��d���)=&��|0��ƽO� ��*t5�/��{�i��I3��_�Gbb�h�R�Q_�ʞ�B����mo�_z#0SꎴS��k��sa�4k�{B+���kY��
�U��BCFJV�2@1�yhO�7�N���vd5�:YG1@�t&�jd'cccs�E�����OQPmpvf{�r���K� {i$�8/nE{���}F���F*���7�([�HY��R����Zg�"��	�s��4=H#�%Λ2�}�p�rE|1@���.E7��Y2SW�[��o��Si᭨��'�X@O�-g'���-��w�'�S6|u��%�͜�������(�[ )9>!~�vj 7�<ʴ����<j�OM���2����p���ߌ�_1 �kb�tQmy$�В��\�RS�;T�]M�^���+^)�M�H%r��F�����$�����j]��A��mYn��1?QB��YoDe�7�Z�ᾗ��+:���y^*�*<��]W�2bLߚ#��l�7/r�L����
��.�>Y}��AC������/�(�|�H��ʀI�p�93Ѭ��S�o ��H��"fz��)�0.,(C�=\Op{O�O�A�����nbH��q�.K~�;�U�5	�e����Go�~�����ا %%��7Q��)]����0P�loQ�H9��|�Ͳ���*�N�@ Q���8$u`I��j���~����s�6���N���>f)�	��#gu�fD�1a��d���"]>{����j�:+�����\lb<�tm��T��{݉�}@�s��D�y����0{���P�|j��f)5+��W̙���j�=@!��^��@�S���'�B�\N�\=�5�#�(�w'a��q�SD3��(V��<Q��Ղs1}j��v�d3�m��;_JJ��&�Ĝ��l�L^�i����q6�� Ʈ�S���3�Jvh��zI;�q�#�8,�'΂���(OH��ۅ��rR|���!rvѿ��� ��},��Biuv�c��k���v��{	<i��Y2Ca�[Ϙ��D��`�t�}����Qt]�(�]BW7L���s"ÿ�ԋE[z@q�	�d1� ��bO�&�e���=;v[]H�Y���?��nM�0�Ն��B������J"M�p4v����ǅy�Yܷ��!�_�i]��Q�D�t]�����W��������u���`b6�s�S_@MBi텽m-��G�9]�PMiO�y�
W��H�]��>���D��u=S��]��R�Qꓞ<��~L�4ݯ� ��X���yGξe܃�TT�'��j`��I��l��Q���&%}t���)ezP�t=HH��4��h,�K#�%�!���z����d�� q��U쪆�2&tv�a,�(�����|�e1��7�������;�yJ���x��䰞�7��S�X��>pwz.�?r^BQ�襗���*�E�(�sP#mar���(F�y�K"�Q���e�T9��3l$�9���cY�C1���BW2B�>�q�K( \��=�͈)�=3!�Hs��g�J�&KW� [C��f%ݏ7��cCl
�/G��!!�BswE{@\Oe��R��}W��n>�|I���?@�s�:�f\���	J��iYw3 �6�\<K�������H�
��y�(��\Z1vL�:��Z��&��:*�XJ|6�%��B��o�0F?����S���<"q��2r
��a�4� �\@�f�E��]���:�)U
d��_�VY��s��:4�?Gn���8�h�(�I�g+6x�I�R�Q	P�7��I-�?q�8B�R��pm+D"�o�u�֛���H@iB������e)	�S��%��O*My6]����?[���I���$HF���#\�t�~��M�o;
�=�k�����*DtQ!��~#�����ugӤ�(ۍL�V����*�JI/L���5�^����
;�-gx,���h��8�2���f\7�:��e��M>�7Z�m֏5��o�|6�)ץ�ndm���k�_���+���=�#�}<a�X��_0S��r�f���B?� �����-I�aϗǔ��\�R�
	��1��l�r�|6aL[fly�����``���i�O�44:��bg�ly��Í��#�e��T�5�������\��g��P"$I�v���R�Z���5��o�!}�B� (%�W8�(������+���g(��h{�o���UW��~k���>��~�|�X|���%f9��=a���C�J�b-F+L��Ο����l{[f��2��P:SC�`�Ձ�/�����m墲|*>@qPHN����M��E�U-4����A�"���-w�K���11�e7�i�H��9�dD�@_�������&B8zO}lA:QD�T�/5�LK�J1(���<�?�1�_�^��)���R�����~#؄Y�p��=���%O�:�Q2D�p-n��X����!�Y'Ka�F�e�jխK3Cy&ڊ����� ��aNKև��'7=�S٧���j0����F�K�2}��"ˋ8��Λs`���g���A��'i��w��������Wr1H�Ec+%��q��Om�;=�ejh�����ʙ��2��g��I������ݲ���Џ��'�7�p�h*�ɼ=bXKR*��ت@>�.z0W>��"�>BP�R@�_8]��t�n��|8NRܨ��mi�ui��B�:�A���@��g���gJ����u��A�۠�),�(�:����\E�n�v�G^v�.�W@h�f���Jf�)�( �Y��[*�����Y��ƚe���6�E��?�gs	��	]��G8�(�7w�����{�(?�O-�I�~s��.X9�XpD!��&�!,�fN?fvǪ"d��@z�̌f�
p(�FB�ɧ�o��X5V���w�uѕ���.�12r^%�N+���	]#0J�X��08�[��+rRe��$��%j�����iw9en�p�͆��H�%�z�8prh��IG�e�4d*��-�C���#x��Se@�@mf=���EM�M?4���6sAd�1��H�6�ӫ������ش�
�m���X��Ҋ�۲9�FĎ|�]>*�g�Cɕұ`ݍ�o��8��6�����u��IE�)�\s��݁P�����-�oH�d+�ʼ��e|���N6�Ѡ�Z�IRCm�g����s���|�����0�
#B�2�O>�C��#�c,YbL��ˮ��`��I�$�2B���}lxS���LSG��� @���$�R��!���,�qB�
�H�� ܠ�����%L���c��:D@�I��ԟ�R��A���pYd���C���ײ��?D�VF��+wp�1щ?W 0���F����-�1�@��⌧
#����y���N�GO����unpt�cȍ��9���X��O)�ts��ȱ^4���D,�C�s�*/֖W�3���9��=y�	��;�]A�$3���\�t) t��6z'򎷮�CIes<dY��D�q�J�k��ȳH�ݟL�����i�6���1����r�b��������7VMvi|���g�~�C%�bKN /�w�J�"�[��~��8~��X�J��8KΌy�g-b�^5�{���>��O!G�Hϭ1�-9l�C&Jۗp�}��GJ�D��&��Ԋۊ �d���������!�ܾ���]�4�U���p�G���è��=����D!�bЎ��X��
��w��i0h��K�����N'�{*)���_q!�	�� v2ɗ�?�	(�c0f�F�NPK����e�o�i��L�k����;c�Zl��n�<�.B�䶘�S�P])hi���j����R�Q�Q*䔺g
3�79�je0��K�yeiSک��Ŀ�1|��	�yRU��*qk[����x�M�Sc��vw�����2XR���U�z9��]�حW 't��p�A{�̔���}W��!3L��&̓�:���#�:M��]Mqpm��3D��ڥ���B�!3Y��wO�������c�Uy��1��
2��fCT�Hƭ�l�Y�:K y~[^�Ji�Ttk��`ɮTR%F�(��S�3}>E�7�>���=���0��������9B)F`{���=He:��GZ]a@	����]��bT!���S��$l 5s[{8rǨ��퇘N�<�Ɗ �Tb��P�VY��q�v��!���^��/�R��c��Q��] +����މ1~����	vE�8��c��r�-�J�}����������½���c�Մu������/B�r�r��`(��C�����L�e� 1��-�h�$=�Z�!����meia`�K���h�ϚE�z
���s��E�T��l#��?������l<�8�m<')�Ԗ�Vs���*k�w1Đ�p�Y�^�4D?0f&h���vfì`�H�6��<|�<������@BK��#�v�^���W���\�a��W˔�yK0�74_O������"q^^�6~9����#�A���C��������:�����ZF�`Ṟ��G����O�M��t��}_������Єq��������L�旲|-=1���HK۔@)ӶL���(]2l�+-��1E���Y���8���D���R6/=�{��M�	d�����*�>��y����S`�<�����ŋ��T�F�\Q�x#�q��/�f��)h�d�B�6�BJJ�o7KT䑟�u�-���mcϪr��ް���ݶ��c��|YI��5Q���P�QȍA"9��N�C(�E���M$�����]�3��`|w����}+o��y�#W�oԭx���!ѭ���N;	��y�E��Ğ�~'Ԭ�9 D���0�?������X.`�O�꽏�H�"�f��( <ԹXj���I���� �)lYU�8%/�ޛqJ�t���0�t3���3�Oa^��裍'D���o1˜< ���]��N�SE��=�Ls)�&-�a
����u I�Oj�b��A��,���VN4��do�g�9J���1���LiohV���G?�W�<rj�6{��@���{r���*����V��Ύ�d�����^<S��(�U;�I�"�2�5��Ł�k`�~Z�8��0��[mk�� W�y�
Sv������/���q�s
bRP���c��P˞IH�X`�ۡ�
�=l�ʴr
}�EL]h���yޛk�Gz��;O�U!}��ppcB�lsP�bH8.IZ��p#�kԹ(��7]�5�]',��&���tr>�m��6\����Z?�E^�_�M|&���%��2����Mzʵ�ē�M�Jj�ٽ|��t��I�K�;`ټ���|{U1N�SՏ�(2`=o#�0�JF���|W�=L����Y�6n�`�H��x[�H�ƽQxHy�{	�W�,�Y'�[����;F�.�RJe~��<ó>k��O�%�����:�.y*���T\��s�[�X�
�su�s5N�b���/�T��y_�� �I�`c��c&�L?]0��}j)��c�d�mVH��~6�H��] ���"-zݔ^n6�;���Ԅ��
=�
{���n���
�o��T3�5s3�~�bO���B���B��:t3zQ&�N@�hj\����	�A�._x���\�%�ֲrD����I��8u�u�5 )��"�
4y��A$���|v!��9�C�� ;�m����\�@h�(�����h>�2��R�A$���P�{o�X�ժ��!�~���U�34��?����$�7S�Q�f�C6B����?��F/�+$>�S�BG!I'����zHe���(�M�o<<N��d�=.���u��ܷ�S"�u�6-"sl
�RԃRo1��^?��p\��+>�����͈|n�&���]|�Oz�>���*&^�ue%o�	W��0�W�d$ uQ��vÙ���T���Ŵj�jY�%�O*�Cwd��Jz��q�l~�[�H9�#(��hz8�P{}K)�_p��(�
�X�M<D������}�#�����00��a_���@1�:�9Fe�o?��|��n��<˂��)�����t��~HB(ˇ�w�B�~���K���;���Ri޽�G�v�Y��%���J�`2y��ܢK�nN������wT��.>�a3�Q<2lM��,]��� ���L�kL�� ,T������9��UYZN\:�"edK�mS����;DI{:܋�*� d�뇪ǋj�kPWi�$���UW��'�h=c�h��V�y��T�Jx��� _��+�ǒ>��8GC$X���EO�0�P*h�����~v�P�[;;��o~&+B�M���fO^�y�n�O4~�d8��pP���K�LA�d>��y��K�f˨�(�h/a�x�Ás��P��A����N<�N>%�>1�.xyDI��(�͋7;��Tp��S�]z锨��&��	~FWşϲ1$�����;�Ĕ�d���J�%?p�p���>U)�

ɨ���p���z�ۈd�k�fQWܩy�uͳ(��Vd�z�/cǜnx��Lč���� ���n׳zM<?�Pf ���{��z��9O���i�Ѥ�V�듣<�$�
]QZT���k\a��a�f�G�Ot��R]����ݹX#�=�����h�\�Xֆ�"È�'�B��?�0w�����i�̡u�%��]$g�0qR^�[��=6�Fyo�L33�榆T�e�A��IJ�3�6�X��S֑��GV�J�0�rpe���8�@�e�>���Kۻ�!7�J�\�<��IHq�Gɇ��"a�������b�������Z*�)xI���!ѕ	����9�R5�e���'"\��`�6��g�%��-��{+sjR�w�ܭ?��&F��h�� �k	3�_'p�ss�3���v�pTA�r^�	���kJ�����B-'YX��[���u��$�'���ף�N��J�U"˥�$�^��F����dF�'�"i�iKh4��Ps�쵢�g��
������Z)5��ݬ�����<�Y��!�Q���ynQ�kB�6NF��8����G�/���?�y"P��kimn�����R)�6����8�:��:!�S~/A��I�0�$��v�|Wng]y��N,ݬ�e��	��q�p��(5i�3>y�<�r�����k/�^�Rhon�W%oD�sܦ$ӯMc��ɯ�8P�] [r�!0����G��Y�OBC��8�#���{ᕃku;Q�ߑD�:߯�'?>YQ�O�nH�c�A�&�;d*�4![=��6O��b��[~�Xc�PVan&��F���j�x�~��'���5�*�[8^�(`�9�
�;�-��^Ϝ��+����< v"4+c��q������1,%�冕*0�"���t��r��|BߎՇ1��
�o$�Џ���Zm:5]<vڌ�HiL�p4���&E�R��ll��JR=t�j�ugd��ѕpJ��� �t ��q\q���ߕ&���u���%�M �Fn{ �E�Zp����yqҕ�J����5�w���iԀ� {���Λ
%
&q��%��LY�.I- ��Y��{}eIk�ϭ/\FF&"��,�a6ೱ�lf1&/6����bX�旎���f"���c�:g�Y���^�(�Kg��\}�{���� �����{P�x!��yl[yJ�~)�a��d��lZf���O�S�i~f�n����uc������YP��հ���n���Au+S^�I�9ڜ�T��,�S�˧A�ѩz�g��]���z"K��\�D��ҼS�˞1K��i��a��au��m7F|3m� %�)�O5�zxYH`�/q����p*0_�M�B�^�����@�ψy?���`HT��j�9:��� å���v$*�;_���e-c���x�Z6��J��������^Xҩ�E�f�e�䯛�������2Ig��n��Yѳq:.{*���I?=��|h��=��dţ{J�S��&M*t�r��W9��b����I�#tf�k��T\�" ���zi���y<έ����p�m�b�}����W�I�,�rOl��A��1Rwi&S�V����=_��~���Evօג7/#̗��-����:vۊ��ZZ'�Xb�ˏ�!^~j��
�d��^��C��Wca��qOσW����z��~};0h	݉�ۈ�; �|^�vQ
��g���(T�؏D�3���%F]�A�p�Z�mf*'Û������--���R_�.;g�6�x"�h����ͪd���K��S���bD�D��A��.�K^A�+?���wA�^ݟ�^�{u	�[)~�y����W�#!�����0-5�<N@����&��u����f���^��U>]����oy�P��$83Z��S��oY��.�$S�\��g!:�����R4%�5(�-N�1�ѭ��$���H���&�<?��,=L^,�&�o���|��}���On&J^��- 4@�L�n��	����!�S�t6ſ��~�T����kUc�� �M�@�ry���c�_�s)ݽ������u�X�� ����
/�~v�Mf���wV ����0�S\VV�<K�*\�z�� �cj��>h*�� �R��t�+Ŏ���t���]��)%n��g��"Xa�^�ŗ9�\5��F���,�@ю�p�!�.��w�I�̉r����� r�V�%���x����Z[?�muժ���&1��{k�!2�/I���o<k�l:3�\D
<.����4l�+�������)�H��R�J�8��N�(��^!ұ�mf�;�,O%ъ8�S�c���� ����Ĺ�AIc�q:_�x?� �86N	����}��t��}4�;:~ԇ����(4>�1�-o]6�XaQe�s��"v�����h������)��wQdT�&�a����<Wغ��[�_���6��f�M6E�x��<���N��w�Jp��I�7�F��M֢�&��OHK���c$B�eP�u!)���d>�Xb.��&���zL�+��3���Q�9fF��4�X.L��xU��E#y�nd/���,�R�O�I�p��u�����ff$b��W5�( �H�|UB���b�����/M,�YtYϺ&k
){�d!�G#Hoj�H�1��NR-�8���*�����߄���XQ)p�ķ��i��������gDX�vDG^�̊;�7v�h�0qнS{�]4 �ɂ�vt�D�]��	������	A�p�� �v�o������I�bO
��,y]±������F��[KԂ_�2���vA�|�Iξ��7� GR����[�KG�5�Ф��D�����/�%k�Thq�6,�)��5KyhM�w\�I�db���}�E]vLMSj��<��.v dr&f��3{�VL�Fe�'v�����т����Y���o/����f1S��oy��ٳ��\����&:\?�n�֒�����@!	k>1>m3#_��'s{8ަoˇ�14��	��� 9�������W��+S�X���(�P<AZ�4�D��1t�˓����F����o+��b#\rC����.��N��0{E���ʃ D	�"6��:���D����Mo3��É:��� ��ܟ�W{�"�c����I�����ګ�ܡ);�t�{1�!���7���
�� ��b mw���|t�/ơ� ��?[+��A;(ŐH�KK��)�M;l��wb���]RY_a<����{�9�3S��ޮ�J�^�|vHS(>�F���t9�w��=H���ﳅ��t�GWB��B�S����������u[8mER����)1s��#�D�Ћ���s�F&��Θm����x'��sWu�r��Z�?�>��;��b�m��D}Ͻ��t�6� ^hő@n������!$��LA^v�t3.��VF�
�)Ը��!-�EB�	��Ÿhv��YTi�yxss%��:<�^�@W���ޛ�� h����ր�Tl�� ����MȂ$;EcS�cڂqd�ш��2���9e�����.5��-/A�A��C�H�/����.��b`��W��Ȑ�`LF㘩ȋ6��@=�mz�i*�Y���Uc��Ѵ������1ywo�`�_b��j����=�U�5�*v3iv��!'�'؎�lBI9O��!�*}��H:�
�#�.	s!���M��(V,üH� ە��㘭�/��V���u�T��X��+g����7e�����}�D����528Բ� �k�鑞�	��F�f��>ΟIŎ�D��i01�I�N:j"���lyq3r�����Ţuuk�/U9;��g��=�|V�x_ʩ���).��3�]W�4�9�&
S4��2}-��B朓�Y[��[��k��<�r�]-�N�ju�ph��?�H�<�Eg-�ʓ�\�s��֫��:�iG�(?U�ũ�Ja;��*&�u	LN?x?��)*��~��~����!Y���Z���Ó���h+��c(mt��UpNr��a��6���Ғ�F��Jp!�"S�d���{���`��?�	��Ж��$$��{�� �+�Ҧ��@YD��S�0�R �)�z)���^	wD�dNzծK�ƀOO���	ftxR+j�9]q�"���$g��\�.Z&Vt����E��O�����p�^��T߅�R��-�����wJbW�+ ��Б,�aG�MV�R��{������Im@�����C���{Qӟno���E)b<�s��AMz#{V:4)�^0�^!�-݇�~ι������_�V��[yL~�re����ǌZ`1U
�gu|H���Ɠ��������:�m�l�u�Y�1���h��M�r�	}m@jݎ$!]��ɤc��@��"���� :��Q���a�,d�kHi9^�n�-��$#�>o#�=3]1B�ͤ�z5�6�)�"/7�d��@��W�i�eZT��K�s��C��É���	��~0�a_��)W���z=�RԎ\l9r]�䡝��ۅ��o��K��&� �E��mL�`��Q�D[G�N���yh�$�߄3�6�*������k���{�w��mm��y�2̈��e^g7~ư�X������c�P�T|��dq��}��Zc����9*����睞�c��4���̽)�+��Ȅ͏T�י�[.K�0���H��ӻ��v�Iv�Z/�w����|x��*,���q�m.TTD.+�n�� �^������zo�h1�0��~T�Ď���%H��R�9L�j5�	��qPj�z?,��O�h{κ�}��r;���lu�]�I����H�w�}:z�G�����$_����_���p����φ��إ�W��״R6���=�MZ���f�	�B	���c�N�@ya������2b	h|��kU5�	2��7�S_}q��61��@V�n��S�]��o��I˰Ss��2<��B����Ȓ/�&�-���B/�pG����LY^g#=���kq���Փ�={`c2�����3� �Jƛ�����m�K����e��"�1daкV+E��ŧ7f��)?>F�����C�;�%�\Z,���:Q���5K?&�-�K�\���Y�:I��=:��H	���(�y�]j���G�P��=�l4޸���#�9գ�����4h�`���M\��$��GE N��>��R���Ʒ��=f�T^��,��\�3�$U@16�Ш�E�@����<�K��u�S]L�e;�@��#IN�<ds\�?�G���┒��q�	��3�X*J�DmmYC�a�� t���0�!K܂��H��D�|����n,u9�
���Edl���-�+�Ո[,'G�Pѱ�N�(u>~g64�]���}�KC� n{��Z�)�e�t�����"�s(��楼;]Q�g�7*�ˉ��k�(�YbU��uP�j}w{��R�� pc�c:�0.EZnq5����\�#�J`���X�:�L���<G���e�9p%^q!�o[��7V��p��'.�[-.�8� �TrN��Z.s���cuz׭�e!��lc�B��BW��b$�%a��1�DPNjh��ԫ*佸_��9A,��]*ZUQ��W���re2�c�Ʌ��3����Lʝx3E,�پ�p6�����Cf1�7d
��#�z���Wn�)�:ݻ�ԕK�&����]Q,�:�0A�7���td�݅/�I׷h���/���I������M!&N�Ufa�[ ��g���� �G�����7��ۈ��pdUW��M�T_��JXNVB�_ ���ui$2����SM<p�Ԫ"
4��ec�}�]��չ��p�E\��C$i���.����)�"n�đ��X`�\�.)1�,w��������#n����JW`�����_:�Z�F�'��,S� #2F���U��{�հ�
0�M[������:��Fa�&�O7*|�o*�,w�2����{��I��7�Q��ĉ����j��WZ�����J���#�5��ϱ �_�?�o��Np�o�o�c>F��mX�y��m��hqA��kG����������e�o�ߨ5ֵ��ȍ{�$I����jĶ�d�J�L9�&g��Fd�Ǵ3f�3q/��d�~�ji����dtH�=eJ�}d6b��ÁY~]g�GH8��$�Z+�g�h���r�P��B��"�㈴�=���b�+���1�)	1��.�#:���i��J̚ ����pƔ��3�XҞQ	Ϙ|7��2.P��OT��6������r:���q�>�(�s� G�iޑ]*�J�����Eo�y�w>h�4�T����i�F��3�E���}^�U�"��8�����b�M�����^2��b+�Is]9��/9H7�GaJ�c���T:��*a!�Թ���]G`'�/
髢>��G����w�^L��ew<}�Ӭ��Dx���T�!����Ɵ<e�Vi�5�sh���\ВFI� ��U�����Nf���9���qeC��&NV��_Xo�����b�ⱺ��DT1�2�@f�}��EID�V  ��m����Wd"�����x����Z�jV�����.QX��s+�w��Ca^�\��U��@3�dEfm̚�%�%�?D}0_d�a4Tv��~�4�K~#��5�;=��j[$��Μ��;�"Tk��PD�<�͋{4+���$�c�K��ąL
wH�k
N�2ܳ�؅���J�9���
�*dE+���&D~/Q��z�$}ާYn���
*�j���:�V�z�2#�f�yK%m�PA�P?��u+T5n�_�������K��<���z2�;�h�~D5�#a���|�h�!��^�#z�ʂ{ߡ��:���૴w�#������cЉ�+�☱K�D��U��(NEn�99=���NKxD��O��qsII�b��[E�˱�R�z��h��`BodF��8=sJ�,��r�Q�ؽ�De�\d�*׏��m���X��(F7��3�G6�m���������a$t͞�h��8hc�g1�dR�o��ϔ�'g<6�zy�S/I��ME�����4K� �VW�Ӝ���5�������q���E�pG1 \G�	^�N��<��4�����������/�p	�t��Gq�]��@{�O��8:�}�@�Ѩm��+)��#[uu�l������S2q��B� ���2�G�/�U"ϕF��Jٗ܈�^%~��Zs���1`#�S�6tY�)�����]������M�����.�gcWA��b��`PU>H*h^�R�uMv�L�0�`�݇��@�����=E��)6N�s�l�s���n�'_�_%u����h��yr���c�\��ܕ�HQ �}o-Eޣ�C|l���ض��|�(Ef���E��i@� � �ܑ_��􁴊p`<����da����:�1uh�Ȯt�K01,=��C�'��k��Q���|����@w_N���sɐ(�r`s��RɃ��x��N��fi���
��"�N�Ifz�bT�(��f��K�:���`�ߥX�B�^%<�J�����a��+cQ�j~��2Y[��z�Aei��Ј�:��B��%�H�vK��buEJHG��8r���6&?�2G�z����g#M�L�K�t�PX�D\��G��;KL��*���L�	f�=�&�n�>
Z��;�_vǣ�{�ₜn�J���W�S����CI�>�c���h�f&�!zR�ο	ӳd��]�1��,GMn��D��ѧ���KiWf"���M8��ݧ�_8xx��D�]D��SX�0��Y�=��o�C�~�꺫���Q��$��	�F�x	_a�M�9��� N�#���d7�`��Å�L��g]Ά�(��(��:�o#�����8>�Cȅs�G�t۰������qG��?O�(d����߄������js�-@�t~�3���H�5{�cXm���F���.C�	X�\&�DF�0���}�{~��C�/j`��<J�!#+{O~��KA �;���(������R\��ƍ����ɰ�P��%0|�g7 �u�o�d�7��!܃�]i�i$ﾧ�[ɸ�R/Y;�~���>7� yU#�͍��(�'҆ۢ���Y0��:8�dՠ�t
�#}��+瘐?���<����%�W� �6:8q<כùB���Q,�L�I
B���#fY���ek��d�������G��#�)�-6sfz}{jIzr�|�[��M|ܰ��=�S�I [��M*;���<��	s8\����Ț���*ҳ��檔x�8W��65�b�..��}9��b�!J�㱜��$�?K�����Л���Fڝ��'|�;n�I���iO�C-c�d��.�v�ϥ�����������q��مw!d�K�$���mS�C���UL�ĳ:�)�Ⱦ�u�U%�|�Â����6d4�[l:;쫽��8���S�)����Kʨ�����������X�~і8)�s���ͥpY�=��������@#���Qk����ޱ��]>8.pe��+���8n��������*��k��
�Z��Y�7�7�C)�B�J�O�Ͳ�����a����c-]��$ j��0z�g����c����;�T��+ "(���`�W�x���WP�H�1��9����-O�8I(�eʙӨŖ�-�h�QM�ָ�0mz_�'�S����7�x��v�j��Yۼ���ǲ��X9����Bh/�����:z�uRu�n(��Θ.-Y+0I��:R�f����s��(�꾂��k�B�bOfs?�8���L)��"v~��˿����y0���&>��F,������"MK�aJ��=���v쳫��N�[
���C�ɟ���:=����řjYz�������ʽ(h�11R�S����{$Pn�����;�k�4�������*�D�-��2v�t�=�H�R��sl���nu���aW�}���}q��BW�v��@w���,D��D&�tp#�bBMH�=`q���'1��k�w�%~�_4R�N5+M����7�������3'�я���\�	B�v�u�#A��L<U����'W�#3z���7��_��%��2�ɛ���Y�;3�"B✵-�&Q :	)�\��1����j�z�w��_�6�<�92��0,0�� 	��\�8���l��o��*�ԤiS�3ԻP=z'Դ�b��GS���l�mV,����TS�ܶю�k>6$�&�+Y��;j�E��Ny��d�蒙LL6?��m��8"��w�Yv�q[o�%y��� W��{K"������I����D�?3�7zʅ�/۶��9k�����Yt��m�S������B�G� 3Q� ���{x��l6?Q��gΚm!�r�k��,Ց���X��\���ssP%O�A�Q�)*o��ǵ�FD3�S7t	����9�Y�R$]�s���~�ԁH��Js�� N��s�\fH�E�d7ΚI?y:�;߷"ð������Ƈ�������Qd�čQ�S�p|\�YTma�`����ZMZ�E禗O�z��Y�;*� J����sK�W�ۜlnG ��W�d�B�.�H�<'���k}���%-{�Z+���ޕ���PЏ��gC�s��?�f�u��wz��i����p^3ϔJ��	�x�>�.�6���ełq�c�ۭޟ*xpF����䨊FcZ/��d���m~l���lq@L�Y�,V?��H���ѳ��ֵ�L��+o�=�C~ �����Ӳ�7�$�6�rMg�098 �:V+�������Yu��m����qWk1Ư)}�P#�@�ƪAod>LzZ�%d~��v���t��*�O��%�����M��,!�<?~���Ѳ�)G���x�*6��2�){��?��.�F����^�D��j��i����s��q��l�����q4DS��ski���}�D,8�����A ֠M����3j_2��.c^��i���^�+^�T}+�!�AU����(�#::���2L-��i���J4R [��
r4i1��F��f��Z��l��AH/{"��݂���o>�[gߔZG�H/R������=��tԒ Ѕ{����|mN���r�J�C�w��@���9��:6��nqy��"�14�����	�_�6ٵ!0$�:�����Z�=z�����;A�e�kyqh���n�w�{p����ܻ�cwu�+�^��^y�H�Q7�t�V�[G��;�-�g3~��-��A�-��Q����ǲ)�i�*��(����H�Zf�&��Ma�a_��K��/�J8itȠ	#'�޻���@|O��=Y/O�ta�&����QM�	���?��{c.�z�8]��"�al˂���;��u	�Bv$ئ���Ik��du�~�!����An�v���*E���f�?{Ѕ]O2�X8<i]���/�o��Bp~6��oa�(m`�m�!��y�Ҳ�+�y^�zlD5�x��Z��M�0t���mea��:N<�ߵ"x<>,��	�z���3�s��Jn�\���8"1�� V�KG�'T�[q"�=!�Ys^�!#w6}��}��0viK�ۤ�H�m�oJS�δ��G��֗�FO�x���A��nw��;�S��E��7�F��J}Yș���(�ΐ��f�͟�eNJ:sQ�|��yܵ��{NOa�L�YI,7�x�KAK��e���qT����¹0W����}>Ƞ+�t������5���q��cVm埠���Jge�19]����)p�=X�N%/:�&x�+Ñ��R8�T�:)����5u\�	�6�r���^���G�&w!�bZ��/���V�0�o�b��Z����5fj�O�άD�i3򈦟�`��%s�goZ��ߊ�7���:+���~����:����y����u����� �I���R�Dj�֓�3dC���M�\I�ta9;RW%T\.�Nl�ii������.2�����]��.Y�.p�s�l.�Pt1-���Wx[9b������'��	�0����Q���y�f;h,��X��։r��S�,���	�W�q|��wP�����*F7i��Ǔ�L4K���$Q���OZ�ץ����`Ő��Xy�D��P2���l;M�S1킿¾�U��n�4�3{^#@���6�5�U�R�@�Y�PߦWBy�?qk����ҕh �U��\�a�-�q�O#8�?�>$�P(���c:y������ʞ$����QV�C8T��v&�e3�j|�3B��A�2j'͏���V2�R��g�[a娍Q#���紻��_����R��J���!0tզ����o�`P՗��-`tO�S�ў�Q;� �<3)����9��,�V� 6���Ƨ�S���X�=d�)��<~�w>4T}���u�?`��mW��S��YF+&�@��\�M��(iR��Qm_�u��o4�)4W�XH	��@�~CX�Q�"k��e	=k���
7��N����z��)�u@^���x7գ�ry���D�}E�o���	`55���s��;��7�{�`�r0���K�P���XUh�ޗL\�n��`�a1���1$[
8��M��Q�O@���>H�t��mQ�dsBMH�kЇ���k;����y�\��iH/���)� ��$�-~mxX �'�S��x��Q�_Z��+.u[o��}�f��n6�}'=_7�E***x��D7G�w���5����d[2l��]�ˠ�f��i'wt�|��gߺ1�lQ	�u�W�V�����f*]W�?�?575�\R�����oš�v�8C�/��#�6�AlV�Iu�b�56�۪|C��ϳ[$�F�v�GT#ek"ϔ�R̸�"DԢA�K,��M-yL?�8�[vf&���Y-�so�hj��т�q�pcvʶ���c���"M����.��^�?�����b4���VKO�&e��2��!�f�J�z`	l�X7c�%��e��);���3��|+_��r�/}��b{4X��_�L:d��!7q\'�~�0^ ���������FU(X�T�E3��`���1ui�|���P����6rE��`�<�!���w�z�~�~6f%�W��t�Ҟe���xJp��E��e���ƪm����������Y){���v�)}7�����<؞	l_�%��Ώ!JZ#)j,�kX�i���j�w�ĉ� ��s�뜸E��.���d��^�yՠ�96U4�#�k���IK�=!)�hH��x}��φ˞ܓEV~�#h�j�c�V6�
���D�)�'��^�vg�$!z�UK� �j����gJ�^Ǩ�J��� ��`�t�h��8W� e�T�ǣyz�|���k�%&�g��g5�����8�+A6��8����ȽKE��~b������g�X��R_P��;�Z�U?^�rG1��6��p�#�C����~s%RT�x{�R��,��)zk�V�%�p��>�k��ur
D��ugѓS�.�$:�S. 5M��� ��L�m�����?�?Ȳ'�yl�!��o���-�)J���^/�3HT7x}�k-�x�Cl˙s���n�?��|��c*���C<���~Լ�O4.���r
$�u�zw
�G�R�籅����d,�������z{��!��u	�*a�����of�1�^�̣Վ����u���V���R�6��h�l�?��U�|��}�k���B���*�����l��2@�]8x6��G��|8���)�`zI�?��Jj��@�L_g.<��n����*����4\����v�Vc��;RL�9��8V=a��K�9z�Mm==��_���s�\�b�O5![?� �jz�C�N�a�wn��i�p���#��Iȷ���w"�f�V��^Ooᰕ)KzOpȹm~��k车[�ZW�Jf&e�������x�V�a5��ֵ�y�={Yj(��LQy�`��0����?V��I�S0�fR�^�)��2ɣeWIr�UL1G��!��bѯ�2�	4:H�y��D��Z�D�M2�O�~����T��ik���J��8
��*gj@���JNu�Փ� ���6�~:���l�� 5�;��wv��K������h�B?�f�+w=q��V��v����|}7��D6arv亷���85�%�9������ϧ%g�� ��%��:���Y�_�LjYX��kM���VD�R�����̐�J�j:�{�������`�����ȷ����P&�5�x�
��w��g�=���1`�@����7'�*C�W��GUAq�N��-�PM���(BY���2i�X@�:e!�T^A9�]���9-�=ٲ�Y���ЊK�]pY�ɹ��kE��� � [$�	�w�ї{w��!.�!�g���c�(�����6n좩�O}�6��`6i�� ��bKi5QjC�tr�$���eՍ�)���d���]����n��1N$^ǰ�^E*牢٠c�7�(ʄl�b�	X�Ġ#�Z{��ҽ�`���l���E�Au�E�hx �}MF2�v	Ax�ާ٧�7ə�L�}�[�~�Wf'��v�YW�Pt <�["�RCy��Q���;[�;̋�Ekg�m-�iCf:nu�5��3��l{Os)�=2 ���*ŗ�7;L[W�㛞02���|`���RZ[�e����� ����^�B©↼)�b�I�Ee��hf(�$�餛�'���	��23�|E��v�B��+d�/]�G��9��J�+ן�w�9�j�߯���A��j|�?����:{|8��
��!&V.����=ē3�c_�~��^���m�~�*��'�W��]��deS�pť�W󂵒e�pE�4U��A8�fݿ��f{x�✹�_���2�gv/��Qe���<�����[I��������v$�� W0�J+4�䭙Q2јd?�SU�����?2��k܉�H �=�#�R���E9ΩBM��ư�1��~c�8������jwƦ���7
�V�_���`�
�+d�RORM^t��*�(",?�!vO�->3��l��n/4'^��2�e��xb��.��B�5{ z��_�����'�A���P=C��wőm��Kn+}J�9���o"�K����k�&	_�[<+���
�n2�iy�V��M�8w{+��Y�]E�"�J,�e���<��(��׏O���������?F1U��5� *��DhP�ޏy��c��v���&�q!V��g��"�JXp��N��@$|�#����G\��beNWU���9���?�m�P�:z,���͔��c yw�L$ޚ9N��`�y��0����0"t>��}X�N!�R���ݳ�b�5:�B�Ӽ���g�Z�ky���i�FwY��J���9esŻ���/k���.�pMɚ�R�w�2��	)�V�C�v8�3
$b��'��@�_K^s��"�L��G\tu�v��؞sK]EJ�U�"�L�kDP�N[�������P�D��O��2p0�Q�7��mJD���jBD�z׼#[�2B���"�%^n-���#h��4�~��24�V�zF򞁸$�u����xh�K�VZF�GZGQYW��z�I����ԋ́��zR�<�"�kZ�����v����؉��6Q�h0���O�R,b���!����~<�c+���3$�l���]�D#���*}in�~��}3+O:#L�*$-��	8�f��#,�g�Ur�$@Z@bᡏu�aJ;�ڈ=��!��h�y�mb�h�5����=���ޑ�L�S"v#y���ڏխ����M�f�"�%#��hL�������'��R>0�B��D���i%�X���;�V<�\_%l�"�9����U;6#��ꕭW�[u�J�Mh]�[�Sm\��5�,��P�yE���%���8��N�G�`�0�C�I%.����x���Zai���J�&%g�	��нJ�LK�G��&ݙ�)g?� �R8�)݆f���V��i����U?��vP�T�R���=�1LJɩys�Ӭ����`�a��ʙ�]]�����So%�B��Y��`&l�Y�*���k�w��uN1��Qǅ��}�o}+k[�G饻$Mb����8l�~\]h{�D�5[Ы�5�5�Aa���ԛ�lǫ9�DP����W��l��v*��+oo�G����@^!SM�ю�Yߎ�S{�=�9�kny�9���N���E<�.o���*�B�|`�*"�8[a������Z���L�|�!��-_��δ@[�vւ߂st�i�FjR�$�Ξ7�p�!V����a~Sݜ����Gj8��F�E(1e��	��J����\f��6!D���H/�[˺B'�N]oMLhSM{�.��q�%M�p�Kvz���L^��^XQE2
s���w�g�<����#4t5A���媘yZ��c@�/޴,}��b�H�4D<�C��@��b�4�%n@��L�e��=���	��po�,��U�-e�?3��D��	㤶 ���5�n��9�:v��V��Er�	ֻ���P�!b��{���
`��]n���NY��۱J�P�mlp��c1P���Z¨*D?���Z�	!�6 _*�+��?��8r�� �cQ)�U������%��T�A�����l�n;�Op�V@ge&����vG�U\}\8O����R�Ό�0�:�7��ŧ2��	F��7��-Շ���V���%N��n�