��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��f�)C���s��#<^�"r_�ׁ��!�	)����-�j�v�1U�_\ïL�Y�Y?��2!>_W�<F�d�du�Ǵ��q����D6�k;_�;�.�n�^;ܺ*
5y�d��<��	]p�ԟ�X�(m>k��`V�ic-�WYj��CS�ì��{��l��A'�����8+����SK�ΜxR+`@];��a�O+
z
��ο�,Y՜�ᥖ�pbn�m7;��6��ǐ�8Z+��@y�\X�{��q�}���cc������[DG��c�N�݇1���fi�5+��ӹ��n|S2諸{��A�Xɟ9Ajj��k(���h�8%��S?d}�ܒ��Mk�j�֧c�����{�̚I_-�b�oC���h����nt�%%��%hx>��@ky=��$P�6���l4*(1�K����=Z�i,d�����H��m�N��c�����j5��LH����z|�y �Iᜂ<�� #)��1"��U7��Nk�	�(�\��XU�r���b��uԂ��e��hɊ�Z�(8^�./]�ڌ�o$D��)�,��u�^Xk���"5�5����QŦVd|e#���a���!��K�᳏pA ��PR�G-h�����Ngz0Tv)/e��>���o�O�F�|��(��J����q�lW�9�g �^tmum�_!̓��X)u�� 0� ��<S���TD�_g����l�+�bo�o��5U�G$���u�C��7�p�eT+�='P�$�UG��]����c!E`����t��x�.��/۽��5�6
`�H~�>��ɾ����4@�|�(Ǩ8	�@A�o.ڇh����h%������yU3I�)"%f2�A�.�����t15t
PX�	
+���Nj�oJ�&[���t柆/hD��T��WE�
{t������iRΔJ��D8���q���g��!G�
XC./�5���W!���X����(1!�A^eU�	���1'if���o�j��k�7C���ҁBD��=�M�A������:۠�!4�{�Z5�5��7}��Ok`'UT��RX�Mt
��G���@��\HL(��A�x��E�d��=1"X��0ٚp�v���65�k�9ѩ�2#9��v"|Ŭ
��n���7�����UU��k���򎝹�
���I�����t�L���� ���g���bND��{nLb��Vr#P3)��1M)�Y���.T���I��u��I��X]R|�qc��a����[4�,4�v�fB���g?"R���sm�%������������4�=�������_��M�W�YG��l�s��FkD *��(��b,g���b��l|�g��~�Oj�����S3���3�za�R�7����ODBsO�)��5i��7RΊ�
3�]?'b-�#�Fb��>��>Rg?�C'
%�Q`n���Q��b�V��o3X~u�HS���L��R���	�U��p��K��A��U�mapp�b����g����9��"��z9�I�$�!���PՔ���<x6��L}[a�͑0�+����!�F�j���]jJQ7w�+#'sqVЮ�k�|��X�5]ɋ���雩�WpM�Nϒ�	I烨L�J�q��j��N>��}��cC�~��^.��;M����}V�6*�yAI�5 ?�7S��9�������p�W+	m��	JPh՗�'�k#׳���6c�d6�J���*���I�b6�A���LA�0$��H��\0̽�q*��~a��G`}#�H\(� Aߘ�%'A��+ӡ�X]�6�f�I� �Ug��3���Z��*�݅?�����{D֠�?���r�[4�V&L�֬�#SnO��b�Q�E�(8%a�bᷢ�'1�|��r��]��WU51����3U|��<��8���/Y�J����Hv�N=L�Ч�'G]Ф�0�{hi��}fYʶ�_���vE��Ө7��M#���p]��̡�V��H/P���ǥ��\U=�GD�澕8����B�K��)l��ޫmz��cXz����D&�.�lA�&6��C��l�u��_���`l\k�'���_ LR��Q��P�;8��M��=H�6�2���9��`���RXi���dA�FK,5(�v��ŭ>�� �~�&���g�tL����"	�����v�ۈW�B��?mG�;�1�N�ܬ�&��ގ�G���LQ=�R���&��b��E�9hU���PB���Y�~�Q<����ʹ6��J�"{�;�l�f1��>/0�5�(��c9�Pl'A�j�u=��q]�r�c�[����Ƀ5���A��Cw�/a����@z%w��6Pv��-�~�9�W��̠s?$�\���>C�d�kImr�3M�]f��L]�'�w�6�����K�^�O��X荨�G,�6�龥�X���5�Ǉw�v�����!�W��I���c�f� Ky�����~	���VHni���`E��{rڷJ�Ғ�b�������s=ם����u?n#�'E�L����jfW٫l19��v��"p�7�"D�ьs}Cbu���. ��]?�������a������Ϡ�:����讀b]h6H�⣻��MG�¶���I;��3�=J�v<MC%����N#��a�*��
���8�D�:�24���D���3�'�/7��/�g".�͸�����&����M�ۧNۂ�s�k�g��W��#=��\�� &8��E�	=��T�����D~�]�y�\�~��V��=�_"�|��TV��drYؤ�<�O\{>�v�=7X\M��rf�'�B��&P�k뼾'?)>��X�t圾���&[�t��4׌���o]S;t��,�����浬�}�>,�����h�=FdʥcjJ��i�:�O���4
�
�*t[���L����������������KaØ|�S!�N;����r����W��ܷ:9j�$�b����fy��%��/c��>�L�ñ�.���aIJ��"5�c�w�;Z&�2�)�=q2T���o��N���J�K�a�2nh�O�/&�p�])5�	��_3剙:�h� �\���|����j]��%�եVލ�{f�^�9<F_O��>%j��_���*��/`=ZJ[�]�������ݮ�4�ȧH�0���`���+EA�;N�jV�`�S�����2�]�YW+��g*�֣�GuH��'.���a��y��T�oC\uaeP��m�;�86�8����3�6�v�^R!���駕N���[B�:� �ji�/b\Mg�l��q��'�(棽0����v�!���8�AUGu"/a�K��稊2����g&����6 ��	�ԹU��ӯ��U�jo^<����	Z�ZidJ�������OJ1`��2��WVdTqZ�S�GY�tN�9gB����MCɥ'�?j����>�ګ}���6�&2:zh�gVO��AXK���Ǚ7�.�D� �%��D߿Y��O�9��,��\��䊄�'���ζ),3�+��&�q�]6�[����7.	�̂�#�K�!07r��3���������2CtL$7��.
n��0Mɗ��I�#S���\Е��`�?c��$/μ#�*�%e��pq���b�1D��i�*���I>b_��������t`�Q����:8h@�k����n��(q�\oܷy��ϔ<�.�F]RrȜ�v��l�lU�zִ�#�{ l,���A�ty��bkPq�/D����Rҕ�0^`�
�Q���d��*>�qܨ80v�fq5P	���Jy7Vɒ��U��u�����#�4���oa!��,<�xI,@���u�o��/O��E�)~=u�I��􋏝4en��!�q��������p�OCW ���~ȩ2J�2��K ���bE�����TٯT�~Ϩ ���K�D30gD��;o����K���/ިQ�/�7L&���e��c�6�9?O<(���~s�F�Az�����C}�N��Nb.�s���9�H��T(?����Vͳ�=f1�5�����2.�tQ�^j�S	���5��L�u@��W�X:Ұ�C��c
��"��93o~��MhiF �y�w�����H~�+����D�݀a-.WzYʈ���ל�\
���7$w�[�۵o"�i�^����m�����F%;G?X���2#G.��˔��қ���Ȑt��KL;�Q�Ӽqw3Osף�l�?Z��$����.��%N���t-.3�n��"U�:쳱��h9���X��̒aKb��_���d]��$��ɛ�3S�)P�\�_4o��
ߧ��U�4��I�����[��^�+,� U|5N�19���Six9Һ�V��*�xGl�.M�)����Dxz���_m��\A��&�6R����¾W�!҅�:?�+�X<�W�qϧ׭Z]Zq�挣�X�c�nE~�o�M�_Ơ �t�x���ĉe}TQ�#U�;!��Ɯ���Y!Hdq��\�9ڭDva��+��2�p�?>��^�R��?q�R9U�aK{P �����9�`i@N�A�*�m�:E���.`O��sd�d0|���(��~%[k21):��+SQ�f�IՌ >:W�ZӃ���4�LX�V�-0{�(�ZHHZo�(�<�#�>V̘LP���#"�Vl�6����~�-�'/����N3;¿%�u�b�Pir�%Qk��\:��&����H� �����Y5����Q�%� ��T_�����v��-�'>��"�a���H`�'.��C�)R�Itװ(�=AD-f]�cݻv����]�mX�I%Q��sQ�$Eh"=:����ɒE�~n�?���Ep�L.��C�����D{�>����jk��<�f+�1�}���47c�Dn�����;�4��kl�ߚ��Ϫv�)��Y`�����-j4��\��f����}TJ5/��0�)��@�A'�7)q����i�&��M��V�C�����G������*B*����:�M��k]���(�I�c���N_��
��Zx,<��V�s��"����k����L���/�llO�3���M'3��[�'d� �"�AF��Vx^}��uC�Y#�|�	:�3F��m��ո�6j�B�p!����R����o9
:�ަ�h��zjoyO�������B���^�
��#iiy��oŐ�rR�'	���6:}j`����]��a)�!]{;/KP[�N}n�7J�xe@):"ƃMr�����6O��;޶����s�]�����E�h�����i����h�BnyKL�[��"��o����	�e�"κ�Pׇ�aK�f�G>�##�7�4 �hxq��u<�x�p���W�ܒ�×q��g)�!)�1���3�_�� k�D:Tu�T��m������9�s�]��_2@ik�?�X9�f^��P��<@+��w�����6<�	?dI�?}i���ڰ��"�ʪ��j^z_�6E��/l�&��ҦW�r�Ƴ=�q��ӎ���+��r#e&�	������`�`�+�P��ә�T]�����~f�>���}.t�m=36���wI�s�t.޶��׻��Ԕ
�ѩ�<�lo8U����%�C�`p"�9�%~�P����[� ٭�w&��WVx�/�v�ݺwU��r�T�4������)�;�r��\��FƉw��-rҷ�(���hН����i�����Ft_}���Z��MsV&Y!�FB�'.?�3Ȍ �E�8� ���L��m�;��Q����O$�-,�f�}����>e��r�%�^��LES*r1��>@�O���⛛e^��``��xI���_j���I��{��p!ײM^$q�G@0��,��)�c���xx�)�i3��π�w~f��]:XC������/t�`EX�R��;f�x�����SD��W2���4��Z��ӚpC�(VԳgSV���܃<#zk���6��Zr���.+�