��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��d	�%�� ���,q?=btoX�j|����P0ܭ�a�!zbbI�sݻ��Jd�i�_�ϗ]mʪ\�ڌc����؂s�V���t�:v��-,F�c�=�E�����@t�^�|�nc[���ܬ*����qTd�������LT�r��&���J�Iv��_n�ib�y)x|a����6��Q�#B���a�{�{�A}� Ax�y��B�-^�+ʡ�7b��TX����:�-[4p�?s����D��b���ŵ6��K�i����Q�u���|�¢�)=���]�$*n>��g��ф���9��R�A;�iE� ��1�C�.�H�h^����4��#�n8�m_��S�Qu��[<P(\^�m}34j%��4n�yUk�:g��II��~�S�É�*u�JE����۳�/(!:�C;̖������K�п�@��MI����R��>�5�c���,G� N�i���l�q��bB�1�p"���5z��E��Ή��[��]�Ǯ�4"�=�]�aA�)�rf�]��6a�ߺ�0'Ԇ��mB#(A����7����ThB#�WTU<�ȏ��!X����_y�Bg�w�I�5�Y.�ZC���f�g�ϛ>��̏����є�u��+��u���6�'�ƻ����Y��a㟸��'M6W=լ��v�1��5ob� !7���4�J��Rx��W)4$/��1�J��1.Ŝ�?rHNp@����J�	�b����Ӯ:B�c��C,�ݦ*�R�JW��hvW9�4�J��c)�a���ܬ�fâ�+��U�]B���%�Dޕ�&���A�f���y�(4e�;��Nʺ(�i_4k����(���1%8o�5�=�b������[N(u4���Ւ���]�؎�֭�'��(!2h�711'�P� �I�.��a��q )�3���2�a.�v�#0�\L���ɷY��tS����ǶM�ySN�v�5�}MFzI��lU�=�Z?��;}8�zTb�c�d4��ؗ�F߿���R)��	3��U����A�-ٟ�B��U�1�<�	�烩:����x�릘��'��B��FƏ7O�EU��������iW�ś�<�.)���'җ��l�s<�e�L'9�$E���˽cm,%"� 4��}j�����\ �����Y��C������1�u���Shc�戰���M ����(�n�l�\�6auWx땲��R@7�x������6�t�m��g�>��� ��7}�W�eAho�?6�Fr+q��o^ ��Hr�٫�s���?V��v�A��<��!�3�.M��$ %�����Z®��ʆ칛A-Rԓ7�7��s�A&Ng�R
����D_�����,ҹ�#��~��cـDZu��W����r��1�[z)�q' �V.���t��C[��;�(���a����D��o�ggV�<d�K�Zݼ�k�#~zE�#��W����^"<H���e�p�e;\�-1Ff��]���Oϕ�*Bp$����0w�6�{�æ���W�����c*Z��eձd���s���e�Sԩz)S(u.�����Ą.>I�����7��j�A\���B���厙�#]H�r�J^F��˭=�Y��[��Ҝq�D[zX���b!y�V������oX�` ��F*X�_&�uo����jʈf�|j-k�WZ���T�nd��(�|��������p o�4��Y8�S	5�O�m���x�J31
D�Ώ�>B.����34k��L�S���gl��
`kfqK^
�b^�J>��JyWs���'��iD8^��]οF��q�#
�|z��C���|�c��'�\��,|���?�"0'oF2tsd+���G�t���J�Xe?�A1�P3��E���xu�l1<.�Pē3]�z�?�0��?⛣,��Ft��U�o��1}d,+up�ţv�M���f�d���� �g�8��#"��7�1���� ���'܂�[v����M�a�xX����`\	3����*dt���y�h�Y�����m�V�Ȫ�&-�r��<�aA�$�'�2��v��0��;��}:�h�/yJ�cҩ>M�:�������� �N���b�m➳j\�BM������ݜ��U���ژ�im:?�l�;[�i_��~���(�j�����=}^+��X�ni�s`����}lY����o��c�g��4�ϒ����\V�Rl@5ř�3���2~9�<<����lji\4��=>�� ��Um����eѹ�%o���ly�+��.��e��0:Iq!bJ�S�D��jG �J'�5|4E�衔�RS�N�Z�EI�~����m�	j����� ��B�M}bۂ(�OR��\~3K�Y�&�JMr(���8�K�q7��Lu��A��2�$7��/�ۋaQ���L�O�uե�������,�[�Ht`��꺔�	%[����*�!D@Q�n��Q>׼ �?���~�����zA�(�XesM�Q���!r��?fX������h�w�#�X�ij"�M��]N�p��E2
 �/�T��g�g�������������"9f�y�G0�۪�]�)7`�y�g o���~=_)A��~�i-���1Ҕ�4��ia �R�غW�w���䳁*r%�d9�7�W��WRVW���#/�!@?l+��I3�%���/���Y�{�r��yL�(��� �+T���,Ѣ,(���G' ��3�ڣ�=C�B�s,&N�a4��Y�u�1�!՟ǜ~�@��6S��>�9�[��7����e�Y>s&q�v� 1gN���k��{[�T�9s�bC�,K�5�
}@�<dNv�ǋ7����y�z��������6l�ep�R�I��P��̶��n�e�6�������L�����zS3e�Hl�6H�	�ʹ��b�]���g4Z�&c����H��$Y����\�f+�����;�b��p�\4'��S~s�Y�Ē�I���nX�L��⭌ˌ�����+�]��i�X�{��&x�[��){;ToE,a��4T��Z�#_
�������A�B�X=�K�r�����n F��*L�u�B���60%�����Q�<d�Od1j35]�J�o�9S@���R������<i?�D��5����L7�.�\���Z��%#�)���F�8\�X��{�l�����G�8R{��7.(T��k����i�����v�.��S(ks��#][�3r<w::�(�Q���"�-ޣ�@�<���5��'G��P�p�^T����[
e��" �D���q?mtIG�&�D�Jzqg����d�,-c�c:l�7����	���
�P	=t��=���r�^�6���i^�bG_ͣ�'8O���~a�vߙ`��uU��x�D�cb�B�ߕD���+��ë>a��_Ω���6n��b�$D2ܒ�{p(i��Iy��}B����̴�1����9̹�6@#
V-�Xb��0Z�ؒi���O:�tޢ�Ȃ�]�x��~�qR��Iy	���W���+h�/��)g�K��x|j����x�XC/*��hUt~��Ȋ,7�K�(R�$6��FiZ`���T�&{9���Զ���G=T�l?����{�7\e��>Np��觘�$K�� Ӹ�<����#��Mv������9�is�)��=��X
�}�|��BG��!��Cu���D�e�ݽ9�PUfG�{b����8�B�%N-n�N���_�Grw�E:r���P�����]�[]�%T��q��×�4���ܼ��OFJ��מg���ָ% 7� �z��C�B��,%���4K���y�,�n�ke��+���~ ��:Kg����D<��)6O�RKq����)�O��_BSy �Uͭ��.�1��.0w�Ɋ��t (��������!������|�K�U-ہ�\��i��JeR�5%� #��&�;�^Q+�臂��'�!�5Ĺ�cK=�ﲌ!�'(. ~��;���s���Z�)R[�Λ���1��ؗ�7���Z��H�]#O7��ֲ��9��>�{��k�Z  ��U�j�����W��3�bΥ]��;}Ю<'R[~;�*:�������+$�[27�o�ʼ��lɨ� �
X,Gco�u�-�"��#��.����d�ĂJ��.߅{9���4�-y����R�6s~L��%!4���V��c����r���;6����S��g�&�>���H��]�_�g`�JJ64��+�p�my�;��M8�k��� ��(=T<L���J7ՄJ`��k'klm��(�c��0�]W����MQ��`��Z-Ѫ?�t�ɋ����W�0.�Ip�K.��(gp��w�*���S�[�m1�Drc�A/��vq�z	c��FWCi0<S\h��]a^�#T��7_�"q��݃�bP���5(��]H-n7��!E_�e���;����Tzn�3��=����Q�e����)Ņ�/�Z}�{�t`TZE�f�O�6F��`������*2�c0p3a6�ɵcJ���I�f�P�t�g�L8�4Ջ�Ji�"|Z`\���H�o�%K�	ş�d��};�N�\�=���毼T~:A�O�Ps�����z��<׌��&��p�S�!�^�~��X����e��j�A3/�ih:�ߑ��v <��b���Hn����x���;-�P(lD�MÉl˻tGn�n���j+����2^�i^�v��������`'�����ߢ�������l����8�o�vY{�`Lڍ�Ԙ9Q��a�O�gG�g�)�k.�
���%Q��|�/��Ы�[~��r6���w;#R�jycTG�����cg�+�	 թ��8���
�:q��B4M���F%/�j}$��z��h'���!�z���0�}Mon{��?��{<�o��oT� ���>����h�j]>Z��OK�sK&�ns���|���F7��L^��M!�Û߬��2Л�66QKx�ۓ/�}Iv@eO�����t�3��Q����tF�vi��\�6H�,�7��v�Ї��<�MEx+�U�֨��^ygq�Zg�_�62�owO���Ff�4��\l7!�E����=��?���!��n//��L��粂j�M��d»uT`Ż�x�~�扠`�O��>�K��&�!][+^X�B���}2\P0P��b��G)l��n���2�9��N�)'�e�2���?���������� �4*�lܨ3�qT�A,;���g��գ�3��U��u�׏���z�`�������jD�,CYX	 ��vmR�SQr���*�~���h�='�O�W���j��#���՘(j�+zJ��v���X<�F�|p،�
~x��*0��O�A��K�ۖ��m8�
UևE���r`8�}�M��>S�cs�W�F�1h����+�)�#�P\�������>��v@\�F���Vc��w��#�3*:}�O�FI�lU�(F�HL�+Ucu��=�@1(�������EQ��E�-�fvBύ�]_�{{a��{�-���z: 0�꧙uX	�����Ʀ|rQ���HӚ�0�,6I�8j�e vLn�\�,�AbLA��u�~7� N���}!2Q�~���5uI���V6o�q��x0D�ƞL��d��h�Nw������K���T<��Hf��[V7[s��5H���K����Ѳb)��$و�6뙣�\�d���3zڜ�ju�$��0�K�nU�Q��3B@O#�%�@,��|`4�'w#��S�|qp��}�,Ot˒o>��7���%N�~h)�Y������0;j�`��eK*�;���3��HO|��R^N�PI�3l_��#ڳWe��Y�\u�!�xm�Z0zF�X�t�w8,$Y��K�F���+K*�F�lDjn�Y�y�����w[�7�>H,����3�3�4gαȾ6 �D�����T�Y�^���2�y�S3yV��,�x��7n晻z�_�����E�U�d/p$_RS��X"ȝ���䒠f���F�m����R��ʪg����&�����7�5Jow�W��g�P�E^P�H��Q���#;[��˪�dZ���y����@���u�C<�µ.��7B����UOr��K,�m'��$G���Sy��J8Kt l�S�Cr�8�|�������������~����A�w�%ܶ!̻�7%��Nը�N�����V6q��c����:� e�[4ǦO�(t׉І�h@�a�V/��V6-��QH+pk""ha�t�h��*�l@'�'C����(�`�gf�a�h8������-=�W�R�*��û��rw�3��;��D��d��7��uul��Α�w�����TP���x�|�vr��oۜT$�&�<=~�|��ɂ{������J:�4ޟ�����#�!8N?�m/�:�xݧ���Gkw#Ȼ��:�S�J��m:��~I�{isQ<��wJR��6mhaq����pخ���f��dfF;2�[:π���}���OA���/@�J:7Ȯq�0@YO�]���K�\Bz;���p���.���BM����~�aI��@������e3�@;���n��h�R��*<�ꅗ�Ǵ0+�Oʤ�ܒ����[�H����'�7j"��=�]���Ћ4�������I�8���l���ua���q�ھA9��jI�z<Ĺ����������.S
a(l��/����è�#�~C��u�6��O��;��F��b�M�Y�:,:�IX-�F�̐�ǀ$LdnCV���j�c����]$�u��7��Di���K�Qi&�����O��?ϔ}�F� Dt>bA*���Y�d�T�o7�l��)����3�̓�X�j��{V���ك>��*%�!a�O�<j�:�!�޹�p[��k�w�KՍ�#G0 a ��-�}���p*���c`i��v�����5l����>ѯ�&�k1�6g�II�3*��h�G'��5)`��eok�)8��������v�C�T�=(�L_�d��x�)N ��CT��g�S*~ݸ�t�����1��^�xe, c �Q�(�A?��S2��Zu$�f<�Q�e\�Z�L�h� %(R�>F���<=3���!m�_+m �bL�<�s�p��K��b����&E��TFu�yt�v�΀�p��$���h������g|�$6�����h�����J�����T�o���	�O���ː;H�X����D�T��U���6rn���q���GOĂ����9��NJ��!��/wx��Z͝F��S�WLc|�J9 ��K��w���Ih O5G���tj{u��+;�P���	~�����E�v����eRS�݌t�>˃��,�3ѷ9S:���?�*k���z{�[с���>yz�K���O�ͻ���^�C���ta���($�|#������S@��������������BT��O�^�W�6�I�vYa����@����G�m�c�@�c~�ɰ8�\��a����K��]A32̖�M�A�߬�d4��?]ζ�hv�_�ȕ
���x/��5�Q�}iZR�%$�&�ђ�j�O	lł�,��Q �D���)laS�"?��1^�<R�T{�����e�#�=
z���L��wP{��t�_/����y ��Dt� ����41�ܞ-{��ْ��˴0?�7���!���.K�:AN����֓��a�����mj�؋gZOl�Nv�0Ap^&��i����0;zb
0*1YCʙ�}l�����*�C=ES*?�y�����`g�7�;�Q2��-x�r9Ap��rukul����t���P��j��[��v��Q�XH@���d�jN�;z�zZܢH
3�6^F�-؝�KGG^[R�����Y�Y�}&�~|�ta�$�ʧFa�,��� 3g�9��h�0q}V���8��YO��I3����{��F#�іHɅ�4�/v��ƀ�wF�i@y�G>�^8#���*2n"�w�:1���*=�,O�T��ky3?���ϥ�<��?�]c_ZT��</��]|rw�W&Ў����3�{<_�*/�L��_mˠ����G�8��w��_�@aP�!y�Tpq}G�,�b8��_�w|���̒�ʱG���#M��me�_�iY�&i�g��H�b}�k���m� E���:A]k	�)��U:�:�;�K�ie�o^;��$�(���؂؂w��-`�Ƭ5<��
��%�к�V��s�B.�9���X=�پ�1rg�]2��,c")�+�fw�Q_F�X�G��c����RAAm��C'��5 �l z�
��u���N0��N��&`�x��Za|<��D�T OBh{R��p�G�{��JH7[c"�� ���z���� 5�jݯI ��q�k��)=�]�1��R���xB�թ��8Y���z�-&���XJ��g��Q��.�pS��?�x�<$(��kb� ��NKO�;�wO��7�-ߺ,9e/�`o �z�&
5��*O���4T�jZ���.vٵ��,�X���������hL~T��.����wml�ǯ�X_�AQ#3�Y����Uȉ�D��◄tN�km�Jw�|`���Qh�[�����tB��������C3/���������7�K�Ӎ	w��?�}�y�*������T͐iB]ϣ����_F����{W��/�J5�mG��,�����^�b���T�*���+I-����oK]�Vi*��d��� �� �}L�:�:�
L�u(�$.}��Z�S5|�N�L~����"�ij����GW��F����G_@ /+��9*�@J��mS	��[�I�SK��~�����;�3��/��紵��y�K�W��pئE=��O���u�'��<l��lg#���i>�,KS�I�[0w�|B�}�9�8��W������q�d���4�앻�����C)�ɦg��d�&y���a/��PM%Ly:Ql;i�F�"U|e�ڝЬ6�q-�[?3�'h��M be����5�K0m��D�$�U8�vXE~���~p>|f��Q�8��[8\�V���E%�w�܈����I��\�2������ΰuzCY4��6ApZ�LT��{����`�m�Qu۾��l��x�sR�$^{E��X��Sj�}�n<��^`<18J�(�1Ѻ�K�Q��4�M;`Yo�H �񝜷 ���nlYi��~t:m:Z}zA3��l�@��.��ӷů����*RFi�,*����߽��d0�A�`�ȗ�演�̛&l���sAY\Yb�iC�!%}@��5�z{���F�t�X_r@�sț���旃�r� ��r�^5�	�9��8'��7Ť�� iN�:��J�6�q볚v�tW������v�y&�V&��d�����ڗ�
��8�MԼ�M���ӎV
�W�"�M�����(W<L���s�&H	�"Nm������Y�M �Ϳ0���+8eb���~e�XŸ�	HCh�EL�2}�{�?\���Y'��Q������Z�L�ݢ>���M�럒�E��j$o+m@�%HI��m �PV��Y^����5NQ9�R늏q�8�eW�e���;� �L]�5��q�F�u�O#��9C�RR�F������j�QtP��¤�]Qj_w�5��������e2 �B� 9�\�9�<�����MUt'��kri%r��~��;o�kp%Why�8JXHxa��|S��M�	�a��zX���(�g���Z��U��5T�#�8i�~]5��, dR�{
P�k�(���l�Q�������Ide}è�0���.�ot/��ռy!�-�4r��)Q짮;����L6�Y�K��R�b�N���-h�n�e���]`�S�`A�ҷA�=����������
K2��\X�lS;�A�9X�oUF\��V�T � >�]���A�X��GA	�՞�2���^k�Qn�Ӝ,���B�4�P����O�������+A� �t�Ż�����#���0�����p�h�g"w<f5)����K�-�U�76�h�\�0�u�����_k��b42����S}�s���ʟ�d@�Y�l�:E/����W���z����ub���tm)5���Rp�;��x/$� o�l���l�����~OAr�{���F�"+8-�>��)����M�+��z)/��G��s��W���FL�i\�{ʀB�l���>6�%m�Ǧ���s��C@��������6�851��'^qe������C������U`[�tYhv��ڷ#̢7<���j�����E���7^U����&=�#�,Xa�+Pu�;陱{,�$\��*Yo<��	,����$@vj�V��D�i^�N�*�R0Qv���xbs AYt������a@��W{�޳�V%.C90(�[$N����3������QB�.ܪ����$�F�G%� ��� �jz�]c=�[1�d�N��-��w��;~�x���㣸P��j�,�4kg����		�w�:g5�����C2���MlP<'G L�@��h���uv��4��;�OL�ˡ'���M!B�i����Z��x5�cb���Ѥ0݋L�ec�����V���o����\��6Ù�:еfD�_���ԕJ�P�l �G,=c5#Ǉk�g��VCqLL)^C��L�Ҁ|�eh-SnkK��v��~��8�B%��J� �Eu��8nz����ͻ����m��0+XО��@�V:L���ǊV�nk�Vc����G� FT�.{�*ͯ�o����ezq��di���׌�κ*v7��D����O&R�~�)A��W����hc�?)�!^h�J����1��N��cu$<E��4.tR����x#&����o&Z�LMt#�qZ�K"�\s��(�0Wuyd���h��4���1$E�2�w��'�d��0�J�`��B$lU�W�,4��Ǚ���n+ =��g��B�Zhv�������y�[������9F0:���4Ë��gъnՀT�� ~��6
���jL$:��e��9�^������wC0T����E�Km�`X!ɚU#�զdLZd4���2Q#
Bb�n�N���/�+v�y��7����N�Or�%��.��jN�^搈����O���Ŧ�0q�z˲qqao�ى20��w��ųI���U�H��ާ���'�*%�¶�S���ya;^3�
��#P�ʺ�N�M���ָ>�@ \8��4�_��O�=xL�����Q)c�xW�D��'��:% /�O�?hb�8��A�5��Hk�I��4��c������րe��O!� O�^B�xX�՝�*��Z7�.�ꕼN鹇s�M��[|�G�笚��0���5�,�bRw�V�S*Ts����Qq�o:9��U�dy��G|��H<�l�rX��-����S�[�Ŭ��k/n��3�rG*櫜t��h޶ۧ'R��j����p/���`�>4�pv��lG&6Ni��XU�R�A�P,H;8��[����I�p�������*��q��
Bt�>%5r�v�z�]��+�RP�$r�f�VЉ)���נǏ�"��.��p��!0{,;���O;R�8<�}�c��Z0-H*k�_���8}�\�B���������4~�.��4�~�$?W�ێ�����b�LX$�G�ph��e��A{�5A��eI0��}A
��~��dqd>݊)��:ۛ~C��1�>�3�~�z��Ţ���}���H�O����oW���2�������q������5��-"�do� |���L�~eX���N��x\�Cg�[ˣO���T�K�ԈM%�(frԷ"p����-��0G[ at*I�:���	�yD��*�^j�6˨f�ds�����T6�"�. د/'j	��!2 �5�4��.+t��~W�2Ro3����7׳�W��N
����i�O  <5A�T���D f��+�Ƅ3���A+�l��ґ�j�#*���+�Q�����k4
�[=Y�����`c�kJ���'�L:��4/aЯ�;�^{Z�a];|q^��}��v[V(��2���9�Ո�m��MOrk�|<%d��n^�l-r^0z��?As�-q�N���*5P��I�0y\���wCoE�˱Tp.kFsI�q�i��&�@<�U��Yd����p�V�8b����ơ� e��s��V���FC�t��&�E��Zz�q��ֆECE�ΫK_�v@��)_��*um!��ң�ňk~&%'�����4�#��2��/������ft�� S�:�☣�N[y1}��_��b���.��ӂ�����{�.�[����ǧ*�P�A2�g��r���^\ݿ%��>�ץR'8R'���;� ~�SD�q�[�IN��p�P��I�~�`����LM�PT3w�y��� #G8I���X��um�X�4B�8(��5щ���ݤ���xL�L�L����O��HU�s������ɦ�κ���_��0ЪU��/zoε���骇�0\/�8�4�tC���>4X~*Ά�4�iB�~�0�*-ϸ'q�m�:�c{����e��W�V�8ru8?b1���Ǿ��o��A��B�V*�3{�I5Z�4j�6V�ʰ�!��fU�!#6�ʘl.~ǃ�!�?"]��� &���ħ��F5��g�ʟU7�$_{RNm���4��H�L�he�����8��.�j��h�%�P*D%�D"��~�8���R���N9�'.�s�)�