��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`����<�V0`Q��ťɊ#�MwU�P�X���s��j8C��eZH�4�L���M��-oi佴���y�w��KX2���M��f�� rF���O`)���3������Ў��T����.���FN�Oݯ�����U��&~��Ōı�r�j���'���6��`bFM,��g:8���?<p�U+�k|YwIj�F�C�&�5�v�0��c���8�N枫?K���|څ�m�!�����8z���|[�pz�<�����ާ\�[s���J�0���S��f`$�z�>$��>H�{`��s �=Os��a��73ݯ5���N�sx�� &��n��z������t���������n��#/r���y�a�*ݲw��k䥍mA�s�\�ٷع��~�{5q�:��jo#w��AI���Ԃ�j��)w�92^����#g婾�H��i��I��r}����GmK��ک�7�@3ꮕY�	��=�"��`���wOن6��q˳��A	�[@��q�f�M���(��W|N���݋���ť�,C��G(Trzh��:����B����h&�p)`��JD� R��������;Y�o(�mawD$���6Hm��t~�I�����3�&z�D	g�g ��>�?�θf0S��bNG�]�=�P}�XY~�aY�ߠ;��I�
���h�ps�£�>X�_ؽ[ق7���(c=�=R��KX��iE�ݣQ��M���A�m��Q�f�dd���v��J.�yqoy���x%��y̸۷rnC��dD\t��w=�l���q�' fȞβON|I��P��ۣ')���C	�i�<8&���dq d�,1-�U�3�����[d�x�����Ӛ�1�F�i�2ݓ���7�(c��C�f�;R�<�l������{(����#s&Gw��)V;˃�W��v3���b�u�T�"���� ��Ep�C@y��Ѯ����)�\�H� 6��!B�c"j��_���r@�4Jø���-^6#*��S�!3zo�z��G�4�@�fa�/L������ç!k���囿$�̧�-m��9�yҧ� V.��0l��o��\`���[;]S��$�#h�GgSz�`Z0(�p��ȸ�~�(���c,w@!��#����|�,���<3M������tI��Zڅ��,�~�zp؝�T���Ϲ�sM�h�z�)��m��b���mB?u5�.��x� ��i���+�p�ü�%S�/��z�A�lXTPx�W[9�{o�Z���ch����`P��z���ZJ6�%��<�j2�?@�tߜը橠՝��	<�>硛�4��>�����-�b+�,�?�l�7��W���ԟFm.Y�V]]�f��IvM�1�m2�l$gk'�J���>7�%���ЖOv�{w7#{�{�HoK�
��-�����bI�$b^�H#����ۘ�(~�}�yB=ȿ�#s ��ܓ�N�\��M����B���Qf3I��6ݡH����PïiR�z}��@��L0y�56�̺�a��H�ê�b� �P5��N����_ڻg�T7Q�W�A�Idן(�6r� �vm�A�`J㫇m�C��?�_ݓ��-g�r.H0먀�zK�>�s�:~�u$Z2ѓ�C�&����&;_8�	�\b�O|	�Qu�kH�na�d�0���l��q6��J�0��X���r���s��]�-Z �}̽��W8,y�G�̡AҜ*�};[0��k�.�\�G�$��̆�q*�4ڬ�G�@�V�Q���?=�j��c�:9�EJv�ǃ�B���wE��|���}��|���䐦�	���F�%w�.���$i�;a$�S�U�pE*�!�T�1�zI�g_Z+E �)eAş��@�&��3�`��O���MZ�1�d�c��Fvj���0- �T�0q3:�>8�5��fcelٗmX�v�r�ѵ�:)O�����0���?+�wF�<��]sT���Te�b�{By�w6#")^�6y AQ���� �k�m�����ՠ���C?���B��u�ds�#�Ѹ�֢G��0��פI�ѭ��X�K���"�1��8$���ok?Y\]�φ�<xک��T�1޳	F�Wt١�fhYS6Wkd��`���L���m�jZb8�[�<���Aª� <�Å�*�˛ yp�&w� ��'J��%��v�*�G3-����t�z3�^c���cԽJ�`��6�܂��0��Pah�����١�UT<�H2��Җ��2y���O�B =VJ~$����|�b�~��	��Q�t��w;��Y���(!e��,���;���U곬+�#�?R�����4��Z��j����j�E�uP{Dgx���X�3`]u�~w2�1�"qߑ@�D��(7��_=���t�8!����(�b���U�YEY��[:.?5���� �)�|��?5qՃ����u�ZO�d+3&a���k��ٿ9A��j\+�x�K�'X�^�1B�9��(e ��S�{��t�y���^ �<���״
