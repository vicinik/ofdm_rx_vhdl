-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SX1gvrVUQF6pDOqBBoY4ItmObi3C6sFMmGbx8tSQPD+WirR1x3+xcNrI+cc5ACCnPcLbI2p3UqK3
MzIVRW9xrOcVroEqKHXQLmjTxkJ888T9IzuOXkyqoT/4iunOMUYAEfoSHJdAO78rlG5quOUuhnNT
IoB1TjB4Ig8Ki3Rstmos/vD3Vzf93XOfFD3Gavu0WWl3j2N4vHS+6kmSPol+bDVQmuhr0ZSEO+c+
QihS5nE6tpTLHJ7f385JylEdYNj6OnIEcF/0ePC6oCMEl5RJT0BIGapfCj1agcyn0BgCtVK9cXH4
Hf1L8+iAcNmcAz5QDP2YeOuBNpjlVkErWjHoDg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 56272)
`protect data_block
4UGj6FMsRIYd82x/0xAuLuvPra/tdktcjyBYVc0vChSqzIIF98JmdFkuKTJmMQwCRgtyF8JpnwMV
27lo/e3kLwVh1nNt62Hk1Eq5DYNmk3vAros5fD4X9QwOa+LNT0ctmXhFRJSLReKbFbjP5rP+ZbKk
Aa5/xqx2007k0baI8mk3p7MoNW8k7e5mdNtCJ5aHyf1dTb6Z+qvYWZRw2RAwL90bz00yBFyOl3lN
H3Oq/fCcU881VGrmZ+fkmxCY/r06spfYwlDOjHC6bqkhSyRPBm+6qqWWCAEPtWqv1GLFLQ9Fw2kp
BEKIzwOg4Ar71KOqAMki1RQMII+kbJ1C1XU3cKCsDz2Xa6wFDg7/OH5S6IEgLsO0WmjNwmqHhXoY
rWDLjYhHBJ6xyWeEyP9fWkSDXQtMOlHAYTm6JYF13/kY/DNvW6oPBTL11pIRv3RLv2ISXQPsQm6Z
Kwhjf8uiFflNnTU/Y74eOhxfp7MPQFjDW/OSoVCx0FO9JPrYRy2buObmv5FLIhXSycI0V9sjBU/I
xraWbDR0g6hksFM2Xc0YzRNL5yBuHxfNTmcqQhMQOkMQIUwp7rjwGUAey+qvRadTgnXrZkhCo5qZ
qGaXjAqCrljh6atTKcjQwg8dViJbXMKkT+afmnJb7RnIBkZQ6G6SvvJ3kiEJip6JUKAYcWvhC0K4
8WYx/10fYkcEE+aOaF0V7+I6TwpXSLhKldfzQpIHDQWlDtl4vNDoxl2U85WaERFP0OCs7NvTm4uX
cP/sYanvx9Utw6mPKEqsr+i1RIM04CyZ9JzxJ1oyE+0fjSd0L3389HJAOUeq8rxBexYB1f1UBFj3
BDYDlRnSCCAvzzTomQjvsLFZN6PVa1VcCq+8V9HagkaObZeQ7RqXbWoHB5EzBbZdeGWdmNqcGBhr
T+HNriqOYujv8PBPG6higajAYq48fw0IBCY2rpzCbD2F4SbOx5AeRxn9y3kPu+sXL0x07n2UwRS4
8nxJxivEeAp4oYqCpsQd+EXvPLObMWtQlz4ASt/rXhAuyFZ4WBE3h0DL55oifqNm0bGPK7K8S1hs
DkiH8FXh8pB4Hj56AoDaAKKdG6IkaZ4sZKDaVKCXo1Wf+CWhi/RVGYRAjztfBjFfMx/Q/VaUP1vd
Eoy9scKO66RzZ6Mu7rqi8W2eMG3ZAMAq1WJsujp4XYuR/msT6OqibBfAr12kZMtSDChElkGm+urJ
Yx+K6IMmxtJ9OOpQxOU/47eBxrgGYbMLUchO/jKOwPL/U3UA945+li7ClLYEpZa1yC/Owj+dIgEG
nJA33EOC62+yXoNuNqO3utMTjaYk1adtv5W5GEo2EEKLHsDw/EteKTst8zyAlUhr6h5T72EKN/N5
j+zCsRB/Ekn+wl23JVvQrNVYLWKhrH7AUTXodWBiXQlvep6uHyIddn8jCyPDD+padAdOUDx+FKs8
DQSDZOkFbrztIr6IpiZKIoivEgJwE252ZUeVXA9VTSXUFyx1Vdjs8wlm6xGIWyDJRM7C63vsMmSF
ZLiE92MPO9Pxw7OnfSM8HG7kQ41PFKvjHDeOywkwBEZrhlVqDC6bOAG/i6CW8NhvVvjFKJk5sgTz
0mDJ8Pqsg3j4+3duBkrw3LsQ7l6GlMfATWJXHbT0x7lCfFjW31IiWPaTt8XJ7WezoLQ6Vx5CoAgm
t6qTTbAWRCSfYURMd/CZJ+Olhd/ThFitbAe65Eml0rw748tPt72yqUmWaTWMYqqu17AH/hKwfpKt
s0OsNQGyqaHboLLFEtikhGOYhkWizP6Q506txoc6qP01C3XcZzIC2erW4rDLJ+vAgrYit6JMiNL4
+Bas3d1MD6rDLN5bLCXaDp2+sXM9kht8JRy+cBn1cP3JA5vKWuh5ARUREfTNPA1ihuNc5mbFMGw+
86lEMSKoEEZQudP1wC5SCcXMl47yAOb2Jyz4UvGzAlAnWBg1W62wYWZGcuuUa08dNAwE68f1yZST
oNHB4dYZuLqET3fZ2n1EPtnXHh6M07UQzFFaXQpvHO1nouuqGh+sNAkg3wu9ueU2Oet7pl5M4522
5y5S+X1Lq5EtIZXOTUOY1ruKzzmRV6acUVqRgEl3LmFhZ7M/6LtUgrKw2cPxteLrvmR+crpYlm8L
t3vxVRJYAuhbDLlKNzPVIauYpCDpvpNsjyFaxtkCb4kKGL2HatX31o5/lxNaouWhX5uMnB7Cw0Ge
kd1c5Pu3EdO/Q2SVmSAt4tDqC0pUcECbt43rbWsjwf76h0VAAxURjX5/o89KJnvlBTmVrXhm6101
PXOumNSwPsAqxaQRqCmFu3HLIoM5DT3Ae7en4c0RXMCyCAaNDZRWomQ+Xr8pqlgwwbYg4BPGX2pJ
Q1FntunU05iDvtMKUyLJQcf99w5Vp5vxDNAa+xu3/UUOgv+nFKdr1Opx5GhG9eeLxjaW7hX44rbe
GgYub1S5drJbkKSl/FfFm95y8kSNLFljRTBFX/V5loWjOcoeovVrLrHm4Ee7zqjXAijqVKND+Bx3
9vsNYdX+dfM44LvSZ7peZRpOmJNjEjP7AacFB65p3LtZbpFydO9VOI2GFGMSUb93NdtmQnLDXU7v
633Z21JuPGsR3k3qA5yb1Lgk8/F7hcPG+CqwHV9oiQmvwdSypeC5QXjgpmGxF/bU9ZrX4hPYsPgq
Hli0y/GAkTLuwYzuf8rHFLFJt/tZtCY916KNPn8daF6jtV4h3EP39la34HQsWJys/vC0VM21lttJ
sRWczeBe2LBzMiUc0wRS2YmYRlYCrGxY4TewVtHZ0NAB/3a0z+utTeMRWANkH7OQYWfU+n+TS0cF
pWJkvrdVo1zmdLph6Dmy26kvdEpOWgYn30eBNLmA8XcVxKZjDdybygua+4tPy7B9SnWQMycQpJy4
dX6mWuIPMq+Bbw7PieIA/s32m2wyOr3fNshe2iC4Ky2OMKR9QYi/RtglYZ0NV94FDA9qmgOxZYQB
nRggSr9bic4mkulattHqHyCx2+2CUahntqrSMycXxLOWTVYMxrIFfVEaoP5k9i31GE1JbjLU8bfD
vyNKnIca5LzCeOE2+GRaohrYwMIfwaHzGeE+S9P0jO43JCUm8+bfos0oIeOGEe/n8yMox3PIopFJ
A9hGZ7esHR8BbDpfbxgobM0H3M5LJFPtaVZfCkK88fUsIZlN6XXAgoArx7IiOeA0ZBYoxLUgWOCe
UEomabV9qzOHr5mX97o/p5ZffnTqNaY7V7jhvyPIWieFrxJaWQR9Xwzm/uSld29peWYETxCvsKvl
nyzsuzmSXZOhugUk/4ymkBpOT/xRu1EVKD1X4hgH9IB19RsKpiU5LH9MUIodOPNSWohdT4s4TZNU
gF8fzxlVFY18DctkYxT9/46PBICiMJ3Zb7cC5eBH6iS5YqnMfNqnXY4Whkpr8gtG5NN6B9FOY/g6
o0qjF90ZILFdZVCGm/IFs1LJVkxxOG0e0EjvSVMiwZSdGyNphvq8bcfOo6DRZZiqRwYBNAho03wL
EeeeUewHw3ncQNL6EeEqN6txb3BqBdB3q1re4YhcA6n4Slr0egiP8BbaSxaBMNtLVmojdsp+fnn6
YsZiQMYgxdJVGtLXxGFZu+Cz7CXlbgxB1mZv4A2MW+OoTZWI6OgwdUIi6lbPfzgHWv6VS4lWL3Ky
FtL4VZPAe/5w+w3ecb+pzjeduUY9A5vn+E55J2St9s1BRqH7ARqLuZ+cxxOeHx4my0epzrGlx8M0
uzW68f0PZHJ58HaVHxVl4hXzqXuQ29fEx+V9FQTqEWZxof0ibZl6cbSzbD8oHjQQXMDalZt8fNSt
qTelhWSDp2ISn4O5AM+UH3pHgVL/Ew2tKiVhmIX7K0YVs3im1dEYH437CcKaRSwUYIE/gihQkr6S
aVbcldd+3GGp37jwN/uD6u2liMsCOXzTKFa2WLiHVJuXdU8WwJNTMn15ESiohSLOe9j4eHEY41ZH
PK8eNq7X+zreah2XnTWUyPgBNm+Bgter+c4Op++ZKh5fZZNz2ZxpmvLvuVwfbRo4gr02UcLzLGbn
NQMuaoYK1wgokjKsE28Dqdubv6EnRlTyTeditLhWaL6YAG62BpUxv3mxqPmKGhw7Wloop873LpoX
0M1zF2WJ1QzdBtr48lsPtL5LvL8VcGAP7LTvSJc3LBN15CenS6mrAPaoHLF9YTGNr88rmMX66EuK
Q/nR/Phy3OZWDexpdxDHXODAQAqXgMlSY5ZL22vrhBb+qUvXFRxHZVGj788g/+jiMfF6MFYB8rXC
S5qeJ7gowp/ekdApJTZu4Ct8/6dq44HwR8KvJpvXr47aUGPAz9AWOdyhZJCqFtKxHk9MNd3wZCCD
Do+kIENKaf+H+JAK0aQNPmR6EUHSrjgAq5ybeZKm3c6ngSn6ngVMvqO+PRNgdN2ZrCSFGprJnkQa
xQa5u2Yp4IzVU9agv+NwdR8c4gChUPC9LSMZE/Ka1bXZuUkLKHfJhjdJddujB3+VAdw75Ui122HA
GxZTJJDx6kP7KvYi0VoBcSfK4M7Tv6iBzoc0g3h5GUqwyTLH4MEkzfxANqa24arRj4AY8jERs5Zv
mgxQ/20h0sBl4FPZ8nnQdnjDFzG+dw3v9wEzN9aEvBZ7bpPwdBnorQ1KOoaLYqTEm+46qsZWD4PQ
3Liy5Vr6suFHpqYZjGNlu3yy5BJXv4skKbLeOgY232x2orDBF2A2wA0ZjFF1e2fxEHEbZUdgzHF2
HvDGEzhuNRyxoxvX+/7ogdlZeKAuen7vMnPP9tJfVEMrSXWPymy5hTTTQZNjAal79YrTx55Wjkr1
WiZ3LWqjxJFggC2NqxCcEDijhsFAuOjHdY0J0vAIOLkEb2hC23wrDJcFKKQZchjYQkpRXuGbfPxg
igG1Vugx7QZkyWJfcy63HqsUHvLQOzroFajzjEgFUxrVbABWiHGxFQo8mv1ReryZEt3p66rFXy4p
dqK2acnmCyqkKGyZ4NBeH75lU7acv2dsTEkdF6SSaouZp3HvGL+brgIgFs8vDTdoHDJ5y24eabAK
T1cAs1+Z32GQw69sSjtPMslhkF/7Rdr3f+sMAFYmZASQet/uwHzPRCEUSp3lfD+RGq7cI265vgnm
XQOcZwMpYgBf6g2W+cmx+ngHWLoHM2hwIrwtNgdc4T46O2K+Iv7qHC+FO/8yMkaJnT76XWWRPk3F
jcqs+lnHsjYYjnbYwBHCjex1qUY8ZTQ7bdJTuw0VQPXecj1EcxKSpXmBVjoVeucTiy7A0Ds6QfEz
eB+JoR+b3ZLhSjGg8Qhnq1nWVHD7XsG8X1W/hfjZn2S9WwQuNIMJSKsqWwjkcAhLIWVv8n8REX/3
miYw76BShCHVJhDm76hWYssXV3Fs/mV8h6vFiooU7VD6xISIGWwIIQB5XhXjDzdBUvl+/lcaZw/H
PfyLVkK3IGsmroAEQGQb7FYn1hs8gteFzWBOa4f3FXcIIyIqtZJ4AzgqAjOD7r75CqEDMwwcikDv
QCvtCj8D1dOvQhR0TB36iyx7I4N0SwAm05eqnPv+AWWBIZMVSTgPqyLF4VmfQ5Mp+i7tT8y1V8OI
SSYpMX+AYDEd7fX6Bwwbb1CH284g0rz2uWeR9cJQVtKj2hE29/wkYNz1Z3HFdrEdGNaCJuAzPZKx
J1Sq+dNTx+d5wMfkBIL8UgjErFXKqN0tEDued1mikP4qXgYxhWa02FBXB1szkIpNmdYYj36yp/GP
Jc43H+VZtBJP7gI0VBLiTxkT5FOrNQxl0+RBlS6U8PuLWxH9R2/135QxgSBxbN0uwHpOmWnPrX39
5AyNUZ6baewW4laXe4VmAgySSKUkeGeqlZv/Z9guC2jn9z2KxspmTvKY011Is/qLupNWRi8IKRe+
yHtf4RQK4g781m1K24FDanmwfOpI+cpqeEuslki1uuAcweHN0zF0bNiyRY8J0koWn1Bnc1CLPl0q
XbSTJYMlaMC7FUdRC/4hWXil39TTyp1VXRWBK1uwKoErGEsULoxl4a/A8hRlepTmSMngk6ata0qE
0B4PuCHYXMj6naK+8N8sFctXln7Xtg2Ows4t6bWjBSdyznTbHRsiKkmJU5OvCI3OmOq1vW8LmTSm
t2RbLzGpkmao5imbBKjf0oZiGK/EEdunmJaKhSwfOu0XyQl/k0AIxCTvpFlIbD/EjNAnQCHgxiet
SQc0Y1nsla+95pe9cAXNGUKxhEM/BKHPcawKiNlp1hLjDMXd/KKmmG60N3czpD8o/guurDvzt5TA
Fy9qoRsE8SyN3ol/g9+b1GYUBgz/F9LaW7VucQ6OfFW01okOqfUf5hz5qziXyQtO7vKKlnIGIHrb
jZ0N9E+R36XFAPErifVsTwoCc/3ijVtY6t1lg63kzaOxBgo8ox5TvDl8AXTvY58iJbX5XjkxmU1D
DdRPnXl9a78SCF/3EMC00beKKMvFsdywZBMc/ZZYbzH5RvgZ+GenQTO7fewcu17nIaHwctGEnwju
0dDELohSvl3NhaK7LLbZl+yMO6UQwNcs72VHCud9y2SlvZf3MdGcoroQQXfdXrBSXSNRBGaaLXmA
6+rSfcuCb7527HqW9PbMdd6r1ezxa0y6HeSuj0lIdn/h/4DsoGeshU447EFqLmanieLNRkju0pS4
hkU1XZDVCqyoc63Rfkp3CafSQUdEfceoxGgqiwr5hStI1qIAsER6HxXVKIrCAxRqIfOf8/RIrmjY
aw4l+1T5xaM17jP9Hmk+L88dmOMHJotF/ZFm/Df2+hRDku93S+dDHKMaP1DMzcXSpjWpEzGwQF8g
g0Z52o3vNmf67lkHutCBoYWYzUu23zntJ8pRbahks4I9B+V3S4dKSf2hbzDYAb+RaOaqbRN19cUv
nmaPQpnxlwOwxSNX33VhmnLENAwD06Tr4CxGajuIjlQBvr9DkcpC/OSxCeqMv8ZM6lLftgtKtNrp
ZOFZvDggtzuObNgeukeYDhPT5o7d+mXMY3O2UAKIu4BvBtoVEZRI/pstYCBmyh8xhJm9zwaF9Sgl
KFirQbGlkKV5C+L3kx9kZqhQmLgRJczif4SUn8RsdSrnqx65C33v/Eexr+1GlaT15erTlf2QkZuJ
RM/NQISZRzfZEEhRKgZgX3LBzTbKYE3f4XfbEQFY2hdk4M8nm3y3+rw3r0KRAzv41AFnv2F6astu
SJVTwz2RvLhCzIy/VEagJ6VLsHwT0h5qw+Yn+9bqtHoO1qffUhhcb3u638DT8mypn1CfdEZXOV6O
rmKFkkTLBfuhoDgeiJ5KA973K5eeKU18YCvhF1wt6hggCdVJGzlbNhrQnRT0+W7cqzbxHSLtzmWj
XV+S82q45c6ukZNLjHs7TTiSO51wleukhjKX8cPA2V4ntBYcVDW27ioEQGV2fGdTQDzNp4U2cfWW
+u4+wPlMafQvvCRgW2oG6hK6vTJlgv8c2KKU2UbmwmcA5N1S9zkJJrGa3wIcX7XqYBo7vw8mGcTY
e4LYCIWPn45187ciR8lWwmRS7N4yduJOAASjB7ozZFQ83kYyAtJ8eiRbUIq4qERbBDMy64O/a7dg
DMZFL4JQcQJ10rxtbQtvQD6KS3NGfucu+vxhgI9kxwDrCDnRmr07zY08Tg95ZIzwAhiKmn2eQ8h5
xedfo+IzPwEof+zoBcPI26GAF8/wZOrpAzwu87+n6KBnjOnq1W8cFwEjJsKRLv16CelGPzrme2YM
rPCGJNOPmfA7gopaRB3NQhEb1FtwM2nzMmCANdt+/Jqgr+buz9uTjRGoF5IYSJiH8yat1X8M/JLd
iI94/qvYmy1qdUEVXFw58g4Bup9zq73P624LZhbw6ZLovn8NIxarIL+yHnssEcMiFgsOlO89r2JC
0qIBpmMDXY4seGfuIcakZH6OVHYIutChCoaWL52MsccquhDh4izuPAMxbsVA2qH2r31xJLZKkFdV
V6n3nl/RcW0VxYMhDxOlVnywQYczGY3avyw7kitYQq/Goyluum2agANIYf+z7avUAy5YIUp8DOej
kLNFMZyO1li1MVVri2DaCUUNHty3uJPcx9pNVDhqahPmYPNoVq0da5sBGaFiiHsaKkcEGGgXRddr
JC9Wh+RwwpCvZks4r3GX0bbkW351UiiYZpU32iqs0zymbVp3SLTz/UfHQVDkLTCgOfQ1WZf4vl7m
QvcWChwwJ0OFwUFY+hWbuvHxb7VMiMXuIVp6r3L+uU5p2omclmJ3Z9muqgJmWjMG5mNDFa+m+1Oo
3m8sNNBz6n7rMuSzreqtbRH7OUcsv473QgnPcw5ikSe27W7CNsOeSnL6/HpqE3KUVHUkvi1lJryx
SO066f+hx3Dj434P+wimaE5n5BP1S8dOLTLVVs2ffU/w39Le3F6Ov9tXKmAIHROv9GIG/X9X8Ooc
lOeMzVRG4zqYMBitQ79R9UyoafCN4DlGyydsUGzn3/vCYTJWw5OlSHMtNiohCx60Be2HXBQ8/vKy
6dvu0UQl6Ecx2ylbBxZTQdR50x9AjP6u03U56KJHjMVRl7RAWchnA2Wh402PCY/twds9t+gdsit4
wnniJ4CTTVjTF+WX4vig4V8EpfEmxnkIloSeUCnLPF8lCImDiRnNP89nyiCYzi/9188LgTBom16k
d2u6AiGqMVbVnXQuSIgo0Zb0eMXBdXI0RcnvJPE1qDWjU9QHaUl+m3R91EhZnXOfaxiLT4omRpBd
TPPfn6/TpE7PvOvYWTmTtoJcY/ils5BE6cI668ZBo4hzFoLCnSQxCyqZrTVy2uSoZLfHKj8k7fTD
PjEpklb/6r1RP0WHy5VLUVZN6rNEyYgcEdKyPrmvXHi927qzI9ozG5g4i6cPHCb4SJ2pbZaeSL0a
PgIgauJcTwJb1D6dBsquKklYn/aPMVj9qeRQqvGS/V4UkSlWdQhszcslJRnkhgCsG6bsi5RWHrIn
35ZhKCaOqgCGHN9+hWG60/tuRuw1IiPZeZKzmLmLKOhhSRc9NFXqqxSbVAlqxrni/5Hp8JfI4R9E
a39QTC4XWnWHoH0qVr/+uuN/YthHS79BAydaMF9J04vmIGxqbL+r2WeQHkqx/HpGSvfBbJXmrWv6
57hdZvwW0YdmfwE52wNowb3yMuEf9TRxV5cAf1oKPE4b1YRT4gwp0oQua+VM+jlFH+SESrGgyMCx
yeCHV+Jzjntr8goUGx5S9KRiwaYEFc2/YcjiMrkQdFgl1KFgMNs9pWSlYCM9fbJ4UqDANQyZVPvl
FZ2rNjhVQHn9s+no/EqZHHwy2MpWSE8r4Dzv1DEuCyGFw8V8IGa4ahKV+Lq1rETlGPRt24GGAbc5
oyfrCl9bmd9ZOI8bzhOANg4lXnfXtN2n5RFucgsL2LPniu75KdwA3stKY3sF7YpkzBX+rm96cPVr
2xf0gN47k/w3M+NOMBeBuIm2MESsruNuuYbEfi2eFnow3UmZk4ThPks4QetKZW5hSxTCGXp9b4eW
161lim93EAm1VaxS35lUZMZR3EKqgXQNxmymReLlW0S/c9D7f5xqXmVOezJUvTI8XfhZy6R4SC7K
GPpdylb0OAZxzLJldJZlVlstwobSuc7uglP6O9kxiYsrNCE8SCW8nN8P4NKr5OZJjpTOviPUgbci
2tHysKJKHX6v7RQ59Z1prD9TZgQ8fqWkTcOkurqjeoDHss83NLkZlqpendJeOKlDMYbblLBvq2bC
PY2VVuVQSeLiPfEsjjvynd4jdiLWpNrV2RZ0TEkSia+itii5o/zq6lPjRK2u3AjDTj04thNGoFld
K0FijGllEJexQgBLoJ2iDl/FOneM5DIwU17+ESGxFgrS/afSN4tHi0lSyoQJlDTdJnPBlR9Tkhbh
1Wdxu39cxj3VCuiPIiykeyAPF5xm22qBwnP5+OMHsICSWgFVspVnkWfZ9Qi8vIcV+Y/Kuz8Rpzbu
/2uHFEchYwZqQTk5otTz7ZqHJRdnlF49mZDHk6ctslEHLp2etYIA/Brpma7vePS3IU/5QrM1nlpu
DT5X09tMqSMk/u+BGkWWoHFdonIaQKcCmf1VZyvE2UC89nu/ei8XMzoyp2Z+PEOGbC0KPA8lRdEo
7QeScaxAcDsJcYb7RruZL4nchfnf6sh/lxZVyoiJhHQZQb+7cWgqLos6QcHf/F8dmy3/RcrC23ha
T70SYv4CWNt/WPNwh8PLdEXWfTGhDEyvtVZughjGyqO0ngFPogu6rp/exfmGoCEcxlCrQWeuBJW6
7zmbiisTHI7rjHtH/KREMLkck8X/EelGU1Fux08ezrNY7fTF6g2QVnvMsy5r0aidAvx2zxGdHKrg
yYcnPoyst1SpxL1+cWvZHHgxsU1LkqiVws5ON9Wx/GUj1Mcl6YJwCBEd2f77/uKqz6wsR6pBXXDH
vdYa0QLA9vuaqc58F1pUCHnVd2l9fl8EJkZoL9S43/TeSj6OQIr8wJNLiSaVLdS2k3WLcGOKdsWq
Sk/k0kq1jffYh3ICQPK0YJ1rbJvVimrNPoR1PPA1JpJ8sfI6X9bLZlWFuRhLoY+AvLmXYc6Sck5W
HOTFpt4uge7OFlYTwTsI2Lln19i/55vHmROnMXoorFS5KrjODoO8eG2ZzSRYeX5GJxxOWtVlC5T1
xXBp/OSjfYVlVOep3HIrma3/O8dYleH/PFlwDRNPTiGWx39auWX2RYzSXlJR0L9xsgFOpVUD+4+X
qBOhLYolvit88zegRFBaUghbNbfmpJefTOfH8cGhuf11UB9FGrLOUoJnA7Z88C7MBrGbNjeDU+o6
mMBjD4WXFcka+YOVzPefh3ne2HYCYJBuoxcTcrSJwVblf2k/sZR1qo5JEfUlfBMvAtMCpWnHZOmh
eInuHgg2ibMYE5CFLhQaEe4lm3gd1M9LQn9u03LxLXVHOGNcXIUj6DasFVsnNrUaJ2LzxQ1MmjD2
Hnv+NV5xKqJdkxdtaeN3KIox8vDz/yU6HvsuRJy7aso5B6poNo4kFUB8EqbfBVWp80Ro8y6yerE4
rjxgRzwPrJBgq6I7u5YSg72oqRTdAnTssZsXcD0hlbpfpm8u6BN46JsXokg4OZYW7y9HON47CSaH
ggjnXwLP3gzwOSoxQnGjSIzLv6q2oGKg1wzxKy7Up2Pdsu3cf0vLel77W4+A0XcP+znN6IVdOKMc
r16BVJKiuAjhElqWfXiFHZxazrq7MKvRBlN/lH/EjSP7i94aC/ey6Hd6oU0rBYvVfcMeIwUOln5D
C+kYJBKOjf2N+ejJmNcdGfyhXlecLjat6zQvGH+c/D/g19z10Z2NjlFGk7T6TqAucAfVQ/ju7jcE
M1WhXYy0ac/InGIpyoARDvGX3LWLAmX5+erPrYzpEeJ71Yc2h7xveFPlVmmC4j22W1xL25eUm2ay
7XpqCH4Un+2xfjFLuiCZtloqyV+aUshE+G/ovLcNkz9VT0nMmxUo6+A9YUVo9ktjte8qL+Pql8dp
Wn3Elkx2XwahWZxE5QE4K8rHKEFeN/61jRqEiEIK5VHKOg8CQdKzhXE3Altw9J39WofEUmzh6cFf
IZBx2M7PVIN8GiIWLaTr6QVCVhU1vGGq3afEGhyT7A7ZT/Gt0AeO895EXDISXir617aNP0Uges8K
a4CFerQu0CGiS73F9gWf4XcRMt2lCKxsVeEKCjjE66iGDqgJvvW4GaYCJCAyv2a46UJ8laHkF80v
hBWDvX7VZeXCmdyrV/wxuAkEKNOkSxwVgkrZSZS4JmOJ68durM33I+djy9zo7nzXJPYyDevuxg1H
RKt0E7VwOhKzm2JxPRc9AY67mOb1HO7Ujxl7Kk4gd1a96HrD4KgCfgGCQ/3LBYip57isnX7SipJn
uLIvM3J76ZbUvYCHDY1JIM/8G6He4y/xx7tCoTIjsqg5Bj+GHaQ0UJJhkRMhQC5yeU92NI9ny0aC
CF5wuE2/HKbQB5gh/n42cQM228d4ifEPBQ704gesLWkzJXv3+saMNJ/feJW0PfXTRfqYOUcK7N/Z
DUOLNsxAYlWH1dLTjvB23eNSHBfd5RKraHNRksedqOI1HOfvve35Mgbr8vbQRGbCvdnWW9zDmHnD
96R/xaE2kF5pxkzibNjI0AMPxAgcelHQn70vTN6DTtA6/xQeTLDXYNEHz1asgbUgo0W4PYTP2vDK
21WDIQA3XqhbSUOX1o+9gIWpO56HMofm+yNquFvPEckh18pPS5X3dap1ixL1rDNnj3BUMeIER2n2
ooJW0JiM9l6PAj7qS2azXHKvvuq6xNomgzfKKSLTuUT18kH0NJXqLFqqI10OKTPl6JL3I23/7imC
EICdZBz2EFR7vznZtZTidFVeWAp1rUBjTeJPAY0FIqa+QO8BaaQw3r9SQ0Bl2fwD6su1l8GxRqG3
lcg+cNx4IN6JYJOg8YITMBDaM3p+Oy5zfIixwepT1oGk46lmxdn5UImyIK2IJAKQhPIehNfE2stB
OhpktcPolQHoaQW/HCZVrTUyYHfWSBVajjMRE2ilpfPvKVQDmmrx01gRN3kcD9Xn3khFLP3Wn+AO
Ancmlm4OJ8pwvB2W3z6mIDRsQeEUN3Vj2CJ33A4HNu2yvF1yjBWXDKGLUxM2dBC+57tTKPO9LU+i
q7IvrORewmzPIrOm1rIzuspAnm4DULX0JEu6iMDXOWa4vhahsweVJwq+htAAQfa0aBTgoqYlIy6i
LAbQIuGL9LZvKEsCX4dFbzAjDI5bHyeCjRpuNMExn3AoyiiceOcTQ2lkucWrfIZ/3IPHlelHn6mz
dhY8EfBsGwfm1i3v3+mEo3o1qTGyhap2p/VDDcQpFoqgMcRJVnLSy+elDKJ4MM0nMza3qSi3mTbq
/ZAQhrtBSw5t6dRd0XsNdVZZL9Ce6x8rX/ayrTj0r/bnMc0x7fdM/AtHFgBcqUQ2+RiMVDst/Ttf
ALo8TfJtJw0c/5g2vqxThxkfXD7UgnaW7mwSQhYdNeJw6UMkHhkeLMN+lj/bqWjM2I8hrH6RdG0q
5Nc4zigPdTUvjatdUD6yGpTak0ZQHWDAl6z0RC24fy8JNNYKWBAHWNvKSq+uZcMPf5a99yKpl0hu
vzXDtOsDqSApkKj1NiCdj1XuY+3nE5FR4ZS3qHW/SbRj2MEw9mxOfdUJkXu3qMh6frhpM1msdWXB
LzgX9WQNwXdb/gM2BJzc0nY82yktHJ1CfhxRSt00/CQuTcsHbXsXBBraalNVaOdA1JKyZSUog//f
0XLjrDuLH27hz0jS+EqTMAXFikwqIPryf/PpiGge0ziZkO/6aSVOKlVIw1vJj/FpLHpTkoLQ/L2G
ulkFLevL4IOrblaA8OT0P9PTo+vScYRIMwpRrRShEobruQaPfNFy0Hh6WE9Xy1ZdFh44xQkzRC+K
GCWVzTyExU5T5llKEINn1DIryZX9t7PK/Su5lKSXVgw4zlwHNikB4eYPi8AIUTB51UYkXMfjfbBo
c1vx1g5NcqGNPOiKwUtpwUO5oOMCAY7kgR/P+z1pFLia9SfolNRHgyfpalz7lDYfGk3PaKrCnbTW
IE7b6AIn+9odf3FfYSBjGbvQTF/IpgeA70ifvm04BnEtdn6SE1ZabwwYzUBKnX2zxYHL5VsXLo/k
50tfGD9o/6/hS7wcDMygtKxg/fYEHGE1PtEDJ2xPvA/+eY09fQeghQ23vEIvVt/qpfZ8yYFrLUbO
mdp8F+d+pJ7MBlt01YsZtiP+7qruK35VheGLGKljBeyPYhpHxmco+3Gyww9ZHNrtX+4pJKa5lGwm
yBJZJ41pEKLWzQ8ur+VfQ5R8P3SdJGrcREic4GFy+EeBqjbLUm794Vw1j4P2P/uPb5plhJFPN39I
7xYQXD+6a0FjR8SmPs+4krJ6AbId0rvrfF5i6XAA/NozrAZBIvxD2pu7Z196MuNN+/UcCiOHA1wu
adECGKrTNSYKlseZWmuqSf6JQHBmgPeeVNFPPsSurtqjbQ745mAMFIoxVIFdv+/B1W0zP9nwypsv
+eY1lOhZPMXYUi/qjghXVodIqt2mmNDVs7Zz4/hfr8/3lw8smvuHZgHk3+2a5MjvH2vFaYhiGRo5
t1Z5c8MwCxgxHWglPZ8lmb9kM2DNKIMaAICRDaz0FeeggIN4ov3fiFMkqW26UMuAIzETjFxVHwZO
scTKbiz8tPo9uKb5HL5uPUlHMP+0rpyjisGSfDhdm5ogGtxPxAT6Va/1vZ/qoigXT7/MbaZT7ywi
YciDKsD27+OnpK8UIRIxeGEUzFFyx8CxCjG4k2LMS6bJYCbgveL0QDrBU0abQdp371muPm3PtzdG
tnpE8hOiKRb50KiCfQTRiHkm0R9GJn5AraOEki6idw1wbxTYoi5FDsMcukI2VoPKEpQSqL6U7jEq
5u+TtXjmLot4cTXuO7IkyUX33Dhyqe7Nlb5fhPbyQOwG39eWCQkO4tG979bW3aXk+hwaALXsQ3ZJ
3oDnD8O9WFTxLyzzApq3QYA1Lt5JUxJzziMfP3qFIFH2kIb7qKbRRHB7ZQHctME3Afoy0OJQHHOz
w1Q8K7dLfZtYmCevXV43396KKkrcfC0c8thr5TBTFYNsz6vGwRhK7ZCl67eCZylpypWiiHywVmFP
1US7KOuwim8uAqc4DWabfEPx5gyWW7nQOCSu/smqCJhDzRBGhWHY4JUvXtebz07hrGZvnzkOBgVf
ez/cOLjR170ncwK0ijfRb+nvB6rAyH/kR1O2rH1cGppHxdowTUm0N7kjp4Ir6hBv1UYl/rgGPmTQ
E5nHQQKyQaSH5vHS5LNMaG7TiTj2BGhAHPH551NpTYgRJUgPBerQuhtJimBWqaDUDlnFZEIvWF/+
DsHaTJj3AkT/MmaS3Cf+Uwtc4fSTtU67HpHzvakiX6f3OVXR4NOuf4TbLq8esQl6PnEBv+AjdyDE
Tmr2U0G9pP5Fji/ZjxcUhATMz+kRnFBQj8wXC4u8sPI1BhcxP1iTd2rYgRBh+g4bem6m0l21naWP
pumcNYkI/OmjQ07UAODKuASXgbuMFou9xEoB8qUd76mUMZ8jwb2+8UviXA5/ekUELDyWUA+VpT1v
3DYCQb0zUWcrO0i9SlbJGv6kcBEnRBFpIveST/FUsd13qcMe2nKtvzEU2VM0GzxY7ojcoJILsMWF
024y/XuuMoON3v8IpDmwrpa+1mxPmjS44cVSBOX/97LA7Kf/YtExB2L9Pfxrkp+91ptYcqolALcS
ruOsnZzRXoRY4csormd7ONtYLc4P1eEAa2DP0xyQBquz5cd/0M0l81mWG6qGf8uatpR1NRG7oCal
XawacNTMje1f1RFvHHmX/Nb48ShmMyQ5hgVHXIOnpR8aohN62AYWOsqPwn5JMhRaVjJ932UurZRP
VpzYLRq+EYVZPBAzh24sv9QV0BcxxRo0iM1c3zfVr9TddDGvJSaPh+ra+bs6tlJZ29GVsa/LAKa8
LqpGzlcqHQrp1A6OB91vAGLQa7IZBkcSLEKPIMaU1XgO9bHlDr8DaZS4a2N5NdM+tgLsWweyRySP
qjYJVYK0MAJ4bao/ELoEbl2RBMZI8K1S74/NwlTUd0i6+yLR2IaRQZA5rC4CkdTw7GbA/D3v7Ej6
fxWf2HHFZOfl2tzmrsZLir9PZmCDDWrbEhnF4FIzHSYyyRhP5mDfhMHpnt+ZPfaAuGQi3HlLOnK6
p4XdUXN8Ks8AKPtfwzwcFe+zpj2igPWrIfSSp+tVbKoRQtcUjz1WtKNNHoTI/0JyoboO1/zq2f/N
YUVUJq64oxxvYIrB4L1bMKAcOhXHiZIJI+3wdFXnst491NjrxSGezRH1OmmzrKYXhMb/cURidanz
3nm88cux4bYdculxIHwLq+nYPfqkC0sSFwlLGk9nqo3Wge47ZYNZkH/A3THgnj1b/OwxKghbekLm
1ZN+ZUcz516j+FsSAljVIeE+AlblOUP96OVc46TDc2aNsbkkZGv69PtY5SyENlfwLv32HXHTa8Y+
umuLRgH+BHNxVrg+i7lyhyNYVMB7dIL6+F7izYwRENCUrIyJzhBAKe5xQMxK0Ppb+ZJKBxEnIYyt
3vGbCIpBzkmzUtz8YlmkATrAYsq0FmUEcQ8kWkwMzwjeW89PLbO3iklUC5Ao9hE6FwT+I324JYxP
ob2CajNsRbyGQt5nWinmGNIDW95Si9hI67jXvCN2Vs+LodvL5wIVak1fSCGLxH1ZvwZ8+YaieRRw
B7Bx+vpqoWY3uOc1W0/0jPWjYzfcxlubCeCF/mcu3xIKgui9TWMwpRTX0hHiWHhyxIa2toRkST9B
X8TJq5U7yZAZiE4APV1j993v+MobVWS2k3NADHjY47Q/oCoyNxFP8MDeangknRmVKBb77DqHbZ5h
tu677Gz78zF1QD0b7jIIr5SUvD1xQiKTspWwTHc9KtIt4WMYAvxPep8ilvkdJHQNIuqpsfKeaBMQ
qKmuVS2innlKR0+8i9O1mm5k9V3EFTuP7579PcS0ptUUBKizS1Yo29TrTmown7J22KCTs316Wmhn
cebdA/VFaVxf14zZMsutUM9LcMzU0iOueIFl6OR0PT7WcNK8B+5HW/RXWzg1dq5nCbPU0scREL3s
uO42HFU9emBGmofD/CzapKqHfju3sdNRcPy+cr+BWEm+8OBvIyKbm1vddYOVUIvHt/ENltN4Np2N
bOASBkoZm6u96Su88ysgRFRQgV5ojmQKWNVrhcOsnXXCAxlVm90MPr8iV0r+KePlmovXhq4ybEM0
8ZE+2ZPkmmLL5Iu1n7MaxzXTNDWVbBS6X0HBq2ofszMBPBoer8acD2v3OB94JOEPdC4cJacwAx9s
e7IEWIHTq3UPmARryHwhHKepjkA+EK3NgqTZkzQAzLlZq9zOgDdjRG0Nym9iwsXUCNnPeuR1502v
2UQowh4LaEbzZDlC/Jia0ndB2i8ujrrAtQod2MsNWl3rvCZknASl+eUESL6lh/eboSIeizE1LWIT
XRzMRa1tJo3q9SYaQaLdMu9Vk1S919HlNl4P9H8TSjRSscWvvS86l7bDc9J+O3rGy9kjweX7JLed
N6tLms0c6gVL1wR7DkVWHW2NTlGM2Uz5TDVkCqNuMBPl3l6CF+OUC4Z9xqCW/w6UYrPt8RcujDjc
e0B6B79Xa5RrV0Zf6RD8+0NVJ+c5jOE7mynGdZOAXu8ps0tq6U2+QTAcGCPdJKgrYLX6YwfTuzms
UbE0gtiGCVAgWqV1OLKCva/nSVOCwCyNj6DQ/MK4nbCFboK4WBoGQdU+ASZ6vGpuqAmTa95PoRh0
Ebrc06u0rAhXl8XzG1877K6xWuA62C3M/Ab5pzYxYldYS81jBozSVwtQt7LnO7V5EJA3h+dExWm7
g2SnHb4C2SwPQ0US+lineedCT6+2sDtdNmOsw8HRe2TbHUZYVayTzKp6tt0lK0pA3gRiuAekyvMB
iYCOoF1WDEV2VUsRxsgfBQMGmbGtAvBcK6edRQfAiLfZR7uCdYgUk5/oRdWtwPu/CAzbjHRJ2Tmy
6M9FEMJ+lbk+NCR3U4WMfPoREwyRkguWve7D6An6xLMGRoNHygzQWKQg1dl18M61kJtbgQz3thdP
IZQRaw5+FL0NbhMGp7AyZISK6Z4RCiAITAXAdjGl8HdIB9FzmERv6XcLIKIhqWSQHS2rmY0eb/2X
aruo52Vgq2bbW6urAUZ8NpKv1bjrktiHKySScAJUhfSK9R9n4T+uwYQ6LBC5vWOjv2JZrjqZLWRS
YgVAP+Ccl89cNysJA2tTrPJF9uUSQ6Io2q+niadSTkDKHxWpVc4ojrW1c9tXRTfQc3aEYKl8vC9S
2/M/oxZEZr6gUTxVrOuxZzc7pbKCgLDNe74Pf/UuIOnckq1sEvde/1Db8qUaS53fZcFpATc0YpGu
4X1BMg0IBJWfUYc4XzcWSkOIL37BWSd8UMLpI8p3OYA7fbNQV6vMQ/oqY4HAtbohaTLMEHCWd2iw
sX5Vh22RuN1xYilnI/xhfAM92wSK0OGHb2K1C56VNvpoITaF8RDRzbxZmluyI7YVVKVbYYFPUQFq
ReHpB90kAJP1uGNffIEKzznYdH1nGwPveoupAFZ3u+iaqoqb/UV+7VwSJDBWFHe3lld3dVoUZwLE
Gp4B4Zs8JmUk/B7RHWfYajt13clJdbS5kLurZTtyP0CcxSr5nZX6953NQjeeagQok5lMFHx6OsTF
jx/jlg7HR/u5zuJFo602jP5DIx8mcs7wS5dDttgZtCdeOvlld1Oit0f/ETjp5JiqsV7J/gYAhfwI
yyJBqxR/EexWBnpOZnU6SEj4oi3YIavSEyDLiZTtEzA0OOMiYwIDQYGTuF3LLe8s5CjZqutAk27+
W55OL2Ltom+dSp628pX+wdJw70TUZLgJMdZziMKtwKAMplm+kxkRpawsT3lKFq2UnCdLqgmzQZo+
rvo/jleB+uN9zhTsnsimj1fnHEmsIefyhcKLRHg3o+hJvK53aJ4ii4SAc+7/MqkrLOfqdlrx16e+
Fa4zoS5JgdsTAsNCRKFzgST3+/mRI8c/19P16ppRXPeZM9yGU8z7T1U2o/vcg7Rm84FXWIJaZMtD
jsbhgVfKrSq5U2IWYX7RJoDioZz5Ugl/g6PQrFhS5m3tKZrLofZSwC6VQuo8HcsoimGrdbgIUCgW
Sdx9NYOj42Qq4sJFmziAg0L/wOL0tyED4+MbH1Z2zoH79CGuC9pzsdw19y9FZUnAb7zBTv0vFXkK
Vd6AXzZc2gCtvyizGpzwCsZqzRxxg6J2fLSd4bvlPCC0X9xP0CLcusrjxNsXnbxP40n9/nmuzT2H
nQkxYxLe6SQDjUqyj8deJJK+dLrITLme3lkLRSHyZFYctPawbRITuz8BuEhDveitEoIS/6KZiSlx
TnhUJb4TA4zragiE4j3O59yXnIz0l4gNZ0wPLtZWv8igDQ8Zm6w/tCSIg8Y8SC0d338N38QkZSgc
CaJSM7RY5cM6doYzrLke4X3I96vaS9ANYaDofhDSwvO07gwiIPmEFRGShBOJTQ6sZAQEY5oddB/x
32NMUY99fA4DMADekXHrimDYshMPB9DziZ9kAc0bi3Bu//xsk/DCjD1FbvCY1QnxYInZXKKbNgX1
Oh22kKSZormd0h1TlccPaZal+5KnzSfSBcBANx/72+Lu97vXFzVB2t1of2DEa8TclafwYRZJQ22j
k4tKUQoOYubaiVLbW3w9jyZeK4zJEVMeI/hmtIHtPOocY3UIy+eDi1O+d/Yz1ScySwGWEulOya8s
oBHkqHae9Z3o3T5UgQdEd+f/HKTLuGfNWZq1Hd+qS6iBGUMe6Qsu1A4deCWodDK8xVfUYX3pNsO1
KDtTJvJFKWNIdHzAwGKWdE8JtrnTyActvuqpXyHH/C2QFh1b0ETYEc6t5L0QAEfrdEXDABNIBMHk
EMWui4Irut+MFnV6Ldbn0PqGYzBYVh+CXwPuB3OmN73gHcH5CtsqajkDCcFd8XbGRW7EFgvD+lq7
+U2FQ0MiJNKcg/FxcBdeecbh0WOJcWCC0U9lpLbz2iTuaMFbNVVZjG75sHKJjyFMOddw4YAaOHUl
tm4HMRBZ8sAszG4sVpTrln6jgm32wPq8icXxwAsBL3GDojhIiYOnP/8VW46fcmkaxtuqGrXwLfnk
7wMTCDFCKXfizJE2HBBch9NkKisMpIRjvGyvfHIipnXpez9URdpFA0NhhDmtvS/ByZupmJ23sA2l
8oZ5NSi3UxGVZQkUi/bmZj7XScHeQbJfBpZU+c3OqyAaznRJp9DudlUstp554NAnXvDwDctR5w70
U7cU5qJpDj6ObnWnnt/MI1zDFnpep1EJ27UPvSL+WZ9ffwKW7svpY1LETErK6A5oYluFmKm97AqT
1WgInheFxA/emv5yuz1X3jX++LhgHDPRxkxnr/0GeKivzZ7GrMRcLGnwox4PGpNl2DWQuCnkvdT8
cu/gwXapZHnZ2OQmkjeeFsGwscSOTDDxq9DoslvVg04HvIMrIhLmQDBP32OHHkkQG9TGPi7W6y6g
x/kp/XF90zkYUYe9UDaPishI7KZHwusJHKtj2zE/68Y0F6KsjN2uDnudvVLgky7fFUC+MfyF+hOH
wo5aRf/TmZu83bHwFUgCDQZz7HrDf778S2NAkaBIy53lXBM4y6luwbmq4RlvVSbNL4eU/k9SOquJ
XbJb3lcdMdzLuytXg1/chTzEynisJz8F3Qrsb7nv5TfwgriOZ3NKpp2VZYVMgMNEREfYV8TtANk5
RBfsWJ9yWh/IocH8hnQxXb2usC+sbMsodHGVE5co/X6tg+s0WKfcSIemiEzrk0qTm/UFGxbWx3k1
ISAOq4v+1E1Lk/uWobM+0RqF2IpgazCA412y1gAY+Ny9ixEO84Q7DYtG8oPkAYPdT0OrznZQR8lD
1np/R9TVRgcEsn/zLNWf4q9pcVBhME3gBz9JjmUBE5CJmw6k2TE6r6t0kyVty50Z0fflA2NGOwXe
LHhstwoJ2x8pnr01AM/eBTei2qfShRYXdYTZPPOatdRjnWCn3NbwxMZDqM+5/OVziUepWn1GudAK
sp6lC8sPEBfWvVPbkOO8+HgOVED5tu1sIt5JA5yufvC9TXLH1DJjcxnpJo+PBu/M1u8s43Q9VYyu
lB33C3bGzkXor/aIFQEgp8k/EfQdSv5IG/kPkv4pNI45t0INlvt0q4/qb3f4YMDyg7NkdQ1OKUWQ
apbDgD3w5R6GQP1wvaXzU8VN2bIbrikpkdJSYpxG9zR87kJt/rDU4Va1/PMvuzGGsxhgTRohusb+
EoMtqZIbeHCjp/EhMx0wLJ9Vgm0uC2Ru3BOBOXCqgqIlU2Cm4+hq4+jvw3lbIwn7sRsx4X0BZ6pO
HhgW6ojHoP90rxahdQ2EBOhJwCQn7TqEcbffFIu1EChKaq8AhtbMvwiAvOdFPmk/Qw9OeztDwd2H
s5JcJhAHv4jfe0CGdhcDc+oR4Vzu6vOn30v99hNtSjiS6fIMitDgT0dTho2wrhIAP2ZWrKjxfF8F
j1h2DbLh6OEUN2iZRWtZI3wRTSo69PdguL3Iy9TSCcvucf1PNWaMalgfmQUHosGohn17h54kU2DB
Y+yYC27eeDK9IBhsX2mzgId1Bx8ahVl0iMT5vyFiSdxOg60orVD3U/KH/qJ/zgGUNPIwBv3AdIle
7TBoGs8F17UTZlTxV9/f0C7ELXHTajZwrUXlIQ+dQ4ejqLbGIVsDJhwVglxkVAFBLER+6Gj+TDX6
+UDhqlxMecDVCNp+Qmcx3F9BcZ8iywB3wmchgeTHy11RtZleDBB+SGI0WBVVrVHSj7sfxu93gJnh
hIUrOmaMmg8GMk0zeF+ZytrBTXzP+MB8uEkHh9Czvy6AwCfcday4aMnHP8lAc+zNrK4kCKRCo0Wf
YL9tG/PHz7ec078ib3OHtUawSm3GTFuQITbfAppqW37iycxvf67ToDaZIm1BEXZFzhrSQ3i3yXzn
vE6wYyjN6rnhdbtND11rCPXj0uist+4otJuLHLLMBP3CUpWOoJ4X2wbCjjalFPqTJ44nHKOzjz1E
t4nw+kA00jwV8B3iUTJb76baiGcBdZuXCtLffuHpQQ0EPHMAe3KTdFEZCpPQrPSkHwhqwYZ0ftZ2
QKO/gWep+7QPCsAcPfjrpsfuQ+kvK8nXEOXQQ4cs037aUFAXE+uqdsuUOx8HuCijuKUEtCmPNteg
r2S9lav1LXRy+qzth2hLFDmadVRQqa+pBskHMZLG4iZRkAZC+fSKF6LqRIdu7R6/8YjwSgv4cEJc
kVImAbp9fB41pQ/UOeuO0a6En5i1nQYG9eebH05/WpqOje/6mXFZaHp18dCjG+XY7ib5mq+OOzkE
9ZvlOG6yJuxdFofLbD4wdlKlJutN6zfnWUq2SDSl62fJlOXAG4e3NzunLs4li5d2s0kSlE1dRuN0
QKBfoKThzOFifng76jLaaiwGZjP0kTwwp+XIOilRsNGhpehEsC7WAwwDFt19fV7ra6bGnxeQ/J1J
Zl4oPDTYWlvXteEbPZcemkcygLT7CVOI/SJsPaOSig3iweWRC5UTijfMxiGR0SntaQ+EYwKJiMZ8
qEl5TxJZw1DXIy9YId9B6eIj2HawYGtxyJFGPB4haohHMeS7rMa/j8lq0dHE4UnwOMMy1g71dh9W
KIh2iiON6BK0CCHMKhIh6BI6Kfzz+fSU8Sl/13AL8GC6wJ9vyuaYsKS4WeaVjqjSnC0z4VyfFpmk
JexJvBXzdTE5ERw6Q1OiO5tm2fqOhJv0rBMgip+6J/zkbV4xCt7d1iEZERNZrZzRmEcbTcZXQup3
NjL+aH2LW1PXT7ToPNjnEu0iBwfV91X5PBkya/GwMt0g3NY0CBxZeKaZHS4D2Tmc0APpKTfQMlLm
xOHRTWnQ05SVSLClNdHsm3EQKSB33Xg1qyPh1+3aG+bs14qmkEt0GHu42xKiHOcaE83Jq3SEy/Mp
dfGIzLE4xKAq+2LGKc3oVciWSQi+fHlHpRV+7reNis6DcwFCE7u+Kpw1LGRTC8koJcmAh99SkYyy
x61I8KI4rguTqvC0JOzJrGJjvMT6n1Vdlr6O1fT6jWxw1heZAjOlTC4jb9eo3rck6COHEjxq2DsG
u/1DguP9n9YrriAiASPVjVEDvDvBUTQeAk/ipaRBLOOVi+Ag+zgx7vpeNyHaca6eqLkVC0NhAVYm
enTyZCC+FRPfqdhkD4pE8FUE2ZvH94sjso8aJ6C0aIKbUZp4nW8S9y6uiqGXo4MJaD7IvDI3PbVI
qypUmsm1n87g5mFMTm3ZrpQy3BIuiMJ8nvqoFEhtTk+1QZQ/dIMTtkauskRGJMpGN7qscJZxYyVV
/UirgRjkj7iSs3359Vb/gfPtFOBHoNZdeKib+85GanEbFCz9NzYASwUtx1ykTDLVyC3FcThbBTm6
rNy2Q+jsa9EtEMv5Lo6KWW2HnIwTl76t1XKIKKe9f5M7A1pRlaM+f8j64N1MkHsw63P9tCAtQk8s
Q3i6Sex+/cnTEZkjH1y6FmsWW7+h2r1yfn+V+3iwQ6nEOIztu2lH7DH8ekaZrhVtehseGMcL/9M+
A7dLrXDRIqblpSGxsKHq9pkxJrfKW1O81A7WEgJtPfBUJeRU1A18BmEXqFaA1sIVcgg7gIycVuB+
y3862ogQGCRpCC3QJPWtVGS1Ba8IccLQ3+3ZS+2jQoS8/kdcTiq34J8D//fXhXQkzdJ1vrVAfC9x
bel3dqUM5tPUicMFfgjycSeqyIM8e3EBQ78BQ/7CkQcJaSNaxIkXKM5DX0h5GCrjL7otJdL/q2dI
tqEWYWKJVK5O760lgnHi3YBcPBYoT48l6RLaf96YZoM4mJZrqI4vL2KQWDKw8qwfHc4i7qVLAeTE
PrGiafSDO3X8cLe5l7vaowhBaUK5HenbuEwI/J3U13qrsAWfvfrTQ7Awr3LiI2BT97KoscyyLLNS
5M4DLdOpt4bVWUr3Q4Y4H68PrNc8410TiL2F8mrA7iHWNcyUuBT1SY8Lq1Z/mvA41ljV2MCbQoDj
9V6OEBQFvBUIuv7qb2tJbGczhX+/dum7UesNgSnoGCoGKXkZX2msJvQVBx+W/DZ5jqTi2b1L3A3C
TZg7J+ECL6VEdKgpW7xQ0eML/6VHTlo+xoQwbCL3YAgko6WgE5Y3f6ncvkNMwrc3SBVa2L3m1sDv
j1yxj1DMqCIcolTYGzlSKT+7Lw8OGIjSHfwI9h3uEQb1CLHDTAdEo4roAi82FvJlzfuVrIAvsjlh
4OR3DzkMoq2pjOGk/jvggp98+trJ38iaxL8yvhzn4YXUWrEukytiwOydVY8DVrcO90n8dxx6EG8o
0jWzFaIrXHomyfKUJM6tSeIKLSQ1xECfdOhnBj3WqbrOaUX/XJEzEqKc0kUJDK1XzvBE2SptOBNU
2VLW30Eg0sdIL1TMOGWnurPv84PRqsRde+vjTDm5RAT32fpwEekTL9MMb0Rx6QyQF9NXiISCU7+q
Y/9pquqAvw/zBljW4nAhnWTLDWV7P9SIdkuto0EPq3v9Umy/6ncMnONePA7rwNMQ9R1HKRJy0a9P
WRIvZxoIv6LgtDDLAUGBHYDF/nMwlJqrk7FAPGlYWnloKgNq4Aui99YoD23P7KgfRc7NDwf/wo/L
9vJr4wNWu3eEox+ScLFagEXc/2dnFGzBkWHL30M0e/gN8xGpsIHvnTLVLh8w4pxr6oNKaXEQiKDr
SZxnwpKBiI6z+7yyaRazRTTTFuoPQzm6Rtg5B6mzsCYxFO8o3zIGKKDXQQ7sIhZelprKXlMSX1KL
GzTI1LQvCPNkvLmOxs1pFcqBIheRtbNTd7P/ULyJtwO+gOVHDR81VvsqCU0iD/Lv7qAb3zvuHoWa
SC+AJSUWVoe3gej9OstdGqrW2VlDDO/iVQtruqkl232OPGs2DVPNMQlM3nhK/GVsQCz65/w+s1Gb
Iui3i4LbBrZVJu5ncNPyq7RIDBw27thEQvrZXwrAmBOJGZIkbzoaoXApeCYK0rwUyADZ/DWWNiRT
huobBnKkqBy7I60wE+Bf8Pi5iST+SZd/lQdo4AJfZp0+UUVtXNM4kvJZ10bTy0mWu0SjkPczcJRF
1F0KTFg/mlmgEUEB8tSx5rHFiEylHJzQNZjtz27fg+jvvR09/rSjICLAk/fnNM22Nrq1U/rpBXzD
mxBM8hVRnJP1Qf1UUgDrq5B+Z0u8cTJvNGpVTFZWGeIL5Y59tIJumRpXEaAlfq3tbzlxcZbsP9gy
HZWMYU8On1HvWFvMCYXEhCghqYeWr+F+cEAfAjULdCECtTGTbHdqQAMierv+F8XN+1eJwwWCDFeh
XNrMBzQluEegH+7rH9jt82/6r+W8SDZKi69PypISqaxW4Cjg9sJ0oLx8uadcFOWEghcBHY9rhLCR
E7bXAgFLmuMHVT4rchhaOrH7bgGmlb87K0gQz6Odtm5d5BPK7wEmMaSrplzHZjoDca/9K3PDalJD
mx73maFtWzPuLIap5e/SJYFJDzpSPRNuaXpTvbFkAebbFEix7EJok5ZT7pVZSY+f/SZsiFPJytzb
mHLr5Ku6U0tv5Ig0ypSb+7oIwO4BzB6E0W9mUkKOVxrpyOEmJBW4Htyaxa3OhKMWV74DM6bgJZLQ
oKfytBOFprk46szuaH4cMe/FEYmHRAeiadYZ+CcliR7p4pWykbTftx3X9e3/RT5jj8nP5eMWTJ5m
kxJY3Kn+JH5o+6q5B4HlJ+zauRyeWPH6egR35SOCLTf/C7Mw5fGR88McN8SEBbcs8s5MyEUfZEUm
VXXISUeeRq2u1vAR/uZTQdZUFPBSAPdSj3hWiXRa4UL5GKL69XudN/CUD1AVWFhwtRA+u71+aCGb
pJ16dJphD2oZlefsHVFUpiYcUlcee4GNyuGQNuQ/yBSlAjV0H4/ycb1vFiGfIooHJ3S/52mRr26D
1VcK/uq16q4i6n4pTNnkOfrja/a5ab0oJ0bdg3aSNEJASGBoSYU26kAerFNiHtUyDiMBuWvfeyK4
5FRBJVbotOSM186VSUNaBWY01YLSKhHflSAT9xbk6vFF1Ts+pczHT5ANFEGek9q3h0CyMobaoSMC
HvDwEsR2Wuo2rQOVAJnLOA7Qy2up+WLK3jgRHKl0snHWhd4fWuNjQ0MNsbjWP45zdsLhBxA0vxRV
L/A/+CFPVhcHJcSGsrVYb8f61siSFweFTnYMv4A1mk3Nwlt7K8/XXHG4r237abzcnUDACs4GxYK2
fZrYWyNuItkurcNf/uoyamzGcNSLdPDOykhRCPUcSMm8KlyILlYL4gd+aP/vcmQ2tcxQ9jl43N5D
H17964qd3irhhRVSOe3VrnG3QiDt7wgIszoOLxv+FYnhNJzSLRg5IdCmb9oIgI2x5/r0rj1ZboT3
mGWT/4j4FygwsgjFBkg7Xm7GrgfiQ2rPE8jUq8sMfYuY/GK6AmzjO7gNYGElL4FrSv8hVMnqXDpj
1tro5wazDSdvFNKPqTZ+rbVD90nrXWDkEz4Wllnvlg/pqIAzOwOswx9MA47JJOraIeQMG5hTePNQ
vxX8CMDAg4Jt5PyfvHG0Q6uFksNhLSNKCpPc6peEJIghv6690+yZAosb4wd1OdIB53m287UFv5hE
sOQgJ9ZkrnxvIo4mwWNMx0Hoc8KatwoRegdF0PPT7jj0eNyoqN05S4H7WxT3ju6BRkq40vuJMCQ2
8YQ/tqjAhXHHwFIj+X+AkvHdyPSQcufKnfq1hSLsK47T8KHtL7nxsKdf8cbBcUYHOWptKXBmGJ48
APlNUxRjilk3ZRvHGe1TDNvTG0DQY3K9ogq8FIbfsG3GQM66U5wpjk9C59HZxNMKYrmBHA1DLv0V
AxdsjWWIk9JW3CiEEzOddO1lpLmTmX6bQEDsgJEtk8i8Sx2LIC+NMgg6FlH3RQ1J1uF98rbXOVG1
Z1wAGbPOi9guqRgVUH/JGb0F2h2fSuRTzR8WmPprQECKsR2mI1+SWdu8qJE0UZpJHEPdAD8qsYjV
3Cyn4aqxKoi1bkMwdkxgKQBqFvH1aTkBogWh+pUrqWKs90UHuw3au0SLmOprGjLIZzJbtTFX9k2A
FKbZU7IUrEcoy89ljuRWwzYR0fr1vn0+K2nXXCFMQcMOVq/BbF6tGejYP5bNYys86uQfZmUMEfUQ
ZQOUiCy6rHfMNAgPJwmMQlLetSrON0t//j1hbZwc17VPgPqxTNFcsJ8T7jc8PYnwlpE5SRmmngZH
wNtzmO8yoOPW9mx1UGGhfiGnHnZrjkcxdhXBT/+4oMW+zOIQOzE/gAO8JHk9E4lL9NN8M03sDKL9
ZQ1NdpCVCY9AZ6s1j/lp8YpskN45xHZ9oGhk/rY/vZS7EPH/vcJD4WEod+BlknWi6Z6qLPMUadiU
12fEM1gy1gS84vIwpCbdvgbSTDB8qgPZmroHfKcCE5xWetIDaol4dAi7bnspvl3Qi7+OMxxZGQft
Qb5HcdFqzj9+FEYjpg2Jg6d7kJKw0DTBaNv0jZsOuBiePjWW5rXH8pTFgweMt4v6g8tWsiods7MY
dMuusBK6GKbtTTWP4YzslUMq4olntFjHxCR6rQNEAGjlOGWaDel+N/S78xhoytgV07xgDHaxtbhR
cFVEmOu65916jBDNj6dPruy8E4V9k+MkDMYjmdhetUBKcYYvAHjm6rh2RTQfWrvLh2szrZWPi3A5
YgJVjzRLySqZ4crLP1xAuZ9NDdngVw2gqDSwnn4ad/QNGq/D6tKlZEUb5xKt4Y8GEfm5uivJs5Ut
SxzCVpRA6rIVvYyorpNPNYFsNLei8C0LAfjmGWWNY7n1okj9T72qP2OMAoG/0qbB4axwaIM+H918
svy7QjUtH/oj7PBde3n3EHGdIDID6xDIUkbzFHwLORl81FSD8pYSxU3YN9EsTVulLHCtVNQNDY7Q
oFaSd+dABTtuxfdvC0RvB9AAj3xJ74zRRfz/Wxo+kx/b25Sq2IiGftkOGVv0qjY5T9NzSShhE9Lm
ppF5PVtjxVT2+oH/xDPZF7Z/P7l4ak/wYaobwg5Vl1r++AIDomiiZhvQaLHG6peylaIVuD49nd7y
cI1iuf/bwpdwyJPhQrTLMKBn6SjBBETJ2Gxp8lcKiYtvRq+fU0RUXtcyEtPAnMhqQ0+z2aoJUS56
55qNZwI5B1I9u1eQRFlZgFxFhViCWtUL7S4EUNX8mHDBG4pg9bxvNvyLb7R7Nfe+FyAnzLd0GHow
uv0irIJlJXCFl94IhOFBpcSBiWhkjYeZMzfUBEIL3fCIid5BSzGm3GVaib/dkDLB7TYIsW7H9byZ
kp/zHbOb8u0cv8Br6UN9rEhHPpsJuzs5Ij0vGaBEXZ98iorMFFQrMsUyx4gsUW1boHd6/dfPiS/r
tFv3fQow7HQR/ZlSXQWEuIsOZ46kZe/j2erCtnHi80X9VpbuMJyKBe+4HPsCpBm2uaxojQ/hdCLs
og60FSD1Qs6C6GHUXikoBKAVOoE1QY/sPXqH5hkS5n7eonIMiMEm/2zKW3XsziLltKQ7NhKne8YS
V7RqpozGuXzxxW6K58NpWu64/MjLAyV4AlLWZ3Ytl4Sn69PRdC6IvPhbF0eCyfq9/+NIsEegh7Jw
eYBQ/VxV6ID4No7TO7tGLifrOXPFiW2KgRNE9MN8pBOH2/cLlKkCcmaqqQSLdG6vba4Mf2uXnNPw
V2R9e9KNr6LMNi4xRUPvM0+MR2r3SlCv8Jxdpdg8Mve73ftH+Lm+cf7pmkaD81lFZ3OTcdw5JrlU
rhHf1I1nu9frsKEMGNTJDAQq/2CaxWuK63KEICwQi1vyWeIsobPgeODIo+UF+CwZC2GdjmcA942i
iHrujiUIIqr/o/RaXEg1CUAFWjpbEgtDwN8VAz/0RX2xx3JwuCQSp3Lr5b+zsZ1v/rYnCWu8rKfW
aLFMLEPVPlZX1rYp+g9p0xTMGCIchn+SGMibu8CfOnPQAAWTw7CRYifbLDMRsSkG68b/IugPgYlr
CyYXRW3EREjAXuFTPEEFvmduj1O0GrjS6LRL9gA+lZ+SS17dMCegzcDx+5WRLQ8WZQ7k4CLe0bYR
M6doq4geUYSmsJbY4yknhhJLEMsCMmyGAekacKGzP4R3dE4axTItEcks8QVD1muGL+tONJJZoWLW
ZPHxfVEh5V0QjKU9Dewd0Nw06s5lqykl6jIF8IlL1Is7eeKyhtuHpkyUkwLSRo4dCc8hOxDgogzy
khvIFNvvjoR3MqQCGQzPb8OLhabjl0f6WP1IvolCJs7wNix2AMEjNLDM1oNiptTEdU5qx1PUMzzJ
bj0vW1MFrGgXMJKVFkXKohJMn4DOEScAc+O3Xh/NbrdiH8Q1rbHAP6rcWGFI7GXY4QAqw+AgGlH1
N7FiteXI3QHcOXy2t7uFKpqJskXv9UjCHlb7eH44B1McePUFHQmdycTzTRJu+Fk1LP+ufD7g9iM9
bizv/5r7htWQnl55u+A8rO+bNCkfFoQRGY+ggSDZpW5wVMxOU85BBw1hwOvr/N87qE1He3UHY+ab
udfQ2dIPrJ5Bb0mv1VegstgEIEJX6p/vzrxItJPwjeC/Ply79iOi/W/OLflZFBmuxjTQCTCA//DM
88/xysyauJgGR1wSS9Lir3D3/NiWW4ZfDER7O3lZK2bnzqOvQ5HRkI1ggfyd+4nprAHVGSk0N+P7
FuMOY01LF3En0JHlShU9Knyjl6iwRThT63WUo1bFAuYGe7oTdAEuhQe5opBcp4T1T0UYr9F+HS3d
hCYB7owrx5lESXGXsDsbEMrigc8zO7c79iHOzSHuNukbPzwW7l3YTuXhgRUXXrbkyjKEXmJUEeaB
8JO7AELFdGG/52S0ihIReJ5sWnGAMWnXY1gq5ycxgKeouqeX0tIDSf4JqTDgGhNTBZAIS0G6erzs
r05NLVPw3/8qg2Vjka40qj0O3YOX6NBShK6zCzGbOpoWU3q+CZx/JmJ13sEzYRSnSZO+5lujTdRP
gvfThA/lpqLSBuB5gPXkYVoESoaVkNVP0ePmHkRAa0iXPMht6MT1W+nhkyHR8c7G55sHdWToKwG5
ko9kkOENqWzhNgBLfEktcFrMArq0UfrB0UenhgHhFcgMutXuTw64mEARlVGaZaqJVL5BWXCM9FH2
04Tdo9ghx5pg3ILOXUxv38ctCoHYbVEDGPH4c/UhkY74zX4B//vrO9Ed1K321TW/jfii/sgVtzEL
bI+bxEjcm/w5KcVbtdeheQfy/BeqLnOtvbdudaR32RqCp4EAaImVqi9O9d+wceENMirZ3Oenh98F
ldGznXMm2VCXQNCJW+y449hyFBmDedj8qjmR0edWFkI+NXJcJRyeb6/uAmwfftBTw/Z82IUDNv1H
sC5Cmo7O/ctvN16iyWvRgaFz7se0JoKxQJce+ChHZznAcGB/IOx4F7dO1mcLEFEOwYk/qoGYUful
nt+TI10Ludk8hm6Z0Gnmz9ZFZAYmxhLwn84e4bb65fgKkkJoIVG2vft8F6fsMgrZJJJ4UIr9BVa4
ef3Zp0Dl8ZyX5VY4inaHc3jzieffk6vXpledP9kGKkUT8NVBvP6nfVh+aDrkpH3TQ+BC/qnBci4r
z0l9uwlDeK82PXmCtH4YZ+u9S2OT4OhOdQsyPTQUvrSOZYtBG+bhNJx4yhiUX4ZQx/7/LhGxrjke
OE6EhF/2FzS2t/wTvkuZot9C1h34y5GM2EVw8pe6SUBuTEHRt87U+M0wA+X1p3aQ4RTj3wGdZfsJ
hUcmC3Ng0s7jxEjwgYsE2NvqHEGRfHl781G8xggQOBYGhhlMi6tt+Yl+zYHXE32z+hCRb2DkHQFD
OlyAjn+MKvV+hlo9rkmsKwNcU3dkoql5Y3MP6af+mtLXUtQtZr/vDkTtc6z0k4g/bUupIZoJkTH8
IyDia1TvFGHL19/YhQyxelfbetvTv8IIkhddBJnxST2sGgQmcs7By5iGnQnIX5j3UL2jF2l02q7T
Bb4wZ9I7+Ppx0srWAj5c8WrILhA1YRoY3zp3NZSaUpe0siCPjpfFJTq/GBTbIrsz6R0L/k6QBXki
vieNL2KvFpmDz0p5jkp2JGBs7iqmwue/t2Pq0LPju2UpJXbrR1an8OIydEYgD0LXItKWuQ2pMtsu
p0CElubsWk4kQuurKl5UL9ToCiKWZRYAYTan1YNGeTfMcngO1CdskY5gnZcQQjkoh9S9pA2W0R/h
qIQuDaVeyKIPeFYydn7MQMlUf+41tnu/nokECoC/64PEfDb3BoetWnRnPcmGWka8PTkMxVs+X3m1
FuBQKHYmfIZ/VJb1CN4Wf/LK02jtfiyuzLtFrOwZp9k4NQOO7JTrBPZU6ynxJ3l2TcmLGg/cef1H
kO86xHUoF7VsKDX3zNcZBsvD2TLCGwl9gwAIikTPlI48vGblmxghz6Pl+E7tA9ccz6eUBvmTDbUu
MN8Ualr5G5Kz+CIawtqtiyIzCEcCVHOwR34t/7gYR4atO+U0TnjKFIIyBmxhO6w1oy2Pp/nGFWJ9
Vy/eFGChLGUNkDFXurQCnR+TFEH7qFe0yHqIagpvgicXZoTnpn3IyVftMFfWQ5b2s3iEIWbFp12z
StBx+TjV2CgSYkTmM861pEAJDdXmd32p7JrK9oVgfXKAkuPM1FXx5A5BaVUIRX1GuF4MbE08VF9W
PsOOnJIrFb3pxkE8IhU8rtDAUgVbEr0SAMX/mqOU3LoIgOEZYzfKrS9ZGILuL13bOIY/UFlTu+DJ
/04/ULeu2nI0gs5YHal/+iOmozKs+cbb87TEftoP/hXCOu/G54Dc5XILq1WNeb/hknQnPdjFtXFq
3C3oYJ2WQtq2UV+TM2f5kXppyjNgeoW0bT25F35cyXP/9tqJndvk6Pf02iNlfa3+065ZSR2Rn0VL
eJSS2pECtJpyQyPo8uiijtmOCbsFC5UIAZyCuWbbabuRydTFhgc7jCFIhYpRjhRpUAWWc2/vUJqn
fgsLIqPN80ozTk73aFw2/D4ag6d3AdFi2CiKddGxV/0G8kvLfxSadGH9K88kWG730rsKXxFrhhCO
auZIP2NnrACMe65QI6cca2ZLxHqoTQdaroKJwJUc2hyGUGwx9aAcqJCVHljz7nEvlwVYr1vbcdhn
fZAQ0FM9CKl68H6nVCWBUSQ8GdZ1t6uloUevTvHb8R66ZbH0GLYwZiAYaAHoCyY9AKyb6z1puPW/
mueqRRNAPLC/4mdaKzDm8TUZG09NIwsBgYBWNxG8qbJvdc2BFLAI03DrVjbtnoWCMsFkFu//GTnQ
BIzdcXyaI93+A0lC/7ACnFV2+jWcEjG8Bqa7a5yhFkJ+XMGJnxAoP2HDtPTi5nj613BaK47gVIGz
T/CHwDlr3JPW0ZFFcF4Qq2LbGAT2X0MojmMbwsrHzOfJNMqTH0XgJeF2lVT1Aqgw1bt3dYRK6wGd
mnA/IvKOZx+R1BvSo57NXLyZpUklhCdbS0kl3rtrlHiO3UIsxcxyIx4B3GLSQC8MPYxMGtVsr1U+
Kk3G7fe33g/OSz2MEYQ5aVtzKsLWPqG2oGJUHwYe/9uxQiGKs4m5MyLTSdNVJl/sJ/uKkEK+1yNM
RXZGsWWT5Nrc3icJAdP9iZCgVqn23QKfiPRmfLmR0HOD0SlJY1T/bNMwx6K17rLQEsa6RZqsX3Ks
aEg+EGSifCT0NUh5tFyYpaUz9iBdlkKIytyDMf1bWmbq1mkP4+1JdpfUVuWbgyj0x3EaD/Jpo5kt
DVnVHYcrN7ps+OZOpuBEsQ1dMVDAzxq0NlvTVg16ftYfvwRPgijYT/wUAoX3jVAJ4wAPN1bXjCTH
eKzTTaRqZrpGLeRAPDaAWw7Q/QTt5Mqr58h8dGUiQKsGiwn0E6g/D9KBhKwxUSXzjru0EYrwefDw
h1RFxI2LQXMNHrPp/mrOTQxbAICzD2rjCZr+kH+Fd+bWpxnt1I80A5LAUxcJlHVagtiA2isM4PBP
62ZQh70aQ6QCw/mBpXyXh1MD+d/UBzfMdM6W320gFdGh7Q4aPiGY5TbSbe5GVPKYmLU95olmFajv
T7NKwpOzELZFQ7Vnon7IvD+gfD2j59P1T3Emqen6J5tsanSZl6z2enAlstVKqd6LpISXFw4yrH4N
tmTJpLdGpOYHLbgtydDMs+7UwsjzJykBBD3YcoXq9DKJyBmWH/HH5iFgWor0Vh1qheRVtYxu6JFC
rW5Q92YaGdRIKLPT2Sxmqst8hFj2RutIPq9vFqqF9m+S1QtPsPUaPiDr85AQ2/RpM/akoXrX4ODE
zY1prtu+rqZhK5fbD8eQkIzvYiuQM59LTC65dtQDFtab5SYZEY9CLR8VWpXD0yzVSHtcKzXeOd3+
vWlkH5lOcJGSnjz3XHuj6GyauuGo/hTM8wXc+PbpOJsHY6Td2R4D8Dlr7zTfLSsWcVHGiai2RXAa
VXK7l9Z/Am2LkJdn4QuZW8oZRIhOZdeJQpQDX+wYx4h7fwsDgpTnjoDQ8CZWheVGQaCIjwrqDcyn
K/oDEpbDyIHjoOoQJGiue8+IOACrrpop9hE9JyhXx0a/4+W1IHrhrRQv2HfcQtvXSggYaaxu9k+p
Q1GaC83x4TUVB0tSw8OxmuCp4nN2+NmOjcPsXQWybWyTr4GOXQw9FfdwM4KPk+mOZ0gvNUlm7Yhq
9QK5GHJxlf5ztsDSATFax/TT4De/3EOky32ytkBnGgey6WbVZxjxAksHWKmeow8nGLfNsOuL/HmY
UD2yagJ9wQvnKo4oy/F5AXiOoXuxZvRAJyqwlAwcXTqftZDQmC7HqWHNBfWeCL/qDG2xRafgPbBw
4J3ikMxH2sFk9NeWYgu+21YnC8G93kZr5zMnFwJiRfetrafnD0GUPHwDxrgbq1Wg89YhCy4+zaK4
PEHcOsRRPAvebM31smlOwCoJW1/dEUGQ+ZvpSK42wkdfkF9YNlGqq31mUVLRId0B0o0p7B08cvc2
cm924N8C50gW3TxfjozFSVdKReFepXSuEPvn/LjJB7xBwKTYew/CDnuMsLS5Df/xSJKRoCG7zR1Z
s7UtgL7gz3F/I7lCS/pDHj1lKSvPOmYq5BlQNJ+w87x+XUMrhk6//0qqNGOY9l46H876Kcj0ycgU
Wym6h9ydXBgflR5NI5PJg8zC44a6DNB6gh5OmXet+9q7+VM1VUDBUBaoGc0nCO0geTs7Oaw+ujM/
VlBpPWpplzzbIFGaRyYHPH92eCbpZQa1IsPbwIlnbHQGUKw8ruYaY0CIfwgzDUO5ZRrKxxCzb7AY
LnVtmLHj7/eZE+CNR1ARgUpV7x5nLiiHwl3J7pVGZMDonvkO+mQsDNiZJt+KM/DA7r/CtZUC1Iio
gv+k5VSQZARSSkpL0HRmu/2r0iIVJQ0lUrmdJbVNqYlxc2gRm/Xg35uZob3DIRC8yrYbEHcjCbW3
kmTTIeSzetyfV9TI/DE6DAHxqzvftMqrPXDNZ5/qQvrNzFuZHBlH3+FAxDAQRmRaXHQglsR4tdno
eDMLLFvvYC4qDsNxgiyKOxWJeG9DUZanw8bcnef/DiqgXajuAVn5g6rihF/rWkOUc/2GK40+4Cnh
9+69+19jJRXWr8+NZuut510C+NL9p/GXgAVewRrpj/Q8VP1vm8QvSl9e5YvnrHuT7pltUZNRxgRu
h+RZQyi4Da2rjAlf5osGeQJbVZCJnpKHGdMZi4Vky8jbe/cYPeYOrRSL8wvHeSQiHGBMvbi6aiLv
AetBiiLICca3wfka7tud9Fl9V7hwJtAZCYZZQViLZhKWoahzCK8gnbKq/8K1VBMDaP5H7oRyHt90
QKLsvWWsXy03lFXE6TwrV6368vX6QCe7Qxp0lmc5KtyTKrFvvpnIAVfgKiiPcDefzlhGk0RY49iE
L2ctPywG58OKjftPHr4cGa3Xfk8O3rH8GnsAq4xCXGm9DKyzkj31lVAqT5gz0sup8QJIc+Fr0lsh
1H6tXxpvZW9RqfehFPtsgVVJQHf4seZLUHJ4UOVnb2QaOSMoHoMkOvwvNB85dRqWlW7HsO/z1yKk
u+6CPIAg3eSuvGwIUJbmseXlaKd08YSA4p+sUKU0M6MFBtGXo6nCpzQGno0gO4pUQCkqPhF7Btv4
LTz9AVwfElFHl6myd2c9f06qgNE85W/NCcpM625wgNqSi2mHsNmDcQbTs+SVSmcKJiEQ7y/UtBrS
NTlfyueWrjl35a69vy+eX6m4E5IFr7WWnyHk25CiQ+5bS7maXUeDbCy065SFP/NuR0OY9DpCMl1b
30IdDY36Y4Mo/VgL48DVgVDQw0DgaCSfpwfU9K3bV2/AIRvIkz0b2aCBpT+DzK+mgENVrFPrlXWJ
B5LRSRsf/g5f0633lCRkZWHvLM+liDB2YzQKF22axRQdlMT5qum+jFH84b34gw5dgoTkrMlkZaAq
XA5kq40gawNA4b+hl/ULEEJ59aObFl/ZjoiCfqlbP9EOcpHZhhKTOEQqQRiqoALfXrGikRk1VmFj
55mCG+CcfL1E8X2SFLD1xXfmyc/IFbaE7iXWsQjEls3nm7xf+38c39HHEWwHRBAHBNPztQ5rxkN7
o2EfekY6Dh3eQ54t8VZCoqCyqKvTxRgq7jjoYfkrsNtJDcPr2e5F/lODQgAMtFVkgMEVhclRTMsq
csGI2H0joOeMqVOcl3GEnIahJldUSptdmbs8QpIVCwBZFdkTyhnC5mLpMF6875y38rGyZ87IgmMg
x1ip2Sd8le+6MgUMabKQywLRLiEm4bgRTEdj22nGIHAJmb1ThZXh0HX4eyZ4jNMWiPdId3uwPZN7
gqD1l77CvA9HLKrQ2jCly+uwP554RWH8rswOQ6ZvE3+Kue6n4LOZGOWjSm/dV8FBPCc4/7AfJMOD
snK0u0RuAhqIjfrnFI2bwguTq50ENxB+tDp9W287s3Mo/5qsTgZ0xZ6CYBT6XmidbbrwKUN0iX7u
dSpnq6DtHFPw342aUTKbtYky2gBko5XnbsHIa+2QTbe647ZXdMwxCGBCb/wNlkPIcQXa5uXetPDF
4i0jMmWp2AksuDc7P37+jYMgFl6X2QNFhspsyl4NWXcFKAWG3nYXSQdQ0YF2FKuakAB9/pLJtvvE
YOambSkYFpz2J5lUejhwAMkktzj8gVmDjmOTG7Qvrn/KnxHuIHIbHDgR+TZgYezK1uEWkhjyuUWQ
dbgbx2r8viKLKIvKMvAvQqgouMYTbb1RgS9ZyrUvmgSg0kQvYOxiJT5Sf+7uinPEYbq8mUYtnCdl
fdo0L4ytqmi51nkLXwWqiNYpq/zbi59XrnqNHx07zBxBl/aKadRg6TDQSZtkcdamLsb/sdUBtuup
hDZAlMtitLzFr7mSFxDPialhEBh7gwyLtUBN1aZ5VZpiGfSgcXgo2i77+lzHT5T1PQ50pMQhmbon
7FMPZjRMvUypbUQYRJ8Z7tLvhhJ9b0milw/B7f1om774+8bKrKTpWgY/cbbVoHlR5VqV6lIW0Wj1
kvRaZNFyxYmEpiNOtYNnVDbGp9+Zd6PoMSdSCAc5zoz2k9QVKDy2if/Kh25mbAxfgCnkWKbNcWjL
oLwcDS3WtRbymQCbMSzyF5zIp8OQ0EONm5a9ZjOhXZZehirKHVIIt95+EK4qHTyVRoI5LOtSD7Wm
d77nR+7VRbAeUoVGKsRNUrZ0anmapmBBdJtPe1F9GXnGgCSOzyqhyaR6sTnmbkjqDCNmSgK4YN52
FbN7ZuBEOwTEvcDFiQ/iL7YWsz91FJiNfsaxFhRafRNr8JJURazW2nnVIerwI9BHt5BUsj7huvH7
+71LUWM/PKRHYdUSyQnSaV3vQ9jRWYyD4NoeoisSobPj1jt1f4iNmvITNB7HjgubVDfz8mRkhs18
NPUIuWHWIK44AKeBHMfoop+1xODjHnCduUtDuZydE4+IPPrn11c8xA5hzUk096zL83xJFDFjAkkv
OcNj4kcCDXt0gm44ErIAAeyeFkUu1tZJMH4t6VekztKwFK2L1q0HiynaQLAyc+fefA6KDYnnm3Em
mxGOfCOW7+oAKnup+w0fbVZA5GHhKwdXJaHyXU2TWISq/Q+nMpxbbe7vPICQiOzwB3rqNmARfLFZ
Y851KfKtthp9neMBrRi2x0WwfdbrUhVkjl+aQMD2CNjoTqPLhbu+IxkUEbX7DAMNEr4p5/FnWkyZ
N3gxdG2Ilrkp3bYTTa7KAxcMqc7B0OflzWhzJlqK3/aA/hu2XBAwLytVyjW3ARv4nkuChIlh+Ssx
RSvHIGLGWtYRY7hibBEuRO6TSZ0jy3f40lwM9diVIV9DHUYK1ls3Q2fVvNcrSNsggb/YsIci4Z4J
BoDf9zoEQgRR/5XurFjF0MXtD6OEt7QkX5dJ97AeYKda1Nxu9zbxDr/KKgUmzwyyskbIsOYu0X22
hfevfnLUrnb6T5HThUxCEf7ln9S+CoURGUTaJHOBpzCKrd4WF7ul/8AWm2fuLTCmX3dboTjAIbDW
bsKcoRd5GjVDlXUXFVjpdBK+iU9cmxpTcLBzuvGVqUX0ZuXKbNh1jtukxIQr85X0UB9GPqwIisAq
d5XovYhtT446+Uh+s+lI5Fk42sB5k+GzmakEoX7+hMEFV3OfN8QqPixwoz2lOAV6Df2BDcDPtQ+0
vQyU4QWdLrsgIIec0NVeWrxFcVJhFTWw4dlRCjjqMTxd/cqaC43KYNqCI8OAs70yyh71w9GIe6V7
pUep9fC0XpblK9mUWfcb4RHp5afjWU9fAAWxZOsPEEfKTiuTPOnBmaGnx6RpnchnWn04vLZfAkAM
ANxjbBM23HCISscJkdPdHebc4yrxItohBzk9noVVqutxXnBIfImYWwMWXYceIn5zTpB/n39bAUnb
vByZQWcZQQNWC4ih9aCybpw26LYOpMzNX6wt+3HFkfl9XFd2QAMo9KYXEbLLzp7EtNexIdpFA4X5
mIwwZw+azHcvLtRvG/zZuPf5TYs1hpdXhpT3mdANp81sUTzlTAqUcJ3d+ORP6zPcxOSJtZThWXVc
mz35TbSv5HmDNuWf2Y2kdnYDksgc9qoJ6Bu+2QZDkJk22uAFAalojPCXYjixplt2XveK//PFZ9nK
K8iEbQ7StiDlcJzV6HG5iF556oZI92ND2/Ouo/q0T0HYtzBy/CgGcNCt9hbzu1sc6tP3KvM+QbGu
LYcgy0FiBZbjvC0u1NXkRAIlZRTHrIWWnO/76voRxI7toI1LiTWN0Kf2Q1WgR16lKp1hqV5Wxl9b
/NJpUQgfija5BEgR4XHACM1EJqT/h0c3R6WQiFKi3ewlF5YKe7j0IfxrjtQ7WPdCunzog3IKkEjr
dABYYlmdJTRROdypp7/et1xmAcoWRBJRmUQZO0SSZ+9eAk9SnlDCuh03W28+N7zWF61TZuzf1Wk0
6sVeNIUED533bCFJcRf4igXG6UxcDTek9qQctM+aoCk3zwlRuIye6Q7wNvVVhmF3bCzLgk5ecy0v
Jxqs03skrGPbBwgzLjPH26aFg9sCXLc2d6AWA2GuwlfnMQgYEAbz9V/bZIEtOQIdIPj8Z30DdaWB
jQnHjIc0/cY2CQ6o5Umza86pHDV5xO3WnKh05pBsy1EDwxPK1A5r8Izm5ngFTH5s+w2xjyc/PrCV
ml6pUnMDH9xkhCqCKVRcjtlXGZ6rOq6Qr713NzHaoQAIG29VNOI60sM7QcbLiUI0Emh/rEIDJhbp
ppmk5xftG9z4/aog2MdQ4Ni2wiFHwZFgSueJ22Vv7hbO0sM3/Lwm2EXSplVez9tUmMUzOhw3Mwkw
OkiQtoGQld9Nnx0EIGQEFbCpr9A27NxCX2qEQlArJyS7ikLynEuoOvGMk4GASL1kwHCKDIF6tEFt
D6fBuaXPxGwdVUx0OkXrBVTc8R4RlnQFW/3cksm5TEJdkDQZDBo15oyPaFuEzVrcUaJ2FrH/Iwwe
EHrSdANPvZkJCb0VmgIozid8esC4SWGR15rUrGdWZ1uuvLhBs6EJd4d3+q/4kEU6N0yg3VoZg85D
qB7pU3TmyeMvFyouocAPqBtac1NNuLpgPZdt/qCDUtAC4ZtjuU2LhQxcnwXccsuwuKL/MOhBy1PW
/AO/ia9Wd6+AUCKHLxCe/NOJX6sahb0lew+M58TCmqFTiEvwpDGQsLD9ZD2UJ/YQQeDJVLY+RVWn
2QQWd24zv4g+yACZAsUW9nw1QaoCyq/ALVAAfI/bOsgv3zSn1iF6HOpF2IUTIUZuQjhAinR8D4TV
Ud9icE/1Qzgq+qeaUi9hKLL8NvTo6Ju9qOymVuDGufCy0jcPME+PM1QGqdeSg+OOdM0VNsi6w7ed
dscaPbRDGTpkjiS5FCWd1wcNlrFEqlkAy5BC7MIRFcamYj4hJLfGPPXF/SMTBbCfogEZ+RgjABBp
0NBczeTV19dpavcK1m/O1COSecmud+MtodG9TRNKOoUrMJhpFcS8Djg/FW+JCHNotxKOmMBd4W7S
ZXVACOu3DxpCfFuO5m8Hs9f8OfESxDn0UuMHVcH7FZ+5BnOQ5k1hkZk3BtSOVrDJmWtH2JEqn27M
sTQaLxFv/+yXceXXJRdmbp4jv0q8M3JNXEM7wIqxGMgaAgJQTROTnGKJHZqvpj4w1cgeWt9Ky7n2
8V/BJSa763uz62AzG6X6Lr0B54IiL6XimXmbbpi3R5dwZOgOQRcsYwwEtx081/szbBz3VF1mi/Ln
8ccUKoUyc6VsvG22xVxV4GDjobKTIeVShunHVOO0pKHvUAhew9YeBmQYEMhyvR3tLenUmDpDY+yU
k5V4HvvMTFPuY+/qyolqQFLTuTleZJef4ZHhcFXMPipxZEef5E1EKz/QuVbOZD9kUewXfKw5sY51
2JRGOLFVSqXDCN9HTfEG5zdji+MxwgNmgPrBdh5D+omgi8nAuGwphtp64Yts0FOU2rjsOwIBg13t
Iprsz9UPz7iS8ZREe5wjUM0a8NiVNLNpZ7gCwouHuRbOFaY0PYiomVll1Yuj65WkVMi9PW2/hvXe
ttLhyZUkL49t5qGvPJugKhLWiuQ+SPsZOcM+utIMN1pWa1qvd9F9lMjPltMXeTwwo2ZTMCFniMik
9w8BhSwI6u0o8ucQGHasKo1aYUC6rlvg0V/80jUjl6H2lArwqZIPzThdXM5Rtn5zCqFYdOJFMF7x
/zOfZqUyCOQSBEGx+bR5dy4eLKPPCphvGwFDdx31YVRRYjSAtdIW8zbQkVYkeUSgocKJJdY5KvwT
aNhRGt2l6RPDRs6girhq1V8i8qka4imDFBZoidCPBHEagBnIo0Qs/QnhQuytxxSt7IIWS3uEq56Q
q04uyuytb3YEzDS3miCeOofAwjNPDDAQ9siGFDmP9UqLwu5HUBvJSrBy0wmkLMf1mYSCF85/Y611
oifSDyVS2Vc3lyxwHP5AcKhwSXXkLqTcWjccVzKguj4EGe7MgiDAzo0bhdgZQ37Z0IDtPewVebDF
xD0hPHMjzzoA/fDgwjny7M5a/tNcUhxw80y03WyQYvlfbvSF6GTnkRr6VvWm9zO0s0wNOr4I54OB
TbXlbiVvu+699hsm5UN20JyoYB1SGUUEi3li/aYeKyj07P4dD+R+hIi0Kkm5QcdRMOEGIUW8IcaU
KuP1IrB4LHShDz7z6t+OLG+6K72nMvWWYy4qgNyWlHbZ4WBO1ne/96AlCrqIiVrb+uWsqlYFmzvk
IgTwNAkeF5YMcz1dScK2frQJ8V2WASb9A5/L7WRIkZIB5JMyL3dtPUSS3Is/zH0QQ5lYzdTsMuxr
SFv7WG0EyYrtZNi8J5/6IW1FtVxN/MFTKkJ5Gtujb4w1lcuRCu7+bZRHWuQvsVbWkg0y1KWpr9Q0
okaXJuD+H0WKJ0pemmLpsXMv76XpuzcQnFN66PR1eZ+Z8ewnD9XaK9heIpxzAq/9LwCFCaLvKkDi
7vlgiLca84CuD8LRrrNvyEKnpAn0W91sKg5aT8vj/zGy2zqIO9Gv7Hh3DkrDbegHsetAoZpCi6gE
O7M6CeUHAdIf0MzhkT7Bf9xodAB7cw9j5w/pFS8KAknrLoCksNsLLT9GmzEeM9vwJ7dluROXgqmP
VCVYmxJpll1+AagD3WrmHzdZUHu7oOfLJueaqlGNbNvE22vyKyVlx16ta3hNEva+AmP24WSdkjk8
fyauon7RqAaYjQf1M1ksBxC3ZPrpQEQ4qysHd3J9sf5MKfy2A+akB2uoBnjgjXqx2FJ6szaO0L5O
ffzTdaoRM3wd4qtCIyze3qReluPLjtm06dtL62He33gbz3O/GzCFhGMH9vK99mw2GtHHLhSk6SFu
p9/LNGgqoRcLAzZDCW8mEeEn5bSHeBPi4S0uk0u0KDiKOomy1ItbDckTiOnye/4kL1iGluLRDUB6
/uOJUp3Re/9ipPaelaBenZXb7+iwmH6yg/ajIHBXDxMZ4cklymRGP7IwxLy3X4h0FOcEDmyd9eIl
dbAf8q3FCB5DeYutYfgePgOrMVBCfH/Kol2kFkgzYpv8xXpN+vxymnLrE/rmsGmO4aX62ns05on+
y5Lv9jGw8p/ypaHTWnNjqVfJitQ5ZhxJSh6uIUWJmcSHUbCm5lFnSDgztdJ7xkWdvBRGxe2cdTTX
N8Se/cViNqrMatU3OTYfejyCIo12JYOL2HT40KzOjvfzzkDaigFzmTau+9dc3XI0YLI13+7MwOaZ
gUmBF3mnqy4QVhDQXpvgX0GVFy3Wxo6bdhFIW67oczlvTpkZSX9EOV32fZqZsmV+c+bWPauY0mNY
XiMBcCxBtwGpb4zw0x/fVOvAbJheYkjJIkgCo1cKq9fJUynBUGLxdlc7JGa1JL3VoaIRYHKiFCHR
D8aLzKLPlWCSEEtymls6/+7CixWA84xcPBBM7VPpKpCOq9bep2zpxC9cNRrv1NhrChygi4dc8ayY
eWg7Lz28JLN0R3Y20U5YyeoNzlAlPpeFWtH+xmAIuta8scHWkX0N4EHjeOLGDYoSECnzPGgpiaop
f7sk1PUPoPMpWvybz2mB5YqHgYOojRKvd7l2/AswuvseRnKEJNm9+72pKulc1mxYlBIkIAQImkFQ
N8lgGp6tKnetDtDig1mP/n+LDK3gS5d82yzhGzBHZjEu3b4e5+SMYtGH6CNNir/NKN+Xhb3gkznX
7/xL2qevfGzZxNKW6qgTGJ3FIyZv779T7gIJLe8xFhvb9/knTRzav5RNtqlEWorakeiEW1NkibbD
2F+/x+2ApD3KF68lVKaIrFOnKpKwX2IhefM03M55N7aPnGY+LQwpuGbsIN4Wu4xXnAal8Q4B7M1K
WkyOWM05h9jLlywFWyH15DAwMv4XsHm/tS/EzJe4oHXaAsI3RS93o8jHPG46xyeFoGEURerExLGM
FNPXAeM2JuvYO1Rmezpd/86nj7X9pRQJ3RGnC283jeCeKXVEoHoxfz9cXWL0m6t+KypYWHzeGHps
01YwZfa9HMRZZpMn/df7q1p8r02zT8BJJ40Y1fz96h279Z/qopN38EU+DjqSEV1RYb2mNz/Otqeq
x1m2WtGoQNSyLQPrWZx16a/M8Uu3uhG6mGcPxczhrsbeOkL8UJL4zNHrN3ovrg8cIx8pmhWBZzrB
dRscsKEUyCfnbv3aDrOjtawP8o8YDrr7yvGU3CsfvgeREktfgyXn/uLa+vXWFTOQAkFAlquBQcey
8AaGoXOyV7hvzMORRHPSxnvP5jm9LMlDmKDlTauimI4sK1bWevvNmNjLSl8z7A7dwlgATPB2/k96
dFOQ3NeTjpKgkvmqOnOqrpgZ4iSot8DdAs1RM764+I+VMadxeP9hVZ0Mk8ti7uPIX1hi7CQwjbdw
ALP065UBVeca+kJaoCPSgQ7vI8FiUPeI9pogNA/JU/E581e9/SoUc7xLeTiaGXF9xKWTzDPTpfqQ
FVzmz6d/oj1Yuw4GNxxJTBNmo5/9s+1/+URPgW6A3kNuadsgO19zLSUASSU8G0v/NitLpR4eHCjP
y9CQ9SeljBhH0F1fDGutRyQkh89wv0R3uFVeGViIsIXt0LBmhk0WBIbchphsCgcRtR6q6a4oEBdS
RKfoBcqR0ZyWAsJK2Bie1Ed5OY++HJFKIwlmQsER1qGVHDBWNFV6aQHc6u+i26zJgPTvgng6KaEH
RX2ww3XPlfM4SwQjqaRRzHRyux7ZnjX1Yct+UkAueXHMVjKpb2FyMtjLVdq+C75H0rEoM1DblEzB
URT0ELRQTmMvG5+KaCffY5oQKLLtLrVghNoayJgL/BxhQnMv3dF6jFME5FJ9sTt68Dqi+PVgQkvL
2jv9nul/bPRCHyISBvmne6hWQZ2XrShonXpKpv6o7lomh+eFei2IHy8EeMm34eKFDARxB8mhsNm5
HXxRNWJQM7UTDBtScgrBL+PwS88BQ9O+0+S69aPZ/YZiWv2ldWbaw9O493g2yFVjX4b/D2dXjU4t
fTzmIQQdX2azHfrbkDa24dy/0EMvsqz0MKpac23phJuLqLGnigaC0SPMd8O6By5eOksknACJeQf5
qj+kChltyVFkJs461f2GieED0nCP2HkH14gQ8FTVvOKypD/KqMlZXnunpJIJrzWINYnkrS2u133+
KaoGgnTX55MgO61KJETrZ1MiMbCg5+7qI6Sz7GhnluzxEeZFmSmDumQVxb1luwSddzxTAPaioMRa
jBklx/VUolwvMollq64pkPVcCVQVWU2s4xruwuFd+T2fkBQLj3IsH1rxsTN+jmOfZEeqAEzVUNBL
M2cDxUf2eL4b6rfmkl+bU2t/LwvNgHyzpG2zRSy3cCc/kRvKfr1NiMkgFjxqQfT++MO06lB6Ws1T
8Phhvn2uMo5Y7nXcqbQ/4s5adErx1DkdKWrG854A232TM0wMhZid4YW9THTNr9ZC8yxeL5rorEnY
xnNE5G7cPE+xbi1OEwae9rMaOGbK+wcddClPaNeq2vkZrETSNyyzDuvi7rIzf6UtEwvfFUuUc4bl
ZlDkRKVZHcd5GMxzbpCUNa9MfFPM4npOxH2i8D+6AqmgfUHC9/9dKxhRWstOT3pPvs4JFiW3VpZK
jbom9Qd8VlFx/jl+gbaCNPG9ETfqLzAv4lD7H0pvQ0seErV/MwxT20hKaAJBpkcJw4LAErZScml+
8iC/DQvJRdaLRlHDj6n+28rrfoUkBeSlCufd4z72xMwmq6QiBoxm59L0r6zK35GErD1rHe4fHnmH
7zwJcs3IrHJ5sxe/n0lMRoHXMwn0a/zvyfcOZ5d5fefeBbZ4585TJOyB/0MMYqL/OrLIwVakG4XR
Y/3wi66SI/5KT8Q6DSX9sMnrJTZezz9GSQNRFy4uSGeFoOS2c56xKcosJ7JADD0l3hGTxSbJDr4V
DvN4IlhYreI2az4Em3wiyNxHNNWqJvjEivnf0MxVLTjAStwyZaNXpSh0FyXNkRLR433GbSWHP7pE
hcFAR2+oiKkkaT3F+tl1OaSySKx/0YThL4q/kpKMm3MDOftf1qp/arLVUkGGHkI2MrpeFiBRInoY
dtjW44GQgAjtf5x7LU4A7GfmaM+Rw2uQbxDvXgkauK9Ny0QnPHUpnWVrbDjKjXna0GvXQhoExfMx
hNa5CVxB8yJG8xCi3O1BWiaf/hM+IiUQThlnHprJEFVmqYrTz3+vi3SQPgH2u0fpNNj6QNTZPkKA
iyjUI3ASRqaCUfnaB08dimJFoYvjPvrfbNhpPl1q/adlCh7jyyGCdJAKUAmtLFTIAeUYWkGgTl9M
qffhPmsJO+jy4YYvcB+i7UIa10XCGNTwkMBrV65lmcpZtJJ+18ions19DhXfjbY7SdrOt8dGzxue
Rjn+4+AsHLIMlVY1VsJQpybWkB8BC1Qb1kMvDcAkDMIFoVCDh8LaQx9nq3RS5praUS/Go5mUkw7e
lI9XfmNDrTqkk16Y4Xkf13dXBzvjJZv2fUCx0cUoCcc0DK2fXbclA53D/fifuCHsZeQ6u+jm2LFP
mOT8Bi0j95eg65+GCeTJWNLpeP6ObHvRFxKulNKPPf/lO0B1Ks6s0+f2zh0XwGlJR15NooL94DAU
KCfpTi9TpbqUsf55T/Vf5EDzjHNlJ6rg+a304cX4Yp1kodWDipH/ZjNppOD8V+YnTo9vaaz2YGkH
4hinRsAyZ97cRjMU80c4Ws99oK1n4pPXf7ajhQmxIClUNr2mTcZFLFZbOfoVcsAh+WbT4doQG2qW
fQMxJPjrcls6h4C0AOKv59OmoK1uE5EkPzRlQEUZQXKTmaYlNqx0An+wzkfQ374DREndHUfKXZKd
rtHi8ZzFSYqy0Vb8eSv6VtLACaknnM+wAO9dZ+g5iAvXJSfPxkSkF8dhPn34STFuM3k3DkmaO/yd
hzn2UU47GSmjxPm+jUdYXP8VRzI9vw333hrPVl9mN3gxV261STVX1UOzVlWIQj/8my8uRIp6LRdp
TEu2ibW+zOmrQHCy7BNE27SQ9gojViGQ16zqNRle8J+IgQ1HBmIfgWR71BZFonTBzIGVQZsos9Vb
qOsFit87/okvVRgKIpyX2QG5zQuj/gfhAA4UYdUvVOG13yw+WaJwpqccKuriTtro+n/fdXu3OGLi
gRJXVzU1jvFQsWY9XnwTiUakQL4yiL1kAYqtWJ8UIDYkRZjT41Z64G9IF0vbQXW/c9KN55vf0A6G
xQOwB76XVrFD+tzoOxVZydy99pHc5wqqzuw+SzjdUWHpA1ypr/VDF8S3ykuuEchIjV/umQu1G/P1
HJ7/a/i9qF0QSAm3gV/oKzHHbghZEaCrvVdVU6Q5paodkf9Yfll05MYl10ecKKuEapXuP7hj+vny
jXOteu+oJoalBWBggxLSmMecwT9Pgyaf9krR13m6YbIegmTntty8qSKYRIdWYxXsFFNsFPBS1GZH
CBkn6I4ezBBaDsW/u4JueLytGmgQxxWRWq4Kf62H4yvp6Ou3BvirPnmQKSrl275z2AQuWNwBduf8
wO8ypdzBGH7VDLmEf9CvV3J6ACe0KlwEkvh/aLQgZeokLfMGRaKw42LyT4qxcp4Q2ddxQw9GcONa
9+QzC/MVJRPCajV8TW2RW5k17nR/u5KORoMl78XJ114d0ndUFqa8NCEVK4D+GF1ZrsQ83DS+0Aag
xvW9LXpTRhWEDGCGIEN1Q+D6xmoJO0rhTHCh6hvcgOFzVeepsYmYyLGkCRhO6aEse+omAjquh6yg
lqeLZSFqi21krscjvlRZATcKC5lKqFtG7tVOIf0AZQDtJdX4dxACWdOQ+kZBxcf46WoWO9NuntSf
sAVmIn27jTTfLStwveC5MSOzweKO/kDjFTUDKxk8vePA0r378P1rYxqrhGT+jhlaxVidbOm7ODcN
n4/YzfwUYthlBKPgi0DVxgegVPOoW1pSXi7PHqqr2gPX1B0qgImdvgI4t7HW2QEcVqSwqYpeEeVU
clZR+50aXQ3iJTtUj8S3c4W+aJT6NBWXnW5Km0wH5gP8W4Azo1Xh8pMZB5JeWuecBbrbdPl+PZMl
ITIdRnQ6aQpsJ2gEK24WpIgoyOOEsPqRBnqtOv07wMJUYKV++zsb1IQExjU0hIv/k5XhZsZKnwbN
tgfGgAIUEM4F2RiVEejtK8Zqe3K3uWRmwH07pcFxTwYrRzPbS8D7HrsBiBKWFGGpxHE5f1r39Jkw
mJHoxYQewKTUWfu7BvRO4Q2CzWcu426Y7+7gajtHZxAZSmSKbv1FhOwfcFQC1YHDg88IdBUcmvQG
ip92CPzktXd5X4W+DSHtLcIkpWpNb50iIKuMunp5wqgvHNimsDS6HOFN93kpwVYRvULKLw+2XkbC
lqKrMSCA/E/touZe9qNo3OCKppGNpQi1xREij7Ult8ourkiZjnLHIbopJMqtUMiv/in7WfcqRaF4
gyX1dbRKkJnJ1YepYt8JOPJOde2I+hzKDoESfhNAo+jT9lri2Pg2gfDTnG8ld1q5F5wljSs761f+
QFgJEwvZwZ93gJkvpI+51+i/PBktD5JWuQwbs9XhHJJsl4rMHbxWgkqvQFGUKGVn5YqDSM6lLWqj
TKLGgoZ5FiAj4BetjYfixN9zFpQk79yELsNrqyUD01yjseI9It67cidutyvE8yb0qPqSZGVqRid9
o65fp/T+BQYSJv/X7QmwmaLo9tUsbi36gBfl5IhACl06qQ8wZEP/WX8PPm4DHe+99dkGY2gcJdT5
99+wILF4v8XgH48WTyF4RzLEFH6yx0RvQPtt2J15tJfspCJqlBK2tEWDdqPYQNV+DvPVpoRlDvTd
MRWpgQAclFnH6ZvlaA/D9zPB35tKWw9avzMk+XTcy64ojTWfYtk6DYLYuDrlz1j6t6Yc2XVzyCsy
4zEaHv1lc5FKuMFNAyiScF72hcSpCa3vsKI2rq9Ibri6DYw4cu94zLMNp/TO1pY4T7xPdpNoOcIE
Pt4kCwplfmv75ZksTWuIUK0ri0pCABlGyQhz9osMKSjDMRI+VgFznvWzlN6w241MuUc/wFlJ0FNH
Nwnex3UHvd95fIH8QwNafad07PmR3iZgiKlW34XSuesYUCrrsVfa62lcNF0NnYY2cJMHOuirLwQF
TF/bbrF03br+vMkbGr9xTvDuLjQEW/tDz8jslJbbIvRYBSi7ozercehkSJfU76S/UUVtGPrZ8LY5
oj8qrwIurHKri02ju3gt0NL4U6a9Wd/WZsPmtjmLceO6DetS7ac/LoZJEL4c3rkFnEDOd4eO3YCg
EW/0OualKMDZQOj/9C7ZPDNBaUdaGgvqKeI4Js+AsuV+Bhq6TaXB4NViwVq5f9x2GJqI3hkS2zxM
nbE/cgeWEmvS6zahOvTV+voBPhGDc2eM8+WVqeTPmhNCeHT01pcoftIO/7K3zd2kSq6DvslQngkZ
K4lA+KuzCPew8LPzoT0IlvcHbPGsPaocSHqGSi/SyzbIk0l0auufv+uMvm7YcWfGNjoGKdSLqzZ0
BGGJmzBuytmM2+oNOPofd9ec0GvD3pC407VHKY7FWhDfvTWnI4jKDMDo53mATGTuCRTRgy5Dvh8a
vYIdfJkkjLaUNmwXJBfZ4eofQ2Lf981wK8BiL3aI3yiUB8XdL9TGWQK7/kK5B+11rT2Nz1oFoN4E
6DIiDOA4jr3m4HZy8YWApR7LKu1OzNN0OVX0Gk7OZvYdbnI1JJbNE0zFYoTQrG27BSBL0VCaIZBe
Smxo+lalwIvMcis4Y+nlisbuDHTmMKBSEsF4Lm3LmD1KUBi4B8GCtluW2ZSNbGnkdd0qnHg2LCpC
T73gCv5J2188j+S9HqY9Ha7plfZOG7dy7fbQiahbWFV5QGzboqeP/J++DwmPun7pLgydUBBQ5D9y
tv1zIqCsNLHq0No7jSwzn5Ai8RwLBr7kQaZnggSL+l4OEK/1faXPce390om1c0GOiDsv7DdMph0d
0Ozch+ijHT+wm68ffHVQIoKj2nnZk21g3yUL6T0MIbMWHoo4ouwYsnMT7he6WEUkJozVAK/UwGJ3
Jx6MlmDA5XCZtzQu+9iOU3AO4MnQ//kX8/yd0MO1o5BSEksSnKTHZGDXNzZ0/RvEczTLp3RQfUyA
2QKBIK1NM9eamYJKKhJRc7DzFenkW3xsJiLrI033T6ljT134x2d5uip5JQ2DUGiZZGHR34BaLVFO
FM9+DwDK8LCN3MYFWmL3qUXPatWVOwXgmac6vGmYRByPziAHin9FL2oHPpG71Do76kHl1QjuaECl
aKcNd2jz5vlTyXNHtKwVfdRLaH9LXNQUJOvybrEVWkpyeoDg6fh9qNRiX14bjKym8YlkuaVRJpTl
xGEH7qAm6Bn456Vm4YNOTWSEo+PMZ6jLNXHKuD23RTL6s19oZ1YOmGEIkm7mVZZ7iNDmSFm0QNrR
eex60i5Zmm+JrGpu0tDszAXacRTyczjFsZDbNqY0WnP6HyPpJHDNhtxWsQEN7aNBu0YjKlfks8Am
t5b4HumRKCFFPaZMxBRZa9IcrCYTF9GO6WoBSVwBHuu4HNNOp3/ngpio12JTHzvfWvt7DrBFaQm0
hZ3Yj+0BGn+9eaXU+Q9IKt58UMal6boeztslGJCEObwgsz3DvRl2eM+tFezxqOEGUtptnj60MxiZ
xhZ7EmwiNOuj/tjqjESPEaL9EeTyDF6vQxYgXOCxZTAw8l44xg5EKFvEIdrCHjAMiQZQhC3dVOmZ
cuBjGMwI6FCQn/d85zDvUpaTJsgOuqYPKhwoXWp3U/NSkmVvFoLZtGd50+67eux4GQ/nbhgE5UTw
614TO6gylHp4HbLgaD0intXVPEzeuydDmNvkrUW3qJYaq2VZG6KrJuqNKbsbvVeAfeWOuUIW7R7j
Zls1gW6QodomfYcHwHTIogCFrEBx4U2HVpNlSoB/SLBk2Ok2/xIa/bx8QHrD+1JtrUuXOzhPVlVH
46HL1VLHTXIz31a5B4oplMs+4U+I3CKw0rfEtHdALOVfdTQGIbs/WspG1grgP4xktbCqb+PX+3Dl
Br9thA5vPNGTlrSVYt8tKGd/Suh3uaxvFVWiqqYzr+h3nl+jSi7fDsmP4sYofKzI9KRjlz1fTcbN
YS5lPujdhLrL8WoSkFPmT8XM9NJfT5waUTGv1gwlxrzMl1s97bDRssViV+mWshsWmPUnvZEiUosE
xhXoJtGgw5ABmkcnlQElsd0V9YZQRhKZhKRwJmWhMDYG08r08zlmGlHsHoG0NfIDxEYH2FqnqXTN
gkptejB/cSkh6/TvnF4sHx2VLNYgnuU/8/qDUMoSn2TMGjVRU5LjlS/leEz5d1u4ESDbPVUeoVn+
jRlRg6zBQ7jxhXW1cRAgu3HrCeJlgr8Svkn5q106Tg9Xr26SZI0LVLf/qkdCzTp+rTwAhO3euh7p
uGh7Hu4uZxm8Wp55LOgm9grHnNlrda+dKGyEJJwXBKJr7ju0xXO7LBWLGGy6Da293OkYuEjzqQ1Q
K0vc5p66kV0lZKxq+JdWL7XLEFJvRwaFgvzIMMpa4FCdpqDOhCSgnT4c+qW4aYr9eVesE0LKAcxy
l6w+gHsjOawBgfRZfik/tGAnK0ySkQMFyFPZZSxq4LYngylpzC8Ngdi4J6aTD4z8Q+fI1DZkc+/A
AZguivIIdPRTaXvEEb2gTCmpDHsSLxoGGy512Ok1uAVPn7y/FHg5QHFCLTc03OK5qd4L6IUluqcu
9xTz5wdKWHDCXtsFmOYEk4hE+zHJN8NJ5u5LPD6yswQMv4Gix7u8bgncJY3eUik6UTCbknMuFd7R
bqRin7k2epSh+aboRBNUVK/ySalLDYVuXYtkc8vpKzPAif4nif3DP9ZC/Br4XWooKfxbMZxYMIkl
JP7PvL7xxOMR+1e8LccFuvYsdC8yDnoZ+kYV6QbC6JRHVs7aUwH1g+NMW4oZjq4PqUKZ6IbXrFuT
JP3EcBl6YUI/AVwTv1J54jSI0wD1k/t35/S39zl37AYajOa5sDPK69/SsiCBORhLbTc1cbh3jZUp
yahVzlSj8NN+xqQy1GaaDwCzBc2tj5vmFPqBGLTw/7IIG+s8XAk1St6m3xFb7nlGAIZf6d91qQRV
SjLuH0PqcvIAzGcvaJdS2SkE4axSbh56nxZKv9d5kr84XmbvG2Hd+PvEeWypqn/9O8Ehxn+qJD1Q
ms3fYpjwMYbmTFGqTZNGbQpifjfboY+MF6FG+5om8KpdbvWAe4WJsDor4m9wAo0v/F9Eoh/IApvI
kffzcLNU2AGV+x31VgiM/GcmaGynpwuuTDtdPSBz4T55zDWn/r/RwII9j1Tw98H0AyLag/Xa0xlU
2hmJnSCpdVxBN9m4tjGPuJkllfjgYUI0a6Zr02lhjiOzTiaOw+/JL4LfRMJxjWjLi3syQ8ZiIlCA
oi99W1wvB0X52rytUz/eksl+aCAOBN+UM3ZqxQZF6B0q645hJ1K1ZrckX8Y4+8SAraKzCtIrPr6L
qTJFsfxwPKGKM5mqMPFpo0msJytcZ2Qd0DBCgdNZ+N3F4ILFlFdc6mEzcmu9dI/JrVaN6vD5qx4p
qVjCzdTSYKgGj92rWyaQFdbbeKjlI+cIrrLb4E8B1BLwKL8ue58OBQa09/V7+l3O9Vg+B4HYqllr
bDqioXa0Gq8vyl/DKFg0P3HBgBcfFACXojB14Kh0nXi0sQ87pEB1ltIclP0+h5ns8qQMJExcVCWc
J24R5PFKWgvI9fIwwMWtvGTwt3pf611gP2YzxVYV/sziYOfmcBBqt/GUh8q+nbmJcVx7GBBXOQZC
Kc+8/dTxPjMnMpvaR6h9J+Sm933jN7iG4Cqcg/TEjYxmGu6ZIwnm4/D5XypLbh/f7P6X12jKmHKl
S6A3m4HNmw39rzhRuGE5rOqph3H1Yn0YJVDD71E07Q8H5NjeHqrADO+ZOwrd+IJdTrujf4t3EYEa
A5YnF9NtPj34Rd4P9jnHijJHofwm6wEyxT+wuJSGh0IW+bPKdazcuqgFYFK7hl/Nfb7OLiHHugXd
Yh1xTRwB57gJ9rLDv40C1/gZ9991+R2rObXodmN43uuGhugAKQYjlpK+bpKKoLtaPtb3kGGasyp/
eAScq3yOnYPNDs786x4FiM2E0Stqf5BPLH389+NLZNwotNjDZOtdUvQ6f8lkPFub1gCbWvL+EPDx
Kg2zn/AXDQiFqB8JCtW08B4Wn2JQYgo9HXqYjmI8Nbjao/LbU3SSaWPir8pMCuzn8FGglE/gn2p/
/REh6xX7K9cCqnqtt/kIpj4Mgyq99OF+E/szuWvm3qa7ncvJCFC1xlvr7dOHv0CaUCHx99c8IhC4
q1+Gd59rOVsHBswpqbJ9OzQGadQXUmNP+WbGUcdWFycl4wKqF6qUNRe2Z7+77ddTO+CPRWZSZRra
a22AzxrIPq0hWK9tcwVTAn2c3w/r6eXr6NONZDy4XoxwQjSwBIclj5BCc/YeKrAPZjKoRXfZmoNr
/utU8HvD152TnRtdoIKjqUCXNwQh8z+hYRv57Lb0SQRa5iEt2V28OFo+FWUWouRYZQMB5YZOf5i1
RyyY92n/78urJYUyva0LWo3+xGzgebuHBjBXYIRVYOu5Dhob+GQN/mSor9arygdycmKGWh7ghls6
gCLaKq+zb7+vvYh+nJh72JajQ9AAa4Sw8UqNQfZySeqH86912lOyW1kbAoD1igrW877CfqMDiSVS
atNOw1RifZdiAIVrvaHTh9JnSiyWJwtM7IZHJI+pNtEs3RAShv1FwNMzJJKtH3YNbPnJcEuPS093
D5v6jDe11XnWSCMUZG95YTpqCzQp+5WK0VmmZYkuUXCUHlupy4Q6mFNMTzGFeCA+esYj7hiNoZKW
H7ugiSfcXFPXuZTZcuqVJFjWCFkWq46tuHoQelCWOLnGBcGpxB1+DmM7tRTP31eD5AMz7/FY1JiT
Hay5i93Eln/ekmEe+paPRlO7faMxRFPmZ6gZPoxrhbfKKPe6qfbJsNc/D3GPaIChY9xVu4iDnZq2
zrSLgcYR2txEdxumtEd7/6xZN6IwJ5hOn2Hpl8wLLZUgZO6GZGOKIjJhvwChhYgC9YEAX1C8lMnF
kUvNiHSc8mNFmW4eSEBkvJT6Irk7B264yICRFPxgBijwcn2Z1khhfqHAr/OgUytSVT5hK9Cdl6YU
bDIII+otP8fjUl0lyvr/4ra/wvsxJUxDBP358r596XX0EEWcgOSwJYp0uD9yw3DTnBMEA31WCOfh
d6gSeVpO1KVRt/mI3qtHkB703f2vHRLboQ/dHt7uqgcF1u7byGF0plyUE2lOrXweDwtxQPOdHH0N
cDDjrpgYSZGwDb3xUqvdFNL55tYvea0oDk6QUg3XHb5t/Mf4B2u/FUiO9ioDgu+AO5aZvjKTZfog
cJMYn+6wbIYEPJbpfST83LLJIL574RtoO6rrv5BCgvQGjCY2+NUorSqTlc+FUXl4Xz5DBQwsNltd
kS/48Qpy6zky2kqNalEXA1eOLr3msAWZa16Os5jRv969eG8cAvmisZ+eBa8IHNFAUZfh/RdxD2AL
iGX+tNVtFPZOSxPA93EObtfJkzbtj4340uE8umnoyML6R30uT9+gOay5bSo+A8Q5ylm5VdCrehrR
yw3SRNlOmSF9g9ptn+8/ZIJtRXKmRZqGh/E1E5Gfuj1Dme/DYHQ5+Xsx3Mo1wDMpC4cuDsotpuGl
dntcgnxHXSiJHMhAXYLMTzuZ+7/aA0aJU3JP3IoxTbCHAgfpVVgVnAGogT2WClokcFY9Q4SRFowK
HIXwsHA3nA9sKeqo4LiwA9IA3HMpXoNqSxwG6628X0MTJsJhWEvk8wupREXFTuGqKlPNbuVlMr2b
lO7Fc9HqvlEkXTAtvc6Ua7prsTuMCofEfZyzznL61k4pD8IF5aulbMLLhDwgalJta6pQ596RKLjH
ehGcaE+wWnBfsUxHa2IKljhwma+QsxqAlBBu7uO1clravkrV+vppR5ZlmexuuVKl5silHZIHVNa9
L1mBA0N8YTfx/sX99X2G341W3zyVBEFn/7J9B2W+fHvmpvNMd4hzvRyuDnqJVdEyUNAhRqocLThc
SXfiz7FIBAUqH3ynIio/nP1AmvPfySfKapLkD/Od+0dpDXm2COJN2yVNqmXHQ89RZ+Wl8/4R4vhM
EFwdj82uurOMnuOsl8ZV+Nw0QvtTaWc9BykSKB78WmbKrzotEgDYxLTfg1VksiDGKRmbYWZHOqoV
7hyaEaoKHL7R+x66CKkOoDtCztSoeUVftwsVK4gBnnlE3uSEe7JVyIaCWBb0Pyo+URRm+UFbCnQy
9n4t4cnu5bk9IQg+H7axQUjniovWjREicibh4+nz+jX6qNd2GipO0Pya3sJFJRs3eja/AQ39TTkO
4Ce4cPAxb0kIarE7Vi8v+yoAvM4KEGe/FVO8oSgsC14zcIwq7AMHScXm8FqUyNn0XvRFv1U4+DPo
bCeYybYFUS0q6/QTMmexcXcHhdUZ88EKiDNimQKjilaF35av+hZetnIeVTjxpxXTutQUGaf7VVtP
kktuXTq9BKQnHlQT0hFVxzFu1sPnBmE89Jjwb5/O8F7l+LZt1ygu/NmdlfZtAjD+gC7U82Yr1Lx4
qUDxxDR6w+uPX0aN4Ncn2J4LeqGSqtt9+GXZi9oDYiGJG90bJU66v8NJT0kASumF/eqipCwoA51+
GnAlLjOWUpWeRafEEnrUNB50jJ7fiThuYzMWAk4LXyDd9kFL136fRdm+vA55+e0v2GOCqVIWB/M0
xIHTBeIkOFQjIQBvJjQoTOllDkIm1O8IqIgc32hrH7OSsWiR2BbN0TxeT1WQ2s97pmAMagkw5Jsz
uqY1cSbQiYUXLNIT7N0zugrrRaxW1G+8wB1kBP3GDHpkl8uhMPQ+YJFmOlfGgng2ji9zBVmFwM9y
KAFUKxMTRDSi1veEqce2b1iPE+5WlJ44Mi7KqhXkHhPO2oAIfRHtJQFOyU8H6lqrNKVUCgXe2SNc
J8RodDNRVBMunCpuduUQ82xUxpMuEgnRFDcs9Y3BxecS03Hyx/PHbLNFK9l8qUHltenDQ5KErruZ
69JzuhANL7Bws7DFI2jceQ/9mJFSUt0vuAR7YIZZULYzH8RGqhzXnlsaIllEOBoGxWhXcUz7gRkY
naq5DaQn1qeMlfXQJUIl/Z/4ym/nBup7ZJnpA+/DHhrbpJIjgC1OQya4Hac3TifAt3p0EoEDbGRf
kVxMuZ6TZFUVTBbW40Axk/191IMyqkYsdG7UGqf6l/DoYHG3J3oCInuVM2CG432+lxNgBtb9RSHl
oJIvUD0YGowCugXtfS/Wk/VRyTA3NJ+G1nHg4D/rwF+L+6lnwku1Y/N3qcFacxAYOHzoV6bRQzdp
QUAB5GL5jXV0FKkY79yuBAW8fpOtRJSOnUIxhWsXuN5XlX08zQ4W3hXgSB15N0YQK8iFejE0fxHz
rxc1YUBYmnjbQ/ZykWDOCKiL47BebEkcSJbp1re0jAN6Tg7SYD+gI/9NbCnYuE/pHC/Qr0PeWvdY
vucMBeOFQ0UCMmAxM9NdOxTA+DJoyhFcrqOgcmQSaAXinq6/uNGFVAhGY/6P1C8Y13uqi3fiCZrA
s3prWzRZP8f0EIbz0A7NKikvo0F67uiy0ZCcl65Lp8eTzedzmQifPTT+lsk66396sPcTtN+h/74F
GvtsHTZD2htTDbFn8KeW1laf3Bej9g0Ep7uGMmsFkuYnVDxyrK6wD12JzqRir0rn70MUYixw3/ky
tM3q/tH+ZMlrM82KhSHEsxtdEeK49iDu7HT1PtUqJwwjMSAHI0QX7Sl32q8nUi6Wsq4KrWdxp4fY
7J1nNws+Uve4iYsnGmSWITRZ51gMGSS65WolhexVh5VqR0jlbP+DLPSltK9NmuSnzCs/QlBRSCTT
CjD7E/TC2q72kRbmMRnooEEAKrBq/zZWRbF7ZxUYDuzLn2rJvlfD21g+c5EY81JnT0WL44ULxTNS
QViPgTCy0JoeLdxJNSSPbieqd2UvmNcwfEcdO1Q1xygt4thVSeWXObFC3omCaO5xBvIrQdRuxJ06
o+74YRL7Z4CmHpK0hyDndyDYydhQyqxVOWqsC48Y421ReZNXxuh0uuj2wr5Sy18OqiMrJDiZIuVc
nIYtOVDTMDJEGn3Hf7Hb4SbELR10L+2skxNYaXAfG0whH/NHRF70GBQGfnWw6at+EfPkoVpuH92t
ENe1AVh1rZ/7hJ4tGALI49vjvooXbPmtU7AIiNv+Ql/4G2q0aXPRWEmPVyIO/DUIXyH/+pg125WV
BCyGmuKLZ25DSOVL7GNHRfvQSHgsS65PcEi3pfjKnt8/kcwjqgf3T1jw6YKwTQyaBPx2eKO4XDRQ
1ssGLl1uAtnOUwSG4ka5Shsd0tGEP4JfGuIz80CrQa1/5i3Zh/TYNj7GoTD5iPtGBoawWAGJXTNf
8NPBZwiurT+QHxAPpf6nA1GKJQtboIIcdZNks519FUQSyIQUlnUv13jNTnhClaZvSDsjzB6j94ZU
Lxyrk3GnnFrUbOG++DzHJ8i4xeZUgJ/R7Ll91QBY1ks2qjKpe9mFe+M3JyKu/nhXrNU/KRGJmW9G
EPhRg3OiCs+iLRQaUAg834I/uO+JmfE822hmkhbKHwuhZ1H3tsP3yFdD71/XKtY5+FZoCyOri9v6
I+69kYbJqi/hYDdGpMY4fyln8Nt5RBsgeLMc+qZg/ThuC6/5GotoPYnePO4LlPNqY4cxYOE0qL2q
fjAJr+yCZRZGwP6bSfdVSttoRqrN4EOZWbAmzaSeAhHG8jTAsHAz4pGCz7jGVc6i+HO6IzsQYCbT
1UNtmvvs3B+VaXBAac85Z7DKxKJOMN903PVN/Yaq0K9JQo2j7tFhZKKvd5dHgXEkWQUechRPmC7+
esKTyyBIKBgUIE3bkgF1VT5bm+tRUMFVvx3QRikTu3IlG7VXicqVada5KlR9wAwsOgRfEN+eMrST
sxnblri/RZQSGYOr0C35hx76XU8hNXiNKxR3G0OIhMNqVk1xRhQe6bML71tzm9gQWWhG9gsMICpK
SezrslrJMc1q8rgbJ82wo0TUpIFRq+eMdlERcNbgz2YjuYdJEQzHcj7p2nFmgWi7qMaxckn1MPEj
Xei1SdBdOCq9NkBTqNTqp5rs+d7nSGHQD0QV8H/IYgAZqP0qL8PB5fhHIQnuQos8cNz3DnnYSQSg
DIcrPgPscPXznkXWb2ya5w8eiCCoaY76+O/WmyLlrTitYRVismaJO1cMgdJbWXXMPaefZi0Q+VXQ
Yu8h4UDFTcOcbgMJ39fVJBmuzArwQ3QiIxC66/QIz0StMTDGRkl/mog6yDcY6d4kH7oJWBv8In3O
Vx7d6LZDM+jjwWR1lvmbHPYDZj0WPIH/0fyhvYP+JytBNviJveNhe2QmpC+DqQddOoNAV9cMz9Lw
wI1xXbNWfHbdNoE9/rEjHv+mzszLjskwWv+OyJzRt2bmBm61+5067dds8g5YrryfJKPK1OOGn8y+
aVIc34kRS6EVUAzmIDxw7GJ9WYf/KOr7EysU1hOHfavJ42oz26bMLqV6U8lAZ8ObDtdJKF1yqEZo
E8tXyW0NjXhFlyBGRg8gmuYFXtwB1+ntq6XemlM8nQQfAcyIQE6+ys+jCktaAil96AHdbA8PPT6R
1q9BYpro0OGFSkUU4OYStsIlouPmfuwFJtEAh2PZFLq5SewfjHQ86ClGQvDEs5krVLxqoLx/3V3q
kYL57mHjBUSMcs8u1rLzAVYUpvTx/bMVWRkykpBMz2UHv663TzPQbpRgkk6PXIVukDpz/n0aNmMr
UBzOEd2NIfPHxjksXEqbAy7jTTsTnN7MMcC5hP81lxIWiu9VvIWRHYo/4FRlWab+hb4CkQZD/miY
1IYGkP8CCUshUTTf9gcGH8sFFP2ZkjfeFSeSImFDoqFRVG2RVMglNvgvBHT21VX+6MBmfo04J4s9
TaxNZ+296wZz+2Qpp4lh7yUN0Ip1k6H9PiclHHIAyxVutxJupbycEZkO1yis9bKLQaxwE7ZVYxTL
GhVq2DPL/UVMjAi/vTtwq0jI9qQrMiQEsBwQ2gPlAhB1IUQK5LobjYXJ+ak/7PP4lOUZzegvbJkO
MrlN/cXSoe2vRRKeqoeiQ3vuz9+f4D8Om6wPd7Xthk6TVCfPSTnQKKG5lYd6wfM/HVPbuvQDH4Wp
ObSRm0IYyt/F97KgNMaidlVTTz3fqWCMYBSzGZsgN5kHmw/4hMjoLaV0gbgOlBlWLPf0EqdIPV3u
wFQdVcYCuX4rlSQu7Ka6HXr1RQQDX/PEtbaRlcXDFV3O2aZZsMiTrqAaUBP4uFHZJYkZLb8fKVZ0
BJmPirAT0g096Ka1NWHHiFc8MnHfbLVC+LUF4feZN+JbrhDaVvoYtUD8ulpWRr3dgHa7IHU7QluR
U/nmcrcrg7AiK1mgcqPiMMRWzMwW7tBk3zXwMZUelGCSNUEIlWxbXMP9ScXY/pCdVFohR0TpVyB4
UvKTMLTm+qWz85DxVlsDsTIjnPR24IuP2Uyx44chwBqfi9KnJ4cSa0GTyzBwHGCHgjceueJCa2h4
QEHbOEEf8oDaOavKUzhkgVSivDo0eMgMS71CadFCcWgrVGM+V71nKnUNir7w3fKwWfApMyqBkbB0
E7B+p2J3G5PzZGbfWOINr08qUecZ/aQVFVFJtqlmrgAcbU1d+yIappBMW2I9zmHmovg62Nm67oXV
u1vQcklvgIrDRWI15pqv0woxNKKt9aIKhlkdlqlNk49X8hnTG64sqDDOPvaud0J+xjwoDuWfxLdb
uKphY7eSA6htOhcp/MI6wWgwoGUk0JcqztVoeBwKpvtOoz9mlSLPs6Tsk/+EOoyyMsGAFAkD76dA
Wm3nVWhME13XEZ1b0m/J/eU/nvnLyWJm+6E6RqIutQo+rf9jeSToUGQZcMuHXo6fSGyZHRPUxLkW
2yZXrjZVT0TujA0KAXaPHJ+KQPv8KLCSG/1C7MIscqvaPXqgyeHP/KvHpm4VVT3xA31QhUU5K+8H
xhw67YxhUmVonrzjkYq8S4u3Comxguy+t3XCiL5i0iWh7YkQ4UHbwXFkmTKo9IHBjCW17uZd3MJk
tT2V3MtBYB/BoyoXtcYlVZSV9kvkJw0VpnHjtQ0PAasPareTwwy/oxe/m4CUjSFnp9bM6lsZhw3a
xTQTHD1nahe564rEcVdlCO30LGlzkFZdOAsVY4aeglQaTJJdT897M1g1kArNTQ/O+SrkAyOFCOwC
NsKUaB9r7EYVv24Q1HhJAIZ8lRkk75hjywCffjlrNiGLeLTPmpmWERf20NMtmArpsJCN8H4/va97
hO0fz9VPFE/Ybt9z2Bs9NIcAY4fs8d8Yoh50M21+h4LqP5vHHGdX4nlo3tZMdhIIi+SEE6SqZ4xY
A94daH3vzheu/AbLRJe3LlXOIwByVwj4OvVqxDC68mlFP7jb+hUXGC8vd56xI3m9LKbnXh3u3cCo
fA1YNjSTl89Atei/vnFg9/V44R3b72RsuWVlSBUEgDgMhapyjiqXUm3eYONw3A3eyhAnzvstATBc
7Gqj9jcFylotVWSWn2vTEJE1FrP7eCXMsVRlkT//2bk1J2vgQcAtHpXkZlPCON3vHF+TPMGHL1Ko
SF0Ww9C/+IuSuJxumsxu9GYtoBWvKVBh4FzmP251lrN6aoWP/92Q66jwesRpvXLgcVYTthYV9nab
KaXuqqDk7xHaWL2wsMGRevTWMBeEWR4/EUansLx23yrwsUcT3P03Bk0CP3qN5+6gK/h/XWKgaFkh
ksSSb5hd6fVIr64yr4x3owbgqWEmCIlLAoOLqi79DQqjPun1SrQRbyON2tHly1+Sh6ozM4YTCQ87
J87YsSijfoDs0ovV75Rm1bgaX9RnJNc6lCrKs6qHH6HsgeUHr8yq/8nT2VUbNZFlHy5Ye2/Q0o+I
BkbijJwvg+ipzDXHWYrLVIMRG/oS6egMYDDNU1FYLLnzDnZ3atX6meyR+KMkdhL1LKExyiBaJ7pQ
XKJUxnWTHV5+4jAfjTON0akQDoawDH8wNOs9wyXY+YuEnmu2zobxtgMUuz6Ujoxmtlo2e/S35aDb
pFGp1EMboJZNJhVpV3Asv2zQ3BGXpJGd88DuaGXcjvB6czSql0CEfYIOyOjNI5+hY3BUnDaJ44rJ
EDCiXmClAv3aKSj4CRwj7llFuFfmXsS6VJ15l+/Tgph2BybmNi5rBlaIlkbqatKTZvF8tCr2v2Bu
Q9EIjq1nvONdX0u+cYTpw5XNyq42cklF3grbW8yy2wIYAKawM0Hhk5/dVNVsEC1KgjUPcFc2tTkz
QgtmENmntJ5G8VpES7HyQivRYpG931b7xgYYF84D21D0thABNMRiMeIkBp1hRoFuDvfGNlkoAecd
heRyfIU59qByFThuxvyJohvLbfvo/dCuL0bU7omf4zZlMB8YqTM/si6x3sPrS9fChGixgF3Hgq4q
QzrXgNrYYtHPgga+HI6CZ9OKiVazivT7upVn4TbZ8iO/1+nGYJfPSPWpIvKTyfgRps5YzL8w7J0q
DRMEsQWStsFUKsZeNQlhqMfehqtC6J/5bi/cAXum0oDv3vga7L0PTyfpgWynDBCbS+X68SZDR+LK
5Ec4M9XhnCEd41vWdjTYnPoVuBZ9UIB3ESJgTYugX2cr4izA1cPUK9CmzvSn34UZ4/Ohf8itLXCS
b4g8wfggHdDD1BqB4TMVSTJU4rxCEri7nQLEu2YL7PA8K5ueDcNruS0B2yjRj6KZ8yqnij93Xhu/
6d1oCq27vm2ut2gkG7kxOWj2pkF3IlzRzzzPQRx5qUfQD4VMtt5bDdgc/O3r0mpA8Roe9J/IkYP9
kQat5rq9Z+IFrI/MVDXW1Yz+fK4UdKT7c9ZuX8PKt2CYB+assNUEBoJ+xuu2ujry5CDVXWT4nL2D
d/VeA+C7syRFFbixIEEUnUWikisiYZaxVpV0MV5MIchscAKyihEyS+wYKf6M7nhxXru1xjMZfDDo
7gYubL8Un5SmwiimocoFRVz69y+faRKFFfs0hYSx3Vyr9ilH7PXapGhBCXMDZj8rCiF19+fufSUZ
FdWD9yc+ZUydlTvW10ACQwa9F30LBUt3/7kmXH584bkYcVzGMG/EvHRMDPGZWPM+bjWsSFqVgUl5
Kxa0ZYdg7chvJXfFe+3FNmm42YS/Z+KlipCBsfjb4TxMXOUhi7TXJ8/2vqeHbIZC2rJWiSfFQ9Hh
sxyu3CHlLfYY/9nu95wRKc0//xGDdF4VRsYAg61UkK+V/Eo5AD9/6b9+Cb3qf/rDmad+u2gotWJU
wG28z57173gfw05/4JSbwHvf9CF9NHn4XlCGXuhRT0iGYkVCkIrzCcw2d+GDzNNk6nXnnBLQc7Al
nsCEjkl9YLf9luT3kO0Omz3rU3r2LrS43Av9Ic/RQ+gRA0KxRPBaZNjeuuAtOXZ+ftou+p3g0bJu
8hsLHbRtXpPlbGkx9eO1K1TnLcEva8C3SVSVyJM4MXw4IPJW2jq8yj0ceVKCBCN2q1OWyuFoHr/x
pYSDdyP0qcEjyo5lfUmwaog82eMZ/5Fp/lhmt4YIYYUG0jjYKGjunDAZ8I23m86EMFRRcTjZN89f
Q9IYJ9yHWdUmaeL2XnL1Zfkm/dE1rg5HMn5g8elJf1NqVoIeVHpvpkn7ehKtaEpgX97K37fEMM8O
JI8/Eku9vb1GHwM9TzQb+zsShnePT2aETQwGaZqnS22c9kY95JvU+GEnwO2WJ2Mw9PWV+BZBzsw8
ekyXAjOm7adTHj91ilwdZdAGs8J0u58dL1cjYby3WAHibfJcYQzN0kR+bi5KUhxVgVL/OBFp0/WX
YL7XbAod5kQmRLEBTP0F3Rqk3PqaczmI5x2DjNzKuwNB63/h5zxGNUpDn/4XKleTsZL/2H2yzV8w
ypI2skPGUkH7ngiGdDYMP64v9P7Ll2juGGenSnj7MVDlizj2TDPZsNWEhzX05B+tPv5juUQP7tXB
asD5u67T2ugRD/Kspp299gpGHN1F9vF1IKyBSFwilz2WIis7rVdMagrKnk+OkPrgiiJOBq777+8i
4u+VHwpe3/RJ6WLmYAIBN8FynMaMy+mjmwIo1tFrqB2sKHLXU3jMZakKhKqSCZ/H/3SryhLXi5Rg
LybMGCSNKwfOHNrTpXlJcfUks26m371wOHT4rdcSq9GncJIwY8KXmqHrm5zt1AsJBCwMgG1S7Md2
vwSvLaMa0YBgFlVbEbUE7m/SEqKVsNwGkrPrqxX7jXgTO9z00wJzZDFNxybcOkvdbAuMLaNwZyPk
xJBzWNN483PySVXuggCgy/+Xw0HmuhHMnCyafZU8m51Ur8dMJrsX4o8jHpO5OZyqQod2iZe5U/xO
53ozci96mOpBXaw4mZag6mzlQws3G9lRKYwGJvMQm/avlIslNWOlqxkWu2hKBVIWPKEzDtanc6Sr
qsew8rCeF6Pm+vcAAm9vYOZ5zPOB5MWZZR1Hj4G+t9xa4wtcJ5tmK7OOV6NQfPR3R8XGW70XH+Sb
Gvi0I+HYvyFJqNhMaoIRFjvoi/5Hyjkc0pmmmXSTkA8Kj3ArqfvHQTsgbdqANIMO2ypRF11hAjka
Cg17eSrN+5ISXpg6tNAO+Og3qRbCJHeFx+oMfxBC32WQjIPBm+c9FnA/66m0rJPlpMMlQK9AUay0
sb2d6CThhz2dA4V4HHiOr3UasZY31w2ebB22dQp4kT7XHGbmD7E7Z62hdFiEEz80gzRxbA2RjCs9
E6SKnCZPNn4iOAvoPLI6A/cvJxmfnbArNgTJftM/HAmLYRGavyrCnV612/54NwkQh0RHXDR+Cgt5
GYMIGWg4667a2oIy4rTkI9isjZ9wt1PjJ+S4gVbq7qbHRvX0x/dmu6zXVQWjyGIQDhjhla/VvjAd
wt1WNENPwZhCvKlgjSMkJNXvNZ4V0RZTYkjUUm6QwouvVZXCVfd3RxbccglqeuFxCllSQi97yBLW
GpW0S9tMbJ9bYdQ6AjVslM4hf1QelGrJmSHWM58BqUPm2jAxRQgkdIPqUf7x94U7Vyc5OlrFaqFJ
ALM5I0fUZKsxrG1oNp0maddmCluTxtSJ0bytvHtAXxkzznqwrWE0/j5QYBkcEgnw4cVio0n+d9AZ
cLCpgddFnIKCp69oRGuxeq/cjk52VBJ9+E+XsGNkBJu7+eN2W/KCxbJQTk3tkN5hstF1MRQhzGwE
teC/wA6cvthAWCWCdvjWTVITqtPGyxeQdnE6UBoJeLFQrp4gehRRGjtto69+VZaV3i7TWi8mIY6p
6n/TvyOHvnDzseqHOW5os5MN98VF/Ap9BBTCxKcktMafMsF6Kv5pQcKflW2ldO7+GI9AY0tBjaIf
uXru4KM5/w5yDqXT2nPgNULgIk5ozeyaduAQuFAcX35AtS0RIqUl2nFe50ilAch90izn2RYwi6vz
wMJTTjnmKVOrBRWPRTepk0A3pU2a+QzTaSji8fGiRTOo6VLjx2yN9nKUpKzdug0/e1R2TdcwlIzn
T7+V5zs8O1IjCRteq8i6v/mkvK0z9i2vdTtoQKb/rns7LoAP+eH5XKxiNeAHFzq0cng8zwcznngY
Dz9xmjblQzvsYtJbY6aJPEms+rZW0M2AlFJvAXQ8biMHnLUvamGKD/1ozIeZZyjInkWWUQ/zNvPL
8EafzSWjLvLDrs8Rt7wGHPDggEpDpyprAqdS+gfGRHDKwP+UqEqDsdFgSr8Cyfg5Qg7993oeHejc
Fxv5Im6eDEL5NRY9v3O2Ly/iBKOxHoXD/Nyo8Qw1rG6fwq0mPXM3Y1Jyn87vyO/iKF60+1IILJdf
OBKfeGUQUbfWpHD5+rDRnSVmYxbj1MvlIqxkFBjCYzYzBGH/LtDDZMe3RuwIUjFc08xCiywVmnpe
Urw5ryRcI5fsBChmH9ejkWT49AbiNzGbFYPqkW3qA2cauKWBoP83QljR7vphkpjtMgQISeomvn/s
rbLI4afl++rK6vy76U7/qKCUKHk88ilSuTyqF0G7ECEpV9Klbd1BXqalBe57NXXF2kLeyGxDvL3l
GNJv+SVbbqBz7MD1I+0WYqGjg9XWSLec5t7GknFZgqogsfhaoDAQJJnYeIQoIxWVPjl1XOJ/gX9n
7PeDiwbrsHAhbmPY6Km6NRkeMdzJSalnygVMG3GYT+UIcESs+dAONDUQ4VcMLdo7hsf+vlStA9n8
8Gq+vSue4qFXgW+r8cdab+Qi+NPTC+If5Ey9+m5kcdPWxEtG+PG1ZMmJW1nQ+FS27MDZuuwCMjTE
p7RC8I315Xjxvi9DZ50xVYn1GIalNjcTdRYUyjgoXuuezfXf/n3XSCGX3tEJpxnaqY6jpkJdqBXF
kwpgKhqDuXU6AGPv43EyHwK27117sTJ0Elp1G34hlGwyHh9FIgxSHSCBWEdzfkDO55Ayq/lEzX8y
+1a1Db3XgjWlPaIF6h8e3cnRTQ5Dbg5kLu10xZoe6RbAU6mS5AbfPNbXRWCjEHAanPlwOQWUO7Nf
JxyhXYuMRyB1iDayjhBtysSv8MIsdf2t8aty+d/zICf6BxBdcTrQ1T9YZFV23fP6yV3pzEHiPgXK
XRVhMrlOKalZ7+WHcCnE0MAI53mgcH24Dd7iym2uCrZTnmy45Vc5fbGcTNDkHycf2ZXi0N0BUlEc
Rg/mDBRZi6JIP/hEv6LXOog2in2/andsS5YvY/ZYiASUaULkuHysp1HfpinPe2IHA7Pj4Sj4+95V
vkHm/oPiXjFnRpg6ORb3/E9Od485ErrbinY/QWFawLldA2QwjsejDDWEhVoaHLDtDGGKMQGqS3LC
U2bgmAE5fmppTeEm4cT+IxDVlduEGejr74F1PbMI9YQE5TR6qXkJXS6mRkKtrB0hQhgdebfk8/Mn
3v1KwlXSXQ06GPick7bLwMXvygXulGfMckeAFV3yZUxDtTFh78IGIUh0NfhcnBMKkfJp4MUxUucJ
hlbbgZN98Rr54HT6jGppUq89uifpHrHn/finj8HuxQuVo0ApVPiUsl+Qkv6JOcXNGoqnGIuXWCO3
SMAgs3Arbp5BD4le31dwxA2yOpomTZjCW0AZEogjj4eZjc2dsTB2xSn5P1WG1TSE37gPxGqKKYdf
dqvJyg2M3l1G5tUpv24aYJu64fbqDbkEiu3C2q4MJsMlyt2hQOGEojB9NlMQx9ZO46GkwRSlh74M
n+LObnimchkMblQUDhPq2rEGgNiIbcvLmFJ9p5oARsPQGNJqj/4Q+wvQARHCf6A7OeWdV+3k+Wcp
sg44ZAllfTMG1MTg9NEuNZFXXDrhZeL5qtWEFI2N1HvSjYIuwG0n5qDkDg+3tkOXwUkP+bosYnX4
+cgOQnjREM1CltnfonYTLkYs99NOy1yotzxToW8wQcjym8sJqefAe1W6rKK/eAnaL5sZ6ZWt4dUf
fipXJk8c69EW6FK76heZZEKCKLNDYYAWndJztK/VYYffRScv2GNnWaRJG0fXrmo6NVqtG52eCRZ4
67vAihnIAm4iutgD45KzZJGQnJxzFVRYur8Hy4mb4xAq+FAkrxe/vrpBVad6aMKauZeyRzQvHqvd
txfzp3THR/PPc3dzsZdg/Zna+fe3esDc6mpO/oM6AqC4R2vR5W2tMl7rZJNwBtx9TpIYdE3QIz7r
57W0GJAw2qqnntWAqKzviRghfxSRF49rgmhR9/KlJ4/JcERhRYsIxp1PasxtXZxvrNIPs6LmSYln
Z3rWDZ7zSGLUB79wupWX96HJp+OECtxMhuUUisiIQfgU5irAmMQeuJKgohVTY1tIdb7yZEsz9Mbv
6fEsBA0v1qDq7tU1RiGzmhk4uwMuc5fdb4b66fQ/M+kCWqb3NTaatSHBTjZfJxb7/1cbfo8ubo9y
oMNzZXP3UHSX75C0QxbIoIf2aYxLvfw3heHlX9U5fcrhT7g8vbuEOnpzIF69OqmR2/VzLWdAuH43
pvvSUt9nFFk/T0BiE8LRWmEZcTvE2ZsbD3eElhrz0ZBeGcagZN+3Z9Xfv2aDoueLHWLwVJj3giPX
4qmwOnKoTvpMPQAnXWEg5loFU95MEdMhyaauJP4ix5tTG6SEUvpM+CT4Svg+UPQtnlOgP18Wyg4N
IitCsQvanpSH094ywM7/S0CiJsPv2S3f4l86KvSzpjzsIsIOauvhinHhY8JTNl4l3B7YYjxKs9RZ
p0TDAeyz1kHVRsxRbUdoFIJ4jaIjOOyjZdIKs1847ft7f7afG9W7Cpxnd9qze3oLj7bf/Y47OE1M
I27Bz4tZGBRj5OY+C0lU22EIT5FhlWT+Fb0RvTuydc6M6+TmuXa5UAk8ow043kkX1aD7fsm/AIXD
od5jhkwrwl7PMrqegTNr7EyatYxOZr0+vK7SOhs1F6JS59mdkCSoW82/9pKZzVORsq42nRw5R5/+
FudpcQZ5o+SQxW5A0lsQEMjao4ts/ay7mEeLPEWXlcuEtaDqmXbAJpnbmESHaTGoeH+cpG32/wUC
nnSH8hMRWRI4vwM3u+4FNv021kmxnIBwkNPbqNEDHWurPgPm9omHWIHVq/URJnb/OCzV4vS5I9Wa
QfICavWDr2Umb9OHAHAfRmvpNfAas/+6n2B+N3+h79DwH9iOrhUd1AvRSEjXCfI5FYYYCHOcKd4g
i4HakURodGr8vuT7IxYyId3YyCow+0SfhUIlNAPzUKSP3mSnx4+slu6dYaSPueuieWrOm7XERvRB
KAyVyjVuuJ93JyM0GXyoryJXPpdg1uWCkQuRbzgisUyhVkSmHsKEjr4y6miuHeOe/W4HtYwKCTNn
kqIp79UVGuHC1hFMKJXy4BMdd+8FvAetRbj391gxTeEupcfcn+o7AzuvJ24A9z5p5AQ5c8symK+X
qlnu4NEvjb2vmrozbK3m8MhgbOyid9ySezJ/obpFLwyOgSe/cw4S2pdi+YL0oLf/4a9lrNwlvaO+
uf3dH54DVNEZQFOg0E6f+WNDvEKLdc7DwL0RN7a2LeuLHx3Pd4UCauQimFBE0DQPCUww7OZHlLPP
GhF6sfpNP0MS2J5HtCrGJYLLlIGWU+a+lghXB7fEtuHJX7SxuOdex5LfsBc8Hnyxo+2HiOmB+XZt
sUaR4uSqkPczGEOafLaqmZ+uCj2IOPS8KvzMQiLAUYcML5NRms/1CKPbTItAJCtOz28FECxndBFT
xDqFejcR4cz1Hrcso0lZpWE8U2N+3Wp+eYUBpcoLQTOAy0QouBlmFUFGtCAOtGkJd4px5UcV0/9o
waLnnnlLTk5mOkMhEp9xCt2fAjiAuEwIiCtaXeA/7XV46f3KilKaKNarW/wdLi06/gHvaqbWzODK
r1Cqwi8D3lznso4jjUX6QdydND7n011T7NU9i3A29Z3w+kf+jy4o5Sj8q6VOxadRKY9X2iXQkJPf
ZQIxJE4lSGdaedro03YO54zpK+y0AeUnILG/VnO9nPue1FtyxKKxSG7P8GzOLbhJ6ShZMU6QxsEw
b3W0Uld6v+uxFsS9pCUfXYcA1sWSpagx17cxiSm+7/+JA6oTDthnLwt4H5W9DjcYaUHQSVYHzq/e
Na0sk2tG0abaUGad8N0OqEmlqmkCyRtll/DOrtv8ysj0MXdB9sixrtQJ8jPuw7En/Homx73RLjDX
ojS6OOQCFu/Bzz5tiQjAnX7pPOPXxPbxIrObooYel9GZKld9QOhmexgSr5n3JLGXGw5r1EHFBZJ7
pqcdbYJMvj01vpx5GKb1ycsQAXCR50fsY0uJdjE2gG29zN/vW7/Pju9A0W7c7Nqp9p1d3ugu60VK
mDFzWy8xMKuXL0MhyofqDEArBBu23k7vogX6KsnA9k1SwBSy76Y86JL70e+x87ARIAHf/v9pRXkF
PrBRlWSXFnUjcElPSbTUSZqN3CXA+o04GALyS+n+Gkn3vNDSN2V/0Kg1rkb8PRFYaxyrGqwVEJdD
W+kx+qt3X5eO5h/0ohweX3YycMTnTh5yea+LaTmNFVIw8Q6vzwSOOQEYb5NRNFCnLQdgZaQR68Tp
oVF7053FNebUHvF1u8QjzwhTQlfGz337Xg2TFSotIq76OdTRkEXPd3ZukhT0Ld7IX/QbvPyWPiGJ
enEKUstYBQ+MLY2aRsyOO051SXNQwVvwwI/qETs4XTCrIvZXcXFIRPHBWhvlm97hAXT3FfJCO+EC
wJiQ2GeW5vWgFLKGFYvMVE/8ygAtBh+MA5TqzEX1B9azvLglMyrqsvskpAvb7O7YTPCvp553RBdP
1huBdb693wExT4EJw2bFbwpiL+1OguNFMIY7SMKV/OjlHUR5DnvdV2WZnXxfmSQzzBII46dGPYpw
fq+E/N6rzw5hBtZP4wPytH3YYTPPxalihNbRCsi3EQgxa9A+o8IEQdL3OgjL82AWpcJiXF67aOrA
nsjz2Bm+ziG2eDkkDFKQsArr8gDhnpd4RSiFsypXvMBq+fchbyNPD5scCIs9YY1Vykvy73p8bsiG
NDzwZ6Xmbr8tMQSh33AQISiuSiK+MK1ehxVYRbt9KH4sl+i7bK3Z8QSEZZ2ajzg/MY+CnU5gFKg3
4VGwtPVI+1zCLBkI+ZL1UUAsDaPFLKlzIO6RnLan7ihE1l/HGlb4hp+8SJ+h6dBLTK0HC/kmtEfk
IOOGB7lEsKd5ZzlcfQ/ysejvZy62aNteXvC5N+gjFmA7RoWDQllfMWTTt6+zmf5BprxRv5pdeujG
q1W2JR858vmVRs38LtcWIUTKUvnFUcUOwP2KJJawntESEucT6Hazvps8bGKE6Cnu3IdMMoQ99lwC
0JD58pQolU2v3Boq6Cg4qef0qE2v0k4jnHeqN4/wq1T4au4ILir6MRXLr67BFPSZ0tx0cBgIp3TO
yHKllUiaegoHpsrgN0HCNbHCK2KqmUdlK8xcjlN7rWco32abEyp8L87gy3mYGFN808mhg53o0GO6
/X20EFrt65Q/oOPUZbk2d4sb/+51zvPPH8BsTyM8oF4yGp9+i4eHls0HmFoaWeyhbYHmp8v7ZFiK
YU8uENPZ4yOubvr+OI/WYPYPIJ3/L7XkHiv5kH72Pai5amxnnp+0bkt2LSRlId6/p3Qi8TYY+7/q
O/xvw3njJhbekeYQ61CFDJh09gmvzdgXt6PngD9yCEZGnXqD2UpHgKG3Av5IKQd2qWAwWK8Mi/nN
n/Ew5ESTcP23EJ576v+5TK1+4HCBBsN6eaZljV/v9QxHCqgPYuRcAtopvPz0GeIUDEo8QxrVoHel
0GeBpWVgfjJLiH1VLV3TUF2XBxP3fIqvhaWZ7meYBPIzWFzyUpwjMFz+WL4C1rPacKSMrsU5rUeH
9A2u9RjzKOA2c/A8gjr/VEbvUfB+6KEL4LPcAQv7+GaE/6Dl2iR8khK+TR7WNirGC5L2ChFTjCCj
7M28rG9Qu/cKt+0ZtM0TwjijRxaovoEFru0pDNyzBXBAl85E+G2INJQFeWy05gdCuraRyWirw4lh
BhwPEqYfh5ssZyK1myqHsoTKDsuePEwb/mvVnX+vbH6nDiPqHZvOlmBRjdDUhgL19wZG1K3einRO
6hBOvp3T9jeCipWFLSg7osOBoB6T0A+4VhnWYy35kLowNbQXsKdDjQM4gsVlkElOFpUL/+k9tbnU
/hALWgSz5Jt7rB3PREUF09qJOK58oTzqZj+xi+FCorxSyEcch5stGcUzFHBFoZPvo4w0rL88OcMr
rYMeCcha7PCM/oYHwQo0zu0wqCXNNwnRvXkDeTYylq72LD52l4zAkp+3G8RXz8NNUbSSysaMx8+K
GDbTefGSIyPnVkyQEvCHTVjhMQ9+kK0zCPrQyh099Yj82qEixPiOwVSid0FbyWr2B6da5BGOYoBG
Z1Ar9B2cL+Jze5dB0zVqubNHcsUXErhYC1qCRv2Lf9Ksl5nFmqVSonvAFCkDva53+znDhcqbwCaY
TuTQngkk1wc0Mmvlk3WC+mIQ0l8212wPyrOR5voSdkZbZLAhlm9lA/31r0Ilx0mYeHR9+qqUprqf
cwdjn9jhAIEw+P8aObN2fbB26iskyXRURRdFMfhwZXQqMr0ITTvleGTnf3tSXYqfTwUINCn4m9b0
yCxE9S9ZmMWEQJKzbR3roO4xdaSbqk7dnDKNnjKT3ZkYGmFoKFqUng1zS3IqMfKB0m91etDz8zUu
TG0BZHlJg/lclUjBjmFAaFobKxRejJ8jRh3GjnPJFoXV14+ecE80gzQJJgvTbs5RzqoaaABoeL/N
+XKoSv//xbCuP6QBspBhPQqLXQOV8JjBi33fERpvY0+F/P5OmRrq+9A5P7PTqaDuxWRJZ6wAWatz
qP9exVK7wEpcX440qR86YGpxhZ2OL/X0Iom1ZRJF++UHcRq0JnOMNZhfSW5vMOVm00wOjX8t5gpw
8LM0/a80qHbo12co04wPahcn5PiHms+Ykx9kaX4HemkFD1QNoPHi99lEo/T1FAokJykkDS7a65L+
xleKJ0umHJEuFOLEtGemwSf/ieDXbe8bXHj/6AioLHkm1thJPoK4sK1FD0AGgg68tj0Dc4eKZvN7
66tUI26mDQelkN55hShm9mVotYydbyfp43ZqC6fuJ2F89Wp++Z30M29LdbWIs/FWF7DigoicsPKj
UKgiXAS8jc90lPmprPppvrdkg0FWXNbVjKg1s4fgn5cYIGT0VSINPmyEwDfwYdvqA/jwampXUO7C
YKi9W8R2NxA/y3+fjfqNpDz8QTEPi82UXXsIaL6rYoc6rTHjv9j3tGQOedXDqNl7E9ISwUloSD2q
tTVsMSwMLmKSLHXK4lSADkqsLbsO0stSlDnLl7KHRUSnzU0rp7HyHOlN/SsNPTuqsrYHURtez+uK
F5b22eBeDLmPxyZwEXBtFzZFYcx6JIL+QTIvS2kRMyDLo4+V5u9HN3NPVQdDVvGe84rClP2vesxB
v+OKnCOCPkS56+LWWD/o7yOYSa8W8Wl3TBwkqW2jQ3vx6LUZ1lf0RzTeA/nsOGgFEcLUZhIQdVHj
u460DmbvYJEosWjMrDbUOgGy4GfPxqy19vYEILoKu1fgQIyaNkQGdzvFOSoVMNaycGHJC0a2n5Dp
aMXuLswNkHwwo/yZkaa1Y1HXPH0jLgsgEtQN6dqm5m9D0tAuQMRnjZi/aAlE0Jhyx87AK/cNdMKu
zZGPIB3uf7BRVd4WNKX/DuIkHdQYinH9Uct6EawhE1W4HksNKgF0rW4Y6LTb5JGGYiIRJtsFMilQ
P+fTlNDenKGdPt7uSCAlykqKulj1nL63008pi8aZRjdH60uVflGIS3+nrpRJ/o+XFZWlJQjvTZgb
Yw5TXL9aDneuh9Ff/GMqgtNCtHbsoRs9AgS3wyoJ+6xUw4dO+TrJIJxkgSLaCabu1lZdJVaMoDja
aY3te0O+GsbvGn/ZenFLca/7/Hru+LQNhQ0rba7Gu4CczmpLzJVKsEA9OxQRhHgskTC5fO4M8z5U
0W3YtMtaCN1ZM/qj2IrV4gQvBTiyZerZK/qhyuseQ3RRXWBuRU6N+ZtO5ysDkUPXRhBViAKe9s2p
y53a6PCwparWlU59bkQxfXAwEV4ySU0F8b7P+pSkD/Wfi3P+iTwvk5kLFO0ckhqS4eZQTzB7mRVz
c7wprv4i8grHmZ6AnAUsQpjxViSN0XoyxHYm0LC/L6jZEM/+RAaLtEk1Nxr7dBm6d3DE2UUPIAbl
XJ32zhEIpZIuPEZEhflYB06P63L1fwDwpzdDeO3ghCbIRNCGTuomVe0iWCxqlrZh0NYOg9bpET4Z
an97q0LofUnmQ/DFL5JwAv41fsLTsqsqBk2z8pjGiN3fHPt+6xBDKLiZ7r6rKw+vPaONH6Rr+YJV
mqUtrXOn41cGAHHY7t2TxTcolsLw1myvRBvq9Glw8qH/Sg5K4hak1G9cSX/UwP8XvcYTK88tGFJK
HIlLzlE3ynMx59TnzgAvBMRJlzYCacgwlL+ObJKP1/F5kK1Y/X+FqI5PnGshqjkH7zjvuaYtQO+G
/YnhlwZA0iOCbXDLo81nH+4BSTP1JBDSCe9/kGN5Zkk8TmEDPrq3bpqBjxrJNm6wRmeG540AdLbp
A8d+ycNE1aQ1dzcaZKy2XnNzaqtiJMMBtrieD/iDomuorU2zQTlfo4rRQgjbl/gz7SDitH/PjISR
ztpTqs9D70e10K4YdMjaxVgPffhDS4pN4XmCt2JHoqNpTZtxsfLEe0JGovveDBqlo73OXrj5r+Nl
MfR5CBW+XYfa42OAWb2Ke1TwQJlkwr9uM2G4sixaak7z58KqQG4b4RXdd8/WyZPYe1m1qu/ihhF+
rbnhqc3VrVXAQTGyFmdnVVfoiZzF8axBSOyDDQq/m4LdXtKogIDhF9lcAgjFRtJ7B2mLmAOs/blm
2iudxsT8Jr+g7VfpgrZtIYHmf2y+Rgp2SqirWyJEQlcDyci+2cJYs/C/cga5QzCbcY0QRQIOcV4w
ewTwLC5ja/8udaulQPx6xOe4IBLIJujDL0xbecDJDzJ3oidn7Ztm+N/2JgJzMmo0GiKhjPkIE0YC
ND/HumMER+uM8WekIvp4/LGXBZwVd2ogk2RsASxUkzPDVcWuVCQfgQn1SogN87ra/BDtdNg9n1w8
+GUS2/MHR4ZNbsDeoVXgVecdcRdwmDF0PidgHjVBWO+pY3r3fv16LT8KZxOHNUcpaOsXC9Lmt4Kp
R73ZyiP75OwcT9eC8zu3X0jFHA4nxWyOSSP9FFNlSya3kLeit+ILsLVcTZNFA6BIbpVPoDVMmJiN
va2GBFJy+rUoGOxv9GEAwkboCICZ62943UEc1SGx9zdb/jndM/2sKb9NKGd/Ms9Z7WxrjENOqFl2
qSqGBZodapan4u2XGDqahb9hws3o27+cPwlrbgiDdRBUtd1uPIdQcC6bjvriEvssl7euZG2e3eJU
+JELIaXunTygNsGFrSz7laWpiGHbAJtGcMjeoDZUOK9LFJQacOAhBm5g05p058ZEaYb5nfRhgGO0
3wpMNxsHChEHgJojNS4LEsogRuyxsiwSPHjR3yKuKjQzkZNgsQi0bjRCZ4n1Ph27d40ddMdJ3FN2
4EIndoieCoBXwF0GhiEXG2vEfeF6q8avJiebtBtaWah2dgS78GVpDYBQoFaMUtAE/yGVY6z+HjDw
o3NhYRgKY37EKZKUAGJxp4rnASGSEtlHnzNNJCf3pCbvDv53JDG4cWEDhvNekBR5Lkx2Kp2md+59
LrvNJyT8WjMIf8o2zDVRVJim/LPQoE2urkXoGpEQAxaoEp3Sy66ppr/L2F5hG8F5Q9+ZJTKJ9rTA
lj3lzN/yWl22mx2Mv4PjRLaihq6G9a4catoTTJEyUtqHROjsSSrCPEANsaWqTb+Ri+iJ2/SJGWpN
/TaX0Dh7KCBy7ERw5iic654wN2uGsPKSiC5f1QS20SBt6rXT7wp9xCoyO+zU/Rzh7qqFizWYvP8z
9+Ftk+gk56ah7+XDjIUJasLM+2eOCVRZnxLaPh6Sw8tSkUp8NcEt9CTrUrbQZclGH4DPyodtK+Gv
c2gJueUYxegGe8rLKU3knwyErLkzlfMZn00gq/eaNwRXGJf15/t4/70q22nBgZAcdtO8ZUpz9yZT
LCdVIsD/y6GbAkSfYkEgp4uX6dZVZiB5vE3Fz8aN9JVCbbRtuD0VSJA476RA72m4UQP255sVv7C+
/XGfwnsT6sD9aPx6FTgU1kC6vA7LkDD9p3v6KdyCrZlabTozxeVhQSgfdQiHI++r343t1azvW2pd
PTe2jxcsZW0k89HAZcTJR/+vMFRDdWqLow3rYgK5cEZ5CZTe3JPJbOMUMqyzFQN2x5WsL4GBQRJD
UL3tMH43DBYkKQ7PFS64PU637uwoFc4DouBr7WqmSNpXrYERZChnjtPPij22m7Cj90OZjP4Wojs0
b+kkQrtNYEIACyZpUYC3MW0PQvhBBdKGiLnAEvuFxieelF7MHS4EO0ltaiYBF+dT54E5+e0A+EDT
g7KZAfAU4ACPs1hNUef44ebPrpsyqUo14aFey3jfu9Bie1MMWIvVgWH/IkzyoyvJoXgW+L/gg2fI
3rtQ3Xbup/g1rml6wJrG+ppfoh6TlqR9ZiNCJuUUluEWJ8sFEyrnAPtBRydfm4Mwaz6qlbQb5wZG
+/7Jj5AIFbysyezkldiwrklHvnieDP/3Yp+u6Vw0DLNVtFHUJuHWPC4dZMqKpadbwrIZ8G6JJ9ul
6UtzB+r6uHhpwBllvU13qIqErqHraabYAyRCsK7BN2xT9wWSy8WbzrESEQHs6Fi08I2kDBtLlBZx
Rd0J9DqE3lsuCZu8thvp3A34QGfYdTRMgH6JXofakr343/W1UYGIinLOeR29sqpItjehb6P1Utky
jQGWxnmmrnM7xj/y4jtn+x+Ut1GUJ2QN79blKrUOTTpofSXU8tLINx2jmTUUTt39TqacL+zmpkeg
leO4Xt9Dr4g1Q4yYwYfUbgR4b6R8QcBkngtGGdUrQ1jx61O5GAJ7fvdofbXf2bq4ptX2SNZpm5KZ
fbpSd1goHjH7mdYolV5ViVsG91hNVEXOcPkCnOLO7z8UfaEipALfkRIjjIXyYUfWqKfpeXAKM6Ld
UiCNj6k7jNcJcDhqIWJKGifE+bbTrweu1S+Wn0bI06fft3ECRbOspB9+BO/wiSg7S59NerrZ/5Zx
XLlRsEeFCHf5yz6/iQzXgXB8e3xWj+CP0VVVlXfeu4Nc8mzwMhwDv9o36ODgSNb3ZcKk8DIkgNp0
Cx5934JKWt7JwtIrelwySYGzxg6TIe9KHHpzLHrPGAEWnfC57N4+Rq5jMpKyUZAao1blIR/n/J1C
hzDJg2McrHIuq9snOioDwzJGMG1Vu24KWlCB4TXtssqIS7b8BppzsL1hAsjD6Jh1dAoapcx02tbx
rxUL5Gy9h1+POYSyjOdJN5P7cpHjxdF9J10yuse1B6Nf7cOFOc6ISkNbqjJBzkz+3d89NhBt+M2m
u0SHlFWRzRMNuAA/3wxoLDyGhBxqSmAgyJrX8Rs7QXW43ovgia6ImfXPcJ2OqcDfGrKanO6EnqGp
WU6+IDm8jWwelQhKzDXlwA8TdLM+mXOfcSw6cUkorFSmrs09alykXXbLWfLlA/CdnSAdPMr/pzpT
dcF0KDzbmCayGmMrKtF7tcX5FDDDy/Ac9Lo7Kz6QvGiL7JbtmVgA9wL86ZCPhn+qvrtmxfPpTw3N
YG/lilwBFQPAmGd1sig/x/53A1lKQK9TGNQ1cX/TPsj5QL+IUH/+V3kKAaKFujdGeg9LOoVzxy0m
jdgq6iatqLS61LrmJDTf7FvOXSeC7pVv//YGEhm3zAsZVlh5ErK4LFEJAdxTuCb9EYyjgMlBASOL
0G1vVEy6wYfxJ9BQflJWD1XhbR2EkadkfcTc3q8GNYEsKny31ReBG+QuliQusEZVevcvC86+Hibj
VH5SlgFzbatpKaaHTQ+cuQkVsRTzFyH0NuQ/xA8NAzq1X1vHcBu0V4VsNl8LXKFlFBbT1Yd1cY7f
pj2F7f5Q+9CVt0jSrXD6aK2t0U2F4TKWvnHj8FRMUbIFzouWiSPJZs5gdQ9lVQbuTEKAETk1g84V
WZt/VEzhVlwLPTDDQpBa3Jh3BDwt1SiV7YZQshvFWE2AVQuDWr4vBvPB52LiGn/oZBiY+0Kvi9A0
vd2beF049Bsg/B26iILfAViN8QhbLBY7tx8263gKBydV9uCyOg7pC/ilGVW33XlhezVGwpW0EKXL
pDdU7+ABp3LrTPvH39M7xcyomwTfn3mKRUCtDgdv3/nV8h1TErp7zAr+GTopFiqCawIEMz5sfRmu
9YJyCPPoWaYNN9GWjgCZRw6kRi3+gDFAW046aN7xbr+LVn6tSNWM0dGWItRVB9lzxASWMpOInO3L
JEAxdt2aSk8a/ioRv0gJFebIiUoAkOl/XFHmDTjfLVzjBW4dUPifUkZ207S6LsltYTyycgcg+Eu0
VSZQwsgO6LGbQlCzk6JkGSwMR1jZKwdGgVt4ncQ2wq0D7Ct62Zmep4bjAK+Uv4JX0BvnRccldROV
mO8eZKp5exn7Fo+LlazBu2F2oSY0ftfuh4AwaiG2T4xvQcr598kvBUpgHhniqtSMroqhawh2v2eY
ro/dhc4HcOmhv0wmFgq/Lxt49hy+iTPddo2/CV+dViQDOrY2tPTxHuKf/3pMCGTlI/Xjra1Bb8Z9
uN/rTECnXYFQz0a0YxeVXQwx4qLYNk7uQoZfaF1iKA5XQHTowyWawcCSXL/PIe5AQDouI2aFqBmn
3ROT8oEq6Qn5FGMCg1Id0OvB3hxs2lHNuJdyXTFsbTCBe6U3H1QUlGuzXhSblDOxSONsO2tw5eCC
/fBQY7/Pv05lV2YONPS/wVFdgLT8/6mqG4NobTgJ/ihoTlkUPVN6uiy4Ub6w7wPC+4ysJ+XsXsYf
0A6KMVoDXyhpR+VXoQ==
`protect end_protected
