architecture Rtl of Demodulation is
begin

end architecture;