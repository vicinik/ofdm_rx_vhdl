��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�/���\����aT�]��;��:� ��^'�v���`N��}ͷ�c���`q�w2 ���V�vy��m��j�#��9�*��q�2�
���I�������{�����W���R��N+�F�VG���+B"�������ئ�0!�?5]����၊!���Py�%e��(�E���cۺ�-�����g=i�c�>�q��Ɛ2��BG��g���Es&��/�?��Yc&�$]��>��Y�Ԃ��_�|����hr3�e��X�C�wꥶ��t_�.R���ر�]�c�W�?3_�u0��&�T��5� d�l�t���o�E!hId,�Q��߶~�M�-7�=uu�Sqۤ�7�r����§T�=�tL��o0��]#`��=��ѭ�!�l���}�}�o�g�(�K���������p~�:�R��i�7v����q��f���W��W��[�H��@>6�b�ڥ���q#�r�(�hTA�%*��K��q���|jk4�t�ky6����킒��0���wht�|�F�m,'@���S]�M���rM�S��DoB7�� �/ ��^/a�{���7�z�/����I^g"��4Է��h��ӳ۳�lE�"��R�`��&p�M$ |����V昉�t�n9����y�qNS��
��� C^��[�Cǲ6���66�<�N��2�4U�����gͭ�Cӈ+i@S�ՠ��*�ҭ�X�ʷf}�����'�K$��g��v�H�̰��d�o��H5��dQ�-t�#4E�������U�:�w!��1�L�i�vd�	����5p�?H��6[X�C�����E�-�Ga��9���.(>ޙ�B
g�����%�߶����@&$}�2R!�X2�j~�����/`v9Ձ���-��J����+�n�ON����@���N�����|K���>K�_"�������2�Q�s�R�Jٿ��c��qѡf�S��?�6Q��c����	�2w4�S�Q%*V�ę�3׸ޏ{�[+�N�EI�v������U�f��'Xz��P�&'��~7����Z̲�=y�:�����T���{Gӏ�D���� Uv[�,j�����+�F����QD��g�d���1�=e���q:_`�kC�;WW�\��u�xafۧE7�S7�T�>ݛ��tn�����X�0�ʿ���j����o"�D���⳪�<R&V�����Qe�1؁}l�t,[��]k��r{F��􀗈��Ҁ9��vA���G�/W��mP.��{�B4C�w����tɒ����.�k}A��9�O ��nL��$}�;-�U��1���`jP��	�-<_���_,��<]���r��H���_�UʦpG�/Ӑid��1oJ�k	O/gk2�e��1�V!T�̈́M����n�{tu�o��C:��Q�G� ��TAf��x3�����?wk��s�>�x��=�fB�>����}md�M�����a�j��X0�ze��RF
L�s̖_hz��7���cO@�T��2��R�pf��sEx[�}�?���v�����IG�p��s���eB�+�;~U��}GVG�i�aB:B��>~i�g�;��l�~�����/A��mHݠ!����M�ư�s�O�C[r.\��8F�B�)�\ұ	���\��b�6腻a}��/>
�M_i�:s��&8 xDMqMs<]�Ǚ�k��)��|TQ��+M��Ԡ���2]�[%]|�>U�S	�h,d�b���p�F������	[۹vt1ɖ ��ӧ(�n:w(q�8mw��{ R&�t9/>3'MQ�к��A"��q�dQ�N�-�[I�������i�Ue���\�$;�'�,��Mx�������[�ǈֹ/��S���šÃ{'#��q��S�%}[�B�vgʍ��B?w|e��g���O~"yh�G@Έ��U��\�M�IKK3�[KQ����<m9�(�Cv�+���?���'j�hq����ߙ�����>�)7�[g��������3y��[V'��m�Rb�8�:տ�ށ�KP%�3s���Ҩ��7�sPb��[�{Vq��A��ʱ!�)~[jLS�!��w�[z�"��ő�A������i<��D����r��ܑ���d��_��׏bfojov� iI�����w׿���ݭ������,"�g@I�a��>��R�6ZhA��?�7��2W����l;�Y�נ����CO��v+f�E=[4��t�1�E��+�֍\G��HZ=꓇C�9#��/ K@�i�jh���	�^��%�A��m��t��J�fM&ק<]�e;�Ң�yْ��%��Ȧ�+�:s `�U*h�B�r| $����D�������P(���j�D	e��|t�ъH�����;{��n�����̥HKȶJS���,���Y2;>Ǒ��	^����������u�l��N���s�8}B�W�=��)��=n^&� ��W��P_�y�֙n2O���ܔ��m�_��s�򗸚D���[l�miH�&�Bd�Q?�O,&����;5��;�}#�aC�MMQ������M͜z|�@�U����a
O`T<�o�����,ͬq$���ڐ�P_��y9<�+��Zs�y&+ ��vO���-�&8�Z�b�Y��-��6�I�_p�x�1g�lT��x	+���{!Z��_�sG�ߍZ5z��7
Qp�s!������$�1c��]��xi�"^���}I��wꑰ2EY�SY��*I��o�}�Ҽ�+���Ι��.<�.���;�`���B~k���?�,l� ߶*���{�Z
(�Z�Va�|CD�|�=ԣ?��_��a��r��Qq�	Z�gl������(V~�]^Xʪæ	ޗǃq�h����ob�`�����P:0
���q�W4v�n
/Ҩ����.�ʥ�߿����Az�y~MX��[��~�-ۇ�Cr���8 0�h�MP��)7�n�6�C�/�;<�xk�6�
/~sU�(�a�aQ�LH�BP�V���t�D)��.A�K=Y�+۾�6�� B4�+���#YBk륂 ���^�fv��nx�XX�.�R��ZQ�:�U,I���f
��F1��B�mQ�s��c#�6��h�9:�4�: .�#��ǌ�P���A�:��Ծ(��׫���2׳v�w1��'VK�
�`��6WmY�����\8%W)wK'FՈ"@�wx�)��}�V |$�	�Z�X�D3�~��J|�6�̣9���>P={���O�3Q�})[����N�����N��J�ᛨ����Td��� ��S�eE�f$�%Uaf��wo����F~ư/��
���6�o5k�ؿ�ǈ�$��(����ZtL��V/�L{�BO��%��f'�ՄV|���lr%� �E��J��8'W�������]ODT�a���ՈE#J�;�ä�c�D�[��@���p���~�`P��HE��M���ڒ�m���]�E
�/�9�_�X���=���̹�\��+#�����8���2�N#׷˻���� �3�a,J��P�BlK~�ͫ���(<L�b�gV7$pL�r?�5�=�"���R��ꐳ���nJ���ұ�6&h�<ܞ���dM(��P�e1-AuhUo7�_�Ѵ�:ʁOc4����Nu�|����<��W�hm�x�(���"��+�݌�̗���E��h'�.�ɳ���	�3v�m�����������*?;ݯ���{���N�"�-����8
Wx�^�cx z䡌I�ݶA��ў��Xq��4�.ِg�m�|�G��N(l��>kق+L0�H�\��@����X�آt
�w%��g�c�xcC�T��Wa1!f$�[G��<Stר�����zd��;��;�u{Y��.Y��u�%���E1�N��d��!�Y:
��<�0/�ڤ~.�,��8�"W�kʖ�gqY}R2@�+��$�Ŏ����e����|����[��-��q�[t8�z�+Tl��CH��0%�����2��Fۿ��f�S�7'o�B�"T��T>���H�PC�v��:kX�c��H4��Y�hANLT��U���ɥ����5tL拾r��
k���P����tXP�
�v@-�'���?���̽*|��a�p�S>�E����^����L�ռ�]������A����iT�{�Tp����f� InH+@dL�ӓ/���e��m���L�Nx������:V�Q���%�J)^K�el*jw�mɬ����M��r��y����@����=��4�L���d�!��\pL�c�ăү�@�q�[�?3���<�f�q����%�Ӷ����%ѸFi����"�n{����
Z�k��U���pw�|�$HDv�E\�� ��x�U>�8��dXV�\q;|�l�ڰ��&"t��0TeA�,��e��8�iÏ���TY���'��"+y�t7����4���%G;���6fw-H���w"g(���2<���yFG��$�R�w�!�����i���������Ŝ!�|JK��v%x"��L�=���ÐQV1g�o`8�Җ]���#���3N�:��r��㐫����p�у��ƌቈ�-���9����"��۟�����2��w��=�y��r�񲏬tz�gڀ)���A�W��o�'�].�U�
��$�[�d0J���[�$��W&�T�������j���Aۦ]0���g�70�}���(qd䈌i"CD���*��
�)�����]͝�@l*dM���$�Ԥ(nߨ��.���m���4��n4bA���C̶���6}H.�����{a{/�r!������Reb��60X�Br��"��+���B)���UR9ol�*u�� k�g�[�%���'�x�@(y//��w�ɕ�s�A����>��~,91�o�M�x�o�@�,�G-P�8%��_��d���Gg&O�Ҿ���!+7�����!aJ�e������`Fc|��=� קJ���gH�2?M�}y�.��Dͬ@n��	� �
��^~���Y�Tm�N�h�0�I�*�`��x�Q���/@կ8e�Dg�]ӾD��+q���Q������z+ac՗�r�p
���ѫ�Ɉ-��ĵ� 6ehDj)���42���2�93|*�������Ǉ2KEKg�;.��md�v&=��uh4���e��"L
��.��!�v�P�kd�|ڠ���Fm>e�/�����)P�٤��	i�YK�̜fH�����C2�O�cE�'xa\d��BuzΨ_\��	7/����;l�/R�I^��57�d�,�B`��segܵ���7UT�-W�ys�V6r�
R�Z�$#��:��$u+dQ=:1^F,�'�k�u�� �����}��$$���Y���3��5+̞&�&�a��{�WcR�A
�C��j�cT�H�P ���c�kV�ս��y�l�FG{?�*0c��Î~��Q4��B_�3]׳�&H!P�>k���o�bpfq�q�����8�\�!��'�Ǧ8^51�]�Eu���w��j�x��'��4�^	dߝce��<��3λÍ���T�R����B��j�f�W�Zg��b��)�]�-�/�� I���Q]���&?�.G�'��z��8s�T�M���EG�b���6��(��Så,���X�_
2^�{��{����P�4�<<��fg�����Uޭ���<?�r�I��2ע:�(���8y�M�t8S/��`���� �o��6��a�����
��[Tʞ�s-��c�o�E�sB�Qgx[d� �Dfi��O��᱓�~{
��-2�c�X�jb�B��o9����Q f���H�\��<��
���抨La�7�L�Y_�maW�.�b��4�[�~��V��3��ī-t1\�9��)�.r1Y������+�t*�d����ҋb��������(	�˜����C�D[-��:��)�Ĝ���`�4�����1Y��pL9Wp���@�F���(���h?�|cAй|'�­xq�����;}-cn��Ɣo���`M�e	���fT����@�`R���oy6͓���^>�`�B�*1O�T���K)�׹�&]�WH" �>/?�_
��(�9���ec�~Z�r(̈\a{�W�R��i��ݵ��C�Q5��b[=Fje,S��a�Hh��􊹙l=5�g~>2��ܒ��1�ِ	U$2>s��{1-/�����h2_@p�$T[Uo�"��<A���#2"�������0^����.��|�)e��%p h篪 ��y�$=|��Sٴ�涫���A�\4Yҩ������/�W �ӵz�a�� ^��%/u�B��=���Օ���vMA�YՌޭ{)�m�����v��v�`�{��
@%#�hE˄2X�@=$ѱ��7���vQTã�j�X�%1dJ~�.�o>B�>:��<T������o��W��dɩ��Cf���n���3�SI�=OP@���NM�&�i��Zl���L��@�ZR�k�\��Ƒ�mzGh"���N@�Bbt �L~�
`B�)-�:Fv'� �؏$g����u4 �4��I���2�は?����򉦋�����v��p	)�]I 5�����TQ`n��Ҋ<G���w�a���	��T��˴\a�Ҟ���m�;�%�IG���Q�!���Q5�pΗ�M�
��ա~�<q�.�t�e{B�8�����8�����,z�aH������M��!�w/ݍ[�:�ja����{��1{8�L�Yٕ��k3c
 ��� ��!*bܫD
��i��2þֳ>���<���y$hk���<oτ��uʇc�c	j��U�&�=��<}����O�����`hQ�=�H�Y�¯22�^��~�b�˨hA���<9�P�۫�l:ѩv���z1e�Ez���@c/�`Nn��n��8�(�N+,z]�HT�Z� ����k�
B����S�_h�Ҟ����w�Bv�1����ov��Y�x���d�
}�����ʥ��_b ���r�!�h\�w��^|f�10��U�	�&��l��7�>�r��E9���Y�����YzRա��?�ޠ����@ўj�V�p%g�L=��q\;N/s��Ehb�B%���IG��fd�G;2q�_ư�2�لĜ/�Qi���,�ý������f��m4	�~�𳮣>a������7<&h,��C�%||��{"e��"�a!j^��j���Gn��ʈ.V
F����������^�,4ڏXby�����$Sm����l-�O}q�ߛ�D(а�(n������j�lY?��Ї���\}������~�� ����]+}y�q����Eع߇��9G��Qjđ]�D`�͇�Ҋ�.`���֜͹����i�䎺
��P5�0�����	�Z̀HR�0ɧȅ��@o5�B�u�q��6�o]�a���r������'r�^m�J�}T�D
�?!�n�l�$�d�h�#O��Ӆ�ȫ/4&���8�Fe�c�F�C�/60���^=o'�����s�(���7gz/�2̬h���-�{k;�f H�m~�2)�L�z�U��ܞ0�_:a���s���S��/Ĭt$�GbLx�| ��K����ɷ�)z�.�O.8�m�<Q��|Ƚ =�k����1W^�}���!Aފ��0JF	!���ġM Ģ�S�l�R'J�g��d�ٲ��	s��<��CR��x��W����*���^Ýi<%�P����;z"�����g�9��d��MO���7����-%�>��g��[��� ������#T�5��D�d���ܳf;U6��.R����O�n��KU�v���qq!2 	��,8��d-�H����(u��|�
�~���&��*k�d��z��z��Wϰ�S1��SZΨ�G��T���5"dSиy��y��Pq!�`!x��4��K@�uS��bat1)�$_|��;���DI�!Є�X}S'h@<ب�̒��È��ҕ���;e���	���l�wK=:�A��������RG"������0�c�����A���ݘ����w�w����=<w�cL���=Z�X��(/�@��0�Y���50�a3ӟ�V�a��<��4.
`E�����\���&�ݮ��k�!M�<��Ѡ�!��˂��;H���_���4��D��GX.�'���7�3k�z�"�C#�dۓ�����IS��52�vȻ~�g�� �o�D����o�U��G�ͪ�c������^���J��{<Њы!��Y�q�}�l���-`�
�l#U��bT��4)�?��-\��w�ڈW�� �p�uKA���/��B�lh���� sd^yJ�)UO�=~�U��6֜�� ��;��*W��P��#���8��Q���J̜i	Q��z]�4#��v�a�hz��gr�*b�^�f��m��gU#�@�U��拉�t+LR5��Y��<�.['YЩ�\���O�"6�;6ܑs���m�צ�`�ֺ}����a�\�D[Ƭ�7�^y"�q�����t��G_��
�떱�<t�Sua��g���E���0�9(�i7Ly	h���K�ڤ<��vx�aɸ%ø��9�y�m�U�#���n���	{ա���s��C�T?��"��0�=��ɺj��.��Z^CC�.�,��#�+1Б� {���&�?�y�@�#��X�hG���9��ɽ} �i� +���=���-{�K�� "����ڷX�!%�5[��<��,N�Y�<*G� ���$�3ߋ3rd�i���1��&��~�1�^+M���_���F�L��������u6��t/�����Qys"���F�l��I�X�T�o`��	D���ZSh�m�꛻D��Vcˑ�Vcu�_ �7 �[i���j3C�Et�um�?l�)��Zi9w	�ŪIft��3��`�bP�q#�;)���x�I������ڌ�Vw3IQ���G�:�[+�h�.��}4��Ɲ�;K��1�s���(>��q�1����'|��̋&ջ\��� Jm�m%���0�3�TZ���&�Xow��B�q��Y�Y9�!_R�SL_���X���~����h��7��IS �4Jy@�l����j/z[��*�?tāBs^�X9x*F�F��8�+`���KQj �!���)��&C��=tV�@��H���q���i;%{BHuG�|�����H \���j�ڟa����&�_6��08ە&!R{����kO��N�>���d�������E!s͜9���_�
7Vw��{�N����*sHT�~�N��Q1�]���߃��J(\��T��lM�g�A���٬(�h��1��+o���ަJ���b@!����]�JF�h;��';��0Ń�j����%��jO�-�U
�ؿ�
+{f�� ���F�֡+�{�ʤ%������eD��Z�/��_l�h�#Ռ��{@i�5����H9�i\�3"�{�M�r��9]�8�T3�"L��J�X���zQ��`:�`�K��˥�b�;A64�6ODZ�ƾM4��r�ҺQs�|� ʨѨ�p���������<Fl(�Ml)y�"��$����P�Q���F**���/d�]�AXj{B�'�T&ğA=���N�rP2>/���s�zra*�YC>OA�/� ���إ���|`(�ū ;����(��h@dN���|�&�?��#�oyB�Ɗ7�9��=o�4�t����)l�9�"��-�N�E�%4jo�P��T#�V�E!#���'[�����H*,�?�c��M_؎,BV�U �2�7�m (��
�X��/t!�O:U�E�vv��i%WG�]!uP��4��l.BUf�(R�u�ٸ@O�6�3�}��к�!�dH�K��֢KR��L��|����GS�ޞ�����Hǿ쥬B�ny�	gN��yEҿ,�#�\d�b�\x�A%/F���V�~ym���4�>�[��ݢax� ��'�{��q1�'I�}�h��ӓ��~�^�IJD�Qf³��-���[֐�F�g28�Z��҅�����H�
�!���1~�.��ywXe�D9Z���V�ύ6��g�_������:4 D�^mX���� -z1�7��0�!�V���<s�� 1ݥ+����*`aX��D�U�w��Ю����w���|�(���qb�r��jB4���7��˫DJU	�R�)��fL��C^�,���/�-"�a�
�AS5j`�$_�Y�o�+��$��؎�n��o����u~�	�	tn�y��-�g/�8$��Hn]|ME�oE¦#&�Y˜����}���Mb*D��Z���?8m'c<"�V̊V!���#����U{*�V����*,�O�D3h1�C�Mtה�R2H���-��M���)JДy��%>f���?KL�䮹��t��$$乧��,^F�����f�a?`��L�;�T6P�
%�j�k��ؕ�kJ^��X���g���`�\;���A���͢�?U�I@f�ˆ<�@O'3/�)��7�z���9����R���*V�&f�
�9M�B�� K���cG��b����0�_�l�\x�N��o��y1�Q�uu���N���;��q`�4���?�Nђz��gۦ|h�×�-��F��oW ���� '��2h	w3Nk@oA�R�_�s�A���l܂�_>R)��=ӫ���Gy�t����C}H�d�&R��A^����({��`L!����}�vhLy瀶EgK��$0I}�H�l�S��K3��_�+����ykr"�}���0An��@��/��(��	�=�Ɨ�5oK	��
�ý_��!ĄD�\\���"9���>/�&�	3�vH*��Q���T�WB�A�9	���v�[��'�6��;kY��m�}"���
˙�u�11ĸMR����z���\�	��i�:�Ŧ#墇����<(��f���/_�97#����z�0'v&񅕊6�\�A�Ot-L!�ɤ�U��AU��dQ�h�=��<Rs�*uznj�5��.���s�
��~)\O{鶹�6>���7��]~�|�,ۻ?!��K2~����5����
f���#�S	���,��]�l=��\�zۢ!5�Y���~�l�0�!ٙI+�j!w�)6<X'y��Y��o'V�U��$��`�\ֹ�J�4�*E������|��ԙJ�'*�}i��f�`O���0�%��~�"���yr��3��]�'�:kW��?�aƷU���_%�m��N<����Q0/�$�S��q>���f���4�vq�cG�5��c�<@��&Zٳ����׍�6,~_�������<Z2*�T���ۣ�Dr�
���t���H$��%)2�lb��e���ʰ'��k����o�Mҧ���� �"5T#��;�C��`�}Ş�C#Ӂ�*H�� �u�]dT'��b�ZC,d�K��ɨq��si�8�Y=�|2����T�c��\
��Eg�ǩ�Ԩ��l6��QϢi��I���4���G�m�Ć�c�g[)a��4���3hG���,?RQlɎD�,�5!z���B�P������n����"�wB�Q,�P{���5 k���	"����������>uݠ�P�g�B�3\��*q�x`}䥭�FM��z��m��Y[�L�*1F�l�d
pLt>�����_=��x-�l=�p�E�~�خ���g�.?(*�Xˍ#�����E�3�%�����5����goU�+3VJAw�'��O����7Il�C��󢉤����/��f���2K�m(k���ڻ�M�}���y�C(g�^e���ٗ�fB�W�і� �R���uWU�o�]ȴ�F8����h�R_j�z!�<��� oZ����C������S��8t��Qn��G>;��uH{DeB��i�= g>[f���RD/�����I�$���(�84�q���֨:$�1m|�M��O��m��A�d�a����O���9���B��NX���T�����k���s�7�_�[U��.���0��.�d9e'Z/���mC�zg���5��-<.t6wfO'7�>�/�rɇ�� 
���T�n)7ARЇT�)r��`�%��Ϲ�v��_��&�2v�&�B���oQ[=_x�e>_�2���9[��jd�3p��8��* �(��-�D}�Ul���If�����������m�d��M�{���I�2U��Z�Ӟ?�t�O���0�Ξ�)R�� �#�_�p�������@�|����+���N&C�*L�����͖v��+�AZ(z�m����=��`��9�\��㗆�O��6�U�����%q�紖��]�Gi��_�Y&��g�%��T�9=a�J� ��=����\��)d0HU!F�e}G�����|a�(tN{���q毋G�|W��MRKK��"P�?�D���{�P3_x�y�ڰ�Ƶ����?N��o�����.�.��kd�?56�G�<N�������-D&e�O���H�h�iok�N��_'��:�0���tH�h[��2|d�S�NJ�a��i��W����ib@�s�,E���BG��_��X^��c���1�j:�$s����%잿��L��J\A�aB-,��-�j}#(�O��j vW_�۷l̐���DP�ʵ�Mq�����K"���������ʨ��"/dY)�>ֿF���Jܢ�h�jS3�����/���*#�ʀ\�껯)�Da��.9�y����ǀc�q/=���R�C7&�٫�B�}M�����ո8��ؓ�S�ʐ�N�o�1!=do�����I��A���c�����B�ܸ�9c�/�.V1Ą�ǆZW�˲ף.��x�=K�u���ԤDn���v/'7�����P������7�-u��ý�!���N�Vr�L:�t؁l����@�T���ݴ,_�I���a��E�X���e>f|�u��#7�e"�w�\�{:�f�q�	U��m��| `��k�5�#��ެ?6~���PxcP~'�� G�#�IEW����ӔQgw�=E�mB=p��� Ǻ3n���ÿBPJEN�)��D��V�r�l?>�3K���S����c�bE��-�����ǹt�aNj���o2sHE�azx�@g���It�>V�cv����Q�vQ�o�qg�(�)t���W��:�+�-�ÌY��nϦ`�P�=*Ō3ˤ�k^��˚��o���؋>&e|����Z��S.5��
?)�����K#FzM�+u�2��l��7y�d���v��b��N�XI��n<��e�%Y�a;c{�Nl�� :@	�O��!�2�����&KV�(a�UPr�z���K��}�(�[F���:��g�P�k(���a�uѨ��gE�#�KN���+P���R���|]�H݃@�ʺ�@E}?���R�cwIOt� i������)��PLA�4^@����þE5*;۫��'���B���;�lf�;�Q<�b���w����4D�C����X�bΥkXj�����ӭ��O�RC�Ⱦ ��d�oLĚ�?l�nqW��2�9gٕ��`M���Rq�i(���*��L@z!���"p]���N���@^i�@M4��g��}M��$�Z\4��7mu��C�XL���+�9�u׍N�Ԩ�!�u���9��#[+�0zڒ���7Q� �Bhl!4�+5��9�&3^U�.d���Le��Ǥ��1�l���h�F����	��#scs؏N)�|)�3R��2��ը����C�L�י�E����Qe9�B ��a�:����a	����B�L���_�����SR޻dc��՝5�:�5��-���+k��}���5��.�hږ��O]�f+���$��':VF�1n�e�씆A�,[�N?����+G���2J������e⏋s�0U�݄�%(4�|��T
ά�	�|��Q���n��"�|ڷm��K�H�-��� ��&|���������r�a��P>�kFq��ZֽV�l;Ӟ��E��1���J������Bx�{�(3a�{��s���6,�c)�������]�hâ���e�E��wT��ЄVu�SfH��%2ho���	��Xl��a�Ope��A�)�L�H>�b�slm�A����3^\H
�s�>Hhō���'	��2�u�����d��̕�F��o'�J�T�Ako���Os��Bse;�wI�w��'R�����݉Q~�L���)G�f]��}2�8j�U���ӾXo���7��)�1mCd��,�����s��B��鷡\|�L]ד�j���yTɅ1FP5�6��#�/u0�r7�or�a��� �a�Gx��+ece���#�e$e:���'�;�|�W�y�W����l(���om��w��링�Hu�k�~v*��~uk���4��=ad�.C�eة_���K$<�$[�;��~�L�R��Py�K挒�{X��KD[	���/� ��o�v
ɘ!��.>uđ��[v9��B_u5�v��d;�b��P��3E�ޫ�V����?���^�a�\3�B���2��,���{�c��m�~���h֫'&/W�� F���TBŢO��Q�իm�B]x�%va�3���7�֎y^o7$�7G>$XB��~�	
����5By���/�Xo�s�27[�0&!w4F��_�6x���t�6��-��Z�k&t��� Ԉ���æ
;`,e٭�����=~#��K��"Fk9��2���>�+&��'��`IUOJ��ݵ��ȥlw�g9)�7g�Ȫ��%��9�b�����!ȯ���>#�7w	��j�y��qjڜ�^w?=�)��JɄܒ��N�
�;CRU������k�W�׌�.Ri#�����Y-������t���S���O��b�F��&4���Kܲ˩q#aȵ|�O���|C��W��U����αXW)���5�_�BMy�e��f�/��N6�e2�8ϲ�VK*�]�]m�#<��j/c@-��嘸��I�	b��~��Uf9.��N�!kv
��LbbD�ﮑi�^*Kz6 �!S��~%7[b)��3��t�ۈ�5����?�љ��5�����g2t�B_�Z=ԷO*K yo*#,iS$d��(_��L�_����+�<b�o��Qc�|ڀ�-�Fp�$Xw	#�:�j
�ܤݡn�@B�u%En��>�m"�G� "�gT��V���O�+ʤ���Ʋ��c���߀�z=��p;M#�+lB��_�b�i��\M
ں�#�� O�bצ�U�1��ԴUMl��G���bO���r�C1&O�48�6�C��g��p0�44��؏k�<Q�0ݔ�ǎ�N�"�-|��=����K��r�OM��k���2��>���3-��0c_o#����u:�+W]�a�X{c��׳�ת*F\�"!d[x2�����t��E��"$�$$��_���ǢC��?j���n��W�[�or��H�Z��/�,�_�� �pj��fd�=��ĕ���ݤ$�;�B�EA�����;,;��I��R8rr������wQ�S)�:������+ԭ��c>�x-� �DT���,yq���G�"��׸h�T�cN!�5�?�P%��c���Ɂ|i@*���kS%���h�
!�T����2{�l��ыn:��z8b1�����l}����{q;�Eݹ���|H