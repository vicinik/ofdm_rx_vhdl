��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�e:�G��PH�=9O2�ڄ��'t��e�����M�O�Ł��"��],�ۏ���ui��]t�.�QK�����ř��3���p?��;?Q��S7+�|\f�]�%�q{-"v�GM�Q;�7oW� ��߳�$ݻ�<��ύ|�dY6�M�G���JBw�t�_�[ns&��f<������yd��kV#ҧ�񭕦:��٘�&��[�_��mc��s.?��n��h����J�Y��o�W۹{"f�'������a�KP�S��À�x����#8�|���m$�Fk���g���9b���CL�	|��L����?#��X�o? ::�w����բ#ݱ>W�8"��瘶=~�p��[pp�5Kt�F57���_ҲCԭ^�Lk}q�ꄍP�*B���}fJ6;G�/u�����O�6g_��B�3��2��S���l�('M��x^<c�?�G6��,P���8���YOţkd�,E=q���s=�ixD�+J�y�sG�d9ͽ���9�B�>S�h�p��Sg���)*8
	٨i��c:�:tۤ���,�
�+_��#^� XF1�����m�3�>�&3�oScB�sC����}
^���R��cn��/#�fJ�w�j!p���e�������U�q�	q݋���V�r��j��s�8��C�ȢO�ޜ��
��hsD%�'ݬ5�+0 J@���p�&м�D�����~�(�1��Y�S~����6��=h�*���8LTS���x����:�f�	�ez���}Qn���6�ZY)�Y�%��VKwf����+ |i�v���i>��zw7ҭGE��z�pa-���~l��%����ƹ1XW�غ�e���V�c}%2{{O�3R;��a�O�_M�W��y�E��+ws^B;&��e>�3EO3��V�t9�R��*�bN<Us������&�����⋜#.X�#����9�z�Lw���6�I�%Qht���2�t���IeKi9����� U+D���!����5���+�lJC)��wm7�S����q�cV)�K-��{�?v�4��t"Æw{O����SE;�wAߓ�;�tK�C��'���H�t�c/�I�-dݛ����xH�4����Kn����C��\����9O4�D)�����hI��U�%�ɹ>�~��|i&x���s��ܾA|c��7��?�iî��K�c�`Nod�P��� �;H�!&V�,{����<�P6#L)8e�.��u�"(����A�ŭ��5{� �os���o���a�Qrl�23��A#��X���V��8�Fj df�UhJz"�X���C���d����b���y�.���Ydd�����ȃE�j�����6�?�˔����ȝ�z�ǭ=�r�^��I�nh�r�A�3;�<Zņ�m��s82�&,�֠��v�c����"& ����k���?\�0�\��f��T�.�7��a�蕅9QR���;I)y�e�|9%�NƄ:���NU�439T*�������hbNA(�ۚ��k4NS^it��
��,�vO1��<ί�!��rٮy/Z������5?0y�@.�FWta�:��hj�1q=e[t*��,��ȩ6�y@|�N�VŽ��R��)5�>F�M?���=z5�B���T�b�#�D��N$�O������X?���x�����G�8XQ0�Ϡ^I���5��<1��f��0�S�@���i�T��gn����!2�܂�� �X�\t#�;�{/؇͙�Ĵ�B����L��!Q�k2m�����W�g���Z��ж1�Ze	"�;�j\;^��8�xT��Tb�9��c����/ ��-�� n��(�A�3t=j�|C�nڙJ���%cO^���@�� 3��|5W��7ãj��MO�/+��(&�>'�2���ǂ��5 �(�u�Ek*��Qm�p��]:�m�&� ��k��5��l^*�a��I��#=9�&++')�ZK�I�������Ġs�F�U������q�㭓0<˩�6��$���^g�^����)�5��fnۋ_�g(�b`�Ô��e�v�����I:��i1:+�cɝ��T��/�����ȒE)��� ���[��s�T���F�5å(8�|%�'�w�2�K)wU�$�Kȟ�Ү������J�s��')*䗳zSclA�iMS�.%����R���C�{,���D�^bYɇ���]#�r�I+D��v�EgU�p"�f�ެ}���։3�[�,�a��.Io��?�<8�հ����28{�\v�<����[��<��n�\v� �0=ް,��k����rޣX���v�X\�D��cH9�f<���):�UwCJs':}�Gd�Y��x)�j�U)�è�Y�Ǡ����T�,�~qI��o0{�݅D0b�7!W@.���6������4D�΄���w�WoV'�O!W�+��8&f��?�/�܃^���v�6�΄ṫ1
��uP(��{��E�AD��F�|ru8L�7����1��7}bG(k�O �lS��P&��
�mC��F����KA�'��y���P\s+h����J�e���<gp��_�S
�s�F���={�)��
_��F���>7���Ή����S�}E3���I��$�x`+�G9)H�f�a�ACȿ�e�V(��`u!�j��;D�;�X��dڵ�V��5��B���L�� /dA�Ed�.�4�}Q�9���?ܜ�Ẁ�m�W�ݧ�L�j\�;p��iCrl����T�أG���ƕ�κ��E_:v.ua'I�$K@룮��c.����_2�.^^�q�@D��3�C'�8wx� �|��F3�ژ�W���5	�.��O���h�|��ٱ�%�V!�#�n�l��0��d�=I]bf�uun�es7l�<��������������<������_e�Fh}��mn�t+�*���m��s6�7+��쪞����t;9u��Ւ�4��zz��X9̅�|-j���eF��Ǳc�`P�-�b�,�~ͪ��:��i�����[_I�� �l6��Ӛ��p����2��?>�=k���i��~��V'�|9�܊~t�~�[��(�ۧz���眶����<٭d@I��}|'���Ru]H�80�$EC0�(�y��T)�W�������S��+����:�$)�)ԫW�`�XܦZ�!\W"�үT�B𿃊/ƌ�/���E��}��b���WEi�ޑn͸t��z��:C���$��ը��V�����|�5��8Ir�V<��V!�o"��^B��`�J��:�a����H�~Q�lINJ�l�r�s�+nn�nT�$\q�e��۽���	����OU=B��*<�:����P��P�#sH�����r�<�k���J�n��ʠ�,��:�m�ި��se���R�l��|n[A��3LR��]��PN D/�_������2{�udxJ�"����}�@n���E5��@z\���Z��e����q�&c�W��r��Z��
��>
���㉁ٌ�#N��.om&�g2]�W�2��?¢5ϼ+�����ߘ�?@xK�	4�f]q�JJ;��ʊ��(\�.��S�G6LoC�$%D��A9�� |�t��?�+&|�j^�H�Y��㲵�r��b�`=����qN��P�#�=v�V�Gׇ�J�aTl�T���=�]Ր?��	#9�� �#��a�IK�Sf�t�yB�[��/Km���S��!1�b�,��D��Ǌ�{��Á��t_�u��c�9��<�o��cY�U���8���U��|���
�¨��@�4�nl{�+��5��q��}L�r�Tc��K�:�"�	�Np�*�c]��0 �ArhW�G��� ��^Т�Fyz�W'^tត�4�ߗ,����l� �/�����y��aM�+)7t�ЛGy�E
�8!�? ,6ڗO�3�T�SqA��(��͛����A�;b&�.eV��w�)����,;N4��O�G:_1g2"ʲwo=��k��u�H���Z��������`�ŷ7g��)C!�`�3R \P�G��!��"`�l[���WH���yG�JA��;����G��;JT�3h�}���|�B~�;�p�����uv���hn���>Q�����,}P��f;xܨ��:�M;�e�#uq(غ�O���x�n�I	���O���;�?A�46dy� y�?�l�����ON�4(vB8�*��g9�����g~L�s�zC!��[�ҙ ��I��HGk0C8 "w����[ȵ�_�X�	.� ������,�B/Κ�S�q8v��[�L��{�6�9�#�<b�g���UI�������f�!�L����S�S�4�N��ll��g���#[,[��(��-JO�ܑ����6o��[!0�6M����B�J|;����G�[ �M��%Q�ծ�:��!n:S ��(���
�M���̜���!���bdFi�VyL�ڼ
{F��IGT�^�Һ��
�%CWŻ�����`���z��|�r����J[񸌉׋	G�{h9̀My�CEHۙ
#��y���pRLYh���>I+6���P0�(
{�G�}c���/���	���ȋ����6��1��e���[���&�݌�G!-e��wO!P$��I����Ȣ#��CX��+����vup
T1�aB;�A]��~��)�9�#}m1�K��ͼ��R,kC;ٮ���SL�Yo���}6��W>�'��	�i]M���'�f-���cع<r$��� ,��C�t.�)O*
��zw_e��x|�7T��z�������:�n9GF*E*��Ep�,*d뙿��G%\��M
߷I���l$��18����n���m����[���e���t�I ���.�9)�µ� X��5��^��w~�&��.�� y����I31c�@|7��
hTYLm� à�n�:�ܒ+NQ�*��uf]X���^��h�=�?l��&fu�Q ���_My��{�n��rx�5��;n>�yǚC �G�:�S1Ȝ�su{?o�{2�U�Yy���j���z�'�>*�H�qY�	���������i�6ml�h؋.PUh!��_
�R��{�}1����&Ǥ�u��-(�k��Kv��-���*�͸�k�˫�������<���K�KVt��6Sk���6c �"%�)a���'��8R-��T��_�^O�N�,�����_C�O*0��}�Z���&FD�����K�	���2�G7J�W:�`?���]\A���C���ͣ�Mj�k����_s��Y
�&j��������r��R�w�l��:��j_����% ^���x�����K���(X�ȍ�.[U�,�<o.���7��oz�v�Ze�/ϙ�릶���i�8�����&��L������s��j��[�TPq�ϙ X�KE�0�|I���N��P|;����<~�~/=��|�m��
���snS�һ�r��)�hB[���z�LV9t�'��'A"=α EFm􎡏�h��=b��� �Z���|i��_�� gI_ƶYqث[�-Z0�8rhJQ"@�K�bYU��+}�L߯L�.�"\�2��P���f�f�/k�0�N�km۴ҧ�p/Y���$|��5���.�u��żj$�DL~���T���b��F�5��5&T#|��38)�c6�<��7�+��G�!��U��s�ǖgNaX����n���������p����Y�W�^3�������J��Y_�=�&�����˔*�Z����:���&ii���t��&���J
Gؒ.*�/���#���͝~�ZG����9<KV��U�r��V,��9����@Y�!�&�gx��pA	��漳w��&��{��QO��kQ�+]ulS�xA�,P;7檷��]Z��3V��$C�}q�Z��K��2Ϻ�l�UEX�w}X�N�zՎo��S #�6Nl�e��	��|�	�Ԧǃx�#���OCW�r���Y�C�"ꙁ��� װ?��D:P����%r8҃�dv���І���]�dGS��5�,2�ɜҴ������n�<����w�?�=a�a�3�d�6�˹%z�5���l�4�����A'��9�ۮSU��N&�B-�}�e ҮmՑ�k�:�Dԥ'�Mp`>�y�~��A�y�S�䉃y8M}ѵ�P�l��>������hwu���yǱ��ct���ǔ�О��&�S�q��v��K��ۀ��驙"�;�����&�xc;�����(t����oՃH����F,P�S�t�htY]��׎�a��CO���[C�0�R%����l�|���F�ͣdw�d�TN&�Ц�2�T���P�AyK޻^U-���e�[~�O	�G��"��C���{O�Y�N����W�!��� ���q�s�����a�����c�ee4}�TY`����<!OUPE럈���`r�d��}@�%��+���!�5Vͻ�<�v�8�}H?�������x�3�?
�� �9a��  �¶|Q�ۜ�e� /����K���b�h���-��/"��9?<��~=G����~=�%k�P�P�-ύ��m�i��1$ �:��sy���'1%�V׽R�`�q��;�(^�� %�U[e"�Ng²'m�8t`��b��mp�Ǆ�"�L_�Vx��"�7J�C�������>Z�O����vF�&=)�B�H3*��]��!�R��n���d���F9��y����\������廡�\=�O��̬fc/�
9�N��x�~^LL����]����06�T$(;M;%ӛi��W��l U/����kPoY4��=�g�?M��VD��� u�ؠ��}
��N�GL�-�F��}�����f���Ơ�Ԩ�,��!�����š|~X�f�����Y��`��گ(Տ�Ա"EZ~�]�=�$�T��Fc�uj���{�a����i�@��M��}�Z�Q�>|X�b���rK�n۔�Sn���Ehǽ���JV�+��v�>z�$����.F�����=�� n��B��D���IEkeH�8�;_e6��N!u�U�XK�E�
ړ�Nhr���ѥ�^��9}�~E�τ���͍���EŠ����y�0zB��B��fc���l)މc��/�ܒو�����J`
�u��v���ff0P�X$Qc��U�0{���t9�ev&��N��e��Q��cy�ߥGҙ&H�%_�%�m����B��AY��0W����m�%/��wh6�P����X�Z���f��G�h'QJ~ &-�Z��	j�1Us;ҽ^��wy�zB�N�]�gy�V����6Z#@��2d7��N?����SD��H�)nc��W�V�D����<_vZ��L��ۋ�dB�7�(��h��~��da[zWʣޛ���_���XA����3���4�o� *h*hI\f}.W�zM}����g�k���S�(;��Kz#���|��j�`�e~���gJv�M^�-L���#$^R����>��Z�E5p����?��h����X�ږ��ِ�C��1�9�+m��1��f����BK4��'�M ��L�����S���1Z[ aX��=��r�j��/���"�ϥi� �,x�u������ݺ��I܁�oøq���Rh00n����HZ�̮OPʠn���M�9w;a�\B�pRV���i��q(2�f��0�<%Yg/�ފ���r��F%y��HdBJ��c�����G=�x��We��F[�N$l���h ��H�$�d�B�W����xK��j��̓��I*�ޅ��-ܾ�a[+��8fQR�h�Ƽ�+��&�A0y<"�����Lm���qfX� ��J��&�l��Fٞ���	���a��A��7P$�dLX�ɐ��8��'ő��
���KQ��x;'1>5�~��p��&	��R|���@�~��WU�����J ��q���o��L���J�r��+�oYS��Sۺ�]o��&�6�Cb�f�Y��Br�g-D��4��6�ԍߣ!�I6;�����cp.\1��i)�g�Y�����E{�`���&�#��&�D��Q��-f�G��_�Zq��4��sc롾�OVH�����xAkܘ24#M����l�g5h�����IS\O��b��io����P��
:����.�)X'���GKl��z^2}~�=�m{6�k�}����1���4�&�5��f�ӑЦ�g�S�ZJ�����%T` �,���F�Y�����O�qQ�w6~eqO܍�]Qi�Ӯ�┽v��,��IM�H�N�'#Hd|^��_�NLi@������x񿤉j�vv0
;�����=��p_�X?�%˞�Ws��^9˴��`�����Oc�Xj\	e�%��u�qE/+2�X|WRf��7m)��./S-�"�]�7(�«%3��l���H�YH�b��@��/oH);������=9 �o~�Y(ץ���+��;&Q\��*��u$k�Y�7��b�X���'�R��w?���|K���J+��4��X��j�eG-R�;+�������k�䷓�gn�����bha*�نT,�u�e\��� l��� Ř���Hk�~��B�{ U0Ӽ�1���K��6�����SB��2�"��eߧ_��hہ�Q`�3C����!���0[Z��7v[kN/
}��sw�9E�[� *{7<~@w闠��6�UFݎ�s��-�h7����m�Ł�h�s���.+�}:�~`ޝ�_���#}�)!�r3`:K�5$[A�-��H$��m�A?���-����0 Q���j`����|bq:�<�D�\��έS,�#�N��>B型:���%7��地X��Q�,X���:kfv[�?�x�x�th����t,�0v���i Q�S@ϭ�+�3i�p_l��|�2�ތ�n�/��_+l$���{)M��>�"!n―z/�5�Ħuu=��y��'��dL�wuj�d�o�%�ڣn�I{Ł�Ehx�N:we�>��v��Xy�),�oe���L����Fv&���#�#$���!>�	�A(��u�J�(X�1�v���pƶt��&:cV�~������e���q�O�,b©�ȉY�����%��Û��!f��$�X�J6?�Nu��5�$�.���;��aӫ�M����*90�.W�Y�k�eB��hR��:/���] �.������%eI8��������'o���i�Y��!�[�G��m�����|�� ���vz���ׯ�l�w:���n�����b��d@�U��hZǫ���o��i6u*�,��e)�&��n��)����y�U�ቂ�֡��+���"�D�D��q�DA�)�of� ��g��d$���a��eX�;��释�4RT�,��1�ҽN8"���ݻ|,w�|,���U4��;j+� )�n��3��$�vxhotlĦ�B���n풩Á�+�sM�k��?5�1|жw���R�S��9e��>�sTc31� ����B]&�%e`4y�m�����ȳ���>�\���0�L�do0�]���}7�S�z�1\㥥�0w��8/;,N����+ܮ/���>}v�ñ�i|����9�!f�5��l��O�����;IH��֣�GJ<�A����`!��F'��9�߉2�ߑ�{�xP�oP������ݦU+�.Ѵ��d��(e(?_/\^�,���� �
�{h���p��1t��Pkl;�c]m�����X.:Zw�hߥ� �$�� �2Th�8X�s�Kl��nZ�����]^��wyA�o���Шe��s�ʲ�"����K�OEz�.� yͶG���}#͚OWF� ��£bB���j���!�8{ ���p�P2!��Z�#��6�8̓CwF.q��;;� ��
O�����}ط=�����ysB����V���y��k��#g��<��E�M��g�	H��*��4�&�G1$(#34U`Z�j�y�N�^?#s�ݳ��3�-x�k�����M�'�jǳp������R6'��$�p@�b�vS-��{A_�l$�WB����Ū�P[�G��[���ݹW���^D�oB.�Q
j�E��,�����,ۿ� %|fy8��fT��IKv��;� ��s�M�&�����(Pm�'�s��]�d��X/ѷA��:D���m�F`�.��[�(d��8���T�X�f�p�������Jg��`l0%5R,�s;���cϊ���p��q��!H�#�V�~@����υ�mh�g`&�B�MW���{3a�FO����������
b6�Z�li�:��(	�
�1�0mS�4#~|����8�Jq�F�^ 'X]�/=�i��'��j���C�3"`�&Z�ŨH�㌊`|KRʙD�&3;,`O~&��A�+���>���m 7)@/�#@`������,�U�rtb���U���m
J���d��s̨�6ry4�Q�D%�u�z��tZ������P���ѳ�W;��uy3!��u���c�=x��,�X(1����ś�"ڞf�����w�O{n��kW2hI��)��>�a��V�<~��h�:�=���莈g��E�f�t(��y6<� �k��1�k����e�����Ԏ,E�#���:гi�|���u��y\Y�-I-�̯p��)@<����ž�f^�ȱ�Y�BD���ɉ��JP����R1T����VA�K9L������w��S��)�Q�:�0γy������p�J��t�=��?�j*��H�I�PQ�{�N��-�s�@�o�n'�s�����j��nrl�Ɣ�o0ڳ�y�/�A=:_^�������oo����4��[;Ш�;��ߪ1���B�J���|ՙ��X � ����KB�� �iD�N��^���|��0���u�@�Q�ieC�ߓ�fLVU@�L���7�DW��7mm<����n��j=	��Nb&�T&i����b�5Њ޴`�V�Z������fE��$x�7RL@"'��?�x���PBo4�{���+첁���@�-��Q�����"�6��8���(\���㢩�qB��qt��m�C��roD�F�Q���\��K
������ú5Jq�J%J�&�.��)�Z��[ߠq�v�A}U�(��I��r�����n�e~�U	��+���ka`�:ܸ@K���dIº Ƭr �3oi��a$��#�K:���@돦�o@�
G�r2�4МE�
}!��P=%A��Z�
�_�Hܥ e�c[|�����M���Q���Qd~��_����!.+����[>��&(�����6���p.;`�u�`VD��8^�RTqA{��exˤ���YP�����٪[�N�qT�A�lӏ�@�1��cu�R?%ǻ5>�Df���ib� ]y���z�ٕZD7��X�"I�\XT�m��zyYRb5�)}�V��m��;%���2��78_��%��sj;���u�}�۰���{Pnؾ*�wf� M�S\���+&qaIIB*ElT%e���p*!� ���ݪ_�s��r����I��kq,�4����mݢļ��	��x�I�
9�bP,+/w���������g�&[�.�ЌoWנ*���|����w}{��$����
P���*He�Q�	|�[K[ԅ��W��,k��9�F8���3G��%��q��PhD:���l��}%�b���;:��βߦ�XD�~��&��X��A���PR;��~�G��V �v��@X�
HV�2���$���&@��G��|ɑ���n� ���9&cg�3�e�"7��p��$�K��1[�]{�Y>ֺ=G^�tn6C>�+D����'6>4Ɉj�tN<�1�T˾�^��o
����?�g��A�R��y��.�@3Lf�ix�bH���]г�؆M�0W�=e��e�n��l������r�?m�ϐ9=l�b3o��F5y�,Ƣ�(|,���Y��L#a�}9��8�h�m
2!?�}�dH?C�G�Z��b��7�=d��z�z"c'�J3Ku,f9%R�
eX%{]0Ē���a@�?�r���D��^�K��f�tn�8sj?b=�'čF%�U��<mc���jSR|�՛�/��tDv�r�e�o���D¿\�?�s�
�0�oe�?�#5��Mm�����O��Q-��BE>>Z2��F ��+͔�霁U��1s�A���`��F~�����c��1-���.����"�����NU��g���)��Ht����-Yg<G���V?oFi��|�L"��;<	*'r1��Ի�^���
V�$B��V޶��(���.~��τ���*�. ;�w��l���z5��$JH��1����0�b|X��-E�?��>�<�G /`��(yu����$���w��o��c.��T�PcU��V��YW�����	�����=_L6�8M��
`ċ���zX����jph���&u��s�`wU\��1����,��+��d�.�	{'�t˕�S{0���jI6���x�����p�r��߹�8½�uL�S(y�s���a����ؐ���a�4#��� �Qm͞	��
�J�):��+���ݫ�j���Lk� o�Ǖ�����dQ�衇+ �V.}Y�p^ٷ��^�;T�纸��=��=r�/ȇK"��0�M\�D)��Ȍ�5���X�Z��Q�!�T�M��i�@����*5起NŖ�v!ݿ��$^6r*vY�ih��N�g���y����hD�Fc�µ_$���c�nEy���:g�e#��TJ+*U�k[�?�����}[��2� � >���ZLn��,��N��)�$"�{	$�;=�MrC���]I܀�qA�k�@/���A*�W�o��*o���d&��A���*��rU�����|�^z?�'�Œ�HYElw������XS
/,O2fX��I��d������� k︑��,h��EPjB�k/N\s[�q0j��h1�F>䞀k&�(D��� ��7���Du2��tT&�we�L��ﰎ
��a͛9\e��:���R�w@8��=�
�ey�8��.P9g�,P\a�W�CR:d�P
\���R �����|�����}�=ߒy��ѡQ/Bթ��n�����aN��70�8��W�J�{;�Oh	Dt5_�P��ь�;ܶ۩�[|�0*"�P����H��0���B�C,����RMv���PZU�q*�-b���:�o5������:���Bf���Y�U-���S +�V�BN%�J�{7�2Gmm*�����Yf�b��-�L�2��5����j�bZ?���A��\�T�'�X��[H{ȳRf�t��Qk}W��$To7��v�iS���nΑc��;r/���q�i���W{=-q"&[���U�k
�F����Z��O�^�|0/�N��5M���iԎ�=TlKY���	��8�yV�!R����I�{��l����tլ+����IZ�Ke��h�\i�>,nw���~v�c��K��9��~�&2u����{��|.�*)j٬Z��/�eQ$�᪾�-�9�}{���o��붫�@mjr�C�n `}C���mB�lY�"zqx黅�-Y^��\u�!�������$�N���(��}r�A���o�a� n3��T�5(l�<6�P��Sު��k��m�e����\1g砦��ay��83�CW�R�9ڊ���+���G@]̞��S(R�0>;���q��0G�}c
���u�|��{�0��R��6�KH�����	U�S�C�,d�1
᪻Q��B�i���~�ܦ9B�!ѧ�U�l�g���fS!Lt�7�G�gJ(��dU��k}۽�[��%X�:rE �3w�)���q��_C�Ꚏ�E�� {��0�ђT�)K��q��}�_ʘ#���;��zɲ����1MdR��;�>���#�+�C�o/J�_}��5ý��e���}m�4'�c���]��!��ɷ�}MC��RZ/���z_����C� w�8�T���7Ik�,��\����t�o�����Fq��L�7��̾�klI)�r��@r�TF�$&���WU��R
uŎ1�ƽn�$�և�*�1�?��hx�q����6�{%����Hȡ�h5&�6x�6�����!UW�_+�ej��u�7`"*3�����P��h��>��j�8��mF�~�*�}Hg2�
��*d˓x�����"U�c	���F�p#Y�w0�i���D�D/j�i�>m�m<���M�a
)��LTR'��g�4�5C<-c;�����n\7J�yZ���a�h�D]b#�?������E�_�8t_���Zu�Z��Uq@aD�ى����.-�=b�@�D����yTi�n��ț���2M�g!�V�Ja>�WR�]�$(��p�Os��W�{+ �Ͼ�=�6'��a��6~\Z<�6a�V5*w!ͤ��a��D�I��0�2#ނml�K�=�����^���AsP�ҳ�	�$nO���&���fO�Ѓ�ӫ�P���cVԉ�{�~���p'tzZi�+7{<Tb���އ���{�PÈ���C�P���<�+�a�x�j+Q���u9H��?\��~���fG���������/V��xIxD+l�v����Ic�Y�p�Ak�f��D�9S/J�;�>�*,�N�CMU;��$�@�ȷ�O�]�A�'���6g���8��e���9(���̴�;~� �.���8��d`�$X4H(�ʢ��q�Ε �M*w���H�$��2y����:�5�pk������d��Rح2!@=b�4���{~(d�.��o���!+�����VT0��躔����}���G~��YW�<�7o���!�/Y;.�m�j�ø)Wgq����|f8�8	���S�߰��}��>��u_0&�B���B��^�<"�nS|zރT�^�d��:Ja��?5�d���m��C�,X� ��p��q?��ׂE�ѿ�dz�l0���laK�b�x���	�W<�'oMd��	�@3�"�q:J���%Vr/��B�9��P�Tjlf*�7sj�� �����."��A�M��S!1��_������8M�Vg��mIp����r���_����QdVܗ��l���jj�M��bê>���!�X�չ��O9��׉e���4η%(�+g���?���F�gJ�Q�>;B�6�ۛJAYd-~"�vmfs_W�����ǎ�H�☻�c[�]�DU�~���"C���Z�%�ڃ�W?���;i�v��W�gCy�C�Qu������4���٫���wU�
��לg�z�����J\��Z}U�E�5\�ד'A-4��E�Z�S��Qg�⯜������Y�ݒ��G�7����O#�����O�J��)�M
$nm��x�J���޺�gg
F��� tv�|#p?dI[�n
	Q�*�}j����ð	����X{�^M���=8�b�jn'7�'-�knDS���W/9�I����*h�)��^7����x�ړE"P*vѶ�����HDQ�p�n�E�GZ���XM~��cQ�E����Q�#!�t}��ΐW��+��Gm�_3���P�,`W��nԨg�Z�'��"����|k�JU�G�b��q���0M9z�?��0<�y�����S�n�lN/Y�@{c��OtCW�^n��e��N�Pf��q� ۱���@�c��9���Q��W:��++�f�{��䕡��`
7Ǻύ�k�c��3χ#H����f.J׶�L�:�W�O(q
Tr A��oin�5Nxf-�Tҍ��|��~����_[Q,xb��er��,2�޼�Qg������2�,u�v]���v���2�NX}������o1�2c^��c��9�z(�^�ɦC��G�~���2����NpW��^�Z�4��m��dJzs�>���.��&�P���3I��7�O=?���?��{�$6���|������lo|'�p>��ׂW5�'3����s��)��S�LN�0Q �� �_����_^�?�j̛�G�ld_#�g?���:�k�q���(^m�#�ıg�R�?��Cr:�(D_�	��fMؔ�X�����Dqg�H�7�?>iL��qk9�Q��Iw��!ø�u��%f�j���A����n\&AX&ߓm��%��3�;|�z��������Q,����"��]�o���$.�~.+�ʟ���q�� \(z��6,N���T�!��d��$�ѡroh�81T�FI����%2�a6�;kLԷՊW�ӷ}�Ko�l�h�
03�v�zi���j�?�R�
� <���?�.Ma��'���K�1�%EX��1�BB� xǵ�����>}��3���}������\ve�~��K?�,���8Y��*!�Z �^G�46d�.�B�`��/M�I��@{p�� ��|�Y�|"Ɩ����q�h	���te�:���7%)Cق}M!(��7��n%���A�ܔ��!�vۥ)@�GI�K��rH��Jx^��0�K��pR�{o����F�-���b�E�l%�Ʋ���[�r�kx,v��'.��n��a�U^�����*do�b�5��h`DW#�M���i�>H���蛳�ܽ���V`�%�+�}0_xL˨l���ZB�;��� �g`/�s2�^���l�%�9�ܹ�M3OO[{�PIL3?,����#��j�ɏw͟>ضQ��U�n�d�^'�خ�`�Qq�"O����Պ��k�NO�����j�h��z��x��[b��A2P+����׌-� ���my=���Xt�c�JhO���B-uȫ�3��{J�73���I\��H|���+=��~";)M^�@��=L$���Yb��|+M)�ױh
w�D;�n�GZ0��g��pMq�λ�oq����Jw�W��0^A���%ɜ�h��ųg�ڔ��L�7�٠�ި��
�HV}tۋ�2U�))�e�2E���})s������F��2 �x��p�X�h��޴.<�ǋ�A�i�>y��O�9G���V�� �a�R1��=-�m����Pv��>FHw���k7����4�{����.:^��I�|��*PT|��0R�},��3�޴��96|4�I��<���_C`M�Uް�JN}R�k>Qo!�ڭ��&�n��g�ԯ�T�N^$Qj���j���|�[��GB�Rx��1!��w}	E*zx������v��;�o_��@��R9�������*���4��#��Y��|��f	W�f�]QT�] �'0;�~�SO�Ѹ��Y��E���eRB�bw�L��v�߱���̃�|�	�S ��8�������%�|���3��Y<%cۿ���:���N���SӉp�Yt� wr��4��1�]�C� [�Ġ�J, ��0�X�4U��ds]���V�dG�hp��TC���Gw�lɪ��#F��.���ʀ���M3��b
�=�#�A�������8��(Ŵ��G��*t�Vv2�N��'	���d�g@����,���1>`����Ld��7!U�� p���3z�CU��`FpkӺ���������ѨZ�c����ܙ��J`2c#���>��G�`AH�~����y;!i�����?a.`@���DQ�Qi@^��I�� E�,�v��8	���JƤ��6�MbS>���@�h :�"����|J�+V�GY|�#�Aj��z����B�ȹ���2�Y�*�&( ��bz=h���_�_�(�V�k�uu*�)��U��>�PaZ~ni ۴�>�|(F��XD�I.����k=��{�x�t�:
��iK�s���C D��oߙޯvx*ta���#���z���C�`7o��G�����t�K?�[��X�^�����{ ��� �V�h�B6
��H��viNN\:/�! Üt:l�1rb�h��	g��0�ƩA���Ky7��fQfEI�n'%
9��5MP&�9WÏ'&ƫ~Ѷ�W]���?� @t{�r8����Uz���/H75�az�aUx��d����`�.�!pz��]퉂|�J=A@oq�����!��5�h�"y�c���a��n�sʐ�G��>
#��<�/{���%��L��^�= @�.r@v5��t;�A����S�qu? �E�-ܿ�k��@� ��,�����i@����/.#���)������࿼#��l�:������Q�z�f��;V�y�k/�g��o�-���J�?)Bt��Q���!���/�O,�/H3�ްJͣ�?)����J���e��ܣHw]>^�,�f�b�2XEMG��٨�Hx4��l�v���5�u٤G���;�=*��� ����uw��9�k�w�Z�בd����!�:5��4���)�2f�8�:�4�O�ͭ��d�$�
Q��$���|_-eY��&%�%������jE,�o��uR��H�|e��?��H[h�CQ��tT8�F#RK�v��f��2���F����T��$-7�����Ę��|���_TI9����$�s�=�ǿ���&�Gw�@�$ׯ��b!m�E��H��Z������i��1ƒ�"W��)�|R�~����?��?6/h�p�Ul����?y��x(����I�ɱ�����
��1�'PAA��|7W�띢țm�,n�BH���%|[@%<<[�񛙼���}��0��z�̤�D6��ysˆ�|'@*t��KK��-.��'=3|1ͅ#�)��@L˕�����9��w������`���Ig�0iyd����w�+H��h�&�-1��J���[�����/��W�Ix6���/1U�D�[�^z(���U��{��eS���&�Z��#����~�:F����������S?�I[,�)��JʒzFl��I�9�'��Ԑ71�'&?�w���N�y��i�c]��J�&}!�S�-�w��U ��g��g���:e ر`���OA�ׅ� NC7��J5}	��,�<�\�P�75�ٛ<UP>����f�T����Y�}�a�1(W�Ue�E�5�^3��0i��=Ȼ��y�iVJк�Q��P/p��}w���
�ɶ�o�P�z�;�'V��!J_Ҧ�j�#L�(��Y1�0��b�azc�K��W �D>}�D�9�s"��ȴ�� ҏ�wVsr@�#�୧�ڍW��@'�Ƹ����1Q�y*ɩy�<e�	˿�Pq\r`c�v��ݽ	�!���W��Ïfr*�X�보�?r�4�k�!&���������tS�����}�1���
c�Of�crN�qE3a�X���$.���zlNy2�GZ)D�����xm�x��596���!EL�p2�T�����T��}����M�y�+v_7�!� �<(6�={j�K�wL��c�〫��AM_�2�6���B�0��[�<v�X>��(cg!hqe�E ���wH�C%�Y�%�ӡo�i��|y�U�����jI�c' s�ד�No�e��.JSe�<Vp�0)��ϙ(3���E�Z�C��� ���e����|-hw|u��T���Y������dEn�^�H�gS��XCX�Ir��k���!����5QƹVw��lK8=*a�/3F�Vx�*�%�D1���(�cn�RU��[�1��q�V��Zc3e���CV�d�;
d�F�#�>ڳ$p}�FK�*\��9�V#|�'7 WOQ%}�-��Z���:�J�1���m6�>)��nL�U�M��X3����L���rT�e�#c�4���q&l��o����߀��m^�7��'?H{�!xw����>��!*`i�-14��؟~���ܒ�C��w=)�o'��)k-�����vh��b�x�nt�����%4Z�K�6�<+C�ŝ��{�Ӽ$E����$�.^<n(/˓㿑�3'��\�Ō�d�rA��L���ǈ�J��[tV�:��P�a=⏳�]g��G��F�"LY�2M,�lp���ڮr�����OK<�����8��!�;��S7���?���5�V����/��=c�L%u d����g�E��m�`H�-A����+��b����w�gD��O��1��z-�8߿QPA��ͺ��6��q;���]�6�ՌY��fL��D�Bk�K��a�&�K-}pcQp���,�sm6~DjBU:K t���XD��=���˲���.���M,������#�
<��^���8��Kp(�*��'[o���0�z���8J����d���":�Q�k~h�Qw@lE$���S�Zb9��+��>��^Q�E@"����ͥR�Cu�e9��?u�����a���[*���:�N��Ŧ�Y����\"����<�83Œ;=c�8nOB�F�ɖ����L��_�&j0*��pQ(���⌃�u,��Ҙ*�#��F���k���U��O��2�����]�ۡ�G�OII��Gr�jd�I�5k�oxJ�g�����d\6�iP��ҏk_���7E
�)0-x0�H���L�h+��gn�n�NFd��U���*1��\�0"Hť�tDN��?�:r�]�<��	.S,����2�6䩨�#Wk�|
��˼�PR�J\�`��+85P�ˤF����zKk1	��*t��,#��`D��G�e&\�B9F&ŉ��r��E4i�C±3Q&)»���eQE��ԲU�?�!U�a��6��&| �6��x��Ej���u��5g��~�_w���9�MU.mҞ`p����/��ĆCy�̔�lr�CV���}5O����b0�2�v6!�t�1~��=(�=��m#_=\�	ؾ��G�4:�p�NP����(څ�ʬѨ#���6qB&�?��-_SX�]�)�����'S����qhC�vă�8�
��_��,� ����grU8�)�K�T����{����9A�����t����E��a���T�\��C��/O]���
���?"�d��-X%����Zx(fJF�B�ۣ[���Y�dw,� �JA)��L�a���:���n�r�t�T�p��
/yAD��+�M/�D�Å��6ԣ;�y�c|UD�c�=b��V�L�>�0+������ƥ�M࠼S�@O��x<F+��eG��� ٫Ii���7�6��d/�h�Sp�?!s�.�/�T���I|�&��ηU\�����{X��p	�Es:�'�m*i汈�q�3N�$׽�d�=#�" ��J�I �I���<�-8PL3���,�	(¹6Ճ^��]Dɪ�t�.�ӽ�$�ͯN%��}K�L�̻ͬ*l�_���2�Ag���iy��S��d�sԘ�}R��_�����e�/����O�p�9�$%�$ _��\�1����YV�;�~!Y(|t+��Bp���WS!)�Z�8���g'�m��*�v�$��Z��������v��|ùW�j��$����3#�Õ�|$�5bc�i!��������O�5��-ƴ�Ϧ<�!#�ݛa��yE	��F[fQ.7	hA:�eWR�x��1�\v���.-&7�yT���.^������+~��h5���.h� ���Q�[r:�\���ū*���K�!X�7� �u߹?����΢��o �۳`0���(j�<���e����=꼣��ۥZ��o��M/pÑܛ��%�����ŕ��݈~��/%DcJGd�Ӽ�\q��(��=�M�����Z�UC�K~S:�^mO���G��'J���F�"�����S�'��N`�˴<�~�����=2¡@�h�kM)��ŭ���>�b��h<W�N��s�m��cT(������Ɏ�->��/�8���cǔ�ʙ��� o�/64ro��6o�M,�+_�u�#���|Bº_N�	���4��d�zr5�^���3��x��-Jf�5])L7��g&����	��A.�opQ��A����������ܡ�6���e�5>(�G��&���Ìj]����y��U�E��W����:ӧՌ�b-a�%@js��5+�k�!��l9�͹���]k�Zݾ߹�0�؞?SO�
*~)o��ړ'���m&X�n�IM3O~��,g�N3�)ٞ��	�"P��aM+�.�,2��r�d��ʈ'�?0���'M���^�G��D�=��]��%����)�Ŧ�����a�8BR�gCEm�$��˕��DmK���k@�K-d/�n4��lfz�׳����䔒cz:�z�N6&���n����Q�L]QT{���5���]�n<cI���]a��'�;&��yn�Ȇ[�fr;�u.$(5ݎ�#�@k����Dα��xk�V�Os���g�Fa!��� �/nQq����v%Y��'�9u�Ɏ�Ӹ�f#�
W������~t�}cG������	0{�����9�I��0+��B�va���x���[��-��۬CU����B��i)ʫA%[n3;�������+VU��F��n��n`��,�������$&�N (�`Ĺ�u�W]M�m��~�t���*�j���F���#z��A�X���iiǁ"|o#ʺ+�۶�}��H8Ku�<��ߞ�	Ŕ�u��,x���&R������$�v7��@oE�
ɐ��1�]S?k�嵚u�Ҿ�e�a��D��^�/�?�N�px���}$-'�8�1_�[sZ�0����N��Ẁ�0p�C��T�~���gLkRW�����~dմ�V�MS"Uh��fM:_���,6c� ��!����m~![�c�@WW"$Ű�Y I� �A�KR�O���� '� ]��%Dk"9��=7����o ��5��}�/��Ź6P�l��E�rݠ����<p�c�b-��=�2�!mw��KQ
��YK#�䵨5V���K�������3�ڑ���C��e�eW�[�n3�����4�������Įr�ƅ��50�D��Q!5.��F[���4°b�̊�Y�Nw�)'��}(=�Z�C$ ��M�Y���C�D*���)�y�07R$,�U>��^��3E)A�[�y��~m�W|i�o��zH'��&;Ǹ�A7��d��y:�A�ǧ������xp+�	�B���;j�G�l�@���y��Wn �%f%�*=F&]a�u!ИTkn
q���}�)A�4��Y�#���DO�U��fmC�Io��/@m7N6�d��J�]��k'ҀXʶԂSNFQ���E fT�X����'ڃ�M�f8����n$n�Q9
��@k���(������s��\����� +`On��+,r�����%F��"8�+���d[����Zb���&=4����h/���bu���A��ya�����T�;RO��(���j�N4��#4 \��l�\�BQA2=�(�(�o��@ܓ's�c�� ��Ʋ� K=���z\d9�K��3=i����ܕ@�W��T#�-b�\*�:���O��銔)?��=��^���8��+�c��R�7(ikj����D����y����0����e��JS���3� ֡|�Q����غ���}Ȥ�nGL�-
4(�j��@,��2N�+ߓPz�c�1� �i���l���S|GR�y���E�è�}ay$ҩ����eAg�?U�*ru8A!��O�%�Ȏ���[�7i&��Y���B>����j,ʣiE�3M���r�\E��`E|S���[����=W��<��&��W]G#¨��K]��S ��ҏ���Dm��.<�mc��W�}�Z��_O@qN�<��˧���n�\=��0QMF�U�"����QVe5L�JR�,�R�b��,��\V~���b��&�&x�us��]�&<��D#/�I�Ϻ����R�)��z[}O��D����4=i#%�@� ������d�H=���{A��)���@UG6񆈙lfw��p�+ɡ|�B��Q0vkA̋E�Nn��B1���m08Ϝ�ٰ�c��x\�/��iRr�?8.�)W��. p ��c���LL��A����G��?�O�=F��dD/#0����5T�V�6�Tؒ�vE_�$��
梙q�-P�\��^�� :�e�cz �l	�el��n?����� �wW1ppT(��v�&���wDk �Re�1���Q{,���I]I���.o����Ӈ߮ �e��q�+jFū��ײ�-4�l
K��Χ���0���x�O��5��^2��=��īhҭ�0�;H[=�a�%&("/hwP��� �	[.*ϼ�g����g�˿L�w����g]#���Fzk1u��QCaT)P�p�ۦ�}r��{�7}�y	q�D���C�>�qA�|%��4��B3�B�-;3���,YS�G�;W��2.T�F=�1.C�/��^��B^�)�dńJ�w�ߋ��WN���-a$���M�1�[|+4a<"��u{?������5��ϛb>F_� (W����8o�'�u���da6W���\�@�Q*�+_	M��G����������@<*b��wo��P�_@�%��G C첩�yPh�P���~��x�ZL�����h_�����/zkJ�2+])�Q�	��O���u�\����OʂD�4!�Y��u�ۭw|ԯk�Ĉ�	�O79?	�9��ˣ�\L�4��Ю?^/LOs,x
0,��'�\b�]0�Ւ�mI����W�M|����gW��8L��I��ŧe�YH����>.X�Av�N�ٛ�BT�o@�̤^������aÄ+v�S'S����/ >�q�8{�2r��ͮ��bHG��7ͦ��;���1�z�d��|�b��J,Gyʓb�G����#�&L�K`��n��ף,�:�܈�҅��Zu`c���R���a"K��y~���w�7�K����{jIj��{j���b��bU_���<I��|�vӂ�ՙ������1��`K݉\Ҟ�b��J"���Z��dX^i�����I�W8G�?�+�2�B�[�X�Zˑ�%������[	&U�Z
j �����\�oQy`��]�#�or�rZKν���+����T� �&w�+�Q���\v�e���Y���}���8�v6�T��Sw&������`t{�בt���<�:m��
�^�ɺe-�?:�$.c��=I�����q��4U/��`2����Xh0��ū�ןڳ`
&E}];�J���~� B3�`�I�I�(��DY�?0�ቡ�=�B�A�{?�U��Mj�T2g��bI��*�0���i��{�� Z裭�l���.הU�'��eV$1#��`�R9[���0c�F�㦕� X�Y�J��_	e�X��}�Ӯ.�2�$�����%�s\o�Mj��k��_���ںm�hJy�
�TC��XT�f�	6BP%n�%�Ș�eD�B�٢�p�wר�>��W�S��p�)���=��edv���TKLϖ���s�a�yk�=$��1�~TtH' �P]�5�+r]��	`�]�D]c��X��&��/�P��=���]�8���l>D��y,��[S"�j��ԕ��,8a3u�mc�R�� WSQPdQ���y{�$��yU|���ַ�GjL�s�2�Ԫ^o6qlu^q��F;�E؅]�>�b���v�2c���<E�x�ZYB�v�R:��\
�d֗4�a:54O%@D$v�=��Gt��{�G�M�
��p���{���&HӒ���ܥ�ֿd5�&�mE%�����Y)cz���zx�!���; 6U�$O�nݡ�΃��B��䖨a���f��E�>���{:���%Q���׼ �_l�@��g
��Ejl��^��ӓ4���R�W�,��L����#eZ�Y|8Z^�:�վZ�*[�椔9� +�My�oyW̉�#�t�({7�IG�����V�l�"e����f�׎��CޭFV�v
�"��y/fݧi�'%��**�W!}%ē����>�>s/�q�K�_�+Bd0��O ���hN��tLr�{�v�2�r�Q�S��rh	ޮ��Lo�)#�$�:F�o�M�Z��5H���2RQ�&��I]�
�Z �~)I��DJu�	���%D�(�r�IGߣ���m��<�n9 nՓ����IN��ma#��#��rY�Y�_]3���E�&�&�<]>���|����
��5�U*�lEh��\=@��� %�$i����z�n��jUy亂��հ�|:|h5G��iH1��7�}��4b~t҂_>�����\�x㛡�@�'V����8|���A͖�d�~��	��
�u��P�c�� |��Y��Yʤ��rT�e�M}6�Ec�ۉ-�j��^Q k	��qo�Q)Dx�Q$�;�-� 6��7Ss�m/��c�� �f�H(�����(5 �ƌ��+���8��K��dٽ��H��#I)��:� ��[8ASf5��^u�֨��4�ީ����^�����@5�w˽�m��;�u˸���t�GN�NeG(0d\��(2�3Qao�^f<��-�`$��[@G��=�
��#�q����/�T^�uT>����������;�L�m��{�&�+X���ƚ2�`QR�w2���9���ؚsod�m�ޣSއ�n \���x�])r\_�2���D�B�76�猪�~u�U�DF�v+�\���-n���z��4b�[�<J���ehLg]��}ڶ�wM7�:�R���G۟z�7	g)�6ݑ-S�'z�WC9�[���UO+f�V�a͏V�Zlz��sy�K�j1�4� BŞ�S�D�h-�,>x�Qt&\�5�sӝV����EA閟�k1�[�Q4�F�a�6�)�u�=�t��6\79�Wh_�&������eˑ�o~0(��O�����v�����i���'�Qʀ���I^|�o��Ǵ��[Q�,�����=���i%�ŵ@h+�f�josd9�JHg�)�$)��^c��S�o �������=����J��OI�MLI�\1j����lsp��i>��3i��/������Q�νʰ�ak�n{wMV����L17�Ҏ�q'r��;§�� �u;fa ����_N�R�>a�� 	���b�l�t��`m����ZظCH���]-y$�ڊ[7�����m�g�H�#�su��5�`�w��$\����{|����Ux߮Ɍb�������$��('�n/���7JG�z��(I��vk8�1���z�)�~G%�}��;�*����1X$w�3��_/}��K=�|F�=�|z�
utM�;�0�x؈�w�������lT�]|�&f��tZG�^��`�(\�JF��Q���SX"�W��b:��Q��m�5�
��j�-���0��tVR}:�l�4�Nך:��$x,LK/�P��v���?=������snӦ��� J P2����f��!�6�ە|� ���zS��������,���t6n�:JHM�v5����o&E�y�&&Χyek�f��I�p�\���~�ϛ,Q�C�N���O��ڊ�M__O��)���#�[�9�a����
�B���@�D��MS�b����9�����GE�Bg��w`�<+���tQM��/6|�gt�a�\}_����g��?��T/s�z�!��& jl����O����ػ[#�_�0w��a��:'FYn9_���Y�?h~Ԯ��UOLfV! �K���u�p/��!:	�vW�I��F��p��Q�3�o�b[O8ҵx2og�@P��RɈ�[˾vd�g�'�|-���f7F���[$���YI�ġN���&�L+��u��I�-< n?ğ�k�/�-E�:C����(���%�9�J�k�m3pg�z�%��	A�ռW昆Ws����n�am�)�t�)����4�o�Wq�T�V�K�̥jK��� �50T)�B�j$?�L ��04�_sW�=�ӏ{da�-_4A�}��"�W�
��wRoX��̦9}#^��H����^:�i!ضk�\�ҕT�]˚��%\��D5�̳�'���bT���k6e0po������X�0���3�W���G�&G��ΏdT��);�=�T�vܹ���<�fh� �.g,H1��1�:�6Cv$�@���ǾU"����>����C�oT	�m�o	%ߒ)4d��z��\;�!ƥKkI_���n�[[퉚� vToe1�!��o���%-	&+ɜ���5��s��,���0�@γH���/~)�Jm�LV)H�>�a8ȱ��o�{�p���Պ��g��,���4V�IQ�y*|[��(��2�㾚�-�m:�듃.gۇH��%�h`�0�]�����f���#qťD������*����Q�e����b@Qn��>�ā9����,-�jm�kZ��q����e��Ѹ�ڷ��4��lbw�;y��`��5���}gj�R��-�R�KWz!��L���QMN)U'�j%�^L���A铷���
hճ/�e�q��xF��k���~���P3��!�;ՙ*����[�<l�O0����qR��M�.������J���Ԡ�Jz����=�nYw��`6ļF��i7kAx��o��]�ժ��H��z�����t�/ �ezy�� ����Y�I�rX 1�]|,��`a�F����\�{���w�	/`��[��N��,tla6���x���E��6������ˤ��+�R3�����T� ��ؙ��>;ǈ(��Թ6�ڧ��k\&`��o.��.ћw>��Q�����F�6�ҫ�)����1����rA@b�6nDL��z[{���-�u�5I�>�؜�ؿ
�FCO�������ճC�E3��Z��_E|��?�������L��Yu�K:��/��E�;1�U��fE�b�T��sӜv9s�zmz�g���s���7�5��ϗ��<2�FD����c&� ު�f�|�4^_Ho��T�CTB�"�<._�(`#�����V��n#"��c.�G1�;=]���02�L�� �&��͹�n�&~�4�RtM��hI�I$�#��@�ɐ�Ñ'���U�0�4l*�%��,��vPJ��XI/m��MkcD_rO�>��/����	��!�Q�sAw��R���lW�2�X����?�!�>.�4�m=�O޵�;�a	-m7ky����~�)��MP70X�8-$�tl���#�wsvO���	�T��;�PmB�js���LG��� auj���`�O�_Ɠ�Aٱm~Jy��~�`�FB���w�::ʍX�˭��
�R�+9bC($�e����P~=\�.�i~!̮�3D�ԓ4V��;)6��|�Y�q;N���eT�g��Z��_��7�622��ڳG��懨��:��/PJ#?���F+:6�������]
���Ͼ���xbf��ʅ�P���,k���RW���^!e^B���� x2r��0�a��q�ʖ!@Zv��_�� _ꒊC�� U 5V��Ci�h�8�쀟*���5�Mrc[�3�o&Cj�˶��hz�7����'q�O>��BI},������H�d�x[�����Y�����$��Q �#�72�X8�:%1���5���
�)�mT��c����?!	6~�]��8�@k�hC��UO���xCWd�'������<�J?qO^&���,ۤDI(�5Z\h���R���j7s� ��Ϳ��o��\+p
!��w�6� 5����������|����Aޡ����>���> ���EcFza���w�d�#]ˉk��z-���p8�La�b��Q���[ʕs�e�n����bj��H
;�z-`��c�P��]:��7���D(���UQ����Ւw�B��'Ə���L�	�O�d�M�����WYf@�9�ͻ�y>�630-�<�g��������$��]���"	q(֮���w		�u�WJ@�f�|M¨*��/I��
�7{�r� ���r�6�v�#x�Ydqc�FR��b��k�e�N�NU���j 颏��ePU ۙ|�����[�R~ �FM�9�Ǳ��G�D�cN�ܴ��r���E�'�ⴧ���۲�V2k�*.Mj�R]�׬���#���٭~o`��uvX��|��g~'?@������/U"#%��)I+M���.��J��UQ��O���)`�*Q{[�	��Q�#jG���kz�&���`�cJ�?{�W>M�A��D��F��
�k��, p0�_��i��Gށ�)�&M����^D���8�\���5{��| l����:���I�I1k��\ #���:���*ZM��+��@�"k�A���g����.���~�]jA���F��y>���oP���ݶ��{���=��g~��S"�d|��:ޒ��1.~�hc�`�ԗ��ql�F�l�u� !����kBZ���1�@p��z�(h�������.�۟��`����K�"M���
J����)~���Nfsˊ[5�l���]�LG)�y/^μ1l	��l�bW
Dr�$��Ř�c��q 	~'Շ]#�l�u����=��Fq�b�Pح)��p��^��w:e�I�e��({���#P��M����Q��
��b^�o��+��6x]X��:������:4(��� a��l�s/#�S����f����0p�5����[;n� If�I�/?�J��vw�~�K�W��豶H�i�	%�<f�E?��p�>�nQǕqK�xz���؄V<$�2!� �����4	k����E�8M�B"��+mE}tw8��^ң�Zs*��!�jG���<�%RZ�
$�_��fG��Bj7��ϫH	NF�l��&��DF�&�����3_3�>�w��}�q��b@��N;+��?���
N�7Ѕ���lGc�������ȋ�p�2��{Wc�ܪ���u��/Ì��'�lc�z\��A����Gu,��pm�!� ��d��k�8�PJ�(ǩd�[J���9H�ܰ�4�����b:�D����}�tl��a���+G���@��a�9��jp5P��������t����W�oO���۪.<C������]}��jޜ?�����'�n�"'�y*(i;��e�g����G��d�]m��%�ۖ�H$]-0���~m~.0�H���_qu>@����J����=�=��B X�q���#o�cj��ﭡ�5�Nk�i��ٶ�^�Er�Or����GE�!��܊���j)>B�q�-���Zn�;�#�:�J[���[�>q	hMD��GT�3�4�I��UEc���e���Ѐ��Ver3.OS���#H���w]A1�{�䏑����y~O��4q{|;6�֧�񦢠?����1�SvQ��-d����N	t�~7������aO� �6�B%ڏ��ΈrA{g��q`v�O������R�_��Lc9�*��	A���,��H ��ISI�!|«�ZN��i�|[�C8ˢ��T��`�b2�\PC�G{�k�\m�#��ն�����Ɔ�b0V�[a�W�fVe���_��Ǡ��h��6>��������0Cp `I�r1�!��}&�q�M�ճ�y��e]���d�qǩ��ݟު��h�FBo%�>U�0>'&[�38��G�p�d9v�gt�?�# pFW2brC+.^��	A�cA-�!��@Ta4�r5��)��ŤX�Ǯ�f����c`[���ﳢ#d�]��p;	�f!��K�"C>>���'��:��ut����Qh,��Yy�	>WH8^:P���P��TH`�[�3�Q�n��q��ޏ��Vq���0�=�<x� t�Vl��F}��n�L�cu��"t�$��UV�?�*O�N���"˾h;���<9�tuw�T�v:u�vM�D`�3�)d1�_c7���F�-���$e B�:�f�d�z�YGA��8��O�6N�D����g���F@�2=�n�jڤ�[��.#*@$M~K�[�`�F���f���Z1��uyXvm0u`%8��[D3�:�S���T��s:�y�@�P1� �p�&!� ���)��y/0ϼ�:.2#h��̂�:@������Ǝ��3�k��g[{�|��Ň;�>��)�	-��N����ID���?j��vR����,�3�zC�V͢��ӫ���e<ϴ�R*[�vy�XUK�aR~��%�eX	 8��v�Z�p*�Z��[X�W&��*�K"�J���ѵ�l�A9���ˈ㝃�����$�H�&�������K|������憵6��u~	�Z�tD�[+�w��W�b%#��~�!��G^h�|��˄M4�hR�e���HJ�s ������3_�(� ��#�SS��0��h��0���q��i>,n�ƘR�V�d��z���t��0�fs�,����L�&�_�h�p��ֻ�z#~b3z/u�pұUi�0ʊ���0���e��5L�/Z�(
������5x]�VG�(3�1y�cӼo$��	_I� (m�с���%U{IT)���$k������u��`C�w������q�{I��`� �/�c1V�$2��� �Z��"	�L�
�ei�.�ta��{z�y�`��+��G!9�tk��Aj6#ҁ���<�=�YԀZ��X��hA�1N���I