��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�`0���:��d�Z.i&�T�x�����^=g���&ㄱ/Smhg��0W���S��/���@�]��X�����d�k�6�F��Tm��Ҭ<���j�N����60�d�g	����0���֟a"��'�7�S�W;�s�v)�X���@�א���>�IcL$��4^ͭn�'��>�ĝm�Ⱥ���TF �$}�c�肇Z��%~��k�Cr%� �1�9ʲ�*�������x~�{�;A&]���&lQRVo���p��(OE��OI��!��C7���]�@�NT�	���4&ʏ{$��%Z�M�ݣw}[c��3B4y�w��V�l�F!븲 d,�k:DK�
"���| �ʿ!e,�ɗu*�5��3�y
��^�~��"�E%����8�����2�����\�%�wk�
dY~������2�AP��}7|�}@o�b
��"�n�Wq�����l݊�?��b�7BW�u��m� .�]ej��0�x���!N�bE� qm��#�6Eϵm/h���n�
7������6O��w��w���)Tހ�i6�1����8;Q��z(�?��A���^������6���G�	�P�2�����Ǡ�qֺ[�M��"OcB���*���gW#�4�˜�I�͋�j��ؓ*+Tfe�0>
Q~�9�@X
��K���'��=��������WU�$'`�R[���K��=K�v�T��!�.7 ���,G��֌`n�J�+<?����xw{C���JaɅd����VeH �� x���ڷ�-僭P7^�S�w������6�/�F�tR��Hj�:ho����'��F�;-�\���W����B\�OGp$�t�ߵP|��B
U��kn�[+�̒�P�v��-�U]������%X.�An����D��܅C��g�=5wW�۷�Wr*��2U���n��ː����W����M��=ŭ����UQ[`��2�����֑&Cs<�Q۳~ũ�<�Z�䍀Z�����f���(���z�	�t���mo�ӣ
��Q� ���}	�^G���,ܿ��s��ͽ���:�)->�Oyܜ��ÉW��]�X��h�����/�c)N�YT�2��E݅��ܬl;v� >�<P�Agӳ�>x�a�[�'�֤���N�T�h�zH�̰x&�6}6KO=����0���fv��A}�EA�s9��]ő��q�i0�DC��xWe	h}$j��%c���R) 9Z�(?�=\�R��@� Q^E�'z0K�$5�],8}t+]����H�n��
B���7��a̯@��$�q	6��_���%u=��ל$��'�Huc�����pv�a�S6�Ү$[�3�8}�$$� s��r��8۫!��a���ȴo�X�|�H����wo����]R�2��@�mH�&d��%>�j3����l+P;��ܭ�1� T��`��d"��@�<�-�M��;|z��-��PR�.A�q
�� ]���O8������e���ɍb�ڽ ,�e.�K���;O�7���vp��~��ŧ����ERb&ظZ�9�i[����g5]�J��aSE�ʥ��/��Y��u�Ç��!G�x��y��2H�b�i>���h"8c:�bs��4��G{��{;������PD�撃��:Ӂw����&��狅�>�i��]�7��$D���ͧ)����@�����������C������G_�3H_[����Γu�(���=W�i�����|#�ۼE��ި�b~k"� ��(	�V��b�c֡!B�h,��[����7��]�oA[(N8���
�$ "�:���f�ٵ�b�T"�B�� @�����  F���J(�S��p��h�����JN��4���̣FbbI-YPO)Ň�e�5Qv����x+t@�Xj6ï�7��������Gφl�M(��NݿX�jys�p��
�\���.�*�y��07';H��A-RY(dB]�������,H��)�"��%F��A>	bR����U������BM���W3���Ĺ�������17�k���q������G����y��r�n�C��Qe��[��H����33�����,v��r��E[r)>x����e��0�����q�OU�M���Ж��\[mH$\Td�/��kN���?YE��'+��d��_NPS�{��zY���2���[<a���'X��qOa��1J����n$�h,������{���!��{N���S2�JĄ0�ñQ`B�!�[�O�23r���Bܷu�U鐆��T�����)�\�k�s�^y�[]%+j�;�P̖�1�+*���D��tۤ�����7o�r�:w����aԴ��P*/f�bu����F�dޓ/7�0���~��%�vC��u�h\�ې?=:)��1�u�c�>D�7:ǽ���qv"�A��=P�T���Ζ��qo3reVnHiq�����!���o2�֟�i�ӞJrǚ���ҽF�K��Ah�;Nx��D�)A��g�:�:^ҭ:�Ĳ!SY�g�}�`W�u�&{����D���b� ��r�ae�;���P�"bm�jk�r�;,�U�M����&�{�����$��Y�x�i����-��m{�@�Clr��,�:���>�x�tZ��g,Q��}=I�|.�fWi�ς�i�	9�mb�Os�~	*x�*=Mʠ�l�M������i�3�L�`Qs�iE��P͕�'nqv����7b�Q"h�d� �B���� �4&�vO	�yȻ=w
�
�f��G��0�@h1i�}D�Db��G�׆��d��~q@N�HÍ�y�M��I�U��(���.>��L�� ����ˀ�Wp�m*���ހ>p�	����.�$�JLhZԜq����kb������ֵw�ȏ���:Id��G�3�\uYMm���^cf P[:�/�R�Ѱ&!�H��9��$����.��=0a���{�*�3���;��)Au5���k�}߻
G:�⛩�m�*L�$)�d3���}s�FTW�$��5�̬�!;�f�!S�KC�׊=������B���^>~�qN��v�d3f���.Ƥ��H؊G�o�OPbJP�=R|x�Q؎!Z�._��c%q��?W��}飴�h�,Qשnz�p���ܑk�<�۵�܅��?�V�/������^qF'Y��O6G��>K+w���*V�O��/���d���;+��� ��؇t��@��W����� p|Cc�97��%<��"nEuS����x|��tC���@�
�N��*G.N�"�̱�G!T����{���H��6��>�,�����_ɹ���K���� �B��#�h2^o;pH�x��Ο*v�]����?߷�y�Rj����2(�|%����+k�eh� X>U�����BNQ#�a�֕U?�����@� }O�}�� ���6��D4�9ԛQl*瓼jn)ۂqѿ�~IiG+��qMZ���2L���\Oo�+L��#@��~�r�z����ƚ��2b0�B��E7�:{j�.�
ŗ��[��k?���w�d���54�w�T�7�Q>#���E��u�ߖ׊^�OܺJ�< ��<ѝγ���̗F]R��#���Y��X~ж�-��`&��W'*�4$�4h����鰼�䯇t���M�W䇴t�ݣ�\�ՙg�j�z��G�j�F���y�ˊ��G��P ��	�>B�Hnwū�[͙�1��gX<��uc�mF�?�ZQR]���f�X�׾	7H��*�4d5�=�'��C�~�tw�K��>l������f�IK�԰����K4�xj�q�ժ�-��^C<a\��W�l��#�D�=^0��J�4-G���S��Z�\���[!���w�=�GuCM��A���8��	���I��~���#q�;g�[��==`l��q ��=p��Rs�9���OJ�Yp�C�N�ډ+A�@Q��:�٨���Ct�"P��}پ�up���
dXP���G�3I:85�:Z;;~�qN�c&5�BHPY��G(W��+Ȩ#��O��7P�M
i���3�-����$f�,��v~'��Y�*��Z���7��*"d��ͩzQ	7Gd;�g��:t�ޣ8W���.��	p�y�¾@}_y��n��_�������ݍ V��֕���(�63)q=�96l�@��8^'��%�0lЂ�本�]*z���*�	��b��[-1��D���$�v�@�_	�K��Im�hrۘ���������;D҈.�D�	�֊x}$��ݛ7ߟF�h0a�U��**���	���Ih	�a���"�m�/C�w<���$�
�&�y��7؜4�������W ����w���b��#{�]�5�\Q��	%�5�cQ,a |t�G��3��\�ə��D!Wd��-,��ג��_�7<S��z_�E���o�ޕ�uR
3tt���᯼akr�"���㰧�P��?S�E��½�<G���p:���V.fi�X��/�u�t���Sۢ��7�h������( �Y�ᓅQ��f��~��eme�à�(yȕfZx�
a�2}:+�+�`8/P�m�
݅B:5���dM������f_��'����Ġ�+��1�����㷏�=�<*���΁�B�7�L�Ş����-q�ře�{��/ҁ�JV��Y����f��2�A�@J�|�E�ܬ�Jt�P+�zLI %���Oz�6i���dL2���qau\��)L�`E����rt�2Z�.����u�T��'i-z�`�� �fr+e����^ݗ�_'%�|�lg4�9v�z$�{��V�/r���[�WA��ڴB���u|;�|�r���-�����'"�)�k ��+���\_�'�P	V8%}P�]����|��&1�=U��H�b;����+�a~�<��I%���݃1hW�{)�$k�m�L�����"��ʐ�GH�
�{���Z	�����H����&��Im26��Z�0lj�M~�߶C<��#�|ӥ�-y��T
�'=�w?bڂ���k#1���1��*�5�<3��`�ޫ��Y1�p\���/٥��Z�ƿk����X�O�]=Ts<#$4�5^��@��Ud>���0���&�?Un��s�}��� Gg{J=/���Ǔ�q��{�t��V^浦	.5)+��RWv��L���CqZ=�a�B�6��m�&�0$?sI�^Iמ��;��[�2�,��.g����A9��> ��I�ݬ���a�()Q��¯��liz��d��]��jCz�2�{o�N�)�羁�ߋ�����z)D�`2����Rџ�4�@S���[�~=�g��"T� ������^KKA� nQ���;4���V��=�H�lj��$p��R�O���}L3�038�8�~ڙ��oS�#�D��ϴ1iV:, �[y���m�zX��	����D���9�Py���,�7�\.S��o���Ѧת��b���c���"�כ�h����$	�Apw��Uf�"�.��?��������?�	&Ϊہ�ce���2�1x��"��F�t �t@����)Q�%cV���֥�Նpe���0��[�7щ�7i��WҘi+Lf����3�����SY���Za��"Ds�O2�ؓ��D?��pz�:x�ի�m�H��V^/�
V8�搮X���S9�R���r��v��sHnf��#�.��^q�e7zsAW/�C�mW�r�r�ip5rya�-(�$ۀ-�]�t{���[\����®kb��V��+�r��/!��I}�6eӣ�D�
������F\�������[څ��X7h���:^�5��4\���ӆ4X%R�
��J'P�5=@h��&2��Z�G
.�6��y�1���<����,������N3^#�F�c�t����5Fu!�k�����3RmQ'��Q��
�V4-D���TA��,�6w��H�-��(6��j!�5t{���@&�/��0�Wxs����5Ef��1{Tg&��X\�ָu�5���(.n]y�v`�c;.�'��'ܑ,�{� ݒSٹ��[��ٹ�d���tr�p�D���#��i����ـ��(�[���"�Iʜ� �:�8ƫ��m��#V�T�WS�D��Rɴ?V�[�Ge�������T�%���h1��7`;��'냈�3�ĳ��W9�qw�U�E�H��]��/�
�)�������H��I3i����U�r���Z\��:�X;�"��"�WWθ����uElhyYr+��v�.�9�����OV���Y�����/	�P#��i,�̑IB�X1z��9��X�{�38R�/6��vB������~1$E�$����5�P�k���r�$>�#\I���q
ܩ�R���K���2����6Dh�v�{��8�4���Y��eMڹN��}��A�Ap/E��E0�;͡������*�g��t��#��@�(~2.� �)e\��L�*M{"�y��}����Z�D�F̰�/��d�Z��������c��q�&��K�����i~�i��
m�h���T��o�t$&��X��;&М�i�	T�L@	��)S��CA� jx���*���u���_}hkҢ�#3{�r?���� ��*���R��lbj��ʝ].u���}���|�h�Ƅbk��@�.\�
���{�5��14	��Q�%�z7��~�=	�T�_#���/�q�ޣ��ANT��iʁ�r�����JV��#E'F�
����ʱ��P9v���C���6*��a�(y�o�_I�un��[pr����I���fҔ��ɑxZ*�ȟ�"��Y�<��`��V�5�6UIh�S	�ﵿ���g�-�g5��U��}֖�i��r|P*t��}���8�x:� ڱ�|[�9Q}���E����G-�/�G��\��SK�&��=�H�r_t�:���";
Z)Af�N�q/�0�� ��8��s9�:ZK�a{K��i�_�����X|�?[k�K���h��x��?H	��hf?;�U�LɎP�@�u��H�DG�xvc��M#������Η��J�������ڜ({|Q��z�+�_N�cV��H�ٴL	sW���.%�A%�݆��~���"�u�lD�̏=DEw���y�'.�'*����07y�)��o��B@oyK)d��{1	�a��]�ݱ׭���o!�R�MK�~B���O�D�`h˵�8��"[���� ?f&rյ���-���4�ִ��ݶ_5��.b(����<8kЎ���3�*�!�з��0��אE[8T�ټ;>��0����y�jsc݇�7 �ū��u|H���Tc�O����Kp�.@��Ӥ�*SJ��Wq&�b�>�W�a>27�����F</pJd����>���["s�����4�A �`����p<G��:��Y�m3��'����=~�����*���,�o����ζ�%/v�����Q�\��`�z�$�$�ضP鸜S?Y�=����c	� N{���}�/�eEݷ�� V�b���t� E� ���A�b}:8�VM��aK���
�D���ݸ���7:���"�@�@YX���!V�xH���� �����o#���M!�blEX������$)�ݺ�jb 5	��8\1�P�E^ M�=iC��`8��<�sy'U��i�L�P�E� j@�