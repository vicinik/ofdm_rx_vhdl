-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VL6/eV1YVXgXicXWQ3XNxLwWEkSWIceXsH8HUT+YTwgIUUgmmHLn0aeRx+x4mCiIRo59/7Z18xCt
nx1e17Mhr8dDjrmtbWG3MTWcyutu5aaWm6GHJZ5aOQyFP1IqSDyBxBnOj1Yswt3ZxroZdvoOrnGn
g6wwCpbY/U/CTtlSj9wBq0IDAnfUL+eRkGkMYBPSU+VQIk2sIIgiqZR2jrNOalwVJMwVN6f4Ab/i
HgfYaTNZNguC4kQowo5rkACgZVPW3xZsC39OiS50fLp2l0T1L9gV7rqHP+uOL+BlTIQdHEz0HUiN
4c5Z6zYKWd4wl/rYxdE8SjuwfQV7hX/rGnT1ZA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3360)
`protect data_block
D0n6o1lSzpNXGU52J3KeXeUGIWjrztSOqmobgspQ1D2XKhfwroLpy8bh6+LNMNCSFsOYv4l5cHOY
YJedQi1EraMEOrJURChvX5V5Pqg2RoyLGnO96Lo/UWWF+2dsELQGbN6uC7kC3d0D457ez4YHP7Ym
Pf3mZUkuK/V8oc3iVgJIupntd/26iE3UZzugeEuoXZJOc2t9M8XtxO8vHRQvqwjkzyF+S/hXqdge
FHKJYmyRvq4jIQ4/QhusAObYKAa3Nk5UOMFs1J3p0PFbgu9GQbbJN/BI55AOt8pAWagDIJmeNXpD
oYcBVnF7b1OkJ/74wmG7UUT+V1Ns3JHpMNWeiWJf5KOtIoPeJUp+FQpmXd1O5vCvsIHDoNBam/za
X3cay7mMe2/uMJXfGkUvis3eOQ0ZQcsyEllTQVYu5bkqZ4XHiNkrLLFGO5J/qVyzHGN+DbiDgbqx
5kcIxUb1ySCuSh3/cSyzPjUERvmLbquRa2EOhVi2AtUzTrppbz/AdWY99N95/dJvtEf7t+nS1VWS
IKjtuBpuzbiAij9zTlfM/4X8EvJlqBsQnMaOoWMp3+KaHIyQ1OzqRwQPMqB4nlQpy9TZ1vRPsgMC
t7e8w4SI6SRYiJ7t6yVSaRwSKqV+fBj6vcGBOimCk/92EkJ3dwZ9IB8VgMb3LJo7xa72STOVZ3B/
Qj08ylu7E1ochA4TsdN4/THyGvq7HIB5K1O4YCta//LJ80baqQz59jtsLB2bgJC3s+hQBCoAhjri
IWHkUivp9sEvUbTSW+2rrgLq3iM/qIeVL9y/xaboipYFJILJX5mSoo+jZQVXCBy4Z4AaVWz1NMW6
l4eHVH1v24wHUJ7hk8H78f+LVxHJqAWO9bxHW99eKzNujm46CpgjPlo3/7S8jdegh77lfUyWaUtX
RFroXzuElF8BitwcFEPtwMvXJ6cStVRZksruT5ZTjOhHleN4d2FoVN0fR8+oJQR5y9yzuoGejPsH
n4nyJWrkgnWZBU2JvJAWoop11ju/Kzyx1Hn8zMLCGKFhDvjmu91P8Rzz4sXGiDPP0huny1bk3KvM
lVsuS9sJKwz8Q1sZFRztoddzjcJSD27WzMN0/aHBjYNkzrydcOSbV55QVVPrBxxZhD6gSi6ZAAqn
aUMBX0ZJsTwSBxqOcZxsoloK1OasEuAslzsruyYXkcXnNwE+Cfv3AivU1sN7+ZVEVrfqPyinHmBJ
AAIgp/ofkDhvikQUfCADEehYlMmxkf7OCd4qK1wfgQYU818qO1fgRCeaT9UZfQGbo/s8f0EHAFIw
m4aOqUYsp1RmZxFiEAddNAz3cod4oKQWHyYjglEn0wCgd+N71RsE0rMCm7dvxb+dMnVuCl1iZzvf
6pWn/Oa++CA3GFrQlMpZx1jXOWMcxIqdtqQpQNrMmOKSJX64cyF28Pa1SLhCREpqr5ampBZ6z5bI
1vO43BGEmgYBG2JNeaDB2AjaktmAgkWgeVKKe6rvVJEvOnxYK/1kulniNhUfrYPxZXaI8ED7As/y
YYHIPr5qK/8uIqGKKTshREO8woNd4A7Knb5BPaxnk+c8wXm7/zed37HsLYB2l8bKLVC3LZhw5lpv
v8WMfUPNByypvQ9LwuRO5Q7Y8lXBmMBnCwDz9dRrXzgZrUvVwGPQ4Czrzdz4gqzCzhWrYCrex6h2
FYqdTlUt5aG9O1iJiznh1tTotwMsTMB7DhhxxY+v2smUVBKKXWopyIzjUa5n1eNbSlGT77LoAGTV
YQmgKwoRD9xz+EQRUJv0Lovzl8Y8xJj25O5TnxbHZpMwK+tK9Xj8gIrINpL8SYND34bbCrkqbpM0
4ukiani6AgrmRcrlsK2STlYn1Kjpc2EcCc25E1XPPKLgeoSZ4pojprMAcmPAr5Lp5E15A216kH0T
LxeIsGMYEpxunFm5fWV3u+3EjNK5WBE4Ic+Zfw2PcZYy+LFel3MNXM7sAkp3J084PM714SSk8Ygx
CSsLjdglwOk17WiIdV/DhvLW/pbBm+Pddl2E0w+VBz4GDo5tZEtriUuXKB+xyKbRTJwTu5F5sCLC
PVWBDF9bLEuADaoXwTdClYg/zzT88rjmCsZu/5nDKryLa+qfUSVRFvxJ1kftQG/QaKvv8b0vZld7
9tJ2QDsns47yfpJPaFYQaez++dHFmkYVYIvtjLBcVAwTgugGdc94+/PVOiVzPf0t+cXXAbLIybU6
SktB/7Erqx2smVLZ4pZIj8b4VtbVGSTO2X98nPgLnUjMfxBATqlcomDaDN/obVAJ/JD0hWxL4BM6
5+WNVouSS8Yt4MpSyQqYhaKdp3fLWVImwDW20quxDF0/uPmCQENaQnBJ/Crd/4El9zCQa59HiJLU
rAEq8AvcVEST+sbQxZ0I4IGp7ojycN2tiFFArxs6K73neLblXTyJifnrixbVKKGMXXIcVY1bKsCk
A2kuKVkMsC1X502ZTaTtVHsDPefxS1yJQ31Vu57Mv9PxmVVrlXP86o0rAju8YeRg6EBOHBvH/J0V
ph+bghz5rh3MnzE185de80itVQ6KZfxFiyGV/NQyZr0CJjvCIyscFDod0mJRvIXglW8yB8hoRkq0
HoaGG9Y/wdZstnQwP/K9kgv30kxsveSbYX9LG06LqQbKRpONxLSC5NO73rVFHQHB1VwlMl2bN+1F
9iPfYbArOcWHp+YwFRbHQrpykT0g7kj8UaxUvdKb/WMohWNOn66laxvyvW0mXfLvfTDywkPxuGmh
vzeZp89s4D7vErBYsuFnwJaaEAel8ePTj8y4QADH+NPrkA08Fl+tHdoL3BLbGIf4ifCMaDIfRi9C
3AfzPjsykM3tI9x0iWSifB1imqYPxtmDdp1Frw13Odzc7lt39T4DxPJT5IYBR/+15Q/Wt1ctMiqN
eDNWYNRBogMWyugcjg++vX4p/IMi0UAKn9XKXuxmHL785SC4SWSEvMgs1FLHMiJnG04FIIg+1yD+
Bbn4UvO3sAyf4wPljXeV2CN9z+2g/FiIiuuVKBrtFI3tCj03i5zY/zktY5cPhxJdF3mdDVfo1lW7
KjbbhBSZfadjWmg7tEYFpb7XCm2RL7c/AXHSZAw/yY7zPkutcV5VhiTeEYXRERxPnMZt2R66hKaN
VnJOAzzu95EUir3QtviehH9DodayJ5JQMqbBUuJkbepf5pYteN5KDGFDiYuuCAq/TJNzHD8izQ+S
hvtHx92IP6zm86ONsrTjylnQm9l6/07pMbcCWrw352fDV+IJWwDfMbIGG7Wh35URQUz6JtBQunvd
JBT8LqN4RVSjbzHmDEHVotLPveYi2Pz+xWvddZTt8xdV+uUb8SwE9InnxbcJ4VFyk13XKSkMo9FC
OIDkW/iTETlKzJcwrKVad9xqSofD42KAdnzN4PLS3cyIgMUpYEiWhgtTyEVgVPa1iAOMRD8IlMOc
rA2h6D6OV6oM5u1gWMPa2gpqh8yJsGSjBLU4Ng4KIUukyBH+qN6UsWVFNHcf/i6sMZ3TwfeBuNV2
XgNDMss9PGrwg8pWWEJDXp7Lfbik6/2cPMNcqyxWBMnU8mJynvn1ktQt3x31QH3G/ZfxQAG9uql3
1+iGRNPKIZOx4CyqF4oliRMgurhBqbPBF6p4EEtKTPHjYnzsD+hxUqv/mD+gFs43PNfCMv1vY82f
aOEOBagPtYgT1t6BO78ImaO4IU+9JrfluKBwe52xn65MpYfDeVUc11QGOUkfV3Vt0Pz1IIVYWyFZ
GraOc9rbfoc7A+VDeNtNXNBUERyq9ld6pBu0qw/i8t2cF1v5nUolUfmee85kqF31l05M9IIr583w
uHtNBWSjzgYUuayX9kM2fI/R5cztUXeYzr/P12J9+aWy8Ybm7XsIHlolUuvwg5hbwb6J0P0gRxMS
tXWpmAqc+neTa94RuTgrPyRz2DOFUkVv/2tAvh2kc5QF0bekTIvagNmuZcNupJsGIp+SeCkcUF9n
6qgBZXYdTie3zfqaoR45i6aQitn0aEtXy9wB7n6ZoVCrKlc8Y2ztB5XWyt/vujKjCqoFTYgjWGri
QSwnY2n6WUZC6eOIhbn8D+cbmGBhznUpZpS3TEiEGJZmQsRtdIylIO3GQS8rctFQeR1K4uUuv3jq
kEgIWTALFqi99xux4p47+e9NgFiFWPW/vfbd9qnVsT5j9Iu2ZTz+E28iboC2Ge5e37CaGZjcZ1y4
ny41c8u3l34e7tQpLFa7RWpSMtcN8wUbluWnyde/V4qSzrVzSq4mVjWlvBagRDSTDRbuniaVLipM
YVlo8KCd6wVFr0qMSvY7upERfTkmN1+ENNjNih5XGd43HD/BwpVIgiQDpS2t/sE3e5h+6H0Rb1Nr
zHcakXXFWKByjOjTZPazDo+cMKt1UAeOGzmnJ7B9yj+6ehcCwo3OzEuagZEusg5op8ZCXJk6EKni
UtW2gewnn3Oz/HvZm/94IH6+gJUiULWcbLae9FTl4eBmPs3xuUgH1ihc7bx9Pwp4xYRQJbT3
`protect end_protected
