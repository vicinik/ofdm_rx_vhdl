architecture Rtl of FineAlignment is
begin

end architecture;