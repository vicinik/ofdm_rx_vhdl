��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��h+Kg�#���_�Y�� ����U�#$/�&�J�5iHתr*?en��?���������b=�Q����9/����N���V$����W�r�s䅮q�N���p�x�,a�-1�5��
_����(���vORv�����M�}b9B�6��1�S�Y��,T�u� M��������^m�om� ���kf1;��0ɟ�]�л3��B��'PV0� N�p�U�}>x�K0�[�0�Q�WJ��P�N/uml"=З|�@��]�w�aapc\�+��:��ڬZ�N�i������1\/���ۅVk.(�f�pb���ǵ����<������:;v��|�&�a.X�3V$B�q ��,l�d�@�����1+�3m���&6�2�
�YQ��te��y�!l�:��}$/�k�^R�}N�b�0�*�������O{=p�-��W�g>bf��8�Es?�s_6�� ���P�#��E�ӑ�L*c�,����'�ѮGON�����)�m�|���׉�Ja�����k�R��n|�5[}7Lb+y�fӸ��J��	T�e�\���_SKq&ꓗ���ρ�m��u;�:�~�"��H�	������j\m䦖��}5ur%�s�Ңŝ��5F-���B�	ow!~W��Ätx��x�6h�Bc�"@.�QU���(/���槽�1:��ŜD\2�O���wG�"	��iGE'ѭ�����?R���ų�r�K��Q���uG�m��J���O~u�;�ւ�5>lo7]�]��zd��V����#�Hx�'�p ��m�M��Q$�\ۘÅ��5������B�v��=������0�s�7�/�'��X� ��nП\�ʣ�b��R�eHp�����!�*�5n��gu����ޭ�M(S�͓Y�v^����^/Oѓ�j���u\��F��Qn��طP)M.����o��R�=��d��H@�u��#�e��d�gh`���^Qz�h�j�;���A��&v��7d߳W��9�W���;��:����ը_k�vD�����K�
 ~%J1�ဇ�27/�*o�ʰ�H�WV~g��+�^@�àN���ud���K
}�i�bn��o��W�-Ц@�Ca#&t~�7�Á|����8(}�*a�U�B�)*�0�=2�,9��9l�����']U< ���T|����p&���
��'4�H���]n����߬��K
5䌵��Of�"�%��9��q�?E��o8Z	��M��)��v��kd�w�̀��d��)`<��%�DKS9��0���-i��F�	m��eЌ3��������ײF�^�����%}�e0^�s�Fk���<1"7�s����z��8w̡�H�������&%���)�_&�@\z%o%�E {uy��`վZ�'#�r7�:�"]����s�:]6K.��O�$*��/:$�^4>�Ak/�r���6�=x���/A^���'����ж0ӊGMԺ����ًj��0��0����7K_�����!K��}^&@d��^T½(SS�r�u ��I[ R�}��ϒi��q�eY�P�QB��̽�<�&�iq��B�~
�
�3�mzj�`�������Bxaj�>e�r y���O��̮-���$;'�7z�잃0���J�Q�u���1�H���s�h�B��'(��!�n�h�ٜ�HC�v�U�sg>�[ӏ�b&zwD(s JUg�;?g�s\D��T���9FWa ��^B�����
f�Eh��ؾ��b&�FS����K��K�=�K�)�2�}�.�l"��7�[�~����IР�V�9u� P}��% L_O9��ֽ�1��I��v�e�kE�c���n�OF���OA��V�ƘO��HT߽=���,��XOx����s�he�ʂyW��6
���:��W�Z�ڣ��g�$�(<4k���c����}��<*ʈ�(A�9�`5��,�ݜInzS�L���s��↣n% ���㇁����z�ӶC!WP��p�r#�6A��\w�K�����^�]3g̜9��pά'{���9P�)�hwYaZ�E
i�Z��'_�yS��Q�.�Ej����wu>�U�����L��?4���G-O62���X;{/�V
@���Ϊ1+?�b7��L�}b��[��]Aи��:֮��9u��F0)�f�cC�+hɲ�4�g�|�3�A����)`<}9���m�Y˴^Uɒ��'qn���Dn�3adTxH=�FB\���!�� ��z^�'�w�&���\��ðvGևu�xz���I&D�'n7��(m��6�q�ys��3:�O�]=r�[/���$=�V��U��2Q�Fi�lH=!ܵ �w!��m�"ڬ�B�M�U��QqB�"i��	���?�6̛v���<��nP�|��>_!x0���؇3"��dΚ�,��C���_��B��鱻���\ +"�����̱��[n�����t�=H�ߛ_tH�b�	���y��Q6���^��G�{-Q�X����I�t�Y���y鹷U�WFa�w&�{8�����f~�qOY����.�:�|�٘��KS���M�¢lywD��*���0%"����ua,	�)�ٿPT&mA�m��n��k*gd���t�Q��|���g/����d�ѭ�d�F���l�B5��!*��7�b�M�tx�poHf����V��W�ֶވ��ޗ?����T_�����屡��F�!��1~o�n=�<<D�1�XeD���ǩ��h��.\o�Q�����Δk�W��j��!|����pſ��m"͎��/xHS���ݒp�6F0�tё��y��#��^��+��B���:���f��qc���rIJT'�`b{c#�(����N��YO{�J�3pt_��{�}����aG!��s���
Ɔ��mzJĀ�����]���%�xU��l۵x���o�(����o6�"\�܁��9E0�:S��^�M���H��Ja̤�P��O�[O_��Ng�
�Q�R�He���&1�Jפ���7}�8K�!��Ov=Ͳ1��m��#_�x$�e) ��{�,��5s��h�W	ņ�;[�ko�}�����R왧f+�s�Ni&:��`W��%�+��C�Dg\�$E��"�8w05��v���|�$r��Ϯ�����3�
a�2͡2�[ݻ&y]���=��4�� ���^�-7�#-�Ui)/#VTc4�k�*�E�"MEZP�$�����׈]�A��O����X����6$�L����+[��ڮ�s�ORr����P�V"�V�6�:����`AѝR�zi���^���Gy�)��{�kicm��YG�KF^j_��)�;�h<���BB*%�\�+� 0u����t��S(q���s�vo�%4X�jPxx����-�*�ɧ��vӍ�#�E�娅YD�NZs��r�e4q+t���F�v�z��z�J;���%o��U��.�� ��B:ub2�}[�D��N�o�v[��ik�J�����ފ���F��z��_rQ7q�c��0�k*TF��s^��e��'�� �S!��8�F3� ���n�'4����4�r^��va��H�7�E&ӥ$�]�K��T� ����Y�:�_7����r!����L��m���e��s2/�oF��j�բ�U��C+1ᒡ>�>�����z��w���E���u���I9�`TTuS�tD;LV͹%�O���Ԓ��_�ý�0:,��OB���[g�!��c*�i�Y��}���������6 88�t���RӞ�b��fp��=�^����*I�h��lq�pw���f�O\��:����/d�ONI� ��@Q��:�~�c�+�ک��|j��sxY��T�}�F�8CY6sΒE���ĿWy�}K�����a,�
����f�GYKkM�Zp_��QX��6/�L�<CQE�R����Ζ��evK�zI*n�iK4�b`���S���N�'H��Y�+��5u�/On��h5�tFdp���0dr%/�=�tc�����5��T�eT�s���4@#��Yc�5q��2�A��Z�{��'�K�<ėf9�%��Y���B.����U?:���[�-������:��K ������h�J��������*qe�.t�ޖ��cn�D�y��G���i�̽O�SѠ�d׎L���Z��@.Ĳx`߉ɥl׈QG�>�;.�մ^����\Y�8��ι�;ċ!���V����N(�!,;�Rj�n�ik���͖����&W�����F��RTB3z�t�2�1��É��d+�3��]�ֻ��m�s�-f�s[�^M�=hP~Mb��an&���_��<(�VL��q�Z�����n�[�Xyw]�h�U�udp٥��;*���N�4R���:��ٗ�,]@܋�ug�G��P��:�����;K�ـ+x��ˤ8��xd�o̬�z�Ā��f�C�8t�Sa~I]���(e�����E+i�h��̹���c��/+���'XN%���!���;���bC6�V�2�}��Otx��"�O*�|1p�ɢhʎ��=Ȭ�Af�Wy��erN'MΏ��\t-�"�0/��jݨ�N�e5קh<����wx�8�������@Q������ň�
B�zy\�ӡO8��U��Ȉ�G.�ux�[>�W�i��[+GN�� ��@q��f����[�d����M&�i�͝��UjIy��a��wd�A�H6��*7q�2�X8�����ōt�;Ev��Y$:~��W�="��@/��]Ģz^���^�{��r�;Mt�h���kN��3�'�=��b����[���G}Xp����|����Ƞ	�bZ(�f|���g�ޙ���eҋ0���&JI�b����VuM�q0֯�~ؒ"x\k��^�[��J&CNX���kڛ`�f�Z�v>P��O�"�M�Se����i�M�H7cj�]E�/�F��T��π*��3Zk��a8�� Z�����H�g�<���f�U.VvX�W�Nrs��)d��d)��U���;s����x > A�m)2�V��N�'���#瑹}���܄f��b����?iןg�6��킦aɜ�$�@��oㆆ}�n#�8q���-����l )-}�1ֆ^=�z�S�'���yζ������!ⰪC4���%
��	,��?JEM����i+!�7��9�������|�T�q+�~�m���ݺ&�)��A�(3UY��@$/	�Oۍa�@�KZ�¯l�R�޲�۽� �"�������w8��;��/Թ��fE�c���W����k��T���_���ۓ�����3Y,.��0�9}h8�t�]�y@�UWD��d�kL�"�֎��@5��BgU/�J�\��e�p`E�@;D��Џ�
�.Y��
M'k�C ���R!r�l���曍��W�)����A���E�)	��)�+浌V'�5_�7��L�M@��)��\�9�`�ʓ�_s��<@j��気k,�J�l7�G}S�k̳Q�k���v�8���kL�*��^�/��
Wh�P9�ﵿ�����]V g�W�P;�M.ϣ?����)��W��ME�T�7�|ټ'�20�J_���R[�}8Z�����4�W���Ϣz����tUyi�񼏺)0RA%�Jڜ�i�$���5h<��s	��Mݗ,��)���f����j��.���W�J�v�qTsv��|(�k���n{O9���*s�S@S�n�H�Q�9�c����  :3;P_|�=�3�}�:�+!�w�|uT �����oL�6�O	w1H��
׵oOx�+�ݓe�~Q�BJ{΂-�(�!��(��Ԥ�*�^��@��G?6x8_%����
��nQ<�lzpG�O�N��k1�Q�]65us��g�]Fp~�1*x3��F��tG�b l?�G@1�U�E�|@%��ORn#��G;�����8��<�!7=�h��5��Fޞ�A7Vj&��c��bO5�H0�\��%���[��-��ۗi��e՘�Q���V�i�^.ɹ�ơ����H
�a����R1|�;\��I������k��*��KJ&��zC�)At������`�pW%u�dT2�Dpa���:C�����s�o�v�6:[6�=��#�r�O��>	6+�*�(�yaoe������@�s#ު`D'��4Ѳ�\�&����w|䇷�I%?���MX�����7ZU� �5�_��|D���(��b���	\���mJ�}�t��#*��
����d���y��I+j^d5�.�/��k�p������i	���R��[���P�e�Ę&Mfg���,ӹi���S[��Q$%T(�&���y�I�%7@o�Y}r��F������W�R�[F�b5TD����UY�k�l�õT��m�����d�9\���R���Q�N*��<Ob�[�o��-{[C�
!7nڳҟ�R'f/-_*�P�yԥa�aސ�=6\q�:Tn5ɺw�����>�y;��/=e�ػ��'B�`@����NS{��pV�f���i��`�0����\�r��@� ����چ�n�A+���k�"�q���i�I����s{y�����ɡ�;�Pq���j��Uwvu���b;Νl��-����M$�;��q�c��,��.���eRJ\[�ܔ����W��^�F�Q�<#�����v_sl��e�X��1�	�\�?Z|јA(ak��u�P�����N1���&�Czs�7�c�s��Z��o.H揜��EPON����K�������i8���9�_�c�<I%� �O��awT�[y!����������~�i^
������NG���rb[_V��S[� `�6R�<f��Y�2%�!t�;O$�VG �m`@v�],���j,Q�#�A{'�]$���O'�D��9h�nzZ�i����aD����Դ��ߵ��NN��� �I�N�\	W�d ��nZ|l4K��aQm�%Yt-�tp����&���mD�7kb�*�[f�o�l(viRy��y��	,h���M��w�
�l����ܹڑ��oG���qk��L6��K)W���j'=�����e����EO��0��E�-g�1ЯP(4��M>R*��ћ��)�'�`�\Ol2WK��s�3]wv�nhxj���- �ᝰ3��b�?%�)�f�:�����jg��H���c�A�\�Ex����r���M��(�yL+�A��Z7íQ�+8!�Т%&U����?�c�� �Jm�Б��L�Fu`KqC���`�YR�<��a;|O:�F�C����ya�a�A♏iF0�;0xi^� ���	�l��U�{x����z��o Yj"�z�l�N�(C�hk��٨g�`+�����ea��P�F���3s�
l�!��uY�×n�zF�;�Z����.���J����.����p�w�\�G�uZ��r˦�|!˜ ���b�T�E�2#�m�PAf#�ƫ�M�@�N�)|I$K��P�P��yao��1��Ur�/���9"��K�zW�
��w�����{V�&(��>����B����H _�� ��@��X8�&�a��^<%�@��-qr��8J3��R�S9��H$y�G�n��8#��}j��(�s�I7j1�ۿ3� ��Ù�-�|{Qm�N#�꯹'����d��S(Q���p`��Q����/���8� I�ﰦ�>ןg�)r�`�l�t�Gϔp��2�㧺�6�e��yyI��Og���bc�'u�b;���@.P��C���)]��3ZwE��3�Ma$G�|u��q�ö�?�>Wd!�Y^��=���lqdV�\�c� '��`a$,q7ה�歞^[q��^�b�b�/)M���oo4)����a��VyL "]GI�VF4Z>�_�e�����>�*�)�j԰q6��r��r�N�f�>�N_�!� �O�]J�Өg���o�T1�Sn�;v*�ZO�s��b{)O����\PL���9�\Á?�H;{��\�ʆ�;8�@�:�G;��X���9�q�#M��1�U�0���;��)�#�;��[�n�;ƣ�x�B�u ھ:��~W�����w���(�j���$��Qߘkr���UYt;�!�d�e|�W׼N�J�]	S�q�h�䖭~.-]Pu��r9G��<����p�U�{8sJ���y��R8�e����5��\d��&\R�u�h�a���a[��u������8�"�Y;��iV�S�}#�W�5��hj,��ex�o�糾���!�����PDN����?�}� q\Da}��NFh��Vw[�ދ�o� �����7�LO0�����h��i��:V7�MO�2�&�ov-
�I�M��C����i�Q	MV��u'�z�}��Ssz,�\�t���4Q���Dr���h���O9F��Z:p�ȫ�����o~``j��##��C�j"n���$�f�����l@%f�O	��N��W��� ��^��������Z����Qce$��zK����:M(����r'��b�h�O�>�XL�e^\����x ��6-���|M�5+��ru�O��ظ�nz�v*���%N︇tY�3�k���δ�!+y��V-�r5uD "���]z�,
{|���laGB��
������p���5�#�1l\�!3�ӵJ%2�+������F.��!hк�T�jH���V�6&w�3�C����Z����6�\,ڀ�}�C��*�c;_�3X�'N��sx�%���{�-[�Tm�����yN;\mEt���7I��(��P��/4
#=&z�z�PL��r ���7��J�i�<��9Mϊ2p�]����tg�g��|t�V�kk��~4,ъO=����À������c�����ƞC����8U��4<1��j��A�[��I�7�r*Ư)�0[pH{A�����w�S�T�@ئ..���T��L��V� px��FG�DXsG�
u��`e$vQ�`P\>�P&q읇��AE.ٙ���ㅃ)���@/����F4^��1�w��EY��	�c}V"`���X���R��8�x#I��ڟ^�� G��so��i �*~�u��r�	v��1Z�?��Γ���'���$�#��v2et7�����^�\(CWio/�<|�߷�`mv;鏧�:2{htnk�}r��JB��t�'���h_/�ˮ!�q�Vy��x�a��_�stG3,|��/ v|�	�ct^~���i�z�|�����:��P�hVWK�{K0����̇�ޑCl��A�����w���ޭ1M�,��/�B7sJ��Om4�,�?�ĺ��CQ�~����77�I/ڟ��p�$�w�J�j|5��/ i���L��|���g�#�@�Cdg���i;:�:�1�~pq7Ng�>Z=U%�T�!�����0��HD ��jk7����+���b̞��x�=�/���)�~_A1�G����&��T�c>�9������F����U9�n����hŹ���y��Y�9���KNo�V�Ǝ�7 XnWNO6���+0E7����廽seG�=I�����%�>_|�m ����z'Ct��*X���}.�Lk�N�:�������)���r1<��P�siL����RS�:Z�^]%�4"�L�:�cs*����fLx`s?��x:|Oh�Fj�>��ܙ��CC�t��6b2��4R��J��Ma�Jɛ����(�c�C���DSQ�'���dW5�=!��jb妠��ӔSp�{����㒠�O��m���w�6�����4�'jdg�蝭Q��W��V5��I	�-���ަ��a�/n��	����Æ���g(Gn	���Qw%����Z�ݒ��g�А+����Oy��Gi�z�'p�b���.�R�(�5p���w��l��eU�f��4��7|:i�Gq��ŉb��nT�Y1COx	3���ih�X.��R:]A��/�N�� ��r�Q�D��le�[QB	͡ᮿ�&�ju�%�ֲ0fv�~�<����b#���4��d}�G,,���@fD���UW�p}f0��X� ��I0#O�QyĮ_=�pGe����u$��ǫ�|uX	{�H�;�尽m�����@�G��Ι|��S Ǵ��Ҭ���󒖼]l�h`���M����ۨ��6��M܁'"��?��K��f�
~��۟T8"��W;��!т���[V�[�wfC���c�<��v
��Id])��}���8$>�����ڞ�-��Ȥ|���r�����;XajqWۄd��e���Qez?�Y��lyT(��?ǃ�a.��`���Y&�Lc`�6�G�-�H
]�3c�E��M.>BC�X�n�߹,ԕ��5�Q�G;���g�R?�s����n�N�I4<�-�>�&=�)@GXWȬ�7�N��)>+�M݉�pe5#Jq��Y�V�+�S^fq�~#2�B�y;�2,�	q����j���Zpaϫ���&3�4}D��l�v~�陫���[�'��"[B=)� ���B63�5��uH��\�d�UG�k�|�� ����e;Ѻ� y7O��!I���l�U����7��8;L��r����vYz��3R��}WG�aH|�&��S��XP�4پ��T�n���z0�tr�i�%$[�Jgzb��HG��z�]0Ѹ�+��g�����Ԁ'��C��t� Q*�g���!k� ��D9�fRg��e�5�����Vj��y�u�*�d����{tNO1���u�x`�{�p�s=��|���z���0���*rO4\�*X|�|I��o�]nt�r��p���,�lz��e��y����"¯6���~ 㡆�V�����{�"�ƽ3ن�jjF����{�5��U���AX��|��{���'�}h��F�F(h{r'���Ċ���F���w��8���(�x�`%E�*���֜W��Bb<�������	��dT��ݏ�6����$}�-N�X΋c+*%��\�+2]���pN�3�:Տ���Ï���C�� |���xi	�a	��`��<��O�et1�ǃ��N��Y�
��!��\�	*�-gT�Š���~;3W�
Xij�����7wC�~Z�Vٳ�B����{6���D�
W�Ɛ�~Z^?/���V$<rbJ�R��|��5���G�\��pF�0��R�i�����k�W|$ �O�ױ*UQ��q��lщɥ����x���j��@&��ۆ��_�u�\��ٙ�R쿷Xr��x�N.:#��F�$����N��Tٽe?�tnN{��&H�*Ο%��d"��A��|�X�"�臄 ��jN�##�w̢x�'�9�����Bu�kFW77D�W|hV����a9��q7����f&�.�N��������V��
gc(;�A!��u4q#F�!�(!{���By#�:"!������.��9IG��5��@=h���B�?.|�溯���2�N�t�.\.��fh��f,��[
�~�H�����U�}�R��y3�����9��{��L���̐���j��3ku v[�V^���`�.Y��vV�^�0�hsJ7,>�F*!`���2[U��ī�#!��WD�{\�u�Gv4���S%h�������l�p�e!�PD���3�s��/h��?�%(�!p����]��^�|�4��s��gh���v�^`�L� �H��\1Ěp�������o>�KrB�V5拉��I��D]�?XF�m���_,���P�Br�K��(ˏ9
'��Vޘ�z�g��HhU���6<| xHn`�����k�et�k�~C�()�;��H�ɪ2��8pV3W��l���ؑ,Ak�c��O"E����g�{v���՟�*�]�^Q�% ?��f���@HQ�YB*)P�lf��S�8��|p_�믠�b��e�D:��(��y$����T~���G�k��#��� z���W�� ��]c�]4	Z��b�?�5���Qg.(�ͮ����i���nڎ�
 eM��E�LE���>u��B
�t�i�����1S]<�W�n�%��U2ˀ�F�%�'��֧� ��r)���o[�����Ќ�P*
&/k`���Z�>�r����=�G(2���)�Ɇ���A7<k��gVI�'���v31ؓtq�3G+4K@QUG٬�M�@:�h��	�gQ��H����hR�:�����"�\��#
{��M�|��ސ��&�],@Q�@��i�GU^�-��}��J�Dj�Z����[WH��I��q�9:q p~W����T��]ɥV(偘=�F�}+%OtؼWB��|�>����jekK���Yr=�T��x�M!�%����������aziu��o�A�l��`%��b�2�O���ϐ)�c�=����x��ct�YB�����[�[2�.¢Z�Y҈�-��Q�xNb�<�܂�Vף@�#��?�@�6������'WT���'��� ��u�7�1��͎�.�FZ�^�����c�l̏̃
�n7�z�VY���x$"��0#\=8C���O��5Z'�.Zw�K�3���^�!����g�4X|zv���qrI�\��c�̫���(˅���N�t��tlQ)��ޙC�7��'7�}�'��D]�W�z�oe�nR6C�Am��,$S��ka2�"�<v���~�����]@0�qF\�>6�+��id赈�c@*J�]ҙ�I܀��yvGg;{v����h��(񬩢j
X�"�Q�>2���K{n�S#K&T�o�=����=��ZP��`�3�� S ,K Bm�7-Xĕ�MeZ�gvr��We��L��˪ǈ���Φę�6n��规g�LK�2�GM�k��j)�{�؆U-���x��u�o[7�1�G�3��86N����GW\s,+F���M�?e����/�<`������g)����u��U{��f�t�bࣱP�ۇ�ɱ��.>`�l��+�B	�+�[�ӳL��ex�N�#H6>wplW`;�c/��ETMq	�~�LT�Xb�����oW��p�p�<�(��<a'sIBF���b��1M���%�ާ�f�FC��rF���1�x�2T�d���S����'��T���WֿIk]Sy�c&tY�+�`G��ؤ�$>� �~,�r>6+�d��o����,�1?{S�hU&hi��D��"���2�ǔ�r����V���>[��u3���F�����^��J�f�`:�Y�(�6��T��AKY�m>vbgt��j\�\�R �Z�p�w�k:-�бM�1��;�Be5��ڗՉr~��V�鸷8���8$l�'؉���f丨����oS�;���XB2��QiFm/0�r�����C0�7`����o��'݋Co:)i?7U� q���\~�B����V:�8�	��
))f�7�B;#��k���A�K�Cќt�rc���J �DEl��@g=��I괆��3����?x�J�׳�~� ��z$_�A?1a��{����c\�D�;�Ų���2y�O�B��=�X-���(�p$��������e��
r�IF#[�$���WM�T���,����������W����'�Z�S4C�4�����=ؙzf{V{�FB̭�q��эl��)���N��
5�*ד�>�	c�'$[9,���r�S�'d�u3}s����F��[5��sS���A/�0��$�r�×ZG��u����r�#I�qR})�ʟ�� ��@��E�E���e߁�� 4��]$ư����v��F����Ij,�Ù!�RlV+�0��<��!��_0`�ixd`�{,3���M�=!�U���
��d�\�a����U0�,�$��h���g֦l��+�x�E~<������&�����/	�y���,�F
��T[r�	��M¾������?6��#�Zz֍baҢ����Ϭ�EU�n}?}1�n��cA<uE��� ���P4%b��lS�E��1�T��K���j��6��b ��(�R%�i4�n:O9A��<a�����T)��y�����+.�i��t������ P����&־h+7�%���E���mZ�9K8���q%�t�:p���D���\a	����6i%�`y첧���(���Q�E�ED����g�����W����l^e��N���:C�5ζ�֌�6� �:w}/�@l�_�G�ݽ�ɟ�.e� b��ܘ-��)vO]��
�^H�ո�QՀQ4 ¥�jn�E��l���sw�����*�)��b�YT-��x��v8z���7b�G���ܽX�Y��F��B^�#]���p�9���VQ�&�(Bқ�M>�H&]�!�kˈ�~<H-�!�!i���D��lB�\�M��
���1���H	&��ଫ)eJ�Z���Ȅ���±�m,x�P��4어Z�7��:��}�:Gik���&�6t�~�e�xA?�B��.v��&�lޢ9�~�b�sx�^|5���D/ѭ���l�|M,55G��^ҬiI��4������������F�>���3�X
��>�~�2t�)RhጱI�\qM��-��rT�o*-_��WN(��ҏ.آ��.˨ɬm��N�	�w�Wa<dre�A��������ݟ}�����a,�}p�]{y�q� P�1����:<��
z����'��<Ï؃�i�5��1})�ԯ��!�8��Ҵ=oϯ&�>��}�N�oءkQ@�ُ��C�6����	)��0�S{q+<�=U�h%T��!	�-ajM,-/m�L����\����D�9�!���j������S|��i^��z뀠}Y}��i$r�SDx��V�i������_ǁ�4��99)�iJ�R{+�J�볒6����,�]�dN��ژ9F�~T`͵��H8D�R���y*Pd#�M�R�U�-��xQQ+�~p��[�\E��Ƈ� ����/U��?-�G�w���<�'Y�?��/�~�p-�����[5�d�˙c�~oٷ�f��Ly������j[�����(�M�2�%,�˖�F����A�XMß�D刍0��]��3"ٺ������Z�����=�;/����bW@������>`�d�W����׃�@]K��h�y����+G��A�Ҳ��<%H^�'hquHdw�
U	�p֛�;�.
�\C�v�9|}Iaܤ��Ԃ|�[zNwF�QW���'�m,]�뫒	��bf���.���pb��m2rz�r�p�`����QX]���y�����ǳ}\fT�����V�5�2�cZ6�H����lF����|��u 1�>�|�ü�=���m���y��9@ϸ �Y��~Np�VeN�=�L�Б��Z�1����m<*�N���;�J��4�D�a8�ջ�'u�J	���ɕva�w\�S5A�d���l��.]?܎Jm@��$�Υ��߇�6�2��bK�Sc8DIϵ���;�쨋�H�������f�ͮ����k��,�|]�[�*ҋ2�������"����V�e�t�kN+�e�
�Ez�v�c��g��y�j4��Zeq}��]S�� �Q� Pq:7�-#��Q��Z�N%c�7� �����
yhk'�F�P�)�f��s�n4&�������_
�����Љ�||����aK�\���\ΌW@��A�V�D��V��G� �H�+�{�Z3�!"�Eհz����l����c�
�PTI�l���c���w����p`�UD�5 ���{�*ȈѢ�,��B�nhf䶧[��m�3!����5EV������zp6ds�?�0~��[;�R�K�F���u��A���k7���z��T�,�J�Go�*P�� (*[������Ů��uj�\e](��U%}���@X1���`Bm�2�jI�!}6[�Dta��C�::J{j���?�z��l���Gu7�f�R�6�r�A5�B3l���u,AþU�-�ǲ>@Xb�?a� \�n|�P�Sy4V��R+3L6B0�3�Po�5<Mg�;��<�r�TgB�GǑdQn(��wUK}=�3��om�bLcPO���H�u.|�g�>���1LS����0vi�����<��X��R��b����#� �r�x�. ����b��<�u�K��IbcÜN~��v�{+2�B&�>�<T5x����;�y_��3c��L�0d7�y�������iGN�Z�o=Bk��P{y��2c�(�Z�T�1+$N�]˝1���>}Ta��*hO�:q�A#�b�:��Z{w`�?�fT�0au3�J�;|l
wE2410�v��������qz����A��.���Y�r�m��)5��l��I�f�ڟ7W����� �Ê�,P��K}G��'�g.��4�Au�4O��7r����EB-�"f�9�Qe����9��5~�K$��ɕk��1��"�,.{>X#���Cz��SW�
%ς�)MwW�-$�}��R�	,�a����\�6�X�
�S^����3b/PҠ��̅�^�|�p���uv��Ój����o��vѕ��^�M��ٝ�c���lqo�����tm��?LW��Xo�d�cnf����:���ʸ]�����
ο���^S�� �O�]\��Oי&��� ��'d|��~������0�1m�G�b[Y�v�d�	vx���fp2��x���-�b6�jf/���At����_��X�禐ϘG��w�fzh��6��D��{�������Z��!A���\m���Jm��Wx��GL>�]Z8qBG����d,Bn zzqO�k4Hu�.F L3�,��:i]�	|#Q�Q�Ѯ��3�W�Nc�I?r�B��Wr�E8ya͛�<<k|+,���ش������d��9h� 6��g�  &���כ]]A��8����gU��fJ#�Ĥ�h��{�P�,F� ]��A,�y	hS����`,���������lb�+�D��Rl>�DX���u.Kl�I���+�ؒ���\r,#ak��=�~ү�KB�'��gs%,w�^��(3�F�%�
�0e�(���$J��`+�|�P���"��fЍ��k[�6tl"�	5�h*%`j�h�Y+�G'�Nµ���Q�_���테�	M��bW���uE�8yŚ��_�hì9�{�h����=�g^!�t<ό�ti�8<{Jo�a<�nEZ��"s���t�_C��<���GʽH�~��"�F3K��;a7pN��e2�m#��h��ٹIb}���k�Y]���ϛ����T�ڃ~_zG�@O�ĝ��M2��#<L����93\O�X�10��+����{��3��Cӹz��'�_ޚ�y�Q%�B,�o"U�@˧k%=M�h�s���s��K�����ܦ��kfA]�]>�ѽ��2��Zg,u�i��PC#ִ�~�=a��ԥ͠���!�c}�+��y��s��A�'�R�ǹ�)8!��+P��C�ߘoH�j���m���i�Ă�������H�'�[�u,��X�tZP�1�/~{Y����4O�&s�$C6��{�4�/�h'�;�o*��k�A�Kq4!��R|!0�S'�j�t�SR�z��[d�d.3^��Zy0������@e�Gz��V�1����߱۫�S�]�	�]7��Ҕ#���r6��sb�ҋ����{��ZK�|�}ا.��_��5�Z�Q�)��J&�+�R���Yll��!c�#M�4��6�U�����̏ܬ�!��1#T��#�{N�7�'c��W�Mh2�KE����e�5����2����� �+#~R;�Z��x�{��f�Cp0����X�����҆D��x�-����5	�`xE��"a��y͘~t����D��:� h��'P��IR��H3�{4�<��ݷ���WC.))�����St�K~���10��k�j��I�u�@�vh���������#����;0�J��'ҚS��Tܗ��ה�ӱq����0!�;pk�]���Z1�a3�������0i��� ����q�E8�v\� x��{af��e�V��rTo��)�Qj�*�3nm��8�sߜü��� d�C����N-��j����
[㙞���I����3��X[J�N�'ׁ����Fϥ���	���@��i��3�\��d^l���0��%�:Z��	��xY$OE��U�G�3h��$�����#��]�o�C��k#Q!�&x��m:���JOqJL�bz�������d��d!�w�,��کY����}��h�c��)��c�[�X5Ҥ5��N*7��� �� `�
I�� ��қIF����&�1������0gOzB�>����'�k>�Jr"|5?�q�"ぬT�D����f�)cA�2W.��iC"3�S�w3���t�OU��%��w�d�}a3L�I0(������z[�S�Zw����x5JeV�ՠ�p�W˧�u�Ah;�xX�e���;�l�N�7I?zi�� c��aa�	�]7V�ֹ?ϑ�d�%b[���e��:������c��G#&��C��� �,�V��]W<7w���h)�<��_��p�[l=A��G�Z�Z��u�������|i ��Jbr(I�!�%�'?uC�8��Ƀb�\��k��2S��!���v��d,�)�Ff�=A�ʧ����4�lS�kn�����~}ǲ�,���񑑘��W�ra�T�i �!kܷ� p���a�`���Ş�LhE8y$���{���y����4�9��P�:��kyp�f��W�V'��z�Gq8��ZZ#�lz�$�g��k��!�4������<�G����y}�g�m�\�����Z#��Ȉv�bv���!rh��Chޑ��*����3[�*����2�Ɨ(v�bd;����ix��qb��f�SO�G�~�����ڡd��P�8��U �H�2�i	p6I%�<��Y�˵;2Z�a��˼4�M�e�_�Η4ӛ�-!���;�J�=�Н��e>o�r�u� 5�C!ط��u�,W����p��#�EsP95R��[�^lz�b���'P�H�	��ebt��m��Z�� ��]��y�	���S���̗F#�fSh�"�.�h?�P���v&(�Z��� Ε����.�"�tO�r�y-T�Y���oAY�T$�5�C�V����ZN�m3�*�ÁD\��<|����A/#;Jڳ�q\@�^V�ǭ��� g}��!P��+'� ��d{}ud]� R�d��D��QI_>o:9D�:ߔE��/
i��@�`
u�2�WM��A0/L�W���E�3�0�*��O)�`Ԟ�.)�DU�e�"27��t\��*^���er��\k��Aڣ֊Edv�t�Rc�y��f�-$�q��H[ّ=��������9���yN�ܱ���lo���mO��g@��4�%)���@/�mekř���OR��p��2Ă*Y�?�΃���3؟�<��9��m"5O�v��$	�I�/ɯ��+P��'��Ic\��~�Qs��X޿K�Q���*� _�F����Wk?(�?KZ��ݐ�j�W[WXD`{Cp��8�zt-!;3϶�O�p�.�0+�)�����4�t��nYͪ?�����F:�ȑ=�-���J4T:OCps�N\��?u�{�aR���$7vg�\úB��-�?*+���'�����M���
������J8J�1����c���D��k�f��}�iP�',���y֑[ޣ���O��m�������W�p�d,@���W*)�$�s� G��/��T�ߞ1-x�c�����r��
\�4L�%+^�Mոw�Q��"+ʓ��!<I��ͯd�!D���؉S�8��_իr���vrk,����0�����X&<R������nS=1B�&5<��B��T�W79�2I�U,��"�Jiro�x;����'�O�1���������O�y1�K�F�U��:�Wú:�� �/����C��ͯX�Z2��������s�}۹"W'��O
���'�
um������n#x'�I[��Z�Y���ꤏ̿��צ�e�˷^m���hBcW2��իϹT�#T?6PG[�Ȱ,eGOo��P�
B���!�ǝ�1?{<��E<�WɮO,�^ ˙�����?��O���6��~�+�tt�?()}B"���Eb+C �Wd�<�J�h`ǈa�.� ���sv�p�ƭ�p�]ZBz���A�j�S��Sk�����Z���p��̩��;���9��f���L}�6aFٿ�?̥��J��~K+P��w�s�Κ�g���F�'62�tr���5��b�r= �w~�Y{�ȏ�������D��y�(-��oǆ�����Bqv1PФ�|����A �	BϴV��B��`~"�x7w�ǀ�ڄGlא��֧Qn+�K����=��sAh8r��t�M��d�ׂ���ۛɥI��U>�v��ԎO<PeW��U_؍1��)&?%#�q��(J}�M�=>�Gd��$c<T�M��w
��e�R6�Ȇl���z�o�3��qDb�Y8R8,��8#�xԔ EȄ��M��\U���
�4g�3��&'DՒr�Ǖ�!��;���_���1��L�f_��xm�iz��t��i�о��'� ]��xT��<[!�Ә}٧'�����bAN�Mh���|x3�>���쳲�ۿ�iNK�?3R����j�a{�>�"Bo΀�M�&��q�׾{�؄h��U�l�X���Ȉ�ׇ��K�=M�[��l/9>��v��
��k>G�TN�z���¶�-�5�A���CB�����1�k��t�'|lVi�~ƕhWV@�4��p��f���3����/��?gB&՞#CsG�R+�6Kk�Ax��t�ݼ�\8!���&A�#*��<�6���v1�p���h�-������Jg�;f��y�;���,�����ʽ�G^5!q�}�:TD�^7g72�Zv'��|C����	qU�x?��� {���2�m�H��S�%w83s	���a�s�/ ����qSWz~�!(K1m�4����̨�4� �aV��O�3A��͐،T��X_�,=K�U�Z3�1�6 ��\��y"S�
�Q��/�x.i�U�ɸ���J�z�0<��+����s0h*��A=�"w�NPr���v��k��'?c���w����!��`�ND*�������g�C�=%� X(�P�JS+b�5�.��w�p���*���o������c. ��BJ�C
�2�#���d9p��9�5���?IqO��>t!٨i��삊�Ų����k]�p|��B��+��p�Riv�$�Aosj�A&9�؅��W���\�>�<H[�P��͢Oz��.��"-Y�I��D����� �7���n	��lw�h�󭚽��$(�^/�Uj����Ⱦ@z��NY~��h���3]�^b�+{�^�Czk�$9�f$���(Z��YP>�|��#e�?!�����C#3-m��[���	x�%��u���A�z5��}�/��.!������Px�	;H�@O�C
	J�c�##�.~��J��C!���� ��INdw�f�.
�UcCC���x:�#�R���������!�C�i�2���iy�*���tv�� ��r��'��������¢�E~35�Pq^/�I�is@e��ŝ�����!>���� }g�-p��v���� N,J�82�љH�m䄣�y߿��F��)��'�/���QR<�B���z����Rf?}7�J� VZ{�S���UI�y�27O�ܖ_{��/Hl�kou���:�ٔ6*0�S�nï��͇7�#�t����ۦk�?��O`���j�:���+�ظy��/ލ?��E�+�$hf`cG�ި��d\�B��:�wh������S/Ek��C�.�thi�,�s�S?�>����
$Bn��}���"O ����h���L9"����-{^X�>I��B�����BH-!������-*��\,�듣vp��렙Z��ו����T�<;�V��I����)����jb̤`��x���P�˧���j��)ኈ��"W���?���p	"|B���s7"N}@���O}�Ν�g��n^v�&Ӕ���U��s���c�~�G�+�O�������� A�D3�i�rh��5+9��UB��/Wb1��+�\���Ҹ��?�
q���*�_NBA �I�cH��n��d����F���)��,T�'��c[a��h�ϑ��]z�=$�7�X��K���I�8`�gl����X�{=�슣ׇ
u!�J#�|_�f��߿C*�M؊�Y���&�r�D}|��Vz��:����04I��.�AfcmDM9z�'�Ƒ��'�{�;�M�s�t�����!Bp����\/ؗ��I���ӹE�ў��:�<��w��T��Y,A?J��Ϛ*M~/mj�n|�>`�\��ԝ{3�",Õ��u�*��ڬ��5�2p�5�[j����:�'%���A㨏�����ݿ��3���F�#P�*��AǞ�m������8�ޥ�~�܀=�&�GY����F�O���fJ� {n�)�g<v���Gv��Bv��l4��Op�*����E���,��]�E����߱�*�V�C.�H.�{2Z/����xj\b��E6�Px�N���,|P���s�MT��O
L-:� G
���^��-�V��%����}��Ԏ�ٳ0�c���`�!)� �I�G��ۗ,�hA��=�BS��6� s���E�4f;����N~c���<8��E#rb��Ή+ѿIG�U�;�Q�cFa*$q0��q�R�s.qyO���i�qu����;�y=Qm�ɯ�S�A ���󃞠��ޢ��~�k��L�1W	Ӿ@��H�+!&���[ԅ��F����@�~����<>1h}d�q<E��4��-���,N�H8��X��;�xp.�%��^���BHۡ�i/�d��N��h�K���|��VF	.u���Y����Q�1Y7����: ׹M��V�Zb" ]� ��h�D	k���Z.��5���3�fo��ȳD�x|
�^�<N��Kk�
�=Y]k��l�6��pF�#DS�TI��9/E������*��3�> �S�2��xf�2�^��v��i�J��;nõ���N	�h	 JJ�JP*̠�O@�]�h�4-�>]v�Y��c�Q+`�ítU�CM�.	@���y��)�w�$.����*n���� a�4�c������
�+�4�iF�R�`�T��yئ��v_��ݕ�
��L�0n�V�����@����mD~A�U�� �6��+:��"-�%��-L��~�ǟj�5�K�U7�����XY�mu�R H`�*`��s� ���@����X���&co�����z6�ӈLL1j{{m�o�G@���?zj�!��c&	�|�%��۹������\D�QA���f~�k��
�׉4.;�o�p�Z9б���c ��3*S\�[���_q_^/���Ζ�Wo���B��X�/㷒��9��a*QȬ<���h�J�P�!	��o ��!��"��Z���d퓻v�X�'�g�/[+�f\_x�C�r��)aFM������U��������in�����f<���B%������3P���󶬛�Z����B��"u\��At7�Fv��VOg�H~�����)��U{7k�p����g(1X8�/�y�R�I�סS�GR�:5w��������:�H�^�j�+'��#1>����}�� �[Ѥ5j����Հ-c;~� H��t`�R���cNFG�8����['HO6Df*;&�K4�ās��#Q�U���Pn($��2��\���m��Z$a�
k㦝ڰ�[��V��q;�q��T7[��G��ό�}B�,�0��'M3G���'
d�|���@T+�T	��8��OU����6�e�u��1�HF��b��?_�R�z�U��t/�B�l-jnGtYc���A��w���DEy�_�IȬ��-�W:�r����ݰRz�����!xTxQ�)Y4�UI�㗚d5be]�}�=I��'�w?��(/�֜6�M�
��>�=�6&��ł$�7^'��v�MN��&l]�Eg1���5����J�5����I���ٺ��)�����6'e�!�X�Mۺ�f�����1n��%.�2��(p�]���gvJ�z5�v�f�����Ly9^��T��,։2��F�[l�TGAF�Gӂ~?D	r�����ЍO� �Ƒz*�y�6��-^m!s�e�<������e�x)
S���I����,�������ȝ�ύ�GDy����)����d{�ۮ����!���y�gհF,���r� Na*�"cM	�>P����!(�33k#�c'�K&􁐤��RE�¡y�<۱����fVuq� 	�8K`��TZ��[u;��!�_��qOAB��7�^��Ի��Dab�$0��6��?$��y
cƖ�����g�Ϲ��o��R>e����⓰�?Ƃ�p]n�9�]��$9�`�1_n޿��]��:����y�kR8�x�;%��g�7[��r����!����s�׿�N�A�=�#��� �@׭���6g����~ �-2iv~�(��n��/�_���??")?a8�z�?�h|�&�_�b]��2
�w�̓����3��s�ٞ\�_��G�VM�B�V��#7�:h�ub�Jֻ#jd��Q�PNE�JP��o0�]wH|7zC�k#)���?gZ�u��<V�H �Ǐ�3�~�*�5��i�iS��~�'�rx20�E�����Ң��⛰ˆ70���>�}��(�Ի���B�Z��a��I��9�����RlPH��J�TPZ�s�\�hK^�f\Vh�j���/<���c��v\Z�^� ��ܞ���'2���XbV<!5�ы�wyX*قL����g8��~������]G�2����dA�8nB6�F$^�e��-�).P-�V��S�x�39�H������}X�<{�
TY4-���1&�:ܭ�8>��� bԻ46HB�'I�W�5�����&3���r�K���� UF2p.���,�X%�2�LOna�Ƭ�h^8��`j)�R�����}ɤl���&���U��)���0�� �I���x������0I9�%'�v����Q����T,�>;U��<�^����hy��OG��V2� ;Mo�F�8��w';�8�+��\z������-e�������`�C*�@5+/���EH���\i��57�_,AK;zן�����B`�M9Sٶp��q��j�v�_��C�G&����.ú�M��O|�8�k��p�%8H��d���d+.&D�Y~ZlA%n�퍏ֵ���
�Ӹ<�6+�^����wG'V:����59�i{��Q ^��o` �g������k�I֬-^���@�]b��j�aRY`�~�+����'a��74+�y��?6e�g�l[�	qd����l1J/L<��,>�I~�m�&��s��?�p�={��ѕ���S6�nG�ȴH.#�$H�q���ه�:Px�⹑��8��__�-�k�w���F��=b�q�qE�^��� ��JڨZ{L[2�m���D>7�u��Ku���i���� ��K�wy��N��n�T��ѻ�X����bN ~5q۝,��ۿ�x[A��o�y�PLU5t���v�hb����Z�K�YK�wiж-x��k�,-��Y�F��<T�'WđD� (��5I_�O��HXO�?,��&*0d�؄�'Q�!J�[�XA,�#���몒�KWx��8�� �'�eQ4|琚�!E�w��d�cy�[ۡ'��!@	 ���D!�i���fy<����m�\-�[7kD}�5���%�����1�dA�n*,��"X����]��_!9J��v]�q {�*�ƴt������v"8�"^�+���ސ Oհ�H��%��TF�ű��GiV�A���9dȞ&�� ?9B�^�li�J�Aՙn�!���&�!3�#�h�Þ,��請q�j�d=���śgU�e��r��R��ng�ܬɎ|b��[�r�;�^�|'�G���3�5pA�򀯝#��u�c!��衮�4��͒���
����H�xD�#��H8mͰ7k�ܪ�4V�
�C�m���D\Dp��'��� 캌'\����1��mJޢ�S�&/*ذ։�j�0���c:X��.&�%�miYC����/�~� 8,��Դ���L�+�m_�ˬ�k��~��J
���+C���kw?�c�>Jn�&mg(�t@A\��e�ۢ	��=��rA<��Pc��?���ғ�}��eP�Bxk}�4aD��l:�nO�YV?���,��Q5���W!��+�XT_��J؎3
[ƍ���r�?Z���j��W}����j&��ăcޮ���~�c���-.�~���X����v'yɢ���ŰXᖕ௣Щ��L�|7�|Wz�L��RQ�T��aH�c��sKga-�� �{��a,G�����lF���:X=5�V�VѲ��M;�������K�Q��%��(/�$F��TK�������w��)�{F�N0��8��2|M���0]��e�z<1=O��SxoLʙ�d�z6Z��&���\��u�5>łG���i�%!�˕�S�רOke�K��I7���:BŤ���s���Lz�b��:��N��fR#�=~�+t����BD�o����n�_"���7�{׹���Vd�"���5�8��0�p[��$[���J��@ن'R�|�(�vx�3]����lI�QL��x�&��g0d�{�P��ypW'F�NKz'��ʗ��ە��Sp�Þ�"	_��Ev>H��ݧ@��&ڋzlH�"�/�%�������ۄ�"Q�H�OTR�kX^��d|_F0�G�����W߾:�Jc��@�\�qTA^愋�biz|AW��
��������f��e�;OD�X��*�`��jF3�������|K�e��J��8;����5+��!�{&R�8EQ{��T��j�_J�*�W�b���$_Z��d'D�4����͚ҋ��0�GV�e1��V��U�	)�|��Q��D���r��c�-|I��L��⦈��k.� �<�x�Iae�Ћ�	�0��<Bc:75����n!u�MoڕӪ���u��^A�41��k�8�;�2�yp6W��c��p�v͆�h�s�h�-�m�گ���碸� ��	�g�Yf�p?iW�b'/�����$�Y]Sіn�<�#"v"�i�GѠ�tG	5���SҶ���f#FE�N��|AY���x�^�G�4�K�G��n�]m;o'���a��<��)޶ �S�+}��r�;.�
LT�J��\[�س�~���?��;��fq;��[pL�������ոR��@��L�*rC����\p!*XpG���8Ƙ��ş���[�����?�9 >�ɻ���*P����5���ۡZ���X��iܫ[�|&���vU����dW�*���,�VH�W]�L5�ItydNd6�9O�4S�@롧A�U�f`�����>D��`8+�"�;�!���8	�@7O��X�D�%��	�hz�9�T�0\[ښ.�%���DR[i��A�76#C� �ޮ�*�Ǣ^�NY:"��q��4Cve�jn �����ֵW��&C���LafxB�r���yĀ U����R������/bo��玾uƖn0d���l��m-�a��[sr!��,kr�Ҹf+��{�R\ѳJ�$>q٭�.{c�?�Q���0�xYI��M��5hy%�;(ξ�@R1��L�~7S��vóD�I�$�r.���i��Ȼ��4^�;p���Af�i�>�W7�+Ч�ws�cv��]�y�m����$�-������ �u������*v����!P��
��!v�>$�zJDk���r9x�/t+Rd�=P�5�R w�{ڞ�Q>���P�{c���՜Z��a�m@;����:�	�s�w��ߐଢ଼\u#��G�ԙ�#�C��@� �|�J�x�*�9�&�1��bp/����4�B��xڋݕG�!`���������)�e��g2mcV��Ynͩc��m����!��W�E"SP�W�-4�N�)��"���6?̳�
�oq��Y�.�2��jC���P"��*������FZ9	��E�Q�,��X~II�.�)��UN��8M23rA�an�g9��9�]*ۧ|��典�%����G�1ɚN�� Ux���kP ��W�R�ci~�Q����fG��	�J�Z��䰇�+]Q8B��d�SР�2�A�Z6E�ʢ�D�dn�0�췳�t��f3�8�<�g�Й�I�� L��	���d��j9�~)�D��o��sZm�' 4��M�;�!�'�6�/j!����F�D��֭����6}��Sz|{-v{���rg���d�z�|�q�9���,}_U�^l����k��w���W��{�o���
&Pz�����1B���!ye�bz��I���N��W}N�"��uM�Q���n��	�q=p��C���v��ģ��ީ�,�YI�����%�־�i�9������7���	\7I��8���V��V�py�kXc�j��=�k�>�͒�G��|���XY�&�"�l�͖�� �[FfG�,�T�����u��\��VI�0�RJ�L�b��6傲�\�Pv�٤�v����?Hl�<��+�[�s]��*�D�K�Pg&E��.��4�S�ڝ��I��0�����jO!�wی��������B���n��+�#�M���y�6�̉��*�,����������e$�V^M�|�礫8����o���691�<��Ip������zW2�X��s�G�#=ž\�F1�g����r͂	Jy���DPg@Bn��3o{0� �Vͧ���s�f�z4��e��x�O+��?����Gws��s�a��=$���!�<���ܚ;������[">��~� Ȱ�������Y���C���Az�ӡKU�X��9�� �����,�
��A�@S��k����(p�98<��p�N���$�=�"@�й?�� j957JV�C�<�4tk����=i,���Dm����,�=��{kȻ6�6��P���������1�9�5�Q�����7]�4��M��.�9.�ܛ�F�P���� �/G$��^�`��XJ`7�y½�ځKT�w���M�j���0|w�<>�Kt�K�CO\����qWņr�zg��-�PAw�2c�,˖�j���`Z����������P8��c�-,Bf��@e������	��Z:[�*���}�����(<�RUׁ"UKc�~�.��_��5��R��h������s=��zd�/��\�}ؓC� �bbi���wHG�-6"���s�^�j~�4h϶Fp �r:��e�M^E/.�Ǌ�V�(�p[�\ɽm*��x�@����#K���[UV��.�I��M*�tJ��joY�>�)�)���#� 9��2B�.�D��M��a�:�4&�I�#�<w�XI��}�8-:ĔU�Q����ԏ�<&Y:P���\L��Dd����{��$�\0�49�#(jO���g~o
31�A)��{r�S�=��t�6��$e�V�z/�Y����,�3��잉�L��c��ȣ�����T,q�6�t� ��l�qxlh�9IƄ���҂���;=K�쀾�|���b44�q��qf*l��,__�|��ԇb1��	��-(dz�e��j;�B����KeݾnPt�0�6�Cz��j�E�Ws]�_�h��-g��#0ql�k���]'u�
q�j�6��J�j�J�?�����h&�U曜�8$�ݑm��@�C=L-�+��Q�Ȱ0��&O1r����~ϗ|�z���
+�r�j���,�n�R��c
��ӊ�K`jIg��H�#���b�����2����y�8��S�æ敃N�5��f�y�����Y@nJv,29�rŴ�к����5����.>�����;�q�pjC[�'<��M�l�X�e�_L�V�_��+���+~�O�%&I��X�%��k�=���n� �"n���j_�pM*��pw�����W�Or��[V��E|,���W2یhk�㛸�(�׮ ��<73��a���c_D`�ҧ2��S�-����m?��W1��ZR��E��K!������|c&}�q�VO���.R�S��߾��5a3s�L���1�jNѲ�,Kz ��,d5n�������A� ���<F���B!�E$�;�,�����şc�!�.j����q0��0�=�C1EY�[KS�Z�y�&~[�p	�*�p������r�����h~�mщ"��I��9���|�"�2�<����W�� �Ty��<��qM�qJG�p �o����1�<��|��ז[y���Br�l���P�(c����0�	ա��� ���Ȅ�9F���D*f�`�H�vX�&>�Q�PZ�v��ߐ��v�%���ac̈́��}�.��0/��<I��N�W����:D3�?E��ݔ��R�L�Q��AQ�WV[��2?o�n��].��^�X3@��� ���4)Z����d0z��g|f�"���Mc�t�79)0��J���ٖX6 Ө�]9���P�`�9��0��8EO�f[��9��)O:�mJX��ZxV�9�FJ�
�� u�����.��'u|i�:����(���BN�����XH�ΟE�8N�x�׃�!�Z�0�&Mo���W� έ�����!\R7�4 �?x-���+���əm�5>�b9�x�k����(�"����CJR�kUĮ���*�(��O��1\��]{�.c��j*!��WB��ʒ%Z���57��5���9d�L�7I�j�
A��f�#�Ύ�]~c��������
���OE�P�"��4��~�D��/>��?\���'|O£͖�н�3xW���a|U��cя>��Dq^���^,������Cd��l�z(�Gr�Z(E��zcԁ�vF �(�.��Av�!S��4�N�q�6D�ޔXv|Q	O��C"箢�jϿ�߽|i��Չ��ߜe&�%�'��O�3JAU�f�썫_���Ù��vN�4�+�T�ڧY�����k���8#����#S����S4h��w뻫a�dF��Ȝ���;����W��\��I���D�*I���
����(K��ѽ�$bT7�솾��I�4��8�_�_
��:�oВ�Zc�j~ģ�Xtg���,�)�^��V�	��Kz�j	����	�M_a���~U7��La��`�v������5�Q#
-Y����<ھ��D�K�� �ؓ�� ��d=�����i]����^�M/Ɥ����+�6�Cڵ�Eѻ�k4��ھ	}陦���7�<E�TG���=�%`	��pB~�1�R=E���|)��H�0�^`N-Z���&0EѼ��I�x��ݷj��聛�:v�2ѩPO�ZN�j$6��+hm��C���Ä�$���9�
�ubjI����|��DvUD��ӟ+@2jf�8b�0�ĤϚ����a�i�'Պ�jB���bW�׮����V�������t^�:���f��N6LE����BZ�4#��S�ꭺ�k���*�P�b����8���H���S΁�f?k��r
V�$� D{ceAY��}O��� w���7e�D�����k$��_���N� S��1�YYlW����|qB�Ȥ{E)�!8B>�פV�;:�f���pN�xD2f�����ٮ��x�S��Ƅ��b��3�߱ѺA 2yxYm?�"���K\Y������>KuC� {�9C0\M���<ȸq�������>&1W�-����i�L ϘR@�5�����5{��4BV�����{�d �
T�i6SGT�D>{޲�s��
b��L�P�~��v��t����Z�]�&�j�W3I����3D�o=�c��*W�00��=��1��/ݲ��Z��f. ���WYJb@>ۑ$|��cq��k�5��"NlI��~�cb�~Y[`&k7~�'6�,u�^\�GJ�߶?��2�a�	\ɔ����=v6$�#x��D�<��Qj��5ͪa������v�ԈrC��k� @�b󊎤�n�'�4ྫྷ����[�} ����̘OR���+R�����Ish��-z5�f���U|����mxB�k��A�I)w�>xʙ����9%�tL���B(�ө�	�� ��m�|KH �
����3₴w�G� ��y��!w)Do�`}��5M�{.��!�p{��h�Ȭ�70f�A(��/��N蕔�tf�3{{��j@S�����!p�sGl)�7>��TT�:��3c��K�sz�nV��l�U;��U�"^3\��r�mc��G�y�Na�.a�]��%���O#�O)����h�<@�����.U)+�^T�	`��=m�߇/�&O ��Äi�(��8���A�f<�З����0�N�M˴`TZɣ�>�J��@� :-����\AT�
^8
X[��=
ij@	��LXտ�Ve^����@�o��.�,�-E���J�4��hu0l��k���x��r�-��3��~��`^� .�~�pj����;�m�f{�����`nďr"�� \b������Z�ं��"["�P�O�gn��;A!>al9���T���-�Fh���_���F��r����q�rዝ�;]l��3^Z,N%vx�F�8��*Z��Y��,o|un�Z�;�b�[�r~�f�����X���@[�	 ��$�*��Ԃ��C��)V�n���fbb��oq	G��%�ۀ��H�C(��_6���6{{ �9�B9ѦOg��?P{��8� r���yjt���K�h���L<+��%����������ɒ�Se�tK�m%��d��u����OY�/P�@����ʹ9���k��	Y�UZ���8��ynpTM��VR0���r)U��T�44Ԭiݒk�ʥ�������J�����������ؕ��\l2��=i�W��Ҙ$����Rʻx�x�@է���'��:��t���Z���H�!-R :����I�ױ������O���ql)^��}����
����������:�r����j��p�����F�| x�է��\FA?�)�����-�pLETkP�i��E�8�Œ�\�"-�~�̥��L���ƚ>�\1���dy~����9��\`SGyWo��ȇ5��.5-1�X�_$��]��(�V!��{��^T'k���]�JiK)���@(Q��Q*�*�4�O[��1�Q�i>�3j�Z{��f7I<����Ln,r�%H$z��E��B���U��[����=,H�̴:T�eW���T�cZ�E�z,[�";�<�VI3\:W=�+�eq��tM.m~`�/S����{�aB������	͵MQ�?Dx��Yb	��@=�z�-��F����x�@�ɯU5���I�儕�6��]D6�r_	���M�Xo-�CULZ��w�,���=0�O�e9�&���F���̓e��
�`�ĲBMdo��\\���N}gkd$�˽CX!`�g8Pm�G˰��ˠ�@%�ԡ�T�1���5�{W�m|Q#{Q^�tC-�1�@�C�w�������$Ua<F�0�IU��ObzF�g����@]��@�	���,w�gӲr���W#�P(�B������+�"��Φ�����Vi�)��4	z��9JrsB���6�<���a�P�ZR�χ��������<������s��^�U�KX���Q$��x~꽧�V�������g��<�!��;u�\?e��њ�La���q�����.��Pzm�p"��e��^�F_�50��ߒ�u£�w����^CU�{Y[/[z�8��f�=)�����A��Q�*^����NI X�q������s�!#xEy����o����#���$��	�2���;�A�yn�
���*���t9?:��
t��ڍ'^��^���)+�&$�u\$blӍo�]�N�R�B�4�ֻ	ke>k�!�J��T6���RѹY���A��Y�|��9��.(ǽy�s�Q�'�x�T�h�a���A����-7�\�<y���0��BQ>���r�6?�b�hc63��wm(6f	��A��mϊ�=aO�����ǩ�{��ūE��n�y��?eY�x��B(y� ��ɬ�ыӟT'p�O�.Y!�*b���4Fq��^(�#J�W��-�'F�c�q�L�x�����e��������L�ܳ����)1�Ph�_�D�����Hf���r����X`H�`��ϒ��FGS��Y(�B%��
�K�
��s'*���g]5�F]$$b7����;Z@� q�n�OI��	�2M�vl�ﴤ(X���)��e0��+��I}���\���&͟���v��"��%E�4��Z�}���)���3�����D Tϱ��o"�}I2n�kV�;lr���M3�yzt�nX��h�0���E%ro�D_а���!��E(�mo�_�E���;�d���7�~-�&�z���R�P:��n�0_������;hKkWQ��ݴx����B�aVp�u���{=ov���(�����g��3 E|/��%���N�2_Cw�/�:3,fP��i�P6b��b����ƙ��`$����G�mAfh�)3k��/�[���ĮcH������3-�j�s����PVӜbD���)��bU�B�s�|���9���HƲ��ܸ,}���ZQy��J%8R�9�$a�	,(�Yr�Y���14��F����p  �Oc�y;�?�����i�G���m�ؽ���8�aa�[�~Q����n=�x�:W�* ��a�_z��E;�K��g���mj;��-hK�5�Q�{#�BF-Q@�>̔�څ�����_��(�oO��:��ބd!j�����{����r\�d�E���3��M��o��d�F �p]Grc�n���Ɋ������P�u*CBL����=���������5NK���}/�n��M��_���R�c�-��ȕ�ݳH�����׾Tdc�yyx`�7��;�ω�H��ɔ]��t4�%�t@�Dۨ�J�N������ ]�3҇Iq6����)��~LaҶ��X͂ �m�v������p_���"�.Y̩����Ϳ>8��E�<e�JV=7�"H�8�4���mo����EI�D����� ,��K�����)s?�ݳWz��.;����v��־P�0ҋ��TQL[�����\ �e\ׁ���H��q�����ۭ����IZP������mA;y�F#ŻYC#��^O�5�F.��&��D�6v������Fȯ` �I���`#2�.���b�.�z�t�N���c���)���^T��D�1��R�F��*�2_���C�k^I�3�Qχ�I��E�Q�$n�Ӕ���-ye�]x
p�rle��8Ы��?!�ܝ��R���ƙŒv!_r�V��beWǇSr]1��j��V�7��nQ�O�YN�#�l�ä�צ�r�2�O�t�O!��~YT~5s�� Sc�P����p�q��p�k^q�E����������\g���+	��qEj�c�JWU{�v��
X��)���^>[�~RnK�[�b6��18(+u������o'l��r��� ��tr3V���8u�A�H[�����eiN�tjv�Ƕ
<�1��;}�t�m���Wd�;��S������iA�����MX��E;�	� �lE/��w��'4P7���ls�V��0��/Θވ�~z�	��M|'����|e?���g2&�5zd8gyP�m��G[Tg��=�Xq"�H��hK�Ij��C�Ţ�mk^=])�7h���% �W}�X�8���@�n�~�tL�����Wԝ$�r����m�t�LDl+?����',��4�7KW����4��!��B�n����<y��U3��4Yn��������Tc� 
��N�(���Ƃ$K8�Z�Y�"�+�g��$�%`�o����@2�j�t�<hK����� �!�G�M�69�0H�z��^�ё4<d���|�a��o���v.;�5�
%S�^�2y��an��Rot��XSG�|�N�H���\���|J^mm��:z+-dp�>�>��B�^{�>�'�"ˬ%nG%�	��(=���oؼJ�5O����J0-�.�|�d!����o��Q��"4�r �׬ȸ����I��QUu��*0#�1�-W8R
����;K�o*��Y���xI�䇗�x(�(�UI�E�W�l�k��j���u��5Z4�Y� ���|������,�-����%�	�Q��k@� �� 9|<� pM�{o�m��8���1_B�<\�Q�9��V���@9�槅� |'�� �Sr<D!��5/�E�hW\np�'
��+�QO����Olp��uŐb(i%�V�̥��,j$2X8bsC�W��2*-Q9x�=|%fd�u�f���$�|2�{z�����5�D�:/��\�DF8~�#�/�ų�)h1���d;x�"Ԅ�M�I̘�3K�I3J�\(Rv�� �i����֠ο��S�Gֶ�{�"&��2��9��)D��.�,�������w�?��x�[M�'���JG���c?\MA6��i��0Vp��Ĩ� ��;?3���@�Ţ��.�qڿg'u(u���V��lF?�s�y�v��tb�Fq+ ��:%�Vͨɉ��h�P����,��&��͏rwaW6���v$�착�`���3��N�S:�>���J7���#8��^@_��m�y�����SV�3��k$�1��`�������M���v`��kz&�"ˇh�G/�/�N9��f�q	2�I�??��g�nD�-���7�Oճ�
J={�^^Pk�U6�O���1���������#?��ۥ���c��[�����t`.��+9#�I��PD�%7>�Q��,o@Nh���a�C��!临�@�Lr�a�{
�@���]נ��!��h�*���N�M#��`���a���3y� lO�!9�`T�6�<���S��L�.���sj��� c�M�t����`��wRݗ�E����f��d<�S]X�,�_��1�����/�'��0����0iA�2�78��\Wä�pW�'Ug�}��iQ��*��򫩶�GX��-q�ۈ\�ɯ��F�l{���e*V�{$"���;��sgM�[u�\К��}��R���;]&.���j�S�:���:���h`�?� cq�,uQ��G=�@$����q,����ĶYh��E��w�*����aX�'m���dh;I �ۤ)��<�B}uw�o*d�m@�uh�W�������,��9N+ >a��otyѳ�3�]�A'>+/Q����\����ڨ��E�&v��_X9;�9�������B��fvAr�(`[h�i|�7�aa��2��\�����N��D4.Q���?�+6��fu�'�;��湊7�Ki�ߊ[ �>Nx�˔�����#Na.5�����U��f:i��媁��M�6�<7`�ɟæM��!/3p���Egg,+x2�sW��]���]�u�G�G����� ~��pYv�41[|?Os�MV�v�jU6+�?��B�[����O�_W�֍��o!�'��K~h��AM����1�����eRX.|ȼĪ�f������z�n���	B���������Ӓ��z -��A��Pυ��ŽD���8�GFT�8&˧�fA���CFK�G7���5��x׌����<�XL�i7�뱵�v���|�ڠ]�����{ܬ&�N�����'�a���bmb;�B[Ջ��;vLz�#�۳�
I���v�\	�Ձb��a�KH�]����z�R��Y��w�s�e��z���֋
V����a�F��)�,�(�8��Ԯ.e�AC��Z��p�?�u�1���6ľ���0�^�)�+�Z~n��6��[4��״�Y����S�`[8�BO2����.h^��I�F7'yh����_�OF�r�B��y��D�X�W1idJk�g���2Lh�x���"�]�W���{�Ī������O��զ����8�&`m��ҤN8Q%�ý��~Y�J�]}Pr4uI�)�U
�產�2��%}k�S�δe���x��D�!�(6@H|_a�CAv�5�B���5�t���p#k������a��W_���8���y��"���g��B�-����yV
z�9�_)��ti�wv�Q�b��k�j�C����v���Q.G��/|�I��3��3�iv��?lZz��P�zĂ��ԛ� �h��J��V���A��f����;�2YX���1U����Wka*wL���؍e���!;���0�.�/�5���.�~!�Z�V�cdR�c�w����0�����"�����Uh�5@�Y$�5�~y��b�F�I��%������T.ɫ蟍!b�ds/�;�R��aXvV���#�JI�䗢t���ɛx���,�pQ�K���:����L"�F`��(����>^��>��Q~/J�b,?��
���D�M;Pz�bGM�u�A}S���0��j�벞��-)�O#��y�]��9	��
J�B̈�c[��y/�%���%��	�������;�z���}��Q7�N���ƙY�}�UP�Ff�z�[��O<��Y�&�p��y���n6��YJ���*��r�Qs,h�a3� �W}�K�Fl���|���K98޳}Ĳ~r�]Б�?&f7�$A7,,�`~�������W!�xq�ñ)�FI#����i "Wu��.�.ڬ�F>8=�	����W�Ʃ��_7:Z#2�x���4�- ��YX+�H�Z�&�w��5��j4������iDgLD}l�ؤީ�[K�V,��~�����Y��5�nvC�p�,W�Q�4���AH,�3��ת�e���%�:�De b>��	���RWyw�;}�f��iH=��}ۡz�OOW�@�s-GYu�5 �1�j^��P}�C�� HC��5������~CB�b�T���z��0ޜ��8WN��\J�q�Ws��Q�X#$��2�7G�l��,ژ'��k/�����KAE["�l�%l1�qW�ř�{��38�M=͐.�0J�X��/�J�w�s4��D��
gc׈�<q�V,<d�b�'�t�o����3�(u;�*�S�YQf�FU��\Lq��&1��+۫�(t����x�(z�w��@g��qW�g���XS#�$�k*w�2�� ��3;��d^�˵1��CrG[Ӛl�Gh7�����vu�Hw���M�]߶c�n}�y:�2��V�7��� �&��	z^&�H@���DE=9[�|^�{ 9��k����� D��Ѓ�LR*�W$�td��	�73^������aAE��/=z
ђ�_ouԝƲ���
�<����/�к2Q���$�_�E�,m���,4�]GRzA��B�kݷ�rsj�<�Gň-� Ɲ�ݹ��o˵;��W�+�XakP��4Q0u�z�pX��R��t<�E@�,��I�C&o\s�jE�����~�����o��Q�V�b�@UD8�Շu�x��P�'�gS�e���>���`���a�͘��;0oƐm��`�!z�������o�,�H�h�%���
;�:�K��pK���q�	ZaU����=oL��~�.�SB4	�b�eJ�( {�m��'3��%n�al8��h<��h��_U�uҁө�b^6G)@��<��1��Ue�&	��vƘ>&]�)��F}S^P���^ҜbK��BC�!H�Iv=���`�m�Mǿ��ׇ{�79�ȕ�x��.UV���]9N��Զ:�4�}�$��{U��8�]U�ƨtpP�%�F�����N�S���{j�蝨;���4fS���V������F�h	"��s��>Qt--�C"稹���VE��f���;�7[L�bֵ*6D��HǬ>�kƧ�\o���{sx`-d�⛍u�xR�F��Ӳ|���c�"�S�T���F]I]����M<�j8,���=��B-̑�������c��B�3�z�i�3��z����O�B�v���%�M_�f�<sg��2;ñ��?���8��<)���/S��I�2����H!N�S�7{����n�Z�k������~j�N[����&ȭ??&�6ޛ?H�-�a)��,�Bh��#�|2�A����
��(V��p��q�n쒸�lA�0ϦlB�Ks��Z���mD��r��`�[8�HḟC1d1�M@n&�r��(=��KF���7txe��	�Z���l�X#�tZ�He�
|�}�+��^}V��< ��>�o*�:mV�[N��������@��q�[	O�0��a�T�'���M�����J[ǈ��H~��c{"zD���4�?Zl�AL��S(F3�����a���f^����Rc���'C<I��_D��uc<�ٞ��p��׃�����T�������B�MWA��,�%�tG�Vf�e�X�P��C��H�Qy���~D��܍�� g���3��o|�B�m �W	��=��^oe�N�M^�/U<^��˧���F�PM֕����p��ʃO@���)�o�ր��r�]51ّ��*�VP��y����8���J*��0���/���=���>Q��G U=���!�TƝ��4 w��%���9Dr��7S�9�K����}e�"^��%��<�l�E8�����&�C-5z_���(rb��y�(gI�-�]��v�ت��K�YS�����֛h�Z������^|���[������È�5�f4�ז�/���YQ��DMhF	E���!pl��O�)u�;<��?� �T�A�w�Ǎ�޿�Wy����E<�����Wї�!��.�m����)&���b߯��70��ؐ��c��.�T�Z��4w:��Rfh��nZE�*.8=���p��@R�G�6 8��v����H��~�<~tV�s@l��ҥ�@�j��K�>f��o��f��������縧(����-{Ɠ��fc�(o��<ޗw5�`SS����J!�m�:-�(r�w[����A���k�m���E;c�������"���a�ǖ!��
���#�f��a�	=dSx(�Qc�!�ita�{c��F*v��F9����"�K~a�{nqЦ�F-��\5��WsE ��*��G�!�"�(H K� M�Ԉ->P�o�9L�����0@3�p����8���!×2Z�v^g�S�ګѳn�v�lE:�FR��K�1��7����I/LZр��2#FY��]�����A�9"W�'qN�6!/����o��]�ùn"��v�:���!�'����b����w�ʿ5b_O�Z��ujZ�`�W��bT�FT3�,�G��D��ZDu��XJ�[0Xcq�e�ͨ�]	�s�靖�����G�lU�x4��T4��H!a�M��G�Pa�]���t�
�̓�)E)7vp���%U��G� �ȃj����i�k��PX���v'����	r�1򇌮2�C)1;�p��4��.σ�:vM�[��D��2�΀J�#��T����u���踐)�sPR<l���cܕC�D���HQ��gKM������{�ϳ��M�#�^���G��{�yZ#<i�f�8G=�2q�&��tBd}^��o6�@V8���E1�t�>�B����#�;���fP���3�m�w�����^p���fZ*Hr��W��9����g���z�|�'͘���=�a40Y���W@����]�'���ǘ̦�?�Z ��/�^�����s)r���p!u��A���~t�BI��걏7�ez9檻k�`|~+���Tє���a���iy��_�%������C�@�k����[�ғ#��������9a�ᗪ�E�.q�?�ԭ��b9Y�~c��ώ�3���2�1����w�žP�e�ג���T����G�jr�D�-W}�����Nw���Wr��Ľ��yO�|�'�p����˒�@�� �g>�྽�H����4����q�7UA��WDO�]˜ �?�Y+T�����C'�$���C5�	Q��z�W�)H�#os_��q����M��Jf�8]]���u����ȷޒ��P<T~�\�CGك��`�ΎmcW	���_V��׃�j�>��Z��v'�s��u�2$.�F"���u�:l*LhwiB�����j��ʲ��+��/�xi��M�l�$F�p�IR��8| �6z��n%0F�~!���53�OC}q�z�xh�&����~��`4�β	�n}L����T"��N�#�`		+.�N��@_L<B�kiO��
^�-Q��W؏e�ؿ�,�q���[Q�+'���[9W����`^sAoe��լU�zN���F��J�۔��6~�$Cϊ�3�m���=��X�-���fs5�Šq�i�}���r�ӈ��]'h���
�/�00'L�i�ug��h�tD�[o���s:�z��>��~�\6s�w��b��X�1�e��y��޽t<�Z&������K�h[~� _Lef��~�=s7�m-�b��E�򺀅�GԐn(9�7*����-g�A�]$Ǽe��LF�{䈠G�[T�r�i�'�\>�e/�Lo9����ǒ/pe�*I����u+����˞�.B��PV��i���%|� l�%�S�\�H���h��{a�s��Zb��-٤��<r�O�u�&�5�8�C�����ĢG:y����Z>���l��c+d+���$?�L�)p�p�K%3�?�b���74�*�(K;!b=��/W�M��nk@i8	�v��|a�3�X7���,M�Jy��j�˒��0X�����<�� ļGܛ`��r��4[���xV@������PQ�bŇ8�Z>��y�Dz-�?�xMz�z��C�>��,�6a��~�/_����/U	��>8.��|h���瑽ݶ�D�p��fH��ӈ,���z�Ђ�Z3��	�fO.�l"����� �9�e���2��L2����s��)�s�N�&O�^���𝯭�������A����,����=X�j�WKdoj����^��PS�t�g����	��t��GF0��"�Lֲ6,,E�A%p�+W���cHb7��4��ݡ+6�dm��㷁���0��+ա����$�o3�x�"����pP�K��m�?�K����B�+r�е���e���P`���
NlA���&̳�Ժ9�ڦ������4�F�@{-~0E��ib��-��	j3s���S�2wrCY�y����xQZ���/M�$�M%�3	���*�9;!��(V~�s4,Gm��L�����]/�h��h�_��Y�F�MUe�7Eh��5�Ԙ	��h�[_TD!l44���H��ggғı7��I;>�I^96y�ˈk���0��C_�E�T�)�>ft�S{�O��f�l����d,B��{?��*�87t�9����Y6_O��ܼq1�Ǌ���Ma�끷ۖ�j�I�^��p< ��@��L���}�l�ݟǀm{���ο��z> ����x�b�&�
;6gT8(�-���?u�_�tB|���e��0��6-$��������%vq��C4��tH�n����w�e�ݦ��_���HhW�-���z3��P��S���Q�q�y�~/�H��q2?C���<�L�p�Q�������'A
6�\�N�ur�g4J��]�^+�;v� Q��������#49.�:E�!��NڢX�K�Ex鮟�ױ�b�`�i�n��)�xW�G7y\p�7��\`�&�dϹ%��v��
d8��!���3!a���vj�+�)��"��Q5��⠛��jڢVO����C�;Nu��Q�&�wۮԟ�t��Ғ7��[ۅ�pf�4Y2�l�{�2��g�З���i�%-BH���Zt7��4��q6�g��9����������Ĕ�`6~@����]�6���]��
��w�}�[���5r�4��4t��W�]5���Aw�P^��u�[���Mb��!�ع�����?=��YXjC�Q�Ƣs�m��#�  ���{R�'2����"Ixo� bG��qJ/�a6�����4��{��n:���Ӽa*�',_���%�	o��_������d
p�G��3#nÿ�f��E0����~h����,|+��C�2����U�ɭ�dOw�ԲGz�g�/!_�*�M���"1��p觮'����@<��0��2���r����z9��V>|	Jp��)!-���t�eH_f�ji����r�;/d��|���Gk�]�O!y=�^3�5�}3+�Q�G��7�J����~��d�Es�żb�¥60���&����r���˝�{mn@
XQΥ(�Z���z��=�;���)�~�寽6ߎ���oU8���W��F���s��.j� P�0�Қ�:���Z��y�Ⱥ�o\	���Q.�#�h�IQ�	
?QNp���
��A�X'��?�6��2�D��$�\%�a���&z5�N��~�Γ��W��D┡��YU�$�	$��jd����{"�6�� �ȏ1�"�*����L�Is��B%d�.� ށ�Xӓr��Q�u��~�P�:耜�b-�v���>��1|��X��(�BE�u���/
��<g��mCP�3�2L����6Tb��4C��X=��ȉ��	��@����\�яN�к���
��Ĕ�:vMw�?��,����Sl1 Gk�J1�SE��[��7��
;G�Ylg��pd�)
@~c��O·�� �e�%���,�_�ߘꝾ��q�\��O���g(���O��1���g"w���CA\'+Ϻ>�P�֠7K���q�}O���|i��O�h�XD!!6�w뭕%�P���lqi�˵F��PM�O��?�8�2�	�/
�#m����)x���B��bǛ��f�S	�SR�D���I�U�5��ȳ8�M:{�����,/=��ZtE��wϵ$\(vo.�\3�50�(��d%n.�l���H����_0������yS�cL>���9�]�J���_$�n_�J� �g�V��ӥt�juX���[�Y<����&�}6U�Y��-�Pl
f�sJ���ή��8>��#��_�)s�_ZH��Ʋ��]�ny�#A�����Gg��7$kPr!s�	����ĚP_bs����J@ۖ�q��Z@g�Ce�X��d.�R���1�=i�qu��J1����je�#���q��xMQ��y{���P�Nݞ^�aF�SU� ��&�J�7v�ܵ�RѮS��=� ��<��Q<���M�	Mo �*#4Qk�Ɔ�Vq���6��rG��zL!P�>��S�WJ�0��������X��s,ӆgM�Q�r3�Z1i�#��H�p#�I4k�L[�0���UQ�7V��]�y�&,_J�4y�%Y'�܄�&uM�|��;�@���܂K��]z�r�K7�RC�4�͝񿳍�P�)�_���2�j3�����˙U�(����P�.\���\�ٌ�ꖹ瞂�v������K���V��)T�3��|�ӄMB�� ��;d������x�:I�f��	����4oƫ��YwۥV���k>���/�3r��+"��-k5�d���:��DC�˞���Sz2�%dȿ$�b�q�8&5���1�<8kܨ�t�*�_���z�(o�dWW�ftWj�k�|�u�vR����\b2���u�M����> 3
qF�`��������߅g3��K[߶�v�v�����	�1֖���5��fc0�q�R�B�ެ���Bf�Cβn}������!��< �O�ܙ2��*¿��{>&��Y#�I�Xp�7�j��UixX�M>��;��P�Ө i"�#��ǥg�
�M�;�)��]X���\QF��K:	�8�*�jT�ɍ�Er�f��o�������1�D�+b�n�*&�t��B��� ��W�� �ŀ��k�oP�$Ա���n�i�̷b�}i����S��B��r��u��=��~!�ӌ�h#�����[Y�ѧ���ʑ@���x�(����]	zh`�bT7$ϯְ�@��j���n.�����OKN�,n9�/ɠQ�R�@9�`����*������[�������'a۹
�ze�*����t܎W�M�����Z��b���yoȵH�IE��\��3�a|��KH�N���J�5:?E�70:��w�̛����WJ6	|Cy/R�xMO�:���N[h�"���۩8͕�=.o���,�:'��ō���Lʷ���w�f�3�!���L2H�+��q�C(q
��%����Ï�F���*�6�\�S���筕���P55��������x�(4쌼��RB��<�s^z;<5'A��ǻ-�LM�*���O����puRj�����Ϟ}9�|�p]|g|#q�d��(�Ap,C��i��DbN@c,��ٵ���8���ՇZ6E�� *��|ZQ���e.�T/�Bv��Mp�l�٘����ś�L-U��^�&g^y�1p�%մ��/�rߞ�$r&�hotW6�J�H�]/��;0��fd�#����Aj6%�qr[�/��<@�t���֟�W��BR8sg��p \��͝�`��3�����W�(�$�Uln�'�`x��Y9g�����S��С�a�u�̈́�<���7���4K�J6��q��a�c���n�B���\]H��X�7�+ܤF��ف�	���?|��Hz��O��]e���RR�eԗA>�� �-V
c �Ѡ� 	�򿽿���]��_����T��}Ђ��DCf?�%J�\�~�ވ�I���5+ �g�N]��c6�{��i�T5�.��(�Y��U-�\�ģ��
�^��:���Y�f������q����7�h]��¶��?�e�w��Tr�<9��l�#m���������};�`?�ا����;���c���C�IN�"X*���,��Ƒ��> Y�T=.����\Ɇ��I��F�t%��	g�v���{�g����ҝ9z>q�(/���3*��#}}/e�kV�W���s�ȳ�.��>�m�@�9�$�}#d��H:���ؼ��3Ř���.�>j� ���Z��%�UXg̬�yl��a0��x�WS��,ٶ^�ƒ�'�x%�В��'�r���&�lY��7�\.�9��)�����2�4�ˠ���6���Q����<'Tօ�Б13��tf���I�a�L(�J9��4c��ŔK�z�?Ԧl���V�ZD[��{�f�?].9�)McP��3e�}Tʊ)�����\i���qI��+�Y{�EF����!�l��BY,�#eϠ���̺��r+^���9Fd��h�% �^_���Pb
I�X�����ӑηI�2��vl� ��[k�6���iMu��M����ĦA�sM7��d��kG�c�@.z��>Gi���k����.HGJ�h�?�G�RF�mD04�afO�/l�p�������	��Z�a��*&��ق�g5�(��D����3l��X|k3�1^ }�����������7�_�\�J