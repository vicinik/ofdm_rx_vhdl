-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GBu/0ML7LsAVopSlTR0uKIdLCj4BHk+eLhKvFAdTiG8nFDvewxoj3pX9zzLE1fTMunkv0BP7NpOc
ePjWTSTwO/oXGBC5lvZs7rcMTxDYjQHXkalDbtjWNg8l8Z5nZQWb8XXwGKT+PY4I4jeM526UJq2D
smN/1p8y1oPr0TpEE1WLyEXryeOrSEeD2h/6XR+551uwsxXlIA7qapE8AWOUJP2tqKra8qnHoTGn
nP2IqqP3r/qhL7Sb/FSbV+ohyOJrzx4LWY3rNLPxqW6n4v4KBIfQRPh7uU0wijjqoJWMuDj45x4m
6BEdMd9RUpws4m310BCgah/OfUvbMwz2+frj1A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8544)
`protect data_block
l1AvIQEnZXS08QeFALL2GXAxBTUzv7sNUMwNrR/0ZV/OybY0p5Z+/cGJD5wI5lxRUx3u6Ixud2gG
TU27CRlkZHzoaPs7NuKiFNkBzqcj1silByaCrdCe/lG5c56bgNSCQKk7pkDWbQL4InNX2y4ySimV
pzxC32XhBlZa0HtXPcK1fKbpBqO9jLk0YkLrrWmASqyLfoCF2OeARkcCMwM2NoCfQfdnGQqAP9ce
UYmWKwEvYxKY+okFGXIsqMZprzjosRBbztCEZoBmGiC0mOX9uHLQrSHjfMmRVQlZx1KIGH6k9TKT
EAWm6sRduNa+BuIVgd8EFqGhXymIVXUA5/EvI/YdHfyxbsIa5FAtQt9U3YISbtmbiWpb2tJ7VsFQ
gt48lXY3OQxloj9imaYpu2wz9LTv5B/yGrlwqJQ4WZ/YXA3ydyNb125lvSYrA3ojvq2eK1Puq1jw
f5Wqfbmc7r5GqBJGz/xpiTDpfmRpUqsfOgtDNTFdc7GCV9tNFSgNImFsrqMfbWrtBOzcqB5x+BmQ
LNVH4Fo3uzlTc98rN9mbKY+8lUm6cyTlW+iAAqH8x6kt79rAg+npBjnbZrxckuc82tttvL6RwQiT
pfwqnaPsYG9Y8AwuvWZX/MX4KC+1j7YW/mzn10IvRLVgv4dc+pOXUcscDjup1HzkiYZSdRMCHqL4
LJ8bLsZsi19GVVrdqgoQxOXZD2R0WolLjiwkLMd0232h52FnNjWkgoDWD95MoCuaZWVw3/ZeKQcF
2duB3hq4BtZ0SIK11VefUsv69Dc4dr0nNiAi9rFcYOcZ5dR7qsNTuqNz7JiqN+7/GRQ+vLkCvYyt
Q8B7IZNVG0IlUdIY853F6gkzZDSoeuJFKQoFtOAFtWLm72VaXHvoAorc0YxfIJDQGS0oeiX7aWQr
TtDquOjBi2RpGX0TgLK6nxPHQwKWmNnqn8/t2U4dgwIfCxgyuDcR4qlRLYKkI9xxENjbL9EuGec8
PfwH96TLtAt/SWWvJ7jn2S+jzpH+i8k8poQHEFBdo+m9S3/rx/7Ez4HUNXxdqZqSWbYsu2PPDFLc
s781AfXg94ZjR6mC1+VU9UzEywLhPQjOCTfDgg+MtKq5eb5kQcjApGll6QvOOpNSfo/2EoBn8BwM
o3DWgE6cOz9Kdipb1juvGYRCAthblkcaffikUH+ZoFuN/6oKXA3lvj0XFxsewckD5izw1p9Rc2JK
Gop/bP6dluRxjXsTbo+esqhxQZdTyArkZvQTu+if9eoJV/ACMtnYRdPusxJcziksIV/QhqUlCN9x
u6rawz76EluSwWaqB9yEmTdV3Wk5RNYtsBPFGwZJq6v1KeQXOcU1EyCNg5FnY6r/8tqIbMVMThq7
P5OZrk/btn6I2rqi7aZyOZ9jf0BE0peiK2ymVptcAypwUIbuS2OOQPoVl4UPRwnUCA8ceJDls+qR
AGRJVdrPq+Z29cMlUByo0Qf0wWK6lmTFW07hn7YCDbhusBg8rn52Rfv+nPTxXJ2x+8UOCpdP6p8D
Y9nQC68cMK1/hXL+8DZIFIWqwGfL1B8CHNVi6Yw4DD1eA7neNtFYT0PwWJfCq7d/F5j+Z4uhEkW5
w+dI590t1CwTJz4pKY2gcnT6cZuXzB/29q28cF5p8+/y+BYi+8rgjy1fkW+lA7xEBqC0ks1uH0sW
ApMk4O9FZbdeQKOGeXtehGDJbYd2OidW1UnfIcK+qtTezWk1CVNrZum3/arr4fcEiTpcTIaKmoX/
8nNxopRHgRe3D4ImQQkT8Et5jwCsXZaeaY7h6Dgk5iJpkOrivUE8RG+xsWoUJ5JAVM4mHWMQM+sp
bbgzjY88e2gq2y/TOZrnsdrmhYLzq+ZMGLS1ajeQt3RLca/YqHgHF/v5Rd2fN0c+7PllZ/Uj4VI4
EDQVurRC9aFNEaquf3OsxsNguW8JfW6gSlWn5U341L5mwQN3sF/K9W9Gv48mA61f7NafV3wKVNku
RPFtMPXNKoz8/xqlJQPRxogPn+WBOofPC//7awNq4g/U5qZwBYEZZ2SYnpuepRI4BshB77hkeGeI
Oamkpc/BYEB5f0zvilZsRv3MmOHkB9WernVgimXYlDwQMuh2nBGeH34rd4BLKhrZTYB+0ky4NTva
GCDu9BdKrAvBMTmyZRluSf3IaPzaqD/cqVpQqyX+PNPIP6jaMnp8KxIPoh6tcXggxmp+rbwvy7Yv
DA7ror+D/OM3tSPCbVlRNhMf9kaASMBN3oCfArDh8IwfBZdM9u1NDeF0J6mP1EzprvMrqfh2Wrcg
gCXibhKxCIAUi47F81BJFuYp6pzIayI94+e1U/K8VIfKeS2rbiiTWvBZiMOsnc9MbPVUGqOjklby
3dRXMwv5jjXEpEe4Vb4VhVVoyRQTXeiHCG1QhQxTQyXJhuM5+x+rDjxco/p/Jw5i8KHrjppPJ87u
PE9S7CfW3sg8y0cDcdCMWE13a5a/tVHL7F6pCzWaMYKOjEvsXbPzEG7NgQbdcldeEKo7C+R7lSAv
jxj7FRPasfYpnyNQUyWWVyG/P0fqpPvAutiLr/kBObgVDGaAQqxr8eKFNAnmAwqTEL6PFfaJYhwZ
cGIAR/F/iOM3+9ZozSd3/FjJcsQsKfWPKYQZrE2p/pWiITkg+3LHvtrDapzbtGqLphbrLgMyREPX
E40aCWv7Zynv1Ny90AdfWHBUvQSbmEeJhULx98kyh9byKPy2PA5qmLv9zRTS/XtnvnInP7034/4Y
Y0ZzqSvDCKorCxU0d2KeYS0KBX6NGMBsC6KLk3ChR2hpKL8AQJDjolwXinRBox9oG+ZN7KofFn4B
HyA5dK4LMcuUoLtUprN1ErrZQFvdew3cG7PyEaIY3ZSOnhWxtyBmX0Vufef144djbCbWE+DorkH1
XK4IaGnGywZTKh0BXReKGNr8O7ycZvqCccPlBHHNL53HDnZVosaBvmRRcAoie8x4TpCeOS7pwnEw
U5Xnqw5OFFZqNFFMnllRJsbVTuqN9P+sDzKWkGVGIutZL37U4gXLMyMzHmc+b+PlM6OpqU9pYxvv
PQarMLyo9cn5Lqngo00ov62/Z6vq4SMkg2IBCTnaNaVvHplM0/4YTdmDD8wcG2tBnIEuH3K0hLKP
+cpkobFuG23d0WhkQzQelurfS84KxEcbNEvDbGHqMkT1Tb/czzJXI8Tfyf+gp5ExqQGD/KybbKOI
DpoZJsNvh2dI6vUoxxj7hmEeo8vPQJj7DhHAk2qEa8e6YMaK410q4At85e0z9d+bsPxpcGXyiRLd
EzOnuUgSAOoKqLSiLudpJzFHbCBfuDmYAdjg1moGMRbni6AAS3W2P051jBbnLymNyJu2Uj21hnY7
bDjeCbPSYM5BV/GjMuUmECxtlmWYQILbU6lvj4re532J3WLrVemRVGjfQrflAXL+VMBCPy5RNfkX
fyg6K5Z9F2Fc9vzZvGSiwgx3SdYT9Y073c7E+mVP+tXv2d/uPvEWPdEbV7iGbypz/CXBkmHSEEKr
pxN0c3rcgEod/Np3pXPPQw9BWxoLuZEGnKnjghVzSH37te0+chr4O/yNaij5b4brMZ53aU0tH2W/
kdYSEdMyrZW+7iBLw6BdrnwEWb0Tr1K9q2TdZ3t+WuOPQAJ5CIJ9bGSUPngxhrcTPNjod3f/hv51
6dq37XAun0cOjWPVOPM5VdvndgvaHMbnGX35iHhnmO3mLtu7fNvliP3e6Z+zPcOOBR+y13TA97fz
2osVKRef7rwXfliWfrYv8LJPX6OHT9x5iTdBv+H8cw6CzfyOeyPFvXVzIVOFTg/Kjp4NA1YKen2s
eAC5hm3Ku0z+qrYbBfksCD3ErnO6Do4W9tlh+Sz4vI9yf7j9rhwC78xU4HX5zLO1S336uMt8Ar7d
OkxRvjhI1OSylUxLMHIExC24/lfyBV/8OPlgrn4uhBeL0JYqigceN0mSeOCIDcqk8xJySTuLSqfX
rSgXineBkMH/pJPtyH8R4+YJlZlZKcEALccOCKaQt60KPVWe1uwczE3IKrHwxmVKQseQ/wNIHs2b
BkykJ1y1wQt1Db4TzbOcEIAuJk3MgqLpsoekTU/egImzO2dcplfI9s+gQW4J4LcavWGsjix8bV/O
tXWGcG1LDuJLlWUKSueXlP+alFwbmMcmQGtUPGxSbScowlY+eXPlZpxjJpkbkEnCxdw/BLI9tAzA
Q1JVQGrmI2E5RSbwsuXGggsHaFt7MO8XyxJEjoXc1P9nLdGYCGo3cfRBTH0flOn+Fm2fiq+xeJaZ
f1sPwwfcyOWvNhEq6maTjQsyWC9wE68gDt4CMnumIIDxwD3tIlMAxlc4T6blO172CTkMvrnI25Yr
fvjaULECr0w8oaJppPipF0JxbyQFeAYa/VLeVHnjVljL45Bfs/m0QZkBT49E+gzOdRfHBPDYx6u6
tDxmDYHw5PKmVLRDiW0zFhxjpMT7W78GAJLyfDlcBoY5UMj/uECiZlJf+j1Ba4dghx831RQxCG+5
+biFnLY8Pbn8OiEO0mYKPXfAxDLdvMaGf/Ax/9JFh9O/NEA/9SO94RtH30+7aoyZofm7Wz9/TR12
/chImTp55qWKH5lOeF3WIDSuCCkO6u2nDqC13/aIGr+ot4r8h2FV1/ZTmhxgLiUELhBEzCRY2x/h
K93qEUbUi2dY85Cuijp+EitsG9iwxfc2cQRez1b1JOmS5+KAtqh0Z+oejvh/KDwM/v81G10zgBY0
SxRCojHGgeaWdjgHPvmzCswiYt1gzjAsYNUr0CseJhhcpVyZAdkVl4sg7d9N4pEfvdZgVms6AW9Q
Pgda17hNK2yjhJSAjelBg7pJhenXD+ISODDJcrAYdm7vOXW7n1qfjvVVdEeuCjtTyQVw7wzaBD6X
IzaFam/PnTedlGINiufFndrkZIEL583D166IeafIin2M6DYnb5EhqDDMuphxrOpb9teOreKiqX0v
H1qysBNmPTYvGQHCrRR0rE2SKr3miTX/UeVEeetnMSwUI+yUYuBGmRzWzXUR05iPpkm+OoEk+T/5
hu6AyTLbKagAzT7R26lETeyW0MWG7R+gySjtCrWofhmGcPgYR2xT6U94GgnjEujtKK/hqepGLk4x
cvbq379/LbKhNrksBWwe3MPsfRDVRZwDqevVXXBqwo+3lOGNBkG1XekoCJ6UgtOz6G6KprsvmVj2
HVmkNOnYV69iTu5sQnDNa4/G3MYAGJXlyWcU+ej9a5fI8bLRSEyyGNw98KNuLQkltGJ/6GQ7U+ZE
AIf1C9mmkf0B9H4CU/NsjSlgX4t3R5XmcC/oo2v4HTCZb4LCWqD4Ao/sKLFHSI9wMr1Wu3ZzBwzN
P0wUEMF6MNCAlN2YsQ0Vo+2Vf40JcOEHKHGEkkqC6j+JSSPLUU+GovCJ3NZcB/wa0f974YNCg69/
ONTv0iMS1s5+iyLwADh/j9KpTI+NQNmpjmHAiR6cdNH0ph/6JXL1JqGgqZhy3rEN+myHYygThPtT
bILBBppU3ylgJTik+Ni68JuvVNAiHCqKTJsa3Rdqwy+i8osSoxDiUH/Ro3GdCIVw5gOmDp5RE8ep
QdOjjmASd/SOmbwdlZ9Iv6EETZlYCFKWYV52Mg131I8jcLGQPuWbsE5VbiksxYSbJR5YbFP1r3Ys
olnT+ciKFo1pGLeEBtp/TBb20BFNk+B0/5vkvE9eK6SehpN6ZvK5U5TnwzN20S6DG2hiCcFNIben
HKypg5djuyNZsh3sMac3KzBlOrTZ8ZXWhbqNFnjSZsOa40obFFFIR4/yNXw02olYDfysxU87QTLD
1IpvYFhwA3Vz3dwBlmiGWvY339NUGFSePY50Q7TE2X5jYfLBQcn5yXdGbML7sawvDgD2o2Hkg5ND
gISG9iN8w0NGoYdhLrmXFv+10yhMAkWPlhHk3qPXbHzXWUpn54vAjIw490BbVokNfyj3BhWmgz/3
FKHatbXUQgpqiuPFXkYONQSvrje/wPKgTLfggfobCscImS0mnuv0QM2Iwrv69pjifVm8ygqnFbHJ
hdQhdN9HFN8JAIl4mLt6ejcd7hRh0oXZX+YrAPCXivvHBFzgSWuJNAXcPxrVpNZv8ptOokAxoQHM
XH3WJG3pAFzMHbrJHO6MRJUE1KtbweGRWKVVyDfGDjPxm4rT6rIatkJeQx6uQrxAUxkU8LMp+oAq
SLylrlrEXLrx72ZII4GtusHVyLgBe2OMgfhr3zJYKyIQWS3SeUdWab+WnSLbrDZpshZT7uyV8IaF
ldKU12H0CYZfEhkJIhaD+mcKEDjpfdhL6XMt0+LEcpFyJ2fzt9BGKTZDf/ZL17e8pN7aPChkK8qZ
vZw1yH+7V4jGbsPRM2rNzx06XZRxP7Na7JA+RUpDHphFVengh7X2PlRBv8uyrP5yaIOCHVCNjlvO
u1Y6qX90nRO0Ibrlske+qWZAtV0o8Skl8CkZuSHxpW1oLZrn0XbDgGRLokSq2PGT4xQD1xW3Wac9
YjGiKflAi+gj3vTXW6le6LDQx+37shj9DmXVQrIOtSh59HxLauBMfJYuscfAa2Gr2G3762PCrVDJ
yNMtTKFBxVxQx2/Vk+vyHMjHyws+hFshXOPY9Wfd942ytxitRU6Pu0tXbgOjL45JsBbt5sBkH4/m
xMdX3q6BmivVaSL6CA6Jvt4FWQ3n/2zjwlUIeHNSVfsTttky2YMTTibnZbWloRt543ReHPviO469
g1Nt6o9lTK4k/IMLSm8YaUahCgpKd4TJvHDWRAn85PiVFal2DNFJnazrMzsNsB419Pcjq0UWjnEi
9oR9hT2LUonrfMfaWG7vtnN2wkQMb4PjnbpNNqZ9gFXB+WBhWANuPoaMEgrPz/5KD/yzFQFEEQsV
KvW7X3fLmwWyY8+szHzdDiK33aO7HL4PHeULJccc0EO4lyt53Tbk5v1gHkGEC0Ci/1jxMP314ZeY
l4pLf+iQkxgKtXq1ttnij4KcKcsowVSf9bJtO28vteo5FncSPOg6tlo5y+jVLRH4y511ZcDE6TmZ
/oFuoMd3ooU4yShcFgOrQRcg52wWdOBhQuqfKtmTe4URcAh28oUpdb7f7dG6MD8IyFXxk4BXnCqj
I0bbR/aFZjvxrrZTHPitmcHld1AZtMcuGF53i2VDhn9khVOpGJYdR18+ACA2LGLEumA/dKKVfd6Z
vRNR3GqiwBvqJydlSz84PBkZ3h/3c8PHKkgYO9piGzKkS5TzZGEtKO7V4O3st1zaVrDayoAne4Ev
lWzA2nky79kAVkKAIbG/x3giG+1cG2tahh4QSmyxdzsOnzg7z3fzDvSrvvb+PU8Gbt9aM8EvJ6F/
gwzK1bbWNbRo9LU0x74PvSQ5J/AVRQ67wXWLj2k68+6nRhzR0iu9jgysW5rOo+gqHV3/2nk94rMv
b4huqE8Kww+OaNViv3gIF0jrjLa7A13NuXC/ydHM8r7utuaNjxz7nJ1/3U+j+Ai/NHg0wnm9n2X0
yfLNIWWWg1XkdDtuA22cw7vW1c5Ymx35Orpgl2Skw6Ld1p1jRuC5O5ha/pbOwvnxQ30tyGAc4mco
7nnRCU7V82PS2dsuGi8FYzBiBMJMOUs3iMq60M9lucsltP185PsrvYX4hifdlONjfcuBgiVFzfsW
7ThVO9H9CTrWILJzt5F3VKvxRmSQ9VlGvJCaRl6KQ9B/6gjVJpgBFJW4ieMLhUycWiUm8jHbZIkF
k+zjAvg6eSOyD/RlIvbFTytTd78KcbMEnlbjA1Cy+YQ4244TtVeJGKNIt5X9s1/4jvfyY7x1bW77
mDeVRQT+EBxvifTe0ZPwzl1PYynTup79mJ/GMAIMvhSdUr1WsYAzK26b+iywTOgXIgInQEIz+/7e
t0k/TgLCW0M3JahFkKgASAjQ53gZrkH40Gk/PN8m0zphfE3mRHdOoWI5IZNSczL/dBBHfreznbId
+sSRyWAq1qDrP2swJT6Denug5w8bgXjBPOJZRWd0FcKD+0P82KMYa9zIeLcsCKude5sJuj48XMOs
zP6OE4nO1KMEgA1ZRcPWROc14KpVald3KYrSJzeiXFjsydGxXcrg4lf2/wWGsmVr6mU1ycpiUm6z
bRnYWw+Am2cYzlV93akfxE92ztpCT9j/Qg7nPErfGh3S/74uYDN8PDoHA5hnvxhJYdsi0pQ4Jmsb
W/+AseP4st+FEbNJvGC7jtTMiT8M0T3SZuvkcVuc6IXHDMF5m2ABG1k3RNUa/aTnxhk2+ZvVyqeU
P42v5qBWLzXB7LP92eEPA6AT4RUkBNQZpiwzoRg3eA7W6I5yS61bw7qjF/R+F/qlA8HTDBkd+KE8
GaIdrAVAmzoKCfdbvgVj0zbrwWyW+t7Wj/Viw0pAu6H3NdUozWvsPd+qhpcQ1snDFup4dPPB/0q7
BT/jCZ8T2g7y3RHB+vE6JL53WdZmFUN4xRyv8fA6kfR4qaxtNomgcwkFgUyTd/09VkB+KrbKWwN+
+bKyIuMJ5A6LsQ2Yv5u4UrG5I+N+a8E1kmN41AdOwtbQpI5zfb4EdqdWBj56S5wdtnbCE2LTdK0t
usRqjFcR5cLbjksid5xG7Ud3qT3xiUIv3jBnPTkJI1jydwm10vPaLXeAvsK+EIAXfmY/SQNth8Lt
H/sqBc3nv4PcLc1VIAP57c8xLvb7NWPVD7zvcYyOHNlHGU2OxNB8rz5k3kqI20sailHfiTtMwQaI
v+xKnp4oeeHEdkV4EtVx0AzcoGvUUZOh8WREFd0EOMAdl4k3/g3/lV5ZKw0Q6Q1+wxD/7q2+Ww3d
/bPm4/a0uJCyOMqe+ujc7p2b3MJykeiEtuo/K/x/ZcKm282sd/F8nozZWIIldfK9ABHb0VyvRGWM
1t35iOtpVHgKOvdxXPuxwwTQ7aRQaNJKvdgnF/2aXQGgGe/VKkintYH2FNHeDlmO9QZ8QcuwegWI
iGCgFjXIuNT4Kskc8lP+OwZ5Lg6Rmpd6SwG6BR1IqSX8bztqjcI7TgzUQ7C5IWh6914ei2nhCrU1
cnauQDDsKPJmPtSpk5hz9YR57X1OMP69Hpw8mNoRLZ0uJQgcJLN+6eeBXUJSk5YgL4icpSbw/DO/
z/lFq1Fa/j67VwATq085RFkBgaS+AXlyr8PrCwnMn4UFhm2GWG7yMwxgIBYtms9lwBV64OWw3vaO
8kCvQp3O0NzSZJdq5ec9vE5ENic+n8nzbFqwfHiqkMkuCmqouCS49LPX6TQ6pL32YdGx+lNzGlmB
Inh1kTxxcku24IqR+ic7aqmfTU9TBYmBReg+BsZtaO/PPa9zG0cO8WYd9QRX3qRmggbX+j7dahrH
u5tm6h4ZrdTeONIVwiooLPDwfpqRjWzTq6exJ6BGz5Jmhx1P8q7L9vsB5HwPWtZONzjK7pdyrB4u
P9b5fudpA+I1UghFElSN6SpXelmd7UbklyQhjcyhcFmBPNV1IpZ3L1XqknUZnjM0wdEmLCAnwLAP
KB+GneNtZ3zBVJpDJXj044gwj9qSaO7V0v3/RlkUL64sto7TSgkjn2zTSbZWUv5fr4kZZ8wiAwSv
ANOD6Jpnag/nHmbsY1lynUpptBCXp3eEgUONsjeqWZpfywKLPJyLokiuRVut6r7DxYJwyLFNQLcB
OF/bg3pda0V2MS4BBV2CPvf7lEeasm1PmBZ4MPYBA4N92aI0nfqV9LgbE3Sat9ByHCrOSxOyH13c
A69t8mpH3+dEG8hpTzE4l4zK0vrKhibQulj/YTp8X2xGmRcwhIJkc1p1dirbXvpt1RNDel1hXndO
MnGKFYT2064oYiQb7lgO3faI4MmClEZNcgZg5emSKQ883EnIyrZIvjzHSBoPFI+fgusirqJbuWJL
QGIQSEisBCDWRBxEObC/LgebmbQwyp1gONE39mFvVeDTG65dSlBpQ2HqtSXzfJDtDtPHetydftck
i98ZfUYCqcxeiZgxAjX5nWgTZT5ejXfW0sr8OXPandWNsXOT7J6lWWxOEWZefJjRDxBJensjbidi
J4uLH4TEc3uMKrX4Nc3z1Q+JEx2JNd5Oi4QSWGx6QfI7+38xe1n/9pfdgquPreMWhs0PeKcsDqWd
KUeVElEHPOJRHxv3H5a9BQTpogOQPlt1Y80T8Pa6pT5N8yNbXT5qPyJApNZos+TAMthW9V4QtU4Y
kdFqgB8CUnauTrerBS7PVM+8SA6sxMpmDNcwg061zfg4CkLAOpZavv2C4cEyqXq3fwSAqmAsOD0G
9TBox2y2CObNdbT5+GqIoTIX8zpuSAIJSNSkXR+occLiGPKVuRaVNGSpZzncs2WVmi6+15qo/Xn4
TQxsdqSZjh2TM3pVUoxoHFWINzYMbnJpIuaM/ydOcnQ5SgSOvR7/uPPE/FjlswCX6SxY2vL2697a
QOw346zaHQuOqsha13pUZlvocD0jkKqVIGqB7NCPqh0IG8VFbkf66UIgCe6rbHoQC0ay/dCiiUhK
dOL40hZbeKeoEKitriBgzKjqukTiQPN88VBytMK6mn0CZ4PMKC4NSL0G6efslhzqKQqy5Gc54pRB
DTUSlLZl5XRtOLuJfh3riIsNw9k2x4gauk4W9XrHPSw8oKjOPajr9BrCdQA+CUygVxC/AlwdqPbO
/XFgYSgZEDeO24jOWKCwVRjlKsn80AjWKmJzFb16xm/talWrR5xCY0HOh9WQK0wNbMg+SOeT5YEM
AJqZ+MbQFmTMaHPZmaVyd6RQEXDRb27KjfKkRfXOsOEUA+bjnSIMkSS5eo2g7uT99fEhGO7omdwG
DR4+2dFjNZWWeWM/47PmXojkJh/v1Bo7YFrOo2JLnu5GD9bFRd/ucHkd/NxUYfy4J/E6R71IbufC
EqtALjQrxB1AEZuN9T5WrqlmWuYhCVTmzSK0NFHtA6onFIJrMS5QPgVto8E2qaWvqfTgI0vO9b8r
LO6hUvZ2dQxy/3RSzgYYG1RERZQRa6YnXdMAU+JG2K427xJXRrQAO2vT/S9XHUr0VrK9AEEXONiH
EjNZTTJ8c5sQ8rb8U3jXBUacJEycYSveoq5rNlOzTpWFk5OneG/LVEXFlqZ6VxsBgym2ov/zwEYF
YuJ2HAwQM+iM+Jf0z9TdN6gnFQr8UwE9hVcXBZCsUDh+KD0Dbrbc3QGXRrhqTHstSFMHrxGaheuv
/2721kPsQPDQ5ZaOnPDxC7OUxKPDCE9B+0jV0xM8Gl5z0BPYOpfTWT/S9L2WiHX5jLWRRDRtaYf6
iKmtIafN8DszDM4ZggbmFqRNx+JqCAGB5Ev7qrJsjR0SwM3Ft/Xyf8lti1ipvbwy0i8aDcH6tbsB
rcV9Nds43LFogT1IN5h3z8gCYwFxrykCLydtoeibCspOnnSuXehUokamsYJs3mBDZqVQ6On4GB0d
QOherJiSX1T/PhXCWe7ZDLdzF5XzFuSbEW9fyv8cvgwV6HbqKoZLLA+dwlGMAw/fptvn
`protect end_protected
