-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sCdJF4IpceuASXZYcM8QBXjqa8qVPqER1uiq7JBMIuMgpk4hjMcUFAoM3qnURg1rERCSkehCZGul
h/KWVbsfmQK3ujNwaeil8/QMl9uO86flR7GtLdRotuhM38oHhPul4Stl0k29VN4RWi/VMtcWonkM
J/7ffNwCpcKlC+S1HY+z+9Cp89mdRHatKozrWBpnUYbzHxU2Xm7twKIkBNHhLqyoy8Jn1RdlRPnk
crdc1MdYW1uJXrS9pjsJR1ExQ7G5IjxTantMftGOCjzSgxT3UnlN+1JV3MQZaRfW+0BtokALaovF
EpfikpbBhXase2yXQIIKK7v2TgB1fWOsPEw2xg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13296)
`protect data_block
rhdsatOH0uJD+3FsHwsWfsohZxgr40jTCQxJptUq98fx1Ts/xZOg20t9BbBKrLMdkxeEVmEj+G6B
4WxSmH3OD+sviTK3n7a0pXjE6J0TgW7BI+oFWCCZxT8RH8sIKETKKUdWYkBDAhiS/+0s4/aor6MR
KLo6Ztm4UGHXxMp7g9Z5J+cJmfNMIu8T5fgG3AwaZjiloW2JH8NpqefMTLu8Lj91/OMbwb0XIxkZ
dC9qxHco+OjA2f30w6u3a+JWripEa3CzDKDB0sIPDeYkFDhMnhK9p7N+8bU87xx+5h3LC/HVxbjH
nn5813CBbt7VGvI45tL8AA2E+l2QMTfs6+pR/c6TDWCecOhfBSuuNykUbLfBARO8ZDDOvUxhfHq1
AmE59tF8iQsx+AouZ/IDVoPGw8feWP8sA6OCaYajYgDyuL3lEr81bbGl3k3KuOEdKXsvDwbxjlH/
hFFptFh0T+0FgxRs4a1ZwBA8THGcm9r236pgWAesAvRCIQ1qoHTFUZJczyioxWhT+4ORI4+4zDI+
W+1vjia2fFClnBhXASmG3PriN9lSaySBvuY7bYuI602wodbtHcV+dhozqxnKCkEiOpJzRrJbUrHK
P91BRQXs1KhG9TczcnQyS3Av0HHXBQl1XjVG+yrGv2bOno4klqf68+fpfqCZd6cCpe9IkAYmFKxP
64whiuAIrL3P6dIJ9mPoQVRsKbpudM48/xzYIEr9YwkTNg0bGkekGx01Br4SFG0NBDhZrvSaOoRF
df7jLVPDnTcK6N1j5FNzZCoslvtP7Gbf363w8UD7UKFL98h6FoUxd0IKV+5V0HTqs8ndYC0Qk02G
83SfkNxqVA/Tcl6aMTajW8A6oRACJ04WjRxnSvGAMVbokIsOvBCrU+2ntStcUivTOulbjvh/1/7W
zOLAaTU59uPAr3uvXA146V43xXUKGc2LIwz7IsBxsOLtkrFVBgcgMv2PTmRv5gieP00RIhKBF+VF
qMLQPnI6Wk6GaM0uAbl4qYaRfySu1OM7ci8nZT+uUjpQIQm0LArWlyfrpnmwJnxYHwY24Te6d8Gb
tYogK2tJavXo02SypV/oRKQ/KO/UUlYolLMTO3EWiuE81wPiPnBIaRZpb1KI3qRga471jozDxQhZ
frdO1vsdkIuFDObHzN6VmI50HP+tmZJHjwU/lz1RZuuMyeKWsn6LCthCg1ZydPKApTS0YTC4FqSs
LpzLRSeHoaoVGdqgPdz42xCt+UQbQZK9rX80haMj5QI2g8vap4D3lOOvokUqOl3Tqmx/2jUdiaby
h/7MG6CQvgz4tmN22OcCGH4RidKDCMin23z890z3qiXrDkD/dK3hIIzqwpr9dg1x4PM8DGCYQkpk
Rw5fp9J6bwOnDHoM2YspcdiwrUblPqKVvdi9WvWqtm7psdFNGbjPKxmaefROzqIbJ6ofrcGnG++B
a8yKPlIq5oPBJQ7HvnKMBP6NG9qHDup0SmPY3CprVXqxPd8WXz8AMR5FbZhiuOjM8BxmE6mdSKn8
AaXwlkodNWE24jioIoUjDvs+ogiXabw/Y0m1vESdRNs71iqjK3e11tHDGuLxxms4KErvff8/aM9g
adqoEZJQFKTksm97Wu49o0+1dE4sD6V9bMVNwaRm+Vp3wEnvAOmT9OcSOI8m6yASPZzWWt7aENkM
fvma6nH2axXuwenLpTCKeBJBQYftU1Fue6GQwph3nJhqgYX8jAmUXTymYwqAmGNxv8ygDu5SCjkm
6+bJykE9peHmgcPzYpJq4C6A/OVgTkCKyswmhhRcMwk4FuvYaSx68aIdQ+PcGG4+K0DdnAyr8G3I
6ifnvsuPbQrP8tOWI1gC4meFbNxLFrhmuZgs9jhe405P+SZaG9HTNa3honx25s1yqNV4dZt3iK68
GUMDM6A2BGT9HkN//dTtnLRqZeUsT0ClbJ+542LrZP4K0IpALf5kfMUP+2mMRZ6lsPNQQtPYKhwF
r9Y9vupekRgcK6ReAWV6VXW8VJoZg/NAGV6x0T6RqbyVYM3ApEVPNf4Dp3KEOwNSnmzriTyxT3Na
SXqOSBZaw202UOl5aJ0PNcB2RcIHF0qsVce8jVlj18QVxWLMkAMPvfVggO1dWQrReMaLfGUbmpAS
SMCxYNm5KupKuHMV+fryk+j4n5ria26PLJTWUipWdCEshnl8+2NdpnLCRzW1buIvrgIlb0Mvmn1L
yHzt6BJmpo/EbJAlgV2dEC5RrPKGXSqG39dr8n0fzHX4BxFMKRz0Jc4Jplmikomw8Upb7ix0iZIb
ZlSJz33B2l/Qbm/0quM/ZpAkwCP2+S1JP/DKpqr6/XJvewxu8LXWs3MrmP9DlIAin2mGyBJkFQcZ
P/blKvpVznglS9Qfaf9vOqbrRiFEX8w50XQToBmnNcIMp46E8jcxkagx5HDU8wJn2fNJKomGKS43
FESEiCwiEDsqRrHwZQlieDtzcOPmXxQq4I6EImZQ0qXElg2l4A6pbT3Uf0OlLyTHw1O/bcNgY2Bw
P7dyCe6k1fEWcGjbuwK5RcGK15oegHoi4XggKxrQQuyeKOunJXe6GiPxQW8qwKaUJj+M2xpDsepU
870e5TvCvuhDvFTlGWhw1o8v9Hw9Qve/YBISNE7hMYHFhmg5yWLna8eznQojBnrTXwujTbowNOGe
wjiG/5FKUQ5fv7Yz/2YZqOHaohUHCkM3xBDE0SnlPY+6QbqimH3u0/4esxtvRdHOm43Xy9dUWxEO
fNSv1Z9xGhE+SKBTooQPu9O0E+VGH6BQUnnmko51xoB0zX3JwsTxIrABMILsXsowjTv9RNhJ1WRC
+WJ62fX5IrnCUqFEbmX6wf6hE7sLtoDqjykmA1PXXwrRvJZf5zhHmWJ/Aswz8i+xwEQizNJlN4ll
kBJUQwIDmj1hcoJ1RUqUsLaTSz8uAQeGCG+BUgSniii04UGwOfc7DZwD1SEhh8PvuAmmkeCxhxJp
RwiQ7Qa0/uzsdrs/CiSp764/aa9B7fk8osmyzNqyBjSXfzfJaZZ2jPbxp5gt0pm92KiwMub6VDFp
up0NMg5EghU79cFb7/Mixub9l3NvAs4yUee6yTHI10ti+ldTKk5UYWIz9HK/bRMioTt4OLLThdM6
ZYaAUdbvV70KfJno7CODB1h8Jmibiv4xzWhI9Ykfcl8r+7ty8i9IeyZJQAFsdSyIQkpPVsOHo3Cr
Vtp28OjNEnU1vIwZMVnw4bRMjCyLtQptlz8t258EH/7T3o8J3vl6P5ep2ktnxrjRJXyz87gWVfX0
us6Lbw3AuHtYbujsosaqxyW31TG1fHcHTdsV6i1itWsMcqs+BL7wojsS0UPHW6UnL0hr3BNo31gW
bXntWda13p0wQdpkXlr0peDOJsq6iV+//8zQMxM9SqkNPTQNVa4rrTbGFjsMbUAw2aDpDH5gJ9y9
k3SIZpft0vDYLiMMQwQGVVzFQ54Lk+sQA1wFGmix8OqIo8HatTamiiMDDwDeyT+qCqtEdt7lnnVo
EWDXCedteG4afJbvrT+8jT029adcaWPUzI8zh40JaOJjJuh/js69vHyFJAlwi7TGc7bnWdAbVJRA
MA5go09BA6YE9ExZK12y3rV70ICYgykgw9tsb7q4kim6Y8oT4DRO6E0uhsM7YHH7wUdAdx6YbW2T
9TLzjYBLzwPoZ8ARyYGpuFQuZP9zVCD321v8slNv7IowObUIN3LDu47tTKfuYjHxMhnO9D9GpAi3
8Pi1e+VT+jLtsTjDw2H770glNbTbjt8fobEbzP85sHN/FL7wKsrggphaYaxcNFUsLMekiuk+3TQ+
MlvAdvlaqd4TlYjOFWsNYeRhoptQA2JvnVqGo82/0vLUlBg4s+IX4fO/dDyCBBp5O+GWa8RHB0fj
JJsSwdJ73Rm/uk4Xac/b8pZ+q54iWZZnVL12DI08Dht5FpROM7IHCu6Iws5c/ZLtEuh+CVmL1kLS
WnDYaOguQc7wceC5qkQpYZAVTQUh+pGJs+ye/zh/cMzXWZwXi2pGK5FGkRocWaUJgQdtpAAQPFNb
nhjClkmc6pqJ3HiKWWNM86XMN4F1KWGYCedJLGsH/+969DCKKlb+LxDXbC1PBYPIL8DDmsrVPGkO
m6whevD57BpVcY09E/k8fvbqYVuql0pGXmZFxGHH/aWOHSr6pJh7KgiKa4FokwMmDTilM/x3GLNw
7k0VFOBGX/IVlnk0pWBt4FTuigvhWQ9GELmWcCBrYWLSzwiMXY7LagwhQOqTwkGVdvJkzeJDos3J
h/g9LNC3Uu1Q6tnlFLtau2fhWRxKqRncJo+IYeeYdE3NPr39Iao5YjWAAYgwn12E5pvjvH20pbwf
b30V3KtqMZnJesfTGjnPWooobXlO50e1AgsYDv0pQNcEK4St+o7WhYhC93yL/GFZIryxa/ci+enM
K2Q19cxafUyZ0gG3n6K5eExhv0uTVBaCxuieguXDCRlmWdV50+0bMzFFNirE/b5J49JEfJJ7wweI
jRxrbhddMVGG0rb8csTzxs8Q/Pw31w/9HOvlNqWIqa6Eh3QtvUUfjMeF4WSQW/G7d9bcJ5Iy83pV
G48hGXrltHDBW95AoZDYmEiLpwmbbF3qHeCqxUYVsx+xQPMCOonsrPDlfrLhgdH8U6R2+poY5cMD
16c3B/3Pvy6fH+9o9In82AzyuKGb0lrSmhGO66phEFE9xdq9EDBJlc/KBJftZDa7LjmL+1ehn0RZ
SY2GuTMyVYLsbPFkLPZqdBQvCngBvsE/9RVukedwXJEG5XEriceyArJUiSLa0kaxPZpyNLF25qTh
0DkNVIK2Zkp9iT3OIQeaggVmHr3LuqzeUxpmKs/8MBdhdS2lveDQ9Csze4GUj9AfAxIiY80cKuDh
mywQlcCOnI327/esIofwkNuSTCbOGvgvi83snJidv+D+rOJhRInbB6SU0ufuJ6y2Ocm3R9ShCE34
ncMo3R7rG117dNrY76Q0TkufUWY2zIy7g5RVIhq/QofyQuALcz7T8x7Ot7HCjV4NVhDarrVJy8/J
Pm79wXWzUTZiLSMKKWBEtNsMaMzmPc4MLkvTvSy+drkWfKRP4i6Q3z+/5CruOPP8VOb7WNUs6s7J
RB+nzLQFlDR2497mKwkHqcSPRZOiN+intSUHtSVzPUYhlHF+aknXVJadjPrbD6bpK/OTlKrlU8hu
9rvEPcNLI45oI68TXzbpWc2YO1VzEwcw5CdHaeeGV0U7iUA5PPz8q6aG3QJySSmqmZmWL9OClFZ/
cDWRCgyxdxW2X0R6RslJ6WP488ba0wdzE0TM+kbgjbq+ftTdlx5K79VLY54M93+5fqpAEwQ3MlAI
Uap+uXfA29KCfTIotI6JaEc+MubTU4IKqpDtRzuhzxNYfLSLl0uIvsDQJGzqmdY33iVexut8bQwc
Cd4ZxGlDT6cXQDVqtsLdXavmmTekMEoyg71Cf2msdBKDLErjmtfInwE/laWo6uxEC+pAHxxTZezx
ocBVUrDpIbHT2kKgehlezzSEWM/iOgRjpwlx8JN/JwpzYTZzL4ecpYBQW+FJ151OJpzvSwQ8akCV
1xeDU9xKmQ3kGIb0Lzm+wPTbSlRbklsG+ffnStiODn5bEW+mAwJ6Hz++9ajD/HPJvpHFBM717iuk
P6gFy79ZNmw8PMb8/4gQaWYSWo5Lrihnj/UOf+a2K638+bAXgKKTrtYar2CIrhTYq4FOs3vuj2V3
s7hNm76Yx5NcQU120dVz37Du+krZlJGF9ZSdJTkCiGDajyJaNunuQCwU/rKyxJ7QhX1lL2sFByFk
aplIC+BS1VBmM0TV24aYKLWv7KvQ8YTMFOCNSTVmBmpUwLTCsZmVPfCWsiR57vdMf5feYO1NrG4a
uN2QIXlohWrId/8faGVl93u3VZ7G+BnU8VK/VGLsLcxFrWsh2JJgxd+CrnU6NPqhCFnR7cZXkEGS
dRx7qpvL8NbmnYVpvi5e66hCUOUDX9kjwubhi7fPGERq9MSfRtp5DMt7p7qA+rNSYyd9tn1npLoY
s0MN67KMmgyTRUfi2Dgq4HdiNczUGLe3NyxSdRjpJWjAacxHyDXQqyGn9jL53f65z3T8SgJITEAk
52qRdFtkrAZh2NIMKrA5GglLlTrzQcBWL9WLqR36iqFLKzAaQJeOC5b1W5U8IqDyxCbf0+DGjfl7
2M7b+iCMfNs4W9n1WMzbo0vmifM5il7Wrx7Dq38cBkQN7mNifOt/FSPSE+Gp8KCnmTQ6fZ5p9THR
xE7k48pezFZuyQ3Een2eLTpwJtAGWTPBUyVRfasJ3PjKWTVpPjHCJaOq6GB2msRS2YDkFMMjiG/j
c81oidJvAhNcFrdwqYAQOeIKES3Ndi6jdu3AJq2JvIQQQrLA3H2+TQ0nTM0HlaGlbimsy9T473Y5
aD4gHTzxcVcuYxEnd/MOzT/zpShXtTj4+n5w04cHmYj1QcZehzG91Ez+I2DXI8yxMotDMLabqIAC
qLyzXlbsHe2eLwSHSSvKwsUSG3mygRiikt3vbO/fPeSOZYbPrSgvBHMS5VN/Iw6Fpnglk0peuO28
Ez2puR+SVoipWCbfmM40aOFZrvLS5aatzwirq7l0W+fJQX9T/vrs3IjyB1YF2svNsuKpHorXv/bX
6A0C6a2PY0kZlAoQX8BhZvhUQOABYzIERydZ9AqlbVPqEJWuHChHsFmW/mzUzR0V/GOKtrrf3wWB
KWpTAhcXxYRYu2i40QmW1N71XsaKMFz8XQRN/Q0M6MH/PGotwna+w9TIT4vjAaRjPMFGruHdDjBA
DfuZRiiV1tml1mFIdfZ4K0rTUjbfNWtLCBHaNFQUroe7VEyBvTTLA1A5fE0lZoSFY+TbE5AC12Io
vildwV0kBM/bWeplg31YRT5O7b65AwsE5xAGRT28eHUAOvvlcbo7qauGroupvAmCRBXS7MMtCJir
hA7k+IlmsiU7vx7ufk4dRxlwlPl9+v5Pi8nO88YNCzFgIE58jqPowm6OCUYXU8KUFOVEjpVQe8XB
8xMKjJhGKZblbwxwVqncODnxQkg+1T/6Oq/4xE/JD7Aw3tapOMVoPMjfADgOSBNLNbwU9t+AI0g2
V/DpzPjMJ2iP1eUEvElm1o/P8mmLSAHNb8oLhQo9QHn+eF36rdvCtef44Qk/58thhGsMGIRC4sby
Ff1TJ0yJKkCVHvo+kNk6ByI8rLgxm/TuLf9dR2ZkS2YW08u6cF9QGPfUj2iDJNzLhW7gLA+1l0Lo
Q83oq6SjW1sR5mtMsqWDx4ySIysQdfrhmmt1tME4Pnm+QzmNv7B82st2i19OwQgH2+5ivxdO9ZBE
9aJzcC0H6/rDz4eUbVjsWL1/72BAR6idfPZC71zf8WHfv3SJ3/KyGaXN4nj3esICqew+lTjETcPz
oyMGNEbUjQD/BccUQkL64VU97GP1bV97ZkltH1JHpr6z3uq69EECaRf+jqP+4ZsSK8xRmNFabkTY
JYqHIy51UO6BtP/TdkWadYoUEwC8YUBIO6BzxNCg1Y/Fbg1u4a5h9j+xq7bN9eL+fPGyVbhUx0Bt
ixCiAiWv2jzwtVCdKBICXrNN2AS8xYIGqJrPuwiyxfvXRYocQAl88J0+86OUlOstM6QIXAeabB19
vwFvHiiDcUfHdVH4TjJUPe54fBtMOP8rQivtXzB7strtoKcsZf31H16jSDp3xWWrXCGyVwplfQUA
PWA9YR+zhXCDgMnDp3JnIlF3xkMXLgAlhi3bq4uaN5MhB54qtXQpaPeYJTZWd/HFlWDnbNQnsOJo
frMxqPZjyeg4ExeV3xfRW41l/bYW3yiWfYyRJGK2fyVj5Ov2dn5Z9mB7oGCNn3UuadX1r1Tgk0e6
vlrG1lV6H4m62/Ang72EoYitaFnD6mUwzpWX/gQM8seXu7W5hkIKuoCujIChHLk9Tdf0aDqz+pju
9ES/ZRlveQW3kaJbfcs1sfFrpyRYNMj8d1LMERkGhkOC4ElJ1BWJE7C9n+NED2Z9WppQ4Gpvi/B7
q6R1BalB03rx8gxGrlQ5kFNguXecF5bWTBrI7/zeRzErMk8GtWVPrYc9EJP8+A+paRisA8Tiur6E
azfnlmiAQMT5XOSSbc1CMT3ByO1hC//kgpcQJuRV3oJBe8v7tEqkZOxFaRX98fEcDitQD36Ctk4l
AcJT43SqFqYBUVTtPX8JfDDkV+XoXmeyHJUCdg8bPM61vWgpbZf6ay33vEamZ8hpKVu5//Npnu8v
5TRWOKOn8bB3nkhvpY4h4BsUUB5zpY9aNCAs+dQjFZR8CsfCO+YHEjd+KnjSmTKJ5aq6v41BZjx+
a5eQGvVgYswDiGPjbxN0HMiWr97LFlPobleNH3o/XPs5dmqiAfMNtPdyi3kLHv2HhndeNzWJwwso
qiG3xT3yXzkIkSgCsuKCmdpgYXiRzOST9FXWfB8n1Knp0o+LBLLpHHPn93jKXh5JaX3uDraBrPZE
cjo8Extp+j83I6lA4zXnJmKUHWDURsNLE+6p9MIczFSD3EXHlplHmlG41rwiwFBP3FVJ8PM3WPIo
amDxQu0WNY7WVSeT+FhNMULJpJdOhVxwGRD5DJd2bVLNsYqidiRPBrhmO/S0ddvzD+eDiOtwX+QO
7WVlXjMf6ajtRbvTQvqrPrRnXZwrEEtGoA/1PZ3hJwfQBhf4Na3DlBD9MprbGm9x0RLbzf2cJXhZ
64V7yvjiTaenLxsPBLEIlHcjHDMTvI7cPk1lksVzR5qsDkjNitrUiuzsQtlb7mDz+Uk7B6oaByDz
YLCiGMVGJpU9+7n8f/IDGjUpNvCTtzHR3t3hyMqZ1RSHYZlBy2A4fEEbVFgRnKsxEM6Q6pj4Ndcl
5WUVC7TLoqiWiCVnFJH+vf189n2brsSPgxghuGF/n2INfzfBk+24XflMu6jq73+jN24Z3RHGiTHc
hWxyC/6kYWrUvhYrtHlIlaUG4C06Y1Xf+s+cdeat0gILQ7l+FJnGPuHzrs2Xi6rWY0XimqDFrOR0
UC3nvgMId10/rlFAft7+Vu7/08086mkRcXTdTodC1C0O6NM51Ni9uAjED9Pvq4yvrYbJOVEi9U3S
nL4mfpemM5+TcSdN4Bnnrx7CVbcwGtETyMFeCp8ya6heTXCy9k1TkVDzZsAJBQlwLih+xwzfsv88
/gWAQC5TGKhCvUGpv0zdVUrsHfu1CLPWY2Z+inLPImQa2QRSMxBAB4hV2SEDfsB6kz3uTlriXV+U
a/LaLGuT4mF4qpGTcoabZNBqnag2QVG+m7gkcaWPqTJ0B9fdUec+6x5tV/0X70WUFiuslJgG2ouA
Uhzht8bJhXIg9/wTqfRKYVz2s3sW0fPRQTKRsn1hHzNa4o4/E4lfkk9eE480sQtZvNdaUXV0epJ1
BV3XpCjRmHYgo1ZyzBtbVtiUYOyhIPCzqxkq3OMHaV5xvGjRH2SHkfVJOTHlCibhPT/aly1k51Om
4RTE1009dvURbE1pwC2nxiYihAiUbjfIPno/x/Dqa+O9BW3Jo/1BtqJKYWMqkol2OKbGEoUNGj7o
w6fUUJarv8HO7zgh+LsdU8IG3pvuTeQb91fJVCjAOYJJvGKX4MRluFutUnpCU2p3VvmJNbc65FT1
0W50gBXf0iYHbB/EQp0XINNcYH+Rok+U9fZp0wtncpa5YlemCLAM8uSoPzSsBUF6TORonm66mYYW
f3wFn839tLlcUQ7fLvmAYhGZnGP5YgBE0bbMF+ZAJz0013C2k+SW1oVwfjbhSVmaX5JTELgY5z+G
HW3lCLtpL7EMHfbFNp7r1H+l8lgftgg1fo7Jlt3bn5IHJjvQ+Ke8Wo0dtMyW4hBNrKg9MvpiuXpp
AOLwhb3Mu7zviI0EZaza/wcqJiKnAV+QEDCRzC8NHLAxzz14ACVegDpNwIK4Gp6brRlkjJrOBytm
TLq3UklPkY7/bM9Qg66cTJfNTsOYuxnljmKInnMYifXplwksdTOX19LHeLub/7EDslJw1Giax7dU
b5BKhpRcKW4Yw2+1JsMGHE7Id6WpZuSUjlYNlsofAa0BSk0zoGjDWCpF5ZQa1EolkSEK24C1D/Qm
wrcOP4WOfrwYawYpZEurtJhoyAfIfOjgc97fMnFgIQq++Ct2orWd6ZtYx1fw/4PlAhxSLhltDetM
+gJob3wfRJBXeVGxXo/3eKy4XGdFHOcxM0Uvk5jAk/YXKeYvLDa87TDOBYgfFkFiO0eCIDPLYEj1
2hLdtDJQcpFDQ8PRlqyPzEFGqx16qG7eJBJB0OGxQC7Oi0Bt39UAaPXinbkyJVnX4FROcJGRecRH
t6z++g4k9iu1HlPrNFMzBNnGj5tvAVk4vN0mEU4zCM2d8GWfceyL7fSJOHeU07CZJ9yDH3Fg7gEu
xD1KpWOJJxylK0chFxSvniIL3aFnTMx7z6bkERvphyZZzTV8orxfidfp6PyZ2fsIdguTbp8QFWWN
ZYq2M+FRY1NLo0bleV/gsIi9vNVof0L8DWrca62XAV0UOogRHd/hzct7TrysHN+BcP4O4BctdGyj
qJeltFTA+yDVLOoB9NGji0HfdtnUIpmuvR8EIxE7aDe9na4iTe++lTf+432LuxtuMs3QTx0uqXBe
SsV21G3mURrEpCWvYvBw39ikJOMscSXKXOqweWecP0QKlxiKrqHm+GvOQRntLfQNGNbiYQyBqjh+
dPMDeqLRKPOKXDI+EW8ViempjmYmyQLrw6nZ8Z7Iqb3Rj2Xxf/lznXNzbspfG040Hsl3d9k2TBYZ
DIbamYO7m2/6tTjpVPR7bkkyv4I0Y2tQD4PDj6SDizZ3BxTRz/ZFIWHaqdwXKeJ06Ol+GVniJEqD
IZAzam2zb16wMYMIpxvd9OScQ7JkBhtDrVazf5YsHCkKZnQ1LPUrfUWV3xOE+tGMuMgm+2Tv93Pa
PJsuHFydeRAithPnHgzC9/ircATRNiihLkBIMCafhS0dcqMof/nRO/u2gOFrICEhmTOyUTDnW4oa
dYt57Sup5i177UHsiFQMQQXCimFD8ZYnflsHku93OX0KLSa2F+DoY5gZH1OpfEjqviokeeeoIY4x
GwG+QW6w1H87zskdAA4fOfVGvFBIBp0ZzQ2G8HbZwx7Z3LHXb+6R/WaokajGKQcM3qb5rKP6xvgI
SX6oQidVyc/EhaUnoUBf2OxO7ZvbJVW4GMlHVbEIdKypuu4N5ZYi/gH39XyQsnVxhKJUupxqSlWS
9BerXuY9o4bUaAH29unH+PDhw/YYQRLUo+A3VJ8kg4zJqZsztpDLU1kc5sS+h+NsKPuK8bqzdLHi
TewFuefxS6KcSfH49Wz4le2wR2PZUNQmzSkD0QMZ9t/Jl9PYS0RwNqTZ2vIVkF+4A0CvXOS/JaTX
r3BBWaYEMqI9GxGUNaO+3lt9PNnl7TK0xjB5Od0kP+1yxk4UJhbkO4DroyhIXwdLFOipFihcNveX
8boY3wQ4r2RqKxgke3/PYIFKBYQzgiSH+xTafWkY8z8jxBNSju26o/BZ/PyvCr8pY0J8ZuAlmDIF
zpxhUGS47q3NLJjDO3mLxFyXrVtMmJCsZ4/bkOvIyqVcVGuECsucDBRi5xOcod9t9kKu9lADnZkd
1r+p6BxEMx+qHBuIWG2+fGqXjkd21DxGEBV50H9xdeFZKkn53s3pVaD4YJMFz5PtjRXwqQ3/lQ7w
I1wjSTNL3voE2jaeDlI2LwWF7qi0421cVhS3gyVWylsTLKJ3c5Q2zH1NrQS/vvbx1BFRFZVDjUlA
eG+6oTrdadktA5hPEBPSCRQYzo3FHcvCqlHo4JnPpzg+ENkadBAb+y+GuOqSV4s6tBW53+BCaA2b
P8eKIkgaTI462ptNSITO5pICyKRhCEJ9YXRwH2aSBX0ZzRGlHi1IhaPU++2sWjZfcTMxHPfN7bdC
2JU6ArgmURFL1Nd+kHkfj3pxhS3Lz08c8MD6KBjLsCQQsYd4dVwJSYKsaOuUaI/Rq2AR3Hitsukz
RVYuhD9nYezSdJzfeU9peebwyYGTYoZCtYiYxoK6udN5Cl4go75FoL8MQQlna9OB2yLNh1Tjc5dy
anI3RmDeVXmZ5SdHiruemvUDbU8NPCg1AosESbesgKzY3yLUXQuFUigPSK88hpHXYbl07gFkhkn+
+5DIjGu45tQJRG0zSktYrixBcbJzqZfxBBv7tGj0DM7z88XoW5G/6+q331rtoCB8zMZWrOwdSgow
1yVuaLCLLlL8atKNynIlGEw5ERdLQQCbvJIdSMJY0HjFI+eMEWi+vTH4cphMKU6b8KFZ8G1SGCn0
2HzMafeTOF0DD/aNKloH7OAKcJHzdOxz+0TCyNACv24idakvkyOW04Kx6oc2dtVnHAKQ1ofgtz6U
vRb5/YvsWkNqFGcU6F+4NqKiLS6XiibUzdzCPPvHLUbI5daT72mFxQruicZkHq0MPLe1R2gjz/nh
zjydBxPFaGfj8h82xrgUVm9lHIEwDqT1jiRnctPxT1mhD2XWbOjhWrdO2BZIOaOxnhbPdtRKz/eW
8EqsHntHVfXqDwNr5j28H7brngVGYH4LvMaK7+V2bc4EDPIg538CSH4GDnmF2T63umTLr4teF6yg
dSeq+UoTi/4jWf6MX+agE/UQQDQYf6uICdVKszUQtUqFMe3M20Fjxsij4+maUfDhsdVPGQsdTz2B
ytwVt01L2kFwVRGR9+amA9N3EJhfa8eHwt2IDLcdzzVCn0Grce72CB5LQJ01OWJY76rEQLB7SJsK
bLwj4VgHGSrtYSFuzJxaSWOlatxrOiEFuFbSbFOHz7hCENkujPWyp7OCLPO5x3OY9FQK+UDzk00m
dyf6If0X0erzF0nY5R9inbBkkLYa786uHQ1/zsiILJAyovAPaE8PPj80aETp3FSb/PfNPzPn6Mqv
nVtdGf5sGLCc4zOwfzDhwnbYBGblQIPSh7gmZfojRhyd5/x72CqHouPkmhfna42Buvo/94K27Ay0
qFIPmDpfoxA0dU/WL/Th4P1Up06E3NLaR/mOeIs2BGaOuSwkEcHQDCI0423HKlSXQPYtSE046D6K
4M+P4kDtgSokINdtMjndenZW1XVdN7CxhMPbBuXqZxTG795CWbGHQ7LwOqkPCDHfQA7dmVL7rQoS
wZc3IUF7dQuzWO6RTF3MWnY9qAmYJay3aj0sTUZOOl8ymyUWC4BcrrwZMsqVia+dX4zbwUhQNk17
A/yxrx+C0g2OrYXd+8PgnHTrdBcxWZ/P+F+1Q5GAT6ePgdfu59vo2z64Za4qmpjr3RikJb19YYMb
k5AgEclCakkw5VhPdlmnW1hOLUHl48Qnj0+IoLOUV7E34/vupM6+OoY1y8U8jzxhcBDFHP2qZ0mV
qgKjquNbCfcE2vpF8rjqFLaC8P9M+Tp44llzjpZuDqXIdAOUmwtHYnwJF/EeWV43AGshTne4FdQB
83zCbzyKdpClJ5S2F/0a3ptHXMqxr5O8RUxg66RQdOKLpIYykYuFJ87vVlm9R3XpkD/4WpN0Z4mx
OshrERWp0zNZ+FTl1jmx58eKv/0KUWxpJFuoE/wMv8VBS9dQ06Pp9kox3jynOW5uAZJXnIRcGh+I
ARItz3J4OiGoiIyyyxRTZUS5vSq/2iRTvTOfQ473XbInNyjRziNDBBGBNrnQfQYi7v0325jLo3ae
Jy//UhHNrK8fSUvUGE18ydCzofqYEWWYxVev49rV3WEUJrZELviNxdc/xJiEP4i9SvXy16Wtk1u2
watu+G1RdKS1ZKhEaBRL7KG2jcGMdhDI4D0v9LBz41FWoz28O0yjM9ffIITwbTTAVEdRpvRLA43e
BbiFpcvLuvhPoQw9eLd7y+bUY5arZxxe6K4MNOjuItinV6u1gQHOarbJOdzqnOP1WScyYd/Pbefu
QGvwG+tdpDVMSIJQPlVz5Pu3Yo2wfr6Est3wWPJ+sl2a87FEcua2yxSNyKPnaag+HRKRWW5dqf4A
ROmU/4DbqQDVWwEe6ftKFw/xqlk6pJsskWlP20+zPxWO6WLnPQptqxYnJUeGaRYU46V/OgHMtzZP
14g+bObEgn4WLWKh62MM6vYiRgcE+Y+OH9uhkS8cenjj7z53H8Q9kfZzAPb7z271feDBX74EAvNq
iUn4wLVycUVVDkLVpYCiwWfwHbCNjUC2LSf1cBHd4ChW/7u+5m2UuccMMs6digfoIRGJm48d59A8
y2eJhCiHd4Hd5cX2790DheySBY/PkaQVNvFad49FuWMb1+3beJqxQ7q6IDRfArM93Vh6V0vHKM2N
Lq5+alMYqRCaUR4MhfnRhFwMjZwqvmf2unZBNQaIiz9xosFY2WRgwmeIGV/vRwbiIoQIki6DLmgo
rLWxsGkUUeFhZydoFhnZLWAenyW3pGGkI2d8fy5K87XEBsbsnFR5FJhYueyUJDm8hgNaGbRwU2uw
PzBYXCRTGtNoAqq3qPnK4/7agjC7sqq/CqOonJmTHpw+b7IwlKDvCshQmun8wHWqkIZwzeT2wM3h
AyqJmABXHkaR6Wua+a0s0Q/d+w0v9RqqhWHlXCTefElUlS8BnW2K6xEf005CETLNYcppq7qe6OXd
/I0uttwWM2YGK+M2aWjL3pCNcjOwJlpNgXkuD861qLZf42aCunj9QVjUimL6P9Zh7WUdQntp7NOW
dgwgLo+lQeL2MNlY/zCEI/uDwXpQ7xbHgGZr48fDtAx/s1cqqsMMUyPCV57KKcvCXoSc3I/jOyfx
8OUlp5s8GV2FLLYDb8LW7DBb9bex3mxu1c8WPD/lEw6xNfIpjFmLrlC6moo+8iCJVwFnOY3VPLSu
KzojSgxBkKvr8UxkwmMlW8J8x3NX8dev4ZPupy1gmz5fq/V89BloKcgCy6e5xJ+1M0gKLY5rWRUd
cPzVxFlJFO2yCQarY6OgiBL7k35Ypoyr6QbjQdekfLxT8IIgKdg33OXRGETaLtFfMN2jkg0Sbv73
w6ywccqDOjMptKJB56xIa+QtxlEO5S27B0eVIN0MgnrcLdNmZD5lZ0WepnZqiW6zuYKa24haSRbD
Akcx3SOcf7a/jrsv0lwZjsd/EF0miw6jEWzHxbAqfYJCekAGZ+XGE5GXXoKEu1hIUI8eVOmPlUHY
e8ZeWI3VRL405jbWngidc+yDS/Zr0PmxOPmrUO0lHLUhFCmpW/qb29sEWL1rxSGim7j67DUc8RIt
zUoyO5peuaYnmACBknvXH7k4Tq4SoFZnQwQtfGV0Jv9nneXR3Ayn27WtT+Sl2mvuSM8wEqrIgHdD
/ZJi08YZvWuey1HmS3bhki92aibQspVQgjWCi+3BP6IRO5xFSciX+as6THy3A/Pw6thklWfy/brq
NO0lsvIZzj6ewK4KtxNms5G2vXOsyNbGFJox7QxNDjG3/jCktZWXvAr2T2v87qpbbc2OWySRExby
h8Nvc37Y+/Jj4nE6qIU0mWV9l//FBxeR2CBFQabAJiRX0vrGTx74Tdizgo396nvJYZB9EsRS4N9M
MN6u9zUjGxfYR0KyBzHz7u4UsTHaqS2YL9ms3P+zA3UhZ0gzEIBvHXaGs9ZWKtAiZ+Jg+PZrt6kh
Y+PvS3H2HOEHEP8JD4lH/XctMUP30x/wWT4Nfy/drCzoZNsamRS9O0aLyfaAQa+XVuZDZFZ1hRaA
j/MyNxxX4XAoUF/Jdn1l47kbk3tlK5YZi8Eh0yCxySbOhtcqg3y9/9wQISjUQzzwO17ksa+2qqLi
f2u3mK15EZM/QxmhQRN6NUeDyO8NkQ9FtH5rxxyuLwCpVwRhDh6wd17qEodD+Z+u3jhOJfVUBmHA
WMX/FSpThrTtCcqv/ZRZpVjQ+wSCjhrQp+NMJHUXNaP7pekGA1vA8U2QSwu+Bj8aH5opg5AUdRB1
LmA3i+w8I15MOP0rm13tgy5Q3m0CD19zPnT3uP9fxtiAUu7wOJKNOro9cAkMSS8vHTn2rDJR8wUs
46IXdDJ8QlQL1hwo54oN76NlQ/kecDzUIIla66A4ikhp1Dm02VB8DzWLQIWcgnI6JbzuQqlT9iPd
Aygp+kqAjHEfWsE/B+ecTHGjImzTMPKJJE9XjEEfeko8iAdQkP8UtTrrJNuJa7wO1g2+qjnGgXHo
ZBP6CLgEiD1jhVjjw9A5jhCO1lIcl/wdVlcbCupPNGxawb+5QFbSs/5SxtfA6aYKhb1pEuftx9gM
y6bXrT4Az6GrH94EjJm9jZ65H9dOmm97DS2Lsw2RkRP5McANJ6p+j7PomarP9Ja4GfLtJaYibLv7
IZeMU/0fAodveIR0YXBaAn9W9Q/bQo9/UvGUQPAfmwtJfzMsX/t29xf5PLPKJhHN6dCrB1kxS6C4
iugNxA6mGOVy8ALK1lzAOF5y9qibOxiRoYh44OI/PgnenYQRew0o3EsVv3WwqSdTpWIOWQQoN6yJ
jIbq9G3xtue6axr76oZjF/YaTKpcryslaz0w3BJIAQ2ycAwr9sR0kfemmBjIO+J3mxT7Vp1Vc7jG
E5mGT8LwfCv61EblxgSFVSO4qcDiYBE1uUOH0ysRo9NPwwomlGZSv732ZpvzwT18ZAMutQZgGq2c
zUUEUWKABAhNAXfNk9HTkKFLQ6CL04h6xLCQuK40BEg8Z2Q+SYXtBPjFlQyB+Gtb9pVSYG22ilMk
VjvZMFcYOl9vUaUhxNaO8I+zwQTjymzCvfVlp4l2lqsjse0KbHq73Ts82weY8pLkwqQLGmKmCayC
zKcv6ChDdkSF0HqeHtB2SY8PZbOmG09/JL+AmKggKR0l6gJDE5G5wS3PuMNsqTok37hD0ypWDos/
CuNFjDBUidelE5IxKFP41scEW+Ys0el5nS9ovXyN269yFW+uG2RnivOfuyAMgAceRQiN+GRktMvc
ef4gLOsuh9XjMJl+xBIpF+kkNyFymF6fez2s0fDTl1bngV//6mGTU9whuXZ+evCsD2gsiGBqxQcI
HoHsgNio2Z5SLZ+9puEgg4M0DFatdjlyqW6px5PHWNKGZIdqrW2Jz1S0SMeMAihjHRzZlSEKveaT
fqn7dsgSrMVHMcU4MG/TYMfrWHC739Z2raHiAkp2iEyVrTiAb5XSTUlVBda6x82HeReofzYW8R5n
TMxvVOrpSI9GpLGBnWR8aGCY9mxX9pypLOhM/5/j6r6+54yIR9ae45pRmCw/d/jty/7fee7iLd8Z
6YL62tSYCBWMZhHP3Bl6rTIdTGYyeu4y4J3wCpfWDER6hwIzjYgq0WDBBNO04SSv/DpBoH5lUx2d
DQADOxx8rT+H7VqoX82KHdR/u7toeGogvDsEQDWtMQm0L+9/iqRsWea14ImsvgBXOC1+IZrZF3f+
eD/lcSUwYDGK+NP5c06YgW6feo+iliFs++DSe0zjrkiJIHw2rcw6zUMH3OabhZyGcFewbMLw1iEd
UYoH0Yp4MO/WGIwz/9za1F4rZH6scG4qAzlDpd2B8G0OPpXVGiXJRqAEmQ3CxSqQD9XN3qqr9Tqs
FlQH3LAfQFUuomQu5qUfYSLxPSEaCOavRpfoTcJ6atASEMTuSuMvzEqoWfdkBMolZM25Y86hnKPE
Wg06vaqihqo9WVd222BAin5pujsdcoOZRyEVsLIpXjzGCRbI9fYVgVnoTX3jtTpN3lKaMobWubXo
znt2sztf1SptjuypjjFRjCG/MbkDZ+O6T1UE7HaEqcpqtW+QOc5DAdLWxG6S9egn5G+CPOZXtmFs
1TohvHNOw77b9EIGKu6qyPEWfXNqnrFrlYHzBgDnITOP0sqOtoOaRfZ1yJxeJqFBZzNFC1EJ4IWz
4mxZ9tjCQS+DhhNxslN9
`protect end_protected
