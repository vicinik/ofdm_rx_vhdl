��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒�0G �q��4˵��G�?G�:��C�d|I<��H���=�[��o{D�����s��+m\��q�ɟ�C҅f=#�җ�^:l+K)ivH�!�ƕ��o�ϧ�ۥ��� �\6���V�GH�u֖ѓ��k�]G��������ߥ���=�s|Uo��ӆm���j��b��"l�W�I�h���J0����v��ʈ�'�3� ���2�{b,;�j�,e\����k�$�7�ADN�}��0�B��L��A�,�IZ�4"�������Ѕ��C�;Ml���Y��|�mԃ��k�I�V��ڼ�a��SB^b���(��yC�9��)�0t�tU:;6�'�ou�'5�;דk	���7-���ȪA�i�/��gRBf|��U������WI�w۠��ϼ�o ]!�6�0��cr}3�#�^��XP ����]�|����c�Шjĉ���y�|O���B&�d�̽��	tDj{d��~l�>�-���}�(P�Տ��c��L~BL�>Q ��!�(��0o�&1>�=��� >�\��wp�-"e\ĳ`>���[� ���$[,�93s�u4�#���Pc��+�1گ#t#�Bwwv�j��?��ehD��h�G�<��%l�]�xxOZk&{u���\��&� ���>!5�LUف"�*
�SM;�߰#��ǐ$�5�ך���mʱi^x2��g�"f\y�If���={�Rۑ�u��~�_�y�����g�%CRs�'��􈫄���`���m��E�J��AXs;�0��bf��>���'/PL���pω헀%����z���&��R�����a�ZD�j�Aϝ����Ώ��Ekh�~�<=^,�k��&�V�f� jc{�<���AԜz�/m�}#)�X�n�*U3RY���珗1��b9!��O�6,����,����#ڸk�<mڮ�5\�e�+X@�mz����C�{�>#SA�Xs�W1�Ɍy��	FVj�\~��<��b��\9a��s��E9;O�s~�Z�EoQ�� u":��A�R�a�S+j�X��ڽ�����v4lx`��ف���?Ei.�ξ؇9��OԺ4�j�iBW�n�`��l6�;��e����ȷ���>EL�����\^��,��L��%��0^��r]�|7�>���E0f��R��%^�\G��,O+l���.�6o�pQ3���O.g�e����:�$
V����f�g3�@�f��)o�;8J�)1�V�}Zȸ�\�9S�'|R��5fw.в�c�k�P0J<6l���'C��I͓��J�Z���	��aJ��2}
	V��d2P��5�@k�_�'��H�N�\Q��q*�����-���v�r<&�h	�g	��G@��|��	賰J��,��/��q��hl���z{j��V��1&0�zE!�|Ыiyl~c,OrS�d �-N��f�?��u�+_� �NMHX�}ȇA�Md�������������b@�3!Ǻ���SM�1-z���˨sXW����a���^��$��"T�xX9���;��߹�idh���}O!.� ޝ��䮽��I	ш�=}�2qEF��A�Io_�#J�.z�`y����{P�;����7̔�nR+.����۽�3-	���=�����m��^�l��f����Ot�R��T"�U� ���9�D�e��J�^Oh�����	�⠾��&��KN�v������Ž�/RyK�
�x�W���D;,�}�\�64AR�j����)^Z�Jq���ޛ��=a���N@�]��͜�УNe헽�F�	��}HখI)?1���j:�*�s0R}h�n���.E�o������.�@���* <v�n�7�q	d�Z�£�*R�)��Z2��Ɠ IR��S����y`��v�s��s�m�.ܫL�A<���m� c���^��[X�*S�ÁӬ縂2��uF�҃s#~�v���N��\�=�UG:�z�RQ:��+�Z�K��v�-t�9.#��l��0�ï��$vm��L-����U�cj����Fp��&O'j���>��x��ƕb�6����C���>�
��I�$�Ȼ�?���~ ��wEGmё8�����Kmv_4v���M#}c�U1y��N\٪�!��!A����t��1>�>�?Z�g�y_��
90�a����5���C�Xߜ�����	������|xѡ�����zp�1��/>���O���ef]��1ҭ4`YkPzI��aE%���(�e#�7�`�M�m�ޔ�s�4�{���T[UV��b�%��J�OS��Tns���Y�Y�;A-�e˓�S3�T�-�N�qy�I_4G����A����Կ0y��F8.{#.�� ?^���6�Xe�����C�)�����hQa"�2$$���,N��v�����g_8�O+g��Qbͨl$0qi�Fʁ�)�pF��JMαF��8�H+����N�(r{}_�F���1�g��k��~#:��	�/|���/��'M�4_�6�|3?-����v��/���9K�3U0�f�D	ʐ{x��y..�w��0)P�LQc#|D�p���kv�QH\�bV0~`��o��CX��u�#���8�YW��Ѱ6ѕ���XT�(44G��bF�1#�$�qJBձ'���4M��r1�G��L�j�B#��L��fH��빦z"d[O�����H�wN�/O�y�sTn342iT\�t`��x�r��v���W97��9#Z�B~�B?5� �|3Q�֏�����D�ZC���7�~�kM�qa64�J�(ȧO#{󷪁�T��
�-�ƥM5-~C��c�Wd�YD�����DϦ)�����̩#塒��Ø�QBM@
��9J�5�rBS?� ��B��kO-��3u11���"f��	���ɣJ��?�Ƭ�%?Ou��q�d���(V���/F�;D�`�8� >M���Tۓ�>�(U�&���Eؓ�?�N���Hq�hr�z���&���%k�%�$M	��o.L��{���I������s����SU�g�Da�x�9F�����;�1���I��Wu��7,d���GM���]�ǿ�c�l���m8�*٥^�w/���v'��wvw,o�a�����+��=�S���^���-孯�K+�&��+���6��D:ZIf ��61=���̷K-���H�a��^J�W0|sd��?�|&��/[�P�!� @��5��ک���J:���Ȩj��*k=���i�B�R�����si���B_�;є֗2�]�|G��v+۪#?`!��ߦ�dB)�9�)M��(?/Ě�^;�W�U�u���aT����״�H�����G+�o��g
r���	 �4c	�8_�>��.�Ƌk�;��=�;�8cY�˨�.0�E���7������]*�u��'9�c��"�;�Y��{�c��$L�;%�H¯4�fl.7u푥��ˎ���u:�Z.{�R̳e#Y(�������F��%u���"G�:�Q���|(;>�t%�7����o�їJ"$�C;���q&�3���� �R6�e��	�.B)ٰ�J���\~��ц��E�'��?� ���F�N_� ��V�����2{ࣸF<γ�B�h�` co�.�`�)��9��2O�������F`�^i ��u���B���i/uAzo��K%e�t]��դ����wo 0�}8M�īp�t~���pVn�i�[���3�(��36��~Y#���l~d1�eލ��E��q4z�0�iȎ�?J32��o��X,O����"�bH2�X�¦x��,Y�
`k͏�z�eo�<�p�'�M��������K�5�7�p�
��[�@�%���S�H���'��)ԯ�a#���#�ޙԼm��'�SEe��Wz�X�7�#0FP����߶�C@��%���sݫ�	i��د��҅��(��wQ T�w:,|����aX-A#+l< �$Qa�8���Z=�J$�\�K]�c���	<n��ҋ<L�Bjk��X�Hj�}���`!ĕ�g%�5�M\��a{�å�о�������3�û<�Y����B	@lg�[ї�I�e�.��8�X� z|@�],op�����̏������@����'�7�f��fW-���!�{���#� x#�ql����T;��l�(2�R�T�WS���d �2�Y�q3.�3�W�b������Do���t�Ћ���xJ������~��`a��}��my,�3.��<����þ.N~}�F�=1v������[�C�1��NPT��`�����3���rK\&��.�!w����7 ��_��[�`RQȓj��9��>G����>C/iIԽT��L��p�O K���|h�h�o������B��g��|��b"-�݈��5�\�������B���ȧ}^a�L�D�Z��|�:k��y]2�p�fG�CY�m�@��Jû��0O|O� �@�tb�^�&��t�=<^M�WԃŎַ[H�N���b�����ax�n� ����)��X�*JXD�h��6��4��,;��Ϙ�)������[r�T�-wV2xA���p���pT[n��WF4y�T��IW�Zo���l����M'.p=��KJ�{���/�-W�����냠7Gk��C�RS��"���b������0��������˷ �)1
�@�Ɓ��v�t�(�6}�og!��ٯ�� [��*R�C:�>nZ���ܪ�~���-ހ�*xK�__�2�S�lpvE�jo��[.�5u��YR������+iN�S�#�5���N���Er_G��(8�� J$P�)�����-��8�O�-Wr�+�����Lܬп��RƓ�8DZY��]�; 
k�W^�?�i�kf�M>s�(�x��{Ʉ�/��lm���{��x[9 '��w���?th;���2�e�IY���y�c���D9㽬��a�"�0<�W�j������P�\|�MJ
��,d����ڻ��_����Ë��j?xAE<��U��oL�u��Z��<im]�+�Il�(�PܭU��r�}i��gϮ.�L�Ϙ%����9�9q�YH��iò�h�����.�$���=��·�r�u��<m��݁Z=b��QC3i�/��X"E�h����W�t �s��̰G�\Vl���i3+%Ds;���ޫ}0M	�jWࣚ�=!k)�놠�E�G��j7���jGFXm5<+:зm�=�֓��AO<�o>m��KCU@A*��g�9Y �m|��B:5B�z� �7��v���Y�ӿ��+h��o�)ܶp*���D�'Ǹw;�'i�bV�=�z/��d\<=���1�}s&.b��9C�c���!F����2zvړXӁ%ߖ ��",$����w)������4��<k~��.��|b�b,a�s�U���4f��?��Ê֖�T�������צ&r��υ9>M#��RH�;�ڗ�6�H���;����N�^�0&�`�~�;��S�u1G��s���2�-�\ٲJi�� �0������v=%0�����T�>J��Sqi��T�&t��Zr�����o6"s.���P�AC=�B���_zƔ�3�`"����S�=��}Y��ƥ܄����Jd~P���IH'}{�ǈ�6�yR��5�r��t�#ʒA�ŘD��#iIk{a�D�q��=��*H~u�Lf���w}���I�_�pGՒ�n��l��9ɟnRs�}�Yr�˳�͋I���n����|!���t;*�i�y�;Bw�B���N��p-����rE��Ds��q�}�G��)�e?��L��9�P����n	���v~	���=�z�=Wk:6�_W�%Y~TyD�f�=��B"V�	^Ժ�5B�G����-b,SI'yh�{u����7�Qec5R{f�i�l����
�FC����}�\g}h�/���ro�� �[��ff@=#8�T�j�#ʛ���-�
Zc���
ǒ;s�)	��I�+���� ����ʁ�����~u�'^P��&��u1�e���L�Ȕ{�2t��a7A�,�=c`z��y�"�/��ȩ�2���Z�Gŉ(���Y�x�O���������>!���P�s5�ep6���G`PU����e�m�}���9r|;�4y��jʶ�kL�>��*�w������ǛWJ��2#H`��=�\tVR>��1Q�¿�RY�����ȹ k��-�����p�R��,pF$_�_��/Ӹ�ˣ��0�\4��"��ra�˚5W�l�!J��Ԩ�~�?�*z�=k�P��}��BS�LٷZ��pM�e�s�^��|/,a~#۴�83�)�(����;�-��P�_>o�`�bAFY����8u���ZW6[v��܍��*|YS4x��@�F�aP�^;ȳl!���Nvc�q&��n�������	$�I�6tM�ə*�@9n9�st]�A�i��Fi
��Et���:�-�G��O[)?��4��7�Ȑ�ΑM�<	���_��\��:�8��^4t[^��z>?-Hz\zR���F*׆@'w�ְ���p[/dXLBQqH�H Nu�}���!�Fo�{���m[�n�.�a�1��؍]�%������4k��a�|Ӟ
���Rt�]0??Qy{�,8�:�c1������F��5.h��c;���k(߹��ct�W̟Зפ�ތ=)UL�S<����!��G�%�=��*p-�uߙ�X��3�ZǏg`+B��n�7��FS�����=ϼԤ��,p�8���\
�G��Rޞ�g�C��o���${�rDN�M{�u`�w0���{ѐ�DWh�,̓Ƭ����nHW��}�@�|��n���X�H���.�!`���p�=�+�hl�j��/� �%J\/��HR��˾��	�$�=���"�0��w�X�t�ʀ㐷���<e"P�]X���[�/�jZ����<=������w� ��j���K���VP�	l��:޿�p��%�E���s�R@;�h+CIȉ��Co9]��E���V�ķ���[)���������E��;��W��b�=������>=^$a�^u2at.*ɦ�J�rs�֦�Q��s��������͌�$�Y��Gb`��3�6I���W��I w���%�Č%k����-�?��3������O�J���J�+�J���&τ`�:ym)Qɮ�-箲y�󓴨�T�;r�������
H�yυ���'�g���ē!Y�x�n��=��k��xv�����#���̎�"�pd�s�3�X~�>mΞQx䴂 9g��3���2�y�n�=	�)�����kۉ1Ęs��ٯ�F���b�Q�NL��H?N��k�J��@�1N�6��,��o<�p3�����BM�G´I�OȐvE����4��:&*H-���)��a���6�D�zN�5�����EWؠ٤�Iޘ�0���� !�uv9������y�}˕P�"V�V��΀L�ʿk�ѐhH��k\!����1)j(�d������3*�����*mM��D (�,)�x�R���vw�"�x���$hѷ=F,h��yU}w5�F��Z
VJ�w<�2ŚA��'���m��hJ����i�5�>�47IH	��	�2�z��<NuW�?���̔�%�F.	|m/�+29k�g��k�s"5�m�U����7{��->�#�#^�q,��|C�.9`T�Y���V@:)���6:i�i��j��.�5���G��`���k2��z6�!�}�>�V�H�B�N�í�'���Ŗ����*X�p�F��ӠZc��f�1�<����g�XID�{� OBп!�>`�?�Q|fz��h���I_�^�p��-=7 �N��3���n�>Xo#�캀��5��\�+U�-@��I�h�&�B��8����\��ޅ:Ľ���B����}�0�T 1L2���/B�I��F8r���KiG�a����l��"���kd���Fa@Ȧ�������T��ji��Eh'O�8�:�Z0=G����f����p��iX�>U���)��z�Z��EZ0�#iJ/Ix ?>�]qص�GG0d�OO]����7@�Tݳ�{���d"#=��� W��]�)Άy��>��_�n�	��h��#"�x暻a6+��Ѣ8s�l�A�:tD�(���S��vLO�Zy�Ej�s2����rP�e
	5��|�A��2k`mEQ�nU�?�A3���T��r��д]X�@��f+�G�r;���?ѭ�񙅭���II�4�c���A��*�{xI�9�H\a�I����$���|�	�U����:���[=sX���ޏ�����Cx϶��9/����0TT�8��GW�����j����nO���z �[�f�o����t��ϱ4�ԀAə�h�E�uT�����~ِ�o�K���-U)y�i�X�r~4_������J���1���8n��
����=s�[2�w1�

��X����U6I�Z;^�VN��7^���p�)�3m����t�2���?�|~��S��ue=�]dY�C� �+�]�'���n(���;�j#���ʋ��$�5i\�Wf� \1���%M3�z���H���Q,j'q�ѐ�|�U���-F��p��we�!�lLϣ�Ӵ�{-��۲��f�����>4q\��50�����r8�6�ԤSOE{��������p���KeZ��4!&5��!Fb<T�<P�zhg���;,��,���>k�Z�&�?����:����~�UĹ]:+i�yN_�v"1��.�Wet<�"�c��iQ6�ބ~0}X�@ؿS 	N~��d�����G�O�y�|���_�ڪ�c֑i=z���&z�J@�\�n�����c*�&&�E��(CG���*�E,��D����Q�E>:2��yњaC
ڊwH޲��"��Hfw)�
� �L�z\֝�5�"�.�lDA�I�/R0'�@���Т���Ve��3�`�쾛5���QT��j�џ�$e[����wߺ�+��R�˔�8�C�����ni�߇	�W.�U����e��_q�Ks�*�]�M#*�=R�cJ������~ 0-�W��!S��>
��C�U�ŮבO��*���f��E�!�ˏ�-��]��J�xDCyB���%�CD�\Ń�G]��3hm���.�W*rM�Dۥ	=-�Ch���ԓ�ШK�X�a1����Xr����OTz�n�)L�nW���.G�XY�B�#`e[�Y�1m�.��Dz8���Wl�ѨO,�\�Åpca�Vs�ź(X���ռ!Z�E�V��+����ʃ#&��~���Z��CWB�Ғ��ɞr�&7���Y鶎�`�R���'
�+ e���-�0b�rm>&���$ߵ�����%�:9u�6O)8�U�ݺ�џ}ރ�/�`����ڼ��W�z�d�~�c��sy�J\\��#�����u�'D'⫕��"(4�1���aɤ�g=���vh�Ϯe�a�Oγm2��Ԃi�/�����]���\@K����� ux�˗�����Pd�^�Ho%x�4�"�����eT�c�H�p=�
�z�R5˄�˦`�lܓ遌��(3zߩ�.�����+�s�B ��Ӌ��E��s��3?�X�:����� �Ҁ���F�ʺ�>�y[��(aX�����ǐ��ػT�N�.�Y�c1zv@���	Ƶ����Q����m�8rV�2X���ca�Η\?�9�V�S+�)m��6����t���r**:�`9y�s�(:�j�CD�niu�Z�8��P�1�.'�5�1���C�d��r[��(Ÿ��f{��8��g��+���W~�򀁾��1�RU{�B�N�l>����T�8�ȽF�d�n���Ս@�^�X����ߛ"0�D��IK�gWEè�Nl�g���I���L�
e�T����#��H24q���Z�ni��N��)�vZK>{��<
�C���}f��d5M��)��i����!���	ƕ@ڮ�a�f��]���6"�Di�*��%�4����b2j	�1��He��6j2��e$��>���߇��P��M���k�y�nW��1tZQ󆸚��������d5��O��#�?u6}e)�!�`#���4~ �r��/*���25����=�K ��X�{MSH��2xRQ�A���������W��n���opݜ�8;ii3ӛ��s����ig0��d���~���VY��5����U	� }ٿ�͓���u�����(�ʽǂ~�jJbY����>���1������*��)89L�H�c�?�C�)���0���[j�g�G��8L)/���U�Z�2�{��rŻm�[1ot7��z!��<E�{�CN��c�{x5�!o,g�s�V�Ӷ���0���,�F����j�N��W�!��102"BI��F��B��Z��T��aR���+S7�	��AD��+���~���� �<����[2�Jl��90�ߥ���nJb�5�V�{}�[��鋚{1Ӑ�N4�e�4���P����L�H����+��y�y#��.Kr8�@�����-�L��d�då�e�:z����$;�ԥ��1@��M��y��Ldd�?���t��2=62�	L �hJ�֧�#A
��݁��'�Ij��A�Ȓ���cK�B�����f�������t��#FH��R���1J�/,���ך9��>v�|\Э�s�![��O!ƣ�1���ȗ ���עзA�=�HZ^b�c164�ٓ�.?;�R1b��]' ������1K���vD���x���}U���/8�Qc1����
=D��;-AւB�?��?�hhF��dJ��F���R�yU���j5�$�1�8��8�3ԩ���#����O �b�!�H<6�� �ʠ�ί ?(�nngޖk��0��Z�k�K/�|ރ%���|� �S��j�e`D��ԧ;Ye	�v�k��I����a �?�u��,����kX��>�>�A!/�����fD��77ީq�s���Nܞ����_�x�A1P,�M��Zf f�(Dߋ��Í	z�/Ѕ��6��ׇJŏ=�����,d�@�7e�{����Wʩ^�ky���`�6��r�%��aZ�}
�&N�__�O�J�6!�r��}�m�*�-$���3�2��ߚ���"��#26�"���f���'@�Vh<P�ف^��x)'�`�U�\E7�Z<do���e�Y�L��A��!s]c#���e+ҏ'�5"���ܢ(y�jG�߫��D�Bߏs��y7ò��m�I"ݽV �>�6o�X
g+��G(���w8��{K%�#ҫ�79is��`N/����l��Vn�?^>�4�%t�Ŭӏ�4}�"�
͞xTza>�%0s�#G��N_�§Bu~ƿ�x���KF�Z-�H?��o��*-+��`���lOIrWZf���J��le��T���5+y�iZY���j���9���I���2�-d�N��zk7Q2�/����
�H�^V$p3~�d�(�+x���K��K[�R������F�1�c��i���,���Z��9����{g61��:�_�.�� -i��إ[œh-��o��U���@E2ICI�x,���h{�0����c���ww�Qt�|�m��ȟ�JD������W.f�C4��{ķ�{0�G���h_�i}Y����Z,6߮�ɽ�y��)�����W��Q<�`��*��� ��<���W���&A���7h� ����
���$:����K%8��.<��]I��ob�	#h�YYgl�4r�U8�c��ëڎ~�Nwf�Kv'��f�B��<�e�@
N]V�����3+��c8��E��v�}��x��p�t1��8-ъ�^3��Bn�"��R����vo�}�T_�M�{�YI%I���.�w~�.vĖ��3��q�B*�O�w[������aF��~�Rڶ(�;y4�*M7	�͕�b���x�4��k�\��t.��)|Ul���t}����\ܲT(��O;��.�d��E�(��9EqoFB���'�2�c���u��J�Z��V���M����@��"�w/^�5�}&�+������M���@u5[9�-�jrs��G�E*'(=��D������1�8& ��8%��s�;�!�ћ�'�I��S�|5EiV[8�j��"�])5�0�/��t�.�0ň�u�؄��Q��|�f�0"�'}�!�V�\�{-�_ wӾY('����+i�jK� �ٖ���0C�-���>�D�±\iɐ~���
������O8�����\�������M���ZV��)}��f6�?�k�J�B�ٰ�:*�J�
���_%��Ϩs���h�O�ƕmmJQ��+b�%Gφ���uk����mP��j��N!k7X�Ss �"�O���m���f�^��6�,�謨�s="�B�����H����x��'c{v�
�N+I��\z\A��0?v�ns��F'���"����L��Q�$�\�_ۉ©��������䑃dg��C*�3��\����u\�$����s/N�u�y�v�]��y~���"�K?_:C����xc*��o:��m4��*)�5qo�#:,��?�����	w���� �X����L<I	E��7݀.�zZ� U�T��.#ָ�M��})����:���{���;��_��5�t}����b�78?�Bێ�=~#����r'��~{hD���^}����p�cq4�#�c�X�$�Sċ�bĶh�>u/�w2�^��dB8�qK��\}4Sx�IQ�F]���; ����tM�Ț�Ċ���}�G$�ѹ��JokV��:|E���$ҍ1u����z��ҡ���O����-1xuy\,l&a�9� #�r�����\�����[����l-���lӴ�x=��@����*�Q|�#�ө��*���WjGK�\��#r�	��w�"�sB1� 9��Y�7�扩���#C0��v8�b;�"hxyY�Zⴉ�O�����B�\�-�V�IY��~z�rڋ�N[d�K�%M�(�ݲ>�L��݆ ��} 07�������KSVj%��HT z�W`Cŋ����f�b�THWK�^H3�7�OW�X`q�J��'�*nX�1�t��cH
Y�h�n����tf��焳HXB_,���Ca�%�n�$��S��_���=�ʺ�FK&���e�)������>M��{ǵ�	k+[Oa���G}��ޖS�Ǆ\F�\�kj%��$j�f]�
�2��<iM�'�nw� ��3�����a���1��9+��~NS�����/Ķ`�S��;��S�s�C��B��-�~�f���lA�e<h�� �PI�?Z���K�3A��o��rxRT[�w��}@�-C�T����E�1%a�9P\$E\)]�s�]���`�BO�m#@��/'�2R�şR�k���S9^�	�>�а=6�uU���I�nC�Yc6פ����7.��I�|��e~[��Wd�Ss��aq���D���,e�d��gW��fǭ�(쏤�F���^�]H "Z���`�tw�!^N%����wi��ж�����ֲ�l�xZs#��78�@pmf~q:}x�V5�h�9;�xs�*�x<7�ki�9;�.�`F����X=�{�s$[>71H�΋E~Mb�%}�9��'����g�g������*xo�ݕ�&g/&���θ�%�ݾЀ#����|-��S�Vj��>�6u�ו5r�z@^�e¸�j���;ս�� ��$F�AH@�:�E�і�ߥ�a�����g�o�;uS9��Eo5��k������������o/0K|���D�����C��î���B;.Et�{��x3�y_l2;��-'�ښq�@�����_����TyDG�t��@�N1��v��|�J)F�$����E��w����iFUr`޷zQ{�˪`G���9��@�gk�{�gWܾ8�pu������.�B�W�(%W1�8?��<w�R��^r����Tݲ/G�W&ts�����~�*�\e
��$�}���?�x�߱^�+�0����'��ÆxL������� @D�F�2���a�4�r�@����\���q(���y�z�Fţ̨Ɨ� Dش�����>x��uFL�V�Y� �o�P����)�^����߂y^^�S	Gf#�,Cz��U]�������;!Jۺ%YlD�)0�8����z���W8�@��1��[�����C]��:_�l��|n���Yi~��>\��T���8�g�h����ާnN��F�@�fqS��;�zֺs
�y�:�� r�{��fU���������vm�vI�,��M�ђ�K(r��.㌑��A��kn�*��7�?�7�[�ܣ�<7G,��f�2n�����qJ���o%A�=���/̥&��؀$O���t�d�Yh�+.���|�w�X�_Z��%D�cO�l�&#t\ � |(��D����.*�d{KAKT�#��&v�%��iCK���e/~U���m L����	��ۿZȗl]��w�[,��L��A4Ȟ5��?ɢAEF?�8ԗ��������E���u��lTP(b
ID�
����'	#uo�YV�^���[�E��X�W��n�i���&�n�g{�}	b�v_��ot�P8�ɏ�s��1<E��Q�z�a>�7�
��fa����K��}�,��u�~U��g5��޿�skL��+e)A0�m5�t+���Эb��k����
iހ�6�tS�R���v�N�v1��6O*���AHi�~*r�M�z1�q��*�3w�������=�MbT1�Ȩ�q1oe������:��z�.�LӁAW	D��&�H�޹'_����{ZRd#��ό�&rW�{o�� 8�G��U��
�ٲ��iI��Q��b����V��Ə�ߤ��ׂ��&��F*kZh�
y��U-���e��օ)���(n����ܡ@�ȜS`����F�D�o+P�\�^s�����w�:<�<�X�ݙ>�����X�G9ו���_�"�!���
,HK�_F����\`�Yy�\��d����c)�6[�qʩĜ. f�UOغfn�?�k2��z������ѠJB�J�f���VJ��8}A�|S���Ȳ�i�->�ą�T�*���܅k;A����N�W;&"j	A����@����@»6�q�MJ�����`$��J2N1���﹓2b+V�D�A� ;gf��x4���6��Y/�L�Ӵ�=��y��c5�z�0�R�)x���ۙU�o�&)�<�z�g:9�(���V�wEd=�/>�dԯT^�J�rON�T��(�'Wi���A��fp��x�)�����/�����y�'�>��׸$�} �͓������0c/6�.Ӄf�*�a�Tx�|�	�Ⓑ~.W�p[1�6�S�E�����tp��9��Y}�jI�&���a���ܤ5�Eƕ+��bW���붡��<!���Me^�9,m]�����CAS<��E�U�b	k�m
��#���TyW���Y1^k)�_�*�i0�:J����SS�N���ƍ h1��X�~�gg�f�[1��M!ĵQ�"�5�|ള�v�,�e���P�G��� �U�*�cPZ��nef��*�O��{O	gcPӲ1oΧ{��#s����@r�냦�Dif\PB��t[��>�H�0Rz�=)'�W����$q�n7+�j�����@����#���˶>U bX�$�fN�.iC��{�t�� @�]$�z���WTbw�h�O�3;$+:r��<wU��^�{�"'�+fQ�n�����h5P�HRX�x^C��wz(O9Տi�?0�E(�h����� f�ë�d\/� �|3����`���Cޢ�i�MJ՘%�OZ��FO�)��B6�a���~4[�;#�*�z�{a�
�&���ؤ%M�OORqBTR�gI<�*�¡����O���h�j�]=�F�ͻ�9ކ!�\��~�I2ʒ��_wh0Ɍr7��A���2u>��g��"�p����0L�֢r��EG���v���?hԃ���ʲ�X�2u��.������V�d�W��	�D����nB��hG]]��G���������M:THM�/�o�J"���V�׺+Bš�'  ��e҂�6�,ɸ7�Ǚ�NfG����1vzJ������~G	H��j�D��l���S��	@�`�>y�K5<�U����`�E�)�)$�"ˡh�=8]��揁���:���&�\��3���W����0vc�����-sK�қe��Jmr���5���X�/�Z6� v�������3� V�_�ӏ��q�`u���pմ&ѱ`�}����4���P����ɳ��*u��n*˻��w+vζ2�Q�As�<�u	6��˘��6�4�qy�ƣ��ZJ6���_(o��ߩ9s���7A�x��R��hw5X[��ؙ�p8�ˇ(u���0���n��[V�&�wG�R�Lܞzmnf��L��	��#aY9��(�(��c���U���3��'%kv���ح���/Ř�2WS��d�ճ㼷��Y����� @�Qsg�L���],^�$���{|�XA�!��k�J���'�:�U��t̍D$ɳi[�n��q�{��%�9s�K�p��Vݕ+x�-�b���d
�ƀ�����/@���d��N��5Xs�i���W�1�	X�VXz���QO��$N���`��iG���$�a��=��c8�h�J���,�~~��S������1�h�\U�� �3���:��f_q=�>6�����Ƒqf��[h�E�F�X��n��dJ�C>p����ɻ�| �B���+�kj6xw�s(Z^��W��K?���Oc�%�텄����FE"G��ќw�q�!�[N��4yU��gt[�ҙ�H{	��*T�U��
o-�2곢��Y���c} 6��M��y���J��q��Z��x��b}�h�4�Q>�H����e�j!n3�P���=�γ¿�ȏE��3��+���iLH���f��n��[5Ɠ�-�A�ң��g�8��{�N}_&_�-6AP�=Sl�2W�ɪC�lZ�N[��|�\.�9����"_�Zq������z��Y��T��[��eV�R��C*�.��6$�qd(-���)�K�T��fq�
88�e뤯���y�P*��){<��$�!M~];7(�)����h�Y�M\�Z�@m����+�] e-�u�^�f[5�p���+r+��
����Ķ��g'�EX�1fvom�r%@�*ko�d��yO�7��aY�ja@��*�F�!M�ĺ�HXTҽ54�T�-����l⾮����$AK�pĶ�0|Z��J㣪N��V;�Wyb~s�\�m8� -�t]9���_L eEL���g���]�
z�A�_�L��	D�,�����p�n*��x�y��9.�ڂ��dϱ����nX!���O����- �h
��c���i@��O�n�9��'lG��	dq�O�>��d5��k׭�i�8m��F@�z[�̺AQ��mZt��O��
��3���|W��4��O���u$A�+c2q�XU�y�S	5��t%'�E��w3�I��>[?��a�)N���s a�֎���I2'6U��Pٛ�����f�O^�:���n2#�i�R`?̧�7��s!DL2+&-�^Q�0��2�{g�-cC׊4����
���cB�
��pO_�ų
�I�G�����\a}��sN��N�k4fJ�s1�s��R�R�/�2�^kq , 	g�i�k��MYT��w�}��%����v�E�q��`�sݕ�r�(c3	o��C��l�G�������O�^s�SdVEk���ϿZ6Cĳ����JT�Gۺ7~� y��6�*3�ߛ�hu�ݧdj�~a�Hj�np�� ;�����0�a-Z:�m�]8�-.�43{R����2J�$�u��;;T�����ǽ�����Y���oΝta>�s���f�K/� k]<>��ʠ�Y!e�a��B��.���Wq���T�����	%�(H*�ñ�*o�;N.����@K�ݨ���^»Ax^U���d����/�Us����駑�_�5�2�
�ϞvV~�c�h��YR�p]�An������Qc~Hr�D��Bg7�ͦLp��-�OV���۬�
��$�g%b�[�
�"W���J:�uah+wuY�(���� j����Ljh�nd�|�U�v��x;���8�P���=H�y��	ᩒ�N�.u@�ne�I�h.�N"�J1��\c�$y��
��Dۼ4;O+82_رR�8T:ٰ��� V���-%�"-{Φ��r���)�\�Ж)��_+�,����B�^�H��B��\��vj�Pyq�����|m���Wz�7�C�з�q�n���d$�L>~mb��b����4H��U�Q�҅����:��|���L��2Z���ج����D�ȿ����~��/��!Z�,�X�cz�b�����|/�v�#�xv���=�ѱ@�~�z:;s��a���r��G�m�Sg��������	-j'WJ�*K(��y���|�)D���1�پ��KY�s�����r��Ƞ��*�Oz�n�o�~���R�XM�A��X�8�����x��&���H�Чg`r�
������E���⮔őG�f����U�B��"R~XʲRD�0�8��7���롅�.�MԾkow=���������v	����
�Y�|��;�`jf�٢r.7:��.�v��DRu�)]�"� ˄�8JI�CLk���7`K�s��h24�'�)�~/<-s���� M�]@h���KztD� uʉ��,+M��=���܅����F�ۘb{%�'��	� ;�v��o6}��?�h?�e��E`��;W��pw�)W{-M�$���� Z�iq��uV˽����dnG���7Ly�i��
�Xa�eIBiZ�U��ʞ���دf.�ШNs[�#��0|�=�'(��눽�.|�	WJ�-b�̓�J����(���s�Ɔu ��|.�<�_.��N��i���������Z��Y��}`������*j`��\K��~b׈	���9�d�)BQ�t�����}�����@�Z���
/���$E���G�!����8�g�`��A�i��b���T�&cR�1+z2G��S��)��HU��~)���[9K8�f����;7 ��O������a�Xm��s��dI� u(�� ��v�&*J��#_�ST+׮��p+ӈ"ɢwŪ�m㶢��2O������u2;o@:9��i���M+;l�D�l6x�1.T�	O�[�G5Nd?ퟏx�\6ݼ���э�����|��t�g��v�2(a���y����)� �P���aM(�"���vv���rG��>[���p�U�o%O���t��"f���V�1����\����A$��k��p`��5��ZK�9ͧQ��+�k}�J ���8�E�v�cR |��?�#L'�¢��}W[�[^k?{�B�k��U]s>��n���y�2�X���1��I��0�T�)1T!ys2�B������ /����aصb��55����h�e>�|������x�ݺ��焪_<=b�7��Ia^eQ<I�l�Lm�E�I`��\���IKj}�k1 g�@%h��ҫ:.�l/�|�q�Y�l�V�ߏ�[^f�ӋE{E;������U불4�?~N�({�t�H�iD��U�!�ٽh�;�����Ɠs6�
�&0�@�(���WBkT��&6J�E�V�;7huwPk��<s�O.;'1���W��2�Pՙ9��ϋ�d-�b߼�c�*����_x�ٗ���%ޙe;�L�VL���$��Ljj�wA]\Ƨ����3~�D��"X"gy�&�.J�@`_�.��`��'�8	��(��;�V�Rk��@5�<4Xܚ�\�!VmO��V�g^�j\�	�/a	�ͬ����*ڨG3�[��GX�x�9+P�%�xP�Q�tl@���Ft����[)��b³���jN�bbʬ2CbAr{KG���
�7
��4?	��Լ�3,ݜ��C$��D��1/$�����S�> zӶ}_nz�uD���}PX�+�t�X)Ď���Ⱦ�D��NJ��Q!k�C���@!�#��ò�lI;u���;�,��%�x�UѶ��6b[h"X\G�ܻԒ�d�i^���V2O����ྨa".��ٟn��P=��e��Hr3d���M#8Ѝ("�<����vU�P֡�N���J k�����,�iIb�?V��i�I27x�	s���p��J`�C���<tBL�GL��5��Ώ��}
�<����ǁ}%m"B�� �<	���F2�?�iH��it��;�Ce�!)lb�Sw��=6�g�e�8�������FP�qwI�8���X��ڟ�}!�'�cdyG+ԙ7��I���Q_bJS;7vD^ԇ��[�y�~ऻ��wd4v�w%V��O]����Tt�5�#)����K"~J7#r)�q��UA��J�$�^o������r`E
pX�QӾ�}�Q��Q��]D�* �{>�y�vM�����3�(�U'�JΒ���'#8ɜz�C>�K��1��T�}���q뭈@\ch�@?���dPe��iٜ�Ǝ�y��v� =�g��&�VH0w�_��׌�(�Q��l~0�u�-�h"����b2[�7��AXB$Υ�ep�a(㐘g������R��]���.&k
:�y�A��N���}��޴��5�YA���f�b�ģɳe�YF����� $9���L���u�.p3�n���������%Y�pD�Ƈ3�Q4�5Y:F�J������-���Y��ܽO̽o�C��g'�(�"e1��uFY��$��Ƴ-�J���Wj�wd~]Vw!5F�c&4���W� k�	Cf�X,B���t	L�0Jŗ^��]v$
{D��gu���]��x4@�Y� V��LE	�Vȡ�ݏ��i�.�>��*�G::�]嚜'I�����HQ͞$ϒ�$8g :���/A4JYL�m�P����ҟ����~���!�1G�QʂbTNPM�@z�����*s��*t2����i�~���B�9�L%��i�Nc���]�KȬ���T\�ğq������ٵxF'6�<i�tB�ܥ�mm��W��<� �|�RO��>�f:'H�*�2L�����z=��pP�h18�]@,(�O7;���~��-��F��=GzY�\��lHU�F��&���ƞ���B��w!O�.�A�]�&,��� �ݾV	�-B�"&[�Y��,�F };�}@m�(=�M�^E�S\���@�4[�R#O��$�L-.�Β ��s���¦!�2C.����Y�E�A���ɓ���×��?�T�ȃ�� ����h�b���v���'!�`H�n�)�YOr������X	Ͷ� 2&¢aq����o�Z�f.d���,��:�rD�t����$�h�m+ML�}:F�%�9������=<�TnY���u��$S!��>֣3&�67�L�TU���A�;�����^n�Bo����>��ctk�����$������v����FB�s�e��Z����9HΥ&Ay)@�w՘��yhU!5�4��m�8�^�vf�375����D`0��-�������bh��y�?!�N��/S��V=?J�_ڏ�_^����*���!5�׬�&I��Q�Z���宮�q���k'Dd��t�&�n�����ru|K~R��b7UK;a=2�If1����yc8�7�+��z����Yb��� 1v.Y�@��i+��GGܝ ��I�f�/��0���hlE���y!]�ȋf��|@�Osw���,{{7a���>��8��6N��D`����r���\�i! �RD��b�v��e�\JԆ����t<��Kщ;�挿�t�{՜�t�NEc�DrU��w�i!�6Vt��aTM�Wt1nK�0�����ރ��%��'�Ed��T��ad�Ez�����7xX8R9L��cn|O���F"����uJQ�^�3�A�H�%�<�{�W�{.�e���iF~��ߨ�1��rG3�Z�r;P^�*��������j&����|�ˉܱ��c`a��D�#�ܧY&�
�a�ަ-�j�׽��z5b����Vf��x�f3[!�bW)%l�Y9N��LJ�5�V��s�=g����7,�r'�*��u�Ѐ;�X��7@���o�nI,�i��uЉN@���1KМςG�c��.'bԐ)��F�~z*\0<���B��&՝]�Ep���}_C>��!K��;�h�������t������id�H��uGC�����|�kO?$v%�⠵�ߘ I~��5s�o�����+ݒ�^�8��悒L��ײz�6��(Z·�X�>�8�[Ɓ�U~I >�Hca?ڲض�u6��Vt��~B��v?¨v�BF��;�e���- ^�&M�4#㟥���[�8�y��,��݇n�Q����ۃx���r�t��|�����$WW_�H{�w���RJ7�QWY��o�m��˿��]S"H���eΏ�x�r��6�ظ�X잞��"�S�q�Oǿ��{l6�������B�\���Š�����U��8>YV�_�>,��Ɲ�L����Ŋ58�΅�3=�����(��U�e�� S5w�ڔl����'S5��"����I�I�hH�t�;\Q��	���.H����$�bN9���]��LUP-�| ��ы�CR"	 �o���G��Z_���.������\��-A����ZMN�t���1*5B���g)i��S/S�*��5�l!;�(��k�]�Q]*2��3��J�h�E!u>��L(��Ɛ�em
-�O�q
�O6���$��"�Q��&W;x|��Ѐ��Bڟp&-�E)�����d�W枯�����O�<�����5��N��u�+D��(*�_�6�a��w�J��',Ґ`�`�0�Pa#�Y]��(�/���r�U�?�=rJ�Y	ea4��'v3��D��? � @��A��O�$X�-{Qc����!?91վ��v%��p���_ɧ.d�-����;`�3�z5��9w_~
����Ǧ|��Wf��y���y �]͠D2:R�&0�����6�W.��9���9�&�q] �,���?�N&R�a���@	��t���ZFϩe���*���"m�(�L�|./���h�N{00�|��t]�s$�J��F�#�,�}��;>��0�>P�7qU��w��υ=.f�x���h�R�K�j��4�[иk�Bc�5d~�-!���A�{g/,��ѝ�Q$��Q]�݄hU�!Y��f��~�[��"�wBdG��.ʸ�yn��-[�E{ x��b�ٶ*���;C=8�M�#�$�1��%��ڸn�©A	�z��w��Gh���RhD%s
�!�5�w�i" �^s.ޠ>��9,��������UJ�KO};5�X�f�<,qSn0%�|Ap�k	��������\x�'�����n*O{ؤo�mȒZ;�DH������hF�U��m��HDg��s`��l��J!W�K�`o��R9��[�T�!�ٗ4�ћU->�!�7�3(�2�wť<*�=��6H����z
���N�M�4��ё@O f�35/t�S�/"�c'՝T�b�������. ?6~O�ʢj������Pl3�K���M�;���/>$;��@�K�R�K�ʻf��rEc�K��Ak������ĝ�+��J��^�k�o^?W�p��Q_8_y�������C��F��L�$6����p��(@]��	 w$O�<��;��L���Bg�HD���Oɐ����T͎��'���j�9�}&ǱV?iN�V�m�):��x}�1A�%>�,�wE������ Q��{S�h�x�N�D��Wq�tVXl��V���/,��;�$*��ʈ �#̞��@���'���8:"Q��6�@��`>�����%�`O6�K�p�;;�*<K�a%�w���#��>��H���b�Ҟ�*{��R ѭ[㰒�舏���j�n=�7�
�s5���s�E1�4������Qe��6=s�㳫���B��l��DZ��o�TH�[��2��Q
��p,P�'�	t�����K�A	I����E���;%x���Ճ����1}5�+b�B�4~���:�z�y�3�I��j	�@'5��J�g�Ez^T��<,�Y��ۭ���_?.���٪Ώ+�c�#���; ����*�t�C�W�{8�i�l�?L���>6V��1u��1�pu�"SCi��늍֣jX��ƓW� "td�#]Ω;��)��ԛ|s���|h�խ.#W������5C�VFH�+�ạ7�ƐU�&tP�I�Er7���͔���(Pg�y��J]��V�{(�\�P���;����Z�ʴ�ǹGF[��8���6*��a�E��#"��u(Wo y.&[ɥ�.�D��Rԙ�R��.��Q}xX\r���#�a�'�-���顼@�{��vҷ>󢢤���'��Pej=P�M�c�(���N:%�g��u"���:mI�+�y�9����" �Yi�zm���k -�,<��L�u���Ks�:gdג甗Ѱ%��Y��Tߛ�t�V��7/�_�$�}�����g|�E�X+a#'í.J��K����L�,�g��5Q�(��x��N��X'�}Yp^�ώ��79�&K�B}.���c��)P�XyDIOP�Emp;V �hI�𠥧j����Lc���]�rr�6�!irs �ޔ��:���Y�9�s S��k��Hc��n��#;�Ę�'2���H3׀Pz��]�s(A}��XL�Y~�K�/����⭭��N���Ȏ�c�d 
'M���[f�{��s�>$��/#��Ņʊ?;�+���Д����>6�ܩP��-ӕ���݃��a�z�Ġ���#�A��Pj��/5dn�Bɷ��U&i�͌p��dU�[՘d�	�J{��Ov	͉��vs�'ǒ��Sa��$j��f�=�KP¸N徐���׮Nq�E9�ͦJ�7e��G�.��xA÷ց<3��u�q���#�_|}����`�F����iq�F��������W�ʢeI�z���mS�U�)}sҌ�՘)ųBt���H2�a�)�x?��M�m�_��5�HZ g�>���5&��g;n�t��;�:�c�;aA�AĞ�%��|���M��2�;Z��2ꇔ�5��{�����Ī4p.Tj?ڂυc���ΰT�p"|}5\�U���9�����<���Rn2��ڵ�A�|AR�VM&%���Ӣ����Jn�r�~^U z�0c��жh+#��-��T�T@<�˸�U����u>~��<��ǩ���8�Qv��S|���d�}R�2���9��C�&�^ms�?�ӆ�dWP�Lu��4��O��ό�¤�`c������S�����΁�����:�w�j"�U�ِ��"�$ɯJ25��p2������p��]���J����&H�$My��JO�������j'����UaH�,6)�z��<�{<����,K�ŀ�h(ߞ�0�Z5�v3o�\�t�|�H��D����em��[(�Nl5!�M�'X,�X	>�XJ3����#�q��r<pC]��=�L�����M������q�'��Z�S��#-���@����$ǹ���YE����w\�i�`�l�S��[r�;?��ɯ� ���P�Ӡ��3�r�����s E;���	�BK��LҦ�CEőO4I��P@��NM�f׹�M{�=���Z�cŝ�P7­k%��H�F� L,_jg���yVO�cN�V��G��H��7�n�4	觳�d��.g������V��E|0�~� \*��1��Ph�3�����9��<"�A1�?Q�۰�%�t�+x�1A7�C��5]0K]� ws�G����^w�p`UWw������SՔ��zT����?Y;?�����*�b֛EbM�a�qZ����6t�u��>�׼���0 ,T������{8�����{+td�����O�D��z�H�3ҷ	�P�f?�V? �l�g
�B ��PE��7�l�� ��[r���<��V��tHK�B�֧�
g&����K#g)C8[P0)��m����ۆ�J����}�Ԥ%+����p-��{�'6��1s�t��셄�׸����'J᳚�#��/����G\�����NKр�?�l6���w$�%��Ie�.�,�|?��>�A)nL���E�H-~c%1cG4>}�>uz�):�`��=,��x��B�m�9�@��'��l��=T:�z9���V��e;�^���Z$m�IP��hж�7��<ޚk�֨v'#�щ�ה��Fx�B���;p���cO+���Q�pr�"Դ� �b�6�	{�i�����f��=��d�ĩ��V'O�S
�L��J'�:�Љ���.���z0�h���zE��V�Oj�b�f���v.�K������TX��}��S���K1�˵6�v
w���]�0.�*��!Z!���N�������ypx��`y�_�NL�gԸ������ϕ+/Zd��L%��x�\
�����j�U}�ڐ����x��ҝ���u��#�������/Zf��49O�X�	��Xt�N�fj|P"��mci���@���7��P��3).��Z�`��k�P��¾��PXI.�ʘ��ځd������>�֥gh��I�gz�&,�?3H~9�G��|Ma	i��QR2^��G/��429�*�8�j0��ۼ�����+����a���!'��JN)Ɣ�ߊ�f���>ʲ�o������_V�G���B�"3@7�Ĭ�h�!�6��(�-���B���ط��5���R(t�4��6/mv�e����vV�
au�"~�E�. ��0g����n+��7�/�%�T����d�5PD�
/�zb#��v�"'ϯ�P<���fX"ȭ$�]�q%����T �R�*�.��^������X�����.���$�
ڐT�r�إ�6`:��G(���qA�?8Z��͵����
�{F�\���b{����	�:�h�IN�2���O�b�Jg	�M�%1<vء(/�Z���	��ܢ�����北��7].�j�A��n��|�T&LjY3��<ˊ|$�?ꤘ�\0z*�B�m-h`�m��M$ZH!uW���������C8�>u��fś�y*�5���{2��!AEp����袕YhoT9o%��2�|� c�Oh��?�ZA�8n�R%��U]/�����X;��z	#{� �a��!�i8��_�b��pP!.���V3��9;�/Eug.��V�4���&&�wq@-#��Ï��&���K��)���l\%5M�ܼ\��m�� �Z$Xd3����2_�p6 �˗FL���/�& ؟w��u�^�j�9��ՌA��D�k��@O����mxcrzXՎ4��-��eߡf<�4L6G�f[�̦��N�;����B֬
�ޜVF�R��D����y�}� ��{���}u�QG\��$��������l�K�����s��2�9r�{DZ�M��������nb|u�*�7,��k(�>�c-�8)���V�p;�:m�93�S�Y��O�g�ƾ���QѺ����G���tm�,�q���6/�=E�܆YAC�(��u�����V���J}�h+!{��IH|��i[aX�86с��yq�A����p����L�)�dJm�E/�n�����j3"�{.M'߸+���2%D�L`�f"��⬄P��EP0h���&�ei�`�:��l�7� �Ɣ-[9P)�5�tOX�����!��n���y�����`.^U��>[��2���%�`�5&�nﺦI=lF/#��M\��ƃ|xm�!}˝�a��$�i1�5;�{���+ �����R���km�,�\��b��m���F�r]ֈ�b/��q�(� <�s��k�H�#�X����2���f�E#�*,�84��s�Ru�M�UŋͬL���;X�nם��W�$T�m_%Vl�;�5��t�˝��؉�6�W_O�{�ʫ��e��#�|J@�3�� N�Z���ѵ�N5e�!��R�s�p�@��&�hk����qz�/l�`ء�dbeƗ�t��QWCk���Kn�I�.=G�1�ۭ��w�JsDD$X5���\v�j.ZIIY'����/<8�ѣ��Ӻ���֒O�cW�#�$�A�h������	�*�T��芵I�|o�� �"VB��6�Q(�PW���6����}B���{<���92�}��`�Te4�V��7H�&���8���z ha$0+!8����I[��G,����Pfwو�:�V�}d�17�p����m����+b���݌��dxA��W�7�*S?�:R��RR	�B�5��D�������Ha�H��;�Ԩ�9��h�d��s*��a��t	���ή����T�z��Ѻ���@= �6�n�����޻u$��:� �t1��=���E�YM�z:w�z�*���"�5��پ��H��ھ�%eF~
h�/������b|{��ܵI���'}ە��sdr������;ͦ�$%	5�.?�H!�ǿ�5l�����������OLB#��!X��Ht@R��QO.X`���z��&_d,"��y��_�`�u��+����{+����Q���=����<_�
?����LXggj���L���p�te� ����Ǳ87VD)���µ�~@/4�אD%�=��\�xa�8�v�6$9D'"Vr��a2t��ˢ�����Z=v8���o�q!�l%����}9�o�4���H5j�~�_&F��*�S��xKo��.���5کӷ����
�o��e!�
@�he:��Ѳں*p��vӽH-K�����V����p|��9ֽ�)LGuthID� %�(�F(�9��4�מ�O��ɰqQ�ˬ�[ƊEg�b8e
�܁���&a�a8ʾ#S�*�2�e��E^�^Vp�SXK LӬ��^�5���qe�E�2\��(�8��Q��3d$P� ���c���/�
L�O��ٮ� �I����o���f�
i?s���\�B�l�q���7�X.&�5*7��(O��Y#;��?�-s�1&:�w�_��^�QQ#A�Ff�/������� Z�[3{��1�k��0��b���h�P[���^�܁�8���66��P��j�������J� �2����e� T���+Ќ�0F�3�VϦ���$��J��oJ1 +������P���Ò�lT��R˻�ϵa�T��&�M���a���j�Fl~��#"���̣����IJI!�"�8v�w#{MX!�_M�
H��Ѫck�Aϟ-�1�3�,+A��	����O�%y�����H���2w<Ε�a���<�n�9����ܮP��w�A��'n����(���Z����<W���"�)<�� l�U-�ǣ����༼D��	�Ro��~H	����m����I��_���'
�W�/6)��.�f�}Y�|��|a�.4N�n{c�T_��K��%?���mz�����o�
Ĵ��IW��l�
���f�[v��"q���dj�n�7~Kz��o�r�Ŋ�[k�F���N�\�:�%����<<���퐆x�5�U�
�Y�хe}Z�q�n�� N,;�"��.�S\���:��?J���b���G&0+���k�;'d���kS	�/��\F�a��]��O�d}���#{���S�:(��$pƪ�y���:��y9�tG���	/�$�B_�+�	֧�7��=��v�Tr�:� ��Ad�̽L��Z�u�}��g@�72�n�4;����I(~�Ǭ����9����/�7&�ե|ǬHE/3fc�-�$M�c��h�M1M�"|?�u<8�8���HO4�,Ԟ6EK *�T|4���12n����"��H�w�q���a�x���/��YJ�r�*Ix&�aY�U�S<�[�h��@��2'�c9�P'^�[Xj�YI��s����#��2���*�V�%tS>%0�']������8q/�/(��׍�ߊlK��{��O� Q`�����x*#��*��t{qkz�-�J�c�Y!��rMH���t�S�P�2��J]�f�0a׈�-��?~�"L�-�G ��f/kV�A�.D�gX&�-���+��e㰾���̞"#7
"q �n�5}�K�ׯԁ���U�H"権�K3ɬ����2���[�!�懁�VEd̈́�+���Lt�_�C�Γx����r};��C/��H����L��1�-1�)���XS����/��I�R�\�f���jI,�y��y�U+V��we�/WQ�=�&��u>���W�*��>������&9m�1^�{�_L���n�M�����R�K�M.~}%��s�;ఙ�*�� �u��F ^�Mc��7Q�ǁi������
����j��d�<�LZEEP2��~V%@D7]g��`��ƍ�������	�;J���U₲��(S�*]�3ɽ��K>�s+8B��m��wk�TZ��ka]��1С�Zt/���Z�m<��3��_>�
IH����+jS)�������r��7RBPE���*��4��B}.�|�b[�ry
)��{pt��*W���7�X��	�����/���/2+�A��K��+�Hr-;M��� 	ב˛;��$H���YX�E������Ny�e��fXG
�%N4�;	�iT*Q�����p�$���Ȥ��z����]Q�O4������o�P8v̥�������^��|"��.�q��CUm?�K�7~�P}�ʃ��x$��3���d����O��<�K��3��X�[j�	��S)��)��]bR �:�1���k�H���u/��+ʘ���L��,��.IU�U�=0 k��
7�O�Bү(<Y	�`ʲ�`��|Ur�z �J12�,\�!~����Y\����9^�T�ݕ2Ƌ����3U�Q�����&�2~�>BK��>	D2���Al�ժ<�.J�5FSIq]R�ͥIP������3h���WTW�V���m�2'���;L�L�U�QI������$�/�F�A�k!g^�����,�A��O<��0�1L`���ʀ��9�����w�}���߇�i�v٣��J}�fh�
fM��I�aJ�<)˷��u�� "O7,l�����|�qGy�7V�2<9<��8�{0���-�#1SP�1n<7�>x��V�� �b�Hخ�2��� t���#��;�/���|Q������
���|Y�.cc~�K�=��q�/����z��3��]M�*N��|���GdD�ga��;�<�j���%���|0��#�r*A��;}��3o�'9rNU��c�A��`���<5Z�-� �{r/�`�#��)��<P��Y���~hҺ����ᑙ��I����É#�dJ�����.ɥ��^��4�9c�^G���|��qNWy���b*����p����֕��+(D.ڍ:$����a�XMF�C�M�WS�o,��ۿMs�J��^���e��/+`�\i���_�\��Q�a�����Mf_���F��rk�m�����b|T��6�'x��D�q�TNY*�d؆��-��}���� i�mj(H�}
�QU��o�	�J��A��ed�g�e�X�fc��ON�!9XG�r���]���_P]�����Q1,���yW5��0X�L��k�U�p����Q!,&$1�2�����T�E��,7#���梉U҈l�UJ���n��<��~u[�su�Fw4X�ﲐR���D��k�F0p7�H	I��G6����E�������Zw����s&��Ql�u]c�:�33e#C����zB)�S�����끡�k���k[�IC.�i�F�l�(b�no���4�W��=᭣'R���;̼+���Q��-�݇@�����Ƹ�a�vf�����ڀ&�e�_T�<L�d��T�,�q\T������M7�_W��HQ��j��N�:%]�������H$���z�7`��If.	Pk6b���e�'�j��mE��Y�=�2�NV$�v�ýt��\�d�
)0�A�$���؉�R2�O�lx*�~�RM��aZ��B��^
n���Y����%D|�Ѭ&��#�؁ x��	�RGJ	�S�Ii����<V�� �ʖsaz2�M�w
�+����*�}%gF�m��@�i�L�x�U��ǒ�!��	٬�h�S{�V��zƊ���r&��!*`9GL��~�`{�5E�X�8y��7�x�`o����[��^�z-�;!�ԗ����Dl=�m
J��!�����3�1�ٳZʇij��z\��l\��~>�t�TSrc=HK�N3�[�O���@��A70��!>1ڕX����E��a��>,����'�!��M�ix�P���1���W �щbO:���� �� Op�..pN��-_��Ч����]}#�$/L�d�>��Om�U4#,b{��5є�є�sc]"�����9��`^��7;y��Ɵ/{
�Gq��
z�P�w�I�G��p�k���$`L�^�Cޤ=�u�Q6(7��+@T�Dr�I�	��g0�0�����,����rN�9�́�g�k��(��up��d����K���WX��,��-F�U%�Y��/�`=���t�EPԕ}1`�/�ӹ�μ���A�g�]O��́~)��.�hi1˩G����(),cz7rI�)0����V��W4��Szoz�+��U����vp���3D;�C>�}O:&r��'�t	�)����\f\�*Co��Ҝ�|�?s`�h��,�ҨG9�n#Oy.��\ծ�Zu��B�����Q���{a8�!��<VyYaw��
�64e��j�u�JЗw�0nݥ)(u*���I?#/N���@��y�C���d�/�CԺ�����넅3�IX�Y_8�.��I�HР�5:���I@[ڟ��.Q+����*e��C
�tM~^	����~tV�����>0@��p��/V�.�����/) (���Q	�m`D[��2+o�>��p�]S�V�;�'8 >��m���ݮ���g�TJ��I���f@9���9�#%�ŵ��96�ֻ�S���H���Ў�tO�*F�y�*�������B˧��e�zS���ׁ�c�<�w�36Q����ʅ}�y���c���?V��;x$=M�'�Z9b��K� N���1�Iە9��O�I�Q�q��$mgፆ�0V,�1�wE�j�9k�%l����,���t:��=�'����s��cFY��nDH�y"��Ú�? �V�c��O����!d�[^��u �6-�����,�)S���v��{���h�y���Bw��:�׃{�\��XYAL:�$��~��p�^�؛�ra惓���0U��_�|�\��t�z8���hq���W n�[�<{g̳'
l�f��,���T�������[[�ŻT���ҞF.c��������(/�I���%~���J�r���#�[��]k��ݠ|=�t�r6\��8�8}�@�ynM���l�k=g��3��p}�vL�,��,���zίfĠ�Ā�b���x����"~�� (g�+dOXH�w9���I �]��9��*ɿĀ`��C�DGӯ$J
}�l*�v٠�V��v��$+2��
�<���̼���~����*�!
������/����c��!}����#���Vp&V3l�,�Ք����ԫ;K��$X�l�u�lT�`AԴ7���yL�|����\�)Y�ϳB��OS�T���@��nZR��g�0U
��w��}^���L��D�siESc�&ߎ�׹f��1r`B.�dJ{��Q*���
}��ZҹHxb�J�L��6�	>�?OG�ؽ��'�D�q>�)W��8ܼ�l���x���^���uU�=�t4�Ce34+CW1)ȅ�<�����_q�?��k�,�t=��!��x(YE�/߼:1_:����e�8��
�?J��jE	%���I��a�RW�έ�?��w�+�CU�I2K�o!�T����!܌�P�\��]h �����RwC�aY|ߊ� ���Q������ �3FQ܆�S��9��H�:� �YE��M��4�Q�!Qg.ߺlF_��k/!��ۑ�,���ypv�IL��،���Hm��NP��Ӑ����9�yV�]_o�ٸ�|��M�A�uTq�M��U�VG�-���c�?��_����*�l4��-�u|ma�g��������
y���b��"�9�X���%*;wδ�ڹ��'|IA����45b��m;�*\�6:6�z�`�]߉w vr+���Q�%𔶢�&A� �`��P�M�wm8[��źZ�����Zo����R:�H�ZL2c�[q�Ze@\�:?�='����ࡢ)vIi�@w'�$�@��%��� �0Z���!�0�!��-ޖb&"S���v�*�
z�ܥ�xo�� ^z3;��z����TEΖ�G�T#��;7E�@6^>�̌�v�7;ͽ��<_"w`��/;,1H7��d�2�(�/�* n�<�\/�G�F���bb�B��꾬�80���U�KR�D~�n�;؅Y���QJ�$蔏�e�	�Я]:��_��HzO����e��a��oj����㡃�{ڴw�穆�k���S�Aĺ#����C��Q'7�����b�g��{�s����;�(b�:����L�\�T��H�#�P�΄-�D�
�;�
�}X̬�����z�� g۪��0��`rh���!�N��!�3�����D����O@<�ziK�m�j��O@{lk�8zY�>ۼ�4�w�wW`��h"�)5�.:�/:��K���L�������t�B�sIo�S/�]6M)W�-0ٖ1��?��G�tW"�!�|�R�ǘ��N�="
�:�����k%LB���@.ˌ^_��Y�<# ̦`�Y/JHhV��I��	ڪ��Y���5�,9���C�Kgh�h�9����t�q�cQ���+?��1�5�chu�%�������^H�kI�A�`�Z���r�Dg�x�
fZ��(-�Ȉ�2|z�	#�B{��
���uA��4 �)���W!���E5���@Vܩ���v�M���t�АU��ؘ��=:���}bɮ��.�5T;�qc��dщ/pۄ�����M�U�ix�@-�Bl��eO�-��<�!��@��-��E��v\���Q��ö�E�k��:�B�9��$��Z�1ԭ`B~�2Yt�J;nː�JC�K�m"M��J]z����}�q��#ۥY/m°�����ᾨvu����/D���2P�*_{�6ħ_�Ky�N������S,3F���3����x3�����m{���f�]����I]�]�e%Cbc���]��)\���/�eo~���*��R2���nھ}����>ŀs���yާ�׹���4bV�4>5�7K?���v|d��Џŵ◱&ˀ�[��%�= q��!P����a:z��E���j	E�?�{)U In��^��g_� {d]29�\}��xA�=,����ձ�j��
�	��*Vr�'�Y���襤��ф��?��&N꿅Pɛ S5�,���h�	Ml� �,-H��DH�\���H)�~=��l��.�X���iS�B��p���JbK�6��%_�S;[h%����V,���H!>�#���� "�g{�3t4�=������}�n�ٿ&,q��Ԁ"{�aO�{���~����9i�}���*E���Y| n�6��̞S95��p����M�f�'�-��s���2�%Z��z�nC�T:��q:g��Ȏ��$.!��\�ۆA]1�	z��m����A���mQvUB9�{*�S��nKI�q¥k��n��ʨ�Z�A�ϖ�/{҉��J�>�'�z��	}�2��T�&n��������y؅B�R�&��ab ��`����Tό�˹d�Ʈ�"q��%v����.ϟ���|�
�^�#ޕ���X̼G��p�z
mWc����
��.�e�yU@j$�"�H��;Ǜ�^��p���TC��_meA��W�#S<iXl6m�����}�h�Hn���}�OJ�"jp�&}�H�,�ְϿٹ�!�$cqh�YQd %�2���=�ӉP}>(Z�.ަ�i
���`���Y�̔��� �{�D��5!n��z���cM¨�L��,6s�V�w�b#��V �0}��^���Q���Jb�L�m˕y���~l�X�x�&
�,!gI_�u��FU�p�nZe������&���|��֣L�}Q��[�V��)�d��8HA��D��su�Ɩ^z������p&��2u8!5cO���BUZ�#�]2$�����s,�\۟�ȷƭ���!�	��݅�N�ؙn��;�^߂H�Yq�c�D*t���`�:��7��*�A��_�m`"N.[���@�6�L@ܷ����]���2<q�w�ϨٛЮ�)8�q��8�<ҏDuF���dyu�d��q�!gPw���?^^����h_(v��R������yd���F��O�5�����i�v֊X��[���,�Q��k�*���m�xܡ���Lﴘc�0[ �Ԉ]��G�"R"���l��1a��&;/�<~z57��N�zH����Z|4��������1����V��0��9��>4�¶�/�K�R�?�Ԥ\�G�.�c��#��G-�x��[��8o��Oh�f8��3V���eJ�=�Kȏxj���A�S�
�XN��;�v�_r�`�A�Z�D�_Ր)O�X	�M�~Q0��t�t�Kbd�jC�m��w���G|"&�́��Ȑ^X�)>/N�ǈ�"�6S���N��j?&�m.��cOĿ�gE,<[@�C�u&y�4�\V���n���/<�LGpb'H̚wpo�eـ �D�g0E��6�I-�f94Z*#6���T=�Xd�}Bj�gvU�@
c��.[ɰXBE0�G��s�{��(ih�Z�/8o�}���m��K���M�Cqlj7KT���������l����qf�<��_����#;W���v���t�Eo��$xN��:[H0��j|�e&�H�r��L�T*�i���P���/�����	Z��YV��N	����c�GyA�D����ào��M��S�Qz��0UC�F-��+��.rz��?�&}�&��w	^�p\�Nm��c��(���f��7���u��h1�M�sF�����Qbv9��r�?t�i܆$Jt���ﶿ���/3��uM�j k��yV֖c�~�N���T���V�^wɑ���>=r%�+D����ў6��
����·�E��GjE1'y���[�$�b�!��e��c� ب�B��f��L�+���L�N��4��i�%e�K{�Nu(\n������	3>��Q\�K������-�6�K��ڤ�6��r>_N����j�]�X]_���.|�Do\(l�]��1���V�a�H�XW�#��?
��H�ϚT!�DZRHㄉS�� ߅ݘ��8�]*��W��O���J?3Z���	a�\X����ź	��g��(ٻ^�^5�̽c<v���`c^����I;�����w<T���o��׊l<[2�fւ���N�(r �G���s��V���}
`�ޝO%L������2����Ghm4�	o��bA���3�i�R�/V_౵4�� sr�sT�������BOu��4��Z��]j���^XN�^�m��/o�A��» �����R՟v��\ڷP�W�_��PC`���s�O;�n�9C/�/W�i��(����$D��A���?F$��4 �m����&<=(w�e�w��w�� ���0^��q^W�(|=�ݛ�F�d�CI~Z��PĊ)c{�Ѣ�{���F)�uN/���*�́sP���a�>;'T׏��{�n�y$)�������r.��7�g�-$X�"�~O,gRg,��2�?T�QsF�Ê��i8S)��ء�ۂ3jA�3��*�r��r��E�c��1)�T�-w�f�����݌�b�0z>��=)�WS��;_�}H�/�2X����S���B}��@�ܦz�=�~z�"G�e*�N���*���OK3 ](�zm�Q�^��c.��f58�N��&{y���J�z�4�� ��\1�ׂ�$��qW�vL�oU]nt�|�C��N� R��hS�M�ȩ8}Q��U�-/�V��;�m�D�K�;�E�CSB�[Ɇ~N/&����?�*�I�E�Aj�{�U�;1x�8\����kLR�nx���ǃ���x*|��n?w�WALb������r�<�1p.�����mґӮ�&�)�!uZ�3$�d�@Ϲ�'�����E|^*"�61�1��P�/�a�)��BJA�~�㰸5�
�aែ�fɵ����pu�sB�Nܱ�5�c}����D����2��2��*�V�)��~�>Ep�u4����HY�X�@b�ݮ�,�ËR������8��֗\�Ŵ�T��0�
S��]�Տ���ޙŘ��>T�����GV�(�H7P��Z�c�/V���5��t��X{vaIt5�h�6��'νB9�{�mf��$�1af���~x�_ˆ���nC���߆[/xAw����r�.V7#�t�r+�����.�u��h��VMe��ZI���\�s>L��v5g۫i��9�!7�;��/CqllU���Y��]G_�;�f��'�*!B�F3����b�Ц9���yb迄,v�N�3��)�4�%b��JH����;v{���^�-	G�c8��ʇ���M̢�9�zsWT�p�L�=س�۟������P}�Y����� Æ����p@�e4��=w�m�&�_h�O*�m���%{l��O�s����05�#�&� �V;"̏Jk�]��f�)��,���t�Y$����$k  6FP${ �ҧ��
G���r#��uN�Zbj�E��!���G!Z���p|q�PZ	%����B���ھ�~��$�+�%�'�������w��#�.�:�6�Y���ཛྷ����>h{�Y�K�� j��+"���S$i��p%%�:~+4��ɞL�g���>aj�M�q3�q@6���`�%|�Y�څ�R��0q�d^�$�*̖����^hj�Ѕr�� u�/��7@��I�mw�~q�/���5Zc�+01 s�gI��� �� [ -��a��y���;��L����3�y�֊�QG�c�.���-������|��<a�Y�c����>S)�ţL<�%Ϥq�^ے$VFj[ɸO����`<�1N�{���>1���5x�5�Q�����N�;�)@gU�L��CO���*���L	��$)Q�r,ɨ,��;�k_�*S�٣�<�4����/]ErE%DA�ǚ����b)VY�E2��l��?�Y�_]�ĵC�hn�"��wP��9�@0���/��C&��
5�+�2怛��?k�#o�*�}�w����4���k������Da��¦D&aKw�a2��s���:��U�������+͕b�F,>w�+��Js�-v�n<�Zͭ��H܌���k$��KKo��Y��lxiH��d���������'���tkUVX�t���ɨ���eҠ�Yi1@�ۨ�������d���ci[a���c���Z�t��x�<1���Ckl���Xm8W&�($�z�o��!�$)�L�y�/���AN����i>$S4�rU���<U���؏�6��0�ݷ0�='��#�$_�V���ѡ�t�c�հc8���p�AW�u�,*Q ��yLN�f�D�λ��<����E�|%��gEz�0�썊�X[��W3���TbXd���ZJ���ޕG� �*���m����N�#�,����N�9�!>A�c^Dm��t���O�Q�?J�T���ݣ���7)��D)o��1@�9�_xO�^�Mp���n5e�W2�tYӁ
7u��y��qD��b�����3(� \�K�U�ot!7����u���Ɗ�Zɔ(8��������C�%AK. �p�6ǿ�������9@��2�|x�)�w(�XAAO� I�qN�F�+�k��7���P�x]�0 � ;��6jf�c�ڿ(+|xk�P�	zK
M{|�m�}ML��ȧY4zÉZ�T3�U���(���SW\����>�,¡���� d�-������/���0d�~��Duq�m�^��Db2�����W"N-�y�f���k���D��å2>>h��Cʇ�ܶ��xv�4	t��r�k�?%v�~�����Eºj�e�1~D��/>M<ҿ;���5������5§�M�ok�O�F�]��h�ٺ��(�,-�_�@�,�G]�e!�B�'ꥌ�<G5B&�w3��-4�z�����3�,ll��?�-�ZHk��w㘉m�P9<]"����X�����ñJ�}~"���.U�*0�n�#^��H�r�Ǎ�y�CsՀ3��h�^��l������n 
�oh��\a��{�h�}�����(�� /3,p��˿�z�3�Yw����^����I3Ha��k��0B=���5*ͭWT(7>w�3���&�/��-|�0S�����3�>I��L4h[[J� �[#�g���Vb�E�h9��5��~��ƍ�gϿ�_��o5�+�	ڧZ�'qkv�Ve,�xd����I"�+���1ҭ��u�D��s���9(�[�n�Bmg�Ί[�X�Sݢ�y���S��	��{��S|maN�
5	�fa��O���>�{ݒb��0�����53*��Va˪d��xN ��6A7n��k��_���Y�P�����z�-m� Cy���mZy0'��-�ͷ;��QK�?qoL�(�p�s���Bg��&mˠR��v�>�ޓt���w
�as�U�������A������OY�S�$l5 �_u�r� M�Qh���9v���_��^R�4�&�l�ɨ��ì�y�H����)"���G+O���a���nn�.�Aw�?�HQc����%��5_�;�O�]<�nAD4-��={R��nT�IannN\����7�\�����aY%sҕ��.vX���`��T��N�£>ebR�4n�8'�m�)��r�ZFҝ���rP(��iP���)ȏ�%�5��zR�[]a*z�`�>S%�-d�gˢ���d&$��⃢�,U�U�{)V�hy:�R�S3)MS�q�:�&�{gkq\�Z��Z��np��][$���ݟ?٪v��χ=�
���2p��p-$���I)��ale�b_X�B �-kU�:TJm����O:�@v����w���KoO�w��ݖT�2cenQ�e��if�;H���!�o���𢌭�C3�i���O�@��2"�"�9�����i����)���p{�]]�Zq��Ɓ0��������N����8V@�ǉj٘�2U��ԱUi��h�9����9��Ι��H���a��f��H{���mA��ʕ�\R8����ԝ@����Q �T;�d(Y�X�M��:�[?m������i��p}a��+�Yf���>�&Z4R
���!�_@��uߢg��tA�=LQ^��uSX#y~|Y�qȜ2��#B�}�.��F�xz��k5�/Z#��.��u��Wf9Z��}�}=�WU�f�NGe)B����f+bb�(�4��?E��ӊ溉���ka�5頮�5���������̗3:����-�:M��km��}�@�^�oLQ!͛��A~� �dR�pXŐ@�>@k�-������}t�v7�F�C�����z��<����=h�[#(J���+�v�� y���f���8%���ʇ���¶�!�)�ۨI���M�k>ҒhX������C�Iĥ��j^"��w�΂�<��?�e�qo�0�#����*����+y9��9�����A��(;t�T�ȫ�4�"4]x�f�.*b��+BI	�p�z�E�!��Z���:�C�v�9t��ԓ��"�r��n�x����{0��-���E����/�yZ����c��G�o��(�"u%U�:?r'	���G 'y�4dp�s�Q��t7�<�ٵ`S:dY(��ܔPB� �� �mg;J��5�D�v��C?)%�5�0z�~-���ؠӀ��S��a~#��`�Y�:���j��M��N3�%��H��!̊t|p���fV$ڮ�68��q/>�C�Q��'ĠP��0�#F�j���`
P�񶧁�kPW��\%�+���+B��1mv��mg;L7��^h!Q���](���N9@v��fjW2��@#���=�+V��e�E�L?��c��G��Oq�V��&��g,�^�U�XH�q$a�~�~�	&��Df�s@}��W^%S�٢WC�Df,�6�^�(}��`L�#�&�1�p�Н�,�~�y#%����23& �P���W`}��2��0��I���dQ�k���lB����>�G�}3��s�A��t��lُDƁU@"�
��zr6�n�l#��s��דH�dM�S
eN��<^�+�x��X.���hm�`�H9�����s�q8k֙����ᳯ?W�5+�,̜6����x�u���CIL~I�U�Z�W� �3�t���q+�R���OR�2����xdA)*����:5b�E��^.�|݂�0��NҌDl��ޑ7�|���5S����F�c��K���SHߑ&�,7VuoH�y+3 =��CsW��x���/�'��ຼV�R� xG^�pm�jaP{����u��$�����1R�T���%Vv)P�BGs�2c��H��78�d���������,���c��z�4�^r�9���]��Pq�Z��myt(�Ft������O�Q͑�,'d��~ y����'iTʔ�X��k�S�S@>z�z�e��lS����#Q�@�>�Pd�2W�+�?���ҦJMvU�s¤�SF��:�a���I ���:����"��7r���B��9��3u�f�k�<Ø�<z�B�(-��1A�r/�[JxJVMPG��Z��0��u������5~��)f���D'x��X=0�>�H���,���x�@}���3ߔX�����	 �*�Z�#*k��W�b4�����1���ݳ��;l�[Mܛ͙-	��hL�71�r�q��\|L�Uc~���՗*��x�o�e<�~�d-+Ve_�gS%Q"���������x}gO�'C"D4F��(��#<�󪃥���/RӰ1� ��(A$���uy�7��I+�ƒV
I�{�e�k������R���q��F~ء>�[�Ռ�{���٘d����'���c���$���p����m2W�F�#=%h�������B���L�D�-CC D��L�5�'81�b���k�+<����Leۄ 0{�&d%�*�F���a��J�O�\����K@���W�L��<��>.��n���@<�'�0�+C΁d5ڑJ��U�hR4���M<3�2�Y�F9ek0�!��c�CI�E���l`���5�xG�CsGR��#��[:F�Џ8���^��H���d*��ps �#i����Af�<�����������n�䜺�.�!Q.����?�S̻��ʻ��WxZ��y۾ uU��Z�D�<u�=�՘��r[գ7�K�6�c5d8������r��o��vT���P֍� R;C"8b�7�K��3L2�^yU�NOX���`���61mR���gQ�m�d�l��YS�����6;�b�O�y:���qV��#���z�R�	e���BЩdG=]׶�ĭ6�I R��:%�*
tk�P/�� W.U"0`#�;J�&
"��%-۟@m�B�����֦�~�/��#��{'Pv$"y]�%yJ�ө��im�b� �����-@؆����M(���W�<��>^��,������]v�:��{��d�&��ϓ#�Y��S[�XB���X�����= "��w�!�?���{Gv� .�Vk�C�����W��=���hg�D��Jkωf���s����%>ƫ}:
��^N�H��k�<<�%<j˶���U8D�Q7c��y�(�}��7g�b<��Ay���������M;�J����ʦ{�f�`�}�ưo��2�L�ur.7�2)��)�p�*���ӻ�Rmz��<�d�{5;��H�'�	�34�	��y�.\]�nA���4T#�`۰q��uΘ>���W��H���=M�78���p����ኽb�K@/?;���=�صA3���KUP2>;�t�Kד9Y;�wzo'B����b�lloPWf_?)( ���MU�?=�(�����ZP:)P����������r�U�#��{�w��yi�t�Ί25�k�+ Q5�x��Φ��9�H��tf}��Y�d��,�s� ��u�w<74u��abK��+��#˸yP����V-́�5 ��4��*���Ҭ�V�ݗ�E0�\�0�N�>����F�U1��p����u��dy�G4�{g��rk(��Zg�d,dC��&DtGg���� �zO��R�cw!}�K�L ��M[`��)��zX����X	#G-vGP@sid�N�h|\����`mKɆB�\#��q�V�!>r%{3-�ۜ�H��W�{ʉ���2��T�����@'�01׫��"�Ƙ@ﰦ��wq~���]���
7$�)L>�7�bχ�h#$�]���1�P^x"���sm��� �Gk`�u��B���Vm/'�j�����3�q6tY�D�+��I8<���|���&��	��W/:�|/�0�*_cH\$ѧ'�u�r�Lk�0���F������9�r�.� �t��	�T��g��Q�k�v�i����Ҷ.E���=�d��|��I�2�=/�4��s�q�3���D9�!�_._�Ou�yX|C�1 Kw�~��t�WO��SMIS|�
9!�J-o�QLP_��d.����y�YeP�D��`��7-s�Xu?X�y�4!�|dR���&�k�EZ
% ���=I��h�~�<�zA��P2M��F�KC:�	�4(}��P���Eʳp�q���{6���k;bu�>h�la��aj�3����)_8~�#	0S�0`���J�qn�N�P+�d��u(��}V -z�Ha��dӊ�	�x6�c6�� n��O�-)_~R�u7�r�%0�ٙ��a�D��m)	���/nc^���V"��'X�wy��["w��v��Ö?���)J��"#��z���5�x�*}v�)ₖ�Wd3�r[E��k6��ou�	��;Qz���W	�����#�z�Y���1����'q��l8>&'��>��yR-�*�!^�Ipi��	��Zk�]akB�0~^�����F+U�e��X��Q��TqF�f.e�MU/��Fj�*tr��p�_�V�/��۵Stq���r��X��__��(��N�N�Ƽ$I�p�/�3�Tr�ɞ���2;ǎ�`L�>���k�7�_O���:�7Jb��D�0�+�ч���"�b���5LJ����o�A!�4����,$R�d��RrL<CQGܳ L�J���^�Ħ����,��W�PFP"�M���gZ�E8��@�qU��CFRl�/�7�#ǁ/z*k�Q�G<�;�8ڂ#�[έB:Ƃ��q�(T_�gމp��-�{C����uY _��b�
O��AH������1=����'ɉn�ۗ�oh��=�I���nHd�9�&'"!(�?�h��ɨ�ۗ.���^5�����C�jsZ�V=��^	�'���=1��@��A&e�j%��fP�f=2ࠐ��J>6lFz���u����䶏Nҳ����։��)r��H�e����Ox��[G(��2������_@����i7J	�g͜Q!5��S���;#/��Fw��'v���K>��Ԁww�)��2�5���x�J��{���L�jyb�'�j�a��Γ�z�!��U]�Z	x�ㆬ��كs08_�8�`����0���B�Ks����&�����(޿)N�h� c��G���_��B�\lH-;�j�t�j*TX������K\��� �6�Zb�E&Ӭ筫�I,���c(\h��}�	�U!�v�3�YU{�����WIl�-�,gO����)����f=f��#���P��=���˲��;��pGz�%XyUGd<����p8��Ko!l�Ĺo�Ch�<R���n�Y+��{��Ǧ�t������u;?�Y
��H���|ǯLʔ���\�S�ʟ!9�}ͮ!AҦ ]��%a��m�e2�������zw�Ly�n*G��γ�J����U�g�Vg#����,�;G�D�fz
�r"�R��#{ڿ�����NHE۾��x���~�xy��FS�]�jb@�σed+񧜨�� ��8��sr�c�	O]E5�2�
C`�ŋ���7��\�m�B�:[p�j]�ϲ�觩�����<��y�3�h?�@� �������Ւ�"Skť'ep�Ÿ�[;�>�?<�Kg�׭����ɼ��c6k�铎�a�$��fg�Ás�^�I����`��A��o���B�8�]C����>Xi$oc�
-�Yo�G���D�i�j���_gvj'/ <|}nb�����U���;^����*�a�uZǝ���N3�4D-piq9�S����U�Z�U���w�Y��J�lNo�h;�wM�(n�,���T��b���4k.?�⠶;��@ q2B2%9@(FTX���i��9�8m߷�5�X���K0�n�8�ش��g�Ɩ���P]���<�V�d�>��ZK�U�$ci�U�[&}wٻÁ��dΰc�����X\�frɧ��\c�Z �����i��켅��j� �Ah`����;0��z�J�p��Y����d�=cr4��Y���(.`4�����_K$#ʒ�&��~�5�mJo�&+����۩8_'3Du1�<ϩ�?N���
W����|���ݐgeߋ|�(m�u�>jn��Ӳ� �B!~Cá��~��焲�e�(:+H;@�C*�L3H#[}	As���L����&i�se����dt�����Պ�]�{��=�����L���d?�`O&L\��4[�U�x�B�!Mk �W��� �܅8	m|b��c���G��A\vj���{Bl���Q�"�$��-P��f>��(<9��ud��&�\��AB� @,0GP�L�����ɼ<)��X�WK��~��BL��:d����6G�'��Or��j�ZmG@~{υD�/��P���,v�#�����]?�����e��_�P���)s����y貒�z&ְ RL )��#H&��ɠ���A���T��x�Gϝ�Ȳ�Nh�y��b�<剋N�/�~7�W�*eȯE��9��D*ܨ�TZW��O��A)�DЯA�Ϙ�u�`@*-j��y���y�s���l�j }֨`�gy
�h�A�,F�Cy�?}%�����ϝ�����ˇ�X�5;m��|U����-�G��'t��'$�Q�L�>���L�#�eޡ,n�Q>�����ꕊU0i��}�h#�p�
2A�!м�&�K����#T��?<�k Nؾ�?�*b)a� O��+V���grd?�M��/��0V�>��I��I���Z�U�aY�c�N�H�uT��*�-]��J�Kɿ��xOZ���E"[[M�-i0���dbr:���kb=XiT������%��7��7U�D�9���5���=�Ld��V�=�K��l�Y3����B�����I]f�ᠦ���%��o�w0�@xX��e!ffF���y��ZU���kxP�;�͡Ecb�)�F
3-?|�&��v�j
�������HBb�!�z����֕Ux� H��n��1��{6c��l>�]�{�f�h�H����ڪ�_M�h���n�ɤ�vI[�=y�j��`�C"�w��5j�WL�����n*�b��_�7�8�uԬ g������d�hL�����AͺB}��'���K�y�E�{s�m�[��l��A�:�V*�rY���8�=��ہѫIC}J�b��JL$'CMy�uq�P������0?ݯP��k����_����T��5���Q5&lZY�vϽ�YX
K����}G�.|]m���8zwsz���&���"�7b�A����Z��8���74q|��� J@$0��ZW(?ʁ��}�_�5��l�[{7N����#k�#b��8�O�:�V,�pu4	�算�z������Oc�ﻲj�lW�.��.+����J�))ʸ��$����� \)LPې�&��o*)};`�
w�-i!�!�4[\~^oݍzK��%��Ŭ.	H@"fh�e�ݛr��ATM����:sb�b���y������7��x��!ܒgq����;�E�_�'���@lt���� ��O����;Y@,�V˓�>��SG�#NUe)Hf�x�1�WXX ��Jl�>˥�w&��&�a=���z��am��b��{��l���Clp�\'C����+�2���z�ČS�ԟ�;}٠�>�ބ����y��������Xaf���1�X�0���]1���)����7�9k�C�_)�!�T5"5�]ݭ�Ac�n�"��v��s�*�����ϲ��%�݃�d�J�+�u�@�����ȜT?![{�\����s��x�w��L+T�}k)�c�ͪ����^OL����!��2�0I�E��a���B�$��\	ɝ����ڥ*�'��2G�F�����{M����l�����y�pB�f�#�"+��aO5���|缲��>�1�K��TdxG����l�n7��E��N����doR�z:���u�o�8���O�|�7�4�$��ًǠLGٰZ�H0a����j�qTف����ϰG�N}(��X�G���}� B<�k ����w��|���M����h���=B{�3�s<��;��D�Z�Z�Q����o��gc&�8y�?�t8	jGg��_���;N���L�P��ϙ�EiJ�ɍ79�7�H�2�Z˶j���Ѧ�׬Q#�Z��vŘ�鞲�I݁�]~u���;��!df�6ǐn�ډФh#m&��E��< ���Qp�=�B�O��d�_��
���ܩ�W=V��k�ibO�3;,N-AX��ɇk�	|��^���W��2A91K��g��=��U�{��1�w㪕�{"�(�l��pr���@l�`��Y������_���/�'	��#u����/���Iam�'�q�yX�{��)zf�';�o�*H	0M'���0K(���5�}Wi%�RjF^� QnhX@L�����g������ʨn�T:�2|�7�&�]  �;Jnvc��L�]4,�T�G#�;ҥHn�ş)[֣��҇��k�gB�A�:����]w���0B�㱟A������).��5��'\v�ӂ2�uⱹ�%�%焉%�'���d���0<+�t�P�,&WZw����&�%�0_��\d��C>��g5cLMVQ��W���`Nw>a��C�yb�U'��l_|f������-��;�ca���ߚ흩��Bt�f R4B:� �O��Yl���~����T�������o�p2�Y�z���)lY�9��j|H�`-����?�x<6�-�ś͗��~P�N*�<P$��w0/F'���*��u(��gB��m�*�����g�#e�����w6���[Z\� ��y�"��Zt���a�# ��������f{�?L�E���m���a���Z���5�)f�n7\V�j�Ԯ7�v>�_����G:�/b05gJ�k�Wc��zJ[]��%S��SG)`1>��D����G%w���pL���u,0��,Sn�,���s+k��/Gݧ�+�%if�bf,N��U��(�Bv��7�IF��kc��w�.�㻌����7.%���&��K) B�t�ni87Q�4�����#���/ ���b4z��?�T�� ��D �4�����Ql�>'�1"_L	$�*��&?O� �r�o��Q�8 -]�&��*
�@"UjN��NoG��Z�,�d�.��S�wVy
�W	�l�a�6�E �d��m"��ex�4�{�)���ӑ7�P�%��������;ݻ�)��3�q��NɆ� �����Z*{v,ZB1��.���ę(�'�*���q���,5�D�ٱhg���;�..PJ�Ǒ.�E�d�(�R���S튟�yi��rZݦ���c���ؓ�򬈪��-���瀔�i��6>�<�z�j=��}r��bQ����zv�^�끇����]���vH�X��;��xf���[��#+�=;&f�8z�ئ��S��Z�S�d��df�����=M��A���zK����L=q��E^�/�Fw�LZ�51U#�"c�L�M���h߸��Z��+w&�~�j=�DNR�-��"�Ƹ����CT�6W�7�	|���VI�Ŭ��x~���J�6�L��o�Pg�=��<�����YY/���Lg��f#(��ʡ�,�t��`��u�}*���H����҄���qE��PieF�}��`���W���A;�tw���ȩ���Ts!��a8�x0�R�b���o$�l��4]�񞆢X��u��%�V�i�zH�6gf���'R�����T>R�«FBm�@���=�Lq
�k��/���7E�ݵ5�ܺ��2IF�2I��'%�x�Z��c���:!C"���f\��3�p�������%��@Wc�X����a��қ�*�o�0����u��aM�r|�7ѾKfC]Sg���|4���r��f,u�#Lɴ:��F�7|��7ׁ�ϣaSk��6��	�J\��A���v�����l�ZD$ʲ��Di��� 9�܎�O����"�3�<�(�_���ꢿ~ ��E~�G�t�G�ݍ��s)U"���x3ʯ*�3�`���d�Y]T����o�u骥�X��&mNvEо)J�?�ZB��h#\�ʴ�:uk�<�.0z����/�ygWH���{�����KQ���[�-�.Ho٥U�n-�y�	���q͹��Ɋ��ƀM��en�iݭ��)�b��(�8~ ���OCU��?h�]��Bb��PͿ��G]D��:���f�����3:~���~���Gb�����^�x��8 jc8ײ�ń��O�������Yv���L�)�PLI?�:�&��Ϣ���w���d��N$����ɣJ�I���*�&^e�cy���t~�� nh-8FJ|��ut~�#�A�R�$c��eE+�{GL�r_i���}���ci_e%��ѷ�R�&�]����&<����۬i�5�ϭ`�����¥��j�R�u�D��3T�zc��a.
UĞ��y�x�R9L������k���� V��@�Y�^_������"��ToMg�o}���Nv;y�h�|�v�wv$��J3Ц����7x���G1.�'8�i:�O�{ܯ���ڧ��9��K�*z���Ĳ�u]�k����0�ݬ�9U��=�\r��9$:	����t|i���d�#��v�x��J@`�f�ℤguP�����<8���BV��-��՛b���2D��>r����{H�v#Kn��B��� ʀ魽U�`|��nY� ��#%�Ӯ�Bj�7S�RK�g}���hċȠ�f	Ѧ����񧓾9R����@���G�n�ii��zi�T�MB�xHu@����CF��fpf.c����9�UGA���<���� �J߬��!����J�Pļ]�i6�s[�h���r�j�/yoak
Y��}��^���}Cz-��Ӵ额0�����ߏ�g�Pm��cAQ���%�ڞ�F�������@R��-��T�����f�둜���h@D(�?CC�cv�M�	��A6(��:�A��8��C8s6*�����·ɥˉt������~�J��6�Rq�<{���qȗ,��Wb(��Tr�=!rZ0����akE1K�>��J�<�a��
���n(6�q�/
Q�H�����T"?gO*��c������������_���m�*����}�
�r�e�	���U���Ƈ+)aED��;���#���E#����W�?l�<>�S\�v�D��}��a�ة��#�۵����T۸�|T$c��_h&�W�/����������o�v���Y��Hr�YEX彨�d ��)�/8���fR��_�v�dn�]}^�	�r��b3��P`��{�����BJU�L N�ENW��2�o$�,�z9��8J�dټs+�6���W�rس�
�0!�H���.�[,)p�`��~ �����b��w�xH�7[`x ���O�H�i/����@,�|Y�1O���{���v���*��j�x����Z��13R�Y�+�g�����T��٥��	���CiLsG����y�H�͢��o�z�*?��x����Pٮ�x���L���?�5��Z������Nq����Ɩ� 5�v+�JIܐAsp��=�)�>&P�!��v7S�����o���n��|"҉��WP�e��Ed|��^����Z�Jn���$P�f9�aL�q4��B�G��01t���GPj��ؕ��tS7��.���6T�,�c��D�AE�o�Sô�9������4�9ٔ���_ب��k�F�m1R��z>��A�H�y��V ���iJ��d
H�y񥕮�jNX�q��<�Qo���A&��A�n���=�aܰ�־u���~�s�cZk�ۜ����O�Ou���R��D��Zk�֧��M;ڧ�.��9D�ƙ��;�P��g�9�"U���$�t�}/NӇ��{�T��tA���X�nz����[q=戒]��%v�ocT9"h��U�Z	�M\H<@�|��i�70���2�Nc�ə�ת�B�����{v�7��
��u�`��Z��2��|w:���CN�?���m�w�h�^�܁{���1����e�5�۱��,Ý�j�(����Z�,b�Hgk)�����TQ ���o�}ImU:�;�w4zR�\�TL�KT�:7�+C�z��$�Re��sCBa�LX0��������<**�CM�Ғ�;f/W�K�/<��f����]��z�ݵ^K�Zf?���w���^��$�F��֟��}?�BTYH�v#x�5J!J��ǸX�w' �H�ms��ǋh�'R���_�=L#*�maA��x{�^�;�Ȋ�J����]B����'�]f���&Ҙ�jD�f���Ll
����!�����{��x�o��be�	T�PtGp�&�y���i������
��-���N(��,`��*}F%�W�<�(���<ҙ ~{���6A��͇ �'���P���|�� �e���f�"N���c�=9⒗�j�'�)��/���-dJa�*$�!�P��7�"sǲ�".d���"VuT�B�-=8{�X��7ͱV����L:���]QvnP�����?�Y�hw;��&��U���G���U��iNEE���A<�ztp�P8dۜ�Í��&b��{<�2]� q'5�5������򚮐oX��S*�K������6�N+���nWy|�$�!��@'��g�+S��ku�Q�m�zd$X>�.F÷��hYns6��Y��a�[08�oo���Zl�
�M���/��C��'vRjg����J���"C<O1�ԽkVg~3e�M8w��9�V��-I"�)�=e|wN�\I�%�f������W��;�#0�'�ok�F~}���bZk�-u���_GԮv����Z��d2Wh�n�e�c��v+g|�n�Cu���*��΄��B�@*���T����TOS��#��3p!�tQMv���m���~Pq#�o�&r��Ȭd�t�(1&	ІBe�Ҕ\��������d0������(�!�A��J���;:�J�ڏ1����}�sDW	eL�@�O
Tx"�D�.�g��mp񁬦ѥ�Lb�ހ���X	>�)�Cz��'�H���y��?�ⲣJ��/KU�i5g�΋���k~��`��z$����u����*0Dr.����:2*�N,#��U�&��9T.GY]HpۦY �<7cΠ�z=���ņB���~6���ED�)�\ 7}<hi�c���kE�_r��H7���
G�xm��4���h���>��}@qg���y=�(�K��f_M�R>!�j+��ʯoֽ�+D������$���'�wfh��E��=���/��6�,�X>�x��0j�X��)���բ��@��52E�𖈦���%\dwi���0TW��y43���T���ȝ�|�������v�%Y� 5�B�e���r'�Qh�	.vw���+oD���8�[jm�2	�1<�tK`���6�������F
 �k�I�� ��2�ZT5ߡ�Vԇ��mj*k�p�ج<�4˿SU��+�������t�m׳պA-�n�PX��	7SJ�$ڙ��Z�fU53�F7���.���P�ܼ����!��/����� f�<:�� �B9Ń����&�j�ȣ�nyEH�/v-#�&/b@1�L���l�8�x��N`Nwh�m� �pF�m&�ʍ|p�4�d���}6R���/8�%$Ja�pYr�B&���񁴀~ձ>���/�Cs�*@3���q��B��Q�����.�OY�/�m��v�>`ßz��D,l�(l��Q����dk2������9V��e_�g�h d����zL�s��N[��(4
l�
˥������7�q�����QV�����	��}��.��R�·?�V1q�؇��<�IH�J���H���3��@�Zn#~�U�u��G���U��{xL� �n�ˣ�m�k�W#�&ίb�H�p�^ux�(:"� ��{7��������由`d�v������h��7BI؆�,���6�t\vu2��X�-4�� �B�,��y�T�S ��b��[��.R�×b�թĸ�8tr��srz�K�x�A�T�M�[(*�غ\��e� �@�麀�$Q����dg)1��0f"�
L��@�qc��=d,�I�����b���[n87���gGG�k=M/�-`Xs�b|).`Bz��U]�Іչ�1���x�{�g:K��j� ��Ǘ�S��G���h���T������㬰�`h~4�*
��Q;�J�Hg��u`K`\�/����/ߧt$�zfИxX�5�ף���[|����3��H!j��C��c}s���=^RG�lw5����E�U{G��b��5�� .���i#.���g�V%�z��3�>��ao$_�yy��_��3CJ�YV�I9߬-z��Sm�^�~���E��q�k�����qm~^�/�	��M�V�4��N͙�	<����@=��uY�P��5�)�������n�{~Ns����ĉ��^����/��	m�C�SK
;w�cWJ�yV
��{���lS�3Ii�\�ȕ2v<�8vZz]�-�O���PP,��F`������i�ti�ٮ��L�3��.<��T%"�L9�>��,^��d���"d��yԲ�bCݒܨ�:�"���:�`C}����_x\�Xp.��<��� :4��;7�O���'�<2Mޢ�n�߱g%�c�{����iv�W��AM���$K��b�!-b��U�j �?x!��iq��_.�a�N�֪ѷ	�wŤr�H�Y��4޷���ԡ��gS��=��r*	�X�^׷�N,�q��Mt�#v-�0����ir�Ru�޶oJ���/y)���ǔ�~�m�@g9G����!ϊ֬�s�ҸW'�UH�!�+.Q�_�����.E�,+���{��ǯ�Z��d8����Me���SՂ�w�ze��H���iMs�5�˫400쟒1�>�mC�T�N�)<����L�4Y]��!������K�S?�<�uJs����n�ߞâ�6ع{@!�\ȴa��Tn?�c��(�TUb��Ja�#�������X���j|\�Ux!@O��Sᯚ�K�G�:%�v�蚯����	�����c����#����N��0~��.{�iu�u�e l�X�4�.�e����"�Ӣ�ε9�$V�e��ʅ�ZL��G� +�Ħ�(��'YNe!#��(r��6M�)��!}���z1��l��rb,�0	�L��z&��M�=����@��ZgUe����D=�7��ݣ��D���{�a,��՝"�Z��5��b�.x�D����+��N!,�Xt��ØJfn�9����.�N�l�O�V���tu�6|��2�k�u�W�$!^�U���֎�؁u/aV�-U�� /ʻ�G�Ш��hF�k�,�4����	�/�s��^����rI��;2�Q�g��w���7=��~;���Ev��j���;�	��������R�����Q)�6�o�^�nڹ�q��c
�ԙ��6�d#��5�-��G�c���3��^	܆�'−s{4����>��R�P'�������x��C	H�Yx�
0As��D�ч�eDre=�p��+~��k�����s�/�`#���C?"U'!Fy�EE�������n��/N�B��A��߃+�b�� ��egټ���GP�F����t=���#ĺp�6���m�p��ܦA.0��H�?q�Ioz�b�,�d��=p�;�}l@ag>P55��^o^h��DH��U'�4U���A�w�gA�.Qa�7�O��LZ�QN��	h���=y5�;��
��η)x%*h�)�zֳ���I���U5x��,ʯIx(�mBČ�g�[�]_)�^ψ�u.����J��	��!z�W5��r<�`�[mɪ�-��dnگR|�`&jSjj�ʌچ���|z��{��'�b��g'����I�U��[��V�iPV���mz�j��؈�s,���虣F�:�Bϼ����[�]���#m"��VEb�s7�R�b"�oҾ������ww�����(�n�B�~�RA+bd�fx�)�#������4e8����f�,�����l0���s�Jw�^>��y_,�;O�C���u�coo2���
S[ʲ�F�?5h�O?�f��>�	��|O�n�[dl*��RB��P�
�Glf��bl������v��V��%z��'��4kK�E*�}�R�%q��g�a#��դE��x{�(�4�S���?G�ճ�ŢB�m==*���k��Q��5�f�����?_�����Jg��@a��]�g�q=!�����Ȋ>�	�U�gF��O:��6���w�#	�I*���piK���Uoz� (��@V ZF�́��Öt����E�\f&�A��uR���u{#6�y<AT>p���]Gc���q�pW ,�^O�_����@��b�ڲ�Q�t"�o�E@<�[J�<K�܄�}-�o.�ka:Α�i��-,�Űт�����������	�?�9|0�%��+�3������7��\Sx��x�C� 33
�X\�t1y���GH���?=
 �{�t �ч�a
9fE����2�v(�H�Fi�A�@U`���ꌋof^���5���P]�l**4�mv�
�D6��h���q탥���i�v��'`���q�L��"��7.��\�C �z1:��%M������&ېk��O"��ޤ�깶3�=�Er��4}��i�*փξ���_�h�ڨ���Q�G
���;2�G�,e{�3���$R!{_�Up�R[##D���ՠ���]�v�0TɘQ��-(fc'alW�"��Fu�y!��9�	���s���q�C�q��91�Ah��|��(�\�����:�Hr5�N܂�>��Y^L
hI�M��~<&W���v,*@4���-��1"�9a,sh0�4CU]6�S�� D�V���{���lm+ =>�>n}%�	+�����;����9��n�/�+:~5,=z�'Nۜ:w��Q�ŧ󮏮Y�|���8��q�֩�R�ʻe�e;��1R���R�N� ����l.��(�p0�����fH.�{@�g�Ԧu����	����'���2.</�d\ʏ��,���ԯ�(���� b�C
S> �Up�U-�'�
�C�_�6 �!B��a�j����I��S�z��/Z���Ӵ��^���[k@�R���M��ɹd�~�I���!U`�d�81���F#�:��
���������sy��� �ke��;�f�I������r8���H���+Z�+x��l�w*1Ƿ�~,�fo�5�$Z{Q�|�Ś3�_�����YU�5��k _.p�&3?I�D�{�Ʃe���4�����0���'[�#g�a���xl܃l>�Ϳa/e�;ί����مW���(��F�~d<��mA9)J�\*��r�j���xї��}<,Zi��_e�	[��7��&X:�_�qg��D�A�YV/�t]���Yx��L�jw���x�=7��@v3nbN�_���6�葳0w+�~5�&'���f�s���҆7bc���
wt�6˻z��2�I�[�C�̾����a�4y�R�Y�ܲ�*F��\�,�`"��X]P�{���<$��h�"V�V�s�F������:�S�պ`^+%�â^�S��G-����X�(ߗ���[P���~S��*%�4wV �ِW������J�����&)��:l�Tr�;�ŹD�l��A���2s�e1�I͠ �����E��y�o�
��ˆ�[/�fd:�v�w�B�|��'(՛��\�E��jKG�Q�D09#�b�bM</��:b��q�+tT)�`B�Y��*�X��rt�꒦:cx&�3r)&((��d��k+�s6|��0|��sl���䪋��"1����Lz�B�d娉j*A��y?ɇ@�������Og���_�a�����Is��+]�e�k���m�����}6e!��"*5rOչj`�M�~a� � �=��������ž��s����A�V��%u׽嵸k�ƥ�^� )|kb%�>]�F,~%��]��L��}j������8�ᠢV��bϙ(MN���[��E�fVj�'�8����5�	�?MLoe2
n@P��E)h�P0��@���yo�[+y,�bCˌ4 c�%�-C�<HBV�G"zx�m*�`M���%��\�Yu&���@c��&���X�6�q!=����-x�`�0.B�:"���o�W[�{E�gDr�47c9�uer��pJ臞	Kz+0�w��BB��?RI)=��p�5�aR�v���>�̎�&kN�$$�G�Q<(�{Ha��T�����'���.�[�A� �w3Ϣʷ�nm��������i ���7d���w���t���MsˇIl|���ϷL|Նp=�$������R����~ܜ��c�l����|LŁ���2O��XEp�!��s��5La���-ߖȪ]�g�o�1��MC�\
`d�9wm9Z�e�/���������&6+�R|�@\i>a6�H��\x�-��6��w�2��qɭS���̈�[p�-�]űW4{�2����J��2��S���x�*7_
|�2� �wA8<�-�E*���V�ܝ��k��x�^=�
��X�O躸K�I�h[�"��C�
&�Nӳ���x��I���F��ћ�����i� xUM&.�A��z�r�
ֶ�� �.R�̷c��H�-Η�l�ð�ЯGȪ���y�ԑa��IP��-�G��o_^]h������w�Ĥ��?
r^*�o����ߣ&a�p9M���3���eh����>�W��� ��w������;��=��٪ܖV/�~�MH�2��.���9�B&�w{��Jϊ7M�CI$�6�Ⱦ'=�ϗ��
y#���t�`�Q7����X��
�=D��<#�N��{��%i��Q�h�o�z�R��Zt�;�6�.%��Cs-V<���l����w�0>���}.���Le8z|v��?��<n�{�_6�Ȭ�I�w(%�������D�'��l��s���U+��A�ȟQ:��&�������q���A�;�]�f��J�X���ܡg�%+2��U������Y�����v{�}^��!��xݙ��؅���8��3����M�!�u���=��Y�	"Ѩ���Dhq3��F�a��ŬOgP��m'�:�N�zg��^EJ�x�-*C:��$�q9�t�O|3�Uw{��t��o�eW�OP.��Ș6'Zu]BS-�H=�02�97jg lwL��T�a�_N�������]���(/�=b=-DM޽��_�GR�Jަ�3��=�A]��<V'e���B��������} u��Ǳ�Sܷ�U9��~d�����6ȯ��X�\A��mL���a�W�Rv��FYG_)�<��w(!�q��lJ���� \�v��=�܁}s!G)��q���/ռ��=���7�֒r��K6�0�U��p�k��{�ǅ��zN��^P��-f&t\�d7$u���HH���o(e4O�*i�5���@j���
ŋ'�`h�g�An���]*�ZFo�z�f��h�**�`
p#;o*%�J��1@�<�4�����vp'�S\A�ai6l���sZ�|C�e�)�з-Х,���D����S��%G��k	j��Ӻ�+�u.���Uv�yT'5N�]����C�C��c���:��p��E�r�}�.��� �.7�R:mzg�$ϢS]xO���p�mf���iNR�y�7|���z��H��؎�#����+��������;��`�ƃ%����}��vA@Y�W�xm��t1�tb�m䵮Uߗ��|�^�I�X}Eo =E�qU
�fQ�U�@Hh
��N�}�X������M�-
�DCL��wV7�V��#�.��S7��Y��C�����2�{"z�:�)"1u������ a"�#g�2k��u�]�ܰ�5��7j��bM�>��d�!봲_Ql�C��-3��ph������ێXv�4 r�l3�����u[_�/��"Z�=s��?�Em<��|���-l���4~Vܤ?m��wO��Y��c'�(�=��]�g�j4��\ʴ�_aF\���,�i������R��LiT�s��/�aAvM���ُ &>��ް4Y���| N�x�W��ǣ��_��ڋ�6T W������	&T[roT�Q̟@LQ�r�1�0S5�7��"\j�a��>���@�*�f�ވ�����ts�����93���-��r��>��8� �<�7��3d�e�p��|&(���Z�Rm_���
��A���ҭH�� a�*�q����^]���*5+��sBQB�|�>�}�V���_���jÕjɱ�5�\Z�K�Pi]�NJm	`I��B�����8f� �KZ�u�J�5t/�^���#5�ڝ�}���Ӣ�B#�/�!}�j��7	S�X0M^��2AQ�*s���a��Ž��|��a� �.�A(�( �LRr�?D~F=�o�∈�����&f�&-��Y��kq�M�Kn_jA���c_�q����Ǿ��F�B-Ԃ{�)�Y'���R���} ������Ʒb��� `k2���Y����RT� {e��[�a/	B�	҇�(tL�,t�$I)��;[�	E���!.����ݑ:w�>�7L��0}Xmr~��H4��Z ThČQa*f��-V#��q�>>����"�#���@WDoge�)���{���vԹ�U�YmM\}wM+��� ~��O�N��ҝҟ]�!�ZC�B�ꣴ��C��)rv
�6��O��uW�d>`�OW�V�xk��r�Հ�u�>D
d���^���v6G&y�LR�l6�;<&���d}�蔛�Pq�lN[%ڷ�X�2�Ȯ�KB#zO�i�斆+!TJT�]��#�dO� ��6�2ӔAs��72�Uv@���擽�5 �t&�H�dw�҆G �dm�G_-i�Fe<Z9�v�����⇬�
�wղ��cx�C>�XMJEXW�T��|4�|�PÌ�}�c��J����,1�5��lC��(�[��"��_F8��e�|�UP�v?�ה�Hw��7�Ҋ[�U!���h����"S�o�6�Υ��Յ�)�e���W�xP?=5��ơ��)����g����x^}�XtwFhC�׷P��*q�w6�d�䧏%lc��� ���"�^�����w0���]_Y�!'�~5%��[{+ϝ���Έ�^�Hп0�nd�b�i�P�P;X�=ϋݝ�z>W���,��o��8���xtǃMQ/TXw�bJ>*E!���� �HE�;��x� p�CV��WY$��o���_�(5� ��U>7���(�1�e�*b���w{$�� �J�
u�|��Tm�tN��}����P�&����Hq���L����D�����$Ƶ�����s���{�h�P�����1L�)�'3���tQ� �Rs��t������^ɩ��o\�_��3yy�O���������Ǐ�J��j��`�\����8�#���9aL�2�SҞ_7\"�"C",^�q��e�^��l�0�9�8S��:bda_scp�o���=�@���������P\��'|&��C6�AB���B�^;�����U=)2��0����eӺA�ǃ���롟,e� ��hE֙�m��+f�Vڥ-=PST��W>*5}�>������\m5,l���o�0&I%����^GÉ���eT?W�$�d��$S/��gB(�{�5��m~\Hі�f�}�$l�8H��sw;� l0���=�+�ցgz?�+�jjBv�s��+�W���@J�O�i.�~��xs��S�J�=JI�p�A���i��8�,Ƴ��3VN�Y��f��`\.�Z��j2a-��彨/��C�;u^�u#��}��֏��cm�y�ѣ���W�E���x��dk^�ե�~o�O��q�!^DD��-���~�]�#��2x�xw�{ D䓵d����F"�?$V��5�s���{a#a�ս�j���&�vcQ�r�(�~�!W_��M��J��4�S:G>�~F?��6�L�g�[9�l��T�i0^�t��Oa��8d��k0�:�ֆGdGb]��$_\
�XA��V�u� MIzq�;����C���K�$�̈́�Ұ*e�o��>4�;�ltr)�1���ܨAz�VBW�9�y���=����t���$�U�[�\�<Հ�Y^Y�֎�r!KߤA�(��1x �r����E�v}����`���I>� ���.��V�����΁��F��~~�^�r0�Yz�㯧��/ �Q���f���H���ڡB�4=y��@n͹�S۷2��i�^b�?��j��ld�gɌ�$%S�����`�
�2HE�`�0zq�c�vB��&���q�;�=I�� ;�8ɖ����� z�o���7L��S�qJ``�]���`ma6y��[d�5��t�,�u�0p����&���\'!��=�{A�22�@�i��j��^!���6^#]�G1��H}�#I�����|�Q���׬Ǝ� x��R���#%�2�A<@���)�p֮��DW���ȭ�ǚf'�
���cf�CXI[�v���C�ܤܗ|!�|�곦6����4�_�%��\���s'0�X<��Q�����)�f�{�\�S!�>���je�I,%��2���c`��g���D���ː����N�:љT�-��ɦ$�a{!��H�ά�ar�rG ���ަ%$�K����:�}6��tR�ej1]0D�i���^�f��ʈ�qi���r8.i"R��}p�4�J�*���rrK���J}�;8%��w���"!�o��?b��~��&[z�H��DrD�_YC���:�[뷍�L��T�N &@��Q���X^G��~~T�%YG���@�B�4`=B�k'���0V�k��[VY ��1�ۯFՌ���;��O�T���j����.A2�d��(ڎ��������1/�=r��d�*���4�����!�Wy������g-�� k-��X�N���Tt	wٽ�[��t�-+�6�Y�C��D�<�OBN=������ ������B�K�n�F,w��{w"0@$���J��H��(���x�S�o��7Z$�S����x���0�뻰B�&�B�&8�x1�>�n���du=6���*Cqخ^\�sel��o� 8^�`̋x�~J��m���a�r��o�E���x�k�F Oӏ��pO��@�D�9h����s0V�~��+�[Cn�wa�%�A�L*�>������X_�![��-�,*��a��Z�� c&��Z�,�I�\�j-nu��+-�zǸ��3�"l�6}+�>�����D�����!������/XMr��%�cڗ�� ��pӡ�9��:���3����B(pń���l5�m[[D�[ـ>4�d�)�
L���~)]�Kn����4`�ɞ�}H�Dʈ�'���D(l�}8�H�uUE����������7ޛ,�H(}g�#@��Vx�@����g��/�S��]���Uk��[Yp�D����r�-��
'Ck�����Ϩ{�H���RW7R��,i%a��L��ۗ�~uM��������CV��sv�I�&���a�_=�_�����Y��zi�� [�.�iO� �7���0��������7�~��ľZ#ܪgJ�ፂ!�7�t:�f�5�)�yE����5�XU<!��j���?p�XX1V��Zo2x�I��5
��=�nYYp��g�d��ؖY�����,;�1��LwsP#'����K�s������I%�P�aw^0j6_�L -�d����7���S>���!��=>d!Y��*��Z6��-�'����ق�A��Z�l��	��FD�N�42m99Ԧ��c�{U�;�0v�:k�Ú����]�v��%�O����������I����5��=y#�?׺C?Ƿp`a���F�է�22L̸�ΪO7 #�����A�U4��F7G'y�c���'�hēv�ޠђk���6���vݶM���Ȟ�~֔��_y���|�ry�\�a��av�U">{?V��Ŧ�}<��b�4`�Ľ�r���A��O}2�e� ���n,�g;�G�8)t�����]8�eR��4��OU���\�#%��FC���Y��(�5 ��_�ڀ��"����>h�ũR�Z��\I�O4�zeK�R�o1���֪��6L�.f�͖bVͱ-�L%��9�RO;�6�=[��d�&�^�FW��|m��0J��/��#�ڰ�M}@����C	�RS�U�]��9�S�^o��������w��"J�t��l���D߁�ߡrHNI��GQU9���;c"&w�bS����D�_ј��$�S�?�f��_<�8���m��O@ud���Ov����~�����7D�u.����o��I��/ �3�v��#8���ݒ�:-r�΢�W)_�f�r���� ]��؈^�*fS~�����uS{�ĳ&��UC;�`�{ik���jjQ��3���*z���
���l=�T��Q�@M[�Y2��DY��/�?mQ�(Ή�OVX�3C�e��Zb��C(�]�=>�ws)_M)�2�:r�����l��Z�N���j����
�&��Ʋ7/�E?ź�S
�a� �Ϡ�*��L�?�0
F!	.1BE�c'���m��y�XQ���zx�S0�Zk��	���7Y1�ywI��˖Uh�9-��] ���ٙ�, ֒w�$���C�-a��R�NQ7�S+R�/�bo*O��R����S������̠�����yy���܀�/3B!>6�O��X�[����vP�J������%
d��9/�"p�  ����|��ì�#�JWJwQ�%�4jYG}K���l���*�Ͳ1ʘ\c?��ݧC�H�\��sv���C�yK���j��i�^_�v	/H��\k�_�ݕac�@�WH��N�\Ϋw�V`�ĳw m�Z0�!$�D�Z�iɠ8�GE�����x��G�z��ى�=1�b�~ǅ�Ҫ3V�T(pB�����E2��)����8��Ѓ�	��-� ��[A],�ݿ��RL����>*x �~����=:�_m�Ƶ
��dz#�K�y�9R�l�y�� `'C��a�( �ϩ"�D)^!�.4L��*�H�X�2�:>�),�/�ɰr�s[[P*�>�I['*[L��/?91�U�S���uF�A��g���;i��3W�Aq�D�bپ�Z�)�����<#Ѕ���B�(��֫g��0�?�y��7?Z$��_8����,!{�v5*$�g�">u^�Y;ʏq���W��Jp�u�~4
VG��D&�	��:m,�ˁB�,|���(.4�� ��h��fl�
XH��0E��O��X/�Xx:564�aR_�P�k��SxA虣P./tf�ip���E\���d�������n#�7Ồ� �ba[����f%�S��e1E�9��Ah?;��l���}I��
��$������Xg����������М��}��saO� ��� �6��4+��Y99U�ܖ��7��a��L��D�O��8�-"�A���qZt`�Q� ���O�w���s������1�����y���R�����G�S���o,ۑB�~(U���2@Cg0K��/��`���L�^]��pH�v��)�TaV�+ş��/~��%��L\�vO�5�0���E(]�ڙi�C.�t�Ƭ��(B��
����M�o<������^�����ˆ��q�u��JC��M�$��E/}�4Y�`��*%��qp�ae�f5 ��ڦ'��A��b��U�[���b�����3�*���jd"N�o|�qI���Ϊ�����gQ�����W%Y��X�X�e-aW��?�q��`�B۠i]����w��Z�.'��~`6�u��a?`��]�YI���n�Md��=(c�C�Y�P?���̟brL�&Xh�yQ}�L�DP�ķt���D�N`�9L�j�C͒���v\������P�m~�8�W1i�-�	֯:�E'�h�R��8�����i�N)VНS��V�@��P%y)-��	�H�4
ΊU�w�ى��g�÷������ ����
�yqAĢ[7�A�� �(��uQu��F���t�Mݯ��l�(�����CU���~���A�t�d|�'UZ�GrEU2�Wk����:�;�3�\�k�w�]��I����|�� ����]�Q��P�5Ao$��g^*�Wd��}���#2�+�����L
^:F�.�M��
 V�*� s�mV �j@ ���u'c9��| z`Kio��@I�����{ �WW�>���XSM=��t����Ǟ/�ݸT�I
I�d�9�x$��_(�!S��`1`��LA��[�@`OQ�+[�Ԭ�шjC�	mS�v�\�bOO��
���Bʌ�Gl��sӃ�2��*A�ݛ椃�6�@'��]���u�:D�j�%� pBw��Wԅ��}���BjΦH�����}�#��+�	W�	�X��
`pCŚ����i7n ��W�k�U�l��K����裼� W�|�����N^\�Q��J�$��WK�h��Yʑ�,�Q'���Vrp_~ܒ�}������L��N��Oa�CY��������$o��=����ga2)�H��Y�t��P�����O5;,�X�	b��ڵXt^��8g�N%OS���n?/K��0���2��u�Yb���X�割��X"����2Ƨ}�J��{�
S�3���$\"h ^m� f��׸����O��M��	q���n�q����8�xXp������{
X��^Qp	���	ղ��8��楕�el�mX �h=\���ʏ��OMZZu!�7���^[I��:����u��^��*K8���,Ά�f7SvX٠�>1���P�27pН��<Z<|���+����!���k��2�8�^���ڽQW��a�I�"�26 �@k��2������Cl�����r�Z\�oO�~F������Zjͩ!�~�1�(�qw>�����sSbm	�9��$}��@w�C����U���Ǳy�i�	��z�
֦K[��}�o���I�9��n]���!Srۯpu�#�����ոS� �ϸ�GX������Pr&��95�l�>8��O��S~��]��vŦg'��^FB�懐@����B�a}#>B>��������U�����N���m���Η��N�t��uy��l�@\�)���hVz�޷C>d���������y,��@�!�k�}��W���V�B'	�jEߪ���`]j��X�J��F b����p�775��;+�+Ձ���q���d8q.�~K�}%L6��+�,�޵��OU�g9��m?�BlQJ�L@cFxyb�K�}��7N��R��m�`�_�P�:��o̿M�3#h�ciX3�xt�¼C+����5AyF= &��]���.�M�}��cd#��+�>�p�v���1U�E�xfZ�u�l��d�?s*��X��7+�����r�]��y��0PU�k�~?�DF�K��dS�ZD1�+sj���|�R��@���P���w��Aɔ��	8�f��b�ٵ4Z9�&38�tk�M�}+-=�f�1�D���@��dU����quo�=+m����59��W���ˍ޺;Y_s�;��(j��[�;�e�% P&�j���C��5����1�|}�gO�eڝ�~��c��]�߱����*M9`ڌ ���h��5�p�J�@�S����:���1��FD"U���������8&�G6�~&��qK��{�f?�@�'q��
�qFzR�f=WZ&�<���ٴ���G'�f��.c$A��a�:DRJ��N���v]zi�We掄�U����s6��^v�%y�C#��J�L��rհ"��q�����6����WB/�He]f|�_6@�+����T�	��ieҺ��b���m�w�Gf�B� ���A��&�����(���䶲J�����H��<�*i)3b_^feU<����Bc -�8`��m��]e�!Q�{6=B,����V|�icu7���*�O?����0�W�_6�K�+�n>�D͒>[���^�����f��'/=	�u�9��-��j��C��tJNmP6�H�5:Of�?r��~4�s�\���������4��2.�U�1)���o��"`o��ajᕜ�FR�r�Ϡhr������.\����I�gw�MP��H/3jͧ�w)��Kp�%��2d{
�^���V�	�G��)D};�e=�������B�!�0����eҍ%w�t�#`�������u� �[��ј0~n�:���yj��a{�y�m)n�x��y�K�#a�XpCQ�5�/�q-Ⱦ,ߌ���/�%�[G�Bg��[�2�x�/Xb���D�愒�͝�qbdd�E�ə�ts�ӊ���$_�i��]�=�u$�]���N �[�/��/�mh�R�u]On�Bbb�,�m�H�BMTGQ!��t^y�_f����z����cl@�}�K{ShZX��GrE��*oE����,ʡ����K(���p�Z�\���`�u�I��PJ�*�7�N�cH�\8-6'6`��r:K��[?���
�%i��hZ�����Ո�i������=��4w��-+�G�[Ŭ�Yyoe]��囟SڸEib�
�(@�+ZǷuv{ fdVz�&� �V�#���k�����h�C��@	�_�4�j���̘��ǎN�I;��?��� ��&������r݃��C���$f��g����B5�f�D2vY(���Mln�8�N8:��������ǖ3|k�ma�9��:���=��%A2DRc�ä=6�*~�Z)��+�Q�m�iqoL3���Ä��ymW�:�(]�h�znok��h{�']�@��Fȯ9�H�;(6�ˑ�����Õ��`��}��z�[�����<��n��cbv�������2�b�Wo1c�����d?��}�2�6�o/�#������Dhξ��\�?-�� ��o`0��cE/�����s]_�ȩHϗP�u�����U���"�� z�댏WK��hn~$���k��?L�qB?T���vamQpp��#'�'a���2I����bWq3�o:���u�Pppl�3Q�L��ǳ(-��YP��E�M3���[]��i;��2E� ����p��';c?�υ{`,S��AX���h��b�M+��@^�~ ��wZ�/�^u�p�H��9T��"�g�z��V�9�|�s���~J�q�nT�C�+�M��]��Џ���O���FۧR��y[G������D���
��mQ���z�|�i+w|KJ�wF�B�b t�6K��/ue�����Ƀ���kT��縌2��>�£����7��T���k.��t��i��x/�f�ͱ�l�_����ty�w)��eJ���&����zχb|����~4XeU*�3٘��=����)��P�j�R�`��e�ި�;�8E��m�S���{�օz���H���$���ut��uq��=+ϋ���m0���-QX�OƱ�H�7�kF��J�]^��m��"���.,������?=�ʥNg���So�=������2F�#�`����yud��r���؋��4�r`wL�S�;{2�H�n �z�E�)�J���T���oR�&��N6�\���]�Gҷ���k���s�߀<�zv � : weq|#�i�q���Qq}�O�S0:Ф�9����25�Vz�)�4�fT
��w�f?�뇆u���yr1%�輲�j_�^�`����>|J�0r�*JlK9�a+���'0k�����;m�vt
�+�v�A'��l�|�޼��d��#3z��sZ2���R����@���ui�?����X�%�Ϭ�Ab*+��Y� �G=r���~��@��AhV,�8��֞�7�(~���	ඩH��+�-�0��n�oGӱ����SK����I,�0��&��c���Eev
��g�HL�W�2�r�bҌ��Г�(�����{!�o�E\����zo\.a��oj ӥ/�q����}���X�>.��Y� �j^�����r0]��G$��!}�"7�nYҎtx��TJ� Z��`�侐�*�?,�"�C�ԝ��;؞.kΉ�-0l��$G �`��20��o�	����E��f�?om�&�C�p�Ƌ=EI�,�u|�B��r#��2�R�����2��"G�X?E@�	W�1't/J-�.>��pbey�ܹ5��Ǆ)��s�~#��d5�L��=��@��,�����o2�1J"_<�������5Bq��	��zI<�OO H��-����}�ɨ�AcƠ�A�A��ɋ�$�WE�P��)�B���.LO|�5�ˌ �#q����S%|�}je���Bý�[;�^G���̚	���R1
���D�pjv ��"����a���nv�?�����Qat`�v`}G,��DP���C�~*��_nٝJ�blv.��x����೟3�F���Uo|�"S���%���*Qe�����;fl�}Υ3R���_>Sp��<O��yp������LHtqMV��{� w��o\'07P<_�����=1V��n���@wl�~�l/� ��	�����������C����a"喵�ө�s^P>��W�D#;�VX{1�ɻ-��@C�<�ݰ�ߏ1�����|��NI�z�I�����t��e��.�zV&1�g�mL�A��<� ㌹��l�4��Mm��V����RhJ�3M�� �k�̚��*T�n���fJ�g�R�ܾ��T3 �$+�D��d�1џ�,�ύ2$1�>K>\�*���ί�K����kM)���B�KQ�:Q�iߪy�G,�u��;>���w�<��ã�����a)��=��",�mTu�Q*�"����hM$���ܥ+lϷM*�k�醥�x�܇<����T�Kih�Է��_J����1����8[�c���Q[��f�Id� T�)޺��������=֩*�S�ɆU\�Hr��BJͷ��T��z44�fY��U��o����NCA�A�`��	Z�����!��>3��O�o|Nt\�x��G������{�/�a0-.�*�;!3�&8��/^k�o��<�5`8�H��ݻʴ7��x�\*Gd؈���pWe��2��
���G��V3ܨ��f4YF4TQd�2a�,���)��?�2�u����^���U�b`���Y�n��o� ��g����k�t���h'��`x�z��qm�4��%B#g�E`�j�9z�=I!�d�K�C�[ˌ��n�JTU��c�����_$�Dc0�p��?u!�Ҳ;��I�/v�U*4�NE�m}�Y) h�ꇗ���HF+Uzɍq�����8���'W
���*�X/�����2|���-1�� #W�l.�g��9x�w�PJҩ+3��(Ի�Yϔ1y����J�����'�I#ˣ����������>�wO��ٿ	�3#���@y�s��T�a��j��p}�^m��������l��<��*�
Ҧ��0���u������/,�u>����~�m�?���[��o%)T,p�B��T�:���rTVE�,�jj����D��q�x�h�!�m�@QL�r��F�$�b"{h���:�&�Ɨ�|�Ym}�o8�h����'ڒ�JU����r8�!<`����D�o7�a�CNb���l�n<^�)�s&�g����I�� �K��۶�G����&���*�!�� ����U�����N�,��]>����B9�fLvb;C��tmG� c��]��"�kB7'jG�c��Z��9s�� A*d�n�	w]r����ֵ܂�(��%��C	N賸H��֬ޡ�-@+��ʨ�MJ��X�5���Z�̼���F�h�		nC�,�n����t�Ԙxj����Ҋ�@Ş��^jY]<QȪ&DOh�k��|p*�KY�_�O;y"h��绨#�&be)�L���ws�p�U��'�|����f��寃�
+��(�}��m�2�C��m��2�Y.���w�Y��i�M{a${z�;�B��v[x�'|Hl
���&�z� ac�M�4]�E��jiG��]Q���8��3V*������~��?PL�j���5Yh�� orm |�x`
��C�.Ė���/$)/�hk4���Ry����4����,��0K�m��^O/$�����H	b�e9Ga� �+�!t�
����b�v�۲ )#R �(�,����^Bv�L�h��G�+�"�v�?���:ѿ��W� ~�' 
�4��!��Ƹ��T�'�p0�������"��(A6"[��"���Gj�(�UZ5-^
�ե���`kYA�E����|�JR �8rO�n~�feǖ[kܤ8�������;�ouW��=@[�X�ʣ�J��AO���}�j��e�'Vt���!��?�5�Zτ�9N��R�M�pڢʇl#����.�˫.��%�������x]��Rw��#��.��`@��UGT�����΋z��Y��H��ǩ��W?������l//�8�'1����&����u��~�������/|Li������ao�t>o���[�����鄸���R=&}��8=�䬲�a.�o&�����p�h�d����b�xJr���֘$y�8 !H�D:�7�֓��
#��QNT�c�ֱ��q�ݳ^߈+�s�c�u���e���z����_�{L9'���:!�8(�xDYh����Ӧ�� œ��Sብ���Mg�& �r��2K�H#?�1I&����M�~�N��,e}K,R\_jh�n0��m=��_S|��T�W�V��H��B,1�u��ۭ�1�S�9�3H�iܲ�I�9H>2ʀz��{�Ն���2���/���f�\,2؏�*$��J�N�6��=�ɬ��֐����j �:[�rt�G�
�#ga��ŀ��+�GvqWVa��舮x��-��h��%'g���Yf����i����E|`q>B�m�#YO��2�Qj��\�������-����j�D��.c�����[P�>nػ��e邢m��]}����zT�e`�=6ܟw��vY;mvf����V�!B�������'�hK�Q;ɹ�m;�O�k��j��y���Ϊ�:�����R�~UL䰋�1+9�}�7��%�)�szWkϘ�i�<�jc��ܳ�^Gq%��r�������k����2��w_�/�ٶR�D��B�$0���V��[���]W��T�$�F�w+Z�g�gL��H*%Y�V��Ք4<JrqF�+��"�J��Se��N!�����F��}ij����_[��A����n+��ߏ�� |�q[�{�ќ��;��%���z�Géd
�~��tb��U�+�IKC��Ǭ��0�
���]�����_T$��m@�`E��&� ߂��ڢ���}�bKN�F0�6���Օ$� r��ܒ[jz�W��s����޿2*nn�N|�+���r -*|V/�$�KT����<n�> �mx��������4ދLo!a�]E`MLQ�\N�n-<��=gM����Ơ���Ѻ�� �n�}h�E�G�np/R¸��v�o��P�*n�_���,@
s���6gsOnT��*[� ���*[�M�_)�6���uM��+����m�ŏ����Υ��UR'ū�k'N]�4):D� η���3v��8-�#YZ'ĹTkxkO_D�ɛl�d�ڭp<�{4h�����?R���^��}��V���/,��-�T~b4�'�ˏ0�\W�5�倐^�B�Mg����<�Pu�����#�h�FI��֗+烱@~�R�+���;���_�҅u�������H�D��dd��W[�Q�RN0RK܏�ɾV���Ѱ�����ֳ�*�B�HB���"�+�Q�S��чڥޑ�D�}��NF�����;Y�Q��l�NY~�LJF�Z�K������UR.�W�K��\R�m���6������@N}�������w�#��[�Q�P\��� v��@���(�?�E�7r��۠�I,�<�NX�{n/�+I���̿O���씪1T�	`W��;�c��L�����4C�R�my�S|�(#=(��� �QC�������7RZ��F��"I���eB^/�?"juy��C~{@�ܳ�C٥��B��� �-�����ARh�ԥ7!x�l[�Ks���,�j���ˉ�g��%ٶĪ���~u�SCc9ȱ�՜=��Ij�������yXB�L��Iz9���)����dM=�BRp�<fj��27Q��v��k���'��M�-��+KD��b|
Csۮ"(8��?�x���Q����ۼ����ۖjh@1�+俗�-	L#��F@�"�����9�fEH��9AZ@��$�Ff)��S�5���4��7$�@�;���O����d.�"C�-��->[���|� �j�=BD���w9+�_l	B�����x{MnΤ�����Y-��T�ǐ��h6��,����$1w���^�ƺ+��x�y0#���R���iθ��sGc���M�C��Z-�K�%��-��F�"�n�����P������
�>dL�i�C@O�}��nC�㊮�/z?���h B)�T&��o6���7-U_V=D��D�cD�<nv��u�kv5�@N�j�P��>0�D������%�i�"�K�R�Ί��5��DE�zu�f��rm�Y=�é�?1b�#M��4O+�L;M-�uH���������=�R4�aķ�+�1�?�,�����vҢd;�~�)���k�er|�yv�+'G���o+��U����}��L���l��lo�pai���F0���	º�+P�D�d��������j���ٽ�"ܬ��&ɦ�a���Eɥ���z:\��>��Ʃ��O}^�����Sh���0O��ns��z�*��~;C�z��T@a�]�q�� ����{J�A~ƭRE����/��h~��"���唩Fx6�p��1
)��P�+��|1�oB`���PfK�5���^�h���*\ʇ,�� ^Q�K�X��h�>%�ky+����ں"�ө�CJ A(�m��*���~�K��2ď�������"���*�"	�&�Q  ����C4:ʑr�X�/�Q�0��NϚa���ZQn(4��c�o���6�#<
�
�s��������RҸ*�D,FLcHC��Yy8-��*d�=QVpH��_:�+���zC)V"]K2s�
RL� mK����!�M��"��s�v���׉q��A��ϧ�s�����a�v��N��\���S��X��Ǥew�cƚoq�wN_�Q��\Q#������AI?�=��#h`5ә�6�H�7R��9�!o��A%i�뙖��p���텭ƴr1����s:7&j4�,?a�#=�&�H2yU�O�?�%�4������e)@����)���g���E~ܭ�͟��T�����'�oﾕ��C�����l�� �~*O�����u��j8{.�� ��t�%��U�Uc~�@��A��h#5�����n�꼨,��<�����h�[oe�j7︳�?ɿy=o���Oc���}"c��Gwp�>�y��0��&�;M�)�E&�|�\<���Z��3i���\��U�	07CM� �$Ϸ��ޙ�w��@:��z��A��r�yR�Fa.���>V�
4վ��K���xA�M�U�	����z.��¤=$�?)���	o{
̟LK�U�!(D�m��h�:+���;�;_�5��8��5����+t�3!�0�p>qQ3�*G�X7A%r$��|�(=[՗K�k�^�bBd��+\��w�F钿��U�S�Q�{�_%���j_Hko���[fa_��Y�o�lX���NH��6�������_>����}�GL�h�� o{��Ph{h�&I������B�,��P�{#��T��b2֙���EW�Ú(�����T�!���s6���FI٘���o� ��[zXm��w��B�fل�6���;K0H�og0���Aߟ���o����3�0M/�s�`�N�b�B!�S��E�W�s/�s�E�ٟHԃ\:w����\^ր�*1���k?�ȋ��&�=��&Յ��A���8<g��ٞ+��%T7Շ�).U�^��voA���|�;���E�D�x�J��:V]Y !�%��?`�Ƕ�Ҽo�p�nОuan�{�p@����ʍ /���m��Y0���z	)�D&8��(��`R�z��jp���ݍ�ς��	�ZX��Yz� �M����u;�v�'^Pa�3���Oˢ�3"/���3	�g)�;I&�ܸ�8{��+0}����1O��T�P�z��T�ʧK#�2,����Bl�i���v=YhfM�!&��n�R��쇂�f
�2�7/��"���j��Eܺ�����]L�����T�EΑD�QK7[�{��>�o�q�*{�uN!�ƹ���`F_�=��H�ܧDy����%�.?�U1�!-9��o��
�C�$���#�vԪ��oB�~�����Ebّ  ۔^NC
�&��f��|��х���˄>ѻ,���Wi���!h~����O�J&��q��ؽ��A��[����c�,=q�}�|H���MCTT���"��vE�,Z]�Z��ɳ�Xҋ�c��Z�R�L�}��P鍾�k�"�7���o�f(@�*u�����%a�gO�à���G	I����z)o�fЦv��2^�"�岶��`լ8��xӥ�{�7����
�<`�h��a�?vP��F��B�~1���(�VM�ҒG�/�>��igޜ=!�dsj�m�4Ȋ^ϔ/c�s5���_��8&��`�3���j`�՝� i�w0��XF��M��n���ݣ�� �7��L\���Ժ��5ʴ�NR�������+�,-I˝޳tGq,�0@�)72�=>���J8�:	(!1t�g���.�tc�^��Q	��ƫy�Jj4�:�&
�\��[������+0M��4����I��!�G�cv_�T_D��@P�=������&fT��i�����|Z���uk朠X�v�*~�`���b��O���}x���!I�TD7H~���?�5�(��z�ƒV����,�t8R�K!��`��[�[��lu��1Ժm[%���s�ͷL��"����gU�[څ͊�'���&_ �0�+�g��_�K{��-y�uY��%�7.�Q2L<����cƭ���%�_��7>��-6�ƃ�����!\�A�i-}��Zl��7�9Ǯ>��A�P��>h#�?���j� k�h��w�r(�!�E��\:�DwD$��;�*�E6�k@����*=��b�E�N�^@+�܁�S���y�k՚�'z�t�*�͝�k\2��3��6B�$��d����W���X���Tzv���㿘���hQ��8/F�Bi*z�+y?�1ȭ�j�IM����c�FI.S�$��j�8"���y�3������/�1�����ok���[��9A�#��m�Z���=��W} ���1y>`��vl���S�Pv�c�H��8@�2�8�3�\ �yٸu�{˙!�-\�z7#�NG!'6���i�hZ��[3�C����+0w��2��n��5�`ޅ(�6�%�Vc�H�y�o_���"��b۬$���+	R��&��w���&�c�Q��d��_h�A-h(�N�1*76D#�Z�#��n��k��O�Xq+|�Σ��y���wR�K��||�g�wJ�}�:�(%~�6F������l����=e��*�o*)ͶƐ�C�_�J�
%FȂ�p�}����Z�N1L��X�$�t���-�����~BPev"@�q� �X9;�/�a����ύO�D�h+R�M����ɖ8;��=b\&�n#��l�	ǀ�y���_ݣ�;�g5�	�<���Xoz��1��k�-\�ȳ��ȯ�f��śE��a�\���zX�E~rϬ�G0x:0]6��hM;f��^��[�Subk�[�e���(�*���w0[	e9�/�&�G�ܿRK�y�7�Cs��͑�L0.oW�l�-y�hu���ݑ`H�t�*�x#00K���˥E�;HJ����8�M�Q�m��=��l��-��
̜_����D\�YLO��[�*Oj+ ��k��(���C���O#��h!��lJ%vT����݀�@�F�'� ?��	ύ�@�e��S8Yx抬�JK[���j!֗���"�.kY�z�]PwW˭HF~F���l��Eh�A
��;!�:��wC�:��������{�,�(G�x�U��'K�xMa˺�����ܸ{ ����Du���8�	J6�����LK#&����ٵ1��HnՔrf%cL�Lf,�1ͻ��$�㌼c�G\�U�O�Ș�,n�� �M "�@R��>9��L���d<�ѝL�-M��(�����h�l�/2L~Ո,� ��ģ[����	���ŧ�l�O�o{�2�K�H2  YZ��uTC�֏-�2R�a!�,t����5���s�ybh�M�#�����#W�w`���D[n�خ� e�l���N�����NΖ+	 +?�<��2�E�o��Ζ���D��2�2���j%��<E`_��e���_T����a~�Tw��g�3�k�W� <x>(�+�О���p��DR�q��>��5��`�GV�����ڗ���5]�4H��j�������8��U@}MAڣ��B�Ȇ/� ��9N�I���{��TY'@=<��PyN��� xkd�˸�HS���5m̸�,dv8�����NK�������;���K2i�6��T� g)E��e�ߒ�O�����hϝB����(x�'���}(��<����v�!(��v�PeE�e̎ޚj��Z�u�~_2 ·�=J�OW�t�(��j��J����!%_2�ZcR��C�o}rBq!f��E��H�����!�7�x���.��O�@+�Dx�����s����O�XM�f3�F�4z`\��8`�o-�}e��vu9�w���]�̈́{<��]����<	�[J��AX"���R%lam����,����ohZa��������|��)�ϥ��	�����A%/��z�� �in(�K�QH����`T���/�|b�q1]a�ޣ�*wU߯pV��%��<f�M�G��U�`R��&L0���4^��ݝְ�a@R~�2��<g�Ih,�=�g��u���9�S]I�B��t�M},����=~0u5Z��sΙ���RL��U��q��9�;_%z�+1���U�?wٳZV�SP��I)/��n�$j�4�L���-���q��M�0솧��`����t��L�̦�sɰ80V/�>���hDla��)�-,5�_5d���}��K���r}c[�daN�-VK�i_~~%����"�,ֵM)��IWp�д$�DT��d��UZ�i�A/3���{~_����X�hY:E���7���]rfq�|��a|�h�R#I�~Ee�h����(�j����{	~XE�fX��y�W=�Bx�nQB<�R����?����v�ZkY��]�I�ϳA���X�El�Er���Іj�?>{��;�W��>3�·`R����Q`}��̷ߝ6[��_��ȤM���ԕ�b/��n�ֱlA����c�D��\�M�Bc$[��8�a��WD��o�>1&�9��>�%�����tp%�>(�eU��e�X���vrxv%�*�"��}���h���7�_���ѳ6u�4�G?��6Q��m���l�5����t���w+�X�w�h�|��v��W�[X�U�K�F���]�8���U5LC��r�a[ ��[�&���+���L���c����[IG�]Zҟ�%�E.���3H��[���CY���MɪA,�+UF ��C��9}��V��섊e~,�fU
P ,�o>��@�P���<�X���?5t��1Ɏ��f)�B
��5�j���{Lu�CK�\�é�b��L,�8P��E�ޗ��{�0�!ȑ㺰}th0~
��H�]L���%N�bW��#~�X0��� �0V�@Bl����p���d�?�S1���{�j�[W������J��_�V��a�����tX"�i_��4?61{�|��s�������Ћ�:�]�ߺs��FW?���a�i3&3׺��k'�{P7���ҍУ�����
H�s��).3�e	ir���Ph�q1���}���s�i���q�O��M�m
8f�Mm�ǉoqT�}`1�5(��� ?j-ʾX
�$�ˋ�M���V}{��/�23�~ UB�.-5Fs�`��|�M\gj"����%x�`�{�	�4�IJˬf�r�����+KJxT�(n>��8�_�Y�$f���Xq�>��p"ɉ��Lw�H�xi��Z0��pF�O��lq���pو��\N�;�*��-�u�Ŷl�-��i6魆\2[�		x���<�h�z~RW�j��1�&�� �\6k��M�g����5m)A��'_����V�f��;������m8IV�=��`Yp'-��o�܊{�#��;��y�2*�]���˔��]|���Ɠ ��i2��8eMx��I	��?�Ҷҟ�<��,�1�ت��PD1|I��6cH����E$����{��R�ޙ)ƐL{сԐ��qiʛ%��CͲ��t��_�ʆ�en���gT=1U���)� {����5�I��ڑ��c`Q�>iU�X�2J��v�Re����v&�0�#�������UO:n �+ſ=ME�&${�-�73��̮�<ό�����Ś�,,nZ^*ƹuo�Q�+����F5A��~E#�Z�Vo����C��Z>�p׾���x�D�@+�p}kk��f��Y�p���l�٦�c��V��EDt�b5;+:<�����\��aЫ*q�
<�Q�b��.�����A��z��b%HuCQ�r�Uj>�<Cm~r�����f*�>�V/I����lM��%b��4����a�����Ϲ-�^M�5l݅i�� ��XIɹ��I&X?���<dJ�YI���K__�*�Af��Řr�u�����Fw��͔����e}�!	QM�,tb���h�Z_�+����Zk,'"�&��dnlzu;�_�8���'�9x]V!��˔�T��=���	`��ў����*Ю�J�x8e*��� J�%�J| m:G��p�Pc���c�k��)��i\�]!U���l���@p�&�K6�c�B�O�,���U �n0�=?�0?����Y+��ۣ��'63c;[��5�$_�h�3H(u|��VO��L*��uY5���Љ�{�����ܲ����@O�gn��
��~4�E����W)��Jt`�[��AC�Rw]hW�q���b�2�8�v�r�_j��+$��CϞ�A��w��wvn��wN�R=�_���f��w�������b���v�;�G��������K��nso��	��ثOB*�/)� �"
�0 S��pehdR�0��I݆z=��n��/w!g1�Vѱ>��=g��My�����W�"�Mib*������.Pֻ"�ʂ,����d� �	V /�Ζ�ƣXR����ٺ5)��_"G+�ex��h|�b�{��.5��	,i�h9��7(���2I.5��[T����2(C�wE{Qn��{��Bx2�Wj�t�ڀ?��c��_�>)��DĪu�� P�Q���#��C�i֍��*����K�@���}�\��vwgn���f g|eKq:���UHa�K�˦����n�,^��)���aq� p�i!Lk�K|c2��?'�ֈ��\�:�.��p��H�L�ؘFp���L��)�'����R������#t��L�����(}�|q)�-"�,��Gw�46��>���a��G]�����Z��s�'�gw���*䬭�H�l�o�#�𾨟!c��ʡ��%ύ%�l`Nl�b���C�+��%�b�3;�%?C�6��c����>==2�^�F�� ���c���;�Df�0ǲZ4�����E<u]�{��I-��|��!�Ʒ��0b|J�tjV�D�{pׁ�l%-���}yx Y��"׈�4x$8UݏڽgD-'m�-wy�<c^�+��|�+�h�X�#�`ǂ�.�:� ��އ��L(@n��yas�r-%�E�۴K��%c)�CM��	H)�c��/�=.��eW` )��<:�i��=��`�B�ؐR��4dμR�2�{��i1H���֋���N�m�<]:e���x,4�[:"q��9�~PE0�;�����u��CG_\�����"JwA�2��/���gZ�%볅�	_�7ǰ�F��ͩ~���+�keUcٱsv��WdW ����!��*�zoHr��~lg3ds�\��Dr�[�˳�Kq"o
oOI��oB�MM�۲��8�(��v�/|c�'�vkI�nd�Im#H���ȹۨ��vۤ7�K�K��:����;k� w�&Xb�3:{�q�0j(Y��YW�p�R�ղ��D��ʞ�{D7lb,�$�a�P���х=-$b���.�oPg2Un�I4�~��G��?���C�HU��3i��B�ap�#gu�2=U8���#���yT��=��9��*�u8]|�"���y������Fq�=�m���G��3�����.%R5�O=5��J� ��p�f5n��ؐ�WJ���=0��@T=�.8� ����Y�{j����¹����^Dh�-����̇D�@��T�R����Xja��d���}���v?�f))lIy� 5��!��L+�sޙ����C����e}�����n@=ƕ�V�v!���Db�_;���dݔ�Y�L�=��4(N�_��'�j 	4Ľ�nx���_}'�-�I��8���n9��O�٪�D(m�]��L��?�w�F5Љj8�/��9�h]/��0k^J01�=[�nzIn ��#�>!�s���_=+�F�3t��|2�/�u�_�]��^�L~ �E}�p�j[�^�_Ee0��.w���@u���2���~͹s�J����O����nW}�?��`��<�Ɨ"�\tn�r������A@[!�7�1�Ye�.�!G�Ιxɉ�*�*�"RL�����*(� QiHZ�^el ��@5V~���d��t.�1������ì��ܪ%g�V��Rc?gP"�n��@�����W�o���]��#A��JZ�x)���l�H���T�d�T^oI��"�2(���V\`�F/�Ӥ�K|�+X�n(L���N��e���Po�^��1�gy@�!O�^��I��q�����@�<�}�n��T��AQ'�w/�2Cv�3PU	ِ��m$~�_���8Z]�D�\�L�-\Jl��#4Z�4'�ߞƞt�_���rs]Pm�P��g�����ZWܣ(�d렾'3J#�t��ޢ��+Vǐ�.�VQ�q�4�v���Ӌ�(�?�ϴǏA�e7p͗S\���_hѪ�d�N�m�#X��Ԫ�\�8����W�~|�ï���.�X$��Q#�L����&��HT2�k#���� �	g���sR��q�5=/ǫ߼/ƔQ.�}���xk�.cd�����vxT�zg��@��V@o����es1$ik�YS��2��W�!�r9��!�p%�6�i)Sݮ�qw<zu���Ș�k�rk,��{���R82��<�j���� ��M=c/�Ѿt�+���_���?^��M�E%L�O5�O�fi��z���P���"E�	 ��|�MB>="���6���,�;]�jR ��¬�>�Yn��o7�R�ɹ����ו��v��P�[�-P��I��M��U�s(�QBUŷ��'� �OJ��1LG��:P���zqi}K?��L�����Ce�s����ۤ�ږ�M���kdg�F��Ԇ~����s��a.�����	��ݝ�����<@�������J�_��)��*���	:\�|3��AUl��Z9L����y�>/���_0E���#���*0��7��f�Z���t~E�1иG*ώS�߳��i�#���q`y2^���C��H;�����V��Hh��)?�z�1"�N��jF0�fC�.7\����e��v�'9m�G����A�"M��<����f[IŁ����Py�4|ͯT����"�eʋ�����(uo�4�3|�}tL}��eC�f�E��nk���df�[�i+N���xۨƶ��dΗ+��^"=���l�ې�hi�e亣^:ѧR��\�8w�qJ�]��;=;.�EI��0�N:gY{���k؆�nk3�8B�.[��Y(�z�s�⧑4b�!_�	��M��'��������P<�>՞ڤ��G�M�����3��վ�B�ϫ���岩y���g���H:���p_���m�ͧ��Zi�9��o м���6�9;N��d,��.8	�T�<���"�&S�{������DiBC
�~�w�K*����7����b��Q�X(Q�f>VX�	���]TQ���|�#��J�d�>0$ɝ�>{�Ђ_&gmt�8�	Ѭώ�Zl'q8��}�ɝL���{}��ʍH9"`(jS�c^��2���`��8>GZ|Y����ｉ;�#����"9�B�����ge�_9R| L���]�l���.��tWƇq�\@��k+_r�8��Y�\�O����9%`��/�R�lv�I�~U4fa���jҴ�su
	�d����x%V���n>9׾1�Y�r1r�p�"D���x->t�vm���Ic�:��	���`w����,P*!�8�~Z�ZyЊ:�MK�_d>܃�I�#CR9Nh�5��`���@ 	'���M�@�q�Oy��rv��OR�L�pt�;�T�b�a�nRgҁ��oc�W�o��T��b���[�j���Vn����3����l����.m���7#J���ʜ��1t/PǊَu�1#��������MC:7`#��{�]��D*] ��{�vWu��(��7so��]�p���t���.B�B���V[/  ����WU�o<��AC�Ps�}�gic�:�K�M���"t�4�1#��(g��G�4��aM_�z)-;���hY�k��}����d���-�g�'�Iޥ�I�`YU�N<n�-J��f�v�j�n�w �Y���x��k�+�i��3l�uג����m#~��Rc��7���T���)t!P�"s�\۱B�w �|�l"c��J��Em3᧗���T�Q0h�����f���F�m������I��^�����[E&5Y.uF���݃�9t��7w��閨�8��4 ����{�zG�9 b��F��+����#C��t�0��4�Pi$��b�z�	�UD��ພK�I(u�,��Ed5��J����1��4���tbz�D%^&�UK%e���������F���Q�+E�6� @���V��T����7{���AC��޺��q�P���s @��]k�7��$�%4ᄔ/b6��w���M���a�"��G�1��R�m����EA��^���*.M��$x�0m�-�k�t�I�4�9��φn���wDO��bF:ɃmM{���L���wl�6H���M��x#��=��1�.֜P3�!�ÜlzNL;ZTy�4�o�L6�O���8�,��.~`���ǂ�����
0��y��ڵ	�~�V�n�9[�y�g3�I*��6)�*���16$�w�{���y�.�/� ��X�#i�ڄp��F���xQ�=��mi�U�?ʇ{�gԧN�XN�a����Dx͓t�@�BL�Cݤh/������G4���Λ;��$E�j?���]JO7�Q�H�����Xyd�%��7�hs�����f��I�L�4�@xq�}���V�%�AN�尶_WSEݫ�(R)�E�(�N����(�bf�����`)��^��ӂ�[`��T�Xx
�k&�P�����Q95s�@4�z�.wPn�ڪ��ժ�-�X%7H�W�����x��|p��E���c��_m/kh��.h!2����4�m�#��v�����2a���d^US�Ō��6wf8� w�Y0�4M�ĖɴE�j�v�Dc�BǕ�{j�E�Ju�SR�Dό:|��=��,��tL����M!(s��X샿�F��6Ph�t�@�`/=��d���'��E�I����voDZ�B�G�Ey��g%�2����bB��?JQ�A��m��R�$����~N��~4��zK`;�u�%oC@��I���ܪo�8������AL`��'6�,6�X�ԐA��Ū��j��;��6"��r:�����{�y>6��b-�("	2�j�}~�@&ntY���,KG�ą�
w�k�cg7(͵m!����^��nǐT�#��4��M��d�
��j�~j��D�!���=4��O'��I��(װ�:��p[[�Y�{5��NH�5@��p��;0�4,�xdu�H|���ډrl}<1?[�v��yyHt����܉�v�#V��|��p$�Q#�Cd���KU+q��e��D;ʞ�F)�#�sԌ�	���W����7�f� g�Ԝ��S-��ڙv�����9�o �"a�8�'G%�V� d�vORLɕa��W-b{z���m0ǒ�X��[郵��ܦ��pQ����Qa_��f5��GE�	m�0�N5r��t,�_��=���o�������JV�����OX���S�z��7d���\�	LaO�]϶�N����� ꧏ-6��dPu��]�Y���C�ߴl�U
���ot p�=��+g~}��Ĩ��H�Є����]w�(R�� wx�ۡ'���h���{�b4F���ޣ�cbE��\��H]�Nz�6},�̫�8�v{��Rd*�ŕ_�	J�Z�� q9�Cv@�������L��Cq�ES�T�a΄wB3Q�Sq'v�m	��G��_��"8+厬&�lӉ�����?Bz.���d*x�ެ�����;�t%��cB��I$�G�b��Ů���T��O���i,A��K���۟v������lf�^��Fփ�X�0aFi/-��S��dP��� ,S��a�2H�Tn��\���+�#+�!˻Ԇ��&ΐ���}Z��^~B0�����{�Gm��2qh����al��Y��`�6g��s��U��"Ob�͞�L�5�DF;qDB#i����Љ]'�݀Pm�1�a򚙈����GRƜ�*�e�B��

C����9�L/�B�F�4'����pf��G�q������������^�h��ej?�,���H)-���-���\5XS�)+8o����4E�����b����YH�zc�������e�<�i�P���鿏R��iLŰ�����ͨ*�-��Z��xF�?��X
��ϑ���ٔ�˚�}w�*ط{$�V'�G�6J�9��I�9�j|F4���[�J��D��Q]�L�C��v�}AB�����)[S�ޛ'q@`��T�;A)���dZ{�^�(�.`yG���?<3���p9��e�/�3���`JX�.�&���qz>~Ds��.�ᘫ
�	��f(���.�տr�m��F�o�Z���$��k�y���d*�&�XU�E)*E��Su����|�Bx�Q/��"�yq�ᖖE�>�
߄�@he����~�*���k���X3f����`�Y��@�58/� �=-�
��U�9#�=&D��l���_�oݎ�i�[�	�D�_NY/���A}�f�ֱB!N��
��O�}T��ls]��
�iH�k�&�ȍ�qG[?���*8��t�����FCj���
�q�˔�b]�m5�Ya���O��5~zw��_x�o�嚺c��ov��F���B����iq�(\ ÉFQ5��jۀp���:��K��� ��r�%�����'��SP��+����p�3�U�w[2*j�Ka������s;��wPz��Gl|�鏐�A�-Uo.���mPٛ��H��J�}�ok):gʠӔ^h��P���掿�'<uz�L4�Ð۬�t��k�����7�T+R����%�q���T�c�9W���$X���(p������5Dm����'�fv�%�Gh,*1Ս�i�\�Yb�ۦ&�~�� ��燪��-w������+¶��ٯ��� ���&LG<��(z�}A󽤘Iv��͹�X�6����g�i�Xm����T��f9�3�Y���E��O�5)f��xǎ���rD��.䬌	p���+�n�q�{�A��D�f�r�K���Hb ~�[Dn��������<��&�)���R�j|����Զ��Uva�YkV��&d�@U@ۜ��8[d|�d�7!b�5�x�=��m��JP�c5Q��GD­�c/%�6٧%a������⎽f� g;�����d�������f�@����@N���x�v.3%�a�j�{�ؕw)��-=�~� d����'��t:$�yp����h�O'��y�vaL�𰖒K���x38��B�؇�CZ����.h��:�e�!�/�<��Mk&ډ���db�,9ͫ{����]6�ŴQXb�e\��:Ob�t�1[˼S���+�ϼ��T0�D~RI[�S��7R>]"esV+]����Y�L<x�V2Lz@Y��4����nu�D���## Q�_���4��M�F��c5L�C�:���\֫�M��j<w��qOx>�:��q�8��i�|u�RU%a���o����c����3�b�>�w!FMh�g���34-�}�/_9�P76�
k	Sb�J[��pV��T�H�	=`�{J/�q��Q���g]���EwE��/7�I��	Qr��^`�g��u���bK>*t$c�z� ���ݜa�.K�ˏ�fl�17�A&O�LE.� �+όvM��Ne��L�4����+3\��V�]⎠���h����j�6�;@�����MK��0�X�������}b��|-꯷�3��a�Mi��(.n�G��9t#B�vүmi�����־fa���
T�$#�$�����rϓ�|~C6=��,I]Q�`,=�!�!�U3U�	����6�Z�?aw&3�J�1���<�M�h�>	`��22ٝ)��-j�ت�#��6�������ȟ�Q򧐮���Q��;�	C ^=bc@��w������*��U�`=M��Y��]��F��M �Q��@L����ZH.XZ���1�}�����tb�8DϲO�q��p���E����s��`�X���`�G�C�#�vG�����"��"�Xex��R�E~�jG.�Pg����o�Ud.��v ��ôU4���V{�"cY���r�'�}�t���m1��z�B��v1��{�kC����[���!+�(ʅZ�dϳ�0��� ��\�Gft>�v����v���e��$���9����UJ"���+}�IАhP���~G%H:�,K�7E��\G_Q(��|�#�?�*�1f3���Z�xC~.VW���WH��0�\�Y�"_�5��$EJ��P|��3��ծ9�ʅ.�LVn�0�;��������rx���im7HJ�
?�
F��g�W\r0T�ω_J���K��شC���.��&k�@X��"�g�#5Z�Y
3K!�y���y�0�����n�c�T$@�V��x��Bsx����BCF-��X�.i�&\)�·졍�����6L��J�T)8������ȷlT�$��A����1�"�c�hX99�<̫S�&�a���.��6���Y�27��ou:�r=O��Bõf����v���p���ܵ6"`j��J,?�J��	oR���	e�����c�Ec���;�nUTI���yl[¹>��u-�c�=�㞟��Ij��R��d�+�}��?�rS�㿸�(CՏ��7�ۼ�<�\{Q1��
��@��W�4;��?�pKm�E���bמ��7i�Ě�H���zv?���2'�f�2={�G_�x�>\
(+0;D��1E��M�����Y��yX�1�RȞ��Ao�<-{4��E�h�~;�8%��}�g`�*���\�\�̯9&(i4Jx������(�m(�����5�A��O���=��ivI�>b}�O]'xr3�qH}�D.� 	y:Qŋ���y����Iz���Y��2  6:�B���>h���@�m�oG�W�	n�2�h�Q������O�d?��Tf��|�%�9h3E�aM�EB9[�0��y��U�q�nğb���(~�-sD8p2��;7�m!C2�;����ԇkC��x�0�C;G9s��H��<�j�+}u���Gz@��i���m�$iOKVY�����i�bw6w��s�bOɡes�	{�L?�P8��ʇ޹������I([N��x�~�	8#{$[�_��t�2��U���+��3��*�љ��
��~�.~�
�h�o�|�{O�׫P�m�9�s�{)�)n_��[KR�5����B�l%	1f�s+<�z���l:Dq����[)77���D�e��?�It�z�7Xd:睆5��z.M¡�eK��S���S�0=/f9�&L�=~gq0͇�H��%+h�.��cI╲�"�UL�6���OqK�nJ����)����/� Ƅ�n�N�'�\�	)(�s<=�m��[�N�j���a&���ns<���=��~�1�Y��]�#������H��;�m$:vsw�Z;m.1�lڷ�m���ƫL(K����jth��L�OuC<ֻ�M��*t�v��� �*�33L#�����<��/%?n�Ԇ�`8P����ً�e>u�YD#�;
K�����E�D���q��� ���j`V7:�)�_1���3![]#>�9j�So�h��B��F��N�BE��%�m�svڨ�N_��"z'���PK��Ն�C����y�W�b������ي)@ ������2��J���#;ֿ�B������.b
fAZ�t՝���x�a�ީSm��/�(!r�R�S�X��:��s,���8��5����Մ� ����E��9ُ�/��6n6���yd��i�)kL�m��&/ �t0���5�j��y9>�	��ױ�T��UP���K�I�>��]�*��[:��e��c6��Y9�R���ވu9�E�({�0�~5�9ק
M�!0�ƌ/n/0��
xf�	T�r�����ֹ+�!#x���/�xd��H(>�����)�6[r���p��=zkl�ܺ�ˁ|���do����m�Z���5���Δ��%���y�3���?^�2m�"p������Цٹ�����G2�4�4���s��ۛ#���^9JkR +-��h��������u�
�Yjf�`IS�����~�ϫ͙I-�_e�,u|B�%�9���c��ӪD, �q�0~<�pͰkx�N���4�qw%,�b�C��>1� Ǌ\��b�3��^n�Ɲk0QT�.��W�������2/OXf@�	X<M�`RF��!J�����t4���Z�.U�秱E��A�z��1��l{�l1c��bt�O���cnw�սb�![����C���e<\,(bĄZ�K,z�g�=p�����`M&���:�S��.�����ye=�̉[���6G����C&���zl\�a��S�������0VWF0��OHe_�/Ň�'A����!�T�����x��)&�����؏�Iֳ�- g�V�G	��fK����y��>x�<��%qӚ��e�H�5r�1l����ϖ�Ԡ8Ǻ5Iy�od5����9��^����]�B=���!�0�3鮈u����u�����%{4i�Z�c�j'P�C��YZ��C&��Dc[�Ɯ45��Dk߄��vA'��{z'���e��9��q\@&T�Y��zHۭ�g��,�[�����Ol�V���E�i8�;������
�md�E��rY�<����0,B6u��� �'�0.�R�� �W���Ӕ�"�~�2�V�,9��L�Rű�;s�;g��`H�7�����y$�w��?v��Q�>M��ޣ>�[��9�@F����.]Ar��hV�-c#���kh�q��o����8S�:B����#&�T2�>�KV�/1)~�%��s�2{1aoq��M�h�H̃�~WGuҍ�A5��`UD���4l�,�(�C��5����+�Χ�g���G��:^) ���W�i
��&(Tߔ;�E�{��n;�QgI˕���W�M�g|�B�""ꎳ�쁬ThC�0��T�ؚ��>Gv�l��2������ԦN�!��"�7���*� 0�1>�E|���9&�p�EJ}1��χ�'"���鑰$����z�7�q��yyN�'�I��rm
��IG|⮪�@��t�F -FQ6 ���*^���H1=��pCW�ґE���i��O_��/Àx~^
{��ѳ��1L5��j�i�Mm��-B7�O�~���*�y����{�%�CwE#�Ŗ�C����vɠV��'�w�����-ix�np�H��f��T2]�%b�7��~N%��T�3ay�y�("j��RN��c�Vѩ��ҫ!�������rI��r��o����>�F�TU^���*���>:�{L~��1\��1��|\�	(ǥ�< rH'^c��4�8Cc�-|��lKǪ�� ��RXxFY���)Bґ�J�S��c��u�N�9HP<0�rQV*^�MT��F�+��5$��D�U��ιÒ,��T�Õ�P�h%�#��ů�� ���j�#1��t7�Q�k��^���G�����{�y�8��V�T4瀞+��(���0E������� G����Lf��=0��U/��өɴ��{f�Ik�p�����
�;���e��� Oŏ����JM������㖈���e�vJ��?8^1z'�r�%ƶ��6�H+��uZ��)e��c���q�W{����Wmh�(�+�q�������Ҕ���v��,�Pv;���<+b��U��-A
�6�d�Kz�D�ô��e�80j&��&\]A�3N�S�Q�j���S�Cv�k�m�Wq��o�3�y+F8�_Lv g�#�����d����E+U�A4�P�ZE^U�c�h��*��F��q����C4?ܲ�|넨z����o��1KU�@�x����4��:ܢTd!t�V�~Rئ(�}��(;��i9Ґ�%r�UȁB[z�/�/��	��W�M�6Ə8�b��D��~��M��9�)G�{4B��t5a��q��V�[>M��F|Φ��*+Y����d-B[��v�bAl|�{SjBB�ک�+1����&�S���������g~�Ăf}�o���9҂u^d\�L�!��6�+(�O�{�>3�=�OOSc>C�-zy�śP�k��U�T��Cx�ݏ�ۓ#*y���I�JY~�mS�lb"#��Lxq��a�_�D�� �	@u(��d0�LA���Nf������2����+�d`�����E]�
Q�-0v��Dh�eK�^�"�! E����!���p�����9j�@#i�&�\[��/���ߚ�|%ɼ#5�_� �2�Vu�y���
;BV��1�7Π)���O�h�0�T	1jAK,W���g��f���iW��)��Faa�gy��9o06H玄�.�*�$S�R�����z�����	g�²E���X�mQ�T漽E�n�*��/��%�]�Թ���"��(�`X݋Ut�$��[��7 ׻�jN�2sTU8ѣ�C�R�%7+�I��T�w��j�a�x���V����a�`�ao���,
�H�<�֛�^�~fĆ�&&���.��Y��YISg��x5��H�N�J¥`�5_��)����sBe�F�qM��D1�����Ht���G\l��e�+eYo�M��#���Y�dٹ-��.޸u(�%H..��S���2��آ���w|l�[��(�\�m%�kS@^={���h���?�=n���Zhټ2�N���o`��ݛ�����|����B��H���U�*ꪘ�w�L�c~�#�B�vod��_��wj�;���i`�x��s��2�O���h����������M�f�pf!l���7�eV���J��nry�5[�y{.%�6BZ��5v�+���`&�5IKW�����w�@��]��1�z��P-Y�Jf��5g�3�6�G�ޱ���	YOZ����W|��^0��F�Y�AXts`w^�����MS2c��Y�:3��/��"�)Y�bn5�_:(Z���T�s�K|����[���Ŋ�
�K\ȍ�Ӥ;q��"�G�B~�T�TY(�Wa.��yYa~�vf��R=�Ku9mЌ�0Ea���ky֫t�z�����K[�W�sY��m�"��;	d��4�(������ݱ�d��~��5|F/6N��C���R�qY���V����Br�� ��e<2�K�?&��EjD�)���<<�vR�_��sԏ����*�������f�G�ESTՌj�z�}3D2|�^��>�q�[�� ��_S�>� �)*�QE,��[�L�e[,���j��(\�M��T!����o����~ph/~M������Z�L�����k���Sb{*��s����a ��޽��D@��_�tc/�f<j?eFl
���c)e��5
���eg5�) ���3i=��o.�A�� 6iN��~�i��4�h�2gJu�	}s�Qk�ӂ�f *I��~.��ſ���Ј�M)/ŧ�s�N+��\=�.��+��CU��f�:o��A�@b���װ'���u�;�x6�H��>�.�'����5���ȃֻ.z��3�!�� ]�L58���s+� �5�+ďI,�R�^�aySꌪ�)���,���o3d	-,4�D���?N�E��ү�N�N~m�ư��&:Kp�Ϭi���i�C�Y�T3��[�J2E���k)7t!��8�ş6|��+���?����C������ ܰ�B�îɓ�O
��H�a�E
�Z��J;"9�%E����2���^�~A��4T�F���+� r�ł}�������0�СQ�K1�|r�#�H���c���.�:��=���=���^�^�9Ӈ���R��e�/J���Hh�WjYo��%�ˍ�sf�K̺���4h�UF�,ż���x�sPZ�ѶŇ��fz(��b��F��]�8®	�]�E�P��ܰfʃ�ss��I�G�I�&'q�ݔl*�Ŭo;B���%�@��֤#�Z���'p�᭔[�b��D"��3�G?�)�s�"͖<�k$�T�����~x>���Z'T�Y]���5��VD�w��HR��WO]P�߬�(�ee�¦X�tEhl5^3��� 2�ॏB?�U���u�)�v��Z&C��Cȁ��l�(�3"2O��F�Г8�x�(�	Q*���G��$�$]��q�.>ru���.�H���{�3�u{P�F��Hfy�˸)�y�����j�6�Pc��z�&N������S�v�p�q��?=튕�K��]�et����J��sQU]�b�O�9�Ki�}�|�8�[n� ZK�ļn�n������0��➕�,��DqdZt���×��k����}g@^~�
�7&��� ��+�)��!�8ا��s%T��n