��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�`0����.1CN`��=$�����U$h�Ű-PK��El�v��nGH�a�n%�|�[���1l:�J0�00�K����*1����Fb� $O���#���߼t�0,�#
�~�9��0������8��;��u���U:pػ���	|R��K�����Ì��e�]��nwo�
�������ѡ�q�\�F@������yt�K��0u����nAaX�HjZ4[��;���M�'��9��"yʌ�� m�g@P
����	���6�#+�$������W+b��݋ړ��L�E��������ow=��'�`O���#Z9G3_���0�݈>�4���>9��b�-�pS�	u����}-~��K)�>·Z��Z9
�z�3S��]p�ϐ1���	>��*�d��5ǕxB�����K�N�|�Q�˞�b�m9����OHe̨��)���ƿo^,������-��ڄ���(�mz����h[#�w��M4�)�8��t��V��00���.�)~\�H�dxYcg�V��>��
E����9d)Gb��3gw��z
�]4�CA���O7:��ny^���c����I���A�F�0���ɬ3�W7��Ƴh��݋,��>ߓ-c2G],ǄI*1�پy��خ�KV��Y�/�۩��M��N\aD��������a�0IY^�����XH� R�x4��.R�anm΄�~����R�|���-���Q[��wT��A�<	�D�\�ak�5�$q@4~���/����S7^i�����Ua�LP:d������t�l��-�'I�}���cz�S�u�����w7f�]��E�W@�^��[m��M��P��)�A�  �=�A%q�^;��WTSP����۴Kr��;��~��U�3#2^(��Uf
��L��������â��.[ʕOM9x�a��Y5pg���l55���z�j�i�8���g�;bH�����D�F㽖�v�w��R��٩S��g���*Hm�B�o/̯�u!M�e��4��x�E�k˓Vj�p�O���]�p�l�H�L*+LE�+�t��6
3�h�QK<)���O�ȖR~7N���ԅ�)�dx^Ƭ�G�pJ����(,�Bl� �\��K�D�,N���L}���߉^�vM-���*n��I����-��1�R1��kȮQ��q1|7K���"YB-������ �I�1N~��$���\z���k�OG��i5tc�
e R~Βr�C4�8s�ՙԴ2�Z`�/&g'%!{D4��HQG�or��f���ؿ����i��&ِ��M�*zq���� ͽ�գxT��{��4�cb@;�v>+�Z��+����0�V�p�i�~��HJ�5��/U�_e�z���_������y��*l��y��_��?ki���h���"³t��9�ö��fd���NJ��a�J8�YKh�
��t�d~�\����ė��[o0^����L)���OA49�s�?`�W�)��!��n"�ܬ�3<295��'>]�I'�+�`�}r@��4�8,�v+�)z�_e�Ϣj�C��$h�3�$�,��ȲJ	�ޏb`�u"��P�B��-����*��ob����u��tS����gB���/5A�d��:�����C�W!��j�b�X�ïO�|0��ؑ7e)�A�U�.�y��kt��p�!�C�a�z$Ϯ��ơ���t%����{�vXds~.���2�]��=k��f��W��	�kp{���h����f�v�P�������yZx����'��v����o%"�Q:���<�[�Wk��Gĵ��À��u��
Sl�>Vɸd#��o�T��va�(�v�3�b����*�}����_{�+�F/c:=�̆��)P�n�F��qϖ&�Va�6�W�f> ��(���h����H�D@�~�߮{u(�~�k� C�'hQ8�$'�o���#n͔=YTl���I,��3}��o���n�5|����~��S�&Y/����9��b��c��$�@^a��H^��"F��L*R_yf"CԍMA�F���awJT��P�5���0��S����h0�C�W>�Wdf�l�Z�q�J�=p#���`Y����=���Ft2b2����Z�"�t����ȱ�s�P`��t��2Qv;�*0au�q��q4r~d�n8I���఍�j~�#`~'�{[m��_"�7*o�x�mQT�$Aw�Ɵn�)z1�f����!��}��D,~e7�2=���M�E�����A�I�����%��=v�b�6�D����`��	����Cp~9�)H۽��h'L� dL
o��	G��kDK�]�Lb����<�[J��@��������1Y��QC��¼������
ܤjaf,�x�⭝���ˤhWv�[V���x|�3Pj6#��#j����~�l�[��f�������f����K�y)���&U���	�ވ��(Ӹ2+6a��X�L����.g^�_mF�q��L<��rTOf��|�|L���l��ƀ-'��l���R�bUگ�nA��y�8KF*����A�AmP��_cY�L�CPK�30Jd�����@N�+n�����,�?M�K/���}9����[�Y������'q����2 F��uV5��������R;І�/G�c�r�AF��윇�( Լ��G֒�W^>�DM����V��f�%	�l	kq3u�&�� E��[NbYϖ�����*ZM��RO��K~5n����"�~nāJ#���-{��G]5	�Z�/�ב���z�׼v$��ذ�';��\ƪa۶�N���[I(&6ߗՌX[�N{=��XG��^�Xy�<�I��@1����_�������?�w*о՘9�+3	�[e�R�@��-�����bb0�=(x�%Ȁ4��=��![��6̟m�re �ش�N��U�w��ڗM�#��%�'� �*��5�9?��]ү���ɡ��0k*9�j����gя
L��%�����P7�T��M1�#v u�p�o�e�]A�;j�?%�?��� �C:�=&�����⦃_��:����ű�1�Q�≯�q4a���e�����Y��Z�{V���#IsB�5<x�dtX����UòJ����zUo��n30�=�F�X��q��3��(��CY}V�d f�u?0E��J>Y�^wŝ�	�@)�s��r��$�&���|��ɠ�y܅�;�ҥ���xz�%�_������D6z�\⍴����Im)0��!@���x����D����7G�i>nx/@�8���o[& �Z��l�X����D݃��"�5�k�NW�-��a��� ӷ�5C�+�Է�rlt�yeb!����f�>����R�88��%P)�5�	JK��8�����Nq��@��~�E���v�w��A�D�ڥ�%ɘ�';��ln��	8��4��GTΎm��^��B�K�J�Ğ��W�S+Ѩ�D��&�,�%��	ɨ5�?����X�v})��ʚj�y��&XOx<5��Ly[��&];�R|�8�LQ>�����*��&��� �!���U�B5�֞bn(>�$�g� <燎��(�_�/��+�X��~��i��C� �> ��!��!�2�W�>&��F��Q�X�)2�~V�l����zȈ@2���itN~~?�ifJڊ��Jqu�ļ �`%�g�p�b��Z"�b�赮�n�jEZ�q@2�^��s�|��&�N��`�kޙv�.�8�7�W�3�J&7+�f	���H�ߚ4(����W��%1� ���x�Щj)|pZy�3��\��$�I/^x�'��)�<>=��t������l�$x���̓���ѫ��G͐m�����^����J87E�O��E;�����4Cs���ރ]�	��)ol
�Z�F�V�3����~���� ~P��=KQ����:m�|���n�B|�c׸��i���%q��Y=�$\��3N������8E���|7n�V�v�:+�ώ\`�FZ���M���հ2.�F�A�s��G	F6�,[=yB�_��6���1}��|���Xk�EX��%�7{���f�%�u���M��w	L��u`���A��HQTq���M�S�kT�b�a���`h ���>�$q����S-��5�0!�/�/��4'�!H&�XӪ�m��� =cz\�@J�!m�Or��l��.�]�iE��Y��vKv6�;$9L���h>�$��<�n��D~$$K��[��q6H�P �G�ׇ�������^���/;�[����H�nJ@S9M������h��J&����B8������/=Mb'{�������(^?'w?r�jT�����{������:߈?t�E�c��U�uU�0lsXYK�f���Wd��4D6-��;����s��:�X���COt��Ω��K}d����J`J�\��,���A3x��7��F=�Bߖ./6��K*G�ΰg�!�w�
]��|Ӭ�C =>���`��$<��WL�?�'`>�\\LF�X�=����	LI�m(�/�]��a<ѩ���FN��z��,<��[�҅�����a�Jw��v=��>3
��iE���}�Z�dw �w�?�q\^|��V�A�w͂Rx�Q����!��4��=hnLݺ<+�i-��,��K$��$�]% �O�dGs�ѺI�o
�M���a9
�h���{��Hh�uG�1�^����p�JzTX8I����1ݒ|$�c(�-<�����x������"G��a�1f85�?��l�nr~��e�@G�RR��$��+�aݭ�K�S�)�9����9&��C�/ی.}H�ɨ�p�A���
ئx�j��埽[˷�94T�!��6���� �S�e��_�����Y�W
n���&}��C�>�%o��n�|U5x ���p-{N�W7�tf� ��N�h�?N�H�q	��s2oU��E ��t���z�y�I�){N!��^B �"�j��`v�ػɨrFc� ����S5/8��Iys��Pd2�*��v��g藵��V.D4Ew��eʇ#!��mB)E�Wa9\�� ��淙�WX����"9��/��<�H��9`�#��6W��ie�Aq��p�ҁ���^�4L�Pm�����sU�|z����(���=]�h�t�ճ\C4���	�%o-����-v���P���
Y
f�.\�t����d؀jTh�q&�A�����fܾ�dЯ*w���c��!�Rr4��!���F���ށ(�pOn4
/	�\z��C�nqq���d���lmd�ɧ���=�lb���&�;{�T��h?�UzN��$8�\�*2g8Śp��/�r@�|³�s�7N��e�c������)GK�,N몮Ӡ-`��u�dw.d������~�3�hp.�E���SO+&��T���|C-b)uH6�u�>�M;�)����vK�n�����;3���tB4�aG���K�D���_�%��Z��U����Yrۿ���^%r��
�s*�KX:.�4�'AU�O�"Q�d��ي�5ɾq��D����p�ݴV^���\����w2�(�f[���~S3ٶf�#���'�n;�m��#G��Q"����*m�p,%m煱ڐ�B�<���gţ��j�B�H�N�G�wBO��fUP�ڽ8�36��!x�J5���Y����Z�a |��B��~�o]��h� �)<��I���<)��
�L@�V)9*�L��ʒ9Vܘ�uS�p��I��A`�w��{��T����I\ܒ����(�>�S��U)��BJ��[3��6���Q�a���>��t�֓���������]=������)�1g�m����ץ�њ��{��%k*����.lA���ۊ�]`�y*ߊO�'T��-u�4^2�#PCyy�*</���IvU4�j��=hXn���0p�7�]˽�U� �Y�~yNf��m���q�jUv��1��D�-6��	@.;2��8�,��"����`X�́���:�fOYL�-�@Щ�+�E8�3+���YS+��JR��(������u�n��U5�*:q���e�`�B�vS!�^r��Z_L�P�<D��j���Xd:ZN$|Ψ��Skԓ����93��%3~3ĭ�A��$�d(���Y�J�XEmO^�������y1f)0|�L0,%S�5k������z�����PU��rF���r�i�Rr�S
�ފ3f���e3yw*U�jq��2��w�ÒU�v$�:�y�9��)��"�^i�i�[�m��Y#��F�_�K���Ǡ��*"E��Y�/b|��E�0�Y���_��=��Y�md��t?��J��~{�N�>��V\{�=n7905J�]��2��~��5�N5D��Ȑ-�gs8���^]�������V������/�/Pk���
�G��=�||5ߙi��C�z�;$�G8�������g0ˮ*]d����~"˴�{���Y��b�a|�����;�]Hje�C���|��.!Q�UWZ�)X+��2 �Eȴ)|��m��v�l��p^��a�������d=-P��*q^���S����2�g�йOל�؞�޲��Um��?�L7���Q�-t1��7
A=T�A��Fi��]z��7� գ�qsh�#���a��D؟�����e���?a�ɮRPA�au����  ������<��@md���t5�keK��h�$��@G�A���5�C9ν������[��4~����,��o��'z��)�md������	�S6A�@��2[�;'���'Ġ0��>a~�\k�f�5�7v�Xe)���s���f��hU��(����P�p��Vx���_�,�Ly��.��?_� {��~�q�+�� ��o�\���7�Sxّ�H!c�����"r���]��أC��e�f=�����T)n\?�w�,�&�H��i�<���ֶ��uO���d����'VP�-�����W"<��f؇��]���gkio�U�����O��y�� a��;��^����%.񱵦��<.��x���C��c?����|��̦D��Am,���nVm���C�f�F���F�֪��u	����)3@�is���d�0A��'n/��O�6�|ˀ<�@)�;3�X߅ Hc���:C��7��~�6ܭ
?���iH9SW��b��N�|�����c�G,u�"���~�%���M�~�;Z�7s��no�^�y�_���A�	W�eZ��aB�oZ'@]�S#�O�NF��JTև�?�՛HC���7&��\�}T����(H��`9�.�=V�"Q�	b�=���a����x����$��T�\����B���a%�H��n��u��ǩS�_��{/���&�F����V,ݣ�$�,#�B�{�������.��+ q�c����Kx.t�C?�Kй�r�\�U�%_ë��ĕ&�:_��X����<�j�d�=l��\���>�I33��հ�w>��-�@3Q���q�R۹>��<�j��+)YM����V��5��K̲G-������ND�d^k}ڄow�|{�Sw�+0'y��X�c�n��svy�\4���=������8�~���K�M��F}��YiLk\�����F3�D{É]������b?J�90��� �Mw 6} FB2*�4n��+-�?�7d�2) �����_\���xQ�����'�(���A.�%������9���%:�1:{i>�|c�ɓ-���t������_��qD]]0�7jcPtWA�g|��`�s'q<i0t�p'qu�S���e?!�ёr)�y���* ��[g��ci��T�:�C��
�p���6c��K##׮!���:�x%��Yl�J	F�L}����FZ?�/K�=��p}�X���K#*�X�n�I�7�#�G!&�˅ԍ��`DG���
��~��a:߃�b$��� ��o�Z�����_��Z09�o1��%u:L�K�H�xr'��cĮ�e�*W����L!��+Iuo\�����AC�����됊T���u`��6�2 �+ǺǼЦ��`SR�5"�͘�^}��ŁDY�>c�o�&V��Gݑ�����G ����`?7RC�����$!��$�cH67���G�w���,�v�&'ܸc����^��-A[���.U�u�ŠL9
��}�vikS?h�>���)��{}a]�Z5����<��k�v� o�~��ŀ�r�BF��X]R�/��Ը'���>��I��!��_�,z �����z��ϑE�>I��Ar!z�>]M��!ޭ\�G	��'stIA��K�y�a+kR�I����QE\�fdV�b��&��Q>Z�^�IZA��U9�y�.J?��>��S{��%�sg2�w�͙�t�P=ܴ,1����-�6v$�?��J_�se �nH�Ox��9�$�e��
���{�
'7�,>K.�h·����0&<��+׮*/��c-k�9CX�VR�tG����:d��ςB�}F3{S�.C�D����۾���e�=``1�-���T[��4��)bX��gp���5dfє�c�� W�r�d��
%����K��~ƜH�&s�-��������{��8߲H��R����7v񴮊�j���_t><Yc�F'X�'%�"�y�L1�k"!�8E	��W\��0ć��)*Xo�0)���s����A�lKt��.7���ߊ���m՟��/�����o��(efǚA,�*w�d���t�@��z}G	qC.�<�w:��A��Ѓ�]�dKG!�C|�9�!�;�0�p�&��E;��� )��ӎ\7�`=LSf�E����R������k_�~� �$6�t�F�ȏ�߄
Ǫ��/�=�l���{�2E��י}�x���%��@�1���{l��''�'�tO��Z;`*���I��E�?4.Y���x�����?�"�)|�]�.��9��gL^F.1�שrg���Ed�ف}�dd?JV����qktlh�	OC�f�~���L�&&Fo�A�c�R���8�C9��buw*:�)���+�Y'0���b�g���-�~�����p�ʿ遪aY�L�z2i�^�2�҂m�O.]~�،YJ�cK���_��G�o�8���n��92x΃k�A��8����/�Va.�ư����Ѹ�0K���1��F��;h�l|��\��8�{�h9/^шnh���\���s�|a�r�t����:�u{ܿ��/l+��Q$gH ��k}�����3z��^�W�� v�7��[�GԬ�h�c�]4���b�t��~R�(z�[<��kk�����_���W���� �����Q�_H���o�PP]dW2�>�����=kO�oh���?�U����a�{�lCI����(�Z֏α��=:�A�|L�q3Jq�����oe���%�`V��,�?�겓��<��H���#�n[7���c|��VZue�E!%kM�ę�xa�-0c������I�{���cZ� �m��~5���!�/�l���>f��GnQΩ�.T�!!x�H�oc�����rq�hO֦�vt}�+Ɖ��ڶB���B�L�Tqp�qC���N���3�b��� .�vD�J�1�	���tD=[�ݽ����]0�9��5�)"��&w���%/e�������?�CL�gh3z���ch+h�mF���*��[��*��'AWΗ37��a;f�6�\2�5�}ٴB,ׂ�:�X��=��ʦ�dRH�P�����r����B�6�뾙n� ?qК	M�J<7ix��������&��"<a�����<H�������JUl!��p�j��i�y�QzR�G&��ީ���I�Z�/yٸz\�FHL&W�n����J��/�ܰ�T��:��Yo��9�V�n�=:l�:�w�n��Dq%h��u����/&�q(�FeJ���옢�m⧲4�)�i����)��(��V�B��2nU(�2�՜�[�t��x9C�7]t��*�ͬ���̍�}[n:���W��]�L��;;	�D �a�7R��66<��v��*��r�L�5(x]x�a(T������9]�,��3�������2>�����m
ht�Rp�fT>:�é*m��liGK#%~�YZ��L�,�9���u|y���M���澆	saHɣ<��gx� =�xP���t�5I�-�|�==�`�P�Υ�ؤ�AቁD!�� ����$���ϸ^5*A�B�N0O�L	pL-}��L�Ņ�oj`zD��3GC��ظ��/�I�0��eGh�)]M��h�u�Л�Ď��p����VH�5Hġ"XQ0s�L�<,]G`����]�}Z�����د�B������2�����4c�Q�1����xVĕh,0�8d܌ $���CyS�;���f=��Ku+����[�Ak��Ri��2�%_W��C�c�T�1�})��+�b�O���L��-�r����M���3�$�}�v��ᷟ�uJBE�?x�	u�sO�z����5Qٖ X"�{�2+ d��*��q��8:�Ď�Rɳ�9��R=`Sؽ�h�O�9�
@��h�ȳ�z��c�p����¬�^�ƪ�e�ᾱ]:�l���9p.¬��Έ6��eyx�����F��.��شO���zn/�̢�^1.�Z�`�e�����64p�d���]Hؑ
����'qK1�KbE�e�Y�
�V_�P��ۺ��`6"�_n�^䴫�IZJ���_4X���(��y��@��Ƒp샬-~�.
*UBz��4X�$˳�fuQ 4$��1��[��Fk��QM � p@u�ZL6j�uc��cs����/�i8S7��=P�x��`���	�k���H4���q�{|V��i�Sa��5u�����8�s	�tt��%�,�yOI�\ a��$��Ǯ�ڙ�ůk!6�g��7/ܸ����eMRZܸS�wkn���x���X��{����Л^�V���(Ҟ�n6�A�;�h�@�x6S8�	���Q�i{����9�\�T�G_��T�ױy����!�,�J�"� 31�^�DX����_�0��Uk���(��R|��=�v������e��Z*y�,�xo�����Sb�P��ډf�u�l�6�n=O�D@%	��(��ɫ�$k_�{�k��z$��gL҃1�%5��&r��n��`�}�_LpPs�o��'yM4�)�[�͋3�k�B��IC39�V�q�텶\T=Rz0I���¸K	���KmrM��^l|nI���{\qd��k+ZR�GO,v�5�C�6�a&\�P��Θ"�������@�ōNe�SD-E�=�ʍ�G̍J�q>߉�z%�3@�����k�����P-��e�#+RJ��t�v4�F*؍Azu亟�O<Ic_�jQ��<�'���o#ğ�O�IB:��g�U4Ÿ$�(���9��Gp$Ipj������C \�ᬥE ЛE�*򶫆��������r�r*�D�Р����3N�}�����G�#4>gǅs��M��}��������|�az�I\����1����3��"-���8�^�O��6�\��գ,<8�d &��J�q�T����J��8��$$!L�7-�"i=��b�$������w�:��k3=��Op��ȼ�I�upG��uǿ>²x��(.R������RJ�ʆT�A�E�h����o���M0/ �n:��y΍���G�7P��i}���şV)��k�,��0Ѣ��n��J6ڝ��ս�4r�R��+I�5�
QwW���n����_"A(A� ��J�Ƒ�z7<�h|�!��T=�P��O�7G��hlk��z�g��"DJ��ź^хp�f<���w� :զ]T�F K�
8�q-��ݠ�h�=�ڿRh\W�T�����L-3�0ψ�#�H7��JAR���Ro̸>F^dW�qƻ]�5��9�`'o����t�]��o�uⰓ��G��,��UU��1������Pc'&��B,����^)�?ņ>��p��Bt=�\�_�U/��7�+��B��9�Mj�BH��x�َ��+�|t��xY��ȅ�z��K�Bͥ�_�@L��JB�vTT��f�)B��Y��d����
�$ȋ?<��FD���駮�G�Zڸos�1�ݩ]޳���B��bR��[|���i���-0��VX6n�$_�^"�Ɩ9Ml<v��h��߳�t	&�nNp�}�R��f�3��e>U'�{1�	ne�Q��&K�,����V��P'�o������
��2f˨�1 ;B*TR|�6s�D��0Lu�O�u4�h��'����%��G��4Ac:PoQ�p�1���~���mh��j�i{�~Z|�`=���Sր�Bi�H�Y#��v^�Ȕ�I0 42g�\��?��˶��1����8��Q���\"aW�W]L��[߈������Z���Ҿ)8�������Ǭ�;��hKY�PS�x����?��]	�%��ȃ������	�Z5 ��e��<����o�.�o��� ��GS�+��L��c9;�$���=+q�����G�x�
y�@��N$�;([����~a�נw5N��Ν�	͔z�N��ҩ+��˚t�E,5?�����]�B�������$T4��a-%Q�A���rb=T׊���N�c+�)�>>���0�f0�9/���R�(�;O!ۊ��C���Cb*���ca_�cQ`��o����z9�Y������,����g �)l�_T��?����}@
�h�ʯ���t:�����$���ȃ����fa�e/��������X�*j��q���8e���8܋%̮Cm۽+�iZ�S/r�+���������w5��Ϲ2��:%�W��Bxz���b���b�]�!�����//���g�Y�2�E��R'=��X	�p�U.���rED)�hK,��?�]~�=�	w�C�`�����.F��|G6Sy]}��+J2�roDM��'H_u��/\c�z�� X��i�d�)��Ē%ԮX�H94��r�����\fԒ*��ah�iD3�4a��»�c�zf�5{QZ�0���XP.u:��P��I�t�Ԏ܅m���z7�l�S$c�I��W�͊��|r�J�^E��n�/��������v�_�P�����m�]�J7���[۾�zM��l؇�	����<S��R���y��8G����{�|�W�����]�Z�H*�"�¯�t���5���U��F�W��L<�u�%6hgR��/X\�9?�D>���\L�m����8�ۘ���5i1B�JT�ؖ������0߄� ���W't��ǈxC$Vv���"��wuC�%6:L�|�!9Bc��_l U�)��5ʰ�V%�	����M��Z��Ns9_ bR�ڏ2#&���U�(�6ƫ&�0E���cw� I %+ei��gg˰!���>F+���{��э0u����{^gux��<v�Hτ�dg�Ic ��M�Y�-�G��	���94v�TJ���U�Öẖ^u�*Z
Dv5�/7mʇ���3˴�7;㷩XR	y���Arm^�^@�tHf=�?���<.�2��H5]⁮���/���l�#�A���Q�T�,�o<\��d�O��`����L���:�ޖ��A�F/�"L�z(6Ӱ9̷zJh��I��B'f尡� C��7����Sނ�(ǆ;�����bFG�8��uD*�d��ye%2�@�I��B��6��uM�j����7=�9�?�16�����^��ؾ���zQ��1{�Vu2�Wb�Gy)	7}]zBXX�ٱ���/9�U��u
���ܾY����r(k�>��p��o��@�������=c�X��˃�t3�^��������&I��꡷�]w ����"9D��b���}�N~��Ki�:�La% �Mn�tH[>�z}}����p���T��d��=�a�+��T�_�Y��`�����p�.*��\��^�c�d��$��}�r�k���9
<�]vɌʤ�b��e�:�4�|k.��V9R�D���b����U��Q�!锞�qr�_�����!��Ġ�����E���<!Q���\Q����M|�Ks�Q"�'�c������AeB�����e���GC��Qk@	(�cQ촗�J>�=?P���J��e���c��*s�7�ŗ��w�&3�L�S�=�v��rB��N%����^�������]��b-�a�-Aj�ϔ��;��P�k��'O�<M	^zӳIN+�#�v�l0O��3�����s��c��_�,u�\��E#%[R@ڂ��*]�X�g���y���p"�.]$��/�'n��dF�9(�g��-c�p�;�a�4<�5%��A�.�����н ��ab5{'��9z��'C�qj��g�v�LZ��qugr˝ϓ3ȶ�>��l�,^E�i��!{�WkZ+$H�W�V�x1�sJ�2܃G�'�����/�΂j\Z�P�A��|�	art{1�@��M�V�Z�4D;-�i}��h�[�P�/��ka�GM�)F'S]�'msz�[/=����p�EgĠ��`T��
'�%�V=(�x�K��~P�D�'(N��E�qU��{�v$"")X�So����ӟ��֑p�PG�.k5@
Zc����
���P��)��Ɏs］�ǿ�R��;��$F�l]C��~}��&dwa=\N ������4���VBN��<mJ�wҵm��)�1�>p5���&�j�t.�Rs��i���K�]����>�^����ٹ~dX�s��"�ت���ˍR��j�KYk�\�wᜇc��׼x���a�#��](g:t�:��b�����݋�%Z0����Rb�)zGC٣�����ؾ׽�~q��ߘ^���r��Z�"tuK�]���)�ǯ��a��2y͂��AĊ���Pi�G�3:>j� ���Y��a4D��)�?����~��&���^���w�2X������ oޓ}����P/��/�\�I8Y"=�ʚ�ݜ|�ϡ`w�!�O��LH��\w�B=!5��T�&����A�8�W�5;�;C�lFR��m���L��Z�sC�2�GN.z��T(������Y����%9|����C4����iɩ�U	jy�]�cR�;�O��� ��_z|��I��o�:�J]���3���X�ɤ�A�(��j2�o�}�WH�X	�^ٴ�Ri�āz��X�ꊤRyx�>T��0u2���_�7�ɠ-��ׯs����|���K�"9d��W�o� �v��l�UB�����è�����Us�s�`�ygif\��?�>�_Ѐ�Ɏ$ĠN�`�>u�<U��.�^nuy%���;iH�A���)�A|q���sG[���������6�L��P�n'�f-iEk�U&sU빗�|1�p7ݓ	X��Y���pwB,�����UB�a��D�]���G���$?8���䉔iz>J��*�Fa��>�$�}����c�6G�4�Ey=K��Ą��Db��b�b�Od��!88�q���s�MWI��k�������K��KC"y�.�Y��uGWք�\Ku̳��A���5d��kh(q[e!�����B��,|<^ל������&�78BmRŠgZ��T�ꭘ��lMa�fI��9����@E�/&��R���g��(ʀJ�w���l*���;z�a�]���x�ظԞ�z��"Is���W{��Ѓg��Z~�����w�K����R�ѩ(�PU���������_�B?fg� ҩ��U����}����FFе���t��\ݑ�L�hBeB�,����4�5����b�	�v9x?�o��6{��r���<�i�=~.N���E�v�#h�����Dm��E��R?�
�z���9�y�>�f|������!���o��i�f:{�ۡ\q�)��r_���x�#*w�Y^|�ޅa� ������v-o>�����$E<�0Ǿ\wD��#�=(m �U�$�R�Ȑ1�7�"Q��������U�$�ξCrp����&.�J#
�������+�Rx���0�(�[>��h�
��#��6S�o?ab�I�8��-#�y�Ԅ�t��%I�'�����rN��6�[S1=]�'O��n���$���ig�͛���m����%�5�k�]��L����� ����x��&vs3�4��S��l-�����l�'և��G��!�%�{�[��6���蟿}��,w��R����ĕQ)��7���p�DX�ϐ�R�,�kO6u"e'u�����l�X�Rʝ���b�,k_��h�]�Wk����?�-�۪���QPtx8�3pb�F���@ܗ�Y��+Aظ�?.H"���G��i��5�����a��A{�x0)]�9��:��U�3����6���m�����kەa�vymސ� �s�9��{2͈��JդͶ{:rd���ZA6���'�Z0�i��0[8�{^!p�_�=�lj"des����*�E��A����Y�c�m_m�
H���I�R�/�
"�K5z��-�?�EZJTI��U6�`���TyOFa2N��J�n/���5U�2�ъ�_G�
�]�I�ݐ��.4���GH�`*� Jg`��g^���
"�ߢ�6�[�Ƨӌ ~���g��>	�4|w>���ͳ4	t�h�q�O�v#YV4�̨��&�!ǐqݐɤ֣� e��to�Ěo�f��v ��_�z�ܺ�Y�J���-XE{���	^�����3*�i��� ̦Ⴝ�7�� �҆#�~WE2e0�͈�B��0iL�?�~�6\"�*=R80o@H��YH^�� �*\Q9�A^����p���DȨQ1|e!�>J��J�fY����c�w�9)�G�S�f}���'ȧ駹�cN[��[^�e��k����NA��%J��Mƀ�e�k����z1����[we��[i����iI9�j.�s��B�>��"{��Q�����P(�F�NVc�q�"��:"'�显�*�Ef/��[�'��=H�F�ÆBg�N��lF��\66���4��&�����y��"����\�N��c\��aw=�z��^�_�#t��o�i��Y�(!���ޚe������@���֥����|Ow]P���玞����[�Kr*!s�f@�m�f�*���� a׊�F�D0�E�Ë+ӣ�yJr�K��P��.x"yzU�*��e(�w���W�=}N��̑�r�58ltY��&��A8���mz���5�q� =Sh/w~B�1��E*��3#Nr���Uudl1�Թ�ַ��~� ����J�,����/	-#��"�nm�f��*[����g�6_���<5��D�x�V�ͫ�H�j�*�1��&#-u�V���jh�N�A&��n�d��<3����;u����5�'�u,�94��v��uC�_��-�Cp��������H��!ZNk�%�=� �.�j�q��JΨu��2NoQ]��Z�a��!��	�"$Nb�"f�#
M��Ya��m��,��8.�5�'V&�˱��;E���\��\�&@%|�4�)$Sj���+���M�V�����
G�^��~�tGއ��\��\'������ ���
k	�N��(��x�<�4�q����:�E���Nb)�+[��p=�L��Qh0�Bm���C�,��(C^2�M���x��n�����g�n�� !"�[��,bl���&��"��7��J)|-�z-Q�� 9�9���ԕ�;�[06������D&`�0~$�p5&c��p�?:t*C��ܐs�<�t���N�-�*���.?��Z�p �?�P%��Ã��L�=R&r�\��4��]���."�aZHU«~ P�8��RN���thN��zt����*��E�˘mJ"Z}:
K������hgH���\��
��n�����hІbƢ��zkr���y���	q��	�j�����NM�| �-�`�]�6v�⠾-`�v���x��xDg6���l�].<1CZ5%��^�Fh�ʇ��TL�r�8�d?`m��w��|�Z�]`u�{��e�Ċf��ϡ`�hР	Y&g�6���Aĕ���D�����yU�|�J�$��|at��OB��G�䌢�R�w��O�og�r�V�y^���Y;�2�V����y9/z��c1H4���p�#+*�X�������ߊ��o���)K6hp��J*4�{/�+���o$����>C�	�`h�2�3��~e��2y� �퓲�:���GoܷX�s
��{{��h8)�50�"�%sD�ۜn��tF��7ݮ�R�n� rF�ْ�s�I�J�y֯��*��{�>��r�%OO{�e^���
ջ�A���������8U^�bt`a�@�)�;6B~9�� �|j�����eS%'1����j�H������(&	@�l/��XABޔsG8+�R��F��h~�G��V<u�'�k����V��;�k�2����e�nĂ���/���m����"�1ɬ�C#����o�e;�������� ҳ��F�K�-�����+��Yj_��s�ctodW��:g��}d�FƩk}
�Ɗ�]�S� &0����)�G�ߣ�v�4�(4Ã�t� �h�=x�O��c��R��O�[��X<��M�h?��G&��*b�U��1���U8�}i�D��}kQ������3�*���=������W.� �ϥ����o�2}	5�h3�B������Y��p�e��^B,yZ��Ψh���������0^�}-��	�.��i����Wv��K:3���= ��.z3 ���+�GBC�j�T�l�� �0EFd��_-�C��HрⱞQ�K:��s��S�@p2QqБ�� ˇ`d����s��u����Vk%E��!a���]e������h�%�8�F>���-	���:����m�����ՖX�0��ѿ�~�ح�Jr��Btb��tb�9n��f�E�\x��k���r^�w=pw.�ц��,n0�(�=9�ǄL�y�fMp�PRk�F�z������A�2�5��X����%��$+��[#�̕�?�]OYE�����]�&�׈Ґjo�,�����ō�I���8#F�WYbNQ�p�"��_A�\I�5]�:�d��3�K������[�Ər�Tp��1K/��l�����G�]�P>�%F�I�E�,�^�΁D3z1�E`���{��7_Y�����T�h\�t̄^��|������WE������3�X0P^��%�T�^v_-u���}�t�5F�N�h�w�>�:����2zsyC��t��=�~�NT�+	�ǀg�cQ�9)�F;����:A���=>/LL+�D?��?�1����V�`QE6���CP�4���3P���lH� y����rLO�Ϲ4��Ϸњ�j�[ɿs��}=P���1�m
dw�#��n�t4��wn p"��l1�鰮o���e�0��Is~,�]؉�âm���= h)���t��ez����C��ӓ�
�3NjЃ6�h�񍬁/l��ycp�z�L��*J�������+�\{ǳ"Vt=,{R�s������M!-B�<����t�8S��~e������@'�]M�N"\v	Dic><����A�O�= *J��{L�xA��#�5��\5���PEi�|���߷X�h�K���C��Pt�vno����3�3������mb�X��ɮ=�P�!��ʩ2��5+��-.�g��~��P/�{�� 3	��IV��R$k!̆��_�F�J�Z�ϛ!�>�|�c��'�ԟ�DF�\,�5*Tn5?߷��p�;�Nw�"�
�1z��$A�#�z��/�䆾�
�<�;��<)w�Q k�b��i�ƺSV��z��H�����p<��~Q:��=�gB$�m5_Rȵ7��%r��٩֜�N5fe����,aP��}�|�'�n���	�ZSeZe��ys��b�^.��u7���7�2p+�T����� _PM3�Pf� �#�k������3t"�-գ�\ӧ��:�G4�81���V���k*N=��ny*����i�u���гBG�	ǹ � �`8e6Ww�����Q�-%x�n�����n�S�2����-��5��Ϋ|˥����1Ъ�� ����VdC��ռ�&����T�0�:c��$!U��;:z,CI �0���!�U`g?Il>�eƑ��A�	Ym,O� ���̔�p�����<"&�_�L��	�/�}5�=�'ɉp�&J�Q��̴h�5���g`J�*qZ�c2!��{�*��m�5��[���H/����͕�]KT��ɲǜt�6 �����Me0����\������Ԧ�_��_����k��yl�_���^+��b4J���z\G'��܊���7>A�~[�N٘���4Tq��Éء�S����^~���'#]�Ȯ"E[���Gc�;	�6���eId��\�ՠ��M|@[3�ü0A�EtU܌�䊏|_����t�p�^e�����y:N�h�*��j�j�A��p�zy�5?g3f��)�LK��1�\�NV��Qp�]�#������ڝ�b����0n�� ��͎��DdDTL'�\Yd)O�����}Ը��׀,;_���A��R��9~���T�}�^y@�r�����{����:%��~�Ao�4bC1��e�eQ���O�ږ[tU�g>D�x<��1
���6/:�Xkf���B�>1�����'�{q��f��d/!�:�/+Q�'ā�q��'�an�U�Ը�� ?����bG�-������1NWy�&��lXxG3C;m�o�谙�� .�I�  7�Y�4JH��l%l^�ɞ�q���i'���ru��G"�K4%�j� �?&|�����d^6�~��m7�#*��lO%L�����^�����]_����I��8ZG�9��#� ��XcS���P$%�]�H�+���#�y�4�/���v`P��1� <w5D���r	�p��O�\�J( �&E�i�0� z<^RR
���2��K��G��I��It�XQ��ZCbE(�nҡ�6�`B&n�\"�녪�ܣn���:�
��,ڻrD�6^�eV"�ߣ�i)���{���y�ܙdA�<�uo��W"�c�C�4`5G/�~&m��=|{,<p�D�O�g����qt,ͮ/3--�����S@<"҃4�)
�=,L+�"{�j?v4�)ѣ;&�&��v�D��� �ؼ�L9��L][���ԜV��,*�Z��
ʠ[iF.r���Xʓ�\��rS�����>�A]���Xq�{s}��ME0�EUS�2��)�m?3]�^�����n*���y������*
��;QjX�����e�/����p�%�-P��8���@�[b�z2��}I/�)��U�u�'/�����qr�ɞv���JV�S�7"�|�\U��S�0Ȯ�D����I+�et��s�!m�3�Gr��#4�
�gN��a�0�hv����o9X@NԲ]~`�4�Yq���?��IHpG��"��~�>�U�:��g_㛱���Q�~��O����R+�~&�����Kу�n� ����u`9
�	�ͯu���%n�� $�� �N���>�qr<TE_mAH�� �����g����k	���a���F����l<��w,$���*HP�z��|��\�B�A�%�Yv)1���`ף�E���џhQ��{8��ܨ�8�d��6�1P�X�'%��3 mVJ�"�^����3W�B�sv�Z���G�p	���&d�0��6���X�0�O8S�Y�f�N�R^�A��.�K<z7
e3s��q��m�oo����:�°��❏à@>H�S�ѡ�`Y%�4;�������
�%zQ+���`�]F�v �J��W��v'30߱���)tX��g�G�"g+��H��w�6�P�>#����.���,t�B2�}Z����Yު�րS�f��o2؀�dژ2�ߞR���2ɋ[k�Y�@.(���佀G�>�V�`�߂��~����s`é�N��ڬ�������_6t�l��G���
e}����uU%���%�#�ؽ8�:w�?����8a�:WC�z�#ÜE!+X�R��0��[��bJ�W�'`M�&o� �FQ��t 4�L�N�x.��_����� [ދ!`N&�EM�rj���#�m�d�9sd^s�������.t�K�;a���gjԔ�ѳ���������HDf�;}�@�P᳙FP�w^�g[\��}�^h�9�ZB�5�.~>��ó��S�0`�ȼZ଀0�h^��<0�ÈS�m�"Jx/�1����]�'�]�ioj�:���_�X�3�܄��4��"�S��4¡�;ƞ��Wh�ޣ��U���L;�p��� 9�d:�}��.Ȓf� �,�DƦ����a>������tל!O88K�l�3Ǳ��$����fP#��/�./�[>"��+0��r%�ʰHUL��e�9�{���������kB�>&Ss���;��Jp93����'�u"	��=^������C����-�b>���B����{�!��Z���1�S���jD**o�GTm�#�"�~S/yLf�/��7!����ݟ���Y<_ڔ��<�?�ߨ�L�G�m�n|l�Vk�Vp�gy[xT�`5ŉW 3�m�$S+;��-.;4�T=���	�xWni�kG��
��z�q��̋��!@���#J� ��-n�O�U� �����sE��W�C���ņ9�z�ιF�mI:�ǔ�0s�i$�rgMщJ/�i��-خ�6��}�8y�W��J]�T�`Ds��iU`׹`!$	���l���2��_���E!;^&����Køz�)�����O���m0�w�*W�y��A�0�IE���ADP��
�P�i���0qK ��Od���>J�:�e#��>�uM���]�?��?�� �^^p���|�u��G�L����H�#:ːq�f%2����7����l��a���c70�``J�j�Q�����`�-�A�	rW�~5�am���7�t�����~÷��e��Q5v�S��F�KSL���,�r��c�wf���U�+/N�/�O�#�F�$����ݔc%^t���g/�|����O',����V]Δ[D�,��Z�Ph����E$ʯ >5N&� �noOM2�M�H'֎p������+��*^��5
�Y4=w`�4��T����2f����ײ[B���ۆ.ǈE��[1-����3$�QRB�Q�Wx:!>�/H��f/��!�-�;��CW/סr�ls]Y<w��	A��R�T.�#��E��bg�ZNh���:�<6>�id�ϖ|�l`x��i�}��j'����
8t���׆4\��uW����Ԃ�_�i��^S�O�	d������{|�6K������j`e�*~���'��>V��k�v��o������.Ԝ.7[U['����7��J畇WV)�����kӹ�X
��I ;5��{���_Y�M����W֓����T:n�8��(���ָ�9�/eB��;<����_�װ&9NkDm0ɼR���[b��g��}���vG(��d�<���
�32��EY�@���Es@�<ciAA�m�P=�d��¬)M,J��xx�2��Xi
/m�|s�0�ǟ�Duӎ��,�D���8�	$L�j��~��%u����0�kb��4Ӎ�8#2�6���1$�vp�
)��o�P�mP�����{
~��(+�*a��߳Յ�~~PIxC��;�����
ŅД���C�Q�%$�e�{֯*�<P�@j�]*��
�E��+��#��o�O���{pPl�W����)�h �0���
�,��h].'9xY�y	I��O;`�C�Yw�wV+CB�� �}�d&`eʝ�P�2�w*���+,���/�b��w�`-f��f*�Я�����3��|(2�>\�3_�n����`��e�{��#��NW������؈O� fĲx��Ȩݿ4vՄu �J��B��uZb���i��� �~3���?���Y{��%��D�5�m�/����t��X���Q���}�� :zF@�q1�!�ri��C1~��B�����d4]�/��F�������z6��e�O���t�P�9o8��E�$�R�Gw=5l���1h�y���.�:�DY!���T����|���/�l�%���>�@,�\8�߯0I�B�4���[�~[�d�L��
[[��UTA�<YY���#�m*�S>���d�<ʹߐ.F@�}��Xˁ�6�3�\L(ݫtr��B��l�H�$2��Ǻ�7#�Q�`�[y���9�7� 1ֳ&��c�B�3��%����Ș-"�ҝ���߬�9������P�/��\0R��1NG75���O;�l[��xT<&i��v����CI�!��E��sq�����fX�U;fe�{#r!��/9��ފjׁ2��j:�Ǝ.�%�1�f��׮'(CA�9�B8��!ϲD�)%b�I2�r:��^�\sv ����	9��X����ɮ�w��crw�z�;��,�3�Qn��*#h�r��b�P!�s�v���O�\et�QQ�!�-lM��*(����5lRȘ�S���`[��t�.�� ��{�{G �$��nd�5���ɂ�|�2V�˱����iQ5qm���ĜUd��i�)����O�.v/@q�^�@ز��Z�H�.�3/�I��6�Y�O�{]�f3�:�p�l�Q�(�O�q�*����2���Z�hFD�֪ �	��v�"yD���h�i2�㏩��GS��& ��B�$�|E6KLi�^�K(f&���7��đ��ZF/���	���QQ��Oy.�ۓ�������7lQHQl6����]l0?��sqn�}�`L�dG�����p][F m��<�a-��?�C'ʆ�0
O�D�(����o7�J`Fp!�Y��
@��\m\�׋|�J����/f&�PUb�$�m���L�����a�����c�C�v�
�\��m	&�(	��v)�{ *��DN�d.���E��'�#�4okX�C�9��Qls���i�_O'�����/-gf�x�o>������q�AQ����N�	(H���~Ϻ2��*m� �v`�+�XLs�����QJ�[���g� \n3
�t}�7Y�yN\�M���,��8=�i��h��Z�5�a!�W� 8ܾw��4'�0k�sQ�2��d��R9R�lM���i���r.G'���Q�BV��b�%
�~i���o��:D���1˃��\�G�$Ii% |��]t"Mj5��)WW�8�c���QCz�F񕽻�L�vB�8���-�4��Z�pt/o ��EO{�;�B�F�N�����e�����VIn��(�S����'�o�=7�[e݋�"	�I�b�wlK��Y�	��1�!�<g�|�~[+��N��io�
�*z�(�i�OB$�r����g��7T�o(Rn �hL�\Z@}U+u✍@c�j_��.&Zg��{B�\� ��,wh!��JKDc�ǈA��[��`���#�m�I��#���8po�(�(l�R�7��
�\�3K�ML>Sq�;"'��3����v܌�Ĕ��l��=�Y���|�B��d��X�y�P��V�1s���E�M_��@�Tt��K�x����Mɔ�� �m��|�Sx��z%Q��a�SC}�Xww�&�$vvg�����{�b�$��Lݭ�s������N��%U�/��E��j'>r��v\�9�J��{�\�a�Ee��+�T�1�R�[���*�3xԗ�!�=�E'�/T��r��>r�fy*Ԟ���}��I��-Ċ#JH\Q�aP�q�����(����MR���pB�R��Fq��'��W��ç�!�Qx�n��/h�,݌S�O�8��`�,n�j��wk�#3�&�5m
`PӘ�՚;^�"��^U��P:7ې���0��ɗe��A��O��m In�|�K���+���x���+���EɧɓAeo��h��&���"}:�20x��e�b�B�9`� Er�2ླྀ�$5jv�ٺ�Ǡf6m-��U�g��vm����2��8��J?��G� �յ���fo}Hơ'n�����܀��ӺG������?�Uu6ga)����'5��b�($����N]Ԧp�G�0�����B.GV/�����EU��E�Q�] h�Y��7�T�~���qOp�V������f���Z�ɸ�7SS|܃��x��v���l���q��r>�.=�&O1�-2�+3gk��%6��P�J#>m]\�g�������WZ�fhy�2p���a"��1���d(&P�����Hk�8"���;7SH��lg+'vG��ϵ"oj�g$�D��~�x�U�!w��LX��y4�`���ai�� i����ZwX[P����Y��L�M$RA�G�PK�񆮜��%� �O��zN��jW���������ſ5���P�} ��a���H��V��B[6���T7�^T	9~(`:�GB�8���Fa����d��E�ø��6�7	5P�s#�PoyQ8�9Moх�xBa�t��ʑ?�`*����_z�]�F�{%�CtƵP�������@��~͕	9�ܖ+6K�ɪK`�����k���X��Tg��=����\.��9o���L��A^bwP!H:=Q�ڃ��K��B&p{��,���&R�I�a�e'G:c��@���%��s���@X�����|��K�`J®o�+�eI�)X��$<��2Ku�܈P�Y+����BZ��%\�!L��N���Q�m*B�8�K)Ŵu������t��L��VS��^r�+�σ^eBp�Q�&�B�'�)��^�����zV������F�L�J������ %G)���d'�~�g�)�U���..���s�q���5��b�8h�qKJJq��wLP�W~���:���u�gCLߔL2 O�1��p.�.i',����	@�\P��4p��_1`�~�AO�4��)�u���q�%�"-�w���;T5��}'�{s}��1��u���c���~x����'�B =8D�-��l���К=�l�5��
tsw����_qc��	2��HU�J��Ƣ�}��g&Y�)ތ���bHB�S����Ы��ƒ���J�p̧4��.��2�����0��ʷ����V�ҏƘȾ��p��X�ȍ����W���P7y�G��˃`�7x3�4�� e(m��/�V�md��ӺFP�c�� x�{Z�J}�J�f"M
���ck
�s�$�j
�e���;��Pa���b��]&�D���f�؇�b��õO��!�t\ܐgr�'��$�,D8�:��傢nU^PҦ����i�f��3u���;Ͼ�%��T9Ɵ,����sJ�L�"�NvLʥ�X(�%�AM��"c��si�(�-�y	��_��e��q���h��
 qҺO_�j�G���Q
��7��8��f���[.��+�F%5�D�2B�un� b�.xɔ���\��9��6�Li!�C���6^��ѡ�32M�A��A��C8}�5R���w�y�g�� ��]��D�ymO�4!VSՑ��!�|C�x'��K���B �B�O��� p�`+��!��~��P����w5��ԥ�������t�ř��S�`���.%E�9A�ϓ��u�n����)>wBm
ET��s��d��1o��������V7���}ڪP�f^w�{$k:�OY�:ľU��=j^4�Mix��m氟�j_E`V�tR�}�P�9+(��)�	�4"���B�[�<��1Gi�B�\�:����4#�1e�eW�tW	K��z��:��<c�x� [^iޔO���j<9O�LI�@#\٧�Ѫ{���k:��S���e�Er�ɺ�p�NY��r����Ԃb�٤b�|���+zt�N��vM� ���Ah�����fT�"���Rt�;��m�P�S-�Kx�i{���P��h9��UlM9� �F�H[g�h����G���0r�nI R��%1YH���]"����!�ħ"+���}��!���5�������[�e*nd�S�}�~���AW�|���d�*ixYt-q�C�f�ݷh��ĉBgXt�t�3� ��}��2��������>�l!' N����|RBi.@��|�jQK"b�o��R��ɲ�D�2Bq�`�G8j��M� 0A�*�6�\���A�!=i�����*$c�a������ `Hx��杍{���32�?ʛ�Mu�X�����>��� ���)�J}��j̳ hu����M������%>k�u�]��U!5���/�9��	S����ұ��w��l���V���Jf���h	�uu�8�������M1W�#S����s?���0�U�7�7�47
)Y+k�w����t���R���%'��=4tK����؎s
{���R҆��{|��@'{����X�0�Db��p�v0��V��վ��s5�u5o��>x�EK�h�~B�StH]���U5hV���jt�J��L�pYMu*�T�	S��`c����O��t�q𑫊�Q��i�������s��F�d/�����Vz=R��-�/�ɓ�^�9��k�������h�q���@zij����nD�.j�p���2+^�5KI2B��4�B���X�)*�eM,(�K��	����VPD� �c)�-��eg�PH���e��p50�a� Ry X��o��@I�)��8g̻�9v�����CM�kCr�|	�TE��\�yc&�~�2l�����d�ReO�	�!�g+��V�����g�Ss�ڜx��-�ʆ���>=����뜖H��l?!gD�T1�Bb���Zh=��kB�%��=�N~�=������~��ÎL+�j��yC	���L�y�{e�*"C��w��!7o7-!��u"�ᢔ4�:<�`�68!G��[�uɾ����#���e�phjy8t����J������7�A5�������';�kſ�rd&'��dG���:D�گoP�I��a���_:P�d{�F�\Tt��|����!X��M
d��&�tE6��]T`l�,PMd"�G��l����T��ҁ�uG��
��KV7�>�lFP:+G~^�wVG�U��?]����U����e��	d��nOL�Qשs��8u@�R ��W�9���ۇȌj#�@xpP��������
n�r�c�ƨ�P�A'<Qlqvo�V>S�]{f��z���J�=�L�5��N���MD��N	j� ����!����w5�S��Ј�9NDN�[kؐ�z�c(5/�*6�/��p�@gbVO}o�}�����2�Le�m�%X�AD"��+BP��i��$��E޳l����B�z�`��Y����*z/F__�l|��Q2��ޱ��� ��~.qy��&:���\m���kG�i�9[w��D�Q�/ܬ����LT�"��A�N���z�,�b��
m�J��?saL�ܫ�Vz�Nv()�7��Dsڳ�h<��6�S%���u{�2��`����(b�Z�/}��1h���A�$�KJ����0��d�P��r�ˌ��RV�T՚��"3���|��u�7���=�"%/�=��L(;5��]�]5D��2��ܧ���݃�����i�Ѡu/�-SR�f�����-1>��3����@�f�]�65����k� P�*	��}���=����y�+�α�);x�?�yt�ǖ@���0���a/����>	l���R�n�7?9)I�*���$�~G:$��F]�)'ZTog��Q:?� �qqQ\�1��L�f=8B�Dؿ��E��������cx$���Fa��]��W�Hۺ�-���Ŵ�fw8"��܉���_�:�g�DK�4��Ɉ,;E,�tN[��_���>��\��>�L5=l^�:�f���6�"VǱ6ff�H(|�-�I~�9^��p�VRC'^/'S���G=F�N���!���W1<iًĳQݏ�Ly		���Mk^y�
a��gzE
���dZ|�&>�4���O����/�X�I��Ɯ��VW,�ͽ|�YJւ刑g'��j�(�T����r�'�_�^�?����4��h\閮�Ͽ���QbE���D��`�Z��?!�*d����l��c�@ ���[�B�і2������M�0�gI!�9��Q��	�KU�ꐤ�Ll����j�4��g�	Tk~���0�&T�HO�1�MLBvz���jJK�ar���P�zj�u�U�����X�T@-�ԉ�n��(�o"=�-���E�;���!*(ɂ�/@�R�b�.;SLt-�R���M���{�+�6:����_�qA١p�ka����C��Zs郲��G|�Z�kܛ��5�ֳx�)Q����@�ϧp�r��#vv���f���h|�)���/�qP���W��5�אT]�U�|h=x\�c
������V��i�c��
���6	�=�3 �NênM���<蓝�q;��Mk�T�٪�����q�F�E�����-�؄I�����4���컠�h�P��fjq�re���Z�a��9Ƴ��@���[죔g��a�K�ދ�²���[�,b==��!R�����=2R�AԳx.�/¼����R����1"���)�Z���vâ��(�d�m@:��|_��󤊱I: ޤ��)솕R�5u�����'�hȫ�g���u��o�p�WM�5���Ӎ�h�+����<��MO�]ڨ��B�RN���v�8]@�eK+�y:�lf%vc-{����>v��<�p��@�+��S�!5G�Ӷ�oY5&�U�Ň���T�� i"c�z8Th$�g	]m�G�T}��D?+���T�א����nQD!�ĩr���9�S'x�ж�##XO=S�,e���.ڍ��X"t�X[,��� �F�(ho~H8�������Õ,j�j�C�蠴h�Z&��gi�"�҃��+�v3la���C�7FT���ji2��y��4�g)T��y^Uc$�xh��\.W��u���A|[/��Rb����c�ߍ_�����z��3�'�LS%�(ղ#9��q�̳����l��\�C`�O4�(�E��-N(�V�2�X��&ht���,�Ii�b�� �p�-�6���u��XH;Y��X�7��ybT7Hy$���	��m��Wс�Zܳ䓙iYu���R��K��B7�������� ���M#��5 ;�7�eY�������#�Ł]���U�b��
��%�W�q�fE��X������2E�Z�zy���� ljyh�Q��v�޵Y��r�71:����nv�B!6Hat��ܸ; �uѫ�_j\��e�W���0SH(cg��ߩ�����D+��6��i�S�߶Q����,tc��t�Џ�����J#�&w��)����]e̓�)���yAֱ��	���8�;��=�B<Y�6e��S��=��<�I߰�*~#h�魇9�![�HX����o�(�lf��	EN�����̫��	��Kl�=��:��v\��x�*C��9̲�����-���G�ƪvf��!]���̊ڧܖ�wRz?�t�L�iga�D�r���ÍCg!D7�oy�!G�lK�m9ʄ�t����Q5->���u��0.)޵��a逫E���qZEgP��"
;]Ǧ�W_�bY��_L��yTC;C�\R�C� " �\��C�( �T��D���9�C�&%����d��9�㮀,�lC?�E@U	]g�%���8�5�	�`b�7Y�)9�"K3��2��>Hk~���BH��3���D�C����j��<��^�x��v@pT��$պn��zmN�F���ۀ�K׆�U����_� �D-���������t�����1^7�hf�;ݯ�j
+��ѥ1|���x��T�nh78�a���(�;�qՑCƿ(�K^~� 1���6� ��L�E�Ǯ»d�/����0t�/e����T��:L8�0�J{�V�W�LP��O.=(vo.��c�&�!^m��R�B6�>=��/��/�8����:{e���a�f~l�����W��>o�D/��.$&U���2��.Y��4�/u��|P�|7]�!g�-kH�y��92빃��SK.���L�	�T�=�qꙄ"��+���ħ
'�����ĎY�k2X���IC�<����'�d�9�ߟ��`A�c�'6��v�$n�v�r�c��:����Q����pc5���/,P=��ߨ@:��cڳtL��U����"���2��z��A���w�sX��g�F���i����=��҇�]5�N"GD����¯e��!{��ڶ����H����CH�7iN�ј%�$->S���n=��U��HQ:�ӻ@��J�ĵ�:zn:�/��g�h�3P���r8���T��$�K�\�?�^N�p�XÙg}��^�vM+�9���Y�ВR��;�Eq�����Ѷ���2��4�K�c�Dɡ��ԴԱ� g��\�-/��˞�B�$�)՚=�����a�8�%6�)��h��t��T�5x���)槡G�G�Q�S ����־ә�CΝm[/�Y��da�2%Шj�X.��%�P��] �wF��l3H �����Z���>�z�&�R�}Hy�g_��I�����5?on]��$��=�;q�b�F���B�`D�v���|j�����+�%n��\C�>�ۆ��g�����#t0�]��\W&#p���آ.�}_.t��a�X�߂o�_��@:�YbԐ8�E��bB��wkQe��^����aE�`Ma=�W�!oc�6��g�C L�:�"t��u���|'N3YN�{Wje&����BaJ�x��#�Z~{���V]jX��J��X?[d��~A%����H.�� ����ϕ���l�_p��:���!¦�1�� -V G)���?��:V	(^�x�9FN�s7ϼ�5{zll�dk����V��9D�ܽx{6V\B�Uq{������'��T��KI�NH�~�$���%	78��W~�:/�����׾nNze������L>�K�}u� ���rg8�!���2x&�m�9o5�SИ[��]��v�#��(L��U��t��\�f-24_��KBm�Z��_*�L���Izq��x�,2<u,M���C�p@�>�m��}V���r.;O�6BJfm��(��R��2�h�p��дZgn�3����
�S��v6D#�Ô����2��XI*����_�m�C�����"iHi��H?u,w-`>�IR���j��u��[-���K8gź��w���s�~~.�����<�`�(�c�!RYa�G��-i˿Wy��'��g��c׆i.Fa�딠)Ŷ7�=�.G4����P����\!^��3��r�G@�\ ����x�����p���E�z�n~�O���HN_��YR����VKrBN�����V6��h���8���&���8�Χj�Aբ�������)�����$Gq�8J˺>}�����n5N��|ٗ����2��4й��ɯ�5W5r�4��8�~�����C$�)��)a�l�|K�aOē���������K�\�W��Bm TiquD�ɤ�˅�����S;���f+�|Nb3��C,=Q��b;k'Ųq���va��gi؃�@�T��u�χ�+k�j\7b�wt���NF0nȀ�|��tc�N���о�'6g��Ku:��䄼b�Y84!���g�s�%+�����K��~z�^^�}���ƣr�Q���8�F7��л	��T��� K��ݲkVN;+i�4Q�V�#����(#�Q��� {;(/[�ǳ�����,W�b8�0�J�9��I#�|�ف$������P�4tS�A�9uF(K⑪���҈�*�Ԋ����{ocTb_�
��R[m�9���$�j�3����	��o�s�jT��w��4H�^8���!�@�j��K���~p#^퀡��m���'m��e<�LϾ���I'X6�(�#�&��d���3��ʀm?q[��]6�:��GB;���X��g�U4b*G��fg���b�-G{K\����ݾ��w�Hlg_�j����ͳ�-z0�O �*<s%�#X;���qu뵀���x��!i#��ͽ:��I4�5D�S��1n��nE���,G�A5&B�J�OM�6�ӎL��į�[���+u0�h�Ķش��_e5|q���|�^dN�#Ϩ�Z{�uta;��b`2C*��\�������%��S�����iBL����zbj���~:�)���~v`m��`�����<�
�I�ꑑ!^ɬ4R��L�5�</�8���Z�3	9�����Ҷ�a�ǰ�:��.� &9{mU�MH��/uHϾ���&���}J7r��-j7�?��Bö���9b�i�*̍؃���^#��_9`x�A��GoF,F���|��#-l�FC���,�6�j^u8����F�@Z�W�!��Z�:d�Qn)@,��&�}A��W�����E��>�h�"U0C���=0��G=|@"�$�+2����ݰ,���*O(d�w�֦^L�\��ݱ=���~�N�6A5�g������8�������;���p�D�"W9�~��RRVemV���sW��}g�6�Il�y2��L4�����ɋ!�HP�F}��CL�0�	#�JP��?ƼJ�rVfO�:��d��p�h,0�����@��S��:�6[����3�27>A\�tC�p'#����p�t�l�G�G,'^@��`I�Í�ND���A�A���r辏΍�f���'��g�Y�i�W7M#���;0�]�p�RK��QG�PI��K)�g��K��)���brz�iX^fٔY�
���S��t�W��%\�|����I{�qJ���?�
��H�`Q;�&s

���(O&D�<�)�ʓYZ�d�X�����<Y��a���/��gk�BD/���h�&�Υx�>ס�g_�U��E�K.(T��T�ΐ��h�U1}F��q��k���O�u_�t��ǔ�L>DJ��y��V�X*�ԦX@�e��x���\�|������?M��*NI˭@sPtH��(��?bM$޽���~��m��/f���P���Z@\�Uh;f�f��r;P�=��M�A�-��qa�DOa��Kt�Ý���@B1CX�Z��-������M��#MJ�N������_��ܱ���ݯ-^�ڎ�Y�B�4ߤ}���|���(�W�N�	�z�KX�~nV�8#P�t���-�X�[�`��,E�YM��=3%l�@2�̧T޽p�3�r��RK��gl�iו6��b��
w�S�=2q׋b%�>�@w�tE��֖6�
�:�_���[q��gf���y��T�����Z$�I@2~����~��]�6�X>�����74'�B�D�U�c�����^���L��f���@��������ٮ<@��3��Vf�F(&�ӹ*v�� $LZ�o�zG�A��G)<�qࡂ���7��3Y]�(Pd�!T��6:u�,u��>o�9���^��b�^���3�@��D�r��C��W��&�-cѹ�b��L�C೛��n�� ;�z00�4`·V@8��߅x�<	]���r鐯Ys~���מ�
� dd���!E'�/�U��X��zi��Z�B�B�M!�T�509ks>�5��8X�6�<ytm ��>/��hTH��a9==W#����Z�93�7�'8�u�p3��,
w�������	[��t�i
^��	0�'jM��g�����lò|d��	׌Nk�*�01�'0H��^���RtZ��7�`S8�T�$���(��׬�"å����6��Yq2������ێ�S=���H��k��c��I`G!�^��[��D �/�ٻ������+a"�7"��������~��5QL(,X�f��r.b�@�:o|�D�2��d�`$��H��O�{��P�7gW�G)#�G����g-"���f6��izR3��'���r��Vak�f�ߐ�v�F�B=uF�;��2�:`ӡ
�YG/��Ai��-W��2��3e+�q��I�(`���g~�vI	�Ubc��9��'\o�
L'+Q3�`�#��(�<&k���;g�J�ϒ��P4j�^�u�P;5?���o0�V����%U9�4�I[&
U�Oq��\���q���8��ʜ`/��bJ+��	bo������Wa_wV��]�B��t�`��>�2s#��sO^qCH�c|�7����3�y�OBC��\ R�!]a�i'�P�L��mC��U"��h␜�|��gkX���ކ�yV$4��5VR_`��Vk���I藢�:�c'cT���g��c��5��4���Q>��|e'�+��n�p����A�L�իW i.��A����F(��+釛tE�5r�\��� �%�<KF#�=�c�;�T���FG�Zh�~���8��J�fiP�	�p�㢃ߕ�-��Ւ� �b�/D_[nr���i�V�;���џ�ؠ���׽^�:k-JO"�C8��\va#� F�x��zr�#�;����<w�X2�.=��8w��J"N�����i�m��D��%�c$�Е h��0�Ը�a�2b�\r���D��,��^�WEu�w���2<��jRً��0�?�B���
oO{�	d��l��t��5=}pH����9���`�J�#���7�._�����b.����ND��)�� ;����m$��h�dE/�f��"/�וE��(ևH9���������KL0vۿ�ݤ���T��=�#Jk��v�J8/������s�h���[�!܏���*{"|?��a	�Q��3�j�6��#[�1��|I���Edy3��'���K:���=P!B	I�������oJ~��@���X!�,�ޒ�:z��^�C�f�,���b�!E$/|��c�+Ι�g���$W6*�s��Nua���^q�s�g4�B�����G�}�+�3��������T����F7�����4�A�V�i�c#�R���S�٦�8���a��%} L�D���#:�*���&��;�&��o8�D<��b��/{V�=���Ä��@��%��|w�KF��$߃��|O����M*���de%�
Zx~�t�[5F�0��94.ڢrE�@L�rm*{�Q�9���$�[4M�����p�mf/������T[��N�`�Q9�Gqd�iz(��<6-P���1��������cK����f�/)��<����+��)�9�nq���s9���]���^H�G�J�C�(aP�U�eH�е_o����ң��F\�h�`ެ9:1��dW��c���8��R�	�EyJ��h�r4o��\���C/�:�K�^��r�A �!�!�Lȗ��{*\��ovH��,��Bu%�BŊ��V��e+m�&�[���ۓ!M����:���>(�o�5����S'M���-���{�>�W���&�:�dtxlD}CF�cL�"ZWk��
r�9�ѱ|`�ݩ�9��1�=�/'��l�Q���Ta����ܥʒo�!�t�.���y�.��i��Y5��C�P��y�Un�K��=��ӂn�@.^x��?,r5W*�ρ[����h�vm��qmٱn+5!6���;��w�q ��W�s6��ua���>��B�\��yn/	�|DʯHz�Tf���W1�=�lvL�e��M�|�MH5�r�6ZF��3��<��Ll�f�\#��e�yyҝ�5�A����}�]Շ�һ�I��7���	q]���+�L�LU��<P�P��ÆӝM����WKts�/#��mr�U���n�M`�Tж��RZ��ҜJ��י���<W�I޾��g>zщ�R�����	�w�B7�[��G�	��2ݕQ�G�I��P���F*�A�|�'9��Pd2���6�Z!���D���u�TLz���F/�_2`��| �|v��! �'�IL!8϶�2s�}ɢ��j}��a�;�3��J�Y!�^�?2���Z2C� �e�_^��'��+|��������#X�0i�*:1�M\��WX��5�&Bq�%{ߍ��"��>����Ŋo�b*櫹^h�'��1�&a��.Vcg���DZzI�e��ѻ8�a���mc3{���U086ߛ��ۂ	1'��l]g@j�"����?�1J湐|�>�<�Z����Ҹ�~h�c�S@R>��k�o��4?�k�/b��&���7Q�t'��٪�9uq�/��(#VձO�)̸��>|
IϗjfE�8;ʋ	��NG�n����=���BӅU3	np�'�ѐ%c"L�Ya�@��wRH�bs�����7��R3��v�=֜�4��wtm�i����ჼKx�>4q�&5�Q;��W��!X�gƹB?������2d_Uu2%H�HB:ġ"��U*�Z.2�*�����$GMhz;�T��&����6x(��S����^N��jr��&���)�cϻ�޶�{1k�����t ���/)�b�~o������8�n�2�
&6�0�6AE�Ɋ�1il4�`V�@;�R=}���[�[����M5С��[�ޏ�#��><�J���i�9fq�n$�B�
���_�+�7Ia�%�1��(Uh?�J"�����1�s��#�_|(�v7e5����f��Vt�̲��v7x5^u����������+܁�+�n�G�V��)1m�N����F������t�����jx�7���MB�,�M;i�h���Õ��!���-eu�����!��)�1��w�$�� 9ю��~Mnr�ڇѤ9k/}.������:b�n(v��?B̊e�,~�.Ư���Kg=�����2�fHH�O�5�g�#��ؑ��*x�R�K�X��8�����"�B���VV�r%[X�Bz��� �X�����J��y��1�*(�MJ�����5Ծ�������^�<�mؓ��Z�rY����,+�;V�,��ٟ��V�#/�[L<������
���hjj�UA6��(��GFD�*���v\���͛��[\�{����N=b��|�;�pb��/P�^s����olg��4��-Jυ���d�o�.��$��@G
5Et��~WqQD�0�,}!��5��Y���[�B�N4��?�X���[*NҮ��Q�Bʥ8�O��S]$;�ԠGȿV�¾�5��K!��JV�z�\��5�c�]S�ҧ�Pyih��wv'�8�=�<��`_�J�����P���p��2v�Xr���.�In�(��iH��*���������H&ػO �3�q��#�4 �����ゝڬA��w�	�Dp���	��C��э�B�-�����%�3!*�X�W�s�kE���S���p���T��.D4�=�#�Om�]��kr�xߟ���&ap��rN��6��[<�{�|�OY��!�98���(d4�G�K�In�ѹ���8�v�)8��F6]��ۭtiO��\?%�!�6̉�q���0�!f�Q���L�:�ˇ횦L~M% <a � {�������&���dq����������ݢ��9���,���@��x^�K
��=r5��(�Z	ð��?��}ʒd�F��#5$\/"��������h�H����ǣu
C6���!��-K�ݒ�h�� \~uԣ���f{ɺTD{K�X��d�3����o��yN��]d=��x.����� �/��k��m��C1=�eKK�Á��b!�c��\���Z��ғt�e�7r$�JG3�my8��}��Ƽ'5��
b�:&�Zd"���;�:�U�D��`�CQ�f�c]�2�gj9�׭�An�
�dh�ʞ�n9�%kyь
�L9�Y���@��XV�sV 2��$��̩�,�2���csϣz?����-*�~<+S?C���N��$x}�/��ÛXFv��^��i�f��'3�_�8�*��N��&`5/c��6�+~S�6�9���?����-Y��ɒ��!��x���?�Y"Q���O�[Ǐ\���	�Â�i?�ŷ�1'����X�q?wwxѳoS���vx��&G� �ZZ>�y1$�LYM
�5��q�>�z�hR߯_��_�J��fk�`��q��֨��q�KrN¯o�>8��/��%�|��ҙ\}���\��� l�nv�JrA ��lD��/l� �pE�';�XM�;����#��MV�(��7_'W��WV��a�o^G\��Fk?|ړ2~@<q]4>O�R_As��ɋ� �}/�:ea��/=�ƷU3&k�9z�����"H��v�eQ��n
���aZf�\��)K���%��/�=.�P��ah��o�=�K�Ň��Ӏr��ҹ�2%�#/gU�.�� � nm�MKO���V�Q/`�� ����`���*U�>NW�I���\����I����N4Pr�4	�1s���*�G�nJyϴF5�gz��BI-.^��{����-����U�ޭ�C�8c�;��_����B�U$]�}yƚ�-�	K���&�(��~������fl��VF�rQ��pvI$qWKuh�b��X��<�rA)��+�O�;.d���XqH�Q|�X@�H6����>Lc$�����&��A⛿tq�_�d<��؊���$�
�}��� ��%P�<a'�4�J�5� ��g���2V9n�~H�d�'�x4���)�8ͥ���px����ߚa��c�K�6�:��j�2 �sT�0����U��U/�����Ղ��6G����X�*�`L�c&|-,��˙rT���J{�QC6"�]VP<�5�[KY�0�U�[LuByH�[�%̸�0�y(��c��.�y3n�f�EL�z�J�/��6m+*�sCgn�� ]�`�� ���%E߹V�+���c�O����G�!�2$72�%��>�<G��Ҫ���Z�/Br�u����7+B�}�MG~p��,,�P�^}5>�u�Ϧ��a�'�!ކ:����d���A���"E�:N~ b�5\���HT`�DA'7(�2B=
�<��|M�g�'��	�ĵN�,�˾��z?�F�)є �l�u�1��q���z�曂�? �B�>�a�\��&��7��w������wϑ�?@��_�,���E|8vG���z�8[6W$�]��ǹ$ZD.���0���Y���0��{$n�US,k�]���L��2.:�҆�m��A����sgQ�P�2����o�K,�G������p	ר��8o�����z�U������:�7��W't���9s5�Q )�p�lb�!O��<`��*������+�0�.C�I��b �D^椘�ZY[�pY)��E��D�Z&���ܧ�F�����|�5ċ1W�&�D�#u�����Iv/���!����L�$S1٫^�N��T-/����?-�:,�a��OW�
=TM7��V[c2Eq�ZFvs��
�Q7zj���/��1��/LN9R��T�XL��XO�ﱇ,�q��q_�JD��G��+���N���g���]_���"
i/�b��C(z��t�׈z�NU�o ����߸W��0�{A(5Inxp捡�f�m�	E-�q+��� ��j�l��Zɡt��-�Ct�^z�%��p�7�A�,�RB�> a��L� S�kO��&QaI<�r�Ps��
�����@�o��+$��rj'T�㱅�����+�m��b*y�A�V��$�̻P
�X��ɗV� ��Fu�	�:�u�,]�ϑ���^⊉�]�x��],m�A�DY��{S��UJ��$a)	7���k>�n4y�M���'�a��"Q�I MU �S�{lb�~e� �AӜșD���%�ɶI�iN�?Eyli79�펃1�藾oy`j���[�7޲����z�B�r���ei����9�@�ġv�tUU�Z�<|:�d��V�k�O���l���S�#�N^;D��kZ�- T���<X �>�Vz���R�U*��{m��N�0���u��b>��>��E�PE�N�f�t�<7fi֘�Q��tX��)��7�S�������@��;*�vT��|���-4�G]����}�?�wk����l�<��s_oJ,?Y-Q7\2�����\)�u�W�>܌��RkMI���0\���~�:,�ju����X.z����1������8�� @{�&i\��7�����a��0�t���1���ĤH��_ղ���i�Z������b�e��>R(���WU�xԈ��w�-�|Jat
��Z9�����1�_ߌ˶0p9��Y0�^	�Pz��|�)��i��W�㓪��.X�R��ce½H������}
hȘ��`M
����*������f�3��r�l�cd��c��:L���;3�\l����ԓ^[ӠM+/. �U!e�w�upX���$yEIфs���Ђ�xI�7�#(�Hލґ.��͸#lNU1��縦��rTV��[>u(z�MS��S�\��ϩ�e�0��Z�F\(��bhE��
�q8��R?l��V���L���.�nf�{�U�ߥ�C��Z h���NU,0,��,0��z�o���2�S@���8N��T���m�v�IoS:�=�w��&���:��O�l�䓐${b��[��=��&;B���E��5��$�d�r<E����O�&�1�q`���(j�d]�8��	��Ҳ�II>����kJX=����teä�)��p ��!t�-U�(�#�t���*��}\Ѥ[L'�����?��$�a�0ڳi���#M�!���U�+T��sn�ړ
,"���������T�A�L@�����i��>�ao	�O$�:�Hq&CR�(oy����O65�>�5�
SJMj�a�6^m{1�4O!>�1�m�ۍM�)r�?��L���7[�;�J����h�,�7v 1�T��nQ�Ntd�,���DCc;�D�� �d��Y.xw�t�|nY�%�w�ȯd +w]�OLN���+g�|�T�4��ۘ�F� �/M}��N�Y�4�~��$�}�������m���]�4#�t���$��p��^�,�x^t�AA#�h���d������e4]�?}dCjH����U�'Z����L����6�S��	�Kٽ�͋Z�`3V�8"v�"V�UύKP{ `�7�e[ƹ��8���Ć��
����w'��J�d�m�T$���D7#�;�0���C���,�`a&�jʰ��\����`@DK-6��հ��EdoN�!�f+k�u���^DT�A�`1�cĞ=y���s�]��!p4j�w���Z.,�'�����,Z2{V嗧x1��T��+,�Ԛ�飥}uii�g�b�g��>F������Wd�Tl|��'X���(�UK��P)�Ap�X�'>
�]4�fƿ~��s"�1y&�D�I�F(��h[cGuׇ��i�I5��"_�r��N9��R%��Z^�� ��u������d8&���*|:#����"�Z�x�26��Ғƴ��x�?�+` }��A�(h��{&w�C�/gE�?���g�"=�V�rX���o0�j/��Z�\��������k*"��C��}t}h���h\��)l3��}į`��7�K1��&P���ꑇ��A�:����m�6���0����w������e�њg�XRˠ���	M'��O�H�j�5�|%��A;�pn�(��7�R���ݗ�A���#��@��i���6�uܾ�)ϋxJ\O��<9��ᖽ���I��m�M!Hx��D{�`� kPn}<V^ >�^����,���D��V�g��NRj������ܔ��S3�	�[�3Rl�k�O�
�"�e����3BU���Ȼ���-l�b��`�µ���:x�t8���H�˭}'�4�d��)��D/�m��暏8�����ޔ7:�����Hw�x���J�l�BX�G��+� .��m���=2���s�?���YX��"+b=�'�vE�����)'��������B@M��5z	�]�|������kd�X�Ȇ����*ɮZ��ݵ�.��U,*4������d��9n���ُ�lZ��4����^&ߩ��W&r,}x�����azd�x�}�xovY� �ς�YB)��j������P-)|?4?� �yk�V��c��C��2v9�]�z]r��\^��j(v��nҒ��<�9�����pW�|�S<{�w�)��\�;i�Lz�3|�_$�lO��Q�t��Q�(�oM}�qQs�|s�D:�Uκ���Z3���S=෶�Y�<R�F�?N�v9�����0_�����S�8D`'�Z�~#�YI9y"�����ke������|���f��ɫY`�â]�:��?VK�,��1�0JM]nr�s ���������w� ���M ")`Ƞ����v�47ѹAp���Xi��}�Y"��Y�(u��;��ks�}��AN&m��N�lb��N�vS-��=5?'��N	�)h��_:�1坆 ��[aN�HX��ru2��o�`Ba��.v"�xl3��tܘt��v��$�F��+ɧf�����ds��e���UM�m��� �u]�td�"��Sd�^�1�TW0�|�u�z��3*�ܗ�H�܈u�<̧�Y��åYWp#R�]���H��yO�gr�TB_�C�T�>���m�Fr��ԁ��R�mZ< ����� !iqj�)�j5�{��轲%ܰ���6�j�ꌃ�����{a��-٪?�ؒ�`��~f�J�0(-aɞS��P�G��3��xlr�}QA����_�NҞ�;�1�aTt����~�sPC#a^$�Pj�����D��G��� ��z�]c(sC����c<'���A?�#$���6����ǲi�ϡ�����&�E��*y1ba��K��!g��k �Q��W�9�<�\G'�?Ӥ��8QL����� �rY���'���c�#��&�=��}d��%�d^�z]t����G���:�
2�Y�d����;�#ԗ�!`�i&�Xg�	���ꑾ�l�:�Mr�~�"���qAV9���ui�l���+V-�L˥�?�Pt,,=��~\��0�=X����R���J��;H����V㇍bW�� �-���)M��'�u�'��:�4\�s:M[R��/�՛4�X1WaROb�J�AZ���9���1�"�%���qS������8�7��I36�QBY:� �hB$?���,��B$��%��Osj�c��&���C��9�1Ց�j�#G7���Y�qUA��A�8���@��Vـ�G����рr�aN���v��+��Cx
T�~��%��pm!�_��ؤJlm��aM����ca뱋��.���0Яi_����:���L 'qJ�!p�}��z%.v����΂ �b
&��9�+d`�>&jt�hK-�(&vl3�`��{K�N���P�"�ԩ���9�2a��^�&�9
���#sIQ�XP����)�)�TO4)�J������-�!�?��"��{g����m<�
�2�����p<��@�<J2G'_8��L�H���7��6�����F���],���%s�g����w0�B
[���g�'�B�f
7��-�!�w���7��`8��ӏHr�qP�2l�.L:u�������n��JiK��e�eY�@�2�*|]����ί��Ԯ�0��9>�ӡ 玬5l�#����D>��3��YN��=MÃpˎ����g����溥����L�7S}��>Q|�E���s��*�&�j:^�.�^	gb�Cl��S��Q��W�V�V�z�⌲h�7)��K*��9�Mm!!z�Ԇ��{�E3U\����j����Q!r�q_(4m�D�MXg�{{ʑGAxf�
[�m�_�B]���1�~!?h����7H̀��U��ކ?�Lu��',�2���M�w2ayi}8nUAq[x܈)�ݤ��9�s�t�-�)��m���;��i�
��8@��O���f2a�`��3�3�#V�l����@'9���N�%f�03�_6�I��{x�xg��`A�_ȗ)_EQ�a�8�8w�p�����4��~��LJ��E
�W�n"5�{��U�ajc�o!:��7�����_ ��R�u��)}�����ȕ���B����f��.��ķ}d�/�M��g���'3S��W�V��y�"�^~�͋Hi'R
	a�+�ï��{�b�C��?n�dgx�*Z�in��jG�4�E��H�ߢ���8CL��P�ܓ��t�V;x�x���t�P��� L�&�^�,!�|����Py�k=�3��~L���rbd�2��E7�%U�S�4�a�|��罠�ʎ�z���d��&�3^���b�b|��9t��Շ�-�N�L��L���s1�����DG(Sb+���� �V���V�Q�Rԉ^��Ϸ+xG�0J�r�Kj���*2h�5"va�hg T�����E��V�&I�PƂ�S-��h�|�~R.\ﭽ܇y�#��6j��u@RT�ixn�8R�{	:�)LIsӬ�[�ZͫnD<��D�x�}�S��2�Dtih���l�|�+���7wZcr���S&����m�K��'������{��.��ځ���?�]\8Ցϖ�TaXV��}�� ��C�Aj��"�P�N>b�f�&j��	��?|��`���~4C5���	bj��"2�x�I6 �/X2���zI\�����ʾ�������OB�tn>�����G�6������w�0��j��Q��EW��)��?B�ю]�i&������R���@�����!cRO;p�z��W���(�-oD��Y����h�2ߋ-H���!�F�sH��c����|q����k�D��ӊDg"7��abX/���KOD?���X4�^�ί���Ĵ�q�d�$3�Lp!��ֆ��`�ध�
%�ړ������.�|۸�P���e� _a�ev#Jf��po�/������aF�B�������z�p�%��`d�է�E��úU�a�g7I4�8�%�(8�)^��_�D�:���J���#i�E�wE1����7F����7�M�I12:�m���Tc���z���`�.𔯯���PH�[�|!{��Bq�����E�]h�]�p]6�{9bK\}�����W�o+�� x�w�m	����y�9|hΛrX��Je]3��
�>#0�����a�@0NK8ɔ�5�r������������������(t������*hz��d���r�/���w�tnHr��T��@�ȴ��i�X�I`<_k����q�O��~<�,\��h�Eާ�y ߸����pF�b��Sk�N�<���F�U�z'q
d�%�}�t~\�y<�g�i�~1�xof2�C�C��}���0��Y`
eb��� K{f�ѨB&��5�!&A��������wl���PZ��g⦹+��@t�^�7.�;�$ɸ5x�
��Z���?#�{ҽ��A�u�h-�G"�O��.�!�{��7	��^�V:pZ
�O~N^-�_?]'�/�"W�ٙ_u!?�w��+�\[��_Jgcd���6(IGA��ɚjD��Z�h�!����Ng����P�LJ���w��������I�<�5蝻��`����n�p�����Se��
��t(���X~�:U'1���O��v��<}x�ug��ﴄ�>F�\W1���p�G���s����g?� �,J���{�t�7�)o�¥@�US'��M�}����nˋ
���Y_|dAc�1��Ei�%�0Łd<R��D!UP��aЕ���Z�AJ�r���T@T��@���2v���%���5�͹v8�z� ��o���˸��L�t�7�����<�`��H���{ba�rƂV�r���oi���D�i=v��v�f��B��t��+�.�]��̣�
��І�(��1���#��)�0˖���8Z̚��F�5[�{�*J%�k�D�x�i> ��!4>d� 	_c,���Q�:��뜣���j�0�+�cv ����.|�a�z���w|���)ĵ���v�n��'��i&j7%pt/�9w�Er�Ѭ5�+�͠��xZ��/}ڷ��?T��}I]m��Y<��$oR-�Mw���ǀ�Z{�o�N���}|v��XW�
�[���D����A���̖����i�ɿ���p?��-tI&���J��x����\[����u�
�Ϫ�ݼ嗵���c8�K�S�4:��N��O�& g��í���"D<甡Rz�z�d'Q"���Ɉ��|h��.C��<{&jG�竻�����󂽶i�Eȣ��*�Į܌���£p=Z��L��n�Hv�\$���m���i�BN�����]��<�"($���~�l,�Q���0g��X3�	�ܰ/�~�T<�ϖ�ޛ����{1/�N)�����~2�����ʃw��p��[T,�ʁ�:�E�a����`�eB4<��{vx�c��+>s�G7u��_�A�v�w\�p���&�~ēlaC�,B3Ɯ�S�͕�9�!��Dz�1p����;����Oh�2����+����J6i�_��n��$���N�8O�G�ZT�H��3�/�3��IgV�
����X�p*��m���57��x�l5pW�L�2Q�+���s���s�m��"��K��9��E�jه+>R����n��J������bR��'�ȕ�����3^�jҥz����������>Y�Ťj#��	JޒKB{�ڬ)t�:��qђ&jQļ��H�l5�ha�W�)_�a�v�_#����O�nA����߃\�<d�t�l��C 2��咪�w�y�B3SnؘPQ!���זR�Ħ7���?�~��b�l<�s���A����&�d��5�^j��h\m��)���������zQ�޾I�]�,�]7�<.wЭ�1��A>�'�b4��Ȍ���4� \:��}��g�����P���$7�`G�6�Ov$�����
&��U�zi?�?)%�
����] h��ɷ�i$if`1V�$9�{���8J[�J ��8Yq):�
�hn���\O����Ј��^�b�2�cK��.1pjU�Y����IX���Qk=���d�<�0�M��ɸ��"m�����K�fFB�b�/4�s��#����,_��. M�n[���ʰQ;z��L��ȁ��he��׶JwpR���9R�=��6��}0и=�\G� s��X��4��c��%_��i�����U2����~OUމ޾Wbl��$	=������y�γ�����1� �R�}���0"�|��s����9��/)Sq���t���;��AI���A�%jSY#��`������g(���Н*�ynΕ��c���F�v<}���8��(����t/��Τ�����qQ�߰��1�����o�J�� �}^�Xn�/��2ծPu"����Wy5+h}<�|3�n�8yw5���y���X�d�CTd����7�\�D[��=^��|̛M��ab���1���_��"$L��p�7t��	
9��&G�i��j�q���Y��R�����1�7�{��/]�Cޕ����qɇͩ$ӭ���'KZ���G�oXѻ@���5z鞤hL��6���>-1�e�.0W �zOGU�[�@��0����s�o�B����}���˦M�gX��ߓ��BmUrQ g�Z���6~��o��q]�MM �f�����tk:ƘU}D9/IP���[�?�_��w2�"�!QG���&���E�71�%]��.�J�u�k��\�E��װ��uV���
�5��n���ĕ��A�X�v2�g���n�B9r�a���V��|{�9�Z�0�"�ns��j����62y��GF$�K�E-R������ͦ.N�T>�b�U �"��!1��H�=xΆ9�u<��}~���/]�W9>Q$���8�H�F�]�a'H�YL�KQ 7>�{�<Q�x�Ω'n1�g�J���+u"_�F�d�b�^����)��[wh6��������ыsJM~����HO�P�r9�uZ��̙��0Μ�9Y�>�GN����5�B��ʱ��m�]�N��O�q��mT��V���~>[g��[��KvWT�X5[L2��[�4�0�n_ϭ��~alj��5��V��@�0�c�J�H��*T�P�7 9t��{��/���P�Vß^�.�}^	x]b/�!8N�0�|�M�]3�ffi}U��'/�.x����#�~��/9�C�X��W} vE.>%��&[�5-�K¸x�%%2Շ�9�p?Z��<9?�KW'����,T\��bM����T���Qt'G����$�Ŀ:�9�����������	t3@�s�����i[Nqv�V��#
a�c�q���[5�hu��La�W�
�xC�,����4�(A�@��pI\�"��}.��{_Cp+����0�	��@R\ ��	�~&\�9B��k���6Jy�e���ܬB�;R��vzU��֓�fq�3�b����0��c�:�{��X����fT0�XB$Gȣ��Ks\D�~�!�x��)xa���s)�V��!7��C���Ro��Q��"t׭6����[T����M��S��,!�`P1�ɇ�}-�|��{VH+�{�a�NЄRtp�@�J�UE)m�yk�ղBC�Q��c6�~�?T�E���~�j�o9��c�-�oԓ�6.�
��v�B�vg+��]�/���u��x�zO��/����*��n��\�ىO����m5E��ƧIE�.d�O8x$�߄��Љ�n�f�����a�����D�0$2��(�_D�3˷��>�uHqE�9[�*�\��G�m�G����Q1�J] ���S�d�_e��P��%�J>wt��H�5��~J!�%���˝0=k�>_��l�e}o�+�t�0�������E��������l�eP��9�S<-��T-�U����9�j";a����!dpxZ�c�BDj�fF|�ប���.'�G��!S�g�T�9"�-EA�B���]�?Mf5�u.�;ĴP�29�*��c�0��$�d.k�hX�Jk��T�	!p ��E����|=���Kvf�p*�k�a�/<6�ɒ����r;�Oy���d�#x��^���1?�qQx8�ٌ�I�ˍz紩��k�0������~�Ӆ[Q-��_��ᜇ�B��ܑD��K�b���>Rz�b���;�{�X��x�Ŋ���Ēi���#�����
�΀J�2?��ao�ڐt)8�N�� ��aR��ս�=����WOV�����BO�Q�u�J�/ՃD��b0��[�|x@%i��<�n��	���T�C��W�r�X�����ne�/�j�Khi���*�(�]�I؆�#@���+p4�x���=v|!x�Tq���y/�ᦗ���W�°�Q�T�ȿ2 �D"�a^�-S�f����o�V�N�|��IN�X��b�^~ ��~�;>e0d�>�D��C� �QT�]/$9wA�6��!��b�����`��!2�W=�{x�:�A�8B���q�Ĕ\߳��=�Q%ƽ:Zd�Z��h��L� aŭ�M����$�lhQ	� �������*@E0@�f�l�˵���ʀy��ҷ��TO���ٮ���=�R���[��1*d��HfV��)��착��ȩv0�+�nbУ�J4��+�1F6'E�_3�Ua�D��k�i�/��1ƥ���}T� S�x��%�,�zx/jz2#�"�Y��)��Z�7�j.[�u�@�*����e4S�"%�6���V�>�W������h���'�6�wXP���"|{V��ٓ�r��6_&�d�?%X�x	͝�B��d�[_A��D��'��ÄL��(Đ�p��q�?�z��++����?9+WX�^��X�Fi�w�m�y~ȃ���+�o�ⴺ���Z�l�W�bl������N����Z�]����CYȁM�p-Z�XhZ}m����6^�D�M���������F��gH�Y\�!ߒ�s#�d ���ջ�jҵ�x�.�7a�|��l��w��~.�' PJ�ȸܒ�H��pz�K����שy]LE�ˈ����,��6;]^�� 0�k�;�|D�ϱ��O����� ��,��ڌ������{��+$t��U��{�w�"����ϛ���>?q��*���@fh�L��x�F"&v���:[&����g��̢U���^��@�px&��qgh@~�M�G�1�+���������� �F��?�U
2��Cu�]-hU
�<�Wϡ;r��b�<������>���.�MG��F�*S(��^:�B� }&��ߧa�=6�Tؕv���p�ם�0�����~�Y��cEί��d_�/Ū�����1���pv��抷��<��H"�W��7�	�<���5�"��@�RP��o��e�i߉�g���;i�u�֟�= t�w\)#V��1i��[�m�(8X�Խ���-#Mt57�y��d
���295�ԅ4��>��o���Zuo,̸��y
/u1�h�N|���\Z��Bו�mB�N�fK�� pbp�0q�kpVM�dx�j$�υ�(�!xR,�5��4M�@�;
�<_���)@���j���H��8x|Wy����"C���WS��dH\<R.aWx�>�	z�26��mM瘪p3��_�cz��?]��3�Ayaճ7��w��@X�^��AeGDih-��mu�Tb�!�ٗ�MpUX�Rq+;��#Bt�v���0wtv�&��^����i>�4��9����$�F�(��{D)C1Y�?�~�,]�	�3N�j*��0�}U�=�`٤=�����D�;�����W�L$9D	+C&<�jqG�|̅6������HP���)���cwm�%}$���=40M �]��2&��ى?l]���M�j��\�I\�umI�6_I����CS�¦m�0�wV�:5@(�j�I��M����(��	�s�5X���r�W�v�ֽ�e�
N��>�]. '4N�+ڣrA�k����4f���{������اӜ�  �D#���I@�K��	�	���lђ˾$��{���T�'�T��\FC�6͋� �=ڌ{���϶��W)��8������8�|��e�{0a[���EӰ�G����:dLgʋ�[
v�.?&Gxd3� -�;f�0�}��4Xk��>R{���ކl�)tl�V;���A���#�J��{��"@��a26�����v�);~e�A�T��B{�%1JhŦiC��!��mf��}�kSTweD��P �A�Ҽ�Y[Y6FW�j�_�086�I�?>�U��v��[���gP�WKk�OE�J�Æq_�WW�r����9�"�Q���O��p�ۚ���~-���+G$��E�e?��1+W�����bJ�RǪ���TA*���W�y�F�Ib��F�g'�eO�����N��N[��8S�yp���'+�]< V���o΅�}�J� K~�Z�E�/&����"QOk����΍�.���m����q�u���]�H6}?5�c}�����@�pӫ�B�6�ۇ���VJ`����/��m~���R�7�/�DٛNM\�e�F�q�t� �>��^���VC�܈��D��;,H�n�cƼ����[��>�2���4R�qBU��h9n���9������& ��������e \��+�P5'�Lbc��oʴ���I0�n0ҮR��xb� �>���=
�:Dn�Z���v����.�.���)\Ӻ�h��·$7eu�m��?$^
�� m(,�X[�vVRbM���>�5���q#9n�8q�H�גC�_�q��!o����犚��1G��&!�s��)��	l	�����*��ǌ�,�_r�d�|	��a|�?��8�ʣ݁�18�A���ۃ��1�gX
�]�J�）#��,�nۖ��b5A�J��=��V��1���NT���7�lz�Z=gՑ�������)��Ht*it��l����Z|��"E	=?�{!��.ۛ�hlҞ�iţsw�)��1��RBh9��I���g��|�
�*��4��3�����-��}{8f��s�_롶p�*���3a����bdgO�v�v�]�͑+���'��c���R��w'+kZ�;VrZ7��oe���Ρ�f$�,����'�B$�l�ڡV=��A�W�{�𑮈��'=��������b��`b�(��/ /'��*.��'t��}�-���Z}��_�`��� C鈊}|��$��&?*#4l��0����wyy������	��Q�1�&��Ig�K���q�XTA�y�2��a�|�t�w�<��,��X2Y[�N՗[/�b;���H�/:D0�U��0��h���:e~�q���3��R��F�.s����O�sLeF^�D3�O�̛F5t��'Jcư>�#���'``�ÖJ>���?���9�TV�o9�d],ԏkT.�GwP-9��.ҠSf|�G<��:�[Ž��R��EG@5i�8CAջk�3<������~��
��2������3�_����pEVT�@j��u�*�(1J6O����35Â�	G���b��U#�Z�\�Z�!�{�na�k�n�wߞ�]�J����3xr��4������-V�����#����?��x��e?�k�a�U��S:�R��*�]�W1��z�l<N_P:��	�"��H�>�?q�1!^0>�8ʊ�؜�hLA�C|P��"�e�=��u�#�+��e�����"l]؅��f�����o2�fӡ�DJ����C�)�fIf;�~������_7le��[P\]zX�?�Z>��fBc�-�"����y�H��h�iIn��:���>�m�����*���������v@7��_?�P�3�f]Sl�=C��|=�1:�-�{�[��lY���Y�ʋ:�?���1^4L? �_?yIT�������jw'��ϖ)�T+y��pFI�yB᫊ɘ�s�
�H,Ǵ"%P�[ ��� X�e��e�s:�8���+�V�b��8{�Z�W��t�ؓ���%{ѷ���bͫ�wId������kؐ�}'ˉ��UQH���V���/�H�v�L�d.後�zp�&`����7Mai3��Y��<fq���`+fDz�盲<DAG��p������1����d��f6X���r���53l�{/�r ,
`���E�W�ޛ�6�Wj��9��kU��E����6�ӎ��Y�!�W����[�. S	�}���y�x{0]�¢�{���ȁJm$��iA��|�:��1�;��ʓRq��|�([kt9�4c����k?� �vm���a� �1{��>D��6~N���贋 ��c�����b$�䏤]E2��K4L�-�(^%�B]CL3�M�iͼ���"�7�;M	N��]�B�]�)�Q��5�X�Ay@>U`�5؍ ZX%]Pe��H|+C6�ڜ����O+`ܵ�����%�%S�}VM�Ǚ�juǖcBC��c�+����B�9�弗w�z��g�Y��S���+6��2�;L���A����_�5U{��Q?Ƕ�7��$�EH�Q)D�Zyox����k� ����P¯�)�!�As���?`�H��+��Ͼ �c������w�/�j�`7n.�p^{��q�Y�Ojd������{�:\�C��YxA]!ɱ�'�I�B�s�Յ��z��� a"��B/VaZw�0_��'�o�)��)�o�&�0�����-�#2qAM4ƶF
qg�y��o<��`�Ò��*���+8g(Ä��Ew�ϊ�(N�B2�°�?3��RY�6�cj�j�NQ��e<:�I���O��?&PP�p���ǲ����J�^���3���8�T�E+N�,n�`|c�&�o찭&�����TO�!V(e��F�R�)��z&�td���e�����i�S���i��� ���,F��I=�	��������u1��ى�'���U=m�y��
�	���d�f���(Y�F�W�K�&�<DOޔk������ N&/��R�N�Ѹq�[�k�l!K��9��?b��~|��{�w������mjS0!)o����wiI$G�������1l�y�k�}w� ]���������
���~�l9z�/P��]��W�ci�Η�c3��JN�{g3ɚ!���eGya������s�eG�I�}�2���z�.�o�����gpCH��?�n����=�w��*���&c��]r2����=�⿵��Bgúz�In����3�*+>��eoOw��g�П����p���G��2�3�ml~��bz��/|I� �u���.���+0�3z(��a�j�6���Eb�x\F�G#y�[4�|��Mu�w�����O��Jt��{�q��'�3�K�rǑoH�_�F,"�)�f}]U�G�?|�Ÿ:�H��\hj��;w�f9�Q��}�/o��,Mtϊ �
����p~�ҹ/]p�
�ȠC��gC>���������[C���ۄ�з4����9nΩ�<6+�_����I�:�>ޣA1����X^{�Xh��R� ���d������Á�R	k��$�(�K�j�|YU'Z�0:QguzЋA�DΊǂ�v���νis7�vJ��q�a�Zd.���n�����N1�7�+�W1�,S(m>
� �����^�{��?Y˫�6,�/s��-�Q8���1,d�i��W�V#k����?�1�Y�.Y� �<Z���.w��u�R�	�2��k���A�*{�}8��4��;��8��Z�+-E�a6����p�&��, �k��?���y�:��>����sM�����;�t/����a5���ox�Z?���s��Cq���3<}��T�B�H�{z�8P�IYJ�g���z`4�v�o�J��Q}�8�w5��N O�f��NU)����8�B!�/�5�����Q��yw�M�Y�5㰶T��Fh��̽c��'�\i٧�;2���5%`�8<<�z$R4�����]cv��(�ֳ���?ڀ^F:�>�NW��g ���O'��ļ���N�V�n��;�.�{�G�YL�}��#_Pm@c;����Z�**��
u�1
I�v�C�C9w��*Fc��0�������s���S[��]N�U�&O%�e�u^������/��B��%�)�R,uzFp2�4{�A��/*#�����>��9S�U�r��Zm�����i�j���M�Bքp�{�P�<r*��PJΏ��!t4�:̱�U;(]�Dt�"%b�|S��=�]������^���F�_u��"�}���@G��8�Fe�i>}�i�mn�_X��~�����`Nm�c��RȢ�����dϿ6�!>C�S�	�g�k��L^{)��X�vа�C��T���uQ1�u���	���<�,A^:�g���̀F;�u~��v�@����T~�����6�H�%��t]�č�[7&��p_oѮ��ej$�(�9�1��Z���K�ǴE�g��r ��3�E!�D�Bb�"�t8��,]�o�0�P碨c"�r3��%5O�T ��.��/�-cg�n�m��(��C�\[�vV�DM��f�M�����3B�.E�������%��k�p���R�����I��ky눷�
E�5pq�	ɨ��/��a��E+m�
������2l�s)ew����Ǡ�b
UB.������]q"�N�+���>���P](as)�Xu�N�����b�����ێ�:l/F�M���lF�&�nDO#�a	�����s�y;NKV��M�Nb|�����f��]i��=p�袄� ��'��ds�E���}ʛ�&��;��D��S�WI4e�F���]�!}T��n����I���:'#/$ޚj�l�α�Er�0�2���al2,9��=�g�����+�C���t�Ϩ6%�X����������Ԇ��Ğԕ1οO��ɫgŭ��E�5�4�?�93��Lv��}�J�dP���5J5�}/s�q5�7]U�k����hwXn꠭�����q�Y��-��K�q��!rȅ�P,Q���c*N;��f7�FC�b$LY��/��"�w��޳IA�
wUy�7���t$%Fe}� �m1'gI�&�&-Ӛ�H����\	�z$^��!D�%) �8�����e�s�l��j�r�ێO�"�@��R����U�N���]s��tL0�����'��˶���n�թ�b��.�Z�oaL���W~d�5<�^��� N(ʹ�q�zn��Kn���_P)޳�����w��2���ڟ��t'��Gs$����t�@	�G���0������!��yapw�m��ܠ��~���6��L�L�ga����\�� ���PV�5�����RUp��1�������x??��Cxe8ͪ�� M��Er��XF*���6ޤ	$��'*��ͣ�͹�uI�B�gul�<-9hs(}Zoo�&rT�}�[�?����U��a���hd��%�w���7�7��Q�d�0��y�Ѕ��n̵���w�����OwXVG����΂����^D2�4L��? TH�GF~x�)�I`�:���gu�ão�$�ۯ:1��n�w<Q 7���"�;��̭Īo�w@O����ȫ�B)|Hq��:˝�5���V7I����
8���m�X!Ǉ#�-���V���zp�r�u�
&�d����g�d�Ɵ^�o=7��.Hx����l:�������q�؉2B5�;qM~81�ĭؐ?VgX��������~Rdc/P� ̋��BW5(�>�*�ɘQ6Oj�H`�=�+�`�@e�/���2B�۽�<�x+\�c--Ȍɧ��:���(G�$Luzu�d�A�d�&y�").��.Qc� �f �e��@��G4�>�)U�q �Śj��x���݂$
-����N��LkGR����k����lc�jK�S���W
���mnn>{dRb:�#i���}jk���	h$h����L=m7�R|��A;;��T����(��f�Rx�d& uN.ܺ ĕ��TeW���nۆwK�T0G)k/�?9F���Y#EᓬjĜ8�[�8��gB	{_��;:(&��a$x�¨����w�=�$w�c����#o�M�2��I�o�}�%OE݈���W�#�w~�fC�ˬF�.b��q>:C��5�*��$�6�^թ�[��t�+#�X-�/����U�ҳ���1���̋O^��0�П�P�D��L�����J�S�(	kJN��e7�1��J ��3�0�$�i�W�R��ȴ��\�h6�Tp˦j����CY�� �]��9��"���Fϓv�rQ�GJ^�܁G�i�$,܄`L}ۡ�cwȳ&���W-�L��H��O�/�|@i�K��e�Ke�����zsph��kF!�<��}p�U���b׾=��H�K�v���3Tnt>~;г��r�����Z�-��o����J��@�� ��`d8֫�-�4��j�B�8�ù��ͬ��~���X%����90�+ V"Sf��(�	i�j�m/��&Jĸ:�.� ��QV����E���&��.��m�$���}�o͕���S�U��5�����N�~UB���\^d�8�}S4��K{���ٮ�[���S�\���鋫���AX5u~I�3gI��Č�o>��t��D�dZ��
S�Bq�h�F���4L����9���P$����!��K~sj�_;RR��a]���<n����/Voo�	�Ӗ��w�Z|�{�Ġc��U���0��Ѵ_� 4�`�9� ���z��Ht��<������U�C�O�m�>�J��xV+�l&�+/N\�
���*$�ڎ<�R�*@�T��²x�5=	H)ڂ>vje_g$�>���wƊ�W��>M��C����ӊJ�	���755�yA���A֒1eO�+�&Ui��љK�<�8_��,S6+�r�z+)h�S��&�1�����n)�W�=�HQ	���\*5�.�ϟ�������'V���� ���Z����y�f�a���PR�a�J;�;�+��s��r��>��f,d$i�*k�Ҿ������>�2!}W��
�L�#��y��&�2h�](͕gqz�4�l!�яqs�˫aC%��?V�Ο1ƙ�hh����x�=�
��J�!.@4��Q&ƭM�'�$?���L�T�d. Y�M�-�ވ3@�tCB�d� Q�di\��'�[[n���*����U%o̠�^�����Brǁ������P#�W��A�횃s��E���}Y2{�!�W����Y��*�{'��Nİ�����$-�¾�X���~K�%n7�'(������|�"*K��o�	���Z��u��?�> �Ͼh
�Ҵ����l��� 9ۮ�n�;}���I�Ev �IH�}*��-�4�r(����T�U��s�pO���ЇS��������U��ʭݟ��u�C�_$��b�\�IWiĄ�w?�ֱ��c?�W$��~^v54�̩rO���:�w��;���w"�����]Y4)3�&L�N��@&p}�X�;��!��Es�;w���qTZ��!8�Z�@��Jm �8�/6x��N���V|�Wg��8��/���a&�"���-D�����R�5{��&& ��B0�ƿ�J�df ���5/4@9r������M���|E�KoW���"��ʢ �G�OZJ��U 1�9�!絊Q�9�����9q��]'��hZ]=Z��RO=�}�:�fQv	�GiQ��JY���!���P�k7�{�����u:u������*���pǷ���!�S����EC�S.����+�������jjsK��4�]H,�lʒ8vO:<'N&y��B��� �H@[�r���"�YG3���<-�m���b�	�M����5������,����B���ç��t^�cr�W*��$�:�_/�-�7+�.ׇ9����ݮ�AZ�.�$5��J����D޾Q)���a�b��w���Y4��2̒��:����s������5�ސ�^�� ��;~�Ʈ��w2�*-�6kD�XT��d�(����.�LG[��T�/��ЯnN�@+�������gy$:Ԩ�c����f8�a%�Kh��I�f ؁��4��ڨ��.�zy�aM;�w��m�N]�>|�o��4"K .m�l���:�?�{Έ3��`NFړ+�D���pǀ�DiT"��ێ΀�8Ǥ6�m4f ���d+c�Pduu���T��]�mx�~�ə�1u"�?��pC�v2@��ѭ�㸺�w4�K�kGBH��V���Ƿ���ht<^|�wy-~Sv�f<Y�%p�Y˒���׳��ah����V~��DEE�F���m���b� 
h�D	ޡ�bGr��8�;�� H�kL��Bי��8�T�!�~�9����ˏ�B\~�b�y8��'o�f���-�
\[��_S`Dnc��}�:U㡟��1�h��F��n	")�@�Oo��AQ��H]�Xs�5L�P���J�EUc�8쎢���!����&�#���==�)@�Y�N�*�U���Q��R�b�K���T���8�vˈ֤���������vf4>����������m�)Y[Tf�^��Ȃ�j�i�n��j:�+�M����p��Oe��c�1)�W���d��tv�w����T��{�ua��`��As��¥dJ�M�WR	5�6~(�i@�}�x4��ס@=j'��pGzy��+�r�������fM�'q�ڝ���\�mS��^��V?���f���2�z7Aw��N���t�6h/�v���l#{p������Eɚ\g���<G�8��z�qw*�:g]YtDI4J�![�3�~"���jՂ|�)��y�^}e?u�I�#�Iŭ�n�y�'�T��	g�v��~dO���u;Re)>%�N�V)��
:�U��K���^�_��*��n�?ۊ₇���/F`�#��W��g=��3`��?�`~(���uB�mǪ������<��05�M!���֣9nQ�,&�k]m#O�V�h�a����� E���G�,e�$ׄK�w��JI�Jeg����7����l��e�Ts�2uC�jȟ�0�d���o�L�t��6Lŀo�AOyd_��Ȓ�dw��5�_g&N��ߔ��M �2�$TȤ���L����H�(p.��"p;�����Ŏ��J�n[3��2�mK����u0꓊sZU���=՛d�l��?��R؇G��j�@N�Ӏt��V�-�W��V-V���w�`<�C��5l͙z�<�_�F��V�ӜX�y�Q���/f����e�8�ƚLa��Չ����C�bR���6�L��f�u[;��6_ =R��ͱ]��=z=2�#3:�0HL�/1�M!�BEgeP���5l�~��N��=ٮa��(�P­�?>��u����R߰���������8,���n�H&���6�SD9��j�!�e�jÈ���:ʩ�/:{�V$k�Ns��g�#��)�F�������T4�<��rP�2F	Fi�M�1����q����k,�6�[��^L$�!8
���
"v�?�j�H�|.�ك�\) �G�i��C^�)�g�9+��-��^�$�E��E�{\?}F���*�_���t)7�i�Mr,.�g�� �
������jYiR����3�8#7J:�f��]"���������Z�)���]����4OҽgMOQ��?��c�<C�|ƛEX�˚j ��H2>�T����e�Q�Y�E��]��=���-G��Ơ_R�Q�)'	:|��b 
���H�BИ	[e1*���N�+T����i�&xhK-�\ZQ�k��q�p��5e�| �K4�ax�c|�Qmz�W���J^�SW�A�V�DO#�S�<6ڑ�z�`�}fM[�f
𐁾!��r y�;���[�����ഝ*L��#�%������#� ��%�tG�*p����<��CP��du-YO۳�l�C��؋U���ZEo�@���/2��P`��?c�E�ʑs��9o9�@��?�����aG�^:z�!o�#�X�)]���7���s�jv:K�������5z�ٺ�����N�i~p��s�Om=Z�y�1�S�Ԕ�r�,�O��ڲ�u>�|A�!����f��^��?�}���p���H�i�b$��1�D��0�@>���9��+wغM�@l�y7�F�BZ�KS������&�Ryϻ x�U�/�҉������{�m9Q®+sG�
$��ǀ�nz�m�FLR�d4�-~!��=�?��^<����ƱK�w�k�%�p�������ӧԚ����"ǔ<p�|��-�.{���g��_'?��:�SF���<,�HXQ���t�����#��eC���8L����&�	>X��5 ��s�6�����џ�kz�m�~Oy�J����ޝ*�����$�,����`�
�J�����'y�&}a�*mn��S���6x�w�HZ6N�$3���0v?�?�#�'����F�G=� ��Ƅ+r�|Wڟ�>gK��)c��[rG�>�h��&��Qt�U��Mܾ�6�Hm���9�g�WY����5���]��d���zu\ᑸ��F�����gL��Е�&��y��7�v���ќ����N��kpz���~������ۿ�7�n3F���>����l�(�ʡg�R�`$X��n-��щO�-�T$��s�4@g5/3�Mr{{�7�6���k���mKI9)��D���0T��urIԣd\�/R��n'�������*;]�$���e0���j�~-��V���ɺ���mk޿�u����rg�_Nd�C���f�L�$�c���h���c6�KW�ش�pP���c�~tˏ�<2��:�lW��|�ٰ�I�pc��Z���������L96���;'0��G��G��0h����'�Rޑ�
�T�����Bo1��X�"x5�M_�A��Q���a�Җd������ϧ�����_}N�Y�l�E�Ͼ� ��g��_�&�2�~\�� �"k�7!�H����z�jx�g(�I��5R�F���/t�߆G�J��%#Wi��*j�W���,� �8'�6��MQO�Ƀ�������W��m��2��fc��r��%��hm�|��?2Eᆤ����p���G�S���Uc�N/ �L'ڼj���3�2��la�S	Q��D�N��a
L�=_n9�٬7�㥚h�-���������rX~!����,7,�@^�t�r���R�4����|�)g�����k���v��}�th ��K���-.П��m�S�!bY��sH���0o7>�� #d9v>2��p�Hm}��xBѣΡ�	�%�%=�8_B:��ΔQW�M�\6^�`��q&:�H<Ӟ�݄V�N�w�3��r��'B��w����b�mSe��rRPԯ8���
Uء����b��/�b�4ɖ�$�&�kC�:؇�6��(*o���5Zcp����wivZ�4�uSm�sg�]�.�;&��rV���Iһ5P=%�K�n���3��ay����D��÷ߨ����酎�4�]�(	������+���\�.o��TW�׋!���I�����4�O�_�}�O�V�PP��M��1��M��lM�4� �x�S�#��ƭo�ɾ?	�E\t�0gn~ES��u�
H6Bs�p���o<Cq[�W��K�*��@�]������v��7���ӛ���rqB3__�`�OSb�f;��l R���`YX�zO&���yya�%#]�Ql��[?�2-�"1��%����G^W�4ĉ0P@���{���,��0��.cb8����v�	�=;0��E�����b�a��� �N�ݵ�gΟ�rf#�]�r�g c������#8������Kk���C�Fy�?&I<3��U�b�'���+��Ք;�4BUa�u�E�˃q�3�z��4a�:�X��8��9Wn�Ԛ(Z�� ;���
XF%i]�9�a�%o�g�B*WED���)f#J�'ك��wG�ᳲ��J�ٸ��9_*�CO[�`F���A8�f��
��07�o�0��u���O'��f����(M����o �\~�l�V�㼂3 ^	dG�F�l(~�"�&-bI.I�	Զ��W��ś :P��\����	��h­`x[�v�s�.�r��&3p���dP��|��O2�i�y��JȊt�.f�s�vJż^0ձ��j���r��a��\��5�Z��Y���u'4vT2$��F>��S�Х������I��;B�ާ���_燸I�M��<ߍ�!��;R��Qn`��%�"�d	m	h�����k�VH����lo��������M� ��*3-őB�[���5�n).�����Y����Io-u����<ڜg�O�e��EAs��ŵ�d�Gn}5Lq@�E�1�ǜ^okj<�M?�#�F[�G��?����S��Z� �,C��e����ƴjϐ}>�c�T^�YbUd��n����u<�3�>"��Д"�n�$���/o�Z3(���O8��}�b�3St\����n�ۄ�l�ж�|����T)�n��F	r?i��dSp�D,���]X����*�{��^����]��l�-����v�@���)y�^��������l�� ./":T��9�4OA�6��K�����z[/ R�$:�;ǩ��9G��D��o{��HgY^�� �&���`SV���>̒�HA��C.PL��$X
8��������(ܾ	�v����d����%�6����:���	���!���|��6*��u>�șk>�\0����2H�6}�-��Q�B�#�5Bt~t�xg������FN�MTU�c���Au������L�G
���7�(��p�$������F�Ukgs�$�=���N��[C9)L�ī�M��>to����_eG��H�A���GȭSBH#:8�@(T-���o��������V��@����?�/BF^nr�'�MJ��7/����<�sz��`�D4�ajD�H�8��C'�͛P@8Xbn��y��ZϘ2�M�Na7�(�K�6q�Ω�4�� �_ݖLAȳ��ߠ⯵�"����n8(���!��+$z4��Gب�k��S�mJ�eWPP�QF>��FD��Ro�9��������<�%���?3��pUu��ʨ�H�r^����4.�ă����Bwa���5�Փ4���%ڋ\�PG�,��u�<�81�Zs�ɾ&���D����[܄��o�_�-�o/���U�1c{��g�ઉ�w������g�S��`>	JuDȖ�k��W۵TI�����[5���R?c�k��q���� 0����-'7S#Z���F1:�{�ۧ�F�bzzn�+T�6�)_�(E����RË��u�gW�),�5�닣�W��#���	s���M�x�0 P��X��	/�M;�ύN^�� ?�f�WcM2D9����t�P"��]o�ڔs�P����hPw���y>)�u�k	 ��;<ƹ��� ]���z���7���@c�f��^f�U�¤�ދ�U�#	�	Q#�X�w2l��T�|Pt���c����ć�4�38���p�����5���C�C���
.��ܯ��K��L����,f_�:2�RQ�?)�/��w�l��0I��h���l'��i���f�x�\Bhs�]�ϼu���Q^"wV�tB^��FR�U�A+������S$��+P���gM�Ì4b���賯X���j�N�o�.�bDhITr�-r;�)�8w�>��E��n�.¼r���$}
#a�1����T�&E�ՙ+���v����'/ii��dyKѐ� /oݑ���m�k8m