��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+�������;�bM�o��q��-�ВM�XU�/ q�8��up��ޕ����f:#��Ÿ�QBBf�6�dm�	\�~
fp�3q@�V��e�e�v���u?���H�p�褣��
��?�j�S�X�$X_����UߓPU�'C�l�ر���8i6#5n�鋮&����xO���m� ���?�y.��"ɒʠW��LL��ѐ�<�����V��:�xՓJ��=��J���� Ԋ��@>g���0:�q�C�/m�)�:Wr�-J&v����t͒�}q���G[���ÚU�;�0:_��5v�h��4q��b/�:M8�����˳y�V3\-�o�3�p�S�opm~�s��~�����&��*v�z��?H���@�{�g���Ӯ�)=WN���N�M_�?p9��*��IQgWF�
��7�Gw��.LX8�2��=~�=�����o�ȏ�Mt���Nħ��rߚ���7>��?@&��ˣy0�C:]�J�2�_�F�Q,����[�^h�� 15�@����̴�ܘ]7�M��%S:�U���j���T���K�3�$Mݨ�z<'-�����܈�}
l�~_���10b4����}'7�.Nz�xxn�1E�����5���g�����"Tƚ�7yP#��cCjC�dtd�4�<5L�v�$ƕm�S%�����p��θc|� ��U�~V/�@҆'ω'�G������g
��0�u�a���>��9�����@
�X ���Эa��s]$�t�=�E�--ܬ��l�9����p�;�Ouʇx�!Hf�Z0�����[�������BǄ���\�c�v)�j7���y����a�r^��(,��L���4�W�g�oG�P�D��'5���T�����l�M"���!W>2��~3A�Q��7֮��:�*y��wo)�ؐ��g�ȉȑS�I��6���U�9ݹ���T�� 1S�0���Q4�G�?�P��t����ȧ�	6�.A�؆e^�o΋�XV�yS� �R��P
�B�+�A7��}��pW�^K�C|�,��?���{����������t3�����\u������N�V���%�����M��c=�^�����,c�-+�B��Q�<�G;��&�`�LWN��������z��NR���ُÈ�Xv%���-��۶�
@s��@��5k���Yv~�=��`�P�c,�Fo����)/����`Cu
H7A4�T��i���4jՁ"�)� �EU�^�Tj��G�#��<��<���M���e';S��$���;'&n���d{C�%�KNQ�wfOB�Up�$\+�g2���KץY#0�	�pˉ��0-=���bpm���U91�r�`7W�
�ϕ|�B��WV#�q;ŀ�E-��Nw�$w�؂w� )i�oSw�X����_��Ӟ�}����,��
����*�bb����`j�K�<�Wj�=��K����)>g2�Iv�G�@2p�֖�G��|M����J?�q���i ���yl�h��n��R4�e��}���k蒡�ï��G�4�U3��g=;�lj3�e�J�q�{�@��\�o�;��9
r϶�����A�9-I����~�u�C���lp��b�P�z�٣�5��`o:�)�f��'�4P�#/�O�'/����^(ד����.t�_���p���],�-���A]�^�ᰫ�e·3n|~��k�a����.�^K�.!1Z�o�$�,g4&���_q�?2 �Y�.+��y��.F+�|�ě�44p�g��P4�%�&8��3�AB :�06⮷!�w���o�ڈ_,�	�߃M��o��Jd��j4�j�P�
b[���r��p9�=�hiS�*:���(�&)�8��=���m��T�"���q�F=lF�Q)��o5s��QJG���*?'�g]��1���X�!�=Vk(��3[ ��#�5��`���.|E�jJBu1p ��$F�y|��R��p-YgL����^�4Rb���8,�G<׵�0��O���ެ�"^�џ�(I�<�M犀6g� ��j�D��b {DC�nӼ䮵��Zw���{�l(����4�c�P�7�eL(���(�zz�84�?�c�k��Y��ա5Q�����FTT����3��xa0j݀gby�}� _q��A����}@	|>wZMA������'���L��2�V�e'�y�!|>�^i���=���*�[](:HH�K�R���H_��C���UḀ�
��:�!��$��޶�P��M�+�i���x������.�:�@!��1��_�
`D�P$YӋ�=K���̑�9���l�!UT�#��k�)�C�����T8�������{�v�$��� �M�Ԙ���{n2�yj��{mJ:�����y�nN�j3���[ⰼa��"\��%w?�S�,��b�y�!�2�akꉇ�dT-V�b��t�����q%�����d_�cӂ�/�C�Կ�1�)��Q�\f���Fn���io�X�f��q���+��;~��j�0p"p��I8����*»VY��-�psh5/�G�M�m�W�*��",�ѩǐ���wh�hh��ﵗ�m� Ӽ(g}����FH�= ����ZK��˃77c���z��f��v*�a��pѢ��T���U��2��K!1:����Κ+m`�Zy�g} �ǝ��>r��=~���m�"��� n��#1��ڂ�{���^�"�8TK6pO7C���r��\��qW�����p�m	��4��S8�������&w?S�[?oI��Y�	w�։s�*���=af!�M��3����zVF�z�M�	f36�}��r3Me
�vM��o��Qg�[�	��Fbo���E���A�u�8��(b��E.���7���Yj�{h�P�^��1��������o�a��^v��&��)[��3��6C	�z�m���rh��;��Ǌ�i����O��#f�L����`kv���8}����յ.���V<��S�ٮd���M�ԩP��a1�j��zA����]�����Z3��4��XFpw���EȠ��\�b��205����s��Sq
�=�+b��>�nx`B�=�C��AOw!%�����r����hTT+D�pV�MF{�WI �D������6ApQ-cz�"�[
�O��n��u ��h$�K=���,��^n��֨��%�3Z�Jڪ�:�Pz����O�to���Ћg�l!�����[�AE|�Y,�N0�x���SxY7��Z?���ሀ���?ɾ�#[.w~��:*���ݭ�&:��p ���\���;s,6��b�RӘ�-����hKe!	����_�_����1
3	�tJ::�vLb�n�=G�)5k�|�	!��gn�Mn�*�(�g{��R/�H����ֱ�守�����d�6-�[f�)��G���[���Ĳ��`��6��*�S�K�Vw�=j�S'��3IkY�|�#?��Z�h�)e�rb���Ǵ�s�E�5e^��v2���<�@uC�l��J"��L�S��'�B�	�HlFJEsj�\�*j�Q��Bm03�[��ۮ�;,�?j��(�N����D��Ԍ5�ˉ�~���pԺEp�]dG�b�[�P��_d�e��0)�A�l/���	�(31�p]��[N���[�]��qf��$ъ�GST� �D�U��D�_��l.q.`~`���.�OX�D�	�S�땩|TgL���o&۸������g�ȈW*����)��q�_���ƙ�����!)M���C���u������5��u1��xX�TE������K	ͭ��+����>u:zK;��Xm!̈�# �A{�^�)����)���[l�<\g+2��J�~�)�?����2�!��3f�s�Z&Զ<h} �c��EN{��6%O�'� 6auD����R| ����PROȆc�c���	0�O�̌�O��Y��<N+�\�*)�5�̾y�S�v]%�/��ό
+�;���?�k���G�̽�lXV�>BQS"p\q�>�R ��4����\|����h7��J8���I�s=�9�5*|oy,�5"�xMdݱ.�w�Vf�q���puQT�S��CG��߫�4,��u������jT��G��]�`�xσ���Ҕ�["m*5��\dYH�n�?Ew�3$��5��ǈ�N%8G�d�Nn��-�=��Q�)^��8&�����=����qc�Y٬�:�o<R[�����SM�{?��A�����c��+¡�a���O�<��d��0�}�|��8�ٛB�z�}ŷ�A-��#�9����T��&�S�Id�(k�3�M�$T����k�N�]|���l��o5�X�7��Da>ƈ;}5��D@�}���.I%U��]�9gj����YJ	JQ6��e"gF_i��)��a0a���7S�;.���`�#h��+M�+�N���7���u~{[89�F� ]P鲦�h$:Na�M��<2�1z�1a�ea���}�|"�\Y]�n�Q�b����T����cx�C�G���t�����×���`�(��,r�^5�w��۸�6~Wؿ�m������DϢ�Cb霽6r�_{·nقBk�g���i��ދ��7㯾dwݻͭ��2G(ݛ/��?ʖ���*�Yz�9	�OR��[DN���D��-7@�<�c�DJS�k���>�/�<��X������ �Z�!f�g�q�G�nmi)��'?k���t����z�"m������K�Om�n�Z��L��Ao���&�,>n5��崐	)�J� �
b1^*>�3��)���듧���`D2�NiZns�|5�ZT�D�,��'-�)0Q�:�d�l���O�Jp�&\�B>5�&"E��[� �pA�%KV�Mr�g�蒢J��\.�1��/U�(�3�Z����)����^Qa�≮�c�-}��)y��aH��+&��_7H(Q�_Y�g��~M1�fRm%���f˯����<]q�v2�5w�kn��Ư�6�����iY#/��B�)V/$�����Η��F}�%�G�1��>�z*i���sNG�R��*�V����	��W骈��~Y��.�%+�ۜD���Z���]u���'��������eaTo��1�n�'����5�e"��(�E��?OMh����~�bg\!��@G[[Ff2" x���m��v�@̭��e�Cg��X��~� �qp#ڴ	;QU�>��0�!�ta+~\�deɰ�5��;�+�]�w�wU�Z0796m��5@3Hd?���q�h�������Z�N�Cؗ?�%o�X�<�.%:�I�	�2����ރ�
S	̳��3�����PƁV�X�n�k�[�Ƹ� >!�0:���r#p�Ͷs��;�mS���:��C�cr����d�,���z D&��o�kG��ק���.���#G����0ml���#��a�A�4�u"��ݐa8���}�9U7M7H:��S\�m����������&wI[��� �2́��DZ�T��䞽���<=����������1�Y��FKU�m���R��"�H��hym$Ç��q��gf�X��q��s���&��Tn�Dx���ڎ{���Q�	�H����� {�ʢ��y�/��O/�d[3��wt��nO�*�L��<���ěZ�G�xn�-5�5-�>�3DF����kȨ]CD8ǙU�>��\�a�O����}1#N\��!����ָ���5�ac�+��DM��]��2��N����bsD�o:-��1K]@�('��p���yQ��az|?+�<TЖ�[-hm���i�%e���̶%DQĠP��2(� �����9�e���EG��A ��O׶�K�o�}�Y���F+�V2ޮ���.?�u���
��m���ǽ8�k�y�4����~/��LN����Y������-���r�]���!��
D�"�8Ѣ[�ô{E9 m��P�
�Fi{7KL}��O���{%�	���������N���-���;-�׮���9poҡ�m(�f^T���	Wꘓ����$����"{3�-����R�MV5����OZ��)��ɮ�����s�T�?xN�Y|UG���<��m+����"X�����*�=���P�����/��R6]�^�$H�-I=�ش)�Q�R��=^�-	�b\�I`��.�uAO#$�sژK�(�vz-g9KF���K
 2Dl�1 �*߻e��Q��o�O F��s��pq����I�^���Ґ*4�E�J����2��ݤ(�b\E��j*q�l��Ļ�3�����ٿT0�X�4���Ĥ�\�R�_ɟ����}��a��;��ZU�2d�p�P%�{V�n-k}Y�� K�K�)�>�TY��ڢ�pb̬�u��7����g�^K�1&XJ�"P4��,>zs};|tg?�b����Ŕ]�UȰ
�[x�>{dh����h$!x �%�ɱ�H�݃g�Ũ��$PoC�p�
%�U[��b���] �}<.K�M������X���?%b�����F�Ԅ$Ʃ��������J�'���(K�
�d;��6)A��1�p��1r����c�9�ݾ7I�:�d֥�w�d��ֿa҈h]*'���֎z(�s;(i�ю�8���}!��+��v���{�V�\��4���&t�eڣ�@��³�'��4��Ϸ�I�I��	t��������*����@7��r����D��U!�S�YD/u��-ى�"u`IC��	=��<A�q�s�V��ݘ���M�6[��z�9��a�i�ऽ�M/B�@���h9�MG;�'l�ܾOiL��Q!?���oi�e^�>��EѡGñ�j��P^NU#Y��~H|���{���H���+4Al(�}�h���������$����%ֹ��~#E#���_���	*2t�?�0�E;�D9H�w
%�0�X���w��=I1�Ń/F� ��?�a�!�\�u�����h�P*^tw�҃�Д@�yc� ��{'8�F<����h��2�:/"A�`�:�����3&y��C�Ro�Ko4�Km�����5�