��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��w���GӆӖ��u9A�����&��;��h��6V��,�aXzG��̚.��F�_�G3�j�õlоb[A�Z�#�`#��<�B�q�F�4�D�%;"}/i������Dol!},��d��_��{(牰��์i���ӄ?P"�g�����m�	����=8p�Hl��!(�p�k
�X��jeP��x��k��Ȇ�rY��L�'��OΊ!ӟ���5��IП��i�f�&�)j�lW���QS��~�Iߣ�äT0`�7 ����v�c2hi5����F~�H�B�gVVq��D�1dj�̯O�zMy� �K�}/`��XfЊ� �D4]ʡ���2%��r`����P�2�(^i��<O��z�Wv�؄_�WK�DJ��B��M�M�K߉��	��K'�L��O� q��\m�	�}A������]S����81��;Eu?��Yb�-W t�Z���8^wA9u�����UoR���>�=����RŹ[�3z�v�������[�0yi�}d_�@�#|����Cȣ���W��[�[^媨�i$�e�1�/9�)���: ���"6�9|����@?���M���Y�	���k�9�]�p�L�<�l�G1)�^b�&���"��/W�!�^�R�Ɋ⦫ʲ�j6���7��un숋|�� Av��1$3��Vo�D��<��;��IOEk�?-l-/�gVjp����65�H�ð���t�L]爥Z�w�w��H�1�t���Y�]`�)a��c9�+X���$xv�>)�@8,�Rj{w�A�&�D�?O�����C.tP)�GH���������2�B(W�5���)V+K~܈q` $�|�a�𹏞̒�է��È���-��(L����*��3��$m��:���� ~3T��j5q�$>!�'���mO���#p�9�	c�����y,*_�,�ne�OHwA���RY�G��=U���/"��	
��	!p{�1Q��g����.Y'�f{�J�	/B�E���t��7��o|�T���W̑;����&�X�4�.����7u��P1�oT'�%h��{�>�����[�:*w{v���X�5;6=s����A��q�� ��u;Q���an��-��h.=ѨRZ����>��!#�)����˵e�#H�F����^,���@��޹Fp�I�ЊW�md�����d��vn����=]\s���-��E���]��qa�����2���$&�(32������K3�"�ܓ�L����;�U��"�[ٜ4�Y&��ީǪ�&M�sV��~ �nc���m���T_���D���	�S�;�cP���J�"K桘����%�X�Tp~��8zbPsOX�#��x��VT9�����t��Vl�ϋ���zF��P�Yj�+5�_���?C�z�6�`�G�ES���y"!�"A���pa�.>0"�-S���^
T�*�Χ'iݱ���İ���h#*�n�<,����&!.��yPL��DP\Z>jA��`!�KLzw�$��7�N��9�.J�H-�p���6��O�u@��jqr��O��P8��ԃ�]Yo"�.5|^ӳj�`Y��|�r@Ӹs��幁���� 1ge7�����,3W� �JuR6�������*zN��Q���)�,:��j_�R�Kޤ�^ @�b�j��kpV���y�OE�	��U)�<��/����j�Vt�x	]��r��ly�$xק�*�	|��ݼB<��@[R_�Ff�Q�E�N��,��9��L��k��8�C�~�l� ����jF)�ՂzE����ˌV#J�'}/�2�vJ�I���N�ՈIB@% ��r	��V�FsA����lM=���;���ͥ�P%�������o��������<���}Z9]�5�fƄ�d�����!��ñ��\���\���R+��coG��ѿd8ܙFu�x�5�I������]&_<���lſ4_�C�P|+�'\�q�ʾ-��?�L����q�W"�=Zq�����_����������U-E%����������?#TI�x-u��l��Nl�!�&�={�	W��R]�1TH���ᔟ&�������D$b��$c
\�v8����ϣ�����1ȣ�-��k W�˓�tLV�����!�n�ϻ�D��h���M�v�Bz��}ҹ���K�9�n��9�T��N�@����;�,��V������g�h*תjԔ+�D���.���'uwݾ�U��l&]t5!8�����Ͽ u��sص�]㢲/�v+ˌ7�A��m�2vaǆD��k��h�#�a�!��&LBq��<��Ȅ���:ax�������Tmm�R�R~=�R��C�Z��$ '�@��N�K����l���$����=q?)���<M�3���"�7�N�fά��!S��{ZL�F�I��7� B��b��60v��>USj-��{�n�6�3�"[0^T�o��\{q�9z9�N�k�l�$�����VpS֊2d�`ёe){7ZV��E��z��:��=֟l:�k��ہy�ӓ��>~��j�xM�77o�^�;E^̫�Y���M�-l4����~��9��E5b9��G�Z��{z�K�f�EUM?�z�c�����~��%X$�s��*�^*�uJfLB:W\6Z9G�9��C�`�E�
uQ{�f���ΐ qvT�� f�v����a`�c ِ�)m���I���<܅n�z�6&��?��g����U�v$f�k����e���UR)E�@T���e���V�4�acxo��ы>���J���8+4u���-��,gm�9�8��D����ѳK���7��4��"��P�hc-�ɇ�˪,�ۄog��B��h3��f��ϝ|�%j*�eٚ�l����6 �%�����q�y�V���+
�X�3��vbH������Q�̚.r��F���gK*�vu���+���b���̂͹� ���.�[�2�y�ji�s��`4�qS��{���������a�	737ղ�c��-�9��<#�N��@�=j�\��>��k��%�le|�WP�# �Ų��´f��LOYMٲ����{�Ӭ�(�hYR@�Ɵ��2���J��\�����g����C��s�::�F���{P�Ȳ�7]L��^���&&�4�&OkN�6��2���w���y*��˘�k`�t@�ķ3f�7Z�t	4�����\�݃6�v* ˊp0�/_$j5c!W�ET�o����ɍ�u�ˬ�Tx�Q���REkD��Lʡ�q+�+�=OE�� ����\�匙 <��$ϐ���tz���4K��2��2�P�B�"`f4��n'p���O��\v������m�� ���=��8ͼ���0�ݭ������T":�zP���W�P��Äo���L��N)#�|�j�=����Xb��Q��"�<n��������������|�^�)�	 6����omC�z?!�{������w9�o����H��u�N�9�{�p0�F���F~�I���̐���J)kHw�}RԿ�LL�'�������vM`E]��N��2���D]Bk)Poۙpja��v������%�/1͠���Ff��I�s˸�\FF1B�[�&���p�<�X�)V�T�Ϙ8� �aC���<����G�D�z�|n�E6��G��!�k�bsq!;E!a�/�����A�5�Ƴ���i�Bj��=��up���:�2&Vt���� ��bYGLZ���+�t����=6g =�����B��<C��bx����OA"j"	;x�;���h��7�rx��pq�98���������䈿uF6U��}�bP��j��ֺ[D�)'Ưh~OO�
�˗�,�K�+����h3l�YdC��<4������A�~6�|X�ؓ]3u/Tcߪ���O�����!A�{&�UZ�ɂPA���[�������4=4a���� ���+�����K���R/�O���VUO6�̣���{�H.��zTQ��[6���j�-��Rf}�=R�Ө+��"W��Ge�^��,�+x����7���n�KI�tɧS���%&����r�U:PE2׾��%�g|���*�{��ퟏ���w<͋kg��n~��!!�8l����K�ʃ��.%�w����G%����H���Ȼ.x������/wh�D�(J����]�K[`6�{*�)�����f݌�1�{�A��IZ�kP�*�jҕ$L^�4r��&$���U۠K�s�L�����W(#M�jy(*���֧W�sJH�� %ܢ��Xީr��!��F�S-V�m'�g��)�<�OaO[�[�(0�d�l����ywc�N�?��,���N�t���#�q��|��a!EY~R�������	��th9mJ�y��~�}F��fb�\!}t?$X?���x��o3|�s�J�UH��	��?vQ7��ɧ��j����ɦ<�`\��ff�c=Ρ:<$7�*ԥ���V���;�������QR��U�[a�pj��?�ߪj]��a�
�I.���p���o�C���m9R��m����3�vf��PDn��̐����N���+g�/�ȣS�Љф
R���EH5��`��ygd;��2|� ̺���^.i��8h�6�[kPP*h�\!&�ө�+F0CY�D@�p7Ă���5�[3��+o�w�j"3o&�?r�_���L�1g��B�5*��+�I���^��<��vY`��r�����(�\9Y��) ����AD��ߵ��)�h�/��7��}���׺6d���2o5)��S⪒_Xk8��S�l��^��-���f|�_mĿ|QG��_��/p��(��o�8Z�d�%)���l��5�|���7�����m���3w���M�g���.P_�8�����h@�c;��U�RiR�v_��[M+,�J��T'����GH�'{%NqXV����P�F`)��[+"5�mG�v�ބ�!���s��kW6rW��xØ&���;�q���g�D^��>or�%gCp�uJ���ksQ$@1�Z�U�콶�-�����>�b���Vem���\�wS7��\r��Y�}���fʐD�t�����l�k�.����"_}����,�RBZ�Lۗ�Ծ ��ȡ�aO|vR�v?znQ��;��8}��>��l��q�q7۩Q��Ȗ!��x�F�}p1�v܍̇��Cv9�v�����M�HM��Xa���M�loA�G(wۆ	.o�?�n�a�7H����Aޅc!/�e�ȟU��o��j?�Q5�$�$�|Q���a7{{����ξ��"����0�g Ih��$h�*���^��2�o|C�+^����%��(K�V�e!��"-dr�������&�a�v{-�������v���mO�'Bҧ^s����EF^����0����k~y�}J*_���j�)Dz�̊;)�2�
�5��<�?]�N�C��5?J-�r0�j1��2��S	��^�_ve�T�3Fe��λ��
GxI8��5�h�/.�δS��+��!�9�ư�i*j����4u�|�K��O��|7Do.;ڷZ�J�����Pa$�;��z�o�Ok}��EJp�0b���D�g�:�U�(�/O«��� �^�ijB��D���jb�<�iQ@0���@\z���yZ��M��� ���D�$C�\q}�C��D�*��5M�ր�
1�3<��JhaPh������R{�Qcվ7��@6�����db��c�r7��Ca�����5�~҅����I"d)Lfˏ�^�ھ����U=�Nȥ��	Nb�4�p>�+�8�cA�(�{�ƫs�C#���Z�
[��/%G�{p��$�Ed��~b�'�nH��s�m��h7�uL��8L��`+�l_S/�$�ŗG.8<vפ��t�+��'K ��Z�\xC�d�Y0(S�ue�S	AT�@y�s�(� �l�����O2����F8qWnt`FKɫ�=�w�"�]<�p�N�9�r�vm���R,a7'w1G�Y)��3�h���G���O�?~�PօTo?SQ��`M�7��JH��~G��}KQٰ!�� ~J����H��ߴE��2���BC�=�xm�i_3]���D���l)Z,t���R���9;ņ]ڽ>�w�����d��&��
�?u�訣���`KB~]��o�X1��R��b�B�YЫ�!>(�V����\�E,��~��M��q�#��3�f�m��׀����,bnݲ&L�Ֆŏ p�F�x�!�@����>7��L���d�2�Cŕ<DJ}�eG��/J���j�ϟjz\�/���*{�
Jf� ���}7��BK�Í�}��j縉�>^^p')ؤ�����7
���mis}W�~w�T�i�n�I�+����11���0���R���ml�$~�ٙ�Ȫ	�~�}?� ^ඕ����9�)
�@6�E�n�`bB��'���u�a;	���.��巢��1Θ�u@ʘ�C M�w�s/蝃��U4K�X�gn�����N1s���P�������P��uPpn	�o�l|+��;�Ye��O\�PƸ������&�!B�J5�{N���_A08���ހv�)�M���%���[�t�GU��|3Êߍ5���t 4v!��2� 2z#���(����Ǎ��%J?Ӿ�� �B���q6rٌ��i�C�T�@���g����:.����K������k��ȝ�כQ*O��,�>6�m�s^���ѝ]���~q��*"�����bg*?>L���4�bo4*��. ���kx��X����|����B��=����"�AI��x���
�^3,�2��e�vD�����F�xm�]���GG7�i$�a�|_��|SÉ��u*e����ОHNVv����g��G�oAml�z��PD��J�љ `�{�֊�p������$�B1���q��"s�����P�����<1b}��W�6�l��V�����D���B�"K%��K���B���ݷ��Z��T;CO��E�IG�'zݚ�͆@�!08{θ�����[r_αn�N�j~��E�'���0t�����k#ɒ�����W��T9cj�I5dd{�LVIy��Ĵ�����b�_�B�6��v�>�~ O�/@Q�L[c��R<.i�J5]�R,�	:&4W
�[�[^S��l	��yЁ�t�g���5�୻��PZ)���m���*���7��0q��ή��<� �g�b\%v�t؊1�vH��uO��Z�z���Z��S�?� U20d�u�KtZ���˙���{vH�L����Զ�T�d&Y���'it�>�/���ʩ'\8ho<,��|��@��p���Bd���R�Ձ[�}�p�8sֶ��@�6�l�!jN����y�ޛ� W�R/?.vPu��g�+� �r�����t��Od�	�]����6�&N⊅�B��U$fPs~騈�2�k��*Ͱs�-��.�``�����%����B۹����w$R�LY��9U��U��r��;�Z�=����ܡ-�o��kJ�9lr�ɔ�Lx~���MH ,٤(��Ƒ	Дy���Kd_�K�a^�ԟ���V���ciIy���o�n
�0X���"�h?bxgƟe��ޔ�{�^�)E٩W���\�&)�x67O��V"4�wl�O0Bx\ӝꪈ�@G5���[�0�J߼t���^��Zt7(~�QD�k�Q�qI����g|���1���"��.rqM"/�ˑ�^�B�D-���N3�䆖^��,x$�l���0~�͝��h�6�y����~#�wpǳ<�n(�̛}�%|5˞�R���v��Ȕ�Ղ{��WΎ�U	�j�J��*�k���}����m�͒�}�vOW�׆]w��&���\� ��"��7��&#_���P\��*�eH��v�tM�hؓ/��it<9ؕV.�''���Ag}�?�{�>���k����W'��=�>V�u�=9|v�K�G��X���6��s5��U�7ߢ�*T��A~]E+7t~񄐑?Y1׊�L���bJ�dn�ӽ �6m2�ӡ��I�t�=9�/攱Gqao�<�e���������+�D��ʒ�t)A���6�bS�����e%�8��ǻF��e��C_/�<�)i�j	�Y�{����Wz��H��:=�5�������
�:$%�%��k����|Oћ����<��8�$O8�&���bZ����h�f���Q�ם����L�(�WÅ>��(&R��Nkp��(wQ3ùq 2i,�
"��|���Y��&�#��3n�z�n%�&������=��+>��yk#�)|lP�l_����2����ެ���U0��|\�W�?[1�y��hN��d0�}R��0�*������.�Ph\.�`�rRW����ձ!_G`H�,�P)�� �'r�<��*` ^L���T7H����W6�>0>��wr�z�͆<�u��}d���:SP�(H��~�p��|�!	�r���br;(S��A�Ě�쀠!ڦD�ka<ᛊ�m�I��ג�}W�佲�AY���jQEλ>��2�t���"p4�Ӭf�k6�c��'8�N39���u��b|h���GH�r��s..(�!�N�q2�A���-�%j8o>��+f�����v�y�O���	������M��lM'�i,<��$�CyE��* �]K��I���+b��s����E�xB��e>|�]���,C�ٍyt�B�
��RP�_��*��Q�Ǚ�yLo���!���8H�60��d- Z�ȇ�$�:��31LQ�l�=� �	�2�u89���	�� S�Ճsɫ�(R��~m������?K}y�����4�9�,��3�ⱷ=Fu�P��ǀX���#k|k�!���桛7�KM��*Hz�`��	���R��vaaH6��[HuRg��B�ɶ�-#=���)jS^�����O2����LI��R4d����K˨z*Q$�E��	b�8 K�M@[��#��$����ޯ�/����]O;��"}��eu퉬޷��׉�8Y�/��߃K����ߪ@�(ů֛�@�L��I����z�i7�RTJ�O޼x��)��໷�O$��(-�ʼ��|�l��� �%�ѳ��*�g%���3C�̈́B��	�rX>Y��cż	�bC*�!%�_���t���%�9��==�o�������� �s�2W��|.��%q���(Ҟ��1y=���h���4|G�_���$�ޝ��^ﶕT<8�o�$8��P���s�_e�uN�Q�'-���#�к�<0��!1�%���.Ƃ>�L�+d����%6�y���>��Lߦ0�(�qMc���Y�b�3>wE��$������9���a9�I^o�l�#= ��o��,�3H�^ю���#l�˙h_�l�u�1{ܔ�2v��+���w�A�T�� ��i�q��>�pM��MZp݆�9����ˀ�F"��<��r�*����z��0�[��Wf��?� ��l�����J?�.3�<�dJ�������=H�mkR)�#�<x���G������qP
|�g8)m#:�;�{���lVo�����[(��7�P���wzʸ͞W]|����w:ޜ�<�C�-��ӱ_�.A%]3Y��3���#^�����U`�JF鿴�:�筙����5�N�xg���bYj���d������6r��y_�y��-�
����	/頻zS?~�UdD�_�N��r�`�f��ќ�o�U�iU۔�+����٘St%1�B^�L��=��î��ޛ��[UW~ȯv+祡�����0*��	�T=|2�U�0�Q�΄"�Q���aH����m����Ai�Q?ɩ�&O�8s2��ɵQ��X�N-O*�ٕq\%h9=���?.�Qx.�t�Ҭ����'�;��+�vC���K�F� ~;sae����{����e��f�/�Ew%:DI#� p7��
�vW켶{2��7��-��<��F<]%�_����w�_Q� T�G�����e�����Ϲ!n��W�����˶S�E�7�;ԏx�j`-Gؤ� ���LLs@�c�9��*`]�� ���A�~Z"k�i�`��e}o�=n� C��?X������\�K��ϳ>�<8�B��=i�����A�?�b�������Ik�<F8� ��i��)�A�,/4M��r�#��g��U���-eB���΄g-@X��"߂ȅ8��Z����G	���[n'g��B��q	�$`�h���i�H�#�e��s"��r��de�}��w:ZY�z8[9-���>N�-%��$���ޤ��q����̬���m��*�0ωVi����Ԕ=]�E:�o��a{�7����#���!�t��*_I!SDI,�}����֚���}�?���ʰl�]�1x�q�g �T~�,����FK�A��MG��f%J���WM{`���Ŝ�O_�U��#���'="^�dnE_A���4c��{�b�1ܾG��_s��V\����V�������ʠ5vk-��N ��nN�3,�܄ͳ'�)��/�ϹK�㮟_����P�$��A#'g�Ȼ�@ʛ�v����;�[�7���! �?�?�ձ����Ѻ}��K���f�Eg��<=dX� �g� �� }!�B~��
�u�z�}ﺬݧ�5��8�nk��պV���K�g��a�S�L����U�#�I3T���`UQfN%����Q�^�D�P}�n�t@���ԑ�� �Y9@�* u�ᗁ��y&Ԛ���q���������<�V\��v^7�7�j�]�q�G@�
�=���q<���hx^��i����QN���$=�F� ��u��l��++l<WD$����*a�b=7����J���ҙh��߶k�4w�/P�A��:��g�j7�%�Hh��Ngs�t�ӂ֕���1�r�.u�����AxJG�=�����b�f�9��)L0���"I�F���-��x�`[Z���pf5,�Dַ\�Vkʌ�k��-tK\�Ծ��KhE�"�$�;���w7
(mFإP��o�Z}�cR,��DWÜ f~�M�D��aj9��B(��RZ*l�4N7���DE�5���)>�t,����E����f�c�f�!�o�b�X%ylJ�<��E��U�s�实p���G�P;F�����(nCH��Av��^��q|I<`���,	.߁��hr�]���S�0��L.l��,�:��'�<��R*#���e{�`��Z����.��<*��
cE>ȷ鎻�W5k�|��o#�a�IW*7
n8=��������9P@��N4��òϙ�8H���&$�R��Z�y̶�B�
����L��+q{����T��Xi���3��H�d�ix�n5�qy�֏d��1w��/s���-����aF�.'�"��	�n`�E�I����H�_��&�R>�.@YQ�y�9I��=:a�̸�_���2xz�ֳ�k�	�Y��lrO�?C�A����rYNYWd��HO�����=�BԶb�rR�MF��l�4J|������ ��nR���̚�pq&䣌��}�������y��z��4ZEc�ocG���:R�$����6��(�Q��7l��Y��VW�K�W���;�/��)Σ��% ��d\��lh)o�>��;\����'��H�=�!�ߣa�M��$�'ҩ�6���rtV�K� �ch��)+�G�����kx�Ģ#b"R���ú����l�-h���BnBb^,&0�����xl�wuӅ�<�5y�E�y�<��Eb�3����8Ŷ����K�F،�
԰3xU� ����-5�"�3\ۤ��I�������Ka�vsn��f�!�W���P�����pۙ��#���m/š�ϑ�jF�8�Ժ��k��`�Y��"!�ꙕf��n�����ן��(f\!�Ξt��!�`����
�t]����W3�H���F�?���o��9A��t}�6��VM�H"3�
-����@�c��/*�!� #
f�D��7@(��&G�Z�b]�DmSq�:Z�y����� �Rfi�ǐ��z���aIz���y���Pٵڞp�<O� �(� ��T���ZWL���ɻ��
1u'��i5G���L#r!��V�@��@���؊O�4]����s���ض�[u�W�K��Kt����6@g�?�v �O(���WEH1i�˕zfH��lo�s�BФ.�AS���D��w�����,su�$Mg!U���z�[�O�r3��@�����b.�-!F�hZ�%	�9^��c~���m@A�Ƿ^@����<Uı����e.������.��T�U%��O`��]���X����"�uS�u�:���b1k���.]�X_��=ˋF�� @�zHݻ�е��T��J�݂A��~a�柰\!N8��è��Iw�
k��9�4�Ɗ��
 �E��v&��I��-��
Y����QF���c����{,}偛����*�<I*�X�bf�f����"U�m��L^[��$�Q~ȇ-\,<��@\���S�Ӳ���}֦D�6z���%haʕ)����{�5��f���t�xv�Q�0gVk��x]#S���k��J��е�홐X�����I��q:j�"���cS��r�6G6�ڛv��_��_�p��PSm�
z<<�'�_#{��eŪ�8������Sd���x(����c0#��
���Pt!��Z@a��S�>P]ڿ�8���ʑ *�;ǁ�a�P#��!][�ہ����yx�?D,��	�4N�+���`,Xq�җ9���1�LQ�g�6�+l|�����g���Y�l�mm=ʔ<g^�������-��|�43��`}�A6�Xױw��u�5A��{d��� ��r����x[o��L�7�����e�-�=�O
vjE�Rڰ'�/�ƾ�I!s�/�b��8U.�.�3)�i������Jȁ��&���U
��#��2�"p����� D6�.Jq��UG��%nS��Tڹ�&I����ڄT�¬�qe#�^�ę�;��#���Y���u�PE�ce�D*�U�N/�A�q�����t=�/e�U[	�@%8�����.��zJF�d�!|mQ���8`����&ț�F"zE�K���AQѕ���f� '�����:z�^� �J��$͏��e�z(�)��/����Y��ʜ|��}8��U/J���2��0�^�?aSݹ�gUz	O�&6j��I>>&Ub�Vj�%�:P<�}�&�qe\����x0N�wx\j�ϊl"��U4�;T�x���J���V��/���?XI.#u�������n�XӾ?���l�S��$�.�P�E8P�@�@�՝�<=hn�X���V�D�em_P'kx���#%�摳�8h��S�đ{�)�����I��N->��z<��&���c�M�����`�L�z�F���*,��{����F@����:����#yI�CG�EPŧ4Kv}�b㭴��Ѫ��<9����s���.���H�Q��f۫]��̔�h�-l�Rmu���:U���N��20�c@؞9�LO$A/��$��
�@V�Am�ffwk�&��l>�}�[F����&�.Q��E��؟�nOCz���=ܢ��=e l�z�I�c&jZd�V��Pi�/X�d��b���ƕ������3cPѸ]�x����#EzkGHW.c��UI�m�ޢHW�D�"�<��Z�z�
"�9��u��
���jCV;�5�봓R�+���q�h�ۂ��\Rypݯ|՞2�H޴�y%}i�����zn[��������;*�]���3������� ����ۅ��%C�>Y@���
��zS���ύ���;�d
Y��<�����	���$w]H�:G�f�"XY�n���Py�2���ئ�1i?�a��QQÊjzF�,���;o�|���݆�5��"*w��	�Ut(�ܨ�(�|�Ƽ��kA�����Sl�e^L�U��;��կ�l�yz�!(ԔҘ����g���(�Q��E_X���Y���cE�� �s���T1hj�8��dV�@���s�o9?��]G/��lm�����>B��|vK�
�s����:��ʰq�h���e�b��H�PY&���-�i(��n4J�}�h�:qreO��E� ��p+�G��U�;M�,���&s#��I��J��'w;�6Ȅ���"YS��;�̍f�x�OG��.��K+}nk�J�#�eP1��F�vV�;}��x�U�v�8k�}���ҳS���֍M��rNZ�Q���rx_�G"��B��h84ԭ��M��Ip�h�ڙ '�q�LL=Fr������Vс_���h��Ez՘�!ٝ��/٣c�^�>t>��U�U�/��4i�n��� �.>�b����$�dx�|P)C�y����V��,qD���2�[��ly�i4H�[�+���ʣe�ʭ͘��]�h�3��-}e�`�o����|��(��Z��3KI {���R�˖�|C��@|�"��hֳ}�Z�����#	@G*�i�g����aj"ruMy| r<o�f.I���t�߹�q�;	ӣ��a��{;��>ϰ�\��� ���w��*Cx�@0�~0pv��v�F�$�r�.��
��kҨ3@���j�o����C�$5�0�s�!r�d�JP�ȩ�c�LM?x�][��� �Uj+Ku46���w]c\�S�~��R��`�i<
���ޜp�{ث��"#E��"���X�fcC9*GPh�荾��={�h����EcE�z�h��qdط�t�\T:R�Y�)
����ϋ�֓��)i����h�J[��s	o;���/)*�"��]�慮{E�ڶ��S7��,)�k�̯�ڒ�4��ᢣDL�rq�y�9�'=5IY�<T���&R?i\�>����/>�v=7��~l�3��ܗ}�!��3;J�]�Hh{��O�>~��uA�uO@�� Ґ�ĭ������ck=	�����$��NG�SGQ��x= ٿ�n@%и>Zſ~�ݣHo�D,��U�?S�o�'�B����:�ϧgؤ�c�������X%d���i7����Ĥ�z�.�ɪ̷e����p�`O��������7��!c��2��GAo���0Cy0���QS�hBBfu�ݾ! ~���|l��1V�<��i�:T�"`��^G���!��Vg٨02�ǘo�=L�SS���-g}�'�g7{�����.R���g��I����Ȼ]�vF�3)xf:p�8�:S�隘��S#��N������l?8ۻJY�3�?�U9�4ҏ���W��f�D!�*?�8��P�a�������P�q
q�E�p#����yN!T����Z���tP� �$8'xDOJ��8wL��D�M߬�xp���y0��Ei.Fzi�����v��e���|Ң�8����e�e6N�V���G�!d{y��U�D�c�rUx�," _�2��Q)��&�m��tsR��E{Ov�^LW��fpф�^0��7׭�L�S|}8>C��'xԡ�b����m�*Ζ�l�H��a��?Ĭ�?c~�WC�-��1��=�L�G��=p�6� d�����0�~k��5�h�L�1�$s����,�q�U�{3zu�Ϛ����](�&�a�C����S�K�~�N��Ǟw𣼧_E�����y���å�ɳiO�����9�܏�2���}�֮X���)���+1ET��q\O�6%a����F����57�#ln��h���Z�Eۺ��ȘZo�7�:W}���A����]h�>��]��Ϡ�-h��҅�����3��ò���e����&�f�Uͽ����an
]i�"��f*�	hU)����M��[�5b��RM$E��L�/<dZ�%b�1��@�5Ǽ�N^�	bd���I�E��_S�г$��3܋����ɝ�6psMO���q�"y�3NS�eg��7~�֍/VӾG;�i�=��'IGC9h�U\C+��^_#ȍ�`��"޳]3�@[4K��%}�t�!��<��)ʓ��֪j�l����@�n�� �)�&�1	�R��֙"��@�FC��L���7u��4M��+�S�ef5(2�u���X�`�����P9�ۧzRjeK��&S���������7�+�C�`�p܃�]V��"�9�YƠ����4�|�����.�1�|��UƇ�����Da+����1����`o�g��mYD'�E�1�.T~\��P#� ��̃@��kA�.^,�yZ��}%N�W��"URN���.�P*��c�M�s��{�WK�\���҈��^�[x��u�.P��;���q�1����
�����lGjF(gd+	�/��jf�Lf��ܨ�T��e��ٚ��?m7M���.	����3!��E$R.S8AѪ���:��t�U`\�?�i�X�y���qz����k�ߐ<���ż`����	�J�9e�(�����	����ZR	�@6|�a�g��� AE����_i��K%�����ː���,�ܖS�P5��Wh����`X�J�9#�F��YPM��c��Y����(w��\��ք]C� �+5��k���p^�u/ȃ;"����V3�'����Y;qϼ�ȋPH"�����DB3Ap�����K*z���:������H����c�5_��6��­m�j
�z�������lH�ta-�y�X·:`-*t�a"��\i��p2�f�I��:_c���"��z�~:s395`��w��a,h���l3�Fz�$c�8�ҫNiw_���M���\�vP5��u~�����/��A�}�P���P�a���Q�Z��w9���!���O���ɪ�:��3.O{R7s����"Y� ���\��W��3o���90,�$���Q<����nᅻ�ݔ�ި/��Xr�W�ŵ(��ǹ�jj�Q��=��u��E�$�i1�$}J����I͝��{q��+=��+�0�'o����ژ�7)5�̀���_�3��ވ��UI�s���E�7��L���dڝ-2pV�m̊
ăGt�~�mO���h�[��������&���Zk����3����"�� ���F[鄉x�d�_8�O��~EFԢ�"^[��'$�O����^)�T�)�K�{R6Y���iI��h?f�C8:�ُ5���&%�R�(y�i��{y9��-��P=u���rS{Z��x+A�6Iq~��J�yg�LS��a"8�õ�!�ݭ� ���z���u�7�m���lu�2јx�%���Iͷ�6��[��)�7:-��C2��'L��K��v!�N� 0��I��i��/�o�Nj���5�ώO��zR�Nw�P�J��|�Qy���"��Ѻ�R�Wk��4�����:1���&#K�|��A����C��>.�%�fMͷ
����g��T	#iu��0�L��c2�
�kfd�𠜱�8�/����3٤c�|^��Hǻ����yo�ǤbN9�
�S$��k�eg�o�+�+-��n�p�s�0��[��h#MP�/��L3E}�?cr���u��3l�]��b���D�-�1a �8��,�j�c�%%>ʐ������)p�ݷS�FR��qZEUU��*�!��[��k�ga;ҧv��S�wT��\Q��4i	��$���UB�\-^1�w۾�C��)�$������k�� ˗8ef�����"�	O��]6��a��k��.M� ������z���-�L�}=%֞O�N�è��l��ڧ�O��?Fw�O���]��-��kjԳ�X�5�3@S�+-�[�)���E�tZ���д2��	.�~�Y��,�Eer�i	�B�l:�l���l�i��6�v�!7�N%0�@�kJ#n���_+�| CO�Yx��u���inv����J�������b{f&�x-,2D#a�9Wy�-����gv�"ǥ�&��>�H�����M*�<��q���(��8�/ ���0�yTx�̃�!O�:��W�g����N�=_�6?�&2����OmO*�AC�&X�9����h���'}|J��-&#{�SQ�D�˔R�c�UΩ*K�tl0�$-�onx5q�I����CX����R�+F4F79�*��T�pU�J����Q�,�ׯu"���S�53��$�6(W��.�l�Õկ�X�NZ�S��E{oS��G���b&�q8�Noj�o��|=�F���I�U�zj�����]��������Muu@o4����r�v����X�Ȣ�{��S���(t���E�Q�7x��ԏ1�74����ע/���WU`[�;��fD�Qi՝���e`�Y%�9C[$����d�j�1�M5{� ��M��KBgT�#9V��������e:Ż.-@s/pV�ȋ�e��;�י����X e:T�K��00����$.��ʍ ��o@���[n�E���֊%�2��6G� d��K%4��%�xg�
���$�ߠ?C�.�Ч��I��ZbQl��}�k��vk	r�:`\��$��}��D�%��T�ҵ���]	pƀ2���w�Mz(�9͔v�?Y��!a�^.�E�d�!�m<�G�w��&	���]p�QP]i譄_ǖa4w꨿�� � ׂl�rSڲC�q�"�Ci�>8���?���P���S|Z6n..�q��`��kW�7��J}���i�X!.�=!�aFyN��387O�'�eq��'���s����I7I�Eԩ��G	W�����G�=9�K)��0j�V���/��	퓬��Y��=�lѕ�?Ȁ?�7����  `2�n6h�M!Yl/V-��jw�$�>0�(t
�@AB�k�Ɂ��6��N�md����b��þ��k��I������B^�1��9*��=c������CYR�.«��.��,*�zOMV�<X"���_r��ḏÇGN�� bu%�N�?�I�����VHl�$��MM}�ol�I���xJ�~��,m��<wLi��w�����7�Ь�w�7�5F��}_:�`9�>g���J:�1[~�u'�	:8P���V����x�DT�NK�\�k�������y��}<����7�����Ga+dv���O�]d6�
pT�4� ʃ�)��Dȥp���T2i�H&�^wK��k�.�O��Ĵo5oB��vB%F�W�"������#����/�)���Q����Q����)��˵cL�i��hש���=v.㑲tH��Ъ����k�G14Ly��Rq턨d��3�R֋9k�.��a��R�:����`?J0¶���8��̬�?�4@��^��:���v�`�8'\#:�'4�ښ@�����%n6p��d�.c�����77��n��c�~H`}a�c-�7:�A�d�����3�F���4b	65˖/ Xb7ԥ�D�8gI�U
:"q��b�\U�ޣ�x�����C� /�-��׹2�t,��N+��!|<�qB_������TK�(tm�L�~�t����+!�YR��{�}+# �lq
�g��f�V�@߳��h�_f�ڳ^���"[	�'�GA��DZ�6��dԺ�岣���*5l�	���'Hn���C��$@q2VnXHk"BnXw¾�D*���@s�ڗ�ܤ�i���찂Vj,��7��D8�+W)���{��Z���^T�C8k�4\�m�H�df�(3�z�����{�L̚�S���bv#�b�h����9%�o%�o����&�T88�%��C��xB�C��K1��A����{�&�{+-hZd}��蔺���Ġv��5��Z�sxX�.�]��|���ˎ>�Lr�[�{M3�HI�e��y�c�d�r�Z�5�#� 	* ����ٗ-���Q
Fh�a���0nr���Ƽc,�m���a�cO;1m�����׀�42j��I�T�yaWye;��Q�uu^��0y{Y*�⮢�H�$}Q'Q7h��0���k�K\��)��ݷ��F���$� ��p�榵��n*b=ݶS�?��l����<GD�)KpU�ʘKhE�i�ޑ��}���g�5�?S3�$W�l�8No��P�M��jW:��l*jqN�Zc�:��pSbw�����$&���O��������Ԏ���:eBN;͸b�@N���.�T��Pų5��� =X˔��Q@��8�t��y�[�F���29ɽ7��,��R�˂k	��H�PU�(�l�1�W7�R|���9����Z��L+����Ə9��1m���M*D�Ô�Ĕ�lh�!� h!)Si�,>�Qv���8�9oJ@{�'�{��w����/ƹs�C�>2��'lH��u�dо��g��ɋ��+{�I�$����(�#�Y�?�;�BBzY7�)=T^�4��`KG]��A�N�T�w�;��>h�@�8������~V����`����m6�X ~}r��R�l����
'��S\n� �J	,`�#����0�a�l��X�OFF���A�d<�6��%	ܳ#�N��\� �::]�lkz��e��={jJ2amƩ��Py��z����}���������a��4il�U7B򩉌<;�,'bcZ��>ڮr^Z��bP�O�����k���R���o6�-0l��w��ܵt�q�in(�S�O�m�8h��)�������f]�`5m$*��^e,RϙÄ�r�y�4�ɜ��}�qME!��4�*~@��|�̇I�_9�FV�~C��Y/S�)������o�gZ����]�MakMo�B��6�%@TSeAi�(���cӨ�4��؎�U.Wg"/f�\����/�m�J�I4�,����h@ G�$)
�8��s�a6�ܑ|L�W�0�N��/����zr�5n�b��Jz/Rk����� �6�헶�u�k)�@�iM���KI��m��M�
j��{ -�]�B�A������{d���C�v"����*�����6Y6q<h��a�g�@�!�<;]��7���W��L, ,���na㘇�(IW�#�DUٞ�T9i�tm�q�j�	�f�4�l�#G��t��.�!C�8à��k��O�5����c����d�T���h4>'�*zGb��rN�B5�R���V��b�C<7$���q6�n3�(����|T���f�07�
_)"��!R������J���p�0*M���a05ճ>��GK��RaU��b�a��ff>�Xic��q3.N������]����d��<�q�/��^���lAC�@C|��l�#{+�]q���v�Ԋ���r��)\U3���o|c��đθ=/;a|T=�2i���}�P�ԉ�fp9�/����6�p�l��\���aQ;��AN��&�X("� ���eW�Q� �e� ��"E��I�) n,�h
v\�u,"���Y`3���lά���U��[�!X��}Q#�6��XD����|ۙ�Ct�9�"�%�ͨ��>�y������@й��mo��aY&��U/� �<��_��il��R�?;�{kE�����D�Cb����������s��s��xf�q�D=�nl�	�l����l�"��{^�qpY��<�#^�mHO;I�R7�3�4Y�#�Y"�ՃY
��Sy�l�D#���W����=ܳ�CIĈ
N�
}4�9��������2�7��m�����mV-�G0#�/���x��⳽�TN��Iέ�m�bk̪��6;����P�j��ޖ؍,�[��v�pT]�@N/�w��tFsY����d�a��̶�n`�n�}�P爸���I.��տ���Sr\:w��!L�����q`X0��Ed݈3�T�ع��z~����oK����No���C�����>O;��Z}B�ƠؾB�D�}��+_'<�?G�s�S�*���iv�Q~���)G�(����	#U��ﱧ���f��k��ĻƔ\�w]��?ږ<EF�~��_!�
�?y��iE9����R"z�E���5���9�~�!(�����K���遲,�r|���=7� ˡ7�Y��?��⼺��1V�Ip,*�Fc�m�u�+��pd��鍦�:��?��'ٯ��n�[�,�hAS'�J��¤����RD��q ����4�^�_��_��T��s
Td���q(i��]=|e-S6~9:����L�Z��l�o�W��"R/����*����|����.wh�
��u:�����ϑb,�Whb�����ϒH�"�;�)I>�� 0
r�q�p�&�h����*S
�v!P�E�ilhE{��ަ�/P��,��Q��4M�5���T�%�mF�I V�a��ۗAw{��M=�3h�W@��6/T�m�%ĩ	8PS~]�0�Z�>��Hx�8ԫp$'���א��[�[�e\�!hm�͸����̰��0��d���!*��k(l^��.�l]�����a�C܅x�I��l�3��~0O�J�>��T#7�����ڑ�] ��|(�v�6/�)Xj Ľ28;��>�SS�5�1I��B_������]��;�*"�֒ˠ��ɞ�̗���ּ���cynD��O/ǖ�#�.��&���r�V�|�.��F�|��{K/�� �T��Cp�A$�k]�N�|D��*����@z�s2PF