-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0SnV4cKm0UxwgQdfPaHSp7Nxk8QU82zoog5AfdoydTrV/cgesCNLIEC1CJ1Thp7BlXF7XmFQEg+7
qK9VI2gvbtD0tw0uiyPD847PtbMs2CaQR3W0HJKpnC9CmXFGvGeXg4//VQbILJxxJVQhp70GEsc8
6C4D14oSUEv3IjKP6E1vnoOKJwZ+gbiB32A51vtY2l34KZ7YAmWX6QZz0OkMM8EaTvPiMY+gRSvr
rtr020l4A969pNsP1NImk38LeIy6ty4zGrYOIAlyNK+surZMCnL+hHx+6NMtHqo/o9RrddB80q2F
Bb15tteBDY+f0IPXQeW1FxK+XvDGD1PqJVhn5w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
LtPEHI7Q0WM4WMxKspC8uU0XxDACiqPWKecm0j6EFQQ1Npp+jc6TCkTDjOosl0EnxhmL3NLCsyJO
Sb4BzJ/BbIR8lg3CLeenhvs1TKZ8cJgAN7T2U5+Yd4jwbmKcOgxJf+421eq3nJ1Op5GA8I071FiP
Ks2rImrlRZGbLO6n9HEqm2j3qoePm76Le3jjByR4A4LTj/lROraXfoZTE2LfO5Aglyju04FL32K5
jq51PEbdeE+Ey3ZB8JHw4cTS1dB+wT0J1qdnfJkkJFShVPzgUqzGaPAgf4NYUJpcLFpmuWttTUJp
1pT5mNSd7B4WJfJZcsl8H96ThvRwPe21oiq6cuS+JXmfpravdFcDQbkOce+pBPWsXX5L6GjYTjgs
riwbJ0MmXRhvW14iO6bfcICAmRxy9Jgj1V6aRj+P+lQROoAW/03pyPPz7BTQ+Wdl+ZZjfVjRti+B
F84jC1edAJoroEi9/6ILtb7fnmCmEHE0khnpPsuLtHKZ64P6k//ja1CEhsCkj2YTH2Idd3fJfTIH
V1QSrpJ5j4iQXcSFV9Z0bFCC1HIlMHKPLL7w6YWccgWrzVSEB0xh+i7+pgM224exu9O8KACCjzRg
30sEV2NDVd+nQicJKpTcSSdO7mur6Fsp8V3+8t9xoNtzOHvFbttsyhh2K1mCK1oMm4q0hy6cG0Gi
4tUeJyg7SHaoKfiqLVWvcvF4L1Wo1eZTYRbWpXMIDnbdJTWQMdYNjYFByyEoRIPkKohae8KAEWYx
4qGLGrfLVp0TyQHCufIlWQLZ9YAgkrL0BtQhEAG5t3iajQvp2eFmdvv9CvcStrFFwesvg1KHqxfm
vBqY0FDQi72Jzlke9UIwLZ2UjgWXj9bM02KESSuRWDVReJCAes0ViCZ95eRrc2YzbeTh0Hs039zI
sLO6ZZ93pl4uW8baaTq0KWdXS8oH2MsFkmn7zYNhOfmjDVeZ51kGvTkXyjG9680O7BDklyBA1Sqj
Yrv0Z1Dx1+EBS/hV21Jwoo+BcZe3QQqcvxbEjtNHQG55zAa2ejP0L9DB5a9q1kuPs3hDIkSoVs4p
fh08qHweJMc0ood+Ez6NE18o4LJ6Z7lRaDfqNwFcqNfnGNxrtmxzIJVBlDVLnyFZAIg7zNflJngk
4AAGPTAe+RNNOD9/luTR/oIdlp0DtirJLKDf4CIO5nMXMKxtLBDYxd0H4EiQ06U+qdkLrIa6avma
kh7IWDDqtV6PQ8SEkx4Pn9bphxMGVlN47yHdjFcUWbeiuFLdNgFmH27CaqSlWuh/RPT1G2xxIL5+
q1JiRVJqUj7iQAaK+V3RdNd7hAGNW34IpAS/FaKi5YbxC5UqYvZ6SuxtS3H6LQQOC/vQZoaRrpeJ
ZlQETlCLjot+ioIV8ATjGisTI2PHhCTMNhkQE+tgs+QBq6xUhpURCN2KqqVL2KQvUi5wSqAXq6QC
QC1/oDUGPxaC0+51OR+kv0H/eb1YociRT1OyOBIhBLbKOgw26+NPOFaxppMsovKSBkgY4QB5ZCbQ
El1g+xi7FYVRuFbEBfl1thb+C8gONvTGyQJoRV9jfdkyrydlnON27qUhRJgDkASmyPX2u2kiiIxl
B6jPfaRC5uD92aPUkE0Z7kbGYP6DR0Y5CIhOCsxbVbgZXMT4LjdQpjuw1Scxh/vUPQQcPXs3wGhY
3m4iK43RfhlcWVV4Zvtr3zBovkLWM5ja4oltSgDJP/fKERT/vxZaDBFOq/61Llhzfjvw1BNUaaMb
8FEEleej/s+5FkJW19D6GqclmcHReMFjBBzqeP46Xn3GR5yMzCCSLu6aS+NaOi0Wu8UBx6WDo33a
isHx5qcge44m/U1jjQX9EGJemrVSRMmvdNTNuyT3g8kdOznxgH5kY1qDvLAI709pG2ebG11MI2hH
ACtvUDJjC/kGlEHq8aSlV9RDFiWA5RnjIzRI3KLIEnlatMx2AH/9XOSdEiTCu7pcq4stQy5KhYZ5
JgJ3NwgrgJl9oztlXeyTntmcttynYWAtiTc0WrLOlGXwMWi/9e1b0tGjkcCgIBCxQPRLbfZ6NlrF
zW1b+dEnYQtbv5tjsbmn9DU2TLbI4xSa7kEyr/7HEREtyMBspR9F0Gv5sn3uYUbaezII4OE09c2j
Bz3urqzY3H8dz0XYBtBTfRT1x4xHTha1CGBQt9G2W9+cj5vXy64yNob0EVqbCNxNieUuC6kBEkkg
8A0/f8/fEqxwoOpskepE2MSQuO09j847rzEWvP5FEO0Em5Q+2SHyKBKqRkSJHZCGQ4xKMgoyBYLh
RYliKkJb5vsWT4CKFpvWwbW37oPOcUQd4DNpcA3DWhzTB/sx8f4CdvJBB7nNkKzNyOROlOs8PN4p
Nh0cuYt46zGH4ynT98HuXthn49HNOvLy3tXGAnQArmlZgi4F6x7R0QaSfn36aDYHN5TxUGQW/p7d
fmev4i4BqTz4wX23QqKVloij9JBctLS4Hw5TiVkPFN0vMjzfPGL3JaL6B0qFy2ru2YRa3+n2aeYM
yHGuKYC8TZc3QjQIYX4+21/3qn8B458Go3g+QsxJlszy2mfk0lBZb9/Em1N6RuIMB2ztChl131sZ
Gh5OJibNOnO5AN7R5CI3vVk5RHax6y5HJCGEj2jDjtdIe28Hj7nn5Giw9degsQSfR5wwRV77LKxM
8yjH7E4mqJsGUy46hkiy5KaJx98xCOlfvU2QmjJ4pe1NbY1/GuXkNBoi2FJc60QuCFzU3sdSogeV
Vn0u0QjJEp9Azg+N53PbN8YAAi1ktEwF6l/f51xgTR2QnQxzPCOTH2FD/LZhTXE2fZbYTnyxY2Iu
GRBxpIjLaNrb4Dln9KOI+7GnS2GzUXlgwUq1JcsqzdP/ywInEN/LwDd0ayU+b92OI1dcZuxmGQva
B6/TK/nKwwlGmXOhXExfMDNQjKr1CH2cs/ghLTQcOlCPcVSDP3+IClvQNXZ84j/chODjxpuKybd7
SQFXpvocDI0/XImShOHNTyr5iab+VhJjAc1LshV2M/FJO/gGP+DYwoLib3A3IAnPJn4wPDn72tYR
RzGQCv8ru35xxLeOLo/b2a+4dqEvx90BO+LigFkICUfeeCckjdfJ+hVgcBPbFqhfBFljmvy01edw
AO5rdyCCHfekF1FL/YLBmtmHT4AgrhqlM8w3M0EorWfzqvnN1LeoFFiET5A/P98ymrfLsamC4v/m
fdiiNqz493NP0u2izSBnq+j2em1kA/z5EjknFgROW+WVnH/qScMPkpaxnJ0rUbba5DSm5weAJILh
lBScJmIXM5NWrg2XLpS87/bdLv4S2uIijkPTsv7oPH+wl/gl7p+QXp44k+JafoLkkguwB7lsmtez
OfeUeN1tu+JmUok6aDQP1Ew2YFdh06U4e9GPdW3mkNpv2jr4WPJOla9xNd/3BJQ9aKVOwuob6enU
6nu4Zi4E+51QRsaWB3G7DfryLmZv5YM+Hn6Nx6lIZG2wvdT3y72Kpw9rc/KL0Y9vLkSjGy1tq1cu
PMbpI9/uzZJmYFPjCeJ/n8Wol2xovb/UoOt1kUiklq5tL4a4QH/113K8AXs/a1npDJKLityB01YV
uccraUhEdhB4oWN3ZAclmX7oaxM84Wsy0rWYbBoB0mVkDjOgtGiqkdrAZNE/tUy+06tVOGM2YaRW
mFwgPBuG4VkeEkEN66QF9IArkASqMjEJ+JK+t/9AEL/tZ+BTQWO84fVs82lmcp3rfhetw3bJeTP0
9aCy7riMkHobKeNLc8loZVGgDRLuzATyzMHtREn6HfpIKIinOH3zU0pF0/5iJLEta4I+NwuRXCHn
y/GuWJwssnVAP9I9EPNRMSrVgV7XvTQgvNl4R2lJ3uQFS0bfujoTKR16ord/RG6XS/yjQjGUHt6f
eryVSIPOdYFM6NpuysaB1kjlRBXCHP+50FuDQOZ7kYMEyk5rV2sSh8P5JrhORiYh14bjqarp8Nry
0fohEcROHaW4783ab+GVCMsBMtAF+EflrjwlqRW6IHGdJ3/pyvQUE3XUcqkRSWw7Q/GQ6U68ah54
4+4e6xljMs6NdoNoAFTlqkeOuxSihQaqj2W04QNmRFYl68GIaQPiM2dvU8KZ4sAQG+qtMOhs7ZIr
B+bStuFUBxMrStiXEF9Fw3IXo+1e6Mgjkbu8sIaVJL8jk4kQlU/eHHmL5VUbaEkB6ias96Iu86+9
UUEgQ5eUtHUAmVZLI8JqSyPi2dKg0vC771VY5hSR0S6E/MnwuIQbEq+rrL1eEhoN/NiU4hMLFEdL
pJCPfaJM8YBW1X3NHjJEPRU2394BEJFp2rG/ftxLgljk6Hsi8MOQmszS6mbUo/8Nj0LQy/9+hcTL
EUwxnBv67wo+zZ9oBy4ImrEgRyYl2Ry7VSpX1yV4wLT9bt6t8RI3v2KrOackwL9guBwsYG1tgceA
m1NQTGzl8YxYKzRDwgO2P2o4A7ICxj5obEHYTKfQpMWk17ATcZEgdb+877lU99NfPiTm2qGF8BzV
4ggoOrVPijQxEnyJGi5uR9oX+4uNampbzrdoK+s86IpgcEMLkBRjA0b54BEYuEYhDRPD1GoHHROa
qYT1AuF3bxOc8SYTttwvXhV5woApBssOm4r/U8EyHBli77oOV2NwUFkIhF09FBWfe58zjcuUm4Pp
R+edxWigmV0a5ev6GxedUdyyHOg3dv4+8G8Jj0jQrY0Y7hJH6KLY8JcwWHZEtxf71v+MkILRO4LJ
lllplH43/kDo70VTSZzRz8zlPFqdJlgOoBTNXFAVeiKgf5iGAdkUQLD0iMW8IkPgbbiXu9Uc8Ywv
XB7fJrEkVVQ1NvKkWtXkzlmNfXiwaR6HjYFRR6aruHoWQ58mpD5psCOpakwmOrv33nfG0dTQd/De
c6moevxBJBiQZ4pMFNlYkYSFpOecCtgZsoqZTTazBGwVZ+eFYqctXNBQXlK+fD1ChbdtjenqIh5x
cLOC1qdcmatXoVBUK5RLMe4dEJUX16pPCY+EzaYxRNEZrwiFdZYSObD+9hUtZreLv8fol6Aaboby
HB/O8ut1zJ/AqbQsjXHOPLmrcK3mOJoaJW8HCq0vYmTwdFc05a5ho0ANoeJ6JCMkAd6KIMNwRaLV
Yor3+nFecR6OZpN1GOyAjhLVzfyqDOteYirT9axeI9lFBXnj3Ag1m82eer/6N4pSunK7xlaC3mS7
Cqz2qyWVu39ywiySU+9/+rPSAl26GGNc24kwTXw/Y1W6YHbQ0456iLwd0ybDL4CdBHYTG9R7WNz6
qDWOhWnw15Fvb891+9PSlexs9CvpGsTS3iUhw+zNB4MLc2PICyrre2FeyTE3iLP5rAbnTTz2lfqg
Owv4g+ZzxF81Sylonc7ry9xU2dZrb9tWxo+h6yDyhP9S4q0JA7kgsDFoh+JgVZTl6U+zpbm8tLVH
MZJWDrXZ4zsBaZcoTe4r7I5aCP4RGjIY5uxreStEAzHs59gAPD2JWAumB3+rCiZFD0IpmcUU0u3Q
J/JaUtBXqoYppqNSWkENkVKIhTp1at3f8v5uN08aiCUJtfyqpUjvtZMOcNy/jFd6FDUc+WqkRTSv
ETu0iudHsaHdXyQU3tXJD0VgR9lhmuHqDQ7BqEZZZ2IAmRu2oAuFRL2B8b8HjjXjqXs/wCx91oE6
8WXJykKkjqY1ZG1y72bOtzehajE4E/MvUZdrC576pvTKkCAyia7j8BHc+QzQNDjyH6JWKWRpFsPa
dJhoaf5Vx3yLjBOzifjCPss1/Mu7YQvIABjfVcAB+hnCrckYfvJ/rzxuDEWo5KDE4X6nncWbJeZg
beXtngFrLIbMPPqvRw4fKTVla9xOp7R2KcyteAeDndlz9Xe1OzkNOV8Yr+HPiVArIh2Og2ggNrfS
vRWjl5ecLVc9C2rIzMBq2A32S3fVbXQE5cf5IH8angCp7w9CWFtD6bQegcORQYnAweGsdPY8CAvl
7n8S24rc0XAmJpAoL0rlBy/liHWzSsCcidoWExEkcO+HkxMzmDpaR0DJhRkLayHZvgnAKL+YvH0d
AipNnXoNB6++fOYbAbKMC0utZpxVdB9At4xi/mm//ai9HTtwtZn41LAQkpP98MSnneHtcCn6IiV8
imu+V69XlVgfxgJpApzC0lA3QbQiQ/c5QrNszgDyfJhEk9hXzM+YK3Alq5NFvOwyF/o6c5dvlTKe
n8m5aiW3Sdzu/OHsZZmSCkQhhI+2VrCmDANooyTHPWCKn24XbNPPQrGBcd3WlwDkTTCW59UU4TqN
kTEr4kjx2YX+ism9BB3YEUAjJr+cIinqK0zCaSYlAl09zi5iJM7viA/Mvsd3hWWAnTDXNIrCeGnR
S0/YMkFmmcRn+aVthkd1ANGteuLQ9n4fK+AaEqWV0qFp0qGm/JGXf8Hy4UMhx/pIWyphdnNnSqih
TrDrhbuitFSRrAKib0c74WwJWyueeRQ9/EQC4Z4USDQJg73o6NUXEIh7PzcO5V0BUBUkXwyLhoxK
nKOi6Y2aZmhcmib4eZEMZCN5e4x7WKZwOxTmwm/DcwAExD6cov4/J+xdNlsqdnTwHYZMOF/kPH23
xfyFq6XYqrNEqV4pu0NTvDqjbTcnfJ6g/jJQEc0cqEEfhXLI8WLp0iz3Z1KFHKdkJ+0vTbBJZme5
KDELvmlfo3bjokdi81fgpOnBFYufNJfrjG+SJIlSEgq7jCvMd091Qeg+IiwcRR25IkioQYYdhmQ/
dvwo8eLJedAf4O1GepqzAoil3YUnKr9Ki4QuWW59L0PFgmyMPVM+WHfpOMQTZ/OTVIRwtSe6Xu/E
WZNqF475DyfyEZbzU0aQsrPIVDIdi5m7HcJGdJ993bBx54aWHU7nto1QquYJXvy4soTvYfIIU0yl
2XbA7/FKw1DpHKi77urDgfDA6WUAopE6taP17hNkoe7jL8c6fT3i0nquFUa6tUY/IjAnjE9sH51c
rfzSmKiYNGJiPOIwo6f2/5XTeQ/bmyMkmtxuIk7n/yiyUGeDQRlWxvPpM0mK5Dzdw38YWVzUEx0T
KpOglsZxSe0fbcvnHbO5Crx+Y1n3QKSAL+y7RL0whbQsZWv3MIg9obBeGoaVtthg2aB5A1iK+Mi2
NBAvoL3uHyFRwKzbt4Qt8tOwQ4gYzjhaJnbnYC7hkDsPwrQYBWQuCKuxBtrmf3vny6WACYJTf/sV
r3vPZg9e8b+VDnWaM04u/1PoHAwl83lYWoNFriqZR3b57Cf0Pfz4nJqdfQIA7FxwKE6l8RUryxLC
6Ahe4y0dqPqz8/Dpca7buwdyZ9GLZxviLjdsu6C81N18blpXagC/bplTJ799Ku3hOEz9tbo3hrx6
kGeTaFJUaCvwdJsgXboeE7rcyTMberA7giKDMAxnzsF/+RjoWuDh7CLipM87wRlsorxZOqrBNdeM
EXO0wulRqjWx9m1/ByyHGr1MLA8DKEUCMuJdPWqYfn9c+dbJv1H7FRetxWvdWf7gWKixH1YguWu3
vay034HEuAY8GjKP/t267lG7OAO55X6VFkFxkCfhHfxk/II6ke0fntIks7ODYYufIZGRXKg/ytUL
7sBW2SoExibNo9mVaBn51fJQBlxOzIEPxPRfuhjVJso6U8iBN0VCfKw783kHfFeTgy2eo1rGdrCe
YJ0KIvsOg38xbqWXpezxLVN5czwkDSR6OOhHhfzklvo2XI7TCPKptiTDRsMH3pOZYqgYjout0RfX
GcUVXdrvllkOc99tU25B4Cucl7aX6o6YOoOmiIcE5BSdvmvnXtSfTD04OmRUIAmBhgf3+wLOVSEC
9CQYb59/gCjFl3zNs6sqCiAlk1WkGfhEvQBzSyV9fne9qg/7ZFUBQhTmgdM2zqGXxlPch+4Rwvcp
LLfWB2AsTrfc0eJWSPcOGvAncMlC0bsdyuQX+WscrNz8q3k+a5Ib5mPSe28/lzV7JZOUGlOp3EEJ
aOmkZmW2dhp/X4GUTFC+jI4BZWDig8QoNAnp02RFzCxpTTQ2NsyNnQwhX7DplsULKOsCkRXosQdz
gIbNqt0QFUMgt+WzlUnJ6MJxvGl9rd7m212xvk8nRZOkH0MXkgp0T5jEun8Yd4Lc1551A2PUK3LB
4tS+FYfYyrKlgrcJpzLKNxkYO3IoExeqj4dLu9jXHuPFQZO51N4hdJUjY1DvuWBpzEvnwFcpmivx
9wdO2x3gCTTJD33qiYR2k93DeBxxCIyL+5EY0F4XiOXBYpDBKRHy96WOpafczV8ox+M3QqPHzZqh
AL/P8FTckFUvOmNRnQyUYOpVOjpsfLSl8Req7+vy4h+EryL6JCMheMCzVLYembWyjMoCStv4YmdY
klFAuUnUFjfYEu2afCSmAxU0P3Zt6TgfZGdmCF/tnIbwTbrCVa/byzVwcyyG+Lhv+jv2nVJyuJko
cUhN5+tc9Irm8fqyNWBWGctgZpB+pU7U85zaf6tS8XZdBjF97aPrbbmOXYW352Z6QQFcMwcr6ClS
ZcK34FqboBrsME1GJwUV0q0RQdSGA38UxWQ+eY/asl7xdxff6iiY7wALOj2jBOkXTJjyXYmZFzaI
NkUCUtw5bgcCw0tiwYqUCJ6s8culSCmSm6grr8eQzL6HSZtRKk5tgfvW1U5wG6ZCq+yfCcr6KmkJ
+WOSUrZ2HWRgH0w14kWaTMBMRUI8cLJ417qBUkovoDg0kTKIS8zf8vL+DyrLcLtEcf/ZzKZamqcf
vWueMO/vhfcBxLwd91gJJf4/AdiLTRfhzkPpDODjnnyEpjKhbVL0u3h2ztALY2zZLtV2B9wq1I4K
grdG/YalDziKTtKZcG1E0Ip/pFPuCuWpdbWkMEzunnelYbpqbQw//sRdSsndHrsYvWagIjrQmmxr
5VZsTILLP0fHkH4BJEC8arPvzytUC1XzER8Eg0tgyNgBK9ZcS4EnyAWE098ARG//Dd/OLAQ8xK/Z
IJbgre+PzxpZ2YKdDdDzE2OfGMPhGSFAwERVcW6mA2fn4VI+DsyptLvQ/AqAWxKe/p1uHtI6OWpv
0t2qis/oAoigGYuJjpnXOORw4kafH0+tkGGkXXiHYFTZd4DpKF1YiBkdqZK7JUpsdQTEuESh7qxk
7ccAj5YrlZM9beXlIgBvkTjB044pos5s2F+oAKPgmDjzs9I4+tVUFSF3NeYMolU1j0S2i5swvn5z
QDdffphH1GavEhqaI2tmGf/NPXxMz9yIJCUgIghfLdivKVyh3fzBFekX50vK1j/Ifg9FCw+RWuhm
SsSjwyy0+Fcbrw604/3sPnSlRjwJJ1XCF+n96WOgJHAftW1ThCIN1XvLi5jKO6FMTY7UH9kZyHMU
Xhyt58THQ+B8Jyk3Xq8tmvuUv1W4+xiogkWo3LLkuy0aeXIRost1usB03icE8eEdfW2Zyr9AxE/n
tUVa4iof/eRc+L2EAfLOQ3KKEKvZtoWEQqRVwEAOlzI2uSvSAwzKNInKewTUCsoqjhx3sXQMU1CT
gnSzmNx9gp5XdC6nkQjOOcO/mh/7czNGZ4muIXFENp/7wa/rQJKcN/ujoyuVop9QuK8VCzrRxopZ
iS5GEng64tUAfkOlMbpKpshQjZJXWVHFOWF75bzqFHpKU2/RWH8Xf5i3CtN/DJzc9XC303jTqvuz
2FCjB+WrdxXhKLvWCxSfOcmmTpqYud0gFYDkSNfJxD4YoCpzUV4wIKqcFFiIZXQsKf683xXIuc9E
HZn0NdskCp9GHI08Ui9bAGAggS6PicRCgiIfNYDNCdpfyz6aZvWGojvjK0dkoE0XVxv5hrpN7jZU
ywGaMkiQn8b/hFzKDdWhjKyD0zMx/DphKsbQgGaHzar374pO4n8OALIgoF3564f96h+wiaCiM7Ch
l+bRU2PFjEZQqgAOyyCHW6XJH7vQ8Cjg4p2HFkA7f+vPVHeEIepP5kCHfgVzOfBEwrRgaTmxJj5S
CKmh/WPgl1L4opaLY2j/7hiovcHHeA4CZwD09BP6ZGVhEqc2GPloBbSDT18PXUx6vLaVf7rLDuaE
gFzv/FyAtqRjjAN23zrXrvQQfoqFz4YYWHPjoaHPHMuuQbbd/CsRheYKbhc+jaDXPXrR3vhCR65m
g/N7E01/AIr6yZZd6FiwNUgmhJF0LuvrMJMP29z2k/wWGzEjBQlxyt9gp/vXSfQ7fMZNT6QCrgTz
qpbRSaxzcd5LDVqomyd7MzqI7bonU+Xn7o6lKw4B11B24ATmIWn77mSg5dRmfFrEs+HM0g3J/F7g
FewXVakS3YXi6K36v/T+0c7nHHKLX6Hm5xFg0qfvGDKDZwzcDaEWlVXthOi1kNQMHXxgVci0pF1J
yc9lRRkT4LUEgFgv9v8fTtrYLnrV+nqA012hxlXoayc7iIvuxoXo9/VkuZRfYn1igZP3EM+dev9f
G7GXE5r+lX1f/VgaT/66TeTwEiyjt2sz+dLk/nIP9/EYzPiJnV3Ke3tl9igGrDZ4p82smxuxmD2f
mWlnKJW+P6TOitmt0I/oLd+OTlN4/I+l2Sx9cjJDc9Lb7XbRpxPmV+x80lzkXSwjS5RLAfPT5MDH
KcPqdzO7GthzrAOUKTHFOd2GX2Fje5Ir5INNnOZ2YWjPL9GtHVH6k52RkNHQsWtKDgvIvnDiJNpD
By4YxsAqPJBLCOKjn5rzbga123qLaGtHtEQEPcS/lmZVPCFkOhkPzcWHhAfqc8Nel14ioqWI7DtI
GqSqEGGZxbL3xq7js4lY677vb1EUEwmTzGFOKbC0jUJHaBjBDPmpSdsp2oc9D2jRdBkQ2rmo2euP
n3h8Q9JJIAqTWJOANZ1pZ2oxhA9TbkzhZsXNmr5/ZHJ3OXHpqhtvHqaJ57GgyUPMDNgLPgzz3Fkg
XP+yEHt/RBldNh2HX135K5JThTcp2GXQ2WNOd2A3QQMi6UKLmKjfX3cK/O1twMyvNlkW7ph3dbFa
5FC5uy6ulMcCq8ISA8KUAcEyvm1ZmqfspUc3RM52co1ODChLfrHSxSSECOb3XihdqMz/483J14KL
MZbd7cMoDS58lVmrlL3mLe1okLDcznc5EjDtvPiarIUQ5HK/hAFCFxKWq3dPgcumnsCfrWNS+Xig
grwgYBaOekZMSlGUCXy7do/2cAFKmN7evo+s92k4e/x5GJo/kY5bANmfE/bRDOBiraPKsiDBy+nS
d94VJqEOEgXh0yZTKabCSAfS/gi+A4Q1uZ6RxEXHnY6fCMRgfqJdoxYTDNU2g/Amu0ufiLGFvC0f
gyEnFGoJ8B3dS6eudi2M27cs13xbt2GAfGcWm5N/QphgB/Hw7AYeBiCGdFRv/ofhoRlQ8c2qOv91
YS1+6PFidvdY1UndervLa3nEHkeNm1C38x9Y1soKmpWsRgKy58yrd9lS7Tk9FeovP+vCjUGeNS6u
5LN8uBRoAR64tr1Um6PYEGk06E+A7rhiq3SdJr4BaTl67RFK3LnZsSvGMTyMLo1DOpd/wr+Un2Yd
bz9sh9JyCWXSDawMlO9+0kDal129i3a59p6QyJMrgqnPPLniZQmIQekzrVSY6y9lrjz3Y6H0i18i
lwC0yqP8HYfLVzoP+RpQZYe23PeiLRYVIzDpUnqgYVAWr3MzYzwm+0S4VwbBcgehEdlmR216AuvE
zGAU0vIiz0w8ezxuPikWEM9s/oxqk74m5BRE13NqCJFwosGMx/sjAJc5ywcQd4K+6MLJs/lJKRV8
yQ2dbcfOfeAR9WBA5w+9KjBAbPipgyxY3dHQC0nrLh2e5D6PNp1yZzJxWHaeO3TyEJ2l6Vff65Er
CNPA+lDZq/3t8tF2ZvFTHVJt+BNmDlu2ASGMJ6GJfTWUwotFLrKXJZ0E1R3l65yx1DFLA5aYJm9i
u/88HBfIKzgZcFJ4oLSe4qpArl+WIRZMWGOQZCRi7e3WI3Altm08oa0+7p9QZutNa3ZRbzIFYtYl
MShlhMFZSGSPydUAWAuRD29HyzA+zK4izO44+fhiuS9sjZTvNM3iDidekItcopxlJEWRgeZSouP7
TBwN0I9K5dFxV5AmmEyBGCJYqXo9ZsK/qCp8SPYr7hTJMusiJZDzzp2oqxtQEZqAkTq8+a9s7kIX
4QAytWl0cKKoIzLOTwQoC1Br1Js07bnbm6N0YBrc4bnczUh5RBmyXgLVORpjAywrR+Zz3F+6aGB+
lGmeyqjIn6GUBkWsjogBo0/8JoIiJ3wXEOR4FicD+pbnZND1EewaAqJ3wagM9J9TqAFagWTX3rAX
RvWuGgESBxgi9oE74xOZCLCsNMrILmHb5CBAqiTFG+MeXjo2QuXZnMOCvI2OaeP+K5eBp39kTEse
JLHSfhS0tj9NRJywNPI1FDKYbsMNcqx7YCNM65E61CFjPqhQLcttu5KlJj+vVg2/ss1jkcMmb1IN
IWNopbEdXp5lJA15deS7GymAqOxoVpWE2xF69DMOYbay9kJxBxR53IK5n24L//WLITC7wTD+AqJk
RW68QZ2zLI74QauCQvkS6agJ/cGOus5Li87cADOLXG0PyGVX0p5Wd2rqq7FIlN95ByiPCj6jpyqH
RXFQl8HbTsZX5Z0/OvuQzpAIaG6N9qqYtWb8L96BompwapEs7OQoZgN/c4IDp5UwrrqJ8z1LfFu9
0cT7lIsXLR6jvsD7ojDMu/jqrSa8om2CDzj6Pg21OR83mzGHFu4MiD7K7SPGR/KTxrdSZHu4+IJP
/KKnQM4C6w3oPp1rHGtMMKiXwPmFUPbiG6GBv4Up90VYnGHsRMFFNcvA8DzWl5mdau3WVzps/vnA
LethV0qfCuaCiLcH6MgYDGddQ2UXFcvaCGmeDijQOTT8boNHcpn1Oxhc1PQZbe2meDIf+B3B1VmZ
dAiHCre9WNOb7nVW6ujPhvHBeG4ZGjNuRPccqYW3nELgDjDPJmwPvBgdwVca9vih6fMSGCMoXxEh
HE7/1dmNo3LLiwyBTPEiCENcgaV34P1kM+bYXAmM5aeBX71R6XJZJxRvhn21JWr7yLAHVZuHG4Sh
sccO7l4q4xQ3fctobOXCys+WpyKqA6N8bOJlARgZPKT/EwxGUvcn29tQzzEsCBK5g000npFZuDim
pVcKD4kZ8vvsoAR+Wq4HROGgSPKI/ETYf0BWZxWXLE8zQThxRe65Hp0UDSEraN+tLSqIOpVv9No3
Xoj/HLBHmI3xR9xQKb5u3JmU7VyM/o7xNXyjuHLPqz2L58evExv52/AU6tE9LNZE0OvgrBrokVn2
S0d24nvm5xZ+2AYBU5pt2p/SNdFE/Wrex7Soj9NUzoh+PRFHWMyIMDzTAN4w/w4CeDl/rA5lhFqm
hh6uqAbFaa76m/ATr0PDplb2Azlh+/Q1Gxias+2iWtkcoKE/k7fR+6Uu4BKhDpsiG55EGY20jwc4
4Sd7th3w2CognRgooffPBAUhvPNtCJKFqAAf32Y+jCCTUyIwwcXsxtq372vyv55l1qc6qMX33eBd
Cf+lJHXLCVnntVcfezIczpQXe2rCOfeoC7mW6yq49jby4nfaR+Wr9JoucWMERMc2b0aP5+SjyKKU
KbGbjFIwMj/uf/WED68hqhgOSr+NwjIUMhQqx9nTEbx18bezgat6aBaTWBXB1/18Oy/E7MsoyCSg
rvFiYF/abHT2ZqjnON1wSZB68OA53cjJzH/B+qJCwi/KNMwUDW7muNwdJvZGCn2VViMSvIvD56CY
ur0eskueqFmBCDQZnSCwpG0aZR/29S/WPprx+wnBQxHkZhaQ8isjJf7hlcrNxLhCEjAs4vxFbu80
wH5EUO/cyg/g4Yw12tOvL7A1rFf+WbFjWDbnMquvlfxmFGdmhzPa5meTwb3ahrgePln4x1CLWfWm
Y8bkL4QhgMB6vR64UEtnCNi5CaksYdPIM2GqHVhLzKDnIkF4cUwKcE1yaM/w/5jeEw6vL1UeHyX7
84JTXbm7CA0zJIv1l0GtE2XktDPs5XhUXK5gcWkq99W9ZR3l+RZ9Cnau7Vv1Afw0w/7e0wp10hPj
pOLlvrDBMNG8D/cfNUvA962PrUfIr6naCWXtdPLNvpxc2uFjetxfE9TcwsNALjbrA835guDMm+tS
+uPOIQSZGR8sMfy3rGgCmlirXPxnO11YDfa+/BJJ9my9s4JQRZ1R1d9SqzFw1XVTlQNsK2EH/l5h
DKv/2rtLWg51+Of1/glf+9IOIqFDaixfR8On9xvpcKvWjxEhfAY1q2SmeswcLuY=
`protect end_protected
