architecture Rtl of Interpolation is
begin

end architecture;