-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tRHk8GNHzu9E8bybsEAAeqvGXWFIJdXbx9Ysyo88baTWOnLs84AlRHatg1DqRGMSAK776vgqdrFc
GllPAf1Ze7TIxSsmPbm01kyJ+KjgaiIgA9okaDYehd1NzmpOkrHHbtPF0SUncRbEDOy+797BFQeJ
cr6ZFLzFiWyTZhCSYbPLmFWo6IOCLPZPP4pQIlWNq00qAHbnIallrNKsjBdWAu+56TyzMridTqUZ
6UyQ5LsyohKR5O38/LfsJtMRxR0DF+haOQXa5n7WJMWgZ6uXTcUN4Jv/wPCCLfyYErJ6KFSiLZLq
hcv1IWJ5ozaWjhuGANT8v7+VfRRU0/d9kRdpDg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
ohZ4m0GiBJYVVwngqN+GZQutPMN9EpL8AzhICimtPs6hCpoMNCyeQfPRVF59F+qOT+Nyu9jtn0yt
MXJcH9N2vVDVGrkb0OVh7IdlqLO09PJyK+6qFsQ4Aaiss4Q2YaDNzz44QuJTD4huH2aGc2az5ntk
ySlO7Kqc6py81ZrtNU0ncxkIilvqZnPelhKQqxCJJ9NJGc/mNyW+bK98qUL+TiJ5DZjMGVM7AG0e
kU1LZuhfeRkcTefjMYV70R4pU0AMke9fzV59Ov9fiiH+m27kdGrDz2IjjcHsd4ModO5H1siKC5Kq
ZSA1PQNOpmrysDEbvSTOmheiKpqbR3pF46AuM/f5KjLORISWk6BuJLvO0ghVp/O7FbbXxotaxPsc
/vtnnvRqDyHKFPVbWqLwMGBumpWD653oW2t/2Ht/EAO25hyh+isnd20rU5RLUl9YKSVJAsU0qrcD
GN5NYU77UeBTOF7rN7AW73Q16BUhW9XbBBkspXy2i/Vr9FxTIN2p0HOS/YkHpuKDsQF2ahw2R9a1
lDDPGxnjGlt68OnZ3OtA019fdPf/MSWX9p/kKq2DjDBY2uXSQle2iMFozPfp95G19QNvcbF5XsWU
59wmBaoE3sLcbCp1P/LrixQgiI+TSOdVNANGQPwM/A/ceFY6iKRBTyGsM8vP4wWdvq+MolRHui2L
vdt5kH4FAxK7tvsk1zRIUIAZRcSzXTo44Iue8S+EuLCA6qraejzbbVd+4/QTCVmg+7Dft5iexc9g
jEu/qsh8LEGAXAmutyYLNyaqioTU2H1dh1kIvqGpzaTNqTMCbloolknKpPx6F8hpgLiO+nhyEUV8
+Kvhpn6ALCrPZBEXjQO8j/Un4q5YK84eUMibHw3+b5phLxw5JRtgw+cEAayre3aWWolFKHO8ZuvL
xj8SrYGPlPGTcrNgSKJZn5s9ONJEnAeF3i7ric9IrqGwp+a8mHYMWpV1AEPnPKIQXq05PWbRp/i+
46eUv6utOh4DtpCCbwoXI5dRyInUxXByPJS7PCPgeD7iMc6jloNC3WcIuGiY4p9pqJtVPzfUaLld
SEdu/n7YV0AvHGdUw2WFRJjCoUGyaptzds5i7JPhzxqXeADv2Yqlm0aQKHytlwa2h6dMrFWAQpHj
oyOJ9zpObV2BOkyjSuZbaSxwrR2o2qZCqByTLIjjQB/FLIXNLkgYdpTYyTdvpI30VNh2F8JnpoNh
wc1I+IMY/dumMXGNScQXlsTZA2w4q4ZcHGohaN23AQtIq9vg1hBhh5iGE6tdGgt9wMNk0RmbNc0C
ynIm0Rc5B7KzejE8GzU8gGvaESQBaGmUjqREuieOLy9NMsrc2O2JGgWm2T/ZXPps/fKh92DdWLnP
5AfPM8FqO79FYT4QOwAJPFi0cOPkxHzvp/iHshl7dlDi5oha+anVzO4Qd8TRVTsWWF31G+/Lh9gi
uRRF5QQjHky/B88GxVa6IHnStWGJGf0zzeOyagv2iz1AkWN72QUud/LF3jJH6JMri/b1PP+XUHRU
ue4+qdKZtlwbC1HoWMLcA9FW8bgAp2H/ZpyUKEBOxOEXLOqqkzd0YR8HCrcp7/3SacUoNR07AFRa
OoHbFZG4Jug5sIrgAXmd8Dw2WjHeoPiEFizJbY2cyi30l+9DiIdgixkrR2N5v84hELZTkzwqku58
Ic4g8gC89PRTQCI62MsK2SmoTjOZZPx+/pgOk4Yjk57dJb2mphvTtYcz2Hpl2TzXjVNQJG7qLRRT
CMQccm1esrINadsGQQe3OMgW7e009d+4S+BcHsE0hUH5gSvLSgT/EkHzQqXn6j1/R8ed70usTKTN
AiNwFeWZE3s2/vnO7jVcjmk3qpHXd1WTIdhejwpBOPr0YME0JFK7Kqx4SqjBc/Ds/5ev9erTd/i6
lrdjtw+YX250qe0Euuc4BLLCSgn00b33lCpArEoYfhr6tO3P33/kprmNspF1Ezud/sbMEvT23Rvv
NYb0KT1o/hZc+nsXNP4GZdXrgsT26Jnoo7RWmasSg9J5e8OSbNYxqlOqbIsu//nX4+PPjCTKWusb
ZFU76q297DEPYlt7n/htnWSw3QviZZeP8fl4qih2ToNKrJTZ6mFRMQ1Xng3KNERWKX8JK25WTGZI
7qAIoCfMlKspKTgOBDxm96Ic6LRcMwMsXWiOzhyOEZksErVTWTsk5S4clh3McEBJSLimaAwTODR0
yaaC37zbuHZ27KsWqVpCJvmanzWapye2QdIAgXJ+cVaA28GcFm1PUU04pduv5P8d6Zmorc+aueC7
60aucbvrd9RFTSdOL1Y4pXhp8LN6BZ5orju3ULnMn7r+on/TA1hdj6AQ1i8zwROr4zhk/rC2lFxQ
qQeFpNTeglxJ5Pfw+55Uw9QTmzusYJFuvfyxM2d7c4/c84I7KPTyXFC/UZ1zrY8ZI5I6ueaEavHL
u4BDQdC0c5hYpItMJDdtAa3Tl5d7paVGTy4Urm3B5z7qFnA8ezjhSRqgoOGMfQ+aC0R/H9ftyD5+
tCr3KD+eAk91RBUWYNa7wMskXrzwcK38MCRqjxYcUvGLRcNc2BUgBfdJJPOlzVOSEVGSZyzG/vy7
r2Nq4BbvHN/2ie04xNBmQe3jY8rHhvDb4gh5FuXlitfnSBscJJpwsSGbUy/ZDcA5cZhQv1c2J0PD
fCj7LsEOT93PWaF98PTktXK0dPa17kU75bSxvi6bY52C3L8NsKBBNzmiBWjcbWLnm26UGFizWxzY
8Q7U+EZbyUSrbHK4oT26S48Ejwdc4AmEHx2+frJIIF5aFbh6lNihtlmRppUTrYnQ7/rXsERuqB3L
Wsot4aVYg2Qt4kSV+znVDuiVlKF+rxcrAvu60uI6Xo0LslxDdsIbyonX10uvVZvgxmdSvopBuLkZ
IepKhpkV6W1dshFo4YOSbKQBmixisMcdFEoUu+sSorK7Uk2+q7C1b1x2wZzE0OqNEPsGBEcxGQiD
N4LvzgZk8aNUk90DZ0NmiFs6LZvMAkiJ7yl9CLgIZhEZ+s3hy7nax1RLHw8x1buTA9vk+xoQWcgJ
ZBsMnwGzogcZii/2XscutIeIxGEn92EcgarwVEjdAx3KoWJrOkmW/JcSKNnH6gnuF87Xa1b988Pt
RFvE2WEELBz95UyYaIgCc2ZHOpM05G4asX9o6bFjnUWO/BemFYCRDchOoGa/IkdhB/Nwytc+wgKl
1shfeQBKAT6mlpfwc31LV3FCJbvZNpcB3RHO+BhsYwm9NGf3dOibRyF3ciJsCP5az6SbdNqnA2au
JrxbG7y9YjhKn+03gEAaxzyP6jXxy5cL+hEw5SYeELA8c6kA4TLfZer+sASYwrkZsM+1QWI6mh3h
TTg8+1zpvZta1Ks+HotOJwghVhODlK+JDlUdFAcFQl4zUmrTDQ3oFIuYAkiod7m2YPiOwOdtfaY2
bKCVKMp8904Tv+RCvaBYukgY8LbwljaP81Pp4lV6BbiTj+a+bYXZKVNAj+NnJG8kTa0em6RlFavx
BVTK7pKClMaVB5KIsBjBjKDZ0MIz2kaJ9gnvf3vxQyxfBpiC2Vet/5SI87BdTBRcMxuZI9k6cifP
FBuPlvwq4wbH8v11LTwZTDEwf7rOrXakEkKy86/cE8d/JC6RWPAZJsCl2/OHoGLolpAEjG086uKU
YcIwA6dScPplqGDeSRRpykjcntJbclW6w1v+5KyDsPgR6LpohSFYKqPLaW+HjSKrh+xC0lP3Haut
jVAE1NqxffJqdbcf+SP3f2I3fXFT4BbsZcY78WZ2FORdOjAUxGbV0SSTvDjsU4ZYuxL4GadKgncM
Dvb0hClcWyf8fDtG50ouaiuC40leiok5907HpXPjpcWWF0P5w5K34ZOgSljQxVD9Uiz3770Gv6yf
kYpE1LdAxkBXM87H2ukhjGZKLquXpm04D5DAOOHze5yFiM4NRxFyCNVCQ7YSuBFhwZGlJilCpDnL
p2IzDjgeqtdxWCBu3u/NuUQB6LnOu8r+oqrHu3fu/oRYXSDaHww8TaW7h357x69eMy6E0pCJx/Jm
vhKxI2LYay1H4tDuZk0CsuxM9bjTFZcAaefAA9FnmOZm3mEltEJf8ny3csxgfxUuySCN5KPIFBZI
NTCnBRZoQmtSH9F2tqy928fGLtJxdaZTr1e71ZSz1QEyNFTw5KSBb/Xw+uZOfPVpIUsxmbhXQB3r
OtyFUsGDShaXXtFH9Ipg+oHSa4FK85Wl1BGpnWkD6eruEhLKxBd2Z1yNe0J9QXNNJvUXhVaCPc69
BDXTsdKW1stPVFyORhJAyMDJl/0ANhxrO9A7mvXRrXb92PXxm/vCutLtB0wLPumxdgWh6sFx2aHw
jtpys/OR/J2b+F0hz5TyFHG5mielI9x9meh1wPULqLBKYZrsx02lcea0YyeattuWMssQbPH31fNK
GHe0nmqtCZsfjUpizWMjGVeyk9P0tz4kYDfj6qFmYzJ3dY83xNeBh8l3VS9iQ8AVd5FQwRSpzFjh
Qn35fJwIowtfSU83BAeIIe/s0zNzZg3E1r/Qil6NZcTcJ/DHi+6WW/TFuVj6LstSUfqHRVzlXvb4
TVaHwBOgqBx/lxPAaHhFH0dzswdwNO4HBJ1pCxu2ND3Nlfe9YYTK5deUmZfOh9l5PO8OJQcVZ4Zz
kvnJ7x7atf+sZw8815PLYo6mqCOpu1vtBkiNNchUOF3xpAEp/ad5uJ6G8IFP4nvasmNCgCQXzXVy
XYnay8OU8lC4X3KLuA1c+H0wjODlOgHQpSValqH0sOUf0vSC4zCyhTdpRrDqPExE9CeWl8ZmBR32
RAuHyPhMkvL54ijhPuAz/lPLriWMXBfasMtVDDfdeXZEqYKfvnlUpvc69lgN6rVdLp2Mc7BcJXVv
EMsd76KPz2S/vphJAQEe1R1YHEBWdzqWds3lFemb5BOVWKdw8ia6wPu8f7ZTWxDqjfd7bX3ER7FG
DGTCRStkyFZOHt/W+MmUBtcfuAS4EmIFII/yg8Kj/nqVJA7GeKjciiQ8CZZwkNBA5W4/Ufrk37Wb
xWb4nUZB1y/ef3pe/IRTEsSFq0eMFt0iJ29wi38+efzYpOJeyEmMq3+RoWBYiUwM2zLNiUyiQ4yL
2CRQLH6iGf7iypJcPG31v2XS732b0UDW9ykYQQ6SKKUl8szT/7NRz3fMYjBEgxmNZ/O+b/azJ9Jb
49kX88AKb6+6J7z5Ie1/XB5hzr/IrsNpicwzyNgtk3ptHtYMkmg7WLR1WXZfrL9C1nKi98vFUPUk
tbqzFjvUo/vNIR3CecAC7AqgNJ6X5u/DnQ0AB8qHuvV9j654T5154eIN6ZLH/iI7Uhc8g/IqC06z
j+Rfy6VYICThL7LrwUZ0FGig5jy0wfb27b0Ekhg1Pxa4d3qniaEPUaR7q8i0zI2rTHkzKzRWudxC
0XF01GHZGgccQQXcQnsUI07QTZsIWn4HHcfJ2RPcE82RjzzmLDK8ldUt6+wtjwAztU+K0KakZwF2
6VUoWWCB+z3KBrGyPxF9FvaI3M5YtSB7D2ow6jTJs6jM+D5OiHXtqSUiGpjoT8ANvuOhkm63W1Ho
DuS3mJvqyA0QzdFAtSWAUTU/Buq9f8sHf3+pKQ1OYd98jNZOJdvaXJ9I1bWnq5tI/XGdI6XbflPF
99qZtbusjoYh1OVR1RCjH5TFf0Hq2qIM2nVsWvManhrE34hpm4029PJ+xQLbOsgL0YV7LB8ggUt8
pCDHQyCCgSxKAA/23JyuGgC2JRgigGmNE2csuGl3Z4b19O2cgHBxdPOOjwLi2CCaOvPvVH/+4CBP
pPHCYYa0imIHXTbVt676mwbF7c5AXZzQNcAIChvslcWVL68qkWr5Ty6hk+xjy2etWwhojKOPxIP1
DJNcHIbcG+izKqBEf3BJ2mniWBn8djLbSd0iNe4ufE33HYikgkVbMwS9c0OSMzJviKFwYN94nbhO
JIDGlhYNGDAnVFbahJW7v+2QyIV89BNkO2jOGfHftkEPv+SPO2COsjkli6JVl6V8toE8y59tymnY
5al+RXnY2JP0fjnY1c809SLKGLqZ8B52uvzhMBFGz1l/FnCSG2ADelgsAJ0OAhs/6QAeltJP22/7
S1zvc+mOAwBpUmPobzU5awH4VfNNEQV/qOQvZsf0f8unQE8O9uXcqyeaX4pxTxe6rHlLrJehsbJ6
6RpryT7zBK4R0H0hnN5naem8n32A48Z9x8wBcZdRv1I1jcMQ3MquWmCOcbWhSe67OEEd/TCOkDDa
9ETpiTTElv9yW67J/0WAWuf3eviRWRVELXGdGVXFOhaQAwIgKJg3OHodhjoq3e3pA9JcZ6MT8q5j
9UXbfm4eMfJVDAFrYirsoX1Fz8qtcJ0A4f6ulkrUwMf7JXEZZ97GheR0ux6hBCvuhaJsB1ZSP10q
AvP3GMDUTrfPwFQYoeSzOjpbA8BP0UnED09lyMSKlBiBpZIf7/XYvn5GyqoMxZcrayJwpASCqNI9
yz2Q+xhl0PG80AqLpk2BSPi2/l5I7fIgToIBgQR28QbJ2LIllDbpI0WlVcFZOBkHVPc5NdaW3P/g
oNjDUH8PhaodaYyNjok3o6dqdmLldLOCOtZRf13r8BjHktM/HwdmRCtv456dsxowi/Gug2PQ4LE4
UF8ftGCfO6U/8IDoe51j3aQvJ+shxn0Mu4yoPLImXNiMHcw3uzs5SEgOJ8IXU554aiA8S3SQZ/E+
FjOhiN6AkcdhJCNQ+p+f0FZ32N2pF6odmAQygOsAI99SJPIqIxbrY3uHwgyULUmkBL5a/QeLqr3L
yS4+QMekB4+cKRsI/JkWTcycyk8Fs8P1VHuUkb8VEwDxtzmqh9JWkvww/GV2qE3Lx6HmezXAFezA
dUg2ZNaMg93SEdBcq/5TLHIuuPWzF/QIfhrDzQoMIJYQDuQIgm7R4FmkoAGfZ53tiLpR/doJNJf3
R2O0dPbLuINQICMGKonnHhQ+rLW/mD+lTaTr3Udx8s/2Owf446bOzB41HoilDbV7TMhBLH69+lWp
AsnHO1uGV43YwmannlpOzetjEZ0LsxLif1V84VpJ3vT5DbNj
`protect end_protected
