��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�"���6�$�rܕaic�q�Z�ψ3D ��}�O��7��ջz�\�:�����5n�#l���%�cu���%y��y=����NU����!x�GY�9���U=����2�:6�xՌ�4o��]��i���оU+_-B��M��J���q�J��ua�F�X���E@���(�s]�{����s����(>���0M	Hﯨ�$HyÞ(��d�iV!QV���:��7�,a�
��3L�w^��W��9��1�Q1n�|�*� ��8�g����"+�esP���o�CH�&�џ�z������u��:p�=�?YP��5��^�[��"��p$LN:�dw{Tȑ& ܤ�:3�gɆ�ºU���M��"�	�9]��2:)
�z�����~���(���#S��0�صm*P�Όj.Ȝ��.1m�������9~��W`As��mW���@�շT;*��^VQ��$4��g?)��&Q��i,�'���ꮎ��Tk��#><����7�6`���>k���L��Ϯ�G��X-;�>��R�C?Q?�~��{�M�;Ξ�4�f6S�]C_�Ѧ t!da � d�A��d$�.���r ��'���˦����X��q'�19p�:���k!����۪f�DLc�Pj��Zzh�x�975�.o�|�������"}�׌��>g)�w	�и�b�h�R��?[C�B�����n��b�Ö�&]q���V<l��I#�ϸ�&�m��W�ٜ�1V�9�4���,���y�jN���ۜ�ؼ͢��������y�@�uN��^�`�Q:�X�����S�
$����0LE?K��<����h1
*�ܸ����%�@.q6r��	��ð`&�#r�q�s^�X�P�t��� {
�7��5"� �Ʃ޳B\�5XB� .���K	���Ǫ���|B�S݊�394:F�S�����$����DQ�aHqRY$����"�{s;��r�J�$~�%��l����Z�L�Sx���T�Q)a|�.�x0���dWO����������,;��ν�y+=t!?s���N�"z���p+��n�9���Բ��_���ٸ��l`�ޠA455�V$��qx���J��Ч�DX�T��9�L��YIHZO��#�L�B��Z[�:�GϬ>Ȫ|��;��J����16�PM^��x_�Z��q�>.��3��*��!�M	P;==Vh����=�j?���B�R�dK��̕,��#�.4iu�/�����흢�w�H/��ߟ���R�\����]�Ј���v�L���7y���-�,-@W��{,��G~j|]n���C�Xm�46�Z���;P�1�_j�i�7�����h��������>
\��x�D���%k��Į[�a;U��YH�Q�D��@����/�yʈoR(�t�Y˱Ym�s�_�E��-�!(�R)�p	�.=���?�0X��-0�'h�⣇	��
Y"�]a�o.���Gj����^ԒC�E�L�ʯ�r<���Ӻ�Fb)]S$�[W���lRK5HrP�PW"6�E��M�Zs��$�,�bS�����q������S�zCNuMV?�Ӡ��
��+�"���e�[E�5N��y�5�������k��/��/'�l� ���{]�Ro�H��)OHO�o��g��)>�86X6��ۨ��J�4t�V^�z��U_f�A�D:�ļP$y����(�"��ѹ:#`���ߢG���T~�R1��L	4̼�������	�ֱ�=�ϖFS�0O�#%}X8��S��
Gر7*q��eʲ�%�)��<8��x8��< �a�WAh�>Ԉ��{��1���l�Ȃ>�X��Zy\�w6?0���@�9o�?�sس"�j�1�Q6qPܫa=6�4~�_�tj���u��~3+{bMh�rV�sJ���\����^��T���[�����m�z�E3^��" ����6D��9.:Y���8������e�I�tq�"�Ƽ��`����9@�)gYػ2	����%v��,�L��sO$��m�s���`?Pf���Np�G�?�*���O�G����t�;�e��w8������qQ4�	�(�mlJ(%˪�W {x���L��s����pռS���:)���l���Ic��@��MavB�
R]��S$�e�������-K�6��{��Ma]k����A��L���ݏ�up$7����	4���?ruO�}�@'@$�`�̥�^�D�d��U� H�$KSX��6X?��� �O�j:�o��-��.vUw�=�}J���ZB���þ�I,_���ӵw����nCy��3y7�&��v!O��YgP�V�2���oG'صE?Q�5�S��S�V��K�8�� �3L-�V=g����AFݢ�]'��Rv��@�DM�.'�/N\�#���LO�������P[�~�^Ӛd��IR;���V���1vw!���G���y�[zв�B���=Վ�ᶗ7d<97I���A
�r{V���v�u���5���u;�pv&�]%둏=h�H��pFyP&꼜�Di�ZaR�38�Ү��+am�Q隈��ƒ��쨙��7�yأgA�<	��f��B#�~E��	��I�\P��|$���m�AV�>E8K����ݲ�0��~�l�Ő�Ep���b��첁@=b�dc����RN_1���� ����w�^t��pz%���+��O	�n�6�h���f-�犍��xt��H�-}���*j<����\������Q�+�&[4�܌v
�M�pUz�6_�hW!����FT�P �[>��֩(8ho���!q[Ø����Dg;�8O�dQ�B�س�f��{�{d�o�f��e�,�j�C�\��je^{_}�����"Q԰�Y=Z*/��'ǲT;�K���,���3��C=̶�����H�����*�OF�ˤڛ>���ZԈ�Z8��E{an��T�a�nE��n����*M�A�:�V���%NԨ�v���"�7?�i�/���p^��y�ޢ8�c��M�1����iT���� 9߼ω�ɠĬ����'� FY��d�I�hؖ�����ދ!�;"���օ�}F4Y����0�!ў����)�ׄ�7����K��G�V����~�OZ7���3���	k���[��Ǆ ��s#WNs�\ȡ���<� �[�
79�9��L?='��xdz�2�o��6�cx��%yz0򡖇i!����y<pyc��H�6J��X��.)5TMbf��k���5��&�t�R��C������#��p�o��ⷬ4Z��Ñu�����XYb~�c��U��@f�
*��+y7��`�`w��p��oD8�J�J�� Q{H_��iٚ�fE����K�J�'aND|?�]�0{�Ȃ$3�í�n��5k��2��Y����*D�IGxS9	.��e��|g�?N�ܴ�3�ֈ�z�ذ���1��k�z=v��m#�[S�o��BC�!A�����	�E4U~|5��,ϙ���d�	?W$�z\2�����
E��������(e����ЍCHv�ݓ59�����vP>���H�ܩn����npf��N�p�"E΁ S���fp�6��}ɹ����"��o{�b�x�MF�Y������L�v!O���!
��^w&��[XfC�j;�u��'4A�_�|�� �ٯ��i�:��#�\E� ب��~׹��=�����K����K�4:9��6S����ܷ$�t�B���=<�3�9=et�Ҿ&r��
[�@k���ܥ�G:qF����ׯ��'+����5��.��1L�,w$=��wƆ%/s�?��_�f5i�'o<��C̾f��c�{�����V���E�hp�@S+��Sm~\�>��)��Κn�o:��͞9aW��Z���3�J=��@�U�S�w��R��|ؑ���C��W��rX)Ɖg�5[C ��r����L��QǏ��a��B���S���w7@B�aru����Ǡ�xt��%�:C��&mCf<��7��O��˼���az�y�c!��z&��p��b���$�3�8y1%���v�v���>1mm�Suj��om������i�cמ�]���*ĝHȧ�Oڒt
����8�)k��&�i�z����A�$�mĽQI%�Ԡ����C