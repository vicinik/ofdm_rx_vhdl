��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��Pޕi�2�Խ�cu�̿�����?h�BH�wd��-��ʴ:9o��:�u�զ{rC�wT/ ���f��zG�ܞ:����칋i\c� �*�褒>m��u�P ]Hq�@i�
DF"4�3iH�b�xvjI�%[ln�-ey1�d�!�j���(֧L��Ō<+^����]ӏ�f�nA޲C?v[��@C�S%���=(���Нl�e�Iڻ�3&ӦfB��G�����|�Ԡ�w��) 6���W7@Bn���E&5'Vo�@:"�ЅF�җ?�-Qk�t���]�����DK�d-*��5�`]���D���Z][b6�ˇЪ��3&Ԥg�j�t�B�-6W��S	�VAV,o�]�勵f��j�R`OY'�_�Ђ��i��R|�����Hp>�<�Qh��'	 ŀ1�혫�{[�ȡ0�@[�JR�;vŏ�`��P��f\hO=��;۝�v�A�1�:�p�2�U���tC��H���Q4LIn�b���a0�"��<R���6!7� #:E��r|E���!���ժ�=y�y�,�>$2�)�"�G/�A��4�.jszi�e�n�������5�-TL��u��j3;[g&�̍����Pt���'o�bьA�]� �(�65W��\
��R�p��o��P���*�J�S7�g\�&���*D���7}�d+�}�M���\�ve"xv���BgY�	�J�[ʽ1�F�G��H�[^�����)��B e�0�x͏��&,�E�ˬi����\q�͘�/�jP)���t�*+kϸ�}^���#�NL���AfX'JG!���ޯT�G����>e�o���c� 1=7!����Vљ�S�Qi3�]�����d�I �ds  ���#�:�P�*��wEU��h��Qr3�Gp�D	��g�Z�x��U��S�$��,&p�f�<�=�D�֐�5��*T�b&���8s�F/�˔[bf�<�z��t��\��V�=x��fP2k�"��p��	�y�';�� ��ڄ~�,�[:5"����G�}�����osNa" Ki��3g�#�/SA����	�4X[�Ph���~OX�F��yeA=��;w�9�Bk#
��o���.3�WY�qMh�������`#Ub�����v
/������Ͻ���a�Д��?�=�^_�3'�L|^5�Z�H�@��ޞ���Ȁn���us�?��S$�{� r�]���P����P�
6��7�礆���\�D�Wg�]\q|�P8��+{��:S�s#%Y��ṋF��v��|�$d��1Y�	ouE�d�n
�k�k�W�Q�"3a�n��vyܜ��r� �j��������"K]�X�Y/��/��\I�a���T�!֯��U8C ��U�@J-QN�}��e��Ce�Y6'ZPr���{D���_��i'-�]���QFW	t����5�z^�V^E�^�]���fl�V�w�χ�C�!����R��V��._�Ѱ��m�v�`x�|��L�������;n�x������IOO:��)R3g��1wc�bts�z�E������Ѽ��+G� \�v��C� J��{�n��ze������ ��u��4S��<�v~^Nq�;�I׫	�?�)�	�	�<���.��R���BUq	2LU����X�]�A�Q힖�)���0��`<�?E����I�{�����Ƌ؝���fk=䠒��gmz��Y��L� ��O�6w���.].bmL%�R� �R�Җ%q��v�a�e�_c�Ɣ{d���g��U����q��
YQ��n�K����RM܅6i�r�~���9hPp��,n�j��kh�.b�� X���S��$e�W\L3��EH0����}��o7�.Nøq��7o�8VN�\�V�M?HJ��Y���@`l���S�D�� ���SFQJ�oi3�7al�R� �0��!f����	^Ѭ�{IK�mQ��Fk?۹�z��ص��8��;�Ǚe�U�\��nYUB�N�;�X��3���]�?:d���j��%F,E��DI��j[�ԡ�3g7n'� 3'�U�PWZ<�R3�um���W��:O��6}��ķP�U�#�w'��@V@c�b.��E(��u��8�j~������߳�M����	�ɷa5e�<��Cq�����ׂ�_���U��پ؃C���f��!�ij�X�c�I�g�)L�%>ʈ���(�@��ֵ����߇v�#�]��z���׈L~�@��tȏ9c n�l�	�y�M��~�" ^�#���C|�\�p�w�՛/�`n����Q�O�%ȿ'+�:����\�V�W�n�:�Q�&����H�p���r6�l�	n�A�Y`<�C���fڄl�z�DA��*����1z�O�1R��P��H�'� �0J	}��-)л�;:�1_.WL�)M �Φ��'(Q+D���}�A�DS�&��A�C��Ҏ�7���gM��K�#̚5Z�R����+�P,�S:W��cP j���'X18�q�9ov὜U)�����	�ŜV�����+��x�S��0��S�tj�$�C�u/��t8��&I˰Қo}�]�5lH{�W)KՄ)�_�pei��Pj���[����sf+�ޝ�͡M#a�*c ��#�
��Bt���j��^@$�w�G�{.�9�n�5~]��HE% �adpa�rJ�P����_2�6�^���+���]��	�����^�ڝ8d�X�ʬN�V'�
i��gYQ"蚘umL��Ai]�38��m/Ũa��E��a�{Q�iW4�]:�vZ$͖�"�X��槔7����������
������v�~�	�1#�����\�bߞ���ڲ�A���Na�w�_b'�X��_��3���e`PH�e9�\���A b1���sx+F��+?l��W�(E,3Œϕ�-	�'E@n-�X5:,��Q����˂v��j�}���x�~�٤J�+[~E����'��1�WK8�e�	wk�9k�W���:s�/ũ_n@��=�}���8L�ܭ�J�r�����>�K��@�Ĩw�o�^dx��ݵ����aR
��@��ҋ��q��-��ָ;��6�G*p�e�y�>gE�ð8��{ ٲ� 4cL5I��9L4���l>E���{H��f��'4�>��n:�^0�W�9�IG<M�hv�	�N��F9�4 �IX��9��K�o�ݡ���Ë:	��^������/:�(H)�C��Uр�DGW�����`"����华^Fqx��ĘYY�y
�L��O�@k�G��C�#��0��A��UzQ��L�VDd�9?�+_+���%����)��=��h�$.5��(���C��%HN�rk��(ّ:��*\��;<;��>ld����53���!��YT��4.}�����e��|�<�
�G���S���g7��R�h����ମ#�/}�]�G�\Y�5�<q�Ժ�Rv�~��zt*�i�וapl��Q�G�TT��T'lȱ��QcCoI��u�iN_�V�������7��yhWN����D�{Lwcrd�ų�F��qk��5�[�Q)�s��X�o[�,O�DH�㑩�  ����&?Y�����)�ҙ�E>���$�����֥4%��	/r|/��Q4Q�f:p���[	�=��J�u�L���.<�4������ E@o�% �="�"�l��+X�\�4�()���cU���^Fe�o{I�N���D�u���V�����zߴ�����,��1t����а���,_���Ml�E���f�0�۴��^0!�F�"����˾���!S��cA2=�ECK�'2
�Gk��(�K�������y�5R����Z�`�NŊ�6A�
�@��:����J�
� u�P����0�1�)�z[$W�E�?g8�Ne5,�@��
��2����Pz4�2�"� ��uo�}�agx�7'h�q4�����(Ɣ|�&��O���D��;mO�H���Ff3��1]�� ��J��O�sF�G$WK�ػ�'�J*8��`q��<�3��k�Xj�:
gNp�@47��0��[�7��Y﮸�%%S*��T�G^4��k'+�!���6c0�y{!��a\/T��V)��s*i��3���,�,�!&0/��^�O�����]ݗ2� �*8GL-5J�����u�����yz%�W�x/���=�E���sW��e�T./5�QT���ӫ�����<���qu�G�,M���$eɒ8ҜH(��$�:��
�׏�������J�4
bS�S���v#�3A�fT��Q��3 \�����u#~a�2���?����txV�o��Ե��s��`j���ߖ���(��:�~���y_G�t��c�k���T�����k[c�g�|�?���IP.J(�/%�����4v�Թa>:c���'$hm\���<�6�q��ev�Jn�b`�hS9CK�|�Du�F��sH�!�WS�g�n.K��*P��`��E�4�h$��w �l���� [������2�T���]O��o�������M#������*E@������DQX+ W#UDD�Ɇ�OB_ӬQ�B Q�#�j�J���-����w'��a\����h�ǖ�$i,D���+c��;��O�����h$kYpkZΈ�=L�vA���#�E뀭d�#��ݥc�}zkT�Ώ5�#�L��R�\���/r�ļ�>i���5(&/�'hoV~]�_�l���1Ѝ|��1�����yX�A��?>��5��#�4|O��BK�[��GƉ>��qk/�]�H��_i�E[A�g�_���RF4*��40������'���/�+]�/��2		V��fU�C��r�5�� �T�&� ����a����bȕh������"b��\L�������wM!��=��Oz���9Z��.I:����k&!�Q���L�1�+A���x�`o���+�~[�;˭V���kXlH#���?�[�r���TA�$qo�p���Ӛ�� ^����ͦ���I��a��Y�-j�l���!�l��������7_��"hm�7��b/�@�8?L���'˦�;G�9s�\�"[�P��Qe��st��ϯ�H�i{�:Y�Y�N�@���z%�mD�#T�3��"h�nŪ�UIXj�����v�(�\��[({�����