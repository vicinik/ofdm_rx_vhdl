-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ndoZva68Fq+9IokyR/QT3LAIxTEedRkrN//4DEES8b8QKox7lSKk5zR1jZQ4J7qgot0pQ+YCoebc
8FnYaVdJEJgQc/++dRPeyeftXKFMh7mdpma0XkZhIwtu1RBGzPxSKYs9pE/cqLtpi0BiwE/NEtSF
7EXlpS1+vKHdLRDjB9WiKYXKX5/k67NrCxCEa3Pc1Ub6YMcpWrmv+6mllbIfJjfk7XV+ZoOZodEo
4koQFIk3ihcn94QmmEEGOLTJ0GNdiUBD5P9c8wu6SnrNnuQkhjXfbglCi498shTtG4M1y/pXnP2h
fj2nsYjoevCi05j86X8J92xBC03ZjZL8RCt/7A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18160)
`protect data_block
08c3Ob6jGk1nC1cg6355esSvMA7OJfSAP37MESxny9NQb0oeCwAEKpYhqqZA/eYq9tDY82aGAprw
/Q+nWJsag/NT/zfwUlEBlh0P+OBbjjHPXRiOqKVNYJX7H8yqwYUrzceK6+5FnUMYNLiNU4Xw4n1K
fxcj/plNnSRON880kaDuvpUiJhFmwnwHvPuOJdj5qBWJWCZXA6oKhX0uUWnH5URqVuqeD09xwe8p
fFpxjgW9xAz8UPdqE6e04oT6MWrgNrF3zOraAZphl9GlCO2i09Gp4M4CFANosJESQd32YreRw9ig
RXUlL9MLJ7pPzM5+rSQO1fAuJjX2rzKZdCAVFRMQMbcw+n5R70keCf9w0RctlwSBPJ8vUTjd8fUx
QSsArcZ2MHUBc8Qsz6oaMqz602P4f8h0nxa7lRIhVDX5vi+Vu+H0aUOF3lz9tNqXLPwOLY5FSnNA
Hxtcbn8EY4ADMcYJ/e7ga+w9mTUz/At3HD5nZOALhZYN2paE3idYnbxpRhMLjX6xp1ig7dGv2/Hw
Yf02UqE16vJlTSNNbh4qMkGcXlHGFBGfM/WQHD32B0yoqo+HjBliNpgebjHaUtGgzyp+5R5caj3q
tgtHgDbQ9XoVbByYTLOaBmK1dGD2+xE18uBOvVj77VIy0Az50KpWJ0WbgAum1Lhtp+BFLgpz3APe
QeGH/uqIqNRN+z5PWgqWRwhYc2MhSdTFHp22oxF2EykgXsBDI/Pc0Q2F6bgsFw37S91oOr1cHiSg
tUyattKxhssdj6HZOmn6K5LDd3sW+KfHTruKEWXwf6wwchenkpJdd3Bti7iNi5MVt8BgRqhsiqda
CzxougWQSz3ccShrWlWx337R0F/AFN+Klc6wgVPaRE4TJ+cVIuUhxdoptRmxUiNrm9O547RdGpU+
ENLvBs2raz3XTT1lsB41mlOxDlN2Yupe5+7F+F5Dq979CZrg2IMBBbbF525yprd1iip3W0iU5f+e
/kjJycdKsCDXuKNx3Ngm3H8h5vEbOVsTRNnv8b2mHtufMZ8PPFd+4h52wD7coHxEgqIzeurs8vt2
Ab3jShBuUGduCPK53di2K41I4pp4Cm2e1dpKCrK1pVXDY5qXzCkgQOaFq3KqU1mYFFE5B0lllMM9
IKA6GeTuJhyrCxMfXkZk12lRVLiaAUyVcpstuDl1heuWplGCGllF1pgK9whWfexItVtfwWlrB6rR
snF0g1fGzJUwq4QOUV0LUvnsPJ7HvyMLcj1qHYqiUbGfOWU6BNTIwuF6HU0kWdEJ1fyl3CTVaCyB
g/spCWOqeqzM7ejcBw8gsf5Nz/+2VqsMRBBMk228ojC9SXMJ392FZg6EB7qzY6+LfC4lfErQCTBH
gSs1wuOYafe1LVzlMMPh7EK0+qKIvL/nb2lS7CY+0gkN4mjw5t+lV/15D4o3dWsX860tO/DiVDzQ
iJD3J7nIJmzN6juVls3VqGPvkeimmOjXdWPVnmme7VdaR3uO/bTdgOq17zHtnxHbWUGnGRHU/ZvR
HbxwmbAJWK1V9MA32l2MG0zbP6Dg2Adr7cD2/wvw2BOsV0SnzAsTMCzZqcyjEaHnvMNwcrLCGyHt
IjNP402cHuAKr1TMxu2zxNeRNaDtkm7hyODBVvfUehHLMQWqhBT/Y9zD5OSuMx10raOwcl3j6N+l
bP7cQhse0nIVSDJ51GqKOn1cPih6p8UnC2/1CWsXaBn2hv8jMCK6Oh39bd5QUsyyPNH8PNABMFZP
3H+Mrki8z5rjm9dwxKfHyK+MQAaSu2nYtc/aDWUaA3Y+lJLNRWH4SnBblWvlpznnLJnWnaQqLPT+
TTw+ZmwyW1fZMjjxGuIC5zbibbw/jFb3lrXM62KSBc4QhRCKCsA6qtihXsfEseZUhjVkQJ649uxr
TBGZF5JNFenuu/CxA60TTeW4GOKUnh1X50IHKYSnpwOZp6MKcWcpVMAGCKEFKbJMBnm0TkTmtEC2
95anC2kZRKCVFE7rlkWM8S7Q1PHyLjkL053z6zvWmPA0ynnvs0/9MenvZzXM1SDF2C4XO17Rus/B
tBOAF0DpViiia42zgVWmOXukofM7abYlWGvMVMKHYSVfCcLQV/2vRrW4yuQK/uhG5ZurTe98nrrd
Nnve7G4caAYZ2CRIpv4qLEU/G+8CUAA8shK7lwmz9Aof0nY8azLoMEm5N0k4SGAB5TYoNJ5KihoL
AVGdybcaG9qcVmDK0HY0jlM7LbDFnYL4j2ZK4NKIHLoZpqTHd3cf2F9JL650TwrrD5GucmPOZ5oR
iug4xumvteVI5XilEAwPv9fv3R8/nsZmBZY2VWOuKFB800wQ+l47kHq4G6ejZOeBWxuDZmo3J7aK
0+evz1HtNLunq1SfWbcKXEjo47Xj6fjTpmkJH/7gMEXnm0gkaEKoT/KxxtNqICqeHsR45GzXBiV7
I5EAz2je/CZMHD1vsN4nwEpS+ckj01fcbtaP19E0HYhUeo1a1+hzHAJv4F7rTc0PYavngNlChvqa
cKS1ImOuCCfrSddd65tRfXLkD7lTcElNU0fjq2l5N4T1+h0oSmaSJnwGZyZgV0bEcGNPz5p5ep1+
e1PCOFuWJBEBgcLrcDo0aGOIe0hCtz4oXTs8fkeh5eE0QGyZ4kXMlz+EUd16KKTpHCsC2svicLLb
q/HByf26ydD2sMlbLqoxloCSiqqxGbz/C67kJjwk6NvUYJj1X66YEU7fj4Q/seEPwyi0EM8umaVZ
7g4rjPj9b5zQ6aYkNxNOxr7FqZmVtQxOPE3IzB2YY2CE/dbAiPVNeZy6s/IOzcwxoJMdWfVVPzM/
gvE+FhqWD3FeeiGZ+wPdxbUX2VidsnHYqwoCDL1pIRIEfvzLAExcHUAFhsZpbT4vwZwKyTesAfFV
+59TxBVCXznk+mkbpGt5Z1NptZbgfsk5ApLW7HYFwgBV331tfKy+JPF4AF6uEiAVhZsfwTHJggq2
cPp0Fn8xcJaQNOP50J+WLQLR1kUrtuAa/qtrAw/zKKAhnTCp8tDqO55VOq9zxgvXVsUjv545fkDO
WUKFdKcANDJSnYOjYysLOxd6XSIWL9wtix5Pieko+Y3jlklaze1wryWkAXWWgP/bdY64ujg5NP0F
gnCj5gQ8Wj6XiuMVo93BIL/DvJRPwIr4X71a4/0eiwqu4Xpx4QKHo0r9GZvHwQ9lNMUJ85o8f+Ms
ODdwf6EVVUUnqLoLDXsF2b8+o2PmSMieDap41FW+mMfxgJ5yWMvx+zZ3fBrvTP1yysReWfQAN7pM
uNrwgsashqVLrRGV/mYza4C5v1+7nKcaA2p/pLaRZKEkKf4mpqN4AUGvu9XTqFUWQ1HkGVVmUWdf
9KisDGvqhxJ3O+4C3d/IsGfLnPTXvqXqZ2tKIQ/A8hbG01l89z9ekUoJF1OCXgelH6Dl4RQ73wsf
sImPXI63cNyyTqFnZTH9iD3SE/fp/GyM0CcWJwR1+kY4O7ma1UT6Z+iEhUA0yaHbvQ/zPOkp8FyD
xJ6j38ekG/VDefj2hTKQArJbelmwHToMbuaaZVegDzgVmFeDbaW6HFUnXOm45j3CphGBoNTp5BTC
ON8RpDXQscnFylSW5z3PzBCIfE++xCaa64BLqUOxF14ArRcgLst81pk0rs6G3ugyHHIO6gxme53e
ztxO2duv6o8/NWxmKhvXhzsA3GLDDD+OqFj6woQRxksw/32jY4L7T3pdf3TH5XpQ8imx2l3Lkb6e
wHaSRkVFA8AlZz22aplkY/czRpcHVUPw8TpbPX8QsPEw6o10PSUFB4PMnRtV2vmhlZRyDr3RanQq
t/HlgCTT2tvl3iGaXE25Nkhz4oE3bOVrU/AqKF+4fZEbiq26kJHTcf0/pdmD57xwy5UX4SUtJqCV
obXoCfwEtrEl3/YFa4WDYYKnrp4ECTmy1+vu+b2Cmq574hXfFXB+dLWMMemHazQaxD828E/eASrj
ZxpUs5DMsxRKjwO8rX+LvMDarAEeTUWCM2Y5Y8VH06gaDtJaGxoi/2CfUBaMYp5PBASxOkQ/hQR/
HEqYfp0krE+IxQN4u14KjywgG7dnQLtjfhgkrI16+e2U1paBofXsrC79Zj4J7XS7t+GXXPgLGCux
GgUDIn+piDn7d3gCOuWk/XjSUvcQsOc7A3J6nCHdhUP90mqbZx0/NdCqBNWDXAjDNyTEefMdHXxM
d8i+xbiVkFbtOEvPui9qEGJnBWPjsCezPsZN6K7PN8R3T9vQXity0Evn6wwCjB+l52FijcxnePiM
mak1w0Z9AQ3zYTsCnKeXa1M3EzjsfL1iPw7qPpNvhoM6IEHGM3XAPHQHmQBLKP/bEinDnGwhmocH
tocUp8krmczB4YinyE2kjnPTT36sr0kJgWN/pNr1hN2zKuoOaHuoNHl0haKwb8jxHvEl4Tvv+Jqp
JI4Z/rLcCaoZSLSiQehkvwy781WMNuPaRyrszZ1Fh+jHux8crtryEjCbobcctuaftTVzGh7JnTQd
7V/7agi7T4Qbki/NbzcL9TPlP16Z01b0qnZjp9T+bjhwTW/bJNxDilgMHDp87lBPEY/+kRFqa5l/
XuBmWVjMCj4nwRfHx+QqYkFIJPFOFl9FHTHJvfBXsUcuHeGM+6zb7aTslMrS/3O0dhCUSRwhCaDi
A0IRTSoA1/b+WbQqvB+ZL8g9yo3Nl75u8Lj9JJpB6ct4SCf1zv4sKHCBEnjU36WERg0NjGbtd2ge
QY2dAoQaaPysmr4t1ukcUePr8ZxaUNpSmfTyAqc3aVP2d9B7z0nwA8Hx7ueMVZPFDAXqbM+ZnzQi
gMruohLfwzBXmNyR4jCXDcehRXy22fE2RbeU1QYWN5DZEo6JoESD8oi/WjGSpMRLjmhdFPxp5DWx
5ahtXo1SWNnQEBtPs5H/QtIO89rC9NJPn8pIXqNsfX06g4xUWOvTgXqYzoz7r7ykJ1oLvJwxT8hC
Gj5BAoQlUab7v7Wqqk7e52GyzIczaJV/JIgLpghbfyJ5bGNChh4Ez7oiujAUrsCCLGMivHxFBzKW
921CRkRmaKiv0p1oENnEWvMkKIavsol4roI/kf4hfYzhQonRw5bBlx+4WVuoupU8hjrMKue03Tai
qgSuh9jiEQQWToQ7awto48QvOczk6a/Y5AzNRc0yNdtNVCxiZxmkuUMu2USlivqBa1NiNXsRGpFm
Y+Fwj3t2tIBKgZ50afwtDG0sBPWgMY+Dx4MuRkOiiCh9mGh6WEFvy7UYZks4cK21XZIg+CGGwNWp
aZFjoTyI3h64W+qlgSjWVGN8XRMmw5lB7BcNDH0kKOK/TWn49IkXQzzeWPdZPbIGVpo4SovTsHnQ
5hnjr+QLzBW20b6pJAzoqWzXA2QIDBJhAMsLg7VSUG76WwqLGHD8R60mfuhb+41rwoti5dqn0Fel
Zyw5n7Ocls2aSH836S6hEJm9Mb79ksVQKtTaFbLs5mvKVnJ0pXMuVzWRtdOmrO4elxCWcSKPtuZ7
dFbbmQJtRVhKR21/RGYSeGO831a8ikp14IQaB8ryAI/KH0oAzfyLQQ2/37wp7zxzfuNALZ7ksRS8
UUe2GVigD59wZmebSdKoKKOdpDHdtCs5i14v+8E4KfwUnBt6z2j8s4BooVHwe53s4EJC8FrHb/dj
yf66fa80WmNnqyX+EroDifSqO5e8e7aOyDtj3591/IRzUxgT6YuibyjVja21NFvyLAggk76fYAPg
uK/tzG1vtWQ/iYbqysNUaq+cIO52vbP2Aab1IQ6gyJeuy1IB/vp8gL1Z0NqYLUoRW4rAej5oRmEZ
XymOFYPnGgGiiq1KdbtjawVd3oGLVWRNTvUBv258D0L0YKTuTUDW7JE152pMm4lTZaeqZ7sOBysn
kSFd4OnqFqbBA3jSgqL5pSSh+OKTd9yVtK4g7D7lrWO33Ex/58mZKrUP/PBDjUZm5hB3YByCd3qR
n1ZjDaME6ek1cgfiB1JjchnEOJmmaSQaJax+qGJ40MSvkH7E+GAlZMOmc6RZ5ovD3YdeD7y8WeD3
WxUnUwML3snHM8TBTAZlPGVGDgCmgb49GNfuyV6wl0H4u+xSCmQMbnZ5DELntyNSvssN7L0ZYRUO
GPqQt2v7tdG1U7zXXKEFVoGsiqEHV6taoW5//76OmDpWKu9os8CCxsUrzUNtcXQhH+Y3bhtg78CU
0DPJvlT6tHJVIj3mPNsToORH1NIYEmtZuSSheU3kzfivl9DsFBsCitPpukasXYRjJA/nYQvl85BE
Nfb4fRXMy+SKSlJhziW92LcuiWN3vKj3GHKgcxjpXqBbbLCFTWpRAuc0nE4dSFWOsKpk+6xRGKu6
Ownwo/20bBZe2opp2IzIpkmkZ4Xl/zwuZVY0+4hgM7QYuzACpDZUXKViJ9RU/M4xtjf2P6QcvYnU
b+TGwlDXVlADUmkWLU8ni4EUdm4WlfxydACGH3UpzepYBwZYjHMowzW/Hvy64PtdpWgX2hxVyKzz
BygJUXeY2VzyeP6Y2nXoDZvGTq35jnZRIIuTuniNr9nOVhnTWpy/jQ7BknlSq46zUYNWIdesMFWp
iSKbOMg2TYQ/fexHn9fHSPqQJ4ZI3ENE1rXRHaDZHmMtxRysmLv33GKEkoI+GqmiicsMp5og3N+L
+CwfAYFaQt+LBQdS3IpJhOoxjH8/qutz3BqQSa4hQ9UQsmopgvkvZxQ5kIO0iCDBKxdSpc229nRW
8Qi+ZWHHjh8qq+jFFAeEo6jSTQ4ZupTuMxTIiREGA2Wt2srSQVuEUH9QBUvxey35z5ORqjPX/SKZ
MMT5PEIYmVTkyTqZvI+IixIyyadYG2M3rhLa1+PK5JrJ6hLbsM6qN8J4oKYw0riSnsYm4LFOdDPZ
xfS8t5H7Wzmgaodn5LbQ1PceZM3elF7Ox/cE8UVgOZInIQ6qiKQ2HQe/dOiDhboYqbhQwxxElnf/
Kgb5utH3OLY9w50MLn/8kaq5ZXGm0uMBk9Y+820tyRi0LHVGfPK2FXRbRLOzLsYQSsvwj7Ti9q9b
dHfdBJtbGIm9teD71z4OBzONhj3ddW1xvTFc+GTu8Q0wLcrlLM0zcUvDJAnFD/1awvMfpCWLI7BD
GrSwx+x9wTfqw+gHWZDfGO+MfR4I8uZE2xsNvdqN4xn+SaQ8g/9byIYHV6e1zyHVGhj8vY/8WJxQ
QouT870oHBo9KDqINePabN9FcmLUlr0hrhgOjCZhto+7ecQisFpcy50AN37ckAgEPGGJOeYIHcVf
OhF227euIwg3SUb5/P6/CUedvr208kAgweU/p/CZtHw3bPiufXsNIHIHKDUUsm76/x57X8KnSEVc
9YfeHsFdhVr8xjqct+9Eqq2apngnAgY36OD1Ug/wd1b7lgg4xTccslJ/IIPboBIB4F0GVT/AX6bC
Ks6pt7Gic7NvUMn98m75ea40FaA7Ze1ZWlZpmxq+NKU0wUDyMFtZHn7rs1mnGgmYY8I6dqLKhqU3
wd6Qs8GplA89HK1X5idD6ms+isMj588exJM8zv0fmwCx3JXnd0kECuO4GU9xZfGbm5g2CYZYnVaI
p+t36yuirg1FhyzCFh82s6REB7NCsvpwrpqdBJuXqB2A8CUIgGRcoDaWVSH+drowJDKcsSTt94+I
TNGHphU5yL4XbvtZo7SDVOsY6f/W+X1PWy6YTT/2vXvxeempz3K3W84PTfi2eDyluAOS7TSBueUg
+UFCCSsfUDIEXy883oVzr+r/uoKFa2XW1RtyPFJbvrmbJdJVkUo9c4+DJ9ti5002yU/QO4ppx99n
9otNqODyvbnQJ7boeLj4o3cGkL0ixzHxbcJt+xMcHhs30cFZ/NYFWFJqPsp4wRtYwFDa171yQk7j
ShAP4YJESzx2zabxA6bAXVRWdB2ClDINYdn0PiV/XB/sTwRqnnpDFDBZOAf2l+WXqXr9e9E+/Nuy
v32JlUTDrMT2P5gSHyYLsKL68OkMb+XAk6MYJHhDRxni/7oS7amsIf3IFHXAb4B6hUWYXX3TRh/+
IIwFAqQ7ixPvdNpgxdd2jXq+BiAuMpwiTdmU+ok0ll4Vz5YEAnLKNE/4NxpiPLT6W8lf4/otvmYR
hn5Sasrjur8a0mQGJDHJkNB/V6Fq4mY7Wd9mbm3XKn4fysJIdPQI87ZpjnFJzsL8hTK9J4eDmrNW
RCXT1Iu93q9U5FJzNWj2E5h0Mo2yhBntt6v/awGLhpGVYOs9g0bGdWs0i+u/LJRfYvAd01Ksrp9M
mALbCMgx8xHkiJtquO619BcwPDsmOr7LAG2FJUxr17KYVq3EvWANGNBN9/AulrZ9niS/0cW1CNim
Cz3jbHdIHfOqiIsR7v/vmxCfrfEXaZn+wrur2M28ekLuGzz+CuBzywHzbMFQgA00OAexHIc0yvGM
lV7ulMqszzoQfmVZKuSZjtSBjKbtlgoR8zz/txa7Fak2RQemscE+xRrzSYla0Xpyxpha/ikHDxIo
dsj2VGpbV0R3dQ6PwTNGLtWp6voa7jsDxpVwMi1vDMCSVe+GawVr5qu6dC3evxaQe9EttfSyjiIo
hq0aE8j1AkBXrezkBGIzigZrHOVtmyphIq9RfGcl107AbPNkYyW8O2u08dZnXMbv4YalYgdHKql+
DXqgyceDDYcuKmOtvPaDaXfTCyjQMc9lJfjwVynt+vp7zf4M2z+hRMvUioxcZa0x3F+goEXSLhlK
7S7cOU4vd940SLRQYy3IMGUeowaHy0JT0xExz60TpIIQLZFg974WbsWz7046GVbq6PdyiYRpSJF+
jqJfeyfmM+4EhxWCGNQItbxW0QDr6ALjGTewKURlwmkEUxfP1gjT4vAAw7hoX+hlMUtj6Z1Zu/Hr
F/Yjy9HqYw292BzR/PApTy9kWIEk8JvEySG2iS3PtMA1mWHPPMQrp4No4pcXlqUTm3oAgO/PShDQ
xgarlgMOzwophtuLU+LNwEUfiJqNQieHE+63jW8rmEKTUMez9vez3Egux28+rDn9x9S1xKrGn6MQ
COX0z2KxrMph+tVW+NzQgpxeoYXYEfl/c00GdkP2CpLPnBkJsJ10OgjdEJGqxeq5hRxYsHL3we6M
/nCmfc/ewlOc+3JIr8Ov4oCO4Q78IU6+gwHozNVonvsHAqEJg4jwHxP3criYwToCwoWOFpCJ1dbh
7a+PfSB0Aqe6jzVgAhS8TTml30L/jcvDjn8SKGPu4j66jy6Nc0ksOC+qVA5NvnBBF9SbKPVSeBUw
c46WkPD3+pihEF+NCk/mFcw8n55V6Q67hXWNH05+fYGXJ/p3kLigyngRHFpbazgFl2UlDVJgOXDF
T1dVC4NzOBrqJHCKcj6ME/q40aPTV15cbFanX0Duml/Ys74iAl7uJF1MhqBxmgOFc+0guLrWDD/R
kfef3Kz5t38hy4lJyUQb6gFgt/1X1WWGT3QDrG3aXhZRyA+Q72Blm72D3SwM5qoJ9nf25l1ysiTd
9++cscuyN36ZjjBQEXhlxs0CoA9+BT4g2RJcmq+dVKJi02HN2vCrwsj7sc/H36J1Bb9J+CkLBm+0
iIYlYGYANxH6dwTW22wa/7bOB/9lSdTBzTj/gjI66iY6+2pwTNxxudNmF1axQHqX57h0pkVysn9J
O3kzI1eSOokH8Yn2SWSPaWSErtFaN8LIBNWdzhwAtMLPuzibnBJYCuYZxYpdOx+A15oFO4iQkPjR
nGc+vlp8ZRxs5H29r5IZ70Ot0yCugIk3dhL52m4OurCqZ54Ntg73TOr2LCQ/Wg44uIgHu+I/r+U3
26ldGwTgm4M6bEdO2MTapwzJGsCn7d4KAq7wHptJSJWbc+ollYdEzDv7pRsxtg3w+5tuUyq3t+Q3
HXDIGHh8T0AWauI7p46+/E2AQRgViau698oEza1OYgSMmz9ig3pkEWPKCg1CJ1OGlhK2DcuJjo0L
l50sfF/S7bhF74rd2b9h4YuWaJMY54+OXGnf8es7gWOAbE0OvZWRcXMBDA0HqQc2a/V1m4cTkH7J
jFgRBD4vfysCqHYmG5PkRUgWD2wlE1h+Ai2bocyKnzxbXuSel36+fZsLSwB0WOIqFPAv2o8JiFiY
GvPB7IJgJ5xegGtpibO3MAAosx66F62vjSuXgGlsRxmrmLoaciAcKvG2lF4kpQuIEbQj5WoqyEZw
fCLxeYE/D7+dhE5UrBD6XqXhhpWPT3LXq+ECAH5RsZr+YB4qLFAQEGWAfQdUvUFe9analhWx2bbV
QAaiJhebKVq6ockzg+ZXNo9ZkLUQfEj0OggMOFLoMC0iji7ErALWK/e1HhlLZGWSKOrCRX6Fvk6g
OE1Th6Z0HCDViWln/v+s8VpQjZAyCGjC3NWJpv5JQxXwMd1RIQWnzQep92EbItlI54SyyPuxTpCg
YD+c7qi4ij1DCQTRmA+FOkcbi9/c43/5a/RKDsJELLlPKePlXMnCgMyys/M9aSrKFUi6ely82qj+
klCLzoLC1XDEClrcnUsiIrsE12q6hO77UCgEqNpZuHtMQcYHBtjuQTNfYhYYBjzeLAyDEDi9eaJ+
1qoSXgHQDFUoRorwdFOFDN6K/gfmAiVjoYkRWy0kRnuKdg8MgkL7yudCfY8u/Fe/Y1UISBjsBHyn
Uyy41XP381nDd1Qt5ZVfB3ZNKN9Ovz1Iryu2iHgqvQQYMbYhJWii1CZrk3PHnv9zd/f4Le1rz+Au
Mpfz04qNHxYOWb/rvMqlKqtvoCpSxlrnwKT2mCZW9Ezex6ExWM8zeO7FIHjDPVlIvJqmHwWjJkfi
zxJBKn483n1pt5t/bc9jv6ML169/C5TNV4gDYujXEjcSIZ4gzgIbmwGtxUdYba3l3Ib0+t+NCqlz
Z0ekCdNZWyY+0BVtYK7HvKNXCxwUreAtGK8E7hyfUbvkyfXpxn6ERa9Q1fjNaB91za6rQSv4mFQN
T8UrmOA+G6/xLyMWoTUB5UyN4p1O32c7/10P/fbToOxj54Jkx+yBHE2DRp7mjT3H94WynyreAErC
gQ6YI2M/td/zqZqlSc5Jplxe7+VwUnvmsb14WEk6T5/Ez7Ker+hhVUZulhr6e3F503GrfMznkBhY
x9rSPB0MzT0w1eetZZ+hq5XiPVrbGDijFzR7QzTXw5kV2ZijJ5onHRw8Rf+riBNkt7lDCwIMRFi5
eY6lwp3XwszIzIPcaCeo4JALlZP6W3HBdjSGYtpZsE8gpF8uqJ4VuNmc7quisVvxu0Qu57ayeUTs
o4DfTEadfbdqcEEZ3GW4MX/KAav9DqHliNWxTy0YezMpKoZR6L28l5FMjyua6DatY8zQF2f4sgQm
YsjjzqAg8VBNrjU+olije4d6pe01lAmh9Zat0LsJP+h0eFpSPbeGTljnUqrDBBeQ8LYflf2ed57w
1JRo1XRd9C1eWsrXKg+h0NfQfsngZpoqaIO+EUnqhZd+O4/EvoiCPlryvzkco8nP8ppkR1b+ecx4
pUCEA0/70tyE9gFEn0xvPzg8UAi2ak0uBeACRVgdXxHvKih4ZS8RB0rokGTsIL//+BOOtiE3uv/5
nF260I2I4WdKH2sIApA7uG2tn413hNIIFupnas2r1QhYpSegj61jLwstAorxbnMlH29ffQL4ggZP
ZrUhfIGNbl67oMZQLlzzrrg6qaPxprA+jBJf0wke21bGlAMXABCcikNFp1P6gRZUv4wd8KPvLkj4
QPZjv8p47pXcxJch5Le4jQoSSDAjB1Wu37XoH1NswXMxX+btb2Nw3BleeXTOXucdbdeorwrHdOuv
8ipB5wdALPz8Pal+rNsIjiU4+CwwPCD1RNq5CihSRn8Ye4q8Ook1TTI9JIHYidm7iDB5RDHcYczO
saUZrmsnzWvf9PNnLPIhh29DNOu8oTroRVVoZlFJZaCxytdgODL8S05ME9A+W7XmJQ2sf5sPLrKm
Oo+pyHx3+vblyR8A88J7/xlZFdJ3TDJrUg4Utaw6R2TYEmFJ7EPlO8ZOzGn6yayH641kLHa0OteP
QO74cWCvA7ept82/FNwazpBQnveA4tJYa/C/O5Hg3dMirwdK7fsTpP3RwSjy9obt47EO65zXssFZ
+7mJlH31J2qWTXXJMEWwosHHH4WUGyNZmqSjvJRHdkaTNh7UtngmFdyh2deHISk4YJRmxQPLVBgk
Apu0Aw41NEDd7giWfjJVDjXOVxVC4DFfmb5bxLvbPaWbghAVZG83IQ4bYElvDjWvX5709KgHHFYp
qqIqncHE32DaG/cFoyyLWtM8n218vyp5PQL/k18yEAUHUtUaFMM9t/8yJI2AEmcaYv316ATTR5qX
9iEsZkwyGc+SKRBgdHf76qzMApUDDkktR9/hK/8+y/i16+WbSsd7nvLz/2YLeswx7VT0exGbmkuE
/hxwLWj/3nYcErc3hWFkw5wenIeXERJAUrnXmfQw19NagYde3X0TTmjIfRcndz8Q/zc2kgcxzCki
H1wp+2wbffXITQUahTMyCLzzKq8mkSTk21k11Eog7LkUsxr3I1BdR5Hop10qWVU2wInyiiNGHt6m
k4uYfJ57avlwx/68JXKrvaWxsFMfvRCyar4IUHPBMAs1PEpBCMVS3j4tklkxN1a44DnjPGI2wC5H
8xblN/clKrAURmwswTubHAM9+6od4fsKLluj6TUSr897pQRfjQfJxQ5cbQDPdQvHC7fLcF7ecGQo
3akNlExFMf4NEhxQ0nd+vNgkvioRv2ALUX0X7NppBpUcoJattz8620A5pyNVYuMCN4v43Iti7sML
7XaFquuE0XqnxUNj73P7dlvv0jknOnWEJ85ZOINQSxlssgB1h+i/EKppDaMw18F2QfAMk6mAJrkb
kPnfOKRMWHKaQ7gi6oOPd129WoAoK+vqsCwlGehLKSMdzfuu2ymN89/f0aSMjOmdNh77jmyHf383
mVXMwCG4Rt9U99im6qYA3XhqvEKCSAMQIJzPVHRcP+/2zNe8M1BUdyFimietlbFj5Mx9hrvfbcdh
zc2xHqvC0VCZ1RE+vH+pHGciXVv7mQgwuOiUEzVj27XH/I4laUCTlFC9s4kd2MAOfshlKdrxB/BX
eOUcaJkPHpM9i7V1D/Hdi5K83H96aDtH03ZqNrgv2QHnUcVJO6yaYENsuBIcBkMTlTes1SbNZV3Y
dwD7S/GVIlocMZg/D9V0DwRHCsMgEJqWGhm32oCTlAummwQwk5iWX7LV6JGS37/RDM1kOOYHfNSu
a2XNp9Iy+IyFK/yJhEeleBgjeH6hfq49D+7JRbXZPYXYxUsORjhVy+NaCjjSVcdItzdArLARvK8o
ejMzeZndyVyxrvazUXKDm5rmn3OgnUqtEYyEWFx9zTbb3UgR4itXqDaW6/TcNENFVfemD3KM6aKL
x0BMrVCWAnhD8P+/t0t3NwMsSSzqfV4HPfL8go0qfYfs7BituJeweVLU0FZdMT0ylLtO9ac7ZJ8L
8fGhvOnw6bE3aXdG53F+F7m2vcSqqZRcRNCOKmFI6Jg2aPn1tUIpJJltjqcV2AbpxP5OiDLRFvcg
UjCTmxXPiiSp6eg2TDeYjJOxYPkGbOH/i8F4PjfEy7QUkM2Y8UnyWb7dB4AC/AT3RLdHlfcGpUsB
7Hdg/A9TYHc2I8Y6krJqN9EwUlbWyR2YnhNTPl714MYo44J8EJCBXuxQP3SGpNiHiTMTs1lll36x
l8XIqrANcNe3wOQ/+7axljbx+xGycTgLmq6ZCT6ACnZ2fWXASXdcUOZCFdGkblio5foJ3bJGx/+j
zNwZMPRTC7cq0cu5fggodM0wqzZTDdRpDEdeJbZppKhYxb1+F82lpLKoeQ/HvocUjirHRjbeHCat
Sq5Td5+E1jGDfWKibYtuzfrY/D8a0szrjUBXvO7TzsbATi/p6hIjDkLxeTs0reKq8FUEsgPgmLhx
3G1KKeEYCB++lxRyIFZnSuJm1tFRjVpx08aNySheXSIaKXgMRcrvDbwdRJUYnaj61o5PCfakVGOn
zDtPPvGRAx/NtSRpeemgKbJ4WC7T57Qg4VPD6hBlHwH7PLKVF/BPCpzIyOM0Rk19pYvDTfvmqwXn
YYZeopS58A0A8qhKMmVFVf2e+kY31Z7frpRUolgMxA8bDjyhrzpSPBwUWzIri4NSHyYoAYjIQPEC
NF7BJPZY/KEiExhKRjC84bvZm3z2PFBC6HOAeHVnTYjfMgS1/bDguiXgtAgdeNMauAb5lAQ/iCDD
5Qut2YyGy8SA3p/2bOmaTC7/sHddS2jW9zM5LXVPVlAQePGT/mSREPeKMtBegvIdg8g9o6NH/p7f
34bdENi64cE4Ik5q0f5r0BgT9wNYSQtTZb8DgtG1aQYRVu5y3it17LfvOybfqmKTzB/euyYxeptl
fR/FVvRUNIjcZt8LxuI9ABWPooatQsknSHcCYWZdu1zzOaJT6LABXl60oBx3oAwGQNpOI34tfGd1
Wlfk9emBQhMmjhTZfwz0zmKK8ZO6dx+xzjafYLTG6KXSI9WJzy5E27vhfhGyP31DD2ePcNFdVRmm
vTS8IyBukMfR2CXOAlzLMLazbQUXkY+duTaincQrsIfTtIwGZjPKin1PmjL8g3u7JPb2WTjCsx5W
F5v6NB3ONSUyz/5U/O6Api/ncpOK8wHswL4ditHtt4GLZcSkVbakskMI3HOUuPuaUh782LbZNuEA
val2EaL+wsY/ugkbrZ+4so6TOVjIHNsopX6hyuTBg5J8FCnShkewnlMLHLxPNJu4EgYtkP1Nxosl
BlPMpvR7tJHQQnQhSFwRO4ecGI08BoXjwNOiJh1v+Mw4SFvjMSqYwWLdA3WHGMv9BiuEkR2IUiEy
UitYIirLWjNWcUyLzafWSKcImUTzdxS899TDC+J/Lo0znZFeUDSVfOcJOSsR68e5pDC91UFRXjFo
whCeKPCYqO5aHIdxAk7vzKo8nuYEyjbdlxp52mYQ4+XFKH7HL1iZU5eih6yeg+5MN+MJCzafzFnA
oZJ9m4uexHNLh2W83m8ITyDhSIYEbhtabAwIy3EKWyKdXBqee4tEaczyjQm8veOgoeNsit7n8xug
4XukrCaEBLRPsg3hOD3vtK9z4hEyoVrk19NvomYe2eI20sbQoVvAAElZVyocYBu7nAyFzORUQolH
lES415oCvj3q1vIa3ghRQ//rQ2nY2khCaxCWQFHzXL/sRgxpBXNPZnCTGz7+jKehwT/L9lSuEgfa
u7t8cCerridyYO2JN5RX8kG9H351NfzohJcxf3cfGuSrEIt+gkGg5f6T3M3qf3o98qdv9nDibzF4
BL3jsNRiffIKCN2/65E8kS3eCvuATH1VkPBMd5GmTRFjDk4lfye3yZCDWU10jrf+/uXivV5PcIo9
jRV/ACnjrgouMPLJQN09JozZpBzZq49Huj3wy0ZamyxskdOzEKvDjkKm21AEKscFsCPxi9JVnYx4
6Nd96l0Os4MEwgyfh2Iu5E8lqVsMZVz+4/n+pJx6aWcVlu2hBeQ5dDEYU9nj++HFCErdI7jQDAYX
VCIyURiF4O1Zx4X6tpkITkh76niFTYcTQ9UG7nRUUPUOpTwZHKCupxPZ3UiPKEMuuB3ZntTcVE3s
roQPW9qFGD7ICTrKArv74RKY2smkssELyRap5pcubr1CWS+IdM37VJYcAjAJgQopN23v6stklxpy
XFezQ11yC6Jr6A0iChUpo0N5Kx+949OEtCANFuG4/jmXSIU1hyL5JVZ7UXmhKmKEq9s7MjCJnWDs
afbekO9VVCfnd0ny6CSp5en8ZinM3cFN40ghgspCdw4illba7TXFYA1gIg5gDAwJJwyWoaAYEbNb
VjO5GGx2B7iz8h3Vy+i/VEj7k3gJ5ZzDixqotx+GwK7GzKRoXg+zelnbyrjHPWY0YDlFyJd1+qCY
CWK5TTlZ0YxlkpR/5do/HwhrC/7K/3/BAgL9aeGRTH00o8N4zgmzOvRah6e/snaZL+iA8gYhcSt4
uagsITV9c+pXZk+J8dI1SaEQSDKfDQQYGQOWJw2OFupZ1oGq5HoBBOiM4YpCeflpWYkdhlRfsTzk
svl0YkOlYK/7tvCLtFwZn8jw2R3YSKqLdnLK/OcfNThOH1iBeHVCpFbsaCvSjnnsJfIqIr6ljsib
DpZzn4xvNhnPtrO36byci/rfW+bnWvCIqmCdNdxx/WBFIoQoH6bMiNxHDdgsRWqh3ugnbFnRxvg6
iQQuZImihBU1pNksZKqeAwt1OUPgn5eCxD6fb62LikkpqfO8h0jegrwIXu72qrDcX3BHpkbvbRVT
dX8n3EgskBN8sHMfs9b6xQcBa0NvTxYJIah0mTFFdIfRUZHmZ/qS5iCt1R8aj5WBIH3qhdeGhR0N
IjwUs2FPBLnXLCXNApt3JS450E79pjNWiJE3cmgYdmeR98RCQbsN2Zmnzgvz0DTMdgaoapq/pFdI
jfFo7z4ASfbNag5QaD0iF3DnZMDgHjLN/UbMP3E9JEvnxeqIRWP64HMCzVZMhpMw9uEMYx9qU8PM
i09LNYA+0AUJOhtkX4BE3pzOIgsBMtFmQUJVBciY8cwTliJ6Koi4IqLLuDZFdqPpvCe66fkMuyV9
OWIoO0P0iy92iqIhPX1UUpsm+CMPV0DmkLBpzryo3nI+PKin/eeHDb5YskZXUVRQwdUVFd/OaOp+
tTshLBFkkLDnkELleUixavDGlTLMa/mEtwhYxIUG/wAfD4YxigYVaOlDUMSkNQw3/clV9xhwmOHh
Ura7lQX9ZPe2WDuXrl/cMFP8dq42JUKgMj8OoGichcLJ14KLZK7WcusFNYH9cG/1lKBCO5llHx57
DZpOOTtgMmLCzfEb88HlLp/QjUFzcTLIWhuiZCKdz5w8YgmUhtZniFmt/XmYiASRr7SjB0aqIsr9
v1uYiD1kHJpw1Xj9xKkbrO5VfEVI9wQhA7nICvXHqU1owm7/P7wjI/aQ6Xar6N1fcVd1w7b4tJ07
c6WxQN4we/gWiE//zzPu4AwksIviWLlY9TcbDchDttbrl14HLY0A073OWNlxDEeBOaZpdRLVXMvH
EGvW8MaQTnle/c/pjai63DV1ZSWA0q1xBr59vWjM64XJlw8UUWiL2Ql0+OueEq/PBBQgTw6ikUir
aJrHnICr6FNtdQs+pbRkYveFJ4eNnw3MQd0ESsfX5Va5c8hu7SwlPCZgG8DzIp5aDyDXPTJFXwsn
Fp1dpQbmfIM3IYiaaf1UhFsaNjIOJddf2jh9VdBP3KxUdrj58weRP/81kzyxIfB4LWJtfp4GEUYM
EVxi/NWqRvOj2Em6dSUGhEXCnu7ijCaBCM7bvsi2aozu6S6ddO8Sca3dBFBI/1Hp00K01U0fc11W
IpYNLRx9xl1445NHDZyTj95PdcxSC4rznc7x2aoBnpfhkTKuu5F2uyODnZe58/5JukIHCia4dvOs
bUjI69KwFlVOQmOeLaZusBjdPuk3MOOZiNPkRGoucwZ0hWmGCjWbLm/M0TFAw7hsPS3a8cDztVcM
8NY+ezWhjpO9ATJoRCe0C67jqtKLhXvW5cWHmac0qhCouORlC/hXHhNRyJCc4G6iY+I3uGJxFA1H
XACjTbwMSlPa0xBOiwoHKAqhjE/hv0r4VSYwUXwjCG0ZYxJCmBYIvO2zC/e46dzCrm/zeCrNDvc7
hI/Qe4Y9nj6Vp/fRZ7sWMrY8ePiUwo2tmFgl1sfbUMni4lZ5x2PO9nVG135SMwU2jz0rzJrDifUF
YwrAdTKOj8vbkQv9/9BkEygCMM/+UVZEIsaQmuy0OESWj7aIfaj8Mn8jJbvVvF9RmmufzEMyO/aZ
7jSuIzwZIAWzed4kve3x0omCpdllK2+U1WR1tfudULN47Rb/h7aHmDzraL+ybocS6djaXw3IlFs3
s1NzNVGtdsPa0jsKFFwiFzij+meMDfCqtUs5gXKn8Ua+NaQlN4CuRfaccHSOg5t3cJ1oS+kK4w+0
XaoLKBq5FDHZTmKbmdmeKZmqhGJGj+WmNY0DgLIzwKY36H8e+Hy1qiiEvUrUbMpH+pgrIrN/a3Td
4jiPmhHT8hqiPpfqoK2MHfHa5x+U5sLFLtJVyfZvdm5i/gO4k0kaVY7BpA8x7tG62E+ntUm+Nm+1
tl/wn+a5bLR461Yr2hTmWK3cIpw10NbU3+YnjiyhjgTa1aGcm2NX1TPWLMkDdkbb3prHPk08txEx
neqn7dy/O8H3Om9tNJ3BdOStWxTIm16TebfyAMGtct86wUJU0vUyMvYJEaFBNKgL6WAf6DGPnbbO
X1GMdRo11hErqg0S17WT/4ghd6NA+DYchmCv9Wgbjucp6jTFCjPZ3nP9T393etM7cMPZcnnmzjyw
MErB9TGN5GDFIKl+TpfKXUhiTIHy3Hku8DWc9yH2b1toU3q3teXeO4yFQp3KTatfFXJr7vxFoHqP
UsCcCkVaK2XFIaGb26WwlrxX0ceC/1Shbu8zebeytZh62jbO58u5IVqnRrhOmt+TS0QXdRJtDoOv
Hl5NBASBfgBztUFrfZ5JuBk/Rz9sFN4zf/UezwwYXjfcYGggbJ9jJ/tfrNYAEfURNfMQpalyrQ0t
3XPf4nGDih8a82QpJexvwojPEm06xLYHSbuL1Rx0gI2lCmow/jDmKpiFvfN2iRAum237+iRsjnZ5
e26/dDUYjp/C6mH3kEvBcaQZyJdPWI2sHQdngE7TwEjoa4WBI1R/mOUL7Vmboj+q4bwJ2CUQFOcq
dUnUgax3jvcwXO/I+Sqbyo964znSz30D5whG1kFTIbShemyX3T5q8q5aZ2/LgO0LJ51BN7l2jM1g
IkZ5oB3rVkuqfqDh7UVGcKdpqrj6BVDD0PE8oSuF+MiaFKz2vdMwtDaTJNARmT8NXf5MT3WivPb8
iqZzxiHd7KZK0N+iFTmvVycKijCsy4bwyBks4zuSkw7AQHzja/3AfECKyY/NLepJHdJ7kmWhqJ2e
zmL8gLwejZqCu3Hiv7D+tQHtCAkfDbmyTQk+XtQMFk1g3DXfFiwV14wn/Qwe7ZciJfSr/xxHkW/M
0RgbkdwJ26tDRL9tI5mat+dvmjfV2cZ5+QS7GYdvMHbx8B5s89kvZ4ovOGD6nRGYMSESxglOnHrg
dkh4eQ20jizrRobO0XVaIK74VMld1gwBBTSxeVJAB0z3iQtI6XcWgKMJnxwh0MY6P5TwqFICmcti
bdq8QDGzoyYvRDi8I9fNaVRlaI7iuQQv/+NrXez/oH01CfN0YqUQ4GlzpVJYLmZTt8qtddRFWhs1
VQwATDH7GSJtLc4dU5k2a3xNEWBmdWsM3V8ThOqkz5yoDiHck3jh/B6yhdxmZoQ+9W5XPFXg87nk
jPkcTV0bPoIZCQ4pTwNV64dz2ssO9Bghur4nBJOjbs5SWfhstZ+4gYry5F5RP7JMlLXvwah1gFO5
vfB6wpPAO+DeZBq//p9IFJph/EqPNayzTn43JyscI/f53Kdqh/zM/QbeVVI+wQa9tCvcZyazSsB1
IY17fMALWBlzTyChgBQCzlDKHryaD9Hr69G1jNHY66JApUb8nwV4AycYuTw/I5psdq4VGvmc+/hv
lrO7/d6MguEYZHHpLds6iiYdRau5AB8OmCS9SZClWVLGvcNd3YN382wDQhI0oRAHSVBLH0adNOmL
p9tgvkOx6etc3gDgR0/49AGgTptDi1klwSByGvv/9znHPx/jhIyqh++RmIHLpsz/ToXtYiv4SX5H
+K0ZO4KFf7h6XByECGZgqqb4x3irCz9RuS+H/XtTwjxhX8r1X2RyemWaiLMNCWYq4wd+P+mYPnE9
aPxR5+IMwkn+zEJj+Nb+7+wDfD7jEa8j3uzLHEvBBa70rcGyMQLY5cmWjgcKXsX88pbPQ6j/5poW
cGkePiGpoBGrQt2k7sAohmma0GduHbVXWbV6Z7Q5kNtecQ62cuiU0Ak8QMRIuFTDt0nErhnsBFPr
n9RlHL9eHYBdx1XG954DSyKwc3FqnyxusP+daXLqjdX2H0TfDOXgYmLCBYm5u9SvduSsdNnXjM8b
p9LtWAL0575eAQEB/RmuOZZ+T/0B3WFVULvu+NHKzoYAkVcRAthMIyMGBiH12dPGvLzI7yxXlEiL
/tEDKl8j9wDWqwaWZjPCS6ozfQPmdgIeJ/L3tlGtOwsqUrvIshiNN9c9GCEhVPNIAiVR5IQPFbbk
8bU/z67eoHx/mWsUj/1XQfAiEkIBApYMcxWwG4xt+imTT4u3i60e73KfTueRC1ii8sBL69jmRFYq
/mVziWiwTOxReZAQUW9/pDAadwKHX5jJ2HwK+HwgfJlG6e9+jTPKtr8gGDMO0Pe0inNZ5+Lgbys1
FtrBBSvd6VcpmfOYkBw4vNgF/nTv+5Xp+So/nBHVjnPH2V1jDOXUOHmhJVp6Mhl+sSmCLaPB4P1k
jynNST76x1P1u5EJ5HFkYpd75UzfiZl5vlti4tHIC67zxwq8nPhlKXaeppUwTiKD+Wupt6STcBvq
Y8TfojrPx7OKk8Loyd9+svxhRxPtgcsXfpPqg86aJlgdBcwO+wxmJ9CGFDYYZeB+fAR48SJ/tg0M
+GG3HarTLbEGF6H3mX3NUuWyPqhxMebiKkrlvSafTXbp5D4/xd2DwPZ3hbwwnCbww+8tBPKxY1BW
b20BEn8WOpzNqLx+5n8jl0YivONUM9aR55L34LpBeXUqM23/5IgGNeqRfhgvOt+KV/DFa56mMaOD
oC2xSsT+m/ie9ycAobeZsPmffhtiWX27LTh0r0H2qlsDVNeYnVIgQMg6ct4GGe7L5RSMNsIR5UIH
hNeN+7ddTyPD8p46rB/fBnFIaSKz4jJdB/H8o7LS1I6HkaI7erxVLagW/ebK9eLJyDjtSfKaKD9k
l6MpNV/Wd1Y8MiE6gIYzRrtd1ExHXCB8jrGBWKF4QuYzojyWK/AZTSQOXh3GvwDFnbaB2sDQ/P1D
mN7ipNkyUAPxq0C2BMQXS+qQuMF+h27rlvMOJdfnw7ZWH+iR5+GChrYKA+zx+g8K+TsczO6WovAW
C8kSRg53WSt762AYNtvoiwtwI6Ki32C/xWbAZf6raXC2MsKlB+nfEfOMDRSmqNotx/TiOWcAeH1m
vnkmhmc5WJhfiDuIw3VTur6hQ9IEikKCnkdN9z7GJweLU+8xI/+k0rpxPWiwiyCMMD2lEpdBbHfa
60gXXIBW4HeKyzxGhrK9B+dAMc7t8ktxQ8eHTWa5OH6TmbaIf960coD3pLeKuxHe6+wA6viJvKDo
pRJZxt/ZzW2QHnU/cow2LHtklyonDWhAxCepXcy8et1rJAM6elw2QUSkZkywaLUNLCZoCv2L1jXG
mlVZECJTGMwbe8jn++dJeZXjFQGVEXjoaO2yCOX5JRzGPOu+t53IMKZeQBNxvBq4ZvqtpdazAC6u
km8etOO5q80qgyu+xdSzXba+4IeJQuxQlg8s4wi3qo9AEUCAQbzvJTtmckkGT1/MSwnx72qO2Dhx
D5zlqhBs5ieEphkMu6RrnzOEuY43Ay1z6YOMrcZVSPCbV6u+2nxyv/cZ/87O7yfVN1+8QrtPfNMp
D5Su632J2qXkT3LJq6pz0Novkfzg48fm0MxEcf7TPNmnvDKDaafBpRm+rk3TFgFeZurnFCnC4yPq
mJuKOC3E1MpS7eoAcCqrzZtzXA7Ud0TRAyMM3qx1Ex7Q6DTOZZyddiITjlANyXAzRUGJiwSDEPOF
jI/rmN+dhFjBJHgxVyhBVRoynZ6Iuar/mMab2LDafH5u1o3qjEbCQ2ZsIXbcGLRtZ4cHd12aBdMu
fJNnKixhbVPZlpqTwBI7B3LQjuos+TjK33vpbJkevY/BSaXFLT6mQr6wBEgB8In+44eSR4vIn2ed
HdwDVEPKhk6SSIheSaYSyamqhdNBUXczhAyBiMJjfIJabJmb6ZwVT3GpK7BiBTU77eG9cFD6VjI6
FQ2cRlA7CvKxzxFqqbpGDasU0sli5y1tRa0TktkI7bvKXvFVNMlu4eV3f4UlNzTreDeSSFzHYnpe
rkmGqZmIIWudE8TEnGoyTU4767zl6NdyyrHZtv2y57uaqdhfIFtd5v7tb9fZ15hKMY17iRaL7bk4
kJygg4RezXnH4C3P5f/C1D8HYjNNfFZnOPqVZrLrh2LxICZ09hMp6iCbuWWFvpHiYjDxHMOqtbSX
POrotzUH3WIPbnB6Uua9EucpasU+8gKETmQW342804hHRVlNTtte7QnPdXbU1dvL1HQtM3ibhRQN
L75nLADM+ArpFR5GiceViybo/N1paZsjxFGaP3d2Yu5vgZm7tRwxa/sQerqR4EELTRvjeLoYWtD6
LOl6Qjq+58cUZZdyXP6IoipxtM1j4m/f5G8udh2t8n6qo6ZdAT6lx2VZTqZuG4sOsG4l0efY/oyn
qeU1CUKPSOzMogpIOIlgHJIMzG72fj5lSg+RdjnTadaevY32O+GQ98Y4juv5Z20/U7SpSOFu5JpC
63pp/C2py0IlfxYVEq1jMTNbEvIeY6aUYQhQ/Xvtiqg9qnQeqTCjObDhY9iIrTbbA3l/CjM6bS6h
1vKo/g2BypVwpT6XRrIg9j6SuFwXl05VXhdyj5Xql58QOBxcb+k0e9pAnXo0T/fpg4kp2abmoQgj
sE1Fd364Lsj8UttM+g6HDt8askqtvKcfOxZl9PYyn0/RKIqzP0/A2SJtg5yd1uIRT3TNxrWxLupo
OfZeymcD8khdA847dU8VDGApD+T7ah+IrH8AIRCbRsc0jKcffNA/g2QqmH4TEoEc77wGiZkNIpNt
EYkAGiZqwsLtEc2qgLFI6GW5ir67V1lZa4dsbdtA1YKOSMGRX8gAjLYy9JRGl2lXLiWqz93fOhHn
cUmN6i4f81nQ9jeuz0wagQsZYXGzRIocEadm/fHcjYq6nM7zxErfiBuZ3GWMu9fCnDC6ehGxXiUa
cS1RNlN4uVIYMWK3TxGits0FP5jjw8KZO6DDoBpF1bP8oeF5FeslqVj6k4XLakc3cLMwWSIPeDe/
kdFqKcMgpBj+8FCI13H/f+gaH/jNAvuFyAeg/YlF6/fh56jwTDOj+syriYIKENDmVofEOJnL7+ZJ
W2MTOWVnhGlutkuyEXbRZKD4QV7KhNbj5bHQ1mZ9Mh52m2X324hwp/hz1zgPEMEWqMHc3KKY8dCu
WQFUrCCN5UFL4PuJm0yz0GV5E02cHfeTO9PRRJ5vv3MJtHklrjQdOWVzwEiCmcLb3iHOTw14fYiJ
o09K5zJNeg7mYIXg+9h+IOWiJdcGEN9ptV0J/amVo0vYzcu8Rm6mPnfe7tyk6tz5hab40HbmerNM
KPUGoEgC3MMohCUad9Bu5CuEbYqQgnm4L4/1BbstapKdE5mQnQ4uNaHu4NUS1h5Hl/fi2011/I8/
jUfTSPxEsyXogNGNVC/UCtJ1BykURyEhzLVAIe6YgfOywqWOfQk0mC5Va65LCUc3yIsiLzrfEGML
UuleeP2DxD6BA9arwkdsrnYP1cHzZePHBQmsP9BAenn8ZPnE7t77TqTIf9bL+ng+SqeM6O+MWIIA
+n2UkUld4sGByp+F+fiHRfQBu8kxgxwMep02uqVbBVEI3k79csfIh8XLvTdHcSTSRixhkr0S3N+N
OX40UTsecO/4Sh5xMhbzZ48OAXV5we6tNi8EfWVA7+uTe/bA+WT7mixRMi/feKjWid49RScc5Nj2
ewQvU3Mh7G+XC+cxK5p+JKW9Cpg9X7k5W23DLKbLZEF45S8hKn0ly8SwzSV3cFdtFcDhiBxBTYA2
TJwAULTAUX2gOfeD29qzHQL0ZslMJDTYlKZ0rQ3fpGhBEBvTQMZrRWBzyhfmnHXUeGCPw0O9fOic
bpUh70wWN+n4xPQ3xReQsITQV/c0wfXWDNqtISls2J8BTYrqZjB8MlQ3DTCAJ4ipYgZ+idWg7+An
iVY8+JQ/tL/vczYSzqhaTcYeKLChLWHpew0xg3UG3soRK+T56JebCM6F8ogblFgS7wLaYTfcs3k9
EjvsKDOA5LkB2I9JkBAcDUgs6n+T80+YyOwnJpzsDBbMGes6KXJpJu5voQXM4idyLkI5CuHNJwbi
+ioYi0XzTZ69Sg/51exiEJH6mFZCN1zPeQt237PB/4la5jbSqglhCx5zoeP7PIlqSBCe5hq8lnjb
mdzvWXvuowF0Kzk+erbO440g2tGKOEVniboPTcV+ONyfMPcfKdJ9oyn+UsbiMYSFuc4bIIcXaOan
cAKyFZOAFL+US5Vq16kjjEy4zlDAsaC6ohPhlZ+SwLCgpt/rbwO8m12M9zTTPMfgJPJOtzMf6u4O
/+N4DImZq8G7QdZI+Wd1DgIZSLwtandDuiI8sWWVvPXA3A==
`protect end_protected
