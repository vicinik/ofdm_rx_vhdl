-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tadiosqwzF++DnFtcAgZy1CH7OeU/AoKqMDiDuTq0vh8TmzpvU8+GZF4dIXE/zO5g/x1siX7uRDT
dIMJMJlJ3dKbn33YVf/UDn0z0KTjUrMWWGLX+gJ6EUMuZfMw1Wwlz7bbrTHbJEuzcB2fD0QFSQRJ
oObq7oIoWD36g2gHUPys0bFLKqc1v/V0+c61O2jujgzhSXOw7kmM6p51fNl+6Tp9Poebu3bevYvJ
pJ2kMwsvncFdyz6z8Q0BgFMe1du7Il6ZlQmZRzJwe1Gc3EGHc1GewXKdJ9aBW5pUR6YYpV2MmL5O
tEoJnmyQSlIzsYrSxXOZt2sCK0x0c0R4F+zM6Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8880)
`protect data_block
Net4ELUuxV7SbB/b8osSV0r76+xjsLgwcGsiqYQ5JCgoFIMZPuGIa4OpPcBrPNgFG3bx3c8Syx5z
Rf+6zI7xmvDCpGkmozGdhX6xt3Kc3zw+pdzMde22mJrukJdT/hNhwBlENEIUU5pRifYY4mzgTQJr
IfPw8lpowWsYWcAu+14MOYvkoEoFPcHcaC7wOK1JuCLILsbNbXPam01ZXd5prbFgRHnQOQT62G7C
d8cJbwebGHtlFJmM46CAJaKmf5EgLllBD9tQpIC/AmnG/KrP2iXMaKfECtBgt0VxN+LLt9UAaPkm
QnIRfM4IsIbAgotFKr7UH0mYJ5WFN27gZk7Mt2dR5GTdfUZ4TuJ52Pz2uYfHi/+U93M2HX83pZQP
HYDFm6Qze/kJFAn6RSpqEuWZdBz+89Xe07y/SLDof/T5dMyNhXzuyTC9NCjcd6zYlT/FHNBtCEk0
0x6huQdMX2WNytR4V4FJVAfeT+feZZxXBZUc/R/js8eQj/Vh7dfPH7amZQ3XCnDTRDNOWz2U7PPD
5pgCXw6s3+2t+Is+8h2VLbaq6McOcCDCqdu4h35M7OGvicwQcB5MNuvO6ieTtPyvVg8rEyHo9GMC
uvWe+yIFxPNCt/3rAtWM+aWD7eY1KFoxB9EP3+ij8fQUVWv+bRA3/HqwYLvR+EAMmeYSohDtcFX2
seg8xoktfbNSRP4nWpyJXNuzz6h/5yblAUpOuQchk8jLZ3gK059wUngrwgYu5A4syEJ09nQUD6D5
felVpFbqKxkVjvglOZ7rG7SKhQlIDsFRxTl8HMSfUBMxYli/4Sct68ycLmhueC8ptdJonoIJjvy7
vQDQ3aRuaN+sT6A5aUn09yCO4GB33Ka8nG/97HYDTLMFmlpfp4HDBNVWeM5zJl6qOivNPBC34Gyo
LY5A9pPR2t5LqK9AZcPIyUCateFOHZPrFQpaO8NPr+7sYbWyPwbUwjYh7hATjpv7wZtJCeWYBEmM
X69JZWHvYkZbo2iXhDbhPE3QgwRgieoT7jQI44T3g6cDdGTxQpvh7Pe6BZVHO8fsfGCAKpyeH9Zy
bvB2avSnhbB1Ce+uVLi2OVKB75KAdcIUvLrvxlSL9lECV5t5lcLYP4RZImk1N2um+3+uB/8XmIfy
fFsawosFbEa5yigECOHT+1bpx5DBX9UWt7BXZVNivHbeuFvLWhWCQLh544Wf+t2CGQ99HbMbJYpG
FhE6kfBr5FEzxKlwgCxTpqgnlcKjf6YRVMlz5aCfE9EOaEv0NJkaDXaPL2T8Sdili4jrrZgUASOM
pwQLYHwr4LNJwG+uBShuxmaCZely67Np1rNDNBYhaGivVaJCRIM2rDmjKyyhaSRverQwxsbvHf/m
Cv/i9adUpcE3M5dzja+AM7MjanPUzNFeKD9/MfW9S6+t1Cmy7OKcH5xdlkeOjO/cAdI66H2QNoFN
+kcROXDrI6pYg8ax63XwhZSLYgHjHZ636jCydan5WCbYg7vzUnbWdLdsUBNEgeG6l4DNjO7tkCQ0
99kPOYUMAzXKn9FgLtPYJ+88QQ+K/9N4UNxB4qFgIo34dBdbvPNNuG67OaR7JfzQXx9soww8qKIz
CCxtXtvCG5JkjRqsiYoJavGAifM+acmFYkQ+keJ1sdiMewitUgXktHsY2OUwwVWyEX4281fc0Z5E
ReLfBHE9lKgfxub2fCYPunK+I+clejTRXGvr4rVmozzwCavYnkxRUnL4rEnL8OEDW+gFDqtO4u/X
y3Xe0t28cSAcKa46rphmjfS78tbrLZnx++Q00Ipmx5v++mws5+bZj9zfU4Px4bUWmaxDYHcvPQye
1WTXflnoliCky9H/3FEVNJi+68/Ot34RqNM8VSfuPOgEdLLvLvCYtM1gVXOowWUhSQZpz/QV3K3e
VXUXbPGMUcPwf0qHUz/xpw1twvq9IW+Lo4Jg8+TLKmdb+/H3ZHjOvrZMoW6uLo30rmt4lmXf80Bq
djJj9BJLWEliiKQnZRXrj8EzkE5fvkECOU+G4myqDL+6a+HtpfIxD1dEB0C6y+iL7RjASBzsP7py
jgTV34mSoYSEo4STmS+kC61ReAPJJQVf8E0qNMU4mPsSwEukEwuEy6m7mlRpXyayF6Qz5cfzERia
lQQIbNaDHIHIIgMeLnsleMj2TEJbvLkgzZzvF9z5FpJtoavhGywcxg7RKDSJysVIfKlEYVtz8Kk0
7e7+niu8WNIEddOsw216kzvqupm9yZQadhBM9MmtIUh+LlSGpFgtYkZ1zh+QqiRDt/4xiWHpndHC
ZAmTecVzg3fvU8wAlufSqFLKnRKlquEOV2rRsPZ3omQg/pthdr5SsS2dHIGWGGob0T8mJtY49mmW
37wPIcysekaE3Um81OUlzmKkhUjKBubQUWGb1dlUavQAJGkg9uU7kx3UXBoZwrtxhzd1xAtG+Jbt
taEPo3eCq+e/fouOV9V4OqqYLaWhYtVy/1U01We3vW6+MnUrRJBkrxtIwb1XO+LOfcsXVXGJnRFS
y/N5Bk1cfYZrpkR5CUuDdJ4ogXLpQ5a6aqoTlZNyRskFXX2bsj5vwvqIyC/TwagfCsOitUU+pZnJ
dYwnENOJ68jHgL38WDGoabvq+JcZVTsAszf6/ujrbJKFL6zZ0LS7M84m6lVedYSqX6Epen4XgKer
YPtmmQocLsJCoSpa+cp2ZkO50TNMV5W7V1jo1R+K4s/Ccy3KZj/dynVaG+QZ5hDRW32ui9bpITWs
3wMKlUwJFKdPZTwOPILB3ID7ebJUeTbszQ+9waqJ2Hcqg5bkqz5c0xuK0oIm/2T+lgZlXSdcec19
Az682zifACaD/B4aeb5Z9FB2J6t5TrxGf3Hm23iFD0atZy+kPw4GJuTgOkk5jCLjaHaPCI1V3xlA
uSMfs1verVrnpesu3EEF34zw8fhEQqZ8VX5IaxCa6nF0wVANx+DKy37mTmY8+ITQoO7VgZ2nF1X2
UDBoB5caHvWGnnYUvh1D4PmPBvKiFGAy3QatQTteTdxHkOQmkz6fXNkA3pkQ9fYh75loJ5OIQtF0
pTggZT4dSkkDGwXhYajNXZPEGEllH5cIhUnKepUIxrn8MtvnHy+BngzItFLOFS8wsEPteQD4wuvm
bViEsnR1TxI8guWzTX64qwvWJuMbqZYS0vls4e/L1/Ud+brl/OXPUYPg5v7T0tNkEFsfZVVoox5R
ycULI0lhg5uJ+wFWT5HL2RUL4983lIcBARGy9Gco7SxrPzlcP4JGdvqoguUfc3l9f2i6Tnq6Kakp
3JtXwgpEHt1ZSRf2EUvPDU61MZvfa7LsB02Ui9jWBpdONEhDrlJ2yLl6wzeZ/Qsdlj6/Cpz+Rodx
dYjzSxOU+GjgUcz/ow6f46r/4xI4FdyVqt6SeLoIml9HjqThgC5KjfJ5E5Ljs3hKTIbY/BEf0srJ
zOqduHWmui3pjR5So/JfNg/LyFDmbvdP9/ERs/h1+mmhp7/Eever8sg3/7u7t0WCSupXIl0spo4y
XVd9osxfLyVUJq+YYlYGO8Ak682N/aavJVY2NAvoYh4aSTQeUk7I+1Uf37q/mApqZzf83+EQP3xm
EcIKOJCfhzJXGGTQnYCqqJRy770V86Oa/WTgm/F3fwxH/8Aj+7Orr1FCOQgqaV1cNim2B4EDZ41q
W//AcDUb5D8gw0dzf9DopupvcFMNiJTUhnfnEQvEEKjsTArt37SWQ/6kQ2e6u6hB4iyNWJ23hXEQ
K6MMDYtxPUP3BfCXXSkQNzM/XXeD0XZxYL8Eu6EzeX6o8w+7hpjHBMAAirzhZuy9eDoWjYQ7ZDhr
AZazlgolq9uqmDP5EmfJHqb8KstntaLcxROBZxxxsPTiRhlS547dC1zJ09CEkB8CJ7IKuT9ht3K2
WYaGb7fOVP+PnzrH/qIJdiJKVirV+71610/JKVGO4KFQlnvzh1to36iGxawjpRvjkrN1AW+xHmPB
t73kgPhh3sV0mbUaz6P7b9fXRs11NshJiTy5aD7ETvlijvOTtKjjN+vNbZJT+GAM+CIQ7LnpNrl7
zc/6BYBPk8vJHX0rGdJObZphtKo1GQ9JZjrlydfChmsOUVDq0p3ft0jZQUJU4nB2K2hA9Pkcyzyl
cqHVfzR83HUoSdbiMvVzR7/HHpJzxkHbwmPZ5xnN+ff5PQRVTkPLYfvStrixMZbBoJgfSzSyOlmn
4bQRUO0qKbxkS/Fj74Q9xsHYxLr9FNZoW1mHN6BTItrnLsnC02OcUqgFbogr92u1KHPnGcr9FOO+
Ia4IBp/PvepR9BcDa46cJCo5Ep0jqEIG1rP8+zU3yZZ0eS0y1fpD3tOZm1nPsSgCVzjaSU2o7uVQ
7czzw/EvraGlp+H5d+wHz69rVu1RtXbKEeyg9vR0en8Nt3rFhEz/AqnHPX/x7ULf5zkonJfh+RzI
Lj4ENP1FjUrgd1TUVtwDr6wqNGA+lfeATbgHDna07ZoSZauwxCXKtu/x3mg1ffENqorOWKuoenHV
aQDeC3lnk+I9/gHJxYm6l7hwLCv9DTDZZtXl61ED1QP1+BaqKpc0inob/u8kNbDRR6O2DU+hiSaO
M9I8G//cKIM5zvRwHVjNu2+DLkCZ+obmrC0a+CCiZY8OMoOUe5nGupONul2v9/ZCu514MKJ/ClZ+
lLC5z4bLU4zQYJNULJG1LZnDNxEqstFORGEPIYhNZrFWN0TqzTu2vm80D6DHze2G55kmQPPK/2vo
qz/tLZoKZ7QdDR8vwvYsRdlI9KXWAC9OsYVG9gw4nGjm/xuB9lMN4H8pU9Z5W2WdfebJA9KQcGpt
cTBWYFlXL5Ot4/4JDrnkewzm9rVf8jcnC+OVQ8eny5Mri8GPbOvY0RU8IZkolcb4MM8ZzsfJMRCU
Xd2QEml6d5X8qtHvnuevYUM8Qezp2ZIDkrAirw+OVqPLISxJ7rrPjU2prseC2wX9B9EnMYDbgiPP
1uD1hXC7YsnIVEyR3pSpTmS7bgGt2KtFfTzwwOb10dO9rse4A0D57Y9KzN0hZw7dvGAltu3Uu9df
NVCR9v4HGDRUK5RuhwbqvBdmmql+vbK82/lZAYBMUAVF/iGb4qDvLk1J5/gbYpSzXMk88LxvYPCf
kYtTvW0qU05V2odAZ7jLk6vWoGTkmEWo7rzNuGjzL+DbnznVog9NLxoclMtN0POme8IyMEoxr0P9
Gl1cvnJTUJps81rLMkE5pxubgWm9S/qvNuV8dxB3sXpRbkIIEiMn/a8BrYzxPkeRpJedt6KZVcDI
YwUNQMjEGrTgibv5l4LrnXOFdqyNYliuzO3U0AfokvaXhIcNKdM/WrPzLgL6gcyjS2nd1rYjxyHi
OFqwjDEBBqeq/PSgmgRxkMeDj281/x7xGL2BEF419VwCa2eBrHXmOE0X8TswOhNnZYgyaLEGxrIN
X4IcmEPp6Eslqo97IYLCybMoxzCxSlZVFzUwbFQRPFqd0LN1R7pW7nEiKN39xDRdzyssg1077eDd
s3goC2gisCUzQr4wqIpc5sCU6CHVP7RyMnHkZBI56s5/I0DKH9S7vG/zP3pYeRLM7IkGEoWc8eiE
JcR3QuCBHQeDalXZmXdjohSDhD911hNP/BRIoC4Xp+/9d/FEQ3YJaxzBod89FCKJunpYNOJ6WREM
a9zxXjREalCYEhlofaMT/K+XqGVw7AsA5EO2U5D2v1JYTMxtxFaxDfd0KTgWPJTbUbn8WpAVhB7E
BT63OXAI1SP8Re2HoVWwsdLY1f7efeMdNwRBY5Ik+xFwZ1hNGm6lZC/BBTPeHEwaOp9RCTXnjyhf
u3aGpwiyAyKGwk0zQqUBha/TPh2zim59wadqy/kfxMiPIo7MW2L90aWPNcy8zcv07V2rw81BWXzg
9dW/+sWxu51yaolttJhMiYhfR3+nFB2ENVRaWSxsY9ooMZ9b9JKin/1vXN0183uXSAeYEbeKPQF0
MakaEJue+RG9Jz5gRPy8EUbnkrkb8VHqNqlUjIDD8y0YnAlRDYdYqmviYHjo8b9jas4etVcbN1nK
D5y5fnsWNkK4aJfzugJg3VBJF5wFRE8dWMnFo/rg1wfaXIktnqwoMtYJLXjF65s98NcapSQEXixX
Zr6fv4grwMS/6wI7r7tHlsURrAVhkbZaSROlAasEWZW1PsSHl55VlGsiFLmikS5MXkPBNE6YW6Tm
8bImTeb3RfbQE9Od4+amYPLseOCQgMgZIuobYDbnEsu+NZl8NAbTxsojWUsxWXUUnxzt1c7S8Ba6
ZlWrzG5apmxInCkcuz9KLW7FIzaZiE41LNnjXJeIi+ZfVLZInsHDdxURmirHDaGyOAJnU+YSHraC
JsFaUTaNixbe3G6Gh+EBMAsvCf9IGEqvxCLBcm4DLrIrwnwVeDoJbHgfW9kIDhSry95P1ak4ipxF
z0TEpo0skO/7WU5HrT7tk7C6VhBgayhjJHORQ+BMEurIvMeHOahg3FIG9T2GIVSoC7LxbEHZoQNE
LuAnoPlExuSxe+Sv96OZthptSQtp6eomblmhnCYei7TXMHHrxrkVJbkT8EyEGIm+8pgm/Co/WPvG
keC3k+P4C3XBPbSzmXyQmNoJrli50OjJ/vjZ0S7MZwoFeeR3zrMA2fZ/dwrBvIfZ6zr6J7W4z92b
uywoZqZ0OD6fpoDKcL5YIu09DmZSJszOhFwHeM+uBCcuKsCn2El59+nAo2MD24T+w5ZoFmPqNj2z
ngSaQPljOqhLH50+THxbr/g+Q7rRVmAztwICTFc40YGc4dn3o0miD+WfEgxQCh8fr7pvCINfMnMj
7EBO2VJu2IUJW/kQj6WP6E2pj8bSB+yuQW6Pk+S0WbUmcb+VMhQP+mkBzP7neFSswxjPa8GDHcEU
AxC/9SH9N3hOtRcYF8ytLw8s3OD1G/C1774zjenayE5tqH800w/NO0Vd0ITqgObxkGjnB/BomiDQ
PjCCB8DdHGBrM/PTneQoa2PLEKB4yrW1oZ6L43faZ8SeqxPwzQctVriBc0IOQrlXljDBi9ZNFqd6
fXwqsnDLlqtNpOu626mhWBmWFE7sPsryQFbv4lly3ptg2kTkGHsvI+dXonuTH2AfbfdeRmEypxEq
2a6wvacIgtEoOpjb8Up8oWAbCtV+lNarJj+mQqdhqpIRwL0NYHDLXJJK+zwaU7QxPpfi82EZWOUG
Bxn8UMQ/7yAiGEO5JrKPz1sdXk+KHLX2sOEdw3pdbM30K4ttQvKX7e3gTmEtweGUx08GMFDTHy1Q
Wq6AaGODd8/XBiYiKBzrMzDUytBtvAGOWh+lhqEGWg1GCJ383tOtvfFYD27imIQzRZU4qSCPCk49
+Q6JAbPpkeTwuonRBWg4hWyzqqPgZ8XK6Hw3kHKcGxrhSOcb5wavgtrWTek1ksdBpS2Xwqfi69Ju
LsaAzgimwPKEFcwLNwp/LxiYzq8kpOq9FY5xmn8/dIEbxN/JJH49FWZsl4Svltdp3Xy13PUc4JHB
M5ImFMjUz9LaXPMqkJ3ONsqcGtVLTtRf5RNmJP8DHooDzKO6i7yDr1HK3DMArycHK7/AFLPm/CnB
rM3tcbSGIKrGDxw4jjjjkVY7WvGioMHeINPLnDGWF9uiyZ2f9L5T5EGkWY68kExUaMfAJegYTk4J
6L4+7lA1pnUbnM4WT0G2oJlpGZMnzkBZxnsQ1+TsBMtZvDayJCZaNxR7K76xj8CJpFXUlKgMEmZd
s5CzfPZSKnuQaOWLXpNjsIXVueiJkscIRHFM6TrVana+sessgtRArK2U4bmcYQp9zVXTk/EEvhaZ
L83AZwm06JXq8fIRqnJfWZea3gTUzJew8/PmwAr5qFzYodRzlbmu3hgWTiC2xeRYvAuE432jnTCo
iNnsZJICTo5KXKwlx04NPq2tDezq7FBGzg+LrVJ9JlkPHj0RJP38/SLV6S3KZTZZkMGJxU9549gR
zjdkf1Nkg4Z3jj75NMnGGe/PFj5P7jagTqM3A26bEuYmxw+aT3oqmObn+4GlmlR3usbz0wTfunsD
kSGQyJyCVXQqdruLFdeo2MLIqXD2X5I8ssZgXySqy3QZOX4awXZ0Mp3SmO25Emi2r1pTw1oM87Gm
/3wsj9TOeF3/9XgwtfPx9um/rxzP0ZpH0zAyBraMB8NcWmz9uEH1DYOUQd5u/I4LWarBcI6fCBdw
MOxwVSh30VadrN41Bw2kGBmOoHqWJlradPVOHDDC6prJFhpY9oEBgJ6hyZHvAOl5Vw9tUb8GXqcu
7lU/FecozTz4usnGbE7DodbihNm2rk3prNZrcZrIFH2VHQtaMFxNO4dY4k0eueeaq3oe3nE+wuGE
zVf3UJJT2IU8XuWRcDq/sM9d1cr6CA4i1SjUkghKCCBspw/gzhZTbryxiTj+FD07yM7LzG/0x6Kl
ipjibEoekZsgkIEhIindZq3ZcbMRy2cljwMJf4D4YZPmaUEECgnPenu+g2uh0QvVmKtFEg66kng2
9iEtj5kCYFrLS3wkYF9HBzGTmUlfZtcGK6NKqBn06h7zYvERKPiDCu7z1qAoBO6uVuKmAwHf2/IF
tPS4Oh4ZSGuEfbl588c8+Eud+Mjf+moKs0F35AgYTnbGHM76a98gs2ftXtPe5qcYj8vPHUJ3nI4r
qHPg/ZImsI0yH10ZKwJzrGRyn5n7oMccJepOf58TVS5//3SXHnPjaY/hX7m+LCqmvBbuSeSP/Kol
aa0ybwT/pBX8iW8ITESRteaCYqTuRg7GMtwzo1CbV3wvKUssBHPW6l6XKFL1+C317JpjW+jb12S/
A9BFIhKZJ8n4BOjjI5dOOMgRj+OnM1Vgali9wAV3FVxyHFuOH52XLi90JwloX+NMtC2SVE/Vrkdi
+R8eO/ojWFcVNgARFD/CU39oLCw2Gruepq2H+8oy1q6zZEtd3ErvMMPqDdwNpeAdb9wniVPPOwGO
eZJFwyIHoZu6+otnWm8haYR6cCRjsb3YWvUm5ug3OiRd34G6i7hcZESMEehjTi9X2DscjBl6WLHY
WGhXU8JsCDj2nAKGsQYr1yqAhSiOTv45P7F7g3C0DzEJh7X8EU5+pgy37IV7Aj96VdLQbaiaXE4p
RSk1v6xLZuhYZPL/fOJ7yXO94kIHD0NjZW1SQVHBOMYR7M8TVqYpJ44vykuj6rAv2qy0LiBA+3zZ
/srdKJ145TnP77rHnM7XLdnpkOglBywVcUwc1/6rNRSi16AZ7mJ6DTSZNy/LaQuxrDOGxP9mKh8j
o+JtfZdhypGlAEOVWQv9ma6CD8MK2v0b3tINnhWOv7bmWaHiNv9Ii73tdnQRhCuGmWmehfo1AYV8
RADDDdjWHSrLdUxQIqSNRH33MdYnIrNLpud5oIPqVF59fvc+gzINiBFwO6r4U2z5mwOK62Lg6g7Q
wVUCc0FikT5O7u4Bmgw6f0366pZi+s1l/xVJh2ocn9p+dKGEOKTVY9udff3S16zIVK85egfkiG36
F7zo65QN09b86RuJxmYZjc+5VgSCpnzC9OfRm4cafx3Q1rusMZpC0vu45iJS2M789htX7MZ2QsYz
5gwESl8Iv7VHswx4mHLzkBckZDR6qw2iOni6ysfSnsnNIVYetVc8YvDG/WajD6OKPhCv8gQD/pf3
rjduFZA1a51Mvbddzp4ZusvXA4LvZUoMVz6iZ7LfC/ryy21hdcoWPIzoK+cHNPNQTFEF630U96sS
qMMognWgUBiJ7M9lh/yBG/+mvgt5X9Rztg6kJkicsLXZ9HK8RN5MN06jwFSVo2G/N5QMO5FCRkpb
3Z9cfGEfxwCsHv8V/7eFXmr+HIASb5TR5YoxlECgb0LUBJs0LzrvdL3SBeKPA0o2gRx250XfyoNa
eU42oJwAQqx2tX+0V5el03X8pxBgoJqwvlCeva37ol/sn3cE6W4a/ZfC7y2eYZwAPm2kjkBwM/DK
v1b2EMYtluke8MTCWBb0wHWA2FU+S8hDntPw9oDbXwRtSEKWaghl7ypD7P/rmFJEUX421YbMHzLI
zuQfoo+RodL3Tp8NfNzwxQ58b1tGY48AkeYvIc5hCBzdpJ363Gimn7xKt++4/QlHBuN/68Szz9VE
GA6p2IvqZKPGhnsvbtxzZAypteWIc8x5/5eV2I3VrhRdurlaNb1xqZJdwrk45f1qZNrwwZG29Le3
0ntlyS7kvJaElIHoeEZfOmnRrxFcipPPTNF2hoye5WT33fyiTJx92clxa55/hfa8dhGyqYEkoMEh
9uL7nF7sJeiLvWotODc1hyC1hoUGuRhvx52ske5bz5paXUSm1IlTpOjsXzSyK/B9s7XEtBD0H6+n
/nCceoeNMAL9/P9MXFj/xu0KhCvHmkQ4HdRrgpJJ6wVl+x0q/T13833gvQmsLavI71Ik8F4d0PTz
2tDUoMnHtzrJw8n5xCDfVP7G5WvwF1AfFTvhehvqC/dZys6P8c7Z240xf9kXDlorXES9mPWty8qM
aKEQE/V26R6kjWZnx7+QMladxestO+K7+CgxPgIbeu9tL/+qKeVjqsK3s8X+b4sN90n5V+PhlfMC
T1txytXhOLo+B3UcGbHrBd8bpn+52W0xaZMWZjc2sgjuV4bsCByvcUc+SzDbxtnTTGovTcbl49Mt
8GkJG3+4QeOeGnJv3oXkVahOmsvUtNwTxZofuKuFIcDja6sEjX0tvZTc2G216gwnxXqRLhw6gkkV
eRRWSNQlw0IXszY2MwP3Weep5/YLWVYhEbVEjj8nuJqlSfM1foBprvYfSS4wFIzKOD0ZJLUR+vzi
B2ssKvyIJh3K/SD1gaZRAS1HeKGBvkcl2esEzPvRbCYPzr/7PXUPJ7Wr6/8yQQD/lGqaBQfvtATi
Y+DdtrxJQCsZH1o5HMJ66fj63SVs2abCwZTHEmAvPL02XElSlrhMNfzarK1cz2RQnG3Vd7jx86Sb
YuPjNFlRrcDoRf5lFM+6oVNA0PThJg53q2RcTlVYNMSwum9hhfW/QG2Q+pLLxY1nZychWIpkS8ZB
VZeWMWAXCRvZusKNB/zn5I9OF4WkWgsZxMHLus7Uxs7RaSrrvWu72jfPgcgjiWuHyxBEEqJhYlGr
QBeIdlrqva/mopQRJo6a25Wfm3LEjKVmk3lGwlqR8cAO0rCLrZT4Trwp6aIIHlpz0upnefTbzlb+
xK6CdUJZ9O6jjwQVLlOka91MgBNXJTwzeX5aZbiKZHgWYUMOlNJEXYKzoQ9AJaYqlK4DynHTZb08
Pg800mUrFCMGXO7+nhrVVkS/eXZhUhiCIVuRL9KU34NvyvNFzeJ/rK1pIP4mfMsHDW1szKlrZIaF
0155Ezgjs8rRt0SI8kDCpQeE/I7fXVKH2VCCrXX4IqZw9YoCaxio3nO/yNo/BHLaFxyWT8XBIgfM
xhjhnHV4QykRU1XrpIQfwfMYC8z9twbdwUiRlfBZ419e1sZqD/UQ/otHX1BG2TwMQd1N7pAhOCkw
SDPdoFSscqg4QXGvimVY6WWR8clWiu85jRBiaK4yRbhkbOWmHtjyDWnDyvT22hDKvoM9hllVycVc
fLsfhirbQQYt2T6znoNQXH/bSn0GjHILqCp5Q8Ez4bMYVE+/wpKBRKPlb6/zir5n279jGsSXbpEc
Elzy4yIVB20nW+2EffnsjLf5COmGgFkRL7eo/MumlwzYptVPWOvwRRaSZ1nuhcocCUWskjFmP6H8
Ib0p2qrhfFZSJ+iCKRmkzN5HPDFPY4Vv6Yi3nanOZfgRK/o8UmuqKeA3VuON0gOIm/EM3Pb9aE9M
Oa331I7btoeHd7tuqExMIXnJavD0Uz9Dar1XwlFSzmkkqjgmHc9hHx+VI6H8/REdVHkB2PqPkGiF
SKM9WTJP6tptwXz3AxLOMF8ooT0Dx/bPY0ysU7vBtnKYNfdOKWI+HlG8DQTP
`protect end_protected
