-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K2tadPvTua3y7eUB0r+2qE36dLEUbDBzHsWAykkvHd+XuwkAzcFx8UyRinUCSel4d7svOdhGvYfT
tAP/BQxlL+ywAgHQkCYuDATrXqlZeFnZD3dC7xsWs3uLZMLr2z1onpdqQUbCIH5OIraMTLO/JRu3
dPN5lBfSOjUwWEi0kbNuSB0b+esI0riSYSl0hmSR1kelKUOxgb76WfQWK5WMvjx5ByuQSMX7eqwC
UPioVHPcXkzw88VK8uzCti5KcRLgBUGNgLID5/ZSlf7nm6IpDjyujsYY06gseLGxcRFyodn2B3P1
VvGES18I222Q+JJHfNeHl8KUQ74nGBRMQuo5Aw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5296)
`protect data_block
IsV0JQIGu8QSlNkaORc5GvwFooPlDPXZlFeJPzgVE0mCcTpLo+e1w4BekFlX9o0RRuruIaOhEsd+
N0NoaI2aMjAleTIHe/kKSgLCac4bpcYQuAkQfWYJ7Acb8wOHd/BUxPYklLzi+V4Mqb2nx3zjcPEL
3Dlf7lM1ys8Yss7vAFDQQ5M32sJ2hGASmmRGwU8GYU21yUfQSCoDfARYiK2jKre4whQ0SdcMCkVn
4xb6590fyE4GWcfZwlRwc/PyQDohsRTctDGCSI0P6bCbFUKIgZjavkLAvr6Dzp36FAE9wFcahvHI
OqpJ77AVj48pjFePFU3cEjzxSDn8+axpgIwnm6pYfA8x/JyQd7FfDv+PT0Cc7QZygujBTPLtubyB
IhmZPdjxYlDZ2VXtzfcW/YXYYVWKZJc3ZakB3QZgZ2BWYFlOFGGGEXy8KYg2uolPd87tESd6s5qM
OgtcBgnvcPDVxDgy7D5EWphNO2C+qoibHpjGhWJnG7jjFZyYgivcvW+b9rLsHAwLEracBFy35dEZ
bZ7VALBbDlYsLQwovuzvrFp3bWBmHJ/MbxT+L9+PLvlHdSgNtL+dUISnPcD3cItyB5eKqLR8agc/
Rl9Q5cYaq/qDCbeXA+p9BRCU4sRQSueWX8uTCN9yd6LZJatjdNcvFyqFX6dIw1pUBlhHyBdje8vp
VsOz9Lg1OMNRAulHPBc8xjUhwRb2CqKo4VQwXZL7gq7wCIVYVL73UmqO4NfqtIBeXjuEPd4PCm3y
ow4dLdTIycD1ZEmx1hJgEHumkFL84+gZHGfBeW0NoNvDQkZq+1eA1m9+2K6evPNk7VcaVbppPTsG
QQnCPq1WNyWLfqVXpMtzvWFvI6d+14o2MkbG1kNNmQt7LjZHnqRoejLZd9qtqry3Ik1ZhLMmb6B3
UaC+fhqCntDW1OgJHv1Eb6tFZp7vfYJtw8VzmhaZdiKeCjnX41bSRpYf665WowifdcYHNqwGL7xm
9Q6tffh/gEHQb4oL/EHbQn48omKTVTzubWA3tQlTVYPhOLV39h+qFsm8QK9HN08DjYZokXe69klH
BXAlmwJe2Pf3vbYp6qzvuwWT2yaMi0gH1HcxTqHmSFVVq5DmdVkNNpmxrRduvmRLtyh1n456q7/l
1HzU8PRFzjiZxCnvAHg1Xq0l3DzzP8NID5y9PmreGLWp668mCO3mFo93wFr56/XggQvXjQncawUB
JK/gi7EWgj+c8bbxC2+6uin+yckx9kij+V4/sUCA2E7FmiqQP1zIb41VIoy/L/+nAinLtznOZ7X1
IIg3bigUUzWg0AocLZXuT5t2dFPBZkF9vyE8fcjwI0aLVPyVpihBbyBeKONkwejjNtfoIyMQYu9C
9IustZN7vOqAPEpufAvJa3DO3jbDz54rPsbR0DfOOpBBNxbYkHoLqTy2YelPU4LqOLm41aim2BKX
1ZWwHlKitJTKJgPjS1EbqamOIQb3PCJ9DXCLWMQGWxU8yb5fvoBWc9OARQ/kv3LXSq+92ZXh9Gyv
1UMnTb6rmduMcHVIeKNGuUTr1DpVkjS1im8qeF1/HqtPT7pVygxEi4PBQAh8DhBz2Ba/1sC4OTtw
cu+TtQ0LLEnxRxkL5/u/jHrl2dq+2mUJlGJULLFLKP5kb6Ga1HXwNZySLzhv69aIHLGWh5QVJJEL
g84p6JXdyVyTk+8o4HyzWj4vQ3z1ENWqOcnwJKur9EM8kVoeNUcD96idssQxawDE3/lOukfNBX6o
ReQ37mGiqabp6tQ9LVEo4q6fWrfsusD4603oZZhqN8mtSv5veKkKAehYJgjoTSlBpZbDV5powTQJ
Kr3k+6l1n7pU6gfGRYM08mlLqP1SFcNMHRUBROcNt4v8yO5rMog1oaVcAQ9dTx3nY8Q7WMQ7OrcP
zR/Yb9G+cxGNmtlAdMDKYYwzbgLviGu0rncrEfdSbZ9bZCuto8ITnXe0A8f3K+uEPagrjJrLHGfC
uoob5VYsVbi9BS+ub+wmVTW9gQIRpgBNoXefRgifmrPPyQQYRtOUcifFFfHWT4ShB3DD8ziJhj80
Llkbkx4Gidk0sS0Nebu3ewegvM8axJoN/9GXeCD5jMDUuDS7uEEe+//no+2/aGr+ibkq685TlhLR
CESkF5DYQzZXV0FPbdLUcIUvtZDNNAUKONVlC7FVdZJ7EU4/beIK9IUaCDIdcNmPWO8YxZwrwO0K
0swZIxZYxuHsk58hyDaLjwX5BJ1dkEzUaO6mwKP2XPJFLvuUb0X388rj9DjnAHYky7oU+ZhTH+4s
X1d/k0+HsZRgTuHeAeRKaQTGrBTL1TF223rdUO1Hs1bHyDliq3c4hMnuZVzXwRn2FlFJ0Tpbj+4r
Ldm8UAEWiPc/6uN+62vlaD0+BrIv+nLbLL0Qyh0tiMkAKtL2OhiYjS2Mw6sQ50l+Tka8OGoNaFmV
nlEq4G/XtPpRKmFTi5ThHPqsKlqyE9Qc7mBeVh37Yd+NvHPxwP2jz+txIfxolitNkJY/Hr57TeJU
sG270TWyylgCDOWSUre+PHW2LjQLp1hx+VHzqAG2/Vn9Iwg8ga3N9QZXpMj0TnIPmSQ/oyL5cqIz
QDI1VmcD9RROVs/y+TT8vmk3aDPPaXhZzie9PJ5BD3rROjrMN/gS7UrmBcWxGZlEvhkKq3pobhar
hHgq3ijW4xRO6gkvIrwfa8vAkoyMuaLZAYkBLDUaDvtHjoPupRWnIg1S/4pdOFzA4KyDzR3Ti3mG
g+XhKhIkSx3Oq06hZK8GV0bW4snWOoVGn65yPzWbq1z5ehOFzPm9ZG1PBVJs7BkEggGJEwJaOHyi
pYEU6DGjRiLw1EQU5iDFa1oZXV60+u6lK/WUH5fyt92SOBvzpw1AKTBeumXKzSH2WZo1/HLUUnyr
Q91Hkf4mgaj3rbgOJhzBGdnnt+GfIKARd7d+1GNuUUG7Hl/k0/mVugKmrIkdYLeeCbuVMzOPbUo1
jI8Q3ZSA9IGkyqCsfkO+Ncd12Chp7q+qXyrvqzXyW5U5k1ay6rM3mZpWDwtbnkLKnZ7SOoGaCF9P
xXuecoK9Ul+1iBQagSh4Ibg8V3NGZXKlahS0iA3Tnm8Ae43Y5S6/S9XryYKmnsgZSRBeGVuxtya6
MYRfTmnD3JA8gZN+7AfiXFaZfs745mY4v3tDVxi32X+nSN4ZavGFMuB7P4JXnwyIPSqtKEkpLy/o
vnPyh51+fUvVx/XW6qm1Giypc/cPncxWm5MVMi8H6577vGt0JK8qbALyGQtom7o32aWt75A+hfW+
Tnq5kMcH/Q4xvSddTxrVBXhChx3MzjEgdb+ylMSKKBKzyC1EX6dIcbRp64kLEX7bTj/cogkLio/e
Hz4IMeykBUaD3tkSIfAYaedocl9qghr6gjyn3azIsENq+DrRBm2uw3cr5N78VYelYszFaH7nF9Ty
4lAjpYa8qJfMOG+S1q1BYbGgecepJH27crlvh9Xp4o3NkLvLLBMbiPD4V5+c08cugIl2AAdxFqrT
+uVnJ/9o9bCLu9ihzTDw+1/y6CxL+2OM+3lv1ybNJc8Pi4wbHNIrGbD7l1Awehpj0+5n9QKQKP69
Z9zmfwR7idIeiYmAbuXLWZfviK2EA/8SdaK5QwhTYj1YMCvZuBKuhrL3E2V5YorNwTfKy1DI2pgv
d9vw3KFVWWZCheUsbycYBuUbE7McxdIBLS1ICTldYbLqiEI+8ydY/gdCYauefuPV5waVUsz/EcWR
21uj+NR0A/OD3KsDDuMCJH+QqhORFfP8CNgXMckQfIKD4/79KMOnJWEdu7rUsZ1ogbHl0odlq4zd
dhVxRaRKx4V+SMv1jTvWGKnX8SJYByPiY2yTh4PcpvtVbZ5eL5aaCt7ivOqXHUb/D6+7XnvZUojC
nJ/Gm5qG9RBIMYOUhFapXdFhjVXEQwR0xdATBTDmAxf6CQo3RWmCgJLySOOoPu+alSRYMLu04YZ2
gNmYDZsa6Tvt+62t0P0idi9F3koYBepi6BsyqJNCzCWTS3aINhuIBO7zkpnDFjBWen/arNbJvlCV
4IBLvniAL+N+Nx7y8Pu+YElKZoDp7ZlSDNbJ+q4afmYxLtsf3JZH+MsliGYEr3T+vgniG05T2vjc
z7TngE/JaouVtX7v4SkKxR9z07uP73gJnF3JQM/p+j8+/S/1mStkzcId4QxS6JZbO5Lb/kIYP3hh
K74V7pkgkCbhyuHmC9a0Fm04jxIgyaL8EcvEN5Asj6AADgDGX+w0dou2eHvzi9ifweLHGj3893HJ
C+bGcCjRxAcy9008Vew5SEM6K4GOQRK7BKnX2RhnGYrtaCZBuFjPypIgkxH3+xRnq1ThfGci3kMo
+EEujsFOOpafqWT4cSC2m6WFzu4i2N3W2a4NqKn6ryapT0qBmm1O4ysi3NtuUYabvlZNZXkCnPu/
FGZovHnem+wkHoty13qTzQn5/SXlDGUs5IhzxkX5KQwUjmOyPmMvKTN7MTIEn70G3SmGsqF02dYU
VVT17YAfmwzB/NX4YJDzCeVoQX/kXLXMKVP9cmcPRzoACZ9+QfcXUcPPktmEQsMN8Bsod0KZnj1U
GvqO7GH28DH7GYEP/QWDEAzy3Re8OiaXx+KApOdg18XuVzydlZhR/F7mjVS3QVA4wEmp43bzlNH0
LV5xSJiwt5bTgzM34SbBfYHdUTJr2Zy6842n9jL77H3wpaIbR/KUVn0JcYasduAZaO88Vvb6tIYP
6Vud9EVg2KOYxF3kFhEJnczZHCtTLHCNOxJLua3TgfpBqBlMJ9SfKn3V1jFRXreZmU8MbaVP0lRC
oZN+t6f5JASU7WMey4+x35JlmgBieBbrEsH/LCFDKuVqaVjUc+FAt7HrXcy0tIhPToUzo1LHASIy
vYdILpljaKkG1vaFqztGSBbz4vtnQCGQNQ0Ff26IS1dW3YTqzObAiUf7BjddVMhV7nn34329tIpT
4dPxo3djxgvzBBrNFUgkfeXwWLFuuCrdz0R1Ohl7koIZrPTe20kj3wVZHKX7iKDdViRnD23Gaxls
F7aHlbzdwo43NxuKKTfjeDXvW1pMjiRxLZgUyrNguChheDeER0eOCMza2OXkegrdU+5SfSy1HUUo
uMLn8kFUkH5dLFYgXoBO/18uOAC7Ge53J9ROWNkttNnq9eRu79UXmDqFvTPBm1M0vDbofxfDr5I1
+1Df/5/ZoGxE0VBkVz+rKmwdB8Ww4tF8Tn4If3/4w5L48EaSIQGCEqcfA6igpQlnaBOGgjsCbIHk
W/Yv894pkdDzR5oImrZSUNQCVQJJYzs7Oe/e1ypgfJ6qFKSOlerLSjXCMIhti7tuHHG44W0SRdmW
TjJZC1489OQLJaqDYX1/QES8rGnG5fjFRL44FyNUindMnZT9utQUk4vfRpNhVNsMBNIJj3YgfBQk
oyZys5fjw0CO016XY5n+NNXpfGqWOmXHtoSTedD8kRj6ElSjwYT9S3FtOWBI9FMkGZJMMuvn9Ec4
l+WMtW2k1uPhQkOlV2AwQWap0Rjy+QvY3UzX6swKthHKKBInLIHfPSCFashgDUQQsFkRKxOGiogA
+FACnhrP5Yy4+1iaw0bwuiTQUoFsXXTMqjcKb8WXlNTfOchuge8x5ELhCi/U1VDDNMqkgJFmmpEA
+cpsLS7rautjguljSPrnAYgkTM1V894ObBVEuCXxT/3r6zx7b9LLtjk/8432Z6QBmw9D1OmgewY9
G7qcar3XkCk2bdNyyXJQb1ppz39iHL3mJxUkUohNqWk7HEm/2E5+6m68ruHB5zn7FwoZ2MBT8LCv
5MVzSqDWDdVTF+STMdw71wjfn07pBAc+p2EyHcKGHQTukNr+uDdKRUxd+Eb9CBUmdPahT8g29d0e
OAL4KhPC8U94kiKz1IwHkHmEGJQ0Lfait5tvrG9wnXT526ctF/35NGhWKT7ly0JQlzCrwmxXHozJ
ADyMyi/1jqvw3sMkP5jbMqZR/DoapWIoflKbHGxSnMXpollt56Y5Jb9OD6uGsOvvrnp5UjeCo1SJ
rSgN1lr4YT8VSRoBkWORZLk5f6ir8oZKPnhmugoe4HK/9xKRI4BeLzxtgDyNgxfSSrScbptPl2eE
J2L3Lm/DE2SkPe0oKzpmUvhBOQwevnisqMi+omUiBWMdUbr+4yG8FhwN2psBUX917yH1dTWgYWzk
UqichUnGIosbggOqTLHqwhBlm8beZwf48p30t9uOkYUSHMXsvz0/bykiC9fIyEquV4zO5CvS6aJW
qRv56SwfOEElHZiELBEMxKdC72ob7Qq4X9GxfA116eMAZAtPsOwW77r5MZK4eAD7etofvOxpseMI
Aq91bgMJRjxiDwhOpJmnzaDUyujrjYOmO/DwoKIbkBB9oYKkqmne3yqHSZJHCzXOw+5Q2/gGXPyr
i+qucoarGzuQvsnFKzErh4Rj6q/8qZsnsNaK3PMrF2mFQGN/6sKdvrgC3fCqNuuK+iT1RkliWB6I
uW8V4Zo4dmWJX/T1xoV7n3pOBeo79UrWdY22b8+ePLfOe2vxRpla3DkjNDbM5pEuPKkVdQ8K80eG
euR8MLzQAN5HQfrycGz+5O0luvaPRggivMDC+csLRaKBro3T4g4KbsRVxCF/NaA6lfR1U/dLsov1
pbS25c3ctQuptfjpZ0oMgmWU5WDDPlDkHOpLUKmBDuL7FWEddO75qQf20ywizlSvfh19b3RjvPcl
BVPgcPyE6AoiKICHKeAayZOD03Ref/p4pGiR2/YZvtPM93KXcPFd63ugp123n0e/kEON0a9QP+dF
ZZR5nPGq/iBZJ/4uvtWY/WNV9gZIp/0DWhDmr3wo9N/K9hfuvNsNiTWIpEhZbxos9Nu1mjipSSMO
a8fmJo+xsXAxIqulyBjFnFdst4wPheoYOGmpLFhcXyOLPNh0RvFVUQUdV1hD8JlfH2GGRg36cmjy
PLUnb6MHq09lrnzJHA6bdfGyuCDOGQhSfDotTKtFNdklnH9JMYbv9Cm63AagpOiVDnnr4vaq2sRz
A67Dw96tBTbzIuKPIHFLKLqGMMdFEhQ9FcCr69y/JEGkoCwgWSQOKJPUiI0EJImLQeac/g==
`protect end_protected
