-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
prBQqjwUkqajsU7lS6ObEUJBrjbOkWRjW2tyInInaI5ydj6Jevs53hzJ0Oc2JMHpj9DWKbvDIKJz
Dn9YhzsP2driIXqN9YPmdIsCjkv7a/d10UwBq9edVM4ofrMwKS+BJoNJqPs8u86gchW7kBh+oNko
+R2RlsJDIasIu8kletyA9ezvaZN6SSYpyhJG+4y/ettAKt8jZm3pxl6tnS4m2YzQs4nFmmTEAGdU
APyV82SXBPIl0BDTMUrUOa4+UnFyhwMzZiUlhn2dx9PnwJzKTRhSzTVEm42UzDRmVsBnTPZpg5Xp
8OzlDOWWwFzn0crWCE8EhJEmmdxpXzwHtBuQxw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12960)
`protect data_block
YTsXw2Iw6cA+Ti3005KVPxUszKq+2qah3Lv8I7qwEIOSTEpsDBJLcF5Ey17H7POjRG9DM2/EYIzK
n1TGlJXwAz47fwyTMluT2pgL/oA6VJfzILSbYdxs6HboeIcuwDsohzYsSMlxXrxdvho/8l+aJYqX
3mKYjZGLZtmPYX8PjMP7vY0VjnzOlPE8TL26xvYXqpTLYER6oZI9pXsOKVxHp7O/MMP1xacAbAmn
EqJHdfRYah9habCe+Sxct0YzvpAhTbwvFRBJIW0qXq0PsiWdogKSSYCblNUUX24H6lWrzHUFIZPy
TF5UkCNDA0VG2G+GE3qMMVuebS+Dm+Pfha6kV7tzLnhTVnKAC6dlS8kzcqcfO1p+5zSL/l9LMO9Q
Fjq8c3d3YgmbF5Y57Uw+EBOS1boOAtfpYAwJzpgpA6b1piPo5gO9+KMm3RVFe9W6X6hoDe9t2djW
YQ76MhwWMEGC9sKYVCG7nVRMMg+llpD02Kxv9KoiTVljExKkEVuzCdud3OE/pm1UOVyhEIu+rZgJ
TktNPc+3JXziJb70HjKINGWFXdgs9X03BvXSRbVPfUZuU3/ubSLU3q+ES+oh0n7LgBw8sfEJUQU1
Xhw1L5W+1Db2ge3xGosRVkNPbcAIDGvMyvTqYJDe0jccqS2H6VSOpZGyX41VYebRae4YU+w9gTbn
VU1mRVDAGysi1yfLs8yd3xsfoN24D0+LGxZ7hf2+sGAFpsP5YoIQ/FWPL00ykAcj2E1lS83Skt3O
kuTXBLQKHFKozaHU2UW1ipoyCGZGDNmADGnNC214h3B0Tpo423rEzMsn92X6aKFoX9kf3uDisNnO
UbEVF1q0tf23HTSLi4FdMCALBvqvr3GN1VynTtDp7gRTWQC8CievHx3nPCSD/SJ1vdVXoCQIcjyr
egUd5qe+JsmAKMhOXUyrDTHILnUo755e/3rLKcZdn6JTJFNw01LiDUHPQoSHzE4H3tNXbOHkSfUg
AN3wWUkEXglOYecThsrqKqP7MdwI20ue0G7on510Ehrx8CyZ4fxMacFvkziDRMTBkvPDhZZR9BmP
46t7+WHDoKbVR1DXkHrcQRIcY4lYQBk6ewz+bOPKyGqyOdLDSd12Phy0eb2RYPY1N/juVBgELGmY
zQzkxOyif5uyonxEO2zucLI1vBwwR3d3MPdsChX2A4qykgUKasxDjY5KkjdaE1tamx1SLuWXhqU9
qHaV6rG6IkDmiqC6kkEn+N9tWrsQ0dhloqPQJ1efgL0oifcpVgfWwROr0iVrPuZkLoIKImLyMWsJ
EYUf5lYum/Fh7gsd69p1lyrhpR+Mzxxxq7XaN9UfzR1lRgMh/2IEOFhLkFJNRUrx5TFJYk/okde7
GOECvwhXDbkGwybHp6MHDaBnPW+EBCSHnTq2i5rzRTrbXPIfwYHEcNmA8L06RCA4WOI61dWqB1Iz
EHmBdC3o6rvU+5tnv9bMjAJ4pWAEpeyZ2lCaLWyuD7W0PTQI2hTih9Ybsgzp8oaVhB03KKjXYIsk
kIRxlvbn9E0PmVS9BHH2IlsePKrbRBrP0t7mQE6Sw4pdftICmmwJCmnbrg5xENnevNk1gXyYWqOh
pI7r5ZNNkK7DZ++QBmub5Bb36UTea2Dzd9WL8Mpo4NIndentnPmxFfIXWbbTCX9dgrVWx8LZup1g
YPZAQ81jCGcp5DiqYHGMjJZGTYa02MI89OXMt4lkpPt5ML+/LnIkAObGWHAwgsj/RZNpRDEvnxAV
mRnyrJm424pZXIshotERVYtx0bNjKPBd2pKL+WBOXyOzpM5I3Kcles7i9R7Gs31uoCpkCw8OoTot
eKiB7DfQLLj+GUz1IMF5O6ozIKR7CSSh1r81s1jAD8LLlPph0/0dOpYqSgFD2TvPseOmoEJIdsqQ
JXz7uUfLRoa1ycKYDUzDEFwoiQ686W2MTpfr85wSs7F4eGFW5iu81MVA9gh+G4u3j52N65PTxQgQ
LODsxytZ8tMlRuP2HqXoD5r20NqoO5rmiK99mVwYNIV8KtL+WLBH1pyDdpmj3m3vDjKUyv4AavCS
rudTp4TRyaZoUguHBdN/rdhiiEaceGS+ThEshDU9Kh7xw+sVla77pQiFa/ltkuUdhZzrUGYcs9bY
F/IRYfjTUvMlJnZI5aYRMnZ8uWVrROhEjdQxn6ZadyxYRmJziKN4S8v4YDNHuHdcME+nQOHoZuf4
yZnb1CPa8tsht949NPYZy60Oi6Sl8JzN4/NjfFGy1TY0SLOG9JdntlKuwypHtx/KmQH56MM70SCS
AO/xnWq60zyf1T7R5/l9bNKR9jSPhrWmHQX8+xj5ASjx89DymK5OF9dg0d7NqZ/wi0XzTxwi8kqL
i4epyo5FMD+DWYbh+LAOaRq40ZJqmJXeyyL28BydY6ip6rd8I4PGwC0dOY0iMsuWmkN6tTlC/Ei7
5+naEHJMnxtEiXyAcNMe5f8oOQ6vaY/dzgE1z+6n8h6vYzkRVp86ZVFcaDUJt1hAnZc2XWFJG6Md
2Vuv9Q8ISCDs4ISXuGA8BNx6MyJI4DX0MfgLq/CdIZfX+19VcGF74ismxJbtZmRQTg72V2LH036r
qtacEoabpUwdeWfXwc8sOyr8UQOoMBi9UxrYmvWJ8lf7CMTxUXJZTPy9SoBaXHIkr/eH18CwdK8a
U90iNFsrHOkQwb4tioynCWkpOxIOdwMBmt67EpxPbkV6sfo/3xmpPWgIHVF6nk5fwtSMw+kcEkXS
4E+ZcdTiUWZ+8rl6Bq5PNuxL74hFHaUiwPC9p/75Cq0uf13vy3yftlQFnuq0sCaELDutorEZy2rB
J8G4Y6R0/4dWQ44EypsagTd1I5ISy+cMaGDzZJBwkx2g5pEtQt7ULoJMRvpYX7T8EJHNTPng5hD8
0AU1BrOHc5v7WPD22RaMRdLbBFh3bMlJP6AMTSHcO6plaKu9Fgv6uqD9To0zg8HFAqZ4shtqo19w
eP3DjPh2OLHEuJ+mSNvEwaSFiRV/R4tKBbMsY8xruc6mN/i+29GmO3GanMb8lMBFHL71oIEODzL0
sEUPDpMH2f0Cm1QzjIzXS86oIAkqZ2luWwwoHaosFqeZSkre/NuSlU6tX/whacRnKzyr49s0AcvL
dHvvs8Rktzag5lCq+5AkK/T+tzXo/7jIPesj/FbaEQ82iTODmf/YpHE7eRepKmjl+9SSRwCEi46J
JePdLUhz4aO8GTSg/PY5gvyDeCgERAkUzV1Xvnt6BSu/W2o0gD4yRvm2TWMqULztqo4q+LW9jfRj
iLDtcEzgiqRtWE2nUX5l8ho9c2XJI9cdkWV2FNjz3QKaNw9wa0ft2WkHt2Etbd2PfDi634q1Rl99
lmANjCJuTS03QfH0Ln0sElTpGugQPk6AC0C4MbF4qLcU0nxgnfY09v2niJWCFZkXu+nqp8BvizD8
cVx0UVxc2SyZ+oGgpoIOUJf8C98mYkoqY1UnJ+rULCHvioocz2M32ikcjeIZX7yb6UovTqEXdM1f
VlKTGm3wgir5vSlI2pvIcUkvxJBgGixTAws6aSO5v5acqLg5sZWhfU57BucDcH36ILaAeCPUOqsD
1QxBxlPbQx1wVP+5mEpKhFizfXGuKTx+V1sY+OQifpmzh6MlAerip7vipyVz9WYaCtbIE/+x9eR4
+UAJ8xETABNM5qUrgQcShvJ6roPXPEgcenNzjTpIN3WJaeNfdLlqWweSjuhsw0oFmu4lNHpqQT0E
tzKtdnqP7YGpKWDPBc2K6fZWdpmDJVPOt8sSEcRRLRFJoqoArhUDasHP5QkxFSu1FG0cODQS6vu/
o9EYleyesurjL2DoI4G6SIa4fAPf2vd7QI0IWpvA5PVNcNMOP23TDcEjLf39vnJ02MuQxO6L5gD1
h3z+3WnzTLCxdynGDX8P4vWkdC/nztMRuKhTQW+JhBn/+57aWIAq8RFtycXwE/OdUvw5KSmaFXj1
3neQgofPjYUq68htUAKWcJyVz3N/WInSpDEf67i/Kcim62Kh6JhZWzkfgTrIg9WO//AR1MAGx8rp
FPj8AgwF5xArI7Rni/VXjhZHFBaPY5YAaFKe5RilYWJ3B+IECNbOXUk7uOl1BJhwm4ioJ6FIaAru
E1pWOf99Ds1o5FX9cGsRzMeOWJo+VMfb0Qnd7QmRS5xlJxqWYgiqTWnqDo5mWFoDtM6gE8/Rvcf7
Ag7onFvWZc9qWuxsou6uQD2DOFzK56KPLr849XcCpZ3oHna0xy0+fZptJzrvgATr5Wt3qHpd+CR1
B1NuqwaT3DZdZZs653M+xJpmYBkBs8w/TfafiuV8MU8rPCINU5o++AL6uve4biXRuzLu5NxWmJ1J
UE2mDYfPAVrg9ghUX9zdmBp3pbW3+DSurmwQHFXngNPgS7zM1Jd6KpdAX/yFxLpHIBWOOWp0o+px
N65y01zYxmyAS9woa5wZHEmsz5t0edDV2pCmlX1aARqnaC0JsibXwXD326zksuKCIkR/crda9J+V
0YlsKjMD5g3z4DL5n/SJNQEsOrnxRDvG+Ay2sXfc6e2EvBZsbPFuDgziSVDIjlKPmubhWegfJRcT
8JsnK/II1+sh2JVjfkoAXoP7TuUniGvd7sn4l1244D4hnWNHaj0sO7wjGCvOGRBaTrTOcjErJllU
MHLCgyrm+5uKf0juQqkWk1JhCZrd/cMJ3CS3CtttvWHFYHd+f0SLzgAReF6WlMW+/NxpDoV2Ntse
MrNtfLvH/TLx6QOd/E1C5aXaY7gmy35eqKdbiKRiwbavOx3ETZ4hmt5DioFzSp7puzvMGKq39JGV
Q4MQ+OHsSqy0l6nOyQFRWI/lbdMbUewb+7EeQyW2ThoBMBRCHeA/IbPnkrJHSsHPy0HeVrKwtah2
UHLqphhQgKIAecVeo2vRBKL1/BjfHGwZiLpnSKyc4teSkwiH0ov59KyJobyD/yuCiIgEcWs3B2tp
xCdhRjjxG9BBlGIQqGegDqgxr48XBXV7W+9Jx+uzfQFMB+8RKmsJG7P30mPRqfqmqwULwepRMdKF
w7iGoskcCcfoj8vsg0tbcX/Ex1xmT0sm9zXxREvmtZ9dRW+K4Kt3Duxd0NW2YjxhZZ1cC+oed1Uv
Z7opy7++yEQwi2Yqou8S4N7DY0Lkr78qcWj8FNN11Kbxa+hTH4ApAjaWhbI0XDuBXa+4WWOy0dKf
qy49IsG40nvtPraiVouiDtQIcQdGVThQnGZz8hwbxdivNQcZn9sNeDZ0Vfyv5K3MTBShTG0bTV2g
7JkTPLun/0x0K9S6pu4ER2c1W7QlIQ9TS5EyWdQTOBnRhT4HO5FFxCIh6Td5GrM90Rol5S9R5PcC
Ce9D55BmwFJ8hDGDGTM0oJMvepBtq6w3fAY39sdKSB6iehWn3bDh2SPNr2of6o+FyXsj9ypo/ps/
oWp3fTvoVSHXL1x9eCZUMV1H/4N9qBE5QstgtfEpHUL/cjCX5V/YPB5DSZx5mqmZHThtRofcZPO8
bKJJyvn6sop9qhdY1EIZmfOckYQSWCYCM6Ariy1GwzL0OtL+HhtjmflPFfBXRl55ytZCEYw16Hga
2TwOHLWS5yUpxj1P2BHTz8DgjexcP2l22jtbsC+AYTdDTQtFn5B6k+PsnXQ6e11MrSzpBtmLPncd
2A5Ev1biHUyBCWYSAxQbpMZTaXBkjQF/CanXHOcTFK91ZPaaSojER49vQSrSGMaWzKPl0nRUVnJ+
xgG28T2ZaiQVOcVcE7gQ1BT9NgWFCboVtsr6OXD3qzu7HTPKn4hqc8f2GgPZHSlfDE79eLPfeEVC
HiucikSaDH9dGCMr/vqSY+ONfF2394szlaKiPd5x3EBnp6iKOG6i/BEBmOSAycEZ3WOIxUG+KeBP
CK6sXQYcCj4ZbKgRytoLgyfa016EiNvn2Ll3R0GTHa7RbCGw9fMSqfWP9mhK95y+vwaca1Ou4bzP
mSMMWQSvAW5uucfPdMbkxOXTUOPeXtrAe1wzaalvEbSj9P0WCio1+8G1TO4/5PnsWYbgRdzF2GuU
rxn/zCIEZ2EBFtXNFFcJ3cNDzgPe2wRM4JLOQXheDncJtXB3lMlmIqtoUhoITsWtpnFyBh8v7K6d
r1e2eJeGYQlsnSbo2dj0zkcgtKRhm50bPZeQjHWoOZS2MbxBoauvwWxxZVt1nQ9ZyAjaD4Plg/h8
RyDdA5HShId7W67L7x42O43D+NbpOicwKRcgaVwZXN+yE+ugfv0NBWIYUWmT0m43z6l+vm0n0D3i
XaSCVcdTsWml1YlNeUHfnZPN0/Pfn38v+AVlEwJVFiolOcULuH8NiGtoK6+cHwfJCK75gwOztqxz
n7kQee1etX4hs5NW3c9Hc3vAKm/apY1uwt5z1EiJ50yXtQ1aqmfVAxFKKYbED5Uzd6mkygz9FrSx
zeqLjL6aUxTz8lBMV9BPiRw++ERGWuor7sRts4pX1Gjq4zSaGBpIsbfeiGSld4ZoG6jsM4b9YqK+
FAvts8JT1jipKIJWYH/OUWi/vZN4c/xzDx/95DVzdG9FZXn9k5yDbjxvyRJ2gKnzbvOlbmh6cHGr
Vj1hqBGpicPZTcHbChClF8PAq2jCIe5fHckOsIusMMpDex4IQ9rfQ+uzlbVG0DhCPt0fPcj3QQxJ
n7Lfp8vhmziUNb+5x/6aZwL7w5fNBKzFRDbhnES8F6QDl0l5KdqWkwEZbYUjX+AaTmVuAFkVDE82
EKEVt5wo6baLYPCFByPS4XMRDWEcBYkLfQ10dZ060eEYjfGZc4CzxgJ1Hu/diMoH8qt9yqVAP6j7
3bRRfoi5PxkRsubXux4qQVmqTzG9WYLB24Xpm2KTrN+OHPPuyFaG8hEIAd31LgkLJt/PDuCnIFHG
Ziu6N57Qos94fQmbMqPwO2EYmz4CEEGreDZytAU++ckVpCiIfS7XJWgEgMc/FqSpH1KljHVqZWsV
TFG0aYX/5BSNKS7lJ/705Yfxg6DNEDyC5yVNxIt1JIcij86ZmYEkCAq0p11uqo2h7Fkakl1Rt3RN
x6yxqzljqt6u07z9N2wzJhnPD0w9P6hQ5BygRbIMJ7eZOGZBF8McccBjgitrHSlXJmSUfdbXv9rV
lnJSQDSFe9pFPUpMhPWuSRDlPLFKXtgr6emT6NN9KV1yYxFcuZAI1S6e0/v0PCMxHMFrBKA85WM4
Q4CnK89FBw18fSDGF/r3F+++3LBZ6CyizC188dEmI4/WWLEU+U1FIUWDgXny8LO6D+BWWxN9xJi/
p0ZdwzAfQiOPn+TuoLOXIgjXhX7A1qb/+IL4VqknHum09ZgEjfP0kRupUV9zBZfJFNF5A7n2e+ey
FTh5S6BOiZGpletWFWoWLAbzA9BNSKWDHHjA7WiV9jz8ZTF1HgjrZpGzHhm9HYXvxg/4MZBggCxm
1CoX16TycQUFN4BWQcolseVJw/1BKhF7FjrABWZ2fy/q9kgTzvetaRx2tgVkAYJOC7PJIchYa3Xz
kD0NYoLQuWOQy60GjqYW+0jEbPMWoG+ve3ylkW+47VwXQMaxKVTzrLtbDBvhWme6lMYKotFPGjTA
LrQsF1kxjELd5BFBR2cG9XZbXQQP4rDgywAb2aKrNoUco2qB3SJeDH7u87S0VuNkX7qgERnu2vW5
wwKC4tuRi33elJ95hxsmlplnhRpYIrDKN2nYKVaRUzgkh5P3ZtXI3iqLiUnLdcvKprIxWLiTaTgX
QhtQeXeoG8Ni0vAiNht4PbPBnvcuBQmehmjIjYsiU4y3QbPln+FEOfQpTzdSgN0wAl5ZI2tNv7kO
DzzTm00V1q0GX+UtUdzULYdLgnH3QfdR3vpSYUi+ketUXKhUN7WcPpGi3hJ3ZY5AQlGsUSoBfTAk
c7UHp2mWZ8PkY5ZqCzilYhk4baWI3ptKkfvFSdprceU1w792kc7Lr15Wkqim2aTLQw8Ye/w+Q/SS
fdU2dcv6RHdnLmrcTAJt+SJHsCRkYrXnpHG02Ed01MJ4G5pQY1qB3yKalOEFjpHS9J7pYJ4/td8m
fPG9Re3yb7dByt/ZeU1F0PUP4GTOHLXnULwNkJftmAwpkJfrUhuwmdiKH6th1xUJTONrVeUTqLqQ
ouUTWukhcs5R2dj9Cd079cF6WQptd1CrsOnWglKNFzB/JOVFwsGSXsCt1wVFDQ8oqD3a89Rwu6pj
7gWyH+jGQXGBLay+pZRSauPXQikdi2h2afL21PzxPOWhmgZdQFUFHD4F64ozW7BJalcBVrOREQJy
Gkn4ifXJJqxJgBxg+vUxhcBfals7RHeUfh3USJYRKB2nwgrIIrEc7RdUNnSCIdtSbt6YE3VSI8wj
Hcvdgz4W6O+Rg9x5qwOpClhY0dyrQRbYmtcidp/Ps9iWYXVc8DEEtPMF8ZPFI7sjvZfomv0czUnr
eLwQD9WlW1ZAkk6HOHdDNEtjy5ZHoh6mIP05Bdz8mPp+Daid5Gn116MaKcfpVUkrJXKuumWJFer9
M9rmPELch8FlnwoRy479stpUvHRCn3+JbcexhirIJXsJer99hkl8lLpC3Cs4k8ioMEWXckPo7d/d
ybryU9u3OfU8Wc+H3VseuaF5YB6RVi7JxibSHWQcKD5Fqwb5WVz1xkIz2dPsX1QMQiePbV1eArmi
sSvYKGmjkcf1TdZUliraNcThIfJY4uLmAoV4P8UApjd8TVK1kcXqwHxoju5lUt7Qmyug0yqP5Ker
50Eu9fsrktm52+gYnG/uH33ZLzsTsP5ub5XmURhBNxo3d8AMgm+sw98Cf5vCM6Bkr5noinfYXGZT
lQUIFYvw+ymKBblWi3j7zY9UFJa2PGAXjCOo+4JnPaptdbpkbA5QtnbD6Do4xE1ngSBzAk8K1EQa
SLX28XzJyhYRZVuIyKImcYIyvTN3h4LLFwhWNU4qp1ytMqcvFGc6/RKv9pws+2pog59v5h1S3wRB
RvMSvKCMKtijXpKLIj2oQDRdlCJB76eDfOmD0RyCzJHYxjJqEydnwcR46McycqWNF30jTvSinB8P
+mDRb2a8sTgys4mwjAA39hzkWY/hMAidkMF6zCyFa9aoeVNedVAY1Y7vd/xsW/IlP6YU6WkzWR8d
3vy8a3dbl6S9R7EUInaz3ntBMCJEeCYuvQvbRXIBu0gpqiCqof8dK/fp+eqjVF7CmEdKgULGAUiZ
gBUVb0c31WdQTiaUttdxCVK3CCG8IosMip3VkCYA7AzU/EtQZPbPeQJMT7Z6c/Hk2ksBqmN2LF6u
g42jioel0uScXNd6ye0mYnIct1nYtTzzuS9XHRyzQ/qMBg4ubP5MGdQSYxRpdjd20L1R9dsVLW0r
Y4a5ED/QXmx1wGQcYRCitiPBY9Sg4PkM5C1g9g1X8YMxfUkQnnaSJ7KHDiJKGQ4DvWHQDiHrYwak
6/dwXCvBXGAg4MG++BILfpYYcli8oIxluLKMDDWw5KtiefRloDPwAQQbfL8e4yryLxfLUM9PnssA
xI3B/lMxejKh01Drspm6LOFBQsiQqQDMpKo9olO9LgVnStuRedBle1HR+mOexxN70n+hh3gdy28e
xANn1wxzPUi1ch682jsoBYT70XLaNXyT6v8UJz7SOFYCNqHC13+ks5TaxmQ7fpE6V/mPmvAK5ZIJ
l8Qs1CsxwM9HyvdP63yuJJqoXri4bxElddHaT6l3FwvKJ2nBqayIojKH/qmHri6Rzrp4K+08IGNN
bmb/fW42CIObRHiUeDN/0fm4R1qcp3YfBD3CFtQt8J9bKS70FPbg8qa72jiwrARuoMuv/gmok3xR
Ic+7UhP8ficigGLHq8GEMnvoTe+2A8/99uEJo0A6bZEiXSONvGj/goTl/cLLnWkERkAsUeNbQEib
zPHl92oqYiuv2ZA6bZ4xgH2d4+oCBjDmqU8Uu6CBED2IvpPQfDC+XkmExxr/ngW423noXt0wPs+r
fbeBdiOeyNwWR3f24HDoakdIZkjnAlDpERNBJwk2Tv5YKTRYEomK22Q76gtYQTZeo/Z9JLMoUAtT
R2ZzetAWKINiS46ZduBllHghVrEDNSJtSiMoCs78ZDLE9q3+Qi/dMPrMlzKV8pezNKHd0q7MYwiQ
AHYEQAGY0xGcFaLWqz3M7SKuNhmYnrBFK1349z3IkstqeEjdBgRtkZ3w+RYGWy+0aI4YYKKSa5O4
nd3qMvssLNW3gZ2se9MSLRySYiUmHd+0zm1SGwFqo2OHYIVfc1CPFaEOZHXwti0t9HQcTvIaNJ/d
P4NN3fhas56KoChx2k7cyWp1tBSk/5xKDhsqnRFC+y7DEIE3aZDIAngfRBBhftYwTy08n5ZN9VeY
kulIbsE2impoDHKMqUTe96DkKonTkSQebFZN5SSw4B6u81rF8Cpz0bIJLZr4KpYuRU8B/ebvjV39
qvXLhW+582jfq0ATvm7iGX6aB/iV7nT4Dn8TwasTM6AuEo0RZfRhOsUr5LaNsaBclrEK87IovBNN
T9Go4OaRJFp6GmN6o0WL7cfEVXRW+FlUqetwzgAQFK7rJ2LdF5aODnS+JnQqu4arxNboHd2bbKZY
KiCojJBwHIOSJd/aWYNNN/tCx8m8Tm/gXBAjIlE0KHkzFSa0T0OYeszxEWjyKVXu+p0BrIgVX22w
n4ytR1VO6XNOco2P1leB8+HKxqB0NjiliYQscmRsBdwAtN2TIm0qAHKwQRElcvnOtDrI/OdpLYOr
0j9n7zuNciUG3+iwVb/nh3KXAbfw7Rn3aXl33KkBbFpXUcJKacZnoKBreJ45uu9RfUHIKqzrya6U
39aYhsnJGoiiBa+gJ+9tvhNOIZq6DM9q/52bx1RTbFCHVoKf5E0T25XzWTc3Enzl+iNCkMrsx5Jw
EPdmoffw6zperj0xRQbUfE6a9khl33uvmd+2RVtAk/YA/wNM0kxcqA28w9wdPSQPMauqoJGWXCKD
0zfvO4TTw5205z8c5Xu0PCQflCA65rtQE3FtV9vmgCm+rTHdMIzxxjbH8gUa9nOixFc7WvX8SD+B
9ojGrn9E941eroe5Sq4lSH8KE6ym0Co75lo29SKLs7AUr9C6SWPXV4Z4ck8TUbw33yfy4zN2UtPn
irkyG0voIkoZfp46JgJOENUWlCZ5Y17xnVvUbsk2BbTSN4eCab1l22p/42hIASjVfN1Q+j7nnRWX
vyeVojQj2KI9cQ/qq2MkfPEhH+BJ5dC8Myso5M65TYUKdpeZpY3mjwcc3SLcHT1T8IkGDer9KvHG
IJxCX16NlozgIS+8M70iMvxVdvf/NXaDs2mY9szbjeh4AxzSQkRJS0/OpFiUCavvAk/x9qqEPl1F
Mdd5H2MReI8jb8TQ43XtgjDUYrOGqJKC5DfdCJB6ASgJqS5pEhCjLN6SnS2q+dqc4CMJUpHSKFvs
SHUBCOZKEr+JLgt13cQArlt1Lvt2mTjYVWWOjzM23CD0DTZkB9hFRx7EX+SmYr5Y5SJbKTJ3OdWA
JGqBZU0ceJz+aL1mHBu1UCjZF2P3LNIcxa1J2CFdH5arKDYpgRsZMEWPKcitf7fOfgFoY9EVfmSh
Jbs8N20SyY2A32ily+qz/BLCzwPZJRGQCFgchHEGwFHRTdaCrbuvZtZ5sUDbO/axBalz2UwOiAod
yG8TNLlYBxcubbFdD/yr9dIfgT9ufiXdLKAVSuT2gBqLuJfZBSDfbQUS2YZdg5woBT2ZDn7YtNog
wvXmk7vWzwX6XX9zYJ8i94b/d5uU0fkK2b3p0SATOEx235S30SL7IH9YV8GHQ8mT6sAtG8AK3aqu
3fv2EgDWkk1dU1YOlh2of18rdnAU+9qLlO2U884ya1sWFn5G/Ayt67gRyfFxm7U1c4kXbvSRpqGT
OKm1XvmLaGyk4Jur+KFABGT6uVBc4YSNICi4lILJ+L0Qv++K1PT4QPDnQ5SRtvXa6Za8vp9UnA2U
SA4Kf6YscR6FEywPtNfH3al0j9/Bj95JYrK0jQebte0OJkXwe8EfNd8PKx5jYBE/bulkUe0s9A+i
TvsQx7d6yZ3ecZQUvcMHuDCX8UYI87t3c0P5FghlUC8OR0bJtSQ3RnDFyXcQTrxvcE4xQ7Fr8REV
GPW0Zbm48ultviYcMnDo9516uggUSgaROuRvsLzqDCWEw+TbhC63a1JDNzaXso4FLa3sT1NbWnDQ
UqT/u0L1S6GDr42YGi7cCpwdBfc/C+mcA7XQz/ClPUGK1/TdB5HywANgOKGe2+9M17pzFDBTCXIC
oI6X+vD7I1xlEjA36jseO05NbIQ1LlaE1Xd3iO5LDOFpsgST8UXbf2aimitBE7uEBiTFjpScRo19
kdaUy+oquR3PmyeH0MQ+yvFGEFCB2Qac4Xfcg9U6tmHhmkGSgqSzmDeCIpy5IgrgHcJBarcjO4YG
LmEOyacCWKWt641iIzK2Qd3B0uOWEHs1BCtT2d5PDFsgkLj2Ym2DnEgEOiIC6cbAQqfYkaratoRO
AGZX8uU26jik+62uVjDQjKXdbdbXqlDM/AVMcTFcBgU9TPkkEdSubAdMYYywzcAhfgPFh/FO28au
trOAMOUFq/w4+GvbhtDtQGOGEWKz2ufaDQGPkc7wk2gl9+bKCE/ROqnB5KD8mi777jCoOU6Uc+7C
J0XtDGISsm3RXbT43B/fZ01V7AmvqBbDid0SQAnhojE1dSjESFKwq77xQgw7ppo0d2T/o+bNMiMb
l5HAfBA0TyADhM+ljU4EKqgEWeObKn3+E7Q+gY+V/gxoS8hNWIWzPfrlO/gLTEun6EkLSOY1KgDP
Ju7kxUOkGQaQa/paQJmq4Rk9MG/BzrJSU29imhQHUT3mJKHCsyAmVHGmAWZ7mvYdppQ0CPy2j7b9
MqJDbphnQU2JpQ475Rb/VJp62UiZcEc+vNW4/uJZBtDdyH+XOg2N/MN4M9gQXXs2lMcNDaw8003C
PQZ8gr/v0qEqOYjyACuSGy4uJ/gAOQySGSBzO/Pra0LU22fej/HEZnfKNOhxPNlsZ1kUjo6PHmiU
MmFsbFE6R3YWkPkk6ITJfXxjLV1JdJZSSW5Ytnwqtes4bWpsyXM35NA8iDg2Rsz0Mu13EHgTW246
WKNU7rIvilorl9GZjHD3g/GKa6AiTLNjqBXCSOiHU8OJ7ug+cq9nTYNPljT8PtzP9z1yfuvwyweA
0AmnpUbNu2Sc4EJwHbYl5L2izC2SP4/SgdSq3+vLzz8De1fE+L02GaXuzvnBt0yC8wVbIPLhqhMy
ysZ8BW+OptwDi4Va5IEfoE7amlbsqDLRTppSFlyGgW1vmzc4OxvvPeEhyBZwbCcXIh19vJ4FZGXx
dSvth3r8OCK4VMl6abvFZWY5IT9GjbdosePreP71SaSMfEX6kQtjEs/+5AvsfDeFyrfoAQcb3B5o
5qvHiGI3RFFLCAwY/Ma99Mic2A10A8miQCLZhzzBZXShIbFdDY2PNhizHN9XCkQE3kGQ/qOTuJ5r
hbURS5FKUinODQY7LSg+0fdMbG1kFrsevJY7+9fqyxHa66qMY8o1Fl8DyJP9LvgXb1KzRDIanvIq
1J4ACsdvpH06PEQ0/z4feskjSsIjqK3vETl46NO97u3AmGDReBBsOddpWAfHu5BTN9QSju2IKBPX
ojnyqZ2Wge+Qt58g/bVlp9DJaEFJ/t0cW925bfnoMNjryCXLXyYonYkcvbQvkSPsrNBscw0s8Ysl
a5u++6jtzo1TbL+lwnG6kK+N2yxNXR04mkhfIxZ/t05/Xq8SoKq+gb+im+1FzAbZKwT757oTtoSQ
5/VRx60M5Qe5aAnSfPJ2iSaoy00Hi8KoxHPFxs6YgVFWJsVzgipUUhyRwDudqYNayxMkrGPJ7YtC
6jMBpzUYLR0gj1PwyLeKna7iJHJeDjfeF9wlck0B2vT7sI49dWwON4XoTpBadwaaooBYs/AoaOpP
rJYLqysdiu+1Zc7b0rWal/EDtdpBoFvH/cXCaIXeN6QJ89M5Q/81OfVHMmpjkpWmDpa68kGNz1ik
fdyoEvbHqxX8szB0ViDYOKstN4QPdpdmL5HZy8cW78UJhzFTffkkG6Xgx6w2vpKfuGsD0gaWc2jh
8zNbWPvoaVlo7xJnovcaPX8THgPAKXMMp45Z5cgkhiQh7RLa8jB5CFx/3uwVZbvrDu+9FxNuDFWX
xZ8t7EOCGVbtNIh4Q8wSa21PvobsqkWNTZ92nwwJjwrxDfMci2sagWuW7u0wLxOFwvsvFrr6bCyB
6w18I33GQmTsbFJ9AZLtV7D5qcQTHcwx6lcynO6bJfhyCjhT9Ve3Wg2B8baaXlowyNxI4lmFnk3O
IqaurZEHZ92pReYRyvql9YSu7gexsySPeP6gB+rTkaFe24UNlM9Ct+cLiAUWxFYJ6t/7FS4/xXJP
d5j9+s8copy8tFadLhMTH9Gj6ubEXnMFja4QMFLPdWn1fi1Nv3g1xASoI8FttWhp9d/JLRPf4V4L
thjF6hWlZuBmtUKmheS5cDGbPJpwJuF2NCJdhzX5ZlAzj5mt85btRpglL7gUth+KLI+tDmAHBA/4
AflL2ZG3wH5l5SgKiel9BOYVB/wkJJwr57WNjJElGFriJspn8cELoauWmVWEpKQ8mHy+JJ5mfd4b
OlyKyfhhGh6EJTSo2gSegOyaH0pf6krVHTH1iKmPqpnGHPx8rToeQh7bPv/uzqOiWFYQfenXiayO
9rrZSMuVSWN0upn3YXfk8Jqy3X8uZxL8/sKu/HYfYN2dzr4zsuIptQ87kBlXMtPQNmtXLBq7PrDJ
ywgQZUTPMyrPP1+0WsjB3A3fEZXhtJ5ALu1m7CtU74DmcUEZf/lO+jJG2ZhJtwNmLua8CM+SwMPY
sTeyvXlaoorNOjJx3izEfsClE8088MQTexgpIjho6xEQYWXbFk+sMj37FbKUSMt+iOD49cb6rlTF
W9Koi4UbfAEi005mHPS0UtZB/uIVnJpm6/x3q5lEFIL+o6CCBOxta46ysYU4HZ2hTgGq/gRIUY+J
6Y1CCf1isMHNtLZX9zIeXfj13eRJc5fG589iPgDMYj1jqjpGUEsUSySMN+BXg1EtuDr0lLQXLXha
g1+qGw+JfxcPt/hPl50m20+f3qjE6QokmX+bQr7E52wOtspmTWADrc0j3Dj3OVu8bcIRM1rriMEZ
rpDAJUjfBLsaH6LDRnJmGDqE5nZX7wpWo8fjYsjkyu3c1AASZ/aHeBMmKMT6/QTEer+9PN8p6Yip
IvZhhzYg+W+rA3WLfxJBWKKMS5xEMRtu/+3FaqhhAyg83EPE3rk35IF0YeiUbjbpw6CG3mNIRGNC
4ACmhFskQvk4hNQtTNNPFHTWgOr/rolANCFeOWf0DCETG72/3OdrSQ595W/OCiNaZ9iKjBFFVhkQ
XW2/9fwJw3/ARUYvpnXvrA98tcLjBWvHVn+yNnOyWYFSNZ0jR9J0mvgAI6B42vye1i5uDxB1JVUj
oH1n012Fr+HMrp5S9AbJqbwK2csnsQy8BXTW+7yAHJA1gK3lI7EXa2spc/oVT+Eu8oA3LfbaVPGW
DVBWZeiMWMfM9CM9NfDLxD5KAZuBW5VB7njzuSfE4l5d5f5A4nb+jTpGZAftSWxFojsBbbR7e/y/
ss0tC0viA9N0ngPtfnAwoJXe1Q7uEejuObuKChk+JFLkPKdHjy47Azz1Jv2JUbeWh2HtcKD41Dsx
nDVdPxhaA/usL09MSAWF3nOVjw71bGu2QtVRHcrZjFqhTxmsgvUCkBRmWk+7j/g6eViXCQ+a6D8u
rS+CqHKZQFN3n04D5MQKulEOmWdtPNpC0gQ4tqM3yiG0+e5EPOXiltTdDGt6D22+yldoRiS/gYl/
JzSw6EJNx/lF+YBVq3b7PPUZJntyZ/RW9908zwmSNpIM1l7Nb5+eYq+I5VQQRyZf7IWUcD1CcXlY
9Z1kzNi/tHr/r9iPPz8069gtTLLMxsNXS7KINJ6728pVbmoifFLrOf+CifM4kzf7QnIJWjxD73qv
GC3S7u00miildushuyuqmCVtts8yKq3kttZg8lmLd6FYSv2Q7dPVJpb9BHcbfMMr3TmFJ+P3PWME
t18SZ7mHRe3N3OMtTZ9EMZgIbdR4bdKhuDDQgyw/yqm3QcEY6VdST+nmou/IVGHZAwEZzMwUqDHN
63xA1V6o1rpa1nzH177PQcqAQ+QmDU5odXejuEa1jZdiWoZNXja8EwWtg3zHXxAp+VgCAWPk6ar8
tshRmWwuJVC+FpdGCgoHIMgEDDttacellS16U1jOJg0STtustDs4e6tXEhq+Hce2rS+qTMa2yC0B
gqNKK11jZsic/29OYi1POHYiHWUelt1UMeCqSeUWYLd/NOfbSXfXlf/k6+8vcsjOHTeV+KLwVrQF
ZOyYO+VMnfAIIy3Sb2C92GTdY7JagsyOijvGNwsfidgq5F+9OyNO4Tv7aWkzZBz0t6iwYzarXibs
s0R7exk1J8KLlGxQu/BdUV2P2uUxOZBeJzb51qaFNpFozSrdN8wfss5oByY0EbkRjLmBhpFrbDIj
jiFL58ayPThbTJur1H49QyxVmnZXoktQ7NuYS23Evvk2KlXFqB8Ls92dFePrSQ+BhXLUVNs2j9RP
bnyBDJodMy9I2oUMk1SH+YNUp2y3MKSdcRjL1Y2Nzb9DdgmfjkhzHy5LowDquqCQAlTJlBWB75AB
ENMxnY8oaqAy+bgM376ITr8fvLjLk5BmnlP8o5QFP8rOpqnIkda7wCqJBnGd2WOUK7rD0AJWzGGj
bqUK7dTDwMiYJOmbkGaVgx25zG5IiuY6+zYDJrl95QyufLbYHgu5x6j928fzwY8JTwmg79RHqD1Z
KfFdYM0CItfojb+x6JM7TZ24sN6V5xp9x9qEc+12sxbtbY1+Uh0uIH/tvNuzIcyMOR2l1t8QyXx7
H+/6IuQkeU+dkRRk67TH+i9T6yr7n7Ooq0pbqP7fwKRG0fGSDTyRFY6DBOyJGHfZKyRszShkMIWe
cIbxLZ00198VT9b5zquCNE7WxZgLfbLNGyQlreuNTv5/YnZj6Bsy0TqE4/IgqTyKY8yHCBaTi9/F
ebHXoI0JsZnNikEg5wm4ti5t2nxBInyKpJ36xAhF9gpU0K8ibKsAcUKjxIth0FszcRe0Bc11zAUf
ZNU+bWpy4n8wtcWGasQXTlJ/1i7jJsb4zx3RwaBqII3cq6MijwWa4Jw0jCHDDB046aE4fv8C5l14
53TNPy4snwoNqwI9ze/GBuG5GD6CNWpCPzoeKxEN+GHQF7++MLRUQTC9fwaU8Iw4Q1V1Z8dGzZu1
nuIaYMXZdeImrSgL/zwfKnBQMZ2JakZG4XEkE8CcpIHrQ8ieMVCOTWVb6f/cRyWBilDZ+lSJXhNd
GRHwT7AWrR8LY8d8FeXD1+q8/RYI
`protect end_protected
