-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kly6+kxO+HwrhUf4NW9jMW+1jh65+LpE3SM6K6TafNpbLZjcFaxqwVE+0uodJiUZ2tuy3X3I4H/k
IJRaHkR9ruRpDnTY+32nhk5Bnce1BHV6MwiFCErnnSDBXde3TtdPOqa0ERChI4Lr/gVWwlkF5iKW
RSNVk7KhteRlhT1+eYWe4dTksDgvBNWzFKMB/alW3j4BqsxnPSJYrfA/U7scLEvnyBmkRLKy4gFL
gMW2TRYSr9ciVjFvosYGYwOCs+VmzpdTlv8tSp3iaoI88pLB+vxkkgq3N861+lKE+ZT5vC7D1A2J
Xe8HunBjhhAUhqNBDa0DaLp3aBfcOobG0ERs0A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9472)
`protect data_block
c1gm04GNXIhXLUjZT5b7wMZGAmnVE4axl4sL6U5nZcJwCloems5IL8TXGtu5/YossMj1B6LpuqlQ
uh5CvoBO79N+kRbwiIS78/Ep/ymvxToDi3Qdq0RYpJMXlQiODQ1MmlRKtqmcXoaqSxwr/guI47LH
fEq9tQMV2gjpFC6t1OtAWii8sgc4clMcv//l3+WVoroQNPvSEPICRJy07N4XmPNA9UNjXwiW3GXy
wzaKM4SKqRBTX+LJ9wb06yWj5t05pXImYNluMYSTm/491ze7M9eXeUmRiB+qZEMiiA1ZlpEagL1/
Ac9vXZpMduURlFOXGg4nOTsB41uPMPRRxIYulL/butaxw0rZmOhQBlqTkW/1TmYs4o/KzXCAOQDw
hXeUn0lY70FnmJCw0V0JDivsoyWQxaT7BOHaDVjWxGC6voc4u/0mPpZ8+Z98dyeVjMG82hIUdcri
FDJ9ltPLMRHcoUbsLzhoutzt6tLsVE39CSnJwiq9WpbmS3dHrj8Pn9yi5+fGk7hqonhNjAloeiXq
6haiMWV/HHPZfM7BZ6tiUe6SPZIz8vd77AUvaKei9DaW3qkuFCgWPQeL+i/yy+bzL2tTsga/wxcp
N57LVI2ZcTffmS7wxpcEab2hkbA63uhgpxhR69YV7VjX+bp+l3ywLJRgNgiSSSs7ONJ11mk4W6Pe
GjOUjb5Y431F8NyhN2hCddCAN2KfLhkdKXNFfXVRDHLPRLGd1zpWcm8q5p+/ekNw7X/x0Fqiak7f
a13dPlGm2L3jVcA/fxmXttYLUKwxnQyCWqIEtkLuX12khLErYL3UQ5m478cmAXlquxUksFRVPeav
JJvcVX/L+HFJ8G9oVdRcJWf00IzrfjIVCFwzovdRNdqjxJufSiX+rCsUsE8yYnHdd1Wsrbu45UcC
jnFS4+bECVZ3oGD7dTP28E7CDShBdiH5uC+mKf+ckIBvSYyiqkwEtZHfPjGfkqLRb1C7loR2dIYu
QWNFq+2ZkoqBftdTJjE1CcRcd4R+rjsuAaVpOXm8yNZW4ifcXnEyuGZUOktbxRAqMM/PX/R3OMxb
4fm52ARcDdi7igQXuRJ54PsxS+3gjCo/7FjX5ZGibPehuuIcqHSFcr/UIGwFjIOTP6bpPq/5183c
btp/mNjp5Z7p9B611lRiW+hGic4lBdSsqsC230o6LbJp2KKwKrXlNVhCvBGNPXBpJcnPXu21mCpp
Kwu0WyD0KFVssuUKRYbqg8babnlYaEejanccumtHxojxwRYPxUD3dgAJ1OecXXhNp5VUvXu5twpt
Ob5W7PMuNJKzCudaRYx/rPvrEcG+sru1iIMB5eJIx8JaVujH/gWAX8oo7Xk9kvYgl6SMJ09Qw9YU
rpQp/3uVfxAl7SPic9ZdAgOKuQV4FwMRKBrqVGEr70JCB51+7fqO1BjIhlV9Su0rvUK2YdmV6VWv
n51y3+KDOZ/mX+SIhn3cqy/PVrx4L0LQ6xWRHY5JfT0YKdCZlIskqzGQakJ+c2DbYVRBV8jLWqhY
pXZb4gP8exOQNDP3WCn9QndpZEqXmLhcx5+IkK+Bl1yzbywlwqLCaLyzuRlg2pzoYW+TZuRXFUrm
z83kdUpl8gInJzJfmApXE5YLldXaTj4tHCioFQ8iH9BRjir+B78uK1FAjt6H4PpLpsaojkNKJIVW
doHesQchKYUcZqlnqOXsxAHgX9Br+ruppGGLzYL+sNue1Iy6ZMn7iPDb8SpbX37YKncLCzKBdV+/
QgviwCtGYAazLC5Px+ACKnaWEEvdVfKvCI6qWes0e4AAJIfUtRQo/YLDFShPRj5ywzh6WN7sS510
7vwjpD4zgANjqSzPOSY3+Wz/QxhAlp4/4ldVz4L2ysgraRuYOJ5sWicJMHYBzs4KpQGeuchAg+zJ
BvXbrdvGiLt2tdvj314qx9HEJ50o0seESo8zFn9FJMwzcKGAtZwO3AnZJBj2pYiZcC8boeBsx+bk
5oqRKSd4tZIR6k4x1aF/XucZct33rRpD5OiIWAmTADt/pVPNrdkESSuKD+EFdx4Xx8SYbA2bB3CZ
51gAhMKJoD0BERB7exF52BIPoOqzcYM7lE6jooEcFEqeT7HkLqo0DghkJprWiCO3nTHhzesgfiHX
0pkIhEPLyXF4I6ZQBB11ZRc+1da0X16xqKDbH6mM2V8iGMExxGeSO73Y5wkiHqt1WTHth4G/ab+N
iwoT6dSt8pToGA5GheVzT+UyiMeSp5iRje3Yv96eSAczR0bmnWnk+wPYOwVk7LXJZi4RxcbZ6VNo
o6NjinW6lolV8luAAHMrvBqqSrm5lMrFxfPBTGQ1c2cuBv9ZYnu1VgoaXOlFQFeQVMc5xjzGhB/+
dIzvYEC9WDFr6EfHfmAmnT1hV8svDVvd5Plsfb6caLKerYkp0RX5+GZ82JhQcdPNhKKTQR2hhIBT
kAgJfFbQ3WzpBY/r1jIXR8bpG7ymYZQ66KgBy2EU/2UFgqeSoawnL728qcKPtfciMRwu30+3qWjs
pObQqRlz8XW1fED6paSDn3HT/HsUwbP06lOcObKCfPeO+U8rLgiQdY8ICskeGhXyvHi23OJmhLhP
8cgkd+TCJeWx6IJ0QtrijW6SBICds22QC3OjZld/QfIce+mSyltyVnoHMFrAdHhhCOr/ZqDKcKly
UWp2G5U/0zVJChrSmzYmCzop1p9rqufI47K+WLOuduYOBDY6HOW2scFuk8ne8XbowgDMqmQdDBUD
N/o7mTci24dKH07Nh4R2aQoI4DUcS0pO3bmUXiWAeWum7aBGz5d6PNvFyl1ja8FBKPNwTFvthv4X
YcmyDco1sl2aJL9DsFUfOpU2Oy4nludyHqGWXOoKOtT65N5itd4ais3gR+FJKkLg+KtDKJu8X1mF
BKNRUbCxeadvXmbSgr8pySBbo8h42UuTOLurky6oN7n3eJFtLcVsilfvqBeNcZBgkPYwV8csHTTz
79kIilT8RSgxk+S/rKZN6L1GJv8mX1ey/GCdJULGxpvYhoiCyF3s8gE/xka7t+KAs3qi7ibuFPPd
dHuZeYPx7xLFDCccZrevoHU4WUD4n8CmQ1nQw51pxHy2g17qE4jaCNBQWDI/jEzUJf6o43vEoRNK
lv+oKhMI1yX9PBRty6mwl3hVk1XRFoUC1FnYIbSB/0T4D3ORA3xixO+kvrjxC8hPA/Fan6Q13YSU
rVrq5iHHZugDcBXDioZ2OJQYiSH6Bj69xg45Xclu8Xhdzta2GVJ8faRLWpkLdnfdq7Lyo14EyFte
IBrtcetpnPkdQIosql31HUZ/jK1wJXfC5TdCs7W4ayzM6rdmEsXo8h3GBktOsaUdRT4Jns5tZyv/
LEnMseU8dP7I8q1sc1b8SgWJ4AhCgkcG7gnfVqLz2fEdiKVGX0jmbOouxkXb5BCMwqGBeeLTtA9n
sx1w7tldy7vrlByh/HPrxYTRaTED1GkITCpREtdynoFnDCTYuU6/RYSHb7GDTK5cZ62w/WpRtwLe
1PXMiNc6WsxCQ4XaoKgrVev0x/QzOe8GBbl/RmXwbSa/MRrBuVbcaFP/A6GQNcvZ5EGghSBbgr05
dkSbLcDHU/xKR1EQX+suJrGvjZrGp5WYrwzAzgmWhROsRz8nAlksUO3V/xNr3jhB+iGHMt7W10vI
8oZmz8TxZ4/3TKfSSaO8b0B0eO89zpXcBBJKc9cKThBRHHlPNX0rZQlSSbmn+YTuSI7yngsjJarh
NW+VKt5loTsaQO1YvcE5UgIRIo8Y5fLgtNunMy1tMb7UX3maKtY+eY3VKa1cYu3wcN/O3YMFjvMV
wY74yOVUYQOBTpqRQ0vzaurGa4cGrdb64QeXHRhqmA04tup61YVUoJjsmuA2K8qyK3vABWx9PCOJ
D5AmRrkHLvpYgfAfdC4w5xk+F7vNhc9ir43+fVbyGuIvHBt6Ah+5+5iEj8w7N+qHPuTa5gySq5Ii
byw2Fspr/nfd0dke2Eq16PYv6zEuNRHs5xndOtlyNaEXOrLzPcBFKmwZAwmH2MGWTj4yJTwqE15+
IrxPmr7ML+EAdDtgNPIx+PV/1O2EAPuBS8WXdiRPquS9D5DtlZ8HnqgcpwIqVXKNMALcXRBLgzQM
WOtR6+lojkHqN9Fr/PFPLtUaloqt8Zqz750YFX2nfz9av5D5aqwas/a8sm4Xxpx9sAYBY84eo5Uv
vrGbNFcmcD4VCmLydFsV6P95ROY7fW8yYDkS5q1V8dVKyl1v+gEGjrPiWDvHZaGVww7P4V8ZmaO4
r52GUL2NeKhFc6Ww3YwKGJa8z4TnO8WP1biW8U6aqkaUhPE89m671IzWZsOMoC51J9vlbwGdf47R
2mxaTKywUxuTu/OvnQi0IfAxcgwDXWADgV7zvlAsVFy221tNlD8xeORGIa8AdTt7i/5g3dCruNc2
QmbEmqLaRmtKUhREXIQYsdGTEKcRBeZEPs2KAVV5weEeMv5e1SyObm0ypoLCaHzEzSHgaJYhK4ls
+8i02S2PfnfzHnkMmrsRZ6NMnpOGw4JdGPY1EonNnApp42DWnQO5xKzoOzTz74LRRXHDDz0IIPp7
swmC9XRm7hrGVMpskBHWOsnjXZwraY/zLYa6x10zuXcUbFePiMNlMsN848yX6XHsKaSCFNPa10l+
GHBbgSCkBx76dMPd96iXuPg8U0shZghZmdLwiokWGhBO753cUQcnb/BA7i6NPtHtWwYSZYu37r/+
X/YxK6vUnwhOqxQ7ENhXvhYUk/xzlMUfZPGT3QbJ8ma5MGbmc1bhSbkyaTxsUEWUSmzS5Mmkwhd+
lWYFEqvv1SAh6eC295rLaAO97yEd8Ic9Gob/lNrIThQfuQSYWOoKCO12PBKuux75/xGIXLGb2fd7
32EdXjhPKHO8hKECAohSvX76BKPxl5y2Wwvb+pnN5YufwZGd0nVV7aHWRuJlj7Zb/Tp8a35yYD0H
Fe93mY/FxKaR6GseyscSZPiFZhYypnVaw15apHwI6VczQ9//PoO7vMVgzUCmT7SKvIfj2MI895uD
6+hARgz9rU10MQ0K0Fwr5nsAx+aPpN3YgVCCl6v9cWoZLWg/LLLhS9bHa+TCr0x9/MODmFhvCutB
hUAh4vSMZ+nK1bUCtNVdZHOZneyzwOL01YJ22WloTrEZt9+g+e+MYBnY9CaQBT+/TkqrS4Y1da45
s31mxOqoGEbhnbCpoaDMOUPqjIfh+eFRqy3eT8yA/xnLhlotfmUk1DxVF+CiVG2bwzYc7+En4AAf
JqxyHTkP8ud0i5t1mC7BLH7BLEmM7k/LsvliUmOZMs3VmpiOuXYomGbPyh5TViQ7m2yESX7EsJ0E
ZMqnmlvdOEdwIrTc/V7GNOMvUnLRx262X1QDEVBymicV1yMoIE35nm5GGaVSnQwJ/pi7eUoq9x27
tKH+iUzYNu+eGbQ9515fZ2MFPocVy8qn3AZdsWRYaCJgeSpknyFgisQCHiIMy2DJSh0F6EeWDZIC
t+UXnm9SaJrfLcM3n028/D4FeoBKinwA1oMoZpR4efEFXBKETaNfdW2uEbUDuelijPLFTgucFORz
Z8JcLf+MTY0ZpoPmF/VYLAc9UYqLXII2uQ+uRud6FjvDjzwvl/y+VFCWoTpyvybabbBrSv3KeQQz
HTV+ASfb9t7+e8YkOOE92W+jfskX60z5h2IxZADel5Ai7nNyuXUe8rnJCc+vY/0VSsRhyi9coK9j
2c5ZSaC6De3cSMtIqsQa4gfH0OKnGnm5iPkyWITsGF6WtPdU/EHeX3dX2t1xJGcFea5DKh6U3m0V
Z0og+RJ96qlKH7F4QKxBPrAFmFSoiuUT6w5DS2htd+0ZKzx3tT5cyJVef8YYucSzfTSiHr8BS8q4
VIdQzUjHphfTnYe5pB7C9xuh2iVzmEFikgFLCPdn15fTFJUJF8Ki6uvwBa0+h8MCScnmwTuhVvXs
1ev+WaGYJazD0RxD9pL61r/kYmp/t+9Xj4bKB1MViBzKJnXlLYAwwAu+IpU9ks9RsjS5q1X0QqfV
A2V1LAa+5+skApf9xiCBk/R8RgJzPjqd7NPk1w6qtDXnmmGg7iJftpqugXVHzAFGRd8Vq2Ryd0nX
K+sVh9mF1ikAGHNDK7n2Eo5XqO7OWkR1TRql7e3JSRi1U1U7z3WCR7HMS0qv7URyXofwKQTRSp2l
1KpmXvjg8c064DkhcU6hGcslq6glA6c8l6dhf8RQt90RO9+EFaKcifBYFZbMwp6fAcQ+rRoGCGuv
5SnNa6YXm/qxmkETxYEoEq4074oJdP706dRG0mru58Mtxu5tDUoXqMfw5pcHSxTmP3Px+p+6gVDO
xQwXH+pugyh8LB/KOiYP1Z647mqwbNjqOM987QJ2279Mdgb3dL7kyqTOs409kJXaOEtM+1Sg5rdq
7w697qXlk/i6uvMLzyuwKQeiA6nf/6JOqFJ5Vw9XRTxEJAe+hn/qB1moghobfuo6PRrAQdjqSKvF
3SBhuwQUfBT2nfuzpC4aSaqgdgtshuvXcmlvbGhmhL+meTC9SyfrodHCal8whgSrGsM5n847qYts
eUssDBhVJ5Q/q/Fncab96RqlVAO/+VZ3QO6YSIFvODb5JO7s6UzhELgXOlNvKIgvZPb4YGy01qMH
tVDeoYsEghR3f2fpn1DH0k5bd+GZBWjClu/p+L6LrEDSED2ELC2/9xsAmIVM6XkK4b0p9IWyBKZd
Qx66Xx6VIqWqlvOCTgLWkEiFHP0ZV0MybqvBn/NRVBsHb5zonyBBUbdd694DKLyB8UIBSxhtasqP
4lASI++kCTDAGNvvo0HIGZeYCB59nPfEU9K/KE2oFKcgw8y+HHN84qCldHuf3F0Qjyh5I+HwB125
fTgvjeYlaoiV2UwvrSQzNEFObTiDNMQXfKj3SfWy7qn5hkN8lA7Dyygwd+OTJ1t3wO1p3aZIltYN
+wzrnbva2VjivkND+tLP86wZcz753DtQCA2CjBXMw39FUVGm3GBZ5ROp6e86XtfJRAz5Eh4nYSA1
gTYabMBsTQubUbKweIwaqhavJ4L3qmMzZbWfuW4YsEyX46H6R6VpOn67DDyEnSjZanwcF1CAtx1H
vOab2HK4OmanPHo/5Jcm118i12+o4Rt68VvwwS2ltoc6nee6Rpj1ISQbNjrWAdJbR1Q1AT1aXqWs
EnL4via++wpp+87Q8SNLFoL9IdwhpswynV47LZp+YA0rGDLwDH64u/zDj5CL371A7bOm979UWrLe
8kcjgVoAO5fXcx9c8HOi57dV/kCXH/DkKudMEOKWo9T1+VbJZWZWKAHq5Q9SICOmBkrTUF91EZHj
U/PvvmFZPXe9YtFX+lQ70IPx4DPWDwE9jkgevCYdDl4lO8jIexA6r56kZ2vJ46SwHpE3QY6Hw4ws
eeEvl73NDozrCuGkksClp1h9GD01eHNuuRK1fsHh1XLIHRH5HCnImtGd9Mn3/+SSGUjT0RszgLzD
D4re1X6Fiq/Tf9SLuuxbD+uB1YWN7MseoUs8c3HMDBHPrjAct6k+V0Nx4eI7oqCqmRTNrRlEbrst
S3Eu1dRz5GTyfsFdiprKf8DP1KqQgHD9jGdFH2d/ulAILsG0qQJnvHGzmb2mER1XA/LBI7Kfgxbk
+hzuB87W+8bKeyT3uPhAQdfav8DUIl0GFzH5sCX/ieOSj22rDB2ZXOcrVqwE5ImxJlX9mqhKx74T
mpgd+BvxqdjouzJWMTR9Mfk+PrqHMMjeFBkItiCYjSIIAGgd51zo7ajkRCqFxBLZolFi939T7GEv
g9fVSdB8XsTdPnbIJbQSJ+AZbWteBqEA/Sw0mP3WC6AjyE11yd8IRsFpm75IntxNlRLOKnGbTbWy
hXfHTTK5m8ZqgoErNJkyx3C0i8z6sPed5uei+RtMojpeYgjm/OpoKoj4xaI7MdJsDyIUMHbyvpT5
Mywkk9pW5XjYXfjt/Xafh4M/biv3JYxqed4C4p/+xPTzsuMEOwidqByTccvZ64G82ODZ72dJaGYG
7X2SquSFE1/8e1wyrx/VEQFpEm0HZ8+aOyQm0UMblv+BDPG1gezou5shADpkuTH0+OypfUjR/hJ3
qaxR/zxowf455/BWltvq1lyXNZTqoCiCoI2/+sIsJBJCxgDMBSgkZJheA+e2TFrGEIf7ZlfnuAR+
lcXxnjEb412WWZF42biq6HLdcyp6DD8ZWV48OPVRxS/GJKnPVInhToYBEcBJ08R2c3mbM4T5VQnF
2HGAAFux9nX5aP+UdWGhvRPqas3twjwAWl8XpilNVgjL/EwJ9si1bNqpVBszc7RdWmalLh3bC8ev
qaXz+onF3QhmuseTE+V8p/hcX9sdAaFw7eAxbj654aA+zB7koxbfbiu74yNbmkjYcXkRVyDgDixI
5Nz4ujAMdw+F5M46bHg4GDqPh1KG96TN7zCLOcUinP7bJYnICn2gKSbOmgOjG+kwsJtg5Iy1KL6b
s/7EPfnjww2nyVM1uZGdQ4gw440wwYLAAiOUdHrY55KBqODlBby+apWo0RCxp70pcNT0PTOqCTVc
/LDnR1oeTJL10ta6LX+l21Tfv93Y3uWI4kJ2e6BaJQr3UxOy2WUczzI5vfuW9xbsquW+q89fKhbN
Iddq02mA4YZofrbE9p3EMi2tbaEMz0lUx9ABUm4XVxoUImOa4oTtKz7R2Z5yIvF6EbLOmx9MRrSp
Z+8A8ctUFv5cLu4Gqs5OhB5It3w5FU1B+Tkpu1epD+ToXI6K2ioMcoy2UIUHQB6sPW+8KmMVkNwR
HqOpDh8dk/kmwrU8x27J94t7JdwFuCXrzCJ88LhO3tatToqf89Tcl8REB7nQvf1778/Bk8KBeC7d
kexQ6ABO7zVAH6/wgoG/MeQTieIAAM3Wh2PN2A5Ck3rnzcp27yfFBxCmVwOvHGG79Y7+zGYEgD47
3vvLoIIkJ2GSO9d3LQzR8l3pdS7zfydS2p4MjOXyNi7jBef8O+BvdnFzTJr0jO8adochLaQRfiWg
C0zxLKPjM7XUirYS3+RzUnRzUneaHXNxXWiMOmB2VNGKXO+Bo6AyCkuyeTyz9CCjKCxj48BJpuoB
hK+kjKO7LccYSSLYPrXtNsxOEEugqgX0wEFuW3GAaglxZZmS8fHnq9ER6eMdcUccO9rlTmpBFtyy
JbUJ/Mz63k1fmVWjZJHx4ZHajDe+hu9PBnzPRf7CQNplV1GxMtRCblCEhEAYNB/ZS2UHVzMNIFA7
QLKlcDb245zGKfoM4S3VWGNjnatQPr4ucXBfh8Gr0q+ZjsE4xWsSVM8QIiK/0moCzwCKS6TQGCN2
WNK7NYpPZEBg8YyaSo2kRQyTShneurwWyDlc5RRjW5hkE8eXKrb/Rvi0pVCXrjDZIUfFkf3lro35
H0Mt+2kOz9ZZNOy2OdUIKmulBgDgAFgckulcq6ClZt7zzx/0vws3bLDOIad2LqYYajvcVQ0dy9g5
3kox9bvOTOtGZ4Fe50nPWEH6nwKyc0h6SdJlrMqgakKvAbvlzNUa2RdrwOfK31ysxkqsrDqtfldd
GDgQQ18A9P8Y54H/oTpJRw8nih4OU+P2JFZtWXZIbAdafeJy8miuwDZaAS5KLJUtGtNue+tHjOt3
RAOkDYGn0cVSiip8aQyZql3SH74HiqiDdCqZ/U8G4qxqYIl7+r2pCBc9cog6Ta7a82rA5fQTdt9+
SId8klNK3d+gO2kz1YM6ExwkvOA8vBV3TfSsdq107g5rhnJyZ+z7mv4eSd0DD0pUg75apUV5zeeq
v4HihHiklBSvZwS1pIXM7YcKSVK4ywGUNnv0NEn9v7bwpv3ak3/1k4fZUKjouYSbBTXmOpVtCag8
/v8tjspZB16DYXTpd9K6buj/K0m0htdVocax5npGy39d7+h7rWXsp/oGLKUhhWEovSGRsnXl7TmG
0maFWozoiaj9/AGM1rihzs7sEC9Drhu9USrc3WkmCjMfSgjMmerTN4fKrqmp5qQvN2mbCWa1dshk
QyVSzrv0YT7Rf29p8LeR0G0bKpW6S5sN2jybQEDdtvFuohxuf1Xi/cMvXR7QBkGdM87ac4c52MM1
wNkzdxU4085Y8SI0FNZK0ENKYHoNK2nDDK35NV7WA1lShLsR3tkFz9cfhAhDT1Awyh4M7MrUTY3m
swBWyF40ZnVNunus+xIhz7oZ4THzQJs7OiDthN7Z3+iE+RQuATI+lSICJhznXhFgVUSI8+hou/m1
0aYS6fH+Yq0Cljlrpq9Kz7S1RosSh3zsFasCDJhzrhK1qYZErLN4ISRXghgA1xYEQpFh+RD5jbV2
2YsMJBbSDoOriQO5gxNQySQfEIX0b4jcOzsEJj6/J6naEFREUBj0g9X8VsKekoq5Erj465SQxMhk
lfa4Ko1sLjdQ0NPbS7zCA3Gr0Emzi5ZVJSM8vA4GffTNYw81wg1gC2ZJUpOpCkX24T569+pPK1Vo
9gNSOUbCTh4n/Gv8RgnQ4iZ3pls8AV+xtEEDsFGliaJTFySACV/1xxIaB6VZ5tIHSNHp+0/6v9CM
EMvKOg0UBf3K0G1YqOuFqtmmnCuyPM86NIE8pxVxPFUdexemfu0AWW2qmOcTZENUct/2VNoiQhpT
iIyLkS/xoMtNsE+3kDD0/cG1439+60W8IDmnrBICklrV9Xabp+73TrdKFfPda9Y4I02+GyRqFlDf
an1QI0QENEGuXbQ+/R/L7HiXtzJNgWyI0xmMR2wMyr5VRSMI7Puj5hc3Ebh5VxlnOkX2l57Ev0xA
+9kIoSSqoK9AuDImpmHRGPcBSWDrblrr75XpB5yVhxAhaTey/7KF02KhyfWj2FoIXU7bm/vSQY4c
pt6sXPiSCaXCb8XOOkCfOtGSB8I3Qg6dgkWGrR2UEWNB5efRk1CJybF0GDasosG0bR3rnuESCAK6
XzDMSfEDyDJm8xvl7gdkrLL6Zhn8HpxL0MzGnUNoiba2iaLUxgWMhq3QIYE8pnXwV+PvXvmoIxH9
GJpZ5VDhlQ7FXbfqEe5atWuGoBW8zMV7N84oEPTS+w8WWC9RhcTiEpCBN6gDlDkc66gUm5gE6rgl
OjtJMBowr+LKiMNGrVOUbzlTJdidzWSX/HJxUK8aInygdRn4RYQbJCcZbarrEeXWAkDWYDLb7emM
iS0AvXKv/2yFYDBw6uoJXjks6+ff2lZI6L2KUVa3bSOaFchob7zklV0Ao6aMnYaS5E99T9jAkSL6
MXOyx1Put21/KvBQlATa6n5NYzf3U7Y7IpwveN0QTBImmrPhNL96Eu/IwUsBr1XG+gQIOA/6GtX3
hyISgcU6oC8xb3A8rIgWUNTZVrxjOb3+iynJvn9wZpFeTfFCMJ93R2YBvnBWW7H/7hWsO3qJBRhT
FMTCRJ7gEW7Ss2vrlG7vUQ6Lb2Vo7yDA4DnT/FiPts+ZdHo0QwdHL3A3ph5yZv9qll4+TzT1xHPL
ifcT0Kx4P1tkfmuPPDW9FvYhCVOtoMP8VBXRqldc99brZeNK0CuJTkt3HTG2rrThkg3QpEBU6JY/
qHQFkeR6q+DtJm9i1B63UgIyYLQ3UoIGRGY/CJr8pvNopd9KCJaTdN4DDg3/7dHted8vb2DotNV2
yalL8+ROVjzrQy8AwuwY+PL3H1RIbvMYmWxntv4KeUmnlBWFJAAUtSQqWj8dPWB8RBnrEj7xw+0o
YYQh/+ozHug3+xuvCOSEqlUAC0XYoW1K6pmV7l32Bp269KL2MTzY9mXBMdgJpgEC9+OuQvvI/k+o
wybVDjDeMueILiM8+sGuappTVzoaJ51JVPZeL5sW6fU7HbdG1iCSfH6bYDGtBE82V7I1ciOGO2MD
cU/y2mg1kOWN049jWubudpAlojgCLmd8VXQuIkLQ/qEPy/ydF90fmRCb4/0UNn/N6jfSTRRlEqyV
mVXHkpmhCHCsDBs9Or9HADAFgJyptLsGDeQfKHtbvtPFc36XnqHZcxqTEKDBQZtOoc/az9SdIZAX
ksHao4iNoktfeKwtxCps/CQDHj4rd1wnCBQ/e9EqKKm97zNeNbHwDEY3AUAaWqQvyudS+N0T4EgU
xPUyveMUiNoJT9lTanS7OJYsKH9KmzgoV556HHWEN/QrwlqPisCQN+sShvdxULfQIfVEtcMjjrWD
EV7q/wTRZKSxwzqZsv5Wlu1kpfr806g0VbdEY1bvlWe/Hwg6lrtT9WBEpEaVBbe0j0n9xsiTas+E
BKcTaC3HdIRc2AtRn3922km+vu4SncZ/H8fOaoUxpACMUAjQK8aEBR4FuY9pV+0ndFPFY95b37rb
yaebaydUekQ9aD/1hOUyEBh8YmZxJVJpzZMW6JUSHtuD8QmkkThtlssTvXQ7IVWotVi6y3TKJGLv
VN/f6m4BJffD24nBpqPpFlb9fvcHxJmq5k9ugjxetel3mrt850Hk0ApUxFaRbcvLFqJ7Bfl1HoSk
G3keLuDV/pUD74TTssyq+r+sCiRbSnJgwnrPLfGWTH2Hb47kBjYpTYQtbQSxD/UZGPnKP8LefFi4
7F9jEtwaj5xwQBB7iWCTjcFvNxcX+C/u5wYUZ/yHrdRmsqrvZkh2GuFZ/HVd0aIYnRe7DR8++SNy
zrkw5JNBHOt4X9DfB2GwdYhPWTLAMVxL099udIQmkuEWP2gJTqpHdniAXuo2nqlXx4EG8/VYfrb1
xY0phf4Dx3cPsA==
`protect end_protected
