-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hml8phQP9NY8P0RkQoF6PM6Alm1n0vnxfv7sAeccJSt4RIEzguBvOdbkYH4xBtdtKtn6QSoXVvhJ
WebiWNxyi8g03F8h+G/pjfRXpp+uBWBcBFVETU9GLeDGnYPGinMPAiYwdn1pqjVb85KVkUslyb6T
XklwKDNNep6OkUVmtjqyJclZ3PAtfMu2v/b9dKsvhwUrYdnYnFn5OKsGBacNuBl/xw+FcqQUqtEy
UqbwFDgW4PadWNlkRAYex5zC7/A96lvZ11ZEJdnXeH4xgU+sgzZH0D0DxEUaM6hzVDOfh1gS5B7E
LmY7es+7m+5Nn1TPbLbY6nnbJpdRNtl/5yLy+w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12848)
`protect data_block
PUg/oV8Hcsq6FtvvpvGceKw7hgChYSenaUohhbI4o0pxhasEEuoJ6ZXqwahexSkTy2VsSLqskPHy
cVtN+2kEHjO6k1ijuF4uX4Cd5umH3Q6+DjGDaukr7GPuJsi29qxwv5TjJSX60k/D/vXD+RGXDvsX
xII2KIPKHOv8CfPaZZGNDyfyWAh/aUyyCGkHWB7gRojgtOVYQP7iFgi5LPgNMCqZAgSmyt1OCocq
Ya6ap5c1hlw47jFW7eCJ91/G6PeVHAy/evsc1Ha+mUp10HJxXabAw2Sh+xEnBDkEcObxWx6xpPkd
PsMFBPVepuwOP/WKvPIX5QiqYSw89yQNdsp0WOY2C6R3MsH2Ckgpwn5CmSDg8s2fYiSLfZVCIVP7
BwI17eZBWVFlph3cAvawizFI81PiOc4PlhdmHaWKrIM6PT0V4uZ/t+B1S8Bajz3HW9PA5FjvS8SO
T0kiJmUPZAiAcfjpRbCw9WHevrurkB608IQotwPcng3tgEGUccZHtEeRs+owJIPEJQ8ADtHDMAnR
rrR2QRgDE+9vatOb4C534PA1svkbQauQl5bdLZjc2sI9Y1UWfuyi3sSFS3NzzhqeQoDqhDDCj3Yq
03dsrZf0uNCiFgCMgEq+xrY6uZn8WE7qRE19xqC63y1QFGEtnPemGvicHGIkb6/PNYv/WphKVQWZ
4qUEt9jw+ips1M3K8BER9OSmve3m55bZjx/F+wZsjxaYwsmbhQQHZ7vOPU5G5U/DzKwEPySZCuO/
Q07zhoSk1YcDF59MXnevYyp3VFsqhHYntenB9nZ4ZFsWMkhhhN6zQkjZhOxzWqMO8fRYnBvJ2om0
KqoUldRdtPTao90NVY+0smvQ0vmosBLDeHcWTmCuzeMGNtHJ2ObKdDCrCq+LrnfdCGfWDJ7QSUts
oikV2mz00FzPst6XrVOdH7Sym3FzDfjvWCVDksKc/U5vWLyqK+yBBz1bHJQDvcVIr3XFKkeX5TQo
RqaLBIxz8OUA0TTwddjXBY/4T92r336FPOGgyacFaK/30c/LLskK07aspsy02/1oF7fel0pY1cmm
eEiGgjB8UgRgOWd2vouxYo5CT1/+uU3nVn8TrOwVXLZ3ExK8ZewH8fuicek/SyvIlWTaL0Pkp5iH
zux2/YkE4/R3e3tYCUgtaHz2O49tQGts4CWHLgwiAQmFrs9flu6m6KmQUmvD2gFrhYM+5/v4ky5h
Yo4KN0pmsvc3+tOCqKdvmAtkRG6z5I8ptKmiGX7IS7Fv5og3CJ7rCjK4e47Alh75syD60sC5Owpq
r6UPBrLAy/Qv7muzw9e1Ui1CaRjxc5UuV4P+3kRgYLajrvkyi1flc8HGYT77Q4ld+KFbNRayKvJA
T9OqqGgzMkNJMYbJjDy2t9np05lEdInjQPIQ1ID7I3EM8LzTAe7jO/vORdQv5jipVoL/9NhDk1Uf
EztRtPNmpzhdc9DKobJN/tKmCSmhu7ENw7oqNLBGmp3fDWwLZ38UK6i0CXQI03V8ujEEqFw5DBLH
eF9qN262jMX1a/9yPSJLY7vM30kXmXlT00lEUsf+yaFeDw5JBQOBPqcpJKxU29jGTF/8m4dkKUOQ
ThxM5ZBXALVwe5VvcSL5Ssm1F+tDN1Q+x8DInZfxsZxurlnOaK4bqvdNQSBRWVCWSV1OjfQNuaBz
ElxjvjkCzzu+5TdtbeWhEiqttHOu57Zi/EeRWWcT0iVYqKTU95Jb0dPmgGiIjXWx4OckUXBpWc5w
Jv1P5n6fuVzlUvQEM5CdXgVcnSt1J/Wgk3nI7cELoFUjb4/bCABeYxx12dsB74u/jSWpN7CwsUuJ
Und++FpHto+U3d3jRI/9YYmKpHtaE8m0vPB+2uARxWBPzGekLUILS4jAkppiML3WCya49V4UQ7se
xiw50n8Er27zHZVZfU5Bt1P+ZWPPBkujolNhnvN64RhYGdohdV0HGVHlkkrTH3GfzBHn7Yq+dGQZ
94c3Ezm2dpLS47IMkDd0AHAjEWBPFXGK0IbwXT8rEWbPP2oMo6Ba8zYdM1bu5XzLjeBc4OQVznqG
7XGxb5SIYKCpMm/dGt1On01tezLg1MMFD6kIyXq7bd2kYq3ziqINSLh31Z5TdivA7w86R8UtNDOq
Cxm+LXctMfWgkrrxqYd0QOQvMZBCGH0gBEzmg4GHPwETfuCEs42LnVFUYzuU9Fn/8PYiOq2TLBDb
fN19WMMcMEcHmXDWinVIfxOzdx/h/KxWO/Vugwe+yI1KLkF9NcHLg3hAhkfefkgOThjA4K7ii1qu
kb+s79DfZTgDTErJW73yS48Y/Ow0U3Wkpb3wk3LXl1xMOpvhIFfJAn+VQHLUX1iczcfzExzx30KU
OvC1hBmoNu9+99/i8Y1+r1jm9rplIMVxJJaboU/WCAZ2pWKwQJr9W6ij8AByavJ3A6ynlWgLG4ku
SpPUsW7V5k6DnH3JaSgwcZZ0imSBW4TTtxQ9svqVaIxg/XBsovfJd84V7yV3G1v+CYT7piJb4ouL
zniUIurONUbrZbUGRWytratOPE1Ve8r77iX6S9RpEYo90Y2OV3rK2TMTt3BEaxq7p9/TC1Q8Qe9o
lUB8yJ1AhKw4pg0ipTQDBALUoNou6UeBh1DM/Mzl/ZdAnFsVApVHWXIcYAlKXcX0gwaXvxlqDXsG
Mc8P5OT00PVbiL1g74A8ToXMHCZbyg820SKA5FyQKwu3WBF8PffpkY8zLgcjBNtDtcFD6+2yJpUG
cAe7eD+PS8XLGqZPqRhZ9XBbt60dvJkizjnoI0iTB5ABOYJWUBjeAzvm3PTIP5vZnFsw0O0rrL0c
pcWoFhzcSPBJft1NWMSvUGvHP7bQRNPDJIdRfCfwfDmAZJYQ9jEHWa2aEv959ghOcnBWQYfyckZV
XOU/INZeDhyHt7jXg61uLU3msoX2UZG5jSFsD7JpH8vRR7ojEzPGu0st/+101ptF/yWFrp9d9Pa7
QpmRrG49dzIlZSWkDxeRSp7NvItNTwNJDIKz/e7g3BRvPB3tppqa/bQNfbwS5LP2oV3+Qh32Kwej
ojOm1nr9/JR5ppkLvAif2/r+MXp004tGmtapXGcWv18g8CWOnLH7tOeioI1aYAyeOn+246dMsaHP
NhAMvN3itcDTtweFCkJgAXgQUS+R2uYyo5GSrik6R7axdw9YUItwEtxrKh/N5jChvUc786nuFbEL
1OOVAoRBDJEq4dNrUwmQOd+YVdv60EFBoRwlvM+qTZYX6L9z13+e2J2Z8t1aDia981E0bhO80Tm0
OSckvkBOMLkofweVq9khGyXh/B4I+Pg9ncjHLWY0OTrDvw5Ohq0QLoSO/t52aqi3DiT4F1kwHPMu
ps4BAH1yfTau5p6iiSgGKV0YaZQ+l/SmEp2cDak9WOlMEJA4PtOEKa+5iG4qB0YThWBTfCM50S8O
l77wrIpFqsLwxggZ9RvBg7Mcq1biJfE8tXBF0hS+2gBB96JcLfLA6H0rfnYnBKZzI641Ye/YtUJ3
fMBAROlXPU9iBkxTK4UM27T9nHGHh7ujN+dVTKL2OT+Qy1ahYZtQT+baOnNUm6p0hnAXwEZizaTC
okW0tDA44QeohvjY0ZL4IPqwyUqrOH52wujsnCp8T3dYZ+cQVa1GT4p89S4g9xwpIzIyHvYcOqYx
JD4nDfIocbCDNZAp0yo6clbsuHkWxWX5XU4BvTnyzkXbkwzJuCbeRHBSndDLtys74OOpFSnm1DOh
g2dDpb5jwhtEt7nhO96a+Nbu31AZPWBc3eYo2fxdlESFgwmQo3ULg6BMmeURp62z+hVuP1XUPiRq
TVnoIKLqJdwVEeEXaTI5TrIzp6YJVsZI0Go79LJcdeHd9t2ZQM8n2suLsLTMKlz3jr/+PJy+pY3H
npP14kjBtkY+WK248MRtosdE+rFtvZ8dGRdn5KPoEmUTEu6oCZqn32Wt1J+W5xreDiCTygtHqo0B
0XlDf0XbaLcGxAVebWi9k6VOrf1ZQ30v9a5RoP6V3cqVnADkHR+d3YlDeQ6hZteU92/rAy8f9TO8
QJ8t5DiMNEki3h0ooHEG4HI2eR9OptjPZG20yX12Fa8uxwSpmXLLI/cezOb2O63A9cxadBiRf87k
8OwMaC4W095KHHoeQPR6j+YXqzX/aDnkmvPb30cUSYvDu5eqfiu+cU4JlDB3foxtZ/foIvgiq1tH
ztL9QvWLUTUEXZQzLSIy1tzjX3GKBJXJDLsLi8ZqQvZ3vSbZsjMWUwHN/Wg0pdKArbOKeWY4hwcr
/oTNgkLuR9j9YcSWUPISjOY/clT0BXQlcjSXBtjOclhg9o83tTGcDKMYhR9fovlIeFjrMqBvdZhD
uCA/L/hNm7QNgOIhSfoEGjj0FmtYWn/dac/8PAI8pU7pryPaE8IgJUm9jJprHIp1H/bkqYDDl8ra
HuTlsSA3Y3ACv5c24kBsTh+0xxBNCPBZVb1g9Ar+k/WIbIHXWSsblnBnnlDz47p0YdCQhOXamkBO
yzkYWACZnJrtZJ6Ds2bu1VBge5nMhHwATgwbysVc2r5TnGqfWg/xXZz6emT+DJSK+BeiWkS3/9ly
CJbSV9SuQ+Bahe6ReEI6LZCQ72A9umhKNnOfhwd4dn7DvXl4O3T5qNMRmBhB2IObSxhx97njmmgZ
Khj7yoIWEDO/kACb6JN7+B/QyCQ/etdum19ZOEOERAlcJUayghbKEusl11aMlLmUuSn5B53JeKRo
Dk9KnbVYem1pBuvJfgR7Qsj9sRufYkBMIM9UOmI281WtPzXc0VO3ZZYSOylQo9j8Vgfu9LDij13p
CKc1q+KFWY6qqHpNqR8v2KGcXWqEFdprLuguJGaB6oxPLbrSGgo3YxKPlk9O+5abYNLVGR8aO2G6
LtxQ0QwbwB/RGqq4sb2awv7t/SBw0zE98w3qhuPHWNt1SsOAKWM2SUFefbbUZo4Ht5gMDD2IySbA
X7DmW3O6TI7QRhSFTQTSE8IZmy6qjWPPVuZD83i0rK7/iyksiybfCpBBBJaO9Zrju+HmLPdyo+RR
mE1SuUFMB8MjZ9xAYCo5rgRYeTkaa8x8Jolp/1xMdDZG8IW/BsHyCQu34Ip+Zu9MW+BGxaDwBWXL
y3AA8QhZ76TQheAC7tkz1VPF7O8eANzNl9mMKfLWeXVnYoEJkehYRw1KLY0rEH7d0rYaxiAeYMil
zlBy77rY7pFbufGg52+AnzSe899NRe4OmhFdvK8u7eGSwWygb17FXzrPmpH6oEle5RNM+q7fe0yj
6JR3o4fhzeFbc6aAIN6ouFeIfn3+3f/Ht0sg5xqRd1oqri+6SHNUJe45dj5dE85nepI+RvfWjhC7
BXKTHijUJKz0M6h9A2Ev9fwuE+VgzcWcn5h1yP+IcNKqBxlRgacEqBYixK7mcG2MIrMZWKPmSG9Z
ZDL+weOit4NdNgLXKShWHf85hIfICyA77vnqtxzfo/QASW/R94n5OQe7CShkVPAW44EnO+kSNbxd
5ecM4kMZUe8za43ZoEa57TzbWcDOQZ+/tCQUSiB6dqcEjFAm4utdhQPv8LXPTnXuu5TvEs32b8ZB
MulfBTLfvNClbhKf1I1bLUYJJS/Ew0wnV0zT3N9EHiif91cY4mQfaSiEm0WNOlHIA0VztCVVFZ4Y
MBGVEw8ZwZqFFgezvdMctwR3q6oPuQwOv/zEmaBoO/QfxbPpEu0NBvWsneSVtatFf7VeEuhvbxEQ
txmcKu0p69BXXrey0E1EtgNJ+H5l9NLDzep3ZyYjGn7TunKwITeXMFfFsp/jo47vfTh1UfASo+NJ
FctDQdltLJs8aJeCWYej3A3EHtQ+JvXp2dJKOCQyqz8bgBWdWoxqFfYhOAB8PYo18q81pZcIDtgA
y0c3R8RZxHmn3rvyPrClOmVqjI1Lvz2qMl0sBfHR+9nAuNJao1VqB+GXf8yc92BkA3sbXvtNFKVR
Akp7Spqm1zT/jcBpahaKhmog5u0OJoyeilCzu9VrwnGIcqRQX80JQTg8wzzsue6DguIrDzCAleiG
B+2FIIe9Q+87RXNDhuUH3i5VpxnWakZyt7qRilOxXmdYjpigfSvoVDom3GDx0K+uQJQL8Au5Jqgw
cR4TtaHGh/gqJuM/fchKtiRCgDPQggLOW50CRL3Awkyt0rpaJusJo/T5UZSt4y3K055zbWNo1lzX
g1+/pKfvQV8RC5lv/VSP8umN0A357rPCKuIKj3pwBD1W+WEO30ZcJEF7AwbACHyezm2cSxnA0Nn5
IYkHYH9VoJ/IByhlKg3my2gxFStKtVz5W3LayyBsRUBeBpMpmRssHZUVx2xVHBv87GLgFVeft9G5
hRtkHfHwUy9snCtR3zqHKv0qVo7BTKO6Ryss48flmPKF2DCsgn/2Uh/Ndp0y+UdV4ILivT5e2lG4
ANHVbAFea72Fd38jweTxtuAr3F/PyioG/6mNxMV9CYun1wbBMzMSmdPcZIXT61/8CykYcgD0D7yt
UvE/2ftcemoxhmo0LMo5LGAewWk/MPJ6j4I8W4Ls0jty1WH5+xAy0lNyPSmVK/Y3/9pdMx+9dHbd
vAO3MDS8t40m/tpMpQZ9efS+ZlYqgVjlm7EmJ0/7wpibDLQ+JWtPi3mCcsv5BF7cZGdZ2xRdAuBx
G1mu9G41INdIMIlyhtPuucVPAH/n/bZtkrJnHYH2FRfqtR++s2HhZidVVS4qaCAExnRI9EHigB9x
tMV+IzxCes1EfmLXLeWIg6Yyjz3wpAhGJ4dhUw53yiftKpFpw3gKWuDS+3IFOoCKVj/I7u4OYT59
/UdOgJll5DxPruSPhdH8YDNgXJJtvdKQuvQZzKXPhAOOYU+82NI8MuFOGbfvMayhNuigv9RuPi01
4Rd6Gouucoqm0xcxDt0rT/n/ySktwa0W/Bfw7IlwqvCDdcEhOZTtmYbmDhEuDN1Ty7CXkXqmlnZL
IfONhhUOSTiHIGF/vsjBsea3Mrxa3+YzoJAe2WuPssxQRMqwzPGFVZN7CtGq07T4e1jN3GdzKuze
RJfpy856bo5aRva7NRSllIBsWwXBrqEeBpS3c6dLfcwiz3bHouhlLn9PuP2xFqHgFKqQqF4ooMkA
vw080UUGOZkJ5BGg7z1iK8cEUGmQzF1/nzz/XjAuoM6g5a10NYMiHHHi28j9cyL9thAkLyr+QSbk
GpCZjMOBkwD9hyDRZdkod+tsICjMMyvQFBXkTfWiRvWx+UdVq2dsg7Erlifs0VvvNOFBW6oUXIK7
1Fx780f9lzEmU7AljDH/pducxcTAr8LRzVX5GqJ+VbsoMYgdRJ+7d/kbDcTNUmzJvOzGlajkouIv
mNXjw/PKinTKTnjxiPnkc+W4B4kKGcDi+CARAR9XcCf11iD3DuYNMEzdxkq7YCFl47leqHKnlR1r
n4/t8j3TiNUdz67gWq9epryX9+lyHhXx5URM7MWDHKM37eRbccOXzs3qqFhCtr7+4UCJEZJlsyta
j5ik1mCGQ5dDo9JEsPgEYuy5o7pIWVT9PcmL0EiKkZciofIU7xEON/zgVnTMpxuPdyUCik28aCNi
wORrF8vz3y1xM4ZQJNwFG7itth7ZO7+nG09cGi3bh2utwnZlcGNC2pXoMRicagM9EaGiuzjuEONd
2VVINbmkr+DcKbw5r090KGrz9Z4oRZ2qeUIjMwTRyCE+ecjjhXUx1ly35BVx6hIWzGR9VE21ec8Q
nEuCsc6JWQx3jkWbtmSJ1toQ5m6A+dow/XwPjMzbk40cWMWO3D4MUgxdDVXu+HPAC/sf9bBpiAHB
MfbSuQzFA66p+G6zuN+nyirxL9gBLLkiRB31ES3gi4PGe6Xzlo8DQi3R5MLLw2pDthAZoEpd/JQ+
ZtmAO9f6d8YWJxecSNMnuh0lA3UaaOmxqdjDPMCU0w7ULpucP6vNTxav/E1gEUed0AtnqBAPFlai
2zMjMV85zazMWknLwrHzpMGoNoJWYG1G1qIcXd1N1e+oIK5Jk8F5EfO1ru132FxusqvNLf70RVIi
pali40lQL73ljbmZcLWdv6Zs4S29X8/mCiinyS3MgQu8eIkj7lltd+Eo9Cbcks48Fv8uDplz00Pm
Eem0VN1u6vKSXhQEqdg6Af8+M3JNrYXgmSabBz7ZDcCiEClgAjLY1KyKH0I4L5RUpy48mN0HFGWh
EyHFlz9p7FSZSqprzQvzei5kHw96AkDAJMO8DKOMg6DFqiCQaox0+r8fgA+X8ympHYd1n2XhhwFz
KaY8tr691QH9L/ha1/MHi/u58p+Shg0WxxEoIu+ogAOwo5QqGe+yzOCwm7Q/6SmwRHTMbTE1Lxwh
cMG/3MmIrCrVM3dosK8Ha+XODjYOGn8Cm7s0Banb5WJYIIWQ97kCACCJEs7syFWFvgHuVIQD6kVv
5D9RQtfoYljb7ZtGzBS578iw12XM4y1N30l+xLDsW6TYn6/nSQqc5WzPRF5fSNeL8a1QrDOBwFYv
fuXtMYMp1ZFApt8UcxiOIz51D6tLyLVMDuyK9+QdbYEN4QbM6CwD4gvzaTaYNsOwZ5gfu0iMxktd
FqglNgUrLfUiP4yz1c7xFKEnhiwL+SWKWJ2aWzRgHF5cGvyRjk9mBL3AcB6X26cnfhw9vp1BNGvT
124shfd0r/Ra3UrADtF3mUxfrx7W+b36iWbSxnEGpeGxyLBsh4DIXdbmbFDp5mCM/BqQlLiFmlYY
DdTlUrvYT9EizX7y3QjBFoIM47Aw910rO3j7cea4Lczseds2GZX3bgJroBzJsaYUtWiGc2bhNPLw
++KvmgAWBmSI18DVtKjykQ9dfsP1oE/tXtyV9z1BpYgSX7n5fWH2/vvoB1u1hBGxdrP2D9Aoy7dg
MYCzo16uy7madNfRW1WWt6JKBBKFU4HU0Kltt7fR747QgIfXqGVgrr+O2J48iFn4KqVNCimTO622
28xs2g97hyZIlsNW1Yg7RvfqzrtAOWRoaQI6mrln/tpKIlnrY6D/Q/zazJfAVdNdySvKI74+yGB+
j+P1XiBv6ssSbwgc2G0ekpZEGimKyucSVE6tRc4u2XoWZMCd7TOQHc5TEGXto7mfhqfa2FjiaQey
cNBUfa80g0zlL0QiJVccjbXGKZ+NdwqP8MEa/Wfnpoo97QVPguPBsYzwJot5MrDpuzEnPzG+55z5
GbTkeNKLXIoEQGrkg4jXBGsi/22EG8C3tLDAB0BNBR2x2an3EVjgbpuUaLGtJ2HX+ywUNYt1MM7Y
nbRW1kPriL4NOpQBcFBuhDTGpzlDeNQzty5Awutp8h0KwSgT6UKQ+xwtdpSo6Z8V969Vp8eK+cjs
QUDR8CvZ+FUlOfDJo1pljcy2f+gdGLF2wJ8vLpuSRDWYy7l19VvDTaZgnFgl/QmzUkX0FneECbd2
iHHEEeH1XTllDZ3KgHxW8jJQXAuiPHuQQKz+DWRf0BQVkEqQgD7Z2UiszWslhaZOFkwZSS2KjMbL
ijUWRKyNhsoU4IAfRKMtvBrZX81NETBW54vJnLb5UsLbs/9kZt2rJ8Nnku9fCke/ZCTO+ONCGvUX
H/3dG9+WffqolssqGo+CFMoBPZa8RkckT38KiaC8xH3ba5OUmOFxpecIwpGdKaMCjMGNyGf46W8+
9JgAH7aDb4x1tJE63nnxBdf8Vlk7A0qEyr9TLXRuYhZkxIReAoQdfY6AIJ4p7vOgePmOA4EHXtr8
ZcMuopIahXUn59w7CCAuAx3ao9NkKMEwqwBObfKC0lIUJwLZsZTytSmjOY2PTSmnkm6F2BT8vAuo
yVDuawg/aqoYTtAEFa2pH8mkIxkZwuMjlzdHK2mfeTHcU0jwjB6OpYzDnOyBsPrCae+sHT5V8Z6l
5jYgN9Ipf4oGGU8CNSjDtS6y5QzMJmSgOpdSisbvijmMs97l+Aoj3iKvqWbQDhc2PX7GywPhSIqe
YpOmTycNpDUrnky8cHOOXHD/TatDt1IhoHnXWFkrKirH6weZGMgLSTJoOZH1+MltBw6Avj79ur6J
7N9kZ4mAEOn8fKhrJPngYUTJyvV8KnYF35/Wjks+P31c5dlkKDT90RyOjl0W3BQxgmiH+vWJWbg/
MlHo5Qn6Pf7QhpDRjU8pVEHjPxp3wINGRWI95qBSBvCwzwo6uSNhvpKXKCCfblQVCc7WYirRVqGX
aUaA+NffyPgwAROe1SoVtg8Z7Ij+z8B4LgevKGgmUKg9iFm2dnCjGj7BwhnM4fTEhtRTJ9C27W30
hv8gDG5s60y8bm53F3q0jffaFcAvWXtjVTha9A3STDnmraY8/1FTTgBcvTH+/I2oS7OROjnqpIcK
OTdfDpxqusgu4ksuwrsTypq3r5H8QYOmxp5n6IWZu2aGOzDN9qUNIm1I4dPbF0Lp0d404doRHxNI
saBJA7ZFZ1h6lMGLJT+bZ895pqGnCIA7xEG2a83c0u6SBzp0P9+wUH5XNSAwlRd5vJPljZZQp00j
2xdZU0y6FmLTwgmXt/1/O98HBkqZmC4f0vVSQenLy4VZswfqwx/FJCWmzAL29UBfcNSZX5D2wpuX
ZLe9EFOxi47S7qFb43ahYtKaKyXWghw7UoWNchSfRncnR/GzR11sc0goguHzw7e8oLB1OkgDCNxb
h9b6M37gjd9ZA2EcRJHtQphKo4a3s9iCJMWczb1ieL5KDb28ScD9eS+BotjUxeSIIUau0XcP+ANs
yejd1v7OtDFEu6BM0nGG1oiVswDUUJQztHkau895Xj1jMbHtFeWyMW0FdIuMeyoB+L/0EoRgovQC
5st/P1x2VgwSwEXUIJiy8mFtsYYNz4pX2FCd9ZNdCFjZrERXXDZ9TESh7+chKP3FCzBcoLLF7FIa
ucPvcm95gh/BHUJZ/pFrj2rnuzIs7yHpjaIvfqnius746zqChIsjApG+MyPaglDr0ks48zSJKSCF
5n0efBgC8TK2HtNd2RQvmHno27FoTaaxQO4OZXitv6JjobMkOxF+h3KXyY2sKhBzNH57TC7ghPRO
KoMql0ZVcbncNKfslAyDM4PjLxK1VTe+byEbMZSkX6D3Xo3ciKGKKF+kh0/ph3a5Gg8tSRr9OtJk
+tMSXe2m+Kg2aQ2PCzurJdxDM3RHe7ZZBg3l60m/scTcaAQ+TZj/I++lcfXm0dILyl+0Gzsk8Zhk
EZtOr2aI/LeF0X+WWM0QUgupedae+BqI+ZDzfp01H0phknhRh58VHQMYbr7cdWOTsbcekVv9renK
kZFblxXFTrxJRKPXbN+V0O9Js3EVlB8V7KfieN5XjTPA9tudlcCSL+YdIuwbnr0ySGE8p3wzq/3S
fZZFkVUv4teprq1SHH8xDGAbJOGniyVLghACEnAz6pbtjFB52KBGW58NiL4jvGk7oEDfeUNLeqsk
eB/CPfjV3+vPocvfsV1pyuYpqZj6f2L3lGxBYwF6GrIXT/mnE18d9cE4lpL42VQtUEpFzhOZsVDN
Nh7gTOYXI8etWoLxwoqi98Ahto0PCW/8AXcBSZW77R5s3F4PXBlM0wi6uPzEb2QVKXibknHNa2a/
Er5pAWB7q9k3ZmWMU3ulggM2suodeBykxiIIBQqW698W7FzoPpBlktAtNO+Z9B2OtV8VutkaiCvM
U2Yyo2FiAwbYBKncna4AlE5TsVsvvc+22qHTrr4cvz+x+St/VFbPB2DZC8ZIR94TjlnNkPmdEoht
1hNKOt9NdRXpGDzL/fPNladsLeUrvi4CtIsXjZfuGmUnS7rCWV7Mv3AFlfrWuF3Lprhj1i9Ck7Mr
g0OpOxVTvXBYvbm7wlNkO6ClNFEquM6ue/StYuT5x/OyuKKcKP2nXlqX+2hlD4HSjYAPFfG0Pk/v
B3j8zONoQKzyl6VjxH72nza/CaBjVQZf37m2BXNBO72wCGwhXjCZ87O5XCldPVfIPkrJUUIgtz3V
1bjpPqIJOtvdyqsthyGJQLTrH4Hecp2Jei1oUtLsAwbKNCE0mBvxz/9JEGNR/twF6pXLmVLftqpZ
/4XXRmuvvEnabacKssRBXGW9myG7ehjYsF0VRtGHyA77q4tJMu0TqWC/N9aPUvfHkcyiv7VuwrCT
XoVxRW4vddM/9pwoWNdsq2kEFBPS1eXJw8jbsgXDGAkCB4VJaOCzy0+aBImeycOauByfIhWtabET
lafmyDL0lLNgmLrpTgVp16C8ZCFwHnCs2P+pLY9ITFQL/os69ctm1HtS9iwTMwbD8sngr9XHfsgW
gHwlQNwxHr3Tw+pEWu5eynkpY1fBmu4lr2TOgNrGAxugpVnkqJXUIIgoGJZ/cnBuXcc5NLs2a74Y
WkER0rGF+m2Djr5+WLr4KNYcIT2t1DXSeH6mdXL02+Fw6GPbZpynuethwtkbwqOK8ZbO7Yj1ocPO
LcT8Zf1QwqQrHh4pxBRzILiI8KN+puMqD9LA4IRqMxd7GYGmjrVxArW4URtP0E9IeFnzBBbBqbGf
j80TYkSy/+SLOw8nf9lGN2vO7OpL9kAT50+rYKBQyVv1who4SoNu9/9tKLD98PFtbYesXYe7XdOS
Q5g1XKtqeAQ+C53L5yUCXDbjRWlAH+JMeLZFZL4Nde+1MtluQ+sGzl8xuXrJQGbYi0fW9TRwvt/B
5EhSQOVwK8EbfitWYzShZHqWVXn6HvRJkbrkNaDjlbLNxvrLn3t6kqWKcp0NX7DI5eLPJNcnkfDd
XEfGAmLQCb7VbzgVIw6g1XS9DToO4DboNqKTgMZgZg5xLoRBUhygN9h2ETGfi3onIRDbiNuxLM6M
RpcudETlVoEOOTL9C0pzOXLfWk9c1QWKh+5LM7z2npVpID/ST1N980Yhiq4o1LSVlx4lbWtzT2sp
gVRq3Si7wIfmGXAC9HSXPZa9fhmFAaQNg/13766dzFmPkAvGu6I7S3l/ocT+MkCOihomZkd2oeTy
EA2+8vYCGWiXy9oLjKMQbqaoNNkfRx4nzx0i0XpHUzi1C4UOfAV8mpQFwj09QuJYTDS+EsoTSjL8
hE0yrfod4OzNrcvUNd8TOqF6XQTRa5vyBVjWZ/2m2jLDSwYMouJlXT89tksqvcMHq/Os1fwirdGY
OfrTWdEeXuyq8lUjDKpNwCgSncYAn6h4CNYiiDTx9in7l59nWnQIfvmnXorrTc2uwbwcrriNPmz8
1gIPjJ2tA3vo3jT8Z35Yp30bvZYiZkqXkkuvrFTjhfBT9+Htlkrd7CWPcb5Lym6tNHDOtwEmU+Ae
D5yh1GHPaiADmreJP/H78Nnd9jK+37tNVcWFdb0QolRgMl78Q3FUy+8u8FjL2XPNwlclpOEdRYHC
Z+4ZYApCiWU618TJ7XH3ZC4XUgta6ieYDGNZe6hLLUxJ50I/30G7NohtuXImAy/3O1MryDApCmQ4
PYWQ9emOnw5e1bKH0pTWETsQa/3Q3fiR8qhz/jq8IdIDAq0oANjLT0T2+2p1ejejmNAtA2Gv6UdY
ga0+nioP0k4k9Q7L87fmufOo7DuMdWsolYM56cua6qvPFN2DoaNub5dgMB0z8o1pWbhEEYvdUIiF
1EVj6XDQnJFKFNgx153lMW/4nV+gN4rl0N8+wfbOjZ5KJLRH8YsNlVztrbjsBWU3xB6Mj6I37zBk
PtWXUEXIxIJzL8+xB5NqNTUphMYkB3oLK8I4dv4CQg1RZX09iCGGWtJka6fIOGM/59nSOIouEYZ1
ITHQH/Tj+HBvE/xnhm1/TIcvw61N2qvDREGJlGOonTf8bwSWKQQU1WuueRFjUH/IZMfOPPr3FFic
VknSjSuvi/c63RoWEBC9wIGLYbv54J1Mzo9SBrm54Oo8GCSPF7R+jTWNOqmBCxKwc9ZOBaWDrg1S
ZMHvFeVNL0r9arvfuY69vQ/AK4ygpGKFophOJIFyi1l67sZfNhQfTIUDWaOAI+IsNn320EV3ZuSs
lOed6tJIO2SUelxpw0rhJZS9vkMEHSwOJhaw8BScN4/MRqwI4uEhDSP2aWRf4SFHFXC2NgFEuM51
DFjGuuzMu3pV++S4vGdhe1uwBzh0fSPiMJHKBXibEr1t1G8fEprdOs2sizgDMG7IUZXrgEwNtuNA
Gg1G34NOtANfo7lPsmOx3oqRqbgJ+SePRMCXUJ4900sheOOm+bV4vPJ+x+xOOcqD02a7SZrcKz3Q
g5y7flOC001RsDn4VPNqQZZx4SePHGafMzotmHDi217jTEaftzhc3s2sM/m1mu94A/F7mSP+tr1M
i5XSbJ/Ob15HbMep0tQVTStGyqFvErOUjnxlBIHLD2kzwMH3h09CmNE2fYsS4wQsRLRfrBSb/1/L
6JY9IDfglQVAkeCbd9usWlKj8rjokKbu9HncYtG2PLYL1LIootZXW0zJVlz+wTQe/shScaFpO/UR
qoPoKq7mwBfpQqR3D5hJ9ugsAaYX88twaOok8ocNMAtt69gVcBdEp1wkUcANjY+cPv5yG4Q1JUL2
b0CGX+nUlnkd9Xc2SmUYnINeUAKgoIKUrs1XYkp7ZSaq6TJ0mv7Oo/r6usE8Ye8XEYhL+LZJxoTH
wbIulLBy+76/zuWDknpFs+2RjuBNyZTyww8xDO239l7XVGlTrxCm7jy8mGlELC0S/7zF0lkvICrt
/hNuX574cFTZUhthXf5J+xZ8S+0ZToUGkbP8/6bRBqtaTGRJPJNkCQsXbSrX6qSbzJnLLXwlQ6m8
6Pt0OcCD20E6M0dwQezi9d9HzENY/1ZMCNHrT3+UALJ+2ZwWgxcm1pbLlssyQwJeckLk29aT2b+W
2N6yOgiZd/haIkjt11+AQTdwF/TPRBYKmLNj8W3ICK4Dok3f3ko8e5Bue4spy4ry5lugpYpSf7r5
2fjiF6DsOfiRzWw4QLj/89bdeeUrt09Z0rTZ1CuMXrEeH2L65oF7oKQB63ZGU4u+X5Ffk59bBXDl
V7pI5Y/E387SzWmABW5lDTlaQ8u2/yseac8tSICngDqx9ofRaSSHcrXVQEOfQ0LhWoE9Bdv2YdnO
SMfx9y5bCE5Oh3RBaMiIHTjUy6M3x9fQhkkWnXEP9h6e53odrZuVsL8EqclRK5CA29mIaziiVD9Q
PLRLpi+NVde6bx8bovkj70VzFukG5VQUY6TmIifgZ32KkmlXgcCHN0b369qDptIBx+gB1w/m/uJB
wQcx7KKDZ+URQdyBloygELaygJIXyK0+SubzdASwJwh9pVL24QckG7e9fPweYad2mmq2xsE+FCnL
leLAGjiW2T7++94zh+NYHaczk1nFPwwLeboAFB2vXWQ+FiXyxGsULJV9kBImB0Qhyclg5V7p1Y2H
7ujnvl82f3rmSlNnc7PGSO4hbAVKouwWiwgQCF7Z0VSO8TWLHpGYBTQzV8425SO/VXQJ6JNcrgvU
f7GRUw2m8/9sWwNhhc6nvEIKIyWe3vkYekcs3RCebRLJUkSw1i1hL3SS1zMo6Mkc5zid/LOzlLEl
wziwbfzBQN2R2zb7IbukPqKQ25pgn23ozmjmWRA5Na9DZfc4Oy5Lp9w9Va8aKdZoC6Q7dN06jS+X
ujnViRsLL3QKF1Ok90nuwXtb2mu4gIAqXb8e0NRdvpsHbmUBR9/BrDxjMLwVTklwoc/L3TxPoaFp
nV/1BhfIeH4jMAQhMrY34qF+2lOMqySD/utzCnZwMrDhREPsIbrEcDjfzTLNazYyfj7FJ5GXJRbp
TSjGnkt9Sk2IhqG1MifKF4UllN2M24ScSQ+62xsBG39g1tYSnvI6TJBcMmnJUI4NoqRNjlK/Pq7w
ALbTX6vaxCTIG+3EsY+xADlZG91AgbTEIDJeD1WCvrdlrTDWJBwY0+ILnwTno/21Ba+k8DIpWzAt
UYY9YC/7/mtZidKOosUElAFJhJlR+/A30zZIBox0dU7obF19HC5VNaxH+FGjCzfvU1WZMxVurPGo
ehInK+gNqw5m/+CmAEEJZYzRXKQAE0FQIQQnhf+dfDneHXs9OvlM3Fg4IKDYFAKgDAji9uXS6CNf
NYBly2VEjIXtY3fyR6p5EYnCuDbAX877BswfHfqgesT9nPV759EDsOmhUJwUpiBvbjXfOuOLyKM4
uQ8NiiMwx2SENZU9y+7inAWC+yD03B/gkgTtibYmS8aB7+wv9sQqoypcpv9cHlbAOBjeMJBe170p
P14FDkYY2r2skf6Rmr6YaKsluDITBnk/lGkmns3t+IT1yTpDBpvkZlkhtUqZZR6dKoPFRT0r1XeM
w6LB+g2Y4cFm9QYLm343DuQvx53auZwlRvSQ0Htf8hF7GyiCoEzJv1Op5mei44pp9gkhVToz+EiJ
Oft88NmPV0o0BbIXc5FZDs6mcC1lzv4d8q6xr6R2D5FVYGvv1aGKFjNvSjuCflUH7ZtTGxxRAFzy
yvrF3Ergkfm3tAhD4zqIh/HyqfpF5wb50GcNJrKN3ThK2BPTRow4Ex9pDwmRPzovUZlA7qjD31Cu
hHKMHeQwn3FHcs9faLiCbNKfpDiYUDtiEInwtx+KavXkX7yBYCaNO5xqbyKjpc+JTgbxjzY1kRP9
gXDCZ+ymhh4g7ywywinrt1T1LDDL4Z0B7XLT8ZlN7VEMzZyUibkNJuWy0kqD87kqdbakL+RGm4J4
is8hF3cbPrAbuYllQkpBBGeKPwxoKEieVw4D2Zld52qoPX6YhDwRbIZ/rZPfkRI5LrhnPG6z/u3v
QOeuaies3o7fsEQ/pdw1XnBhGYmPuFBGnbN5eUFbuAXcCmh2J2lSNuGGS2B1hPZcLpVOLs4AzS0d
yGjT9g6QtJQa01t5PANTWhQ0SbVT6rxmLDXsrRQhI8htvWwkfQ3zv2590bwoDV/xeqPUPLx2Dlmg
dNSZ1T8WSCaTib576E7KYIfsWcXgY/Sqtz4u2CSPl1bGokOtk8s3jwM3PXRHS/eDfzLsrsQd8VQ3
OE1934Hd/d1oWIVmHMnyFYFtFQGmham9PxlVStEV7XpqYjV5ZqyKY3GFHAmC8qgU47tOdhVD7nrV
ikHQXU3Sug7QFJXVj6FcSVr1ph8Ia5FpwSrFku/Ah7TaDyUGZpcyifEdSAeAzETMzTel1x/E+rqO
JyJZLALR3S3QUBbxOSWy0qZ3dE29s3U2ACcU8N+Hw4bcA/uAjf1vrgmonT+WnFTRTSPyNIpZeUbG
Trr0RlFJVQ6vHcnmyr8qD4++nkxpLK8K/DEhwbnR1wqgRphX4fpNIj6d9bjRhwCiRyo+F0GLAZuO
Dwln2y5Ky9dlDisv7MwPOt6TLsRQIwY=
`protect end_protected
