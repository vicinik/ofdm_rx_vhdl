-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HS8Hsn9vJmVzKR/RzApyezVJ4aR7ipjOim9F8/D4OjB+2Ny2M0hUmEs0ZOM7cG9YNLlmYIqok+UV
k0Q7JXY+UwDiu9NOrvwIwCcwwf9/jogA4iBgTBr4KR15Kk8MdhWCyNCU0oUPX7hWWyZv9V/TYbat
d6aCyY9tM1O6vLw+EEK55f/lOLIkZ4SISSqLYHczDY3UNfuDS5YlgEXyVeMz8F5scq6+oNihRRnH
2AO+SCmSPCpwIOi5RzXeT4U/p7/kLxm6dR6Yx3G+M74cj3giGS8xmGb/OF/Gf3qw3+v5GuqJdgh4
s0wpZi+sKVmJPAC16ZeinqQde7vDgk+8Lpujaw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7664)
`protect data_block
HW/0YMdj25Ym28qmv+0T6PekvlkVTIQ7v0aw7ZmlA/lfgnCfAEs4+7Au49wjDIJoNel7wzqnFyhc
Y5BsMa3lp/YMy4b68NWVH2zhC7LESe7RLFbaghOmU00jXs90ZBR30nibb0PTwZcguMRmX9uEqNFV
pdM4QHn6Bih6KYYtMRHcatZ9Lx+TOcDglYSbYbmF8izNo9JTyWUa0SdKoIjTwws8+qlx/kyInr0L
QyAMBfIhgL9eW7hwdkLbF0b/ysORTIOzKYueazbn2WiBYpzuxy6wMBnZfIXxq7m+SOmabgC/8ccP
FNr4lmeGGYxScI+xI2WuOD8m0TDoKH0V2TFYK7oHIDwhZjMDBcdRK7z9iHb8uEJi8IL8F4NNCTUM
9Rr6D+AVyocFEEzKufny2iDz+CF7TSZvypeCh0yL2Rlps2meKXl3QjK+q2DVKO5nSN+1iOu+mQ9J
8Cee+V069tlqwzKziN2HCW/GfvX/wz8F+08qJdvhYCF0MVIdDJIeikSmoDMzCYwi3hm773oHr2iD
LAihr/Bdl7PUAVqRP6Gq3oeyQt2gg/FqPRWqpTh76/4l9U7wnoTuMUXQ4YObJ3s4B1uOT3ko94Pr
QgzwWmnv3iuQwA8u01KrVQrDDn0ovdWkPuEtfC4lGaGTvbVFG9Wt97RuE8e/8mGEEzdI0nEWp2s9
L7FVR4HumzdBb/hU5yNDH8Qn0kOFfWzhJQ5/Az5HaZQ+bWOXMDJogan9cE6zp9aRfowbIg83eTdl
SuwbmVu/Qcb4DaMXpYHy0vE5kliVgatgGuTU/xXu2+LXytshu1o+fQba1f+UjHvPnVw7uMUkh1IW
bJF9ytxP9UMSP8CRD0LWHQEyvxzM5Oy1kbKzDNllkrBElaWcwmeFkvKPyRrknrp7gWJLd6eQ7nnG
uU1qdgfOVA6GdjX4m6NIZ2Gjc7G9vv/Wl0euLTs0ESo2UVVlfMq3rDbCWAECH1PYUUmQp3NH683C
0FQzutDMRQl8KMRgfswbbFBuMTF+UCYr+8AVyW9CeOg4LYSj1J2a/nSoeGMsJ6NT1WkM0LUM71Eg
Lco+lzQ9uaJvbMLKFvoI6HY3B7OgeJr8ZG6FOlKb0s2+j42wbPzb772OqNG2gQdLn+d/WeSkkQMw
2KeH3KN/rUA8UOXNqLodAzAClDgixTEeinfiaJTN1d3RcjLtnz37LUPr9ZYoa9ON57YKRpnpspGP
VuXm4gOv36jorxxJhIzQ/fWvtBPe+hqZEIjB/L44waOnhQfYMqFqusyoJqzKWVTFdG0Pjx1Zl3Jd
VEMATOrMnvp0Q+n245PIKDLjJQnL7GVK3T20pTwqJE3eUp9MIcC4jgf32K0yc6+aFfkk45Dl/qzk
PB+F4mTBrOcNSuqG3KhNoewUOeXrO3nVGaKicr8qvhbR02nAZ73ArMiXnUaJeWvI932lF9JA9TJo
0SNzzbB9BNFn2bmd7yFFFC39HoORLZrd5SaEIQkZkmgrqVKo5+qJk4mxZmwuVbbHaah3ix0n1fVb
lyyOz3LyxUeYkdohRhLGfwkkuGINwCRWpvTevJuwIaTY/n3OCpjCMpp2jTrADiEzjPLnsij5n5gE
zRZcNrTCfIzuO4Uhv/4keACGCkK5MUtuaqpTk9ms2mrBDUqwihVutliZluVtrhnf0b2/OgvPW/S1
anicZdVsSoj6nY1YJkC41VYKKHFwpLvuQphIOslIKJJPoeuj4PzRvL2Md2WTOx0WTkoj1MyDlgEX
eDNv588jrNZfmH5OLpBtlHkd3O7RLEb6KnwQ7kxPh4u7VHjiTXEWk4vspgheDf6IORNs6SrFTWsK
dcJwDjNqe4/AYpyuVRfCMpPP8oyzNEx5xa19Aic40aXhvowz8yDbqHMkJ6GSOdfM6Orp4LwbRL7V
v16hy87HrQn3UKxIbfFSHiGhsatfze+wI1b8MOwRcTnFjkrGrEAUBBzmJkc7vNh8V3t2wz/PsJ1c
xz7evnRv5eKDp6OV1Pk1+gA7mm5spLLq38XLYSH+6gftkNZJnG1EzT2XeajwRO49tpEy+i+f/QJd
9VDfa8/SmR3bx8v0vOlvFQw03FgTftfOradAEl5vaooop9BrYfZcCbrqNR81CrARRkWurixN2ny3
5buin2fAtnU5psZuVFyG3VVLFOUC2W/LFug8Jo/ihZ72SbITwBBlfhlRMBIDLunpuSPyGESSn2A5
PcedC98VATajHaOygzUnCESWKHJ5nlJYWsri1zm7jyhYHPcCpCpOUSRmabmMMzoekF6WiPAEPvbs
l3Py3qp7iroApAumHAiQe76bexrzKpa1ttRpNgvOFBT10KOuKuvqMdwo6y1bv6dxWAnTf+yuxr9y
CpAyslg+f59WtJV/GO/qKIoIR0nN2wGAQmTHKKZ/6vGfQuA7LDIxULHxZ/ytM9/pdlmzfjHx8ZW0
LloRceF+ZkU8fQdJ+aVeToXVzpyUqMUq7j9XfeBCwFj6f9I+N0mc+mAsXPKIiSRP0F/6Eu22uamm
rXSn3eXUFHB0q3qbLCmZW241NxMhS+H9aVUwYdruHTIvzOe+NdZFoLWaKvkW/vWNcpGi6p1gTAuI
i8qEgRbCxYJBskpITX9DwiyEc8xDb48fAhhTVkfQquY+iF+SYM28JaJhy2/W8/T8I69zf/mV8Y1c
g31cflV20Ggy6pbCHyTmWFKhPixB9+2uO/A8CHsA8DbrWfHBF2VpQdiJH1OHSbOG8TFySuGGPiou
U7aVGrMuPCJMtdestmdL3pFjNEh4/JIvkrbQAExLboLPaYvzSlmQTleRssNuWb3eFOl5Nosy3NLg
wu4rOTymFunD7AUOxDHR8oYGkTptcAVbrHTCQTwzJJXnvX5pFgbflrVdm9r/CoPBg+rOjsV8580g
YYGaj5GFKj/06SLj5q5/pvRAljBbfFsQCyc3/aOjhbvvbQabrJdozbBC82EXsYdvPlScryJrEAKS
s+mQHtB9B9KMYL7eLKW2hHkFKR6hgFU1wV+qR6JqE1eDmb8/E+iJ6tDY8YMTfNFHnzaT6U1Iwd5w
LlWfN2YArRntda/vYZ2QY6VyKQfaCjdDNbJY1kGKpxjHqouAiJuygoP32dcMspSQpOi5yU++PeVS
flyZ7JrO9wvmilQnBJOZ3shFD0fl3gGC+U/Wrd+s5RHyFdulH9oVDiOnD2IwqtvKmrtN4dIjuvso
IjmD9Bu53vCXj9yv5A+hbhIoeewn2MVLy96JflFwrdLllVTC7x9lkY4pcf+C/V4knnUKY38zW1he
n5fG1F6Q//vHTHKrZzDJogKOADdVLhEdbIPuuOBnRQDiJxu7hRfLT1KMIHy1q3hyybsT2SS/lGZI
msl63b7ubnGuJwCvoSFgj0+4wXv6qn7a0jx75kaQL96eqZMc3Swj7h8cGmJe5UPMrfZu+kVatooA
gWedWYlrmZS7FwuFRTVmgmIRVOjVoZEuM/ez2TLaBlcxU41sxksO08RPcVEd9EfdNDTLfIFWJ1+7
HlwphOqwzvhW39dv628i3ikiTCptkt4A6QZKWQ7xUK0ILkP3CxXI9DpZA+Vpk7ZZmQreuTtUAddT
V4T8zb2E7BKnDyI701hCFbiOwbbj78yF6scWy/gUvvKEBypFJujq2YtrCA20cMpnXZ0tTcou2Qhg
EBY0KKNV+GtxTlbiu/Rc0AeK9k+jo0jZiwckLeBsOGOZzF/PZAbEX3ihbkKVU4ktKGdbwEPg6W0v
8ZDK8oWx3hJR4+AjAAjYChN+0EHvmBSbgNjryoplVjMa8/G+NBRAC2f+jBrGml4Bq2c8hqyTPByr
FdnKhT9pDeMz20x1gDBhPylPjrA0Cd6s9w+UOcA1/Bs3Jcw3xBVV/xzC9p/IlxrH6Mnwico0ASBw
JCk69sZCsDlniycyoTEVyJ7QGDkScqGVFZCxlgXapX9Sfuvh7d5kEdSBF1qv8FcpcQB/0D1cFKAu
1U2OIzbhs8p6wYypGe6LkyORblmklLUJyWfZs2weeo7C2vKxD+T5+OxlgxeaZW/sz9i+ojfdQzBS
n434w3o1vguq2xAjqLV0pkpgPz1pGM3ZkapSOzVHiaHbeXIm7sJl4CRaxeH6SmDq6b+9Nkkyj2kw
Ek/flRlrgLg6tjGMqstCBy9mSCgZxxw7cwcnXGat222py2FovDc2q9KnolHQq0WfOC3Ril2rrUzR
GwXTFhfFZWMmTVLiRrtndiszsBniRgyohaFK+/vIatI2kcJpun48qfgHc3KSXY4CcNAXAS+QF/GK
P9Eb0tz2GBnbpr0fqrwj/9+zCPKsuamASGwA1F2ouoE6XL29HCT/O2bBD6HMulaupqmnE2YigHF5
vBGb4WF3YdbgXsBFh5FnAb3LUj3ruheMlpeAnnuNun+l2Ew32BkZSWF1tsi9Um5cZ0rCV49tj8Wj
wD4RecTMdRLYO/zWvmF1IU5V4fvf8xZ6nmVSuF6Qd9D71fLSS1HoeIJGTplLQHz2pr8k2lqfeHQg
MjRZpF/Qh+4XtcGDoVZgiaMd4HFxDgueF+eiSb2Oq/wrrlOzA+429jsCP/3nUXVGqYf0L1m4Rg7V
3Fa5jdPtS19FYRg6me9bSPeLfgl2S0gSRwr1fQJgXH8siN3pytD1I/ydnf3q1OOBCLdVC1ByBoZd
1mccYOWQ1AkgOsHUYESnmjIgPxbyaXySWktDptOAN0HePguJAoDCYhgCVpAhE515OBeplKz4rpDo
GFW+loZQMKjoOmd7DRIX/4NozFNFjg8OBrTFRwYi+n20kajt3q6IzwFNW0Up2ol+Lk/mN3GcxBA/
NjtdVF8V1cHJ0zkkvZxtne08InSeKN3GWBjPb123JRz8GB0go5uk87SN0d/FIKVj/8syeaoAlYjX
Lk2SHQrOorHSlGwNQ75exyV3Zy1fGxMpckUpRYUt8MkMT6EaqaT42ZZkP+QY8b19Iy3mtzVXy+MN
/WOH1EAEz9+Plyu6DoVW9jjve/FSeOP/G9mRuVU+kJMT4VujOObFBU7SASB7lvSoO3lzmbExAkdz
JbmIZDvyZkvWD39D1bdAZ3p1quQHOrnB9+AJFMK0WPHnxMeZV2iWtgbAH1JumSW0CIBrKBte7xxM
owFp8EicUS3+di/mSKu/u17U33dlHAfOqexb5605XcI0L10e2SLmWe5MTqe2UfAklJPSgYDncF2+
ZZsPwps/hqst5qoaT0YgOHycV48q35/yjeBGq32kUWSKlainvRtn3c6UPa/EeP+oZlNaqkZNnNH4
sCoutVltPgDyH2V1ViTOgiZwTMjRTLtKB37N7CW4ClxgBBsLZkJ6+W0KNnGa+tbJxglRibp+8qpN
u1ZYToz91vz/txYGex9pLiNDOgOtoje75/CvqKGqAO1SHhFtdQAFRVSce5jlwREEcsK4qpjhQQ6b
JUogeoxzuur+xfRvmCUBcZyqWpCd04Ae74+gwz1bBA/w/ibVi/YebzlOzMF2Z2A9TP3fFWnVR4W6
Qz4bD+upxcjy5TBXS0vHtinx0CvTJC+5nWoN/BJeY6KTFhaFn9FSL8ILz/ZlYhG9Cktt5VsmwtPy
H7sRIUMeK2KQvdpyW1jAW49vTqHMeZt02rTvIcLaLqMONd2R9X4zVZdZWt8EGmDCNQ+F82uGeLCt
aPcuY2UkWMs8Af4KIBiJWcbpWQ6ROalclrGRiTZQ7OZfO1lHmHZnryRJRFAo4Ba0RqRpvMSIIpMY
EOCUhEBHjw5vfjhMFlJ99IbDsgREIZFatMOzCLioEE44xkNlJZ3K8qmb6BLEW1JvTuuq9L2n9FyY
TR1OlvlrYco1/JkNHW5wCdTN5JZhHC1um7b4YcVqg1MMvs4nRQ0dMSLlOpq3o97ALvZZIAxVui3D
CEAR3DS+jaZnO5jochjSauxzfV4C4yRks/YAoVq+hBEczzMX7iIJ3pg1OkxGkHxAXkiBGk8KXvSA
VFDpx/Q5RF/ubEhct8NgU2u9l7AvzjLa6//FNBALEHY9RgIfwdGCYz92JH9s3xAKBGeyJu9YTgk2
CFnS5wGSlAr8gWlML2lsgzJFS9iyAIX5wkIXGIhUxCOEiVIdxekCmsh9Nk1PI7ffRLQAK0b8xZPL
930GuHQFRw1DkQK2izIMSBqpTP5H9jVG06SZZahS70BtrHZPboJgDHnFQ1o9K3WafDBPg5IQvFRG
99xvDeMgJ1r2u/uwQVUZoLnmINtKkiWJit2902bhPeNv8Bg4r/SAgzHbGAV4OguWdUPZXfd1Cjf5
9gJujvy8S4noGV7KCyL58eVjNmbtqWwSLT/uSyA4izA6X1dfY1ro2Nuii5XDj5fEJkUJD/2FbNjF
haCQbkn221rdkZyAXtwt9oKYL+yFnaH10mRb7itxq2QFJsnddX9nhXxBB8QnR+IeZxTBpxrD9pjG
mrsqC34creJw132/z0Jctps0WvHvS8zXCxnpteFaL1f+epauh6Zn2Gfo5v6uyHr9W7/BPhw3qSzm
I9rctZDVFxjTZwBbpG2v6MNu7LiFTVdnc8Yt2BSdJG7ITOg5IPfjQeb0z6Eo6EQdT9G6jHmXUqRb
WwApAIzbUgmTcUi8ehhvDd/fo5P1tgR7Z3yAdyK7E1GDfuoPoQUpgc+YwSNW4dw9/cVYEA9xsIAf
YcXCxj5qsOHypotB2xE3ltOf47GlaMDSUmLMj08II1LGlOre0dYuAbVsVIfvu3CFHfyvI7lEsha0
TCzlevFKq6lQ4PgVfQh90D1XBCyDwS0SI3XYycNY3fYr+zWq9csp3ewel/sfUZDfeNTp0szHRdic
J0QG31ORMPjzer55OjVAOxS0MreJLox5FhkvXhYJmmfJxzKgla5ruSPZgwnTU7UqwCwW6/so3F3U
9WyG+mTcnoKal8coMOkeMNOdrM0xDgn7Z+kLFtCvt3F7U3HrHRjWczz5ah27YBYysHC0ZREQ5Nsa
slQbcsX/pV8632Hrt/z1uIpsylScNGC/P1k8XZAZGlci2anYfqTZcVRezxxvwOQWz18BXrD/lVDz
b7+OjNJkLO+YcOCuQOO4d8epbVGJ4I/QR/WDFTaOStdNofiaLIGzbPPZS7fZq6neH5UQkAd54xBQ
EjzQTM1ycHkbMGMmVWe1DBpu2UfVCIhTAE92AlG4iRsDqPZh2M3kbE16TfzinuM+jHk+LbUQJMOQ
gVPt1kSmfmPoEIr/LqOEAgcx47CrVLbIlrV8kgF5cAHW8sGKqnD9LmASi7suY5iR59DnIh658R+T
qYpy8+K8XK0fCRnqMMoA9SLTL4SwZlhMmT+lyC8V8GeQoJ+2QvaLRsPPLQLBLZVxkwxn3L4JZu2O
sIZ+U5ax6c9pmr0snHaqDN1HXWTBoa8DI1TdPqtYqo57g/0J2B1aZxucL3LQXDh2sg8xIKoYJmL5
IvxuTNDlLi1cz2vPZdz75W2SyqIvymTLcdwhS86P6L9kfDnK8+CaDA1CNxppolPhBMtnCir3nkFk
guYypzKAvhvy5uTeZ7WMctjg1DooICrrYTGBjaanXaB4Q8a9paFPLy875kev4SSZ7LuWL0KpTuSz
aWEucbvOuq8UJGbrwkv0DI1QaqAIsChD516KLSc6CfHS7lt/hh5o7Yzi7feoSykjWjfxck2h4UVE
75NOTjVh90bZj+HFnVx/HxsEcHJx3Az+MG4TIa6ia68Zbe74/ZSqteI2EunAxbrZ4A6F01VpuTpR
QFI16y/TZ3mEc6pe8aZP7IiN4UInXYtVDUlmAG3Pd7XTAX8DPgEDnqB8xFHS04i+JfusPumTGSQg
0MCVLc83Q06FLiMHvhVKToDo2vOwdPG637eXISg7s9vbbgkcFl384yT+nKBbESkCWmrL1e1g+cEA
wltQyGNepBsbGNc4NB4aG/w9fMvVBWRd6SGM5+5t4gur6bjtTJGvC8p1FyDpvxvfsk9+Uu8XZ5Q7
uimeUEIFmAPS2Lude95BuuvfuV2BvwN0SBk3e8cgL4oxzjZ6VbFwSF90zscsIlBnmrHYpDo7IewF
2dUZXyem3rDah6x115zOUlkE/PHqUZiCemV4rt2qNzZXT/193/FbO75pW9jpDg1nZdPppkCVxUYy
2nbFxjS6S12h0vGwTpExQ9gnP1lCkflN50bbo4GlSbn1r9MIXeDmZ0wyOWgGC/HvYkdXNiB0SaGF
Y783JW10jI1eVfx0t5WtoMDWFo/wy10Az1cdrD7cSOhO8OXo0Lk0E35ONWcyXHAtLdjRHgCtf36M
oGIRbrDzy191d+cx0dv/qnmi3tnx1jEVWRur3s8bDSQS6trvXLovmTuvnzrFJH38v7/1VQ6nYryJ
bq6cMJwG7sYWmY1Gd2XGuL0GjzKEb1/PSic7GvvPCKwqTbNW+5b0KVR0bu430yZdS7JhpFrKsSQI
/x6FV1dSOZpJ6bPthjDk6MAobHWTHmzMg2spixaEJpf8VvoBO/l52QaZ2cCCXeOErnkspicYqcvm
KrW/+EaGkrtZJGdWqLjattlI+BvFFghL63HuiegJGY8TrivGvJTPYjTJGRC3UleIHIhjvExHJ3ho
duvAOTg+uK9u9pzGbd9aHONd/5EWiB3N/FTd/OPd6TheTVUnBz2PH8Yk4oeop5SFSeNR8rE6S57i
ikbdMPXOcmMd2ez+KmiE4623YTUlD5Lb8gU1GFBtqdeHLCbjmqjDRB+ET8IxNJjGAnn/BXXBdoyr
3JofgcfG52eFUTFPOERiBNcLP4cSnOsxVi/Jo//6I3h6s0w9a9dgoFWIHouPacXsnhXor4b8u9u0
pOVeg7PJe+Pjsqa/J0saS8df3LejKIYlTaWbnYRbhxuoqmgjT8UkT9t3mMB+Wf/4glNGuqJLkx04
X4Co/JllLUlvumSaYdeiKgni0WgYkCtLOx3XT0/bzQgPfL9NjpEsj3aNKxs9r1f8xc+z1GSVp3Qs
VRVmQOe7RcpjH08AFMElWNoxljQET6GQUY/3sNl/KbkLljzeQ0YfJxZ5HyVWSlUU0mD1fzDszdnC
hh6e9n3H5sFqqxDp1kXIVh6At3gRsFDAsdxXsWErzFyyvVkmBpGWZjwkeWFm7h28MokaciZgHrjS
vYvbQXmYYx/N9L7ShRIdMui3cHARCQDeYzhXOaLQ8444KmcrYsbIHuxKzyJbrjZjrispXprMvIgf
qJG8J/i8Gtv0vtVQ/mOXq23DuSq5fxs3mXI9UGNeSu80HL9PtULtouV0dmwmE/H0Uo9+J2GFOMUR
vCZlI7VGBUZO+bJqgvyRzBOTlpypyDehXgOv6Ygmg1CwhmnAR096JlnXjGRgUHNpjUq0Pk0LCadr
bQ9RAqLWgcW/CUZF9cfCJY59dJ4rGf95X+VV3/AdQP4zzeZvdw+MQGRdqcyYQvLNgwV9yINOX8Lw
jo953X1KjmnrxRybcegr38kLIKmXm3EndHGrJ1PgoEwodVRsLbi62jdQN5J8rWgBo/Bu4bO6Xziy
d6hbnE1OmexvXlbPNdI9kSC9SDu+wFMLNmJFGuX7ad175P5GJGg5rD8Udr1do8tWXPZ3qdu6/t/h
jMN8H9ynrVyflL+YDnRAwuOe/EGBJrLEMfenQFZVW3gp7FAeofJpG4+cx4z1h95v/C+KWTsPOoRo
ChBxk8ilRVTf1pIXH9Qa4+IKoFFottE6iMTmyKpCQE7aLMWZ851vTkHUaiPE25FI3+Y3pgNQlUXc
kDaGN5RYLbWzdC1oOL92Hfqz2uY3SnYOl6ZLoOJ2X1rtPghTI6R93O6WY9OzqnAXmIcEuziofoDX
NY/fBkTYIlu8OypVLgJfLeOKikYxUwMkwbCOzr2VXrXg9mXV1OnlbtEOMOPOJruBuVmwZs5cCGZD
QDE3y880we9lP8SAP63pU5pwKI6uQkBEpliWZVlJqMjG9DCR4qfnMS12anYgtcBaaP+4MuGT2mgt
FXPju5OOwoW4s9HARFbCV31ecRdg+fubQDDk1IYXSy8TKISXSiPZvR8PGMa8j0zFMO38Go3hXPXW
feT8bWZpC2IvC9Xhy5ncP2dYsQ46vJa3p2iu/n94oGENDN0N7BONeh0wOXGxVNlC6wrbNFPxIKcD
Si8vvVpxAiVb3F+gt0l/Qh/FMNOpXIxsTZJZVsoihtbltGFexsew2nHYX20+5w4WA9rufl20cGqK
z00ngWsvIxkrYX2r6V6/lBQyCegeX0R87JOwOHd7O8/Tk4zUBzQzTbyCauSmZVbvSr13mrl9JAKE
HZ3XgR/H+29F1cL/9SQmmwJSOsrdm2i1HaM=
`protect end_protected
