-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tckcblk5UEMZYAe+bc+BiQgDJES09GQDr5+UN9g3Fyb3vpyQhW20GEsGBbELelkmS6lylwye1iO/
zLnZgaX90etMSMy3fCSBgX7vLClz97ykV1I51xevEfwb3tBBPjHPJ9tFqapJoM/jOiouRxbEBT+s
l7PWrxCWLo1yfwu7xJiGuFeT0BZ/MSkQuiOGyItbpUIWU7g9DW2Myv9FgASudoexwVTWDmCwkRnq
rOintV5E/gFlnCujSe8/QGE7UcRIByXfYE54y8wJlSCV6iPUzNz2+b/kujJZtNv+Qesb8H9adDE8
uZAtUAOHECBrijwmQNhSllkzhw8WAitA/JrqXg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20544)
`protect data_block
Suu79YPnG9ESkQZN7lbHuGTseSgfme2D0j01QfWsBbiNL+BHpoGl1y190uKa+b7kiAxANS8VEqvI
X5oVrCWyfHY3GUQUADN5JQteK092itMDDd4vVJZBV4+kDW4voqjKovg/gtcSKMghdPUjBEICGalm
9pTiLg5IEn3ooFPrbfVuOqIn5Oyz7c5YXbF6HU+8GWUXqbPPsH6Ikxt0ADfIe5o83GofaFK1vej3
bA3qkakneoNSU0xnEQy/ajLOjEL4Ws1S6TJ3HHAwMJt9rn8ju6z27N3GC4ng/tgKsfScbCGk2W9h
MEFd1nQ1UtsVVtMHwrRsjhf9RT3gWsL4AEC5jERU+cELJUX62a6ruQx0FResxa0UbO16VxGlxYRE
3qIJYIgFYCzjvshVsqErt+XxUs7/92UQ/Ax8ua1w50cdIa2MBGF6MmYsbd6unaL6X/RNop+EZFMG
z66CJkh9IJ0kh5BSkZM6Pkve3TkzbBNaHrXeve9qbyPx/wI+XcliwqxEBpicDjtp+1B0gULDIpDA
rYaq4n0u6jT1r74N9uRcVP8BzKO/FM0RB3cHmuMK5/rJcE/Vz4Kw+58VGHuSGqnyv5cunsm0+5f4
VRGbSe0QHLwgmV/UxFl8MHtdUOP52o25z4asdd2aYTY2WqXx+aJhdYZTlaRTat4pmEfvuMoAnhuj
j4Oe7qOdAxxPVHeWIyGNBfIkfgVe/ZuoIfiyb3oNuRpa2JwpccEdy1jKwxoSddUq88r+3qMHv8o0
5MfcE/Vf3qydR24Vm08+yTEFbdbnjVm7UlbF9tCPIWYscdstWz2VT0iHL5uNAe8mHmKVYfuGLv7d
EONFTkY2AVqrbgXDfQGEL3Zhv+qSK5FCJUuVXqGUoTimAN3KhTxFLzsBxYOSG1a7tx3uBzb+KeW6
dO/1NGHe5/IFNKui4tiexg0mgtpJLrW5upNW7g2VOsHZluOxBAIi0TJ7h614hecxIA51HP1DdboA
SIS9t9iWHb0V+TW8fUkx+Ug4Uje9lybyOIwR4HnV1Kt7RWuVlMDnEbNnh1vmGChBcObz4CHC0ezc
Grkjaxy4OzYPXfIaA291vzo7NCNb4dBMeAbG3xewjjau0lsPBfSu200Uf43OpaTcmmJt+uevqSHG
t2pyoM+8gSrMNTrornVrF5oVsyA0yYJ3m+O1OmpSq73OEuGfkop5YmG0hCJJbg0eWSsuIu3cPRdM
am2SzcWlDI8GezDjHOzGHuXZPoET2bJa5JK79XRUXopRCkK9jWTaZDGjv/yU2OcMuvzops+U9NDw
Bg5DZspLS6AoXMF3FIR3pYN+/iWijfmg+3wGwT2D1tcTjHuzxhCbgsczDK+bWbGVROvHXs0mj6EV
4bBdiRHn++tXWqBl46QlsToMAPw6o+JeOEADsXhD7YZwgzVuPvmFcmy6TLkvo+zUvyescYQ/3G02
FMSN1TYDiOIAWZYTNji0edZvPsuPV7JkY5szTfgSbbB4Od1kvBVJsCLd+HNBfAYJBeenDnBEbOAB
kcCMFXbdjyAWRNFL+5Dqv82pwd8O9DYzPPHjJP7faO/TBnPSwCAqU/nS2PBSQLV4Tknep2j9FWkV
fP7H2sDz5EhBHRG3pInW9pYgbqdw0DLUiQswb37WJFeg5JTxXVBV7UgxZpj3VG9K4n3P/9hQpcZB
Halgft1JZhA+c5yO8IrokofTRixl+f88wogimVcFEC2Tgy16VNi2DTIwH21aphYAKKEfGSHFjwaZ
9CI+pBjAivFHQr3h2hr4wROLzoQNVr/CojFB6f/aVxqgL7Vtn3qZCbYXk7uV9p1tRX05MyXmI/VD
AFJDV1v2UPG+hlc5ZYsNGdB1pexOMpgGXQP4e7agkmGEAjLH7Yb4nDqSCl9jrydc2yqZ1zcx/Svd
714b63BNmnSk2OHdpzVmTYBeXnzezLr01N+Y5dbStKgUv7hcljfYC/7W64gXnC1DAIB2+o0ngHPm
fJRUCLvaDsmHELpEmigorcV1kcXW2xQwYoA5Z14L6thjngTJUs3KzE5d8z05QDhkQbXR7YEjjp9d
x0dMsAeGXdVVL1hNsi2yT8xdFAav+ISwJ2EAhlvmK6F8g886GBJGjgjWb3APSzhRava9M+7hv7Qg
kOunVlt/x52Qkfeugq7+NEYS6AIIFs2A9bSPXX1ja9oF+IselYWHDaF0fUIxpPUZW2nklH1qqYLh
lm6ufknfZLec1eSM1e1IpyT6NNr5dqzhWcUcDyZPBL3olW77rGqleW4xOl8FnTePPtWPBomz9F8I
CaS+J1646JlDATmWYwNDOHbAGyjHAqfKNe+wEbQNl+zx8Nm+vvhdkEzEd5tLjKoUx621OFzLlWAL
YmwNCe7FvWj5fwGCDi3pJi5WHfz3uVi81Y0op0xRlfaMFgM0+RnvHuv5o6i6PTv+eWS4rVqJNlNt
1A3Zf9nDql7xMIPLl7FO0aW7KjpP+nMjJDC9lD7rUe323EFRlbqKTF9PqBPm8JzVR6dpADgbR9wB
E+49unSGuQbu4eSyoIPNMxjoqFR/Tgb3zine73gdqtfrB23plFymt4SzyAMFpgvJvTprJHjDmhpu
nQjpnkGCxDifANF3cJGUQsiBLzZmxOkbGJdGfgF3YM7mV1+HQ73bZw81ka/uHTgwkNu/rfW8DHNi
31DCvXxp/OTCqdJALVtrqymCB/KjL7fx5r/CEe7G25zvEKH2xlVjHI5l/WEspeUXAY/61XrLqJHm
2QBUohomThvWnQ7KVi3axWx/iIy40leA9Aoj/Rgreq1BwPqurp2hwiAJvPX7cbh4I+7GYp7j/XFP
oJnvlj3E/kwv2j4YrkcXQN8r4PqQt/1gSYFP/dKwoHywpdplOzsMMEKns3A9rEkDgTA4jYmniXEw
/B4zH0WH+3SxPWKi6hmMGFd6PHXNZvh3JmiCy4C/og+PZMURBKEH8BoM0zxBrZkryhcXFQhOsoFM
0N9SI6G3n/iiDNfdkGGbc45ItGyQxVvUxwppRahMHPn+oqMV7OOYoNksnjsdYU0kiH1mPTScVwTE
dAU3thpK0wzo3Lq2uNL9O/Mt5BVBU435K3ZaLu/1a+IX1yR5XOiznVcxfy45D2jE/WCSCAeCI7u0
gouFn7KbcyNjgbueGFmq9doBdv0Oh7xjxLGUuD/S5k8Yw688UpGJCGCXi20l1B4q2KHtqR8Vl43e
+nSiJ+78z2k9GDh8dcOzs2b17qAQ1z0veH10wFEUl2Yd1SE0XhhSOvBbO82OPoxGzlP8tifcEgWF
fGeW67eTe0raMgKe5TW9YVCi1/71C7ccew1X0WIXD7aKK51ak6jhHWoeUCUTWl9blvDX3a9eTwx9
V/MMvURPkuqvLAk3ST3cOKmYCS05JRAYo3nVGItCzWsrd2iecpSijo3vo5mEoHTiB5zxXr9LExvk
B3Y0Wmzqhevywr5sPsCBBxxKRhmJrL5hIzdyuBqQWzAFH4f7fLgnyc8d/nknx1nKhqakyTpPqvdG
rKfw8V2dCytComluOfc52/5hqGv7IJooIBBKTui81hAsc86LEuk3jblDrBmPlX0za3qr90n9VRMv
ACvgQcU2gxSyqOLfPdgS7UvbSwTx5jbl3RVVADslA00CArhOfoyvbpqSoYyJOPNB82o9pbXu6i5O
AdJ8xP5KRRUf1wy81JfQF+3IxCusccHd+5ls+Iez38Y8tqpg61lwcDaNFMZ/6itXcznuUCMxKfo4
saTC/Xm5llC4i3syo9AOQw+wvdLvQPLfy2QgWlde16cdMcND/Xx6GrqEgb3ots128fym9wLNKEzQ
cvdG2gzhGnhjNCKJcb0nVUlAgEfEPAYqSB/ZqojnP4qbGnhvCdxtsZJnsrcC7JvGuF4+Pv6tF4EF
J/RnlZoeDA8qP7igfDYxr/5SRa+8jARg7KgFHAl8dIdeR2/km60qopfs+9sCaHG8NfPmFJSUVp6/
pwm6NeUj+EdrR8QZNApejFxCFOPzlFINcO3PfJe0yzabXv1CMIejiXNQEe7wXgfg4eqTlyKMKq5s
8kr160VS/JkeTLsFoJmjh651sl5DcZ2xyL8zyE0SjEEjRTSlb9PUzO8B7QyUCxP78gRACYzW6Zxy
aufLSSaphg0EHPPJClsW0NQD9eiI2Mx/ejcxMq/jl64Vwy/dgEvGN6u/0DJw4X0zowrKS7xxePWe
lA7OoTdBVH8fJzbN+aI2IjVoGBWZBvp7EjiByEBR7NxF2PxLRDy7J/4N/dEN1370GajM+Fh/QlKC
2vD/DVViU1S3kFrwTv0FPKgQQvDp4z2m6ecYUxz+ZMum6CtdohtBShr1OrFj2t1p2nF4BYrE1PHa
+RppTau/v0T0COPEQ+KzIIZDCQaeJDlWbrOIsniOFUUi3K2cJXVZOyVUumuXG8SicRky774Bu21U
vzKSl4FcqT6JX6Cf7iz9UEVMsWxZtSwoIO1qeRlFHRLcptDFzDNvOqmaBkWVC5N0KPFi8eRrVoc9
5rvC7KKC+J7M+5TqIxhZICbXg6gi6SPGBqqvhfCm/7RRWCuVMdwXltR4AwDoZSVWrDEAZdH6KCJx
wEvEUCdKzmO/4mnsimtcBAv9mU8zxW5wsXmRzvXg08t+J0g9PIJn+6dI7okRTRXqVjkCaGANqZo5
cn0P5qQ1idaxxu3QycbwdddGSp5HD8S8RT2PycTjNGIWqSWYW0oBpW1toh8L+XGzwi7ap/UAUFhK
15lmlY1QPiS7rBK2awuFy1dL6c455YV0yD7sv24UA1JEDhDqDaVauhM5ZJb5PGYvN5zvj18igQxg
ejqtdd/scOOe9SXlHIVHR5pmR6hz8zpG7O2RcWwhUbQyeCFxlRuCDV56exK586WGpuhNc/QmYZrW
7Qk6ZXAo9172gReKOlht1py+9VdUYHwrOCuC2ZHzUAxPslx0gXkHLOZVBnM8MtnBncRaRjf3WrfK
BeIzumNGMvu1fzcCvVEyFUCjhbfkmISRfuNY8t026NjVrI3D7hQPYi2EB05HzE0vF0r4ImS5POTs
81v+PXb69B2/SmT3OU2zzK6hDkY4dNTTILIFhdX8MY+sC+VCbVmZ7CR1vdiGMOSa6Rr8IKN41UGe
1+iF1o/Rs9XOslULuUHtTNFqVwIcLqL5I5Kkkeo5+eTOod7sxUsfmFvROIY4wOpV/2Vj+WJLRpBw
79B87PD57loeRv9NS6LNeuM9sZq/knMEnfaCxSMOLryrvWYLRhWRbRzTG/F/RBMvU6cUA2UUz2qI
mjKpDlM0ilfq1N2TYH3zdh+YuBx1oZFoM449pPI01VB3fi4u9NVLZHoMpl1AS9zWJvR+KturPSeB
vMxKSfyl8OudrJhGmCz975s/XcRi/DQoz1WmWNxkJnNgr21TD3QbxHx1xORYavqFus7r3kjHOk0Y
rhjZ5Okktn2zFPzRyWeZka2W5+qWquy/6E7hKHRjlHz0gY1TFbJvq/kS/1wONj+W85ibZYb8AjlL
jrIrr5/+64wSj26tTwkD5DBvMPL1+IdVSvOLuv8DrVOfA0SzuJfh5goDuf1ZbKau3sqz6egvEU9n
cKvDCBf92Cjkw8fRa3XNx9vnFgzoR5tdom4XqpWtcOV5oJ7ob8dbo1JLDwW6c+KAEt3jyJ1oHFU7
I16RpaMB0nq8BlIrhlCAj1Q1LWhoYnsxnuXi8mO+GpqRCYy893AztDJfXvyuzbZ5iWksyxXcnQ3H
GAUj5+0PUE97LoC9k8Xho1atCOYikdyh1dLqlVtljQdUwXRUIJoo6Y03Cdqd3QIssC8M4Z57iO1o
H/ls+/or8+t+dee5jEDvO3cktRtAJWoUAjC/Z2b9QkfrtIEDavAOupjaPxZ91GAq1DVNd3u0njKk
1xmQxrzVXl8/qJmTtT3xscx8qy0WH8esQqL2UGgea4skSWzf64op/aR4h+37p6mO1lz+eBGXnAQJ
rNfmGrLCJ0JLPbfYcwnq965fsdsQ6uAUej80Dv5NrP8lZxE0zn57Ktcf1BBma4GCQ6+jCxTn6bTc
3xPVwE7g+UMxjT39naKalWC+IH0RKog2PntCdiuhbbkfuk8VFVSIvMeWwCi/e0IgWlQr5jA0mD6+
i2LDUnHfKkA8XZehGAif28OSK+Io0yP/XfnQ5rUhrGlxI9ogm12NsT6oC3IPJ/u7+kgmh29hZBHQ
vxwehk5FDu+avVjuCf+UV+VMsc3EbRB0I3vkwNd/OXnxA/zLAdvStHpfsGbrfyOC6aTsH4NNRtyh
YQdJRSBU4LxvsyTTeFYmAloeoL8OK/vjQuMUPpQDEx1Q8XPgFC42sgSC0Gfub0oGfFoVEQguMmJ2
vdSdU2hNsaTtUZhWHFzHNWL7COuceqZfRqaaxY9UuyXUACp1xkd/3HSY8y2GC6Z7Th1i0kXhl839
UF8445dBEfnyB2E96yYY4X4YU/7Op5moya4PF8aXU/3jM/mEA4MV5dKbzpcO1qN5q80+vaVxv9ct
+sCMGlg+h01Rb+/WbIWmIhp5B06oCmEmd423n5Bynud7kKR/BUly4o3eGuqm76yaFBk8T2DEX5id
Nw2kvwrU/L3zgORMUAN/AN0GUKM8UAoGGnM3pMufbj1WV1cdpluRihBF9yD40WNQMtD1Hj+8VAcy
T64UTiQpdZ/TxoGXJP8Nlb27Bnfm+g54Eia2VBwICHxAEpVbHKuo6UEFLXzDf24qKcxD3Ni8VC3s
TILrXUNj+OYxXfFXI3fW5WQr6y4eQjWjAocwb+xbILX52+lb/dGLWwfTUSvRWfl9utPztQgoArMk
rr8h20qZLHWJYrbR6xkdMqXBASb1gDWeUB6ZAXwLAcmVFpZzx4lBiLQZOFUTIpCvBC134Ovkulj8
ACwunEbbhP0AJWaq3P8eYkIFcaHZyOBiGnMmxHyN2LDNcXW4nOKzXoMuilZNpo8+OQMZiCa9wqEL
7JBNYsaIxbSmrJElcNVV/hijn66C2CgfYYf4vtMzW2O3vbbHK+SieJwRcm4Nyr86jpHeraS8XiyT
xJ2tJq3HJHtzsRZmMkIJBDIkM5AqUHZw7HTngY9Dge+Lil4Uwh3d0/6rbpPOiQFD2dk+J4cKiEgj
6jUvoXnGP0Q1CptmnFpkVZyISRYwy6r0TXsYoMfiVxPYHk51sdrI1O49EFyfpGEJcpxLdT9z/CfA
NFy/UJuXbyOJdC8MfndlbFvFzAP3ZW3rWceqgMkJQ2aoOUUjS7Fr9x85K0NVKRrbD5+bNflBNBWu
KF9i43zkNBxHlyIXPPUDgtbiRdGncfSUR6ImPReopmKkaGyXZdKD+HOTpEIc6NRR5U09OvrBV2bY
va7/WUh1zOo2XOqlVycWluVZ7jm6Z8V8yppuk/ggrGriMlj+uiwS+O3fia4NRLsVMsxyKQjtlmSk
FD+Lw2sNBQORy9fyFJ37vFE4wA6P4JEG0kXekySq5ccjyBFh9sokeEURQzVOwD8FbyarRHK3sAR7
dtVhsc3JVql5x8dJ/3zz10OXjcktHJ4Dc4vTypIQv12XKAa2R8AxNzqy+3DJ8qUVOwfsyiF5SYM8
E4lbRRCGWKQGS41j88pwTCvFYa4NBcerKUOZWM+cjwc2l9NrDWWFQFa+DgHNg6OZsBdNmVkq7igA
j85drq5sk4deNLVI/cU0yNlNDpXSGXy1nhfaFlPBl3BG9BVnAKHpxf8iTCuEk9MZPQntk2tP76sl
1x99BZOs2ud15NqbcOj5tmeqPV91bB5SN8te42PB/5VcX933ARag/j6NgWZ31qtU4kY5G+xWA5xP
bZAckQsV7m8ZzJ4FiXL7EOEIUFrsQlGQtvbOf2nEvad2bnPvQEJmhyuXiIQFb1Trv5IOxqD7FyrT
9/lYxXx4yM8splJD51Z7fRcpAkN8QGk+IouajdSCgpjxbFT3mO/UuHZ7u93NCduNdvfez/qJ0dG8
IvfGTh/S27z7N4MQBJvPSVcwEOOmJze+tREkerVk9HmWePW/Xwo/QAkyUadrFhrT0abRfRfGMac2
9vu8xdR0HTx6WQsD6S/a6QW8Xk3xK33blpMLHYXJgSX7O4rzW3OnU9G3N0q2g5mludgi49PlSmr5
lWMk+V8WAA1NOiEiv/L4ZXtIROIFUfcmcz5BXJoZBPX48aYFThcPCPCQ3IudxhnHGuABMeMfFCJR
AQvrrwd2SawXrqzcHHI96tigT6VRXG8ud+FsKMC42Rus6A+gG0/1Tcr4B7E+2RDYUCoYviuezzKP
qgpEdCX8V3aIi8TfgokVQoXCuDutwWELHn/akfCMP1pWhGIMm/dHQGu3MBKwakMEv40iimnHyGga
H9nkVg0TIjMVcnwWtkMcKNUSgn0a0xigpR1DA3bAGt6vJdBSrNisy1SWQxgs7K5sRZCiUJWqi8RH
7kWrbIdaFldCD+5Um8w/BLj6PH7Y1KNzVlIXWJPQmw1gh129K8T8J4tN/7fys1nASQgg7IoDKUQK
w6Z72KjCPZgxJO79JbSBTKY/pIFLYGpAxJhcVwPxXuBYelgw/JkNFE4aQbH9PpDf9ruB5YqJD8+w
qZtbXmCeFoNXUJ8XqAXIWxx5Khq1kakmuGOSkwN7zVHMWXEhSKOw78vdMxl9Cbp3wMkC1oPeLpKO
RinZf6WPkCN/QFcBz2w96yEpZ/aN1nDxOKWHeFrKzrN3J1XT8gzTH4a6Yp4DiNmJdtLVwNvojpvL
m8LK9JuyhiZDAO6sIpjropum4iN+xhjCa4rGnhqWzP5mjml7ZCmEszwoAinmzYTPSTY87cO15Nz8
9bEinNA9oS9o4GQJxuDxub6n2vXdYTIJiYIMBXj/5nIVdWxqgYVxcJolawIvEtUgtv5WG/NLutCc
mGM9I6X09ADfyOrzzsiSCxQLChkiu80acumsM4KsgPFp2306+kfrvLhyXlS9sEYv3W9MiRz+uO9N
5vruaGvUA5d7Hdod8V91ojmJ3Iw0W0amOeGC7R5VnxUZrEQ2+avh/9HvcTirZIyTjDYuJq/ENKnI
YnjwbqlMr2ZxfoBSp+G779yLdxdn1j7L0KmGSzyVxUKVJL+0cyXm9H11vjosEbSGRRPFZ4snP5KL
ElBoxND4G9CjHTxLo2WzuXdPP1F8dkuf1qCgWMp7GV3ohiiotLwOVNO6J983fquHfbznNYlUz/1H
U0nN9NDYD2ztmUG+zgyCw5BrjEFgQuLtDZVHic2pY5nP72GJRb0FVZQxCadYCWusHYxEwzOo0Fws
mUARQwNrWivNPBEAqbo2J5QnE6DU1vFUyh+cfP6Fwdp2p6h953+V6V4kDxnm2myM3puYNNYqq+E6
BOaOcoS5ZCOelhtvtVw4Q3SGanyCOzPZ8Kx8dB1+Y6rj6iOTpy7fUxjJkevP6E2es9LvzRbl87Xf
6CpmOwMz++sQevkl5aTRtf+wMkjgpmTv20haIOlzlNt/TGmkQ0SXQpli1oZp3APRV4HiR6ufuceP
Z7uX1PNeQngk4tFkugmILzdasFEuZ1fvtXfaLRKfYu2H+HZcwymBCaOJq3Kfl53jos/IK5N5s2dm
+GNK0KoA/TLhNS7Y1BYmAeYipl8dAutpfZleiH2YTVtqYkxn2X4hXnoYHH4wZ8eXJiOL3xvOFeTc
LvSEg2jv9JCAJSjhg5RAPSezogVhGPYdV2mKTUfn/+ScvS7/3QB1oyxk73LeJ3Y01q5Lc/numRyL
senP5IUeZrh/rMqNy0NA7Zn7D8grUEoEZAxGYUtiiHDXTrNR97wyVnTvhfJ9/trSi+b3f3JoGOIf
VdwGKjCSCWG4u5SesfLsCMf4a2r252b33hzOJj8UyW5o8HiVFtxSQsm2mx97ko5gInchST3JP7RE
2GpQ9M5nOkSlI3dBLYdEU7C8IP+zMuzkKPGBJBthDC5EJezEVAtWn/qJTNDUzvlAixS9uTjEU3Ki
hdeyVvSdbFXtLO0Ro5AdEkh5XnST79EObbw35rq/tsCIExdav9SzsdlplWmylCh0Icp0OognoxF2
ry0zjpxbP/gNGrqHSmT3dkADN/x3gENBo9xQk3rwftoLNmEeEvE6cDX+O5HGd0UfpkJ7vg/mlF1k
E283h5h4cq2zX5ADg8S1V1+nUpD5gJbQErlEVp8Rx3cB9Ntrq+9A0J6980oV/eqYiYE2zlY/VvLN
xTRLnF9p/56ngDjSGsWraYniFmJiaYiboez6yX/ImEqamBnKBOcPQE48ubkADQSSxse6+CObUQK2
JSBGHKvNti1VRaHl31BcqxHhkBd8n55C6hPxKB6TpEMmOwctlH0pwVtJvd4RjpWRrYwTWx8LkOWG
p05hdszLiix9OYh4z0MfaNXAP1aO+Y8iK58FtqTVhjYEVwE0jNejH4+KxVlPwBVrPd7csKdcCLUS
FM2kdc/l+yyZZGgFbb5UqZB1oceeA+Lxv1J+IYtmo7o5HC0JDoW4mu9QjmOzDN+jD8zKUQBjeKR5
V3vTwLq5NtoEdqEnFf0UvuPOGYOVouK75n1hzCoEKg6fb7NJ4t1SnW5sI1cF3eJzfSlMj+LnlEv1
NHwj1gZRg2K6G7a0lrO+eh4S/PGMedCLNAfZf1pCWHtgxYlW99xmgIT4q8L4SkqciRKffAlZRF+e
kvv87VXw1pcLQEq3PHFJG1JoLbyeh5CjhfvHePu4u6Zswkha0Q98Ii0d4TaXX4Wq4/8daRtEH15R
aT92/1+Ew1z9SiuBrFU947Y68UZaBTyRBDT+xAe/0KwxVb7nsWp5uhYMZoNbTQQMUcRCplYn1Xnw
q6ZH43rwv47GOd6xHvUKpwloZhM34HG5+6DvENdYlD/iCLje0ndsgIw9DccPmQmG2ThLLWlYDLfM
3oeITYL1Y70xKk9EoR8tiTVxJao35ROj7nlR3RvwYAY6oVBoG82dGJqi5S3SEk2pBx7a5LHyRPqA
8KlwfIMvRh/FMOpovcQw912MQ3QdJprJ/fkX0L4OjFpHcK4BCZXfy62KG/C2U7aZIHCiJD02CWMp
tKM/vjzp4QfbGpbRh/qAaNID69T1k8adaXIYsM8dz16HoYSMfXOyOwSAtJ2hxRCwPLynkn11yyyO
rske1VdPg64RZQkhlBX9+BSsQ7UL57BZXfZLphGN0wzu0Ro69s0ygHa3+CoJa0X6HfIo8Uqmnmau
3+tGTSBT8OXL3RYl2qoKH/Lp6MxNXDdza6ntikkrtEQIGdmqmO2/H2wAGTy2p9tCTJzFXweYxLAf
cvGE5zfGN85f6Z7S0WohEpg5uHgQEWXqZ/qCAz42Wi/YlQclBzx29iR26N7GcydoHq6/xouqJHXH
gJz35iP7oMSKjSezPlGGDeATDpN+JDM7Yw7LXUEN2jV8I9aW2SsU5SGYuKXnq214hYJjZQ+tpmw7
S9S2kTePDflT8SvffKFaA74gwOKGcGUaybRYkBYXwugQSZS6BFBvffb/O3yM/BX+VD2JFkewDkUD
G5bQZuxz0mPCNQk5h+kAyUQt/USM9OCfUBiuyG8y3RkQ9B0WJS3F9PADQd6/VL98C/5WL9U7ZHUy
Kx3wnY6Em7h543y3Sl2EtPUjNziOpZxs7y8+lqPB+EN6+Z4qMfpx2sOAKLSKbttyUeA0j0OYn3MP
6hgCssa6nBO7UN2M3OkPrx+dCj4CEvloPvRT32bEysFmo4zcbJbRenAcjk29rdIZlm0j0IY5R0FT
GEDmyq6N/XgjeF7LaRQjambMClifQot7ZJ9hrMUdDVhPuHXCmIZRZU9H2HfiRTZzpFvcaWVvWjzR
Vc9ZsrG8BSgC6N9knm6Ul8DrKY4IwWLLtirxD7TMq62KgRxaaTP2UE6gBf/NxtJucX5V/iuRfvAd
MwO7gpq1VvWRMrisL03Do2xzDM3x+UP1qXWAaU5CS2H5XmWP22fifDD3rYJDHmZJnudGWSaG/tf/
L+PQj0mUBzPBWITiQZENvdIyeEfSoI2BUYGybmojJ3T5pIK7ikevT8xgqiz6j/k6N9DTYcBvMHD6
K/zzyETdpaTbzbnTaMsUnCA5GsTb26xoluhXZdoNqPR3DvB76QO/p61t+GUHqeIz6/bo6WAX33Cd
5qcxcEgVHcRSINGkxD0Hbgy6ITsKVXCHpFlZCjkLBZfw+5rHDPTWCPn3qncD3YWpeZr985B0u2gq
aSv9RUmYc7idZubNqvlaFsNRRs8bswghL2Sbk2LM+J3LmF4Y4HzswHBIdY+7cpKpRByvAL1IrPSW
qbnHYRNP7Od5DUIXqhDAIQAkAs81jEzchF5aO3NnptcBx9LdXV08aNaJi/4KtJ35pGmNaIVXYJpc
+3M9xHcneWJDirQLXOYY7NwGIZJFg6IcP/q4f4IVTQm4HYt5iWdr7nfIawDxkmU84WWGFt7msr6B
hCH8zoIm4WF6Eu4j3al28HhjBcpRL53s0hSnqmTUpGH0V5Vkz6hDBmkiEBHRfwOqpUpmsotySrxx
DxUrkQJVmUprv8AfD49ZImEkKftZfnJHOWxGt1E9BYtmLtkHMUkSDP2utvjC3rgAKt+s5XJtmkDQ
czlbJpGEkmP1+WtlI5nJnOcTtwHPnn82K1YWfmxUSUriGvOx4PMMP1ALXSlyFrj7D6S0CK+ILkVj
ibSiAo5ONGO2ktVZRGzsHf/wnem+lqYOsmz/5iT7/2rrYHjLuh8xn2bLh6fl8+ztl3rvb2n1RYJp
kmnFCd+lu7RKbEdUoZufp9tMZfl6rZ8p8yitITNi/HE3WJrDMbuDD9q0qHOir62dVL+voA3MHt4N
UFoE9W8MO5IaaKXNTe04NbsIRWRb/NckaPE+xpVachMB/1qNNs8NdeEWKfyvR/mBWsI6mU1sn67P
vvbZu+AWV9JKch0q5OPKRFz7TFeTQygrQR1jjVqX/exBqc2t2cczxQxoysQK+Vd64hOKhgfMNZvv
3cTQqorLWXKcORhg04/U8j2Qpdmvuwx1ynscxE0TZBx9jjxzpxeCaoPQKXGDwoTEho+y3+zYaJov
jaVVrix1Iw/v+mZL2de38gyOVRrPYvTJpl7ZTvmcyssYHLlAQrrEgpnwKd2aiQ8+kQ5kO8PUyK5g
I2UtuSTDB/1qXm4m0IkjZWlatSxPaQ7maL/d49IrQn7FYzvaVfm/Y+2bi3nhPnw5S1OytGHMvcdJ
EzjyKD6mJN0Ceh5qzK2Fundrs6QjhirIEs6I69JTTq9qI2R/GmFlpCF1koNgGiku22mwzTkj5mO+
EmB3k1HXlKxCxVownwylpd8BzUYhjaEC77f/p6GGh0Vgkd2t/4kR1f/LJrePUJNWlX++0yq1/gPh
Rvq5zsnO9nt9D2aVSCJJ9YN5nxC347zojGCjcQEUrGAF8/g/AazFPbRuMgh0hBY6qDiXEmjg22QQ
pZ9B/BOyB5dnT/Va7JtH2Wf60KTRYrlaCxrb2VCnfzBeTyHoIUngzkBrR8hUwvkP0LIdRr2t+rbl
o3Fet2Xp5YfBBjLhlZA66tEQCK9jO52k5Mtl3alnM5B/3P9W8CuXfKnaaQTkqz7k3SQu7I3jwc1X
H2FE77PDjZq1zbQq4/oMhsJGI7lvLVCeUZgGeeBABUdr919XCsFNWA1rzsf+OxuNQNXNicnGX+V6
0eqtawLg2eSWib+sFslbyZls5RyEuvL51oH57D1xkmoDBTO51hTHBVHrXDvTNtnpjKeoQqxZTRGI
fDjYLdHUP5Gp7ePs/hm6sbG5L4CYtqTEXY//i5huV/jnSfFdOtPRdlJDv9XwzhxeIER1oLWI468d
JK97PlUSOAsvwNre5FOGeOFVqOtjdqeuDzUYwwEih4CMlQdTehk+OPiw7OiJDmSuUGvHgEENY9rW
1uxRIzjfmmfo7pJsRSFrXXxeylIWrCGvcOkk3TFhYBKMJ0V7EeiyQNIXZvm71QlI7difhDVyt7mK
TDQnMVDJf3153ylzkFwJb7aZG/C+lWm6Et0/0XGvgt7icu9+2uKelnAbgFZ/oaXexoqAkvT0fT41
Kbm7qBYGw7TAW7Frt2P85f8NxwtpvL9AfCgR5hj1pX/0VAZgQqvMZPBC/QtT8kCxeITiqOMGb7ZI
iQ8JG/SbG/I8867VjEObitEDPoQyFqiE+oQ21AlXEUEsxc65NC+uE84PaFFI5CmggUivYOcLZXjR
Pr+ldthSFyw7a6JV6BpufhkI0NfvUZKyI5clIRF4VX5d0cdWvHAOVQsxldpQTrLTcAhxLH9r3Qg5
XW8de+7MMb4qyMZ9W833JPY4G/F4Lvafq2p2HO2v/AUFL9zUfx4F1UTXKPJUw6j75Zx/G/MylPji
HWM84VsVQJSunw84xrS9FcdkrGFYH07H3BVnGotbWxmP01f4OGek6Jxa1GT9lgXNQJVEGwgVsz/r
yv3u4g8mYh+B8g+FTB1t4YhTQNKYZhxtfHRkJGsboaCpsxfXqO1nZdjHoORvJmg8HIFyaTQJH2vM
05H0YTfNl63DCwnRmagVA87av+QS3zlnfSZlRsckGeBB9Htcg+RyFNReSvM10Y50tqbe4T5+GY3R
ptcQIK1Y3RPe5FAhq5SqPAkV8jzFENVwWhil0Kv2EEgEsRUzzeXQJvVoxKgjHNcco8gBU2cWd1Yj
QGg2MacPw1b+Q7uvUWBU2YytBd9x8tWi+2AEu15IsXv1zfIHu0pgQxlHZwFRWQEYWQMiRnRQEyNb
vD0k/4sa+9BlvuRwe1xhzwjiaxFXoY1C8AAO5j0Dxsbj+RQpdI0B9pT5+Axfph9BVy51KzA6ixdE
YCN+MmpAWMpf7BRmgRCb74OFVSkL3lsCVbqRFTT2IcUUktIROPAnY9C1BNUtvB2C6Q/8xrGofuOt
ha2MDBKWpK1tvpaBQ9CdTeoaaTdQjZgz91+Pu3+9ISxB0Jc/BVoU6ydOUG1paEkg+WBsF4ChuSuA
c0BUnRJ4NQ7pseoyR2PRD7v5e/t3b7NtNv0mCRMPmiFMbhFT2EGq4ZhrSy1hSoCxVli5rRTKii3c
juQIdxksMevhPWK+ngava92COayUMaFpBHYwEb7lja9PLyxmDIetRiYXvFQarq0k8KkFld0bCVXh
xRnuR+X3Q9X+nUIt5kbrTb6N4P6HDYMS9SqIU2eph9lvUIzfFRO3/MxEtSL0sk6zF2/SGoZtalvF
y/Nsb2sS3PfQ2pORZ+8TBTW5HHhyMwLNnpgdF/HcZVOET7q08thE8SQG99HgRGKGDjobvpPfHImr
iFcvGwn2n24SKsoy4wNcYm+q/ABXqDL3OKeDd0GoTZCi7EwRP08UnCCF1hBiGtC1Z3AgWZA3oWAX
u4UOng38jMTLSpr9GQSi1vHpjl6PQee+pqzGiOjn82bCte2Q+M9l3TwccjSkmcPDglAx7TEDwUQm
Cm6lowQKeoApGeV84Zzj0KlfxvtYJj4aw8WIjdd0vQMDs/6iDiFFzaQe34Otbpw/a0EoirGWpkw2
rjxzwDVknPCQR6OgpradwW22sj80qEKXL6YwTRpaZH+PqEcgtOhHmoVFfbFzqxrC2xAF80ZPZ50b
s/7duwd4mY9086wboE9GQtfv++c+OQiHM5JT79sjAuESAM6PzV+vr6m/f/gBGgSh6oz/yAwfYpM/
Rv/mmLI/n5dPHpzeonCO2JJ2sUIhxAVQAP8Ypl3kCh6kKR37xTWaXpqoeCkf4EviopHVT5B8tlRt
TlCsWgHHLCeZdB3VT8GVPsiOkZQZM7BbAheaUptSvjD35y+o4/plOh4Ff6i8FkcUMiYmK1TBkeCX
DyTyG386ded+3sOYqJVSdpWjkM1jXE2b/ZgT/WpxI9vv/UReZDtJ0lpDJFO03z5DSbUrz5D2kM4z
xs6bhFc1/dOZDjT+YXxZNQ007vbPYgZ+K11zVldKJu9Fii5B5nbhN3MjtL0HCp2uCQGgDchhnsWZ
i7pZoTA8YYZorYMJa0N0/7Vx4nWOUF286E/Yd1CUYPDOpvM71fXRavkFpI10Db6P9asP4FtJcgp2
wxyhL5RkWR8EvIMaIW6g21jUNF4SuUubN8pV7cIqF3H3jnExLz5vArd35hUMCj0YrvT0OrOUbgUG
qGBQ8OV6eOUtSNVcLbJYXh5aYW0IJIOwE/VS5Yv1AAEDm2Fvo/v7xWCpc3YmV/Z9EOVo0z4kyrW5
AsvvGC16kcHAi3vimjUNX9lkDpcbmi3PEiBFylu+DY02AlfC7wQU8tqcD2EHTz53E81epUFXOC7s
Ziulm1/5goaLQ5IDJJAjhs91nq9Ai93evp+idjg67xABrq0aJ0gH6vPx3hEe6DyV7Gk0YQjtdFwC
j3IQCCwWPoE4uujRrKmlrIg3cCL0YV08e90AGD8OrEymqdXj67CE7wBqCtjbSBdghqM2gpfuiwG1
Dn7Sn3/Cho7v07Eae0GY0oVIGpiz2ZOnNg4XGPiwbva0y1dk/Ue7wlGz/b5Q8FtCatpiAE3Xv/YI
4/0Y8tp6rTKVCSGVqfp215Ix5fiKMzKex0U+hjnfUoTAAIgXhGTEPOl1zdBRFU7Jhv8IXtiDFXjL
tu3bro4Sfhbh5cs7BfNh0MxxRcx5GHBV8h+M8ZiOsUPPj4VwERHVWk2tt1Hg0FFIN2CFhIiG7pnt
DC2RBEMB3clwxfZQWvZqTjQAvc+tZlVwRkRip6Nnf2Zsu5ueC7BiBqxFMCja8r9LQ96x7wOMD8cE
GyeUCDoWzqMv2+uhVuJZJqQBjYZyQAqQeKr2CtyAI5Hyv04+3FVeJBHv+dqxov90t8FfEB9gX4zd
cenh4aGwDW64BZ714SAlPqXFDHe+8EnomWGIrPp9BKpRPlZ7GFUArFppbsQus2TyjefKgj5a43SW
SX1wzrPtVbYXe8b4mpPJlZMwvVJPqQUuPlB4LXqU3JgYHPhCqAEhOkQzxT0YLoUgqNL0s0t9VqCe
eqHu8b/EJnsICH3+zDKtdq8JQdAMvwMe4T4Ui0SiBLa+rTYavR5521+c64StN4T01u2ivU1baOmK
Nq4GRZpBCjzFyHiWLuJ6fEOl1tVxaRv/M/HLLcgw3FESu6qIm10GE8Xv/xBprBbfQ/SQVKoYUtdS
C8SqSWYVi0gc2GgADjuTTC9A4CFBwT+qSK7Q/AN08TRcecHWovOOIgNLptCb25IXc7NmpkKe+uU6
t/vUtllOGr1rT3eRGl2kEVBAv4kw7HP4+XQBg5Eu6wYNYoKFefJqCT3FN1Iqw/b2CI+0tTlFfyhS
xU1UjItS6PnsTmK6cTCLd891xvWR1a9GKavLDzfzJ0Vp+mTlVVQ7/BJSF1UOv23ZsCnQXv3u7JR8
awvU//rWqZyms5nsJ8E+vGO88BpUUsT0zvax3IqINBF84PZcmJPORGygNTy49NTz8A5odc5pLeja
WvgBUkHti1APr1WS/ZDZGNPh7k1nTtojkJFyqjiiw1/sSVxDRHEVWLNSRnHvZFJ87gKacqoK7STK
elafLIfvBIWRDj1SF5hsQAPXZgyPAnQ8AWQIbIOYgKZ+6hb3LqVrIYxszqakGqHVEH49NY3By0O5
wqWDTiKh4B1ZP2jQRgXx1OVO1yElAGc5F83vhndnJYcFh4zEuTfPSrOtpAMBB2sQ/ZXeTyJRvu8v
pSiSlmx7kV6NNNHpZbp3RVPT2DIcyJDgvzOQ5ZX5M/mZB5q8Fr+po7orMtky44GYk/BFlrEB6O85
4jBMx7RsZaEOxmRV/+LpMbrhP/zwM4wr8rq/E6cpkQ4mk+Oijynuc9TvUs+GQ0FjoOryP/jtgqa5
yt1KA/VhaQF8iAmxSgz2HBGVTJmoTIIA2ECoftF6vRNzTscHALU9ihzoiuIX5Hg1d+GwHjdDP2TD
ol3o/nrTgg9ijJAdiDQ3ze7KXQaxEwWR3NHcAteD3459Dfr+LKgCXzE6uiaOo8ylzAipzVOLwdw9
M68HKpDPQqpkROaM1O4f+xtzQqjQTvSOKZfuMejUXdBarIhczQprZDr0EDCo6ijZOqJ2k4aabDzu
DL1WuKWyF5P+z71a/elrdgA55OMsvrRV8yuLSzKbXOeJjIg/gOxnVHcmDOpL88I5cTGt+iPGx1rX
cIY0mnJrY1UnScNIVu6w/h0AWiaeQf2RvM2HDt2EZJvO6DNpGIqAeeUYetBoKzSiYB6Wn/HkUQho
7Am3pz3np0qZGcuIYtr5cqnvMcvd2OXG+EaKDiIbewCg17P9CLXIUtLhOszqwZp0vB2y204OQIsY
cuugGatDlPk5M+LfV39A/KJbcf3E9d9xm6vrWm3yOqsg3wSF4Pn1WXhp3Et+d/HYhib2oTiKhTpn
IhQjoM3ArxC6mrOsnP1mc5N5RToVxU/CFXayEcEiKiRgplNRWHMDgm/9oJVeL4I6wb+QV9ZfgJn6
MO0A3UldQx/jcJ8fHc3+/V6SjhygHc96ZsNbMkHTpy95BxhFeVFcmH+5+LoGWylA/40U+5eEpXEP
CxJWC45Eukwf5KXZ4LGVYYqbeAH3BnkyMAPhnDWLrJfGmE0a1txghLFzk7045nmwoRoyIelNoZQD
iQi2nfnokH37dw0/q3DVw1z82j8sney0iytrR76mNu2S8NVk7jKSA0oRYRiZGwlOtAtBtUPl5GPL
b/ozVLIujnt4SfFGYqlWFsQw/uotFJqq1HGhRKh64zqeN1g2y5sY3gzCzmXifHi+lxV5fjaFh475
dnOXQH+AimSIjIymFh1xQ8S+otI/NkTHCppkHU/89omJpkl042O/aNLuPrMv4Jco7rkhppKGsgIJ
G67i3H6mUEleEc5vh17um0gjAvQMOoHg9lwKgrlzgBVlN2DOTyFyCrFLs+kq58/oE7BFISd51L2T
jXXpp3PpmUZPTHjKNoz+2OZxs/4Z0t0XqpsD0XaJNwwooP2RnU7ABnftHtYugU5VCT00FFm+Ft1o
sLo+vFRfq08BhYvRvg8rUHcReNFfB2JfszDMFNT9R88i8QHDa4sG/jdzp5m0o4jOiCKZKouElYjR
XodxGC4AVGbmNbzQFO2doJfkWsiGnBh66YsvoLMPlPOsEkzLD6tr74s7+z91trnQt2m0rJf8lI+w
GWJfkJLtuxI2vdY51FEtS3wnmb/bS1XEx5FSzsiz6OOus+7xVHJzyrQgclOzCnWbXkOyHlS85A/P
q5u3eWMVaA29pfT7OvUH15A2Xn6uyw/Orc4IAhAwMJK5r+kjHJEzaeiiu56pC6kO0ab23BtOZjDV
RLdDB3ytTQN8cZURIw3NKKNOe6PdezY+0WElZn7qawWv8BjDzAuBd8eWPHsUefWh14l+GBmhs65u
06ymE3rR7nhm7N3vZy1SNR6irXbabN2PK2OtwQsvNWNY9wYE/K0KbH4lbYFuypRDLUj+FnD037qp
NxGDfrlj3/35wulCpccVa2JwIwCcgSoUfSVTASCgv4CEnatkRQdOdcXWVKDFOyMGbg27oTXbA8ff
Wsnh4lxArXpZG01B5SpIyVVWP/xL1DSwiVv1R9dIgWTcn/TgNUDr3GHJQ1VCyKHqo+fP+x+1rpzB
CX4GfXGgSYpCLuWfaPZgDwF+2zhglAokV5DzUHfEjlr+CfmXhx+audPOwPTxTzRSfOIYTRu3LcUh
tgO+GEDxIQEkdFf7pHKuS/iJ8WAg7z7mS98mBPxEQIvUfjhaS6m/b3wmGvkrJ7QetgoaGR5cr/ph
34zKoDJzg2QqeZrC5dIjqg7AfiKnNRMP7gtBVROM1eOZgchQeBr9Pc9fML81e61uloQrO6TV+aqh
DOnfQ/6Ysn+zWGbj0hhi1803n1eIyPAUzRfnzgcPLdBhm34LE0tG3QScqmiP4n5iMVMheITPofP0
sI0TUUFvxLvWhI3iy1EaK6pQ0NcjqCrbgQTyRZEIuHEPJTpjcHNGA/t2V6HBQIwC47XqVMe9QQtA
ft9wrxTFhHB4WpIpwvJjHI6qakBA09U7oImWpFSv8oNXeEa3b6JcfOfMVvXXJNHEiUeMw7M1nY6f
qYBI+gPO31eULbWlxtqJUuGKH1JzGWWRBlz+wiLcOvZlsSl0hnyUE6vtCRovlnhqc5JcTrmOWNW2
Lg0tklYWnU9FhQr75D9/UO1wOKqDm21oScDllGrpz6fIw4Iakq/Ownpy84p/tXixKVpskXxRJws7
Fv69vL0yOuCu2tRdloM579n02c3oJYi4r/pV0z5/y6euduL8lWJIKLqxVS4RAakjj0SjB4nP1FI8
Dn6rP7KU8EytM25nVcw4XxylNAkNU0Htd/yWl1L7Pdf1Pf5t5xolM3emi/cN5DOThWNgQsxjcOMJ
07KlJKsywrUf5y+0zhNqULNEtstH91ESPiqyv7o9gNry2LT8T3lLnzI2BE4oU/M7lzkBOPEIx0d/
slMJDA8QXT2GB/gGJLpcmLcUfBsqu38+AUc/Nn31xxNR4uOiyrLTlvNiv4EiQGKLrKFaH75o5Pu/
hXyu0BH9LGvN7yiwQaeruuPSoPuZyqAGpK4LEf9LCOJinCaWRS/sJ4cdAY2gyZrBhbYu7gqQGN8u
1nOOxLUqMTjOtXqtRWb/BDjFC4fsK5muifhofIwILy318963TlDrcEXOeFvvD3qcueEva2eO/eeF
+kdpkN5eCGRD4BphrZtAKCeKn0KecyoPvzVoS7Uir7LTbKW2vs4fU4yMVo6uGdy2ZXPai6qJiXsv
3EnEgsDkftTa6sLgNEs9ji9lq10L1GmXAmuke8KMr+cWATFXGrRu9QNFgdvuHf4++H8lwjlOsula
b7CKNE7M//yY5dbLNiWEVPr9uj18yRBQfgNrBZ5dMsL4yHWbpLMYBzyQgJMuRT0uZ2h+99RN6WHB
d0TiupccvgyejA7n4H8QdseK89EyfRJewiN+38Uqd17aMxGj/oDvEln1WQrhpjlddmh3HCo/x3i1
S93e2QC5Pqsg79si1cnYSKKFjN0/lN2PY0m+nF/UFv7O0wWkz1Q0725uW4624K28I1BgvytajzQN
2Oya99XuN4N6pWLoWTirP+1tV2rTo22mTyCanw+SnvcJuo8ozcPUTuetBebL77NZECMeeJj/O5VV
CYiRkKLrqniREbHVkGN3eBU6ejEruquEqCYU0JNudZi0vmzMTfgDTB1IB1UZxVSZNQsaVpBTxgnr
J+WXxy2R4opdfloJTlLDcSAVWIAjNjAqdnqeaOxpxVpOci0c2U9Tb7AjhnIkOo0ZzuTHkmk+j5uz
WtlTtpa1uCMbnIhLPrzRTE4SbMvszEPVlwafFWXyAGNXqHHyHD24KojuxH032q9tcGN3nALwtgT7
tb8zk7Pm9q79yftzQEf/k3xakh496M3d09Yi5S36XlXWDYOsxCWkdQpfKXeris7Y+B2Aj1uiWjx/
V8GMfk2Pw1VIlhklz82vFouB+eKG39DsGdx97ze/dp5KPYEFwXg7v4LrjEY7m9IGbTBm16pl4/+P
FL0Ej7TTKy+cJiMYQplEjFj0b3gNPwXN2MDyze2XF1E2AqDsTt9xfvP2JRpO/ibQ7UEbDIkWlwih
lleRyQXCH0+RcpnckvS+xCOkR1iNSCN5c3MamBbtXiH+x7R6CzVQKELtQh8NpAPqoliNRp/hjAEc
BgFflQeUOCFPnhT8TA/c/GTSr0a/NbC6wTcqnGkMb4MKuV/nQa1A6xKb3gNxkyMie2wFhEpe4pH2
jMkJZzuy6DWN2BrUIxDa25Dgx2lsH2tEczLIC3l+iQlYdZ/Q+jc4jtw/+aYea9LLbI7CrqELv0Jc
YSMu/OREbeH3KoapSJ3zIaDdl6jl1HpXzPrnoRAMIgbLqG7ILJqw0Qd2OT9XXNNPI4k0fC4uWhac
lQBSi2z6WB1p8+8LslTmupn2W/I4Pz29t2VqEeIXjIj5HC9eObCxHGrzmTxpSlLRuNyPiYbCCTqY
L3Kauka3/3Qb9/z+Ts9x4M+Clt1bvkGvpGo2WJaN150h9q+ND4l7SHnZahSU4JtR4BS3a2qtETh9
LI3iIgCqLKO2Q4ez2biteL4sPoZTxB2qHy+EnCTJTVD1PH8YJMd0x+sv+hmZpn9uI08dlmVO+2rk
3XjyR8XS5RqzC/enI0IA3OnuDWPrR9Jkrf+D/Y8QM6/9zQdJsz3+FfVl+H4MD1tcR9bQ00WmoGEd
BxqaUVGo95D47LrxECKmjFMhAXQFuefN3JATPuXjDVAFcqnicgFe/8pxqK0tHZhvOSMD9LgQ03R5
CYGq7fjhUN79VVycx7apoaKFZERfvJxzqHNDHIseTkVbdvcP2ygseSM+jUTBf+rw6ma4HY2O+sL9
T9rpDdJm5JL2TO5Mncs0xAyGyLZn/hymytyb2miUvK3MSs0IvU072QsEeTq+YaCIWw7IT2cgfrMo
1a8foPxrLyk3+LY1i2f8A7hQTLJAuiCfy4BNK7A1N4ydrPDfpeFrXw3f/f7m8W3vfc+rrjskDUjY
3DF/DybQyB7ELRPHz50jWJTNjpqEB/1KEqqCYhpDB8enPDMQvR1xlSCCB4lz3MIxVvnc1ibrJJAJ
v77ufWBPg+Y9v5KvjlJvyJ8phwMiFxqJdKBr7nS16cC9m3NIGi4WdcIQxnfHGNoVKpl22KtqUtmP
nt3bUrV0tz2YsCN/OokPooa7zyz5NV0lKQC7TgvICggL+MiGWzqVz21BKg/z8t4GaswGa69ZzDzO
wCMHd20r88v9XcFrhDR8PI54dO181F8YT0VZjPxJ9+tFTeFXHrhlNkeiWTmh5NHzDUls76eKvXqq
CK4QiFzKVAKGXthh8Vo5L21z27DImguTmItghwwssTqIF9CTv/dhhvN/5dg6DbHImF57LUay1sHc
IOJ1HEPvUqBQAli+Rm8narb5kUi7x5RuCdKBv87IWchZXCSRlnZrNI5X2sHS0NXwYuiX7R88jsUT
eUTmVSvt900iW0xz7myroc4hvsYGoXiA//HwYkVvuPCUl7gX4muF2dzNY/V8Au+XNFL+m7n/Ex5O
esAe4r9ccfgP1qJ57PrXt3Cp+lQ4jUc4XdQq1MyoMxVBM0P6STYuzg3Le6r5ONoEfW05Z7G3RFYt
SWW290qmryS3/Dx6ZONwfLxN6EVZ4t3ufV3Gzb/MNdUo63Vqmt0ONhct+S39I4E34DuFQ/gX8N1E
KUEULPttYj1WHOUwxMRj88gaRs/tJtAn9umoKUO/J3PBlER5zO+26W5MVeU2TDmRoBM5rfQs6nJN
6YjYjsYhmkfaXRFAUiHxCGNWbFOYvEi+zL1Jhe7b/JuuS1jL+cqRQ1sihfddAmI2FL4BnAfdsrDB
AuBC6AUyr0ubZ4xbxLKUuF9zYAXpLgFrPm+cg4SEQF5hlPP5yT7eP8ilg6KwaqTvxWKeRFGkOHyL
/zNdCUWkJJQnKwzw4I0+NHTJd/rP4FtivPFVnSlroBf4xdxlQJtJuywQZPb7om6HgR9NA9Dp/R5b
kxmWFSD3uu28y13yb1eCD+2luar5zbWCH/EuExwOHS8/wpMxrY6w8eZoCs1YeQ7R2iQ7oiuUxNvB
VAYnMqmrVU6qaOOo+MSfT54dHr+vY3fYvyiANaN6fFqgf3kTeZ9rdYFUtIQYOvCBUKuJMZk5v7by
iU+xtlZy8lAfuCZAqp6InrHlBck3y1317t4oL3R63uZHxDt6DCdfSNHUITZpwwh4gN3gJ3aKiS9g
ra0OyNF+h6NUvFEiRu8PohdKM57uGE/wK99E+MhmreXWwdonSlIxoxz9NfIG/2YAw37Cut1rk4Ti
w28DdUxM9IHh4DPVgNVLCpugM/HHak5zq5V+a2Rg9eDq/+i6elUk3YJ0WuVgSmf8sf1iD034tFz8
/sh7nGhdWZ7DLN9DSEgPLlcP0pjRJYnak7/OVeS4VYa2aq4XpAfD52937iCgdakexgqJ9OhwolfU
qhok1AmGsvpkg7/wo3+fkuqaz7IOWEUuGU3TKLfvwQSJJ60mm+NLkJPWU7XHkT6ontT+z6qpOYXs
OSOmi1jmELoZE+zrxlMemGNzC0tdYgK7hCxZfGcV9OrMcPt1z9Gi9yZzITQFvUSya26prgkzwoV8
EytQj9FQYTczJp+6J5atpvEZrru/geuIjN0qpbALqxyDNkNnqdU9lzpgE2lPq7UDl+Lq2XUgPHBB
2DsLCh1l7zzbiW+6qPnfAxAQTzmgNuCtdrK4AzbDhubRBARw/i8eSAuKe4FwSAmM7zkRsptzRgx8
nzOdNMZ/4tuKsYZSaOt0+hg/xfnO+Sbly5vZbnfPydgNH4pwcfVEUhEyA0GeQ29jUsT9+PkfRGc1
yLF/S2qr6xFJSvG4+gVAQ0oI3yHIzOL2BQJ+dwk3T86OPXqQnRjIWB5q6BdhWnWHI+DhPhbhXcLt
10KEHVZrz1/RN3kdSt2zEBshROPOttKnGVDmUpYo+8jgbcXDRCvs+2KZEXiDP+Uoqe2vyvc//WgL
Q1TtPU8SEHhAGH0/gFKmC7UVPn4okbzLJkhSmNqtdAV8TwZxDrbKDj6f5pusUSBGXPfIGOI/VZqm
3QNaABNFVDSwtpdX1sXs48BysqOhQc7Z3gOPe9LdaE7InmVz0I7Hta3Q9vmb4XsMbC9VCflwP+iX
L5TbxZ9eaT70NBMlyh50dUXpvxtixJRRLu80ksZXVXXwNNwr345GHWhgbKVEeklP3tScUAD7CBkR
5CIjUWCD86oc5spoMO2DikaEKM0vcwV/blVORy6EYWoOpD1SUEHxM30dXgX0sNfXgwdUG314OqLq
KE91LF8PGTNk9dXU8ZAPnkzO8Nyi+8Ttjskh2U+4T76LT/yQv/SNUO4h3RCz5qLjoDVKC+vJCPac
YEMPKvIriNSJ/Eg785ZrrbTlLwbNYL4+FQYvdXOz7WtjAkwQ+Q6TRRJfHOeFBKQBw1R5SEda/Wov
vKoADHun7Nu8r3L6CrIudHUlU1P68es/I8+wg0eOHWpCbBuiPG0lxAjrpMqmkCAhhNXWLLNb1xcO
149IVETu0ePpHtLGOERxCpx4rp3IMUslkswX7ae7ZOx69jeAkJqATBCitBZc4PfMZqyIr4NzzPqO
qXGnP6SvaT2Do5dQwnsmxtJ2TtbKS3u2KVWGQiMRtaqIPHRbG2xpUS2ko9H1lZ9x9iKbnuOaBGLs
19bsxBAkTwCG7av5F3OjRYchlz2zpDKpyP5PgX1dSxmTd/XFn4C0AGP+VGLPUxHCWMKcAJPY+HkB
eg/kupu14g9pUtIAutZAm+oKUk/4e75i/0otWtIm1DWajk2lb2Y0SqeJNJsAGbQ28Sw/+DEdexBl
y3YHQBiYTD8uh05EP2XuBVQcjsHSUhRl+J1Bdwr9XDBYcIigqrVB8a81kNI5Vx8DS1Gq/O2wLKUL
um27KVkK6MpPkfleZnticI7ccVbgVEUDUCWu2/mZg25Qt6A27dgGEwkyIO/vaLIAhyDiPnH4Rzo8
4hpxrAgg+CUFQdVq1ne/HX8phk3jLsVZq2gKnY9xU6f61/ex1DGejnRSvRBfViteAOSmTUtz/m/c
nuvI77Wf+hvesPVeoO75oPaTEXXYvhDhtaDLhS3Q3TxGEGm7oghBiSlYQSG+sYLC1KBPxM6cROvL
UJsVhpq6uHv5lL4jl9tTOeKI+eodfoJhiTjSH/y4Lxcr01ofoLUs0Zmoo9gGEPcpOXYPEfwIIIZN
mZYH8LW1miK48ECAAUKdvPFxlKI+7tAyJBqETJEkE/VnT6W7qPD7L9gM2U0diNWqgTbiygyWI3xs
N6USUBqg4r6hMMoB03WfEnE4rBSBeDqf84EjQipmC0MeX8zXNLvjMFqlD8PLGiaL2bPVVq0X9ZQj
ogtfkED7DKrJK8fpkbEWx2M05HD35Np5Pjsoak2Ju1XneKKSsAORONDoAJ3Ud31z9s64BMvIarOn
h2VwbEPMRpS/DEsLijP5KoL1NZ1ir+LHCC96SSo83PuxuMtp3rW1V4NQECNcNYX2WgUYaPHbOipw
1oLSn0acWdQGxpFquJl1LmGK49cs6dzrmhBZVpP1UAOq/sRDPpVviF0S+mWX9T3ZZH1haYuYfcha
faNxbFW3qlkOeDuFo+CvXNvFwCqMysud00hws1Kw/jQgUsvgPaw0unmBFcWJsNb8Sz8Qpm/6dXRu
vbjTSDmDqboOjqjd/t/Yocu4QPF5hip2sJfL8isZcZphSUFjtoKZ34EMc7BS50s2jP39V00SCDjo
b832HafmO9V4jOyGH+JdnPNPiBh3/TTo7+mZJLn9vsIIHL7Qc/kgrzdKd1fTLzjqWn2oDMrj87RY
27aNdtTD5g2dF82dv7Q3Ub39CUzjMEeyoa+YItm0HV0hHF7KNK4MymdVOUqDKJB4yj0mMQx2UpBn
6yBvZWP5tgqwnNT6MuY90rtyzRFWwIRXHNM8k+TzvZjclRZMr/UGX5Rpn/G0CnlOxTAx4kVNASdU
FxoKz0oIjE4n879v+YKqWZhsnqFnKy8GQ6MBRGt0bKf2kPxrUJgmBqH+Y+9eUSxM5YPAf6RzXD8f
zv4QzesxwecNuvjgItAXhCk3HfQfxtXRCQbvriAY0ur5m0oJSc97eYEk2/NracY3guOBTjPIddrN
mMnrG9+TVk90nRFw1558KNUcUIMsrN9ZjgG6Nh8y+9oyKcESuf07xVIz+pjcXiXjC0yM1a8kA6HN
xbALAaOtZ2CsLU0NNwnUomAAcNfvGthI/X3hNXnZcXEyz+8qwzmg/B1DzLXiAOUvnCjuf4+i8Djt
NQN1AHzBq3EQcwvzkdjGnf2yjsMlHap0UVe2y6g6d3oYm4V1NIb2kYflSp4Z89bUlLWdmwN7Xw7G
qt/YmPf1c7ynArcvQ2/MlIi/c3hwND56gOa0IBraJBnpU8Rlvo3xFCMpuuxKh5Uya7Sgw4ZhAmif
KAWBlGnERrANBd1fQHB5plJdr+GT54M1yHMxDSSkqCY3T9SnF+jh9Dh58zZVt2ZpRyus+xbo4Zjz
pCBtcyWymwY4T3TOImTcqLI9sY6h0O4QjJ1TlEcjErPWqUoNinezuPvCOfZC0hYWI0vQPIlUswyK
prBul7t4EyrHfGxHcLzKuYc0BdF8okGmsknrjghrqWWYWwdgXj8EwqDi2awm2hyqKMxgLGAPQcqt
UvIlsIHTYjAWiDhmAgnVLZiOCmHs43j/Flb7lXqY/3R1UVbKsMc3RAAxBO5nMA1TONg4kf86+T4x
kR4As9ITMmdp0TNkwrnjOBBZIePGkdPcR3gE7AWq9xc2loBo9XjxcUxGrA/sk4GxU8LIuF9Tec/v
3BXyZLYQBi9zEu1hm1VcMcOa/KQDHeg3zRQD4qKroJ5pvSuLNroKU5tIgtfUmATdrp/QdCRkmgUk
Mz64kvgomWB6S1FGfJ+qBKIVDHJIbqSgiS2h9EHwsv3KoYut8POju1fN4BoaO75A8sEQh9G5leps
OGMHpJ37xqF52PUTG9h8xuHYJSuye9J3FxOqV5dwTfbXSCR6qD8DNttVcSsBS8NKHMSsYb/2DC1D
THyEE3NIGFAMmG629+ZJ5gef+I3k/9vW+h1Rnhr8nYweByixUCfvMTb6dYpC09V1bET835L/OXsi
KkrVHfwhStRWgt/iZpB+FNwSu6V8esqy
`protect end_protected
