-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
upfDnG7zTcHeKLOfr+l6U8DtyrpZa9tMo8MVuF+KivGL175vvDgSgOP3p5eE7pvec+Pk7vdxEAFJ
20nYqJixA82dcz55xN7gwiMxd30D4AwDQyfAhgscbGR1pLWEEewgL4TDNnfWfeNLkbPGFV9HxJkk
bLurciFz1J7haqKs0UQQOGFbeiEYk/AZpuKcmlyoj1jPxoZjcx6cjvIpSrfthlmvOMeNhZu8vUxC
xjI5a8pumU1XjfQY4TjLmM4mgYHhH2prg+5GqelvCBufxRUKXlGik3MtAJOI6U0FJtL3UQZiGQSp
okgpHo8qTicthHP5+Y1OQieXlfXxTN2MjigAAg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21168)
`protect data_block
xdtz48jcvEFFz9DcKP7k4xStN3y6apiFFa2v8aaCrml//cMwyaRRcG0cv7vFhUjhhVSUJYgozh5C
zYsU/X7D2JQQLqoRIHtfLRHQWTpRh6nBpDbUFE16Yz06r1kmEaXp65ZzyyJpfzWTQJ7LFP8Y/CpA
d98dTjfn0/oYrOvGyWfJg8ySVV4u34EZ5m693UgGBu2VRC8FcPd7IPHxK1Uj+GJ0leNli4y3Grsw
mQ6QzGfuNW9YaM4kqb3lD1rJ4UAXvHfxoYb/sEWB6/iN5F4L3E3RutvSYujMRNqeThtZ67d31zXh
juIl7CReqJY902hhhxMtEkmXDecPEr6/4lItcXYrWKOVJMnBtsCqItyrdI+F4O7KorNCsc5iH6pG
PgY/tx59EIa4mfRTj/O69K47qXgXhRgwNzUEyeQhQkzU7ZuVzawGCx9K6IeuK3M0h4CqDvOFoC0I
jLiVyanp6anow1TesVRZmErxuZA8nuTkzaqNNssiqGI1ChxGDQbbh5gjcFJaWH0YV7eH3BbjuDFA
3SR7McSDmnAShyHv2ZRW9m3PK6alccMl3Vpf5dTvJjWpQT1BDSyyjqVNHgD6WLQYsU0zP6u0GOF2
vz73zEd0cIvZzD2wUDCzTuKT88z2qNxevNxuWCnVLVrqqtMV6/x9lKP/aVYJ4R9BbEhNDBNqw+Rd
SQTtlbUtSdDrd/fJUZxHOCmQPvJaBz0SmPQOAM7PiV9r7I9Jv/d5sFDCKUmoUZ9v4dnQ5ZQMCiqc
XGoojshJPzx2SzeT5OGuWg9l/P9wNdYBWJHXmBB5fhTCMDaNEbb5W7gQFswtpMePAyQYGT4K7jHj
hURLbDUHr0CW+3hgFJLcKm8EdCm/QoIK/T37DMq+e7B7mBFmuG0Ar5DmWwq3aJgLu761XP7oBimI
sAKB9OiH3CZj+Utog/NBi/GYx/oTPRGY8WacCW4/lBoY7UmqERW3xeF0qiMYiEkHLAEOE8HqCKfg
AjV5FX8rDTVGC46R4/oEpbiS/dJ4wQLBrc6cpYI+qlzrbkNNGJZ0iHVJNBL8wEX9vpNJAKAuUxLu
wIh4zzow296iue76ImWP2Wd46U2Dk4z36anYmO88ozSSYGno3Yy0A5DBLef0po3wzKJ3515ISIrz
bZl0qqSXHVoh1CYmJ6MuZpI/Nk7hENWXjsJWW2sZcmqUnMpyyQuiCH6bYozKu+DW2ZMwYBrT+LRG
5Hzc9bk3Bz9RmkLfMjKHLXK2FOIqU2VBPt+hq0ST4rmG71Q/vAbI27aJ+p+iJqRewG/sLpbngR8h
BTqisAAP+yQ5csfU+kRk3kS5TMwJPipJUrMHtLXFUOI3+HLQcHFRdAgdeyMsLXCBWI8Ebe+ZPBT9
ZDhy5uxAZIADeChWrsHtuhLqxBlehWbNsWgI4oy8GUCBMf5eXhM7yh2nTcxvAwKI0DegMJ1xENht
WJqquLQ388tv0s0jlkuN5ET35OrtBpCxOZUHWDyFgx22of+QjLLOWmVTggKuegd869AuMRWnt5Lb
h+B2qf6fv8fokeG0R0LfAEgQwbVf9HtwYGViEbdEjztCChYKN9UAoXxjFi5QSMCs/Lqn1kWN7pT+
+by3KKuljPSXmOA3lt/1Dlo01Mk4bIgqKTpKy4XSj/MGaRdmrEs9le4jdVgg56Exz6V5LKYJc6va
a6lSSNw3kZItRr9icV/nR6WsUKwSbLvlZvhRZiLQpItuc/K8/crNcGmaNChNNScBxmKKuDYszKp1
6TajC3uk1qX8TffDnf/U3ooNlKY+kiVczHDY2S5i2nShSQ4yMJEXFbSHqhy547jrUJK1dFOXsxEz
HzDv/2oOJpcgwxpxxy+nRkCMoyarZ/rBNoxbybUTQWJ8dpVS0ZiM6xPv8knOoWGbCCalLSv24a7p
VG7tsR7BjeAcTgACS+/aNZGtntSMObC0WdqG6n1U/M2Z3bS6qsvDMZ0UiZmG9Vg79vYj6/VRW3S0
atLT7HJRZQFWgfy1rIk9tNmLgKGOvF87HjzdQvnWEi2tc6QZ0jHWihSImzgMAslK3nXmLBeCiPW1
ViV+aYmUiUH8YRL1Qcu12Qn4xEyxqe+Y+3gHi3PTLTfeFIibat1lCepDZFzFHI8LoNuSqGbLX1+L
jMreG4wSpY3jJx/psIAHsiOUt8LuNmlTK0LRKogEwMg/962AU3AqMdEadxAeVbTWaorC4W+AwsmL
C/EVXBBelZM1s9/F/nYjUursNieQU8V1ZQYqCzip3hKDClrJnAf5N3ZDDWaD+rIUHqkqL/KLTQPZ
Q8UcvPWcPYOTARS6uSQvPfAJX8rOl0eCzJDuhXQ5rVPZTnyeuMsaX8htv7iLZz8aEx3Iv6VcPX9A
CJlFnSXyRduYIsgcHTWEkqWZ6C4osctkzf/9rFU0K9DLfs36T1uggqpAHpTTvvYSRQOASWAl47Cd
Zczq8o366QJIUedTjpy8M/f8E5uXxMtY7bobrIDybs2L5IlKo11u5kLOaxK7oiNocw60FMSuPl+c
t2ZrsZUYodt6qKNZ/PryySVbfzXzfd75FKSCsmoX2C5Y3mk8Zce0LOEH80yGvOtBX23l+8zxsC9v
IiNokt2+Ofc25xhiycQt3UDG8BLU067sbZEl0BQzvoOp7Kl4CJN/RAQpfwYrMUfs61bM78m7Tr15
upxVL+SHEfSHcfaTMiEV9VRUvCIHZ42S9+tCcrWwtah9WOLsvqzsI+p7L1b/BTFrrn24Q7zNfetk
yEWCIdRQqcJMsEBfRNIHpF2G9Ldi0iAlfFsvXF3cYUaphVjGauXzKoH/ZcC2XPEI+HDPrn6pBqDl
19rtBM3nU3OkCNjurKA826uzVRUsdy/nmIB/jBQhV7O61NOwRFj1BFmVG4WPLPdQQ4oDhR4m6Yta
WMypTiZrzl7YZLU/2Liyo4PWggJhA0aoAZmrLkd4W4y9jJX40PHCwAv8AEod4WRA7BJ1ksLxfYgj
oLv0Xjq0n6DFg8haLThr96nGl9BYXMD56zuapczi0p8egIVnb1oYu3SeGpjKjxYkXX8jc7koD58W
Y2S7NS0UkdGQLMyADPMXYDFGqKR3QTFmN6XcRiR5LCyObFa06KYuTtF8HrQG3pBWAdeLVvzX3rwG
9ldQp58+zhLhwaEa6gq2IuOa8C/q51HAzl3Dz2HUqBnlseId0oCRgDJ79zj1QMarCQOZS2JyM8oX
70052zweL3pqbA1M2/yBHBt0CSRj4AKuW0MmNiOZjzTM8VoHyKBeomA9YffTA5dm7ZFfTtukUM1l
JamYJ9x0iHu1LuMZyZupmaV33kawQ71nvSQyxj6hTKw3aAwRZhiAEdIjUOhlQdyqq863SKTlAjit
a7NdRCuRKcSfvK7Ksa4cfWO7roOvWUfCQuCBKI+PLPxAUvRg66pv+913CHL4BkXnDzqc2spqbFnt
R+r18JzUxTz6IZd8ckrT8j19eIolwTxvInPoncLsWeS3ain2/8n9q1YItdgH7LFjwSq+g+9ehCHX
1hf/xGea4fXHcGYQ6cflSfV5pZnhCVlPT1zMm+eIYGL78TMtNh3q7gALsSNHuWIGuiBLlUCMi/n+
O5iU7IvtTH764BNF7LzzQSfVoUt3FFnZ+3atMCfA/sqKH3FRzoRyrwQgP9Xcp4ugFKibcpyRKByp
2oXqmw+H5xxdNcpuBXbTD/aihKC1I7XFnLn24p9qapoaF9cAJ/8H+hVvY1su0nFkHqboRIGmAa+R
mpKHPAFCUzxMGdFLq0VL8U7CpFwp3Eztyhn9fnPqmwYjmV7VrJXiJRGRgoOMh7Upcptb/8moQ1mS
Nwl9D5akTFqz9zWu4HmYnQA3bt2+kqTvEw0JU9nIn/VP3fD3hfDjAcjaqqsl/bRrI7EeqB5M/CM6
g0V0HWWdWioQExQdu8U/jEeyVdYPL9zIPMUU/nlCPe3VJe9KFqXE659Ce6wo2Cbs4DXHaYdbyaHk
biEYNkbvJrYbrcKZxhhchmxSnQYjqQvYJdnt5ans7BYRkjiauqEML4mizUR9vImnTqEpqBZjxorU
ND86zkTUgAxgVU5icLLyuXYI6+jerPYaQC7d6Ta9qpJSn9Hu2aMUvIPt0siVhF4WFCR5QxNrxt4I
Ka0KISuKKGME823xMppY+/dfCImYpzT5CwebbOZ+nlD1UhEEA6zILzhrslDHHALSD2lD64GnYX7h
zpdgAbiUyCqrugnw3bom18h6rJg61lDy2K+O3IP+ETJwvX5ZtFAnM0p4EKH6CYwJYUeebrZq1R5j
q9WO0K8LGy0h/bDJfBsPVvw4tfShDBDjhwYR13vHDmhfnvrJym039FMf1VsMy9UZ1RKUWgAfuJqK
38b39N4hkua7x9LDghmKM45sHWS7x40gWeen/EqShm+2RS4OAiyvOMELye1Py+Ik90NbsL3tQ/BI
8TU/RHgnIZfx2cuHye8D+bhqCndGfq0OBZrjgTZK2EGiba+kCgAmAItQhXdTOXB8s0lE2atCdmF3
/VDwgfujy9pYd6P9P14EZ+eeT7vhwjjM1piyyx2NTo1zwpiBMxQcoHT5pqyHGZjxqDIHdzLINh9v
HfbSibXpLKDO2b9Fjqa6TUzd5AgApCeBB4+6b7WLgRzlj8ZehIGhuxoU0w414o9GVQQaENVHvS5Y
UaYsRmo7/Fsu5QGBNE6Q9Q2Xq1LW1lnYEfbj95HDH4Z7hYDoavTKRMhetFv9/l2Ezc8ApppNC/79
ITjGI6yZ04nHqdmtD9Cle2Z9xkhy1+BkdNttMHLU87UZ18NepoCeo9UqKZck1i6nS4ObgpWpPn9H
iT1KzAQsCfd0cS0NC9FpcMn/36uq8pc0BaY4OTtxBmkUCaaMZh1VpjQN1830p+R9MfGWZhN7Ki5X
lSi4cFVIFO0Xkhs96SBuPQDUrqbofgpCmuGlQ1GNUB2sjUFeYntBh5WcuczXwITeDccEC8xVpV06
zLmBYEYlKvN0PIq856Jn/aMKbeJF6yzql6hIDXqE2HI3vNnd8Q1XVk8f6drjhQgEjrNBU55V32LT
tJasJ3O6OldIfMKb4syar66an82Gs5eU5x3rKKmqGrHsX/SbG4dVTU6snrgM2jiaHr89bTnFHIwH
WDpdHHLAYwygd71Bkw9KFKC5IZG0pvJ2S6LFbuozV3R2GBQrMMKS9Kvdrfj+MNqIp9BlgntCK3S6
NvbjJWJCUS1UYG1eR3DzFKy2VArrLp3Lm9hKCLRuNqONKmtaNkUhsmIox+Piybw6wO/XsDBBwFPl
MKCbhtIMlq1FIK3auaBYghgpJShhBzYy3LyN4uu3pxxYgA32gTOKWzEBaKaVuAfJWFZBP2oZfu2T
P8Ipd8cL8Xg2QRXX5LGqDU4s61gSxVHWkyn7iPOvkk02vh8QwUK+e8aktKZnABtmMLMlVw2iR7qf
1MkyuW6L+VPm5ywV/h2TM3rbBxdZMDCsXttfsXBLaFb9wrA3Zlqw5VRD5X2O6dvtFRnJKgoCQBA0
1bZ79yPMb8lWSe1y91rExfYsv0TAU5uAj1eCUe8qOdrgr3sUrKmvJAFY44PcJMCrmh8mQG8Ez6jr
0Xm9h0RLFlAmUhHFPlM69H7lncNFkwq+0Jn1b4qTntD/nvsbqe4pi78kIKbjI4FtUTzlafsPkiek
k1dEHaiVrW0rOMeHKLHysd6tiyNlH9abVRmJwwXyPgT9lNccifNqoJ97BxPloLBQh1mUpQTBrEys
dO89/wUsnXL7KXLoRzCEB8sKhn7/zqnF32lAO5rzdTfSiwivWF8ADoObddXqwHONTBzEliYZ/5fs
GtnfhSf5ptr3pwRMZCyw+Zfjo1Gr5VFxYgXbAvONYxbAjyqLAMB6QGISQehbgNIdaIkQiAmI9LoT
OpceicI1LDzQY1SIZhtgziAEEZn1Zy3ZU+XqQGXzgz9Vp7Y//lfO7hzCUysX/e9FgS+APz4x7T6a
pw/Y4wz7F1zL5jauckaDm324bHo9tNnpARJC0bDKILs8HSbH+TN/jMj5O94+eFwiIT6NxU5mIRBV
ybxNw6Em5g3yODGarhVZYjxbgc5vTq3W21/VXzDpnCHz9fjs75GXlgYHVUpfJLRX9btMFyy5MtuC
TGgx4hXHKhUsDufyREE7cY6ErXgRJrQZJrsXXcazrKJFXgL7Qp1m+/5xfCz+2fVRCjyVtKFqul3F
Bug9kue5Xa3ucHAfQIfXn63iuJ1xUpiuxHWPXogY84Kqu6N3oQa0GYSzLZpi4bHpQwkpXWsHbtQC
+7P/ABEx5OPalspUzXon/boUqrnX+fxxa8vN1M9wUQKMyYIAckbr8GxirWDE+D25c0mkDO5tVSmT
Wykmpt5sd6ix6zAh4NJ/xtzTsVPyTtB91R/36a8jEpqiWcq07ZDtpiOR0VIa8xYT7KttUiDpCjou
DXvUTXiaFBjJcrlsXbVXEEjy5sfOnzzQyjIBa2kshFI8RtV5KlZilXEvIk4OduhZd95POVn29F0O
EQFQYoub37dKK3xUwhsGosobpkoIXzRpjjQyeDBuOPhdOlBqeFpzChUS195cyRn6ACyjafidF4pE
kh69u9NIvGpQgg1Vk9JuUrBhoV3GBEYaQoqS5G4zMds3TuTLPcitBU3LZ8ecy6GDzbfitqkG3ne5
P7flQ2438e8tT6vY2EamuLGY4BqJW9QSxWqrVVJNbj27vJT2JT3+s5RQ0PAvX+yPI+KQs2NPzj8T
E9byKgiHKLJR0u7YSFyI2JvwvTSzr4PD4fyiQ2+fnZXHWh7hjWDYG5sZ84ft1OqwfT7e38S8FWba
qwXU+Td6qyihYRM2QD62f0Wv+9K1eKEdlgbHgkCK02Au8BKciEnqoAjnJzNzeOV6X/VNNKxh6huu
rFOI23nswG70RRJNcum9BCQ5pLtadDVamEm6POQwY2B8a7HqHZfK8D63IDgHK33IFSfyhqQGSCJ7
AgzE/FWR5uXxe/YLCrCHqs7+r+21fqf5UPfaaT6sKG3DeR+TloK1toEjw/OjV0AdNPlW8HtD03Kk
96AAUa74E6tVO4VyN449MXTqvk0QjOLazPsNuPrPcIrCzPUUcx0o7TiLcBHi9uCDY+6v7ayHPy9F
GMU9g8A92PMiCpVSU3RK9h/Hkn0vttzZfsHJhpQtD3XikkwT2eoYq+dbwn1H6YRltPwiO5EhGnja
ZLqY+0bDBsQff0VeLaTdWnNFp6C3kL3BF8VE6xS53CdVC2I+U05c44ydWznVPc95a+vyIn3jZ4qZ
6JbsMtRgNmLeRNQc31p7SuUTca9f3j/j1du1dESJMrTX0jB/wo+pB1WO0Jtqr/qCXgI5O3WNAKjC
z483MFJra/bIVzT0IpWrf3UEq/dx+W7f8xni8kLXfotzGQ72MJDxk0k8J56NJPbEjyfEspbVlHKE
Ual+ixSEAd7C0YFXzAMF2IfHqYGPmQg1wsld2TOy9c2w/CZeVuSm9WqKDmQepKapQaZ0J9e3sZfs
sdvWCvS86yQfN0kkeMW3ex7JZMHOEL1UWh2rU51c/YgD7QMYT2AsoY/EUolgXG9U52DI25Siogve
MNZ+a60YpcZLAWiuj5rgEU2Hi6MYUT3NsMokh2tFumwTaFoNC7gvHZtwDG7vIUVW3gM5OXf7WKmE
Iz2mrIC48cbOhgLarOOxhZ7kZJxQaXt0LKJR4YmNeGRbAdPVpwzlCOAyka+eHbg+0f3OkFb5Izbs
SlUY5ZvrW9Fn1fazlw8r5c5ggtT1fmavnOvLzY5sa9dzSXX17q8qU3+yV6RKWe07XJH7Ci4rXI/C
g+3xaP5eGV5JBGX100IMZohTe5qVHkQAMbKEewjb5wSKHeCRi0SPrtkZzJgOWW6iNE0ZYn3anqxl
/StzvP1sdnLxbgWMRWSe5OtE63Jr/WIJIU8PatpIJ+Zdb0N9GkrzPB0TO7sDb2C5PmMwGi8MqUqr
Rzm3HPs8gSxN0kJ/3RjCIz7z9Cw3wVpfdPjpNl258k2IdHt53r0K5ea73gFA3VSZrAPVR1G1qfre
NaGFSoD4WBYUTahfTDFp3fBLTngiz3MZTmwL5qCW2YcGsTrsDS44H8E+vy4NtgLVG+oUHVmjEsjb
9MG8w+sX15IINQVtZYY/7zpn4wcoh/cDuncxoE4EgQWkKGyvr2FijfUqnQSeOA/GR/c+Q3Z69jZ3
4plyY5MYN4VbZV9emORE/YMRhFHMPj2csKiTcuBEXMsnhF0EK/6FSqjvftHMUgE6chkS2hBtjuc1
vx2iEE7k7XDxnjyGvSmT0Td5DsEN1D1x7moRRdBDlM4T+Ss84nc0kQPZ836ecgGueisBrCxWLx16
BkP4exQSSK8aFFqY170dAlzamDH2uc2cEbsZqlz/pHPme5gVo0z7bk8ObK5S8f7wrJvid5Hsi0/Z
jIOUr6ViRDkjwZhxgXUapBtGGwm0gk/ULC4xbuLUrz0UxBhyYu9Pg7akjnVZJ4/vNlZ5N8ukvyK7
hVHoVU9cdEIUTtqpzm4NKWJ0Y4Ghk8o+SnduuWTOXxZZNBNHaQntSdPiWgevV68Q0pS5UkFyFvEU
bx/MH+kVo+TNsvVvMJJ6aOJUCdkiGUlgmrGQ0zz+lh9CxD4nZS5+FyVy/0qKC5s0qDmH3Nyt03Ux
5yzVYsB6WkHIXYFEh0azHbCzcDB6jE49B6/OIBKp/Qtv+HSiXzD+7XV6P4lFmCJ4w0F3y3jZCR6c
hlUdCV6HWsWokH5p9uvqJtQXXrvBm0a5uwZrB/JfDiggFir8pHpmQ60UEPswJyCCJ+TOTLFcsGnG
1Aj5ZIycbl2VthTlEH7+/VuwEj30EHJAxuHh7zvzu9cA0SclVfjKohkULbKT4eqd7BDCJmzJB2HQ
vo7dlKGb1M5gtr47ej0rReDOiE+u+Mic7LS2FfWNUaRrc17s0XxnT8nBa+GMUjXBQELvn34sggxk
7HmqaX59+g9q1KoChZULNB9TdnaYL1IfSFMzGc1tcEWXuZDMAak5I2SGa0i/xS1/4xROe7ULRFPj
7Aqfs49xwhEAXo79eGSEQo8SVviPWBeikk6YMdsbWcpSm0UDNedqcu7/RKHv4Yl53XqUbQSBHc33
gxrZsj1uOzuKmFRHrnmfy8GNuIKLI6T3xr/Fmyh2mHpcMf6cNCSZPOcmcizRsprfACqs0H5QB+cY
YVqqsK/tKb3TqXVrHbL5WpUX9cTe5lNHNhhkFvMIEOk22B9OkSB55jkMGv2LJRyleoOho/QjN7ZP
KAuA+ERaRi3AgButfR/hRgn/BpUDa+tJirUjbMFJrb/CQLyyR+wRHtgHlfYU7CXajM5d2xh6xWQw
g1MOJWnORHLwvou6b96Q4j5auVXe3mYM4JyTUxZB9uXSSbWHr0BSRlvUbtqtXwJ8BmZ3ZIr1vQKn
7d5QIpZL0hgHtIKiVSCkBXUWaheGQ5H+5TlRq2U5A3N4jyJoJ7MSaVy4Z7bncfTfLQHuYcwiENW9
1EL0Qx2IxcLRgf6U0GmxKwrPxmrbHw0BdvZuxHcGq9/zQoaIRyHOxTcdPhBZZtlDgDo1w+0FbrvN
u4rxyu3ujP/6tigPeMLURYjp8s6A2QHSSf5cR33BtfiKrA2hK3Qcy5QM8dRp0hQe01Sk0mPtxN9I
9MosryyUmuLXfjpBEsiaHAeswUwqwGSNmsVX6wvxhYs4O977hlR2tEm0rfEFkFKt3d8QmF9gF+iF
6Krxpwctl/jQqvJLpoW61cy9k30U1VlPyJU/b9bnHSFwncyByj2uDpLMHt4El/kCzvmcPDOmo1j7
ab2+6JXoAbxl5bFROe+VaZBBl3DoLUPPjHg+FhGBpIZC1Xxbbe5aIExCH0euHAuNP3tKB1yjIkjC
LQvtvSz1wMb479lta5YmpmH9DXM5g0mbj/FdzsFRwfB0gDS3fFc6Jw70vN5i7zoOA7y1yonG1N0j
A2ks59mGFGlY5RYF3SDb2pEQF2xYBFeKoTRyWQVC4qVdZB7sjy6PaJtjxLdyZ7u8zOfYjIXC53N0
w1ZCJLKrlliqHoTL0p8qYyXg5HHvp4W7QcuVeU4zGz+sPT6Dk25QUtBJ1roNnb73nWhsh9YDUywT
IWGprmwuHJFVQ6rriazw9Fg+ldUTkaQiM9HXH7ZinNfNtWKwwDslRv7RpPvX7qq/elUO6b0ixGTw
umzuayM+ZTsGoNXpHi0mPlnoSTYQHSfsV+vz1KcD3c2YnkuAtDkbNhRR1iFZThakSdYgiGCewkHb
U5Y2wl8SXqyQPZACIZkq9t9Q5paOtNJYVfe2fM75+vbPzc3sYdraA5pjcF2qjHw+aYDrr033IEpQ
fI/M/1afXGh7vL/O9ueNgmSyBohno7CJJTR3j9JJqM3PsmFIA+5Fm8I5kMWMkQSXlsgHbJGMRKsr
LqEGD2XtinbQVCQaPO5ouD0qj8a6opm+sP2Cw2cAvsd1BEpd9pqrTOzXpj6E43ujfSLYTJDGS2Tp
PEYYTaryfm2x+AYV/gLXykPyNl5RJJJ39m9eGuU8U090Ifmdir2+Rjf7oSUIafwLYaDRDhDi739L
fW50rnNRi7i1Vx5j7E2qmiFyFzqxJeR4RQJ3CUhfJvYAT+jH5FSxagmMu3Y3Oh4SdYATvtWD/SPB
/VzBFNnIvhNTf5FXK7sShvQ8n5fG6ft69DZPDHXt+LuGM6wUJeAORmTVXGaGgwOWD3N+VopJO6ag
opNV/3gQjPfh6YaLiYpJvFrctLWYosgJcI4E01+spMj0DNBWVlbgCBeji+ovoabJXddtDv9ynL64
fRFdVm/QFmkmKoo+RanhF0mlqydba91KI3EpfFf9czni4Oe344pzypykGgsOm3QTP5TsuYZau17e
IJT7eM98qkYBddU7zblbDAAeRe4xbZo7YJ6ixJDh5iSzTglz/lp7pu/Hb0w7XDRvyP7osf1U/e99
tcPp/E9FiFrQ40u/ydmeE8L3IrPE32DDJk33f5AwixChTqD9FfikRbajK+0reSUonI5sQv6kJh4R
CvZY4z4V866tEg/j5pgHV+EGpemSKfKkoAt9EdwZ3oxdpBpohqIlXbW8sBoQP0Q5tNRC7SY/5OWm
JxdVzuMnF5IfX80EZIrkMvb0oWShdWAYxeUPVuxXuU9hw4M0GAYIeYbpW0F0XF2z2HANr504YHxH
Hi8b7KCV9LJLs9Vp1fpy5O/jbFUAMMli5sJWX60Cc/3fDsAR10LrEckTNX7yQz/rlZHf9w1+dgCm
XXtUsP59H8hLzFJOtIhM6hw9yX5DMeGJEYZLfhFyj38I3iemmm1I8aL8MOOMUxcPL9OVZfLYpK1o
BFfcsl/lkm+TNsnsGRnnSAg0aZJVHm3rceglI5uHEuY7DSdgHewdJRzUcYFWj4uMsD15EQ8Ys86d
3+pu/JA+yhWAbypkyekdrb2z0ID+B+dCmufrEenxwOJDnc1ZD2N5yHjkECM2B8AlMGBE0k/44L+R
LFJDp1Y7zXv2PpsUDAI3uK4ei6N2jFTyTKkJx0Yb5w6Q4QfEKl8wg/re4Xp4FMQrjxCZVkpP8qwS
iL21jJbFj3InJ/RsEAtAUZCM0pmcFxJZYhnfNLZGhKCOyysHELpAWX5JECoBo14Qe7IoFPwZTc87
mri976uYTaBlSlsSjcCZlW0cJYRGWQF97OUzl2BHxd+fzPgd6XuHm/hnzLxLAvzOYvEHrSPlxxE/
60PnASp28bzHz3itllwDOlJfQ6XKrZ+xFKjTdxYkcqElLzIDBYmYacS6GGJzozSYnBRFiDdO5iol
UNQMQ35ODL/Q9CM99zeCDbPiEcUtIKEBmYCR74+uIMRRgy6sJ3R4eHq9LGXsTDuX/7hLVBeiVIc8
VEpmB1i6/TyY1I5oiG1+uFoaEOs/z0IxI6qOsaBKvubgqYJVsWou0fBmNH4auSd7PGpwwp27hWxQ
scnrZse+ld5wv2fz8I4HVllJ9ofql2+jSYILsSug4xJcJ6IBw4epZla9/O5s1BgYykUOm4CegZPB
XsTLyczzvibKcRX4uVUmqqvisCDYomck9qMVVieuRPmhfr2OFsDbLtdoE+6gWMDeTnj3mdnQ13B6
pTN9GUYklu7Dbl7U+P/Pzg7do+i0M0yonfDDbkhnbmlOPwn1EWCxn+aTTFaaiFp/ANdnhLqhwbwe
F5aHWaMK3pqM/KJGEMCytLb8DKqP9++CS8vC83XjnJA/UCt/qn/QN/ne7ehqvnFMlBaKxFLg1our
nX8O66X1Jgxu60ybubd/oDQIVP3jE7eFI03pufNe6OUACKX2CkQwSmce08eKIYG+QXMT+jzXoszK
M1O5+x0xqXPiBsomz6uGLqIbzKsERWcqHmTzgWwf4/a56ilYJfzWlQUjuUJSaiWsen1wA1B44/B1
XjyB5mwqFvN4FajtUeTMWNLRgP7npDl72Nuwba6M4tEM2tPEEZnx+EjW9YArkCVhZ/xl78Iy7gqv
8XaSFqryJGNPmZ9fiVT+j0VMMnVol0e7y3yCMlCvX5UMvJIYaiu9jQkbUog27UM0/+AEnl+gNnng
L7Futl4DeQ0j+lkM/Ue3gyR4G8tficnqbqCuf1L7knflxMHgKWkj6uZuUjpL3iQxVO+ZCaTmIXHT
gSZuE8kSFSOM6EloTLMu8x3LaZ0dEFV4s+A47z7qk+hDGsfLUh/fL9mb/lk7uTaC+CLHRH2TDrn6
43hwNiS+25cdlwaE0stS2+tKAuyMDMoJgMJ6TXVHi6sNb4gXOfSZ+CIU3JtnGqMf8/tooZgGHPzK
qSoPXO1+WoylncCY8sbg+BZW0z84cZdhRHKdPUO2hh+h/JnO7ynR2Ax4J7FnXzNVSwzmkXHkLEvw
NngvIwKht3UamNIjJWxTOOx0MJCm6fUfEC3F/NTnVmice8bNyxORQ/aXl1hiD12BY+Xx7VCEjsqr
nkURJK7ie2+K27eGNrGn30wd99hfKhpUMlbdwyD4OVeRFsTPqYgrrVx8eDPtumLnsr6gyEp+MBqC
s4308XQ3ZXWK4MbRUi65x5zkMaJB4irbr52hY2atln22L9J8h3cdF8+jxZ1paAEdMZclZN1hUAxn
C2Ta0wytGX8wALTVyBmllkNemigzX6jHGoPzIAArr7rud6dpqoti/MHyTQsh4kN0nnpnXz5FSMcD
VJbTBYoG9XYqkPeH+QUyIU0wHXXoTGBOH+wTyHbLtGYC6WtdsFlHXVnuMWv1nlo3RX7lFBhXEsXK
Ldcu4ucbtuuEKGhVFG8CAFrS8re4YOhoh/TfntfZeJUOFEhpcE5Xa3Uwf9/uAKpyQ8g/7p8eAVk6
+ngPnN20l4/Iy99dt+SXS4rRFbefFLGLbux6YaMj4SN7+z7utiaz6shECK1UmfZfK8LBY3VC+nnN
xG/tZaI854f4Z3qXDlCnD6FZAr3dBPwNaPmp5dY9iuojrNqt9GGUpv9kGql+Tc/jUTSuEGnVjoXa
N0mT3Lw8iWcYGwKah75J1PNqtZXMQZBxX6N0RMZjDdUs8tztlAQsBfwxrrU/eAV8x+dWXKrhvS+S
ZjiGxHpzm6YlfF00765RnjccTitNWoJhDbl0J6qENlpQULsLCQQ1A2Tovx1RoiQ+pR1dj7fGpxk8
J+0MpCDBhZWwmcaOAq5JTGddHxOY0BxHuxvyDvmqGgg37NHpps+4DLW9OOEt1dApIqrTaUiGzW2K
vV0pYSeZQodFTit69RtCVs5ky8achEYgLIWCfuF0btZJhVsh+YPk3BLP8vteehej2jiiVJ7D0ATY
aU8THgjxCch1Jik5CgLLWtXBiDIO+fPqZWYJv87HfIYvdAhzNXHXGbECtcyJib18/bC7lj1duPER
EmzhxFwrneX+H27IxJRt8NVdBLMXfavvrVlLoE3ImToyY7fyelaa1UPKuT/J4z0T2+9U9YVPNBi7
mdniefl10yhnJWpIn1prAqLjyzEdVXSK2pPuhV0IS7zvYvFP6jWK1f8FVuw13eVjJ5RqEKBp86Ho
5sNauL76+WjAfc5yayP3K4xXBlvc8zVI2mls2rdTuhKE8XYZTuWzPGywjbBGZWi0V+2O2i7ZpsYI
AeQTOIF452spHhp4I6p/xVqRFhKWw4RN64IjAUmLCsmzxV7Qa0Z398IwRF7BU3U1CF0rJ7VvDwm1
LFv0UkrstXiymwPq2eN02aDqDlsYva3a9sXeVAvcDdB96SGeN8pyxiFz5n51YKxQfyHxy6NmpZ+c
MyacA0BJfN31MNmtB0swQREKNd2u++YXut6+AqMtexpHbdqLA736MXgh9+1kEKOlIp0sljWsnsjZ
AS1P1aUA24ZS+9e0iwqJ2xfc1AXnibe15Q0Kr+3licIZOnr1h4TaRewpU2qHRTaCFU5X1k3jJ/NX
B1pCagY40FKKip+cd0GFKeKEHZdV07Kb1O6GiCaeyxBfS0ZBlfSR8Jdg7tQONcGXGXC7Pt/HcqFu
kFis5JpEhQn/e8B2TtcvQq3VHAu6KpdryfkMGxD9YiajnOMoe5Bb8Df4P3h/kAET3Cv0TC53IJ2C
aJcVntquOI4yt24AKKutdYHGMG8ImSSMQMnt/UWAmQh1Hs2fHf/kGwbs4ndPdKbXAqvpQeLM1j3s
It59Ol1c906XV7DwhkcWna4b20XxTaIUD+E8HZDpgKHErQDBkBCMJqs1r2xftPTFBGLcIQjlLvxl
TN7Hzd5udIbmvQUa5zIyxfwISHMmL30OaYL88CCbPL8T7BfCRIGW6fbr+ujOLGvCy6VLcLFwD8Xt
8F5CssqMixEHJfWG63aXbG0/JsiXC1eB0Sl1kGZ6Ac3XY96YFODfPtzc5+Bu+p3hNk09zbV/IRVS
Y8u0D2WUL/UtdljgZvMyoB+hfsIhV/HmT4T52qtiIl4dkMAgbCWLVy5VuXmgPYusn/XR4zUZKnQ/
CDiX62lrqCrKVAa+lapuHq+fHDQ9h6rIdyYNauQNu2lNt4QjrW3djb3zIbA5N1gqdS26+X1idh1H
yoxVVLPCfVKZ2fPCuL4zsPSq5SDw0SfPCHE5wcLqRSegPaTFj/4Q2W06DnKv46bYgcPyBw+UIHIm
3KT/pEKDgnGKvEDhFoZkuiTsE5iyTuo6Z+D0rMD//3ezGLThWc1Vh2YTJXi2JVp6QLpdwDJ581d8
WuHiOt4BFQ56V6wVT5tOkLgq344BkBDIAr6+YtEy6t+RRDazZHkseEYpXICcG0/ID5zG9JDl/Uq3
JuFNriYvLcAM/WWg1l5A/IYEyvb17gQjp3FfVqRWlknCQR+4TfQgUcPk5pI7feV61gfARRJtvAKC
VAzor3nHkJgVfbB+/l36TGygGbdoNIp6+hzXO6OubekExQhnfKGHAiZPeRLh3gPdSZH50/mOSn0m
Zoz0MfEzf+NBnQ+NmuVNU7jI3xhr52MXAh9PVtg33/c59P7Z8v2JAV366UB8ZAZInZKpudoLnpOz
lv0efbVHZStdh+0kpRZt7dbjH9xqYDEUMMZNW/CLALQNvDgAahESNlOmWDgjkuYa8qjw9oanQqNT
KQwjkwhxP2C6I/11NxqwrLDatXwMEJ1NIoRjrIsivo4ebC7QXFrq5doOB/HeoqTFhHZZ1J/A4VHA
n/hmPxgux8aTuKQa5aonbUXO/9KjFeXo6afddNXZ2/+mP0jufjpY6gG3risf9P7zgXTvYi4/0j/x
jIU3iH/3b83df59K2naOhghoDJaLob6dHH9PWj5n5xWi4uQybvvbflA+TwfQ1Vgdm1T1kQGBYmRb
G7+97C5tD+ZbUfrIbP5/imQO50mp8BUQrhH64KkQw6UbjpdiQ4M6kCvtj+rWu2yZIaYv94LXD6vF
E95ushDydx7kFE/t7u/1pU6sRY+s1jAdk6huqNLycyyjp4r1X+f91FQnqwHw+OiCKolNCg4DmPAk
DBF2TpT7IeoFqLDq5M9PbEmHgtTxu7hMSR/oicZ3uSVEZ6V8iIRu+icZ8P97wfcEJoDdGqlcGHnq
AMWsN4u3IE99fD3QLCkyEVWWKfyWEm2GtxpTv0JgY2oQTL9CmSOPIw2YxtQnATfbZ4V3yO4He5Nn
H8AEhDwN7w4WLOLg3WeLiEv3SK9R0ZviaelPFs1NDTw70zPsPfiQr2mv94pAV1H8l5H3HzKVYwXi
jYleb5p0qLnQ2b3UEFiAGz8BIAo8N6yvOySY5G/rMYqlFrWL2mwSwxzIgiTcKL1p9pFbA/B3EKze
8rX/N+WTPaN/GvDecS79AycXwhYRPBdqtqq9P+wyBWHFW3VDll3EP4FcLekjLirhVc3ZUwu1eJGL
IbZd3MDQwbIDDbQa7+8yguSkRD63QMVOPWiwrkzRsIZJ+lWw1TTtUDqUxZklARPV2Vp6El+3QkDB
ud+78Bb7hb9V/XY+Tpl3N4g45lnkutLS3+KU+WlLBi/ONcDPHMRQEe/LacUdCofYOkeDTYsIXNev
ovjb74aNFkDeQ7Nkquhv70qnv04+64XkU3sqsZkV72TN0ZdVPgF6GHcvLKcDvaQvPLyi6wI3q1CA
rn6uOEQg25IYzaU4edHdRVekP3ybEeB8+0Vs3zckNq5zcQDNHp8ULht4DJdU96mDCetcWaG4kQ12
Y3tAqGBuAus+bskDl04wejvcslk4n4Ez4zcNxvApeapxc3tdA0aCR8ycKuyaNSw+811ZMwrZezFz
iZJOxNGOJ3tmFpbB8XchCb1NfxaAnN8LOGUlEpHwwpX8kdaLzKQ7N698kCbKGwBPiunmzcxB2PVm
N+zCsq6XsdxfGhclFp2B1v7RHiK0Js2T1NP9sHlIIcYcEVe00n3ax3/AFWuUR9PMFJtUukOAwX9l
eyrC2MGISzTTZ/jshAWccQV02rbRC3iP6M/OLFFvlIe+oBT0tK7YBxLoQnJ//MgEPxO27/6tTDVH
vCSEckVM5sYlBX8wnDW2KLy/GF9LIOwrH2Dg/NOGCIkaEgTWsNcPEZxRpjquO4dLnWqJNT0spbq5
LBrZcZqca+tT0px5OAvjbHNJWwzilitNT+OpmZPIbJfbIftwSANwQL2Bb7Avqw2wAlwf7KKh+5Sn
D+DJPfLExJu3bygqxnt2pj/I/IMdCsaREu8P8yPmAN/8Re5AZfXAhqod8jWfefPtj9/emNapOWFy
hVdbVTV09JZcU5De/67IOkPaAwIBFODIeM9z8nDvjok0Dua3CqTSHwHjdr4zXj4lu/solWcXTQHy
mB2oVD3E6bf+kMIJLqDzETtnos6Oci0PJz0S4SQGwTNbRP4IiTCwGCNaKYgb5HI4sM5ErCaettjb
XKyYbQjneOeRWthtwtyWSASPWqSHv08ITsn3yzyFDmrGTWkzio+5G9UZ7jlNpjt5Mj0y3/kOeRnv
5pD0TTAuR1j2G0bZxHKmnqb6g7d2xV/+BzAaUF79pGsR2lhl/OqVaVND8Q47VSHbVC1tYg/ajjD9
x7XQCW4v+8tgzOup92c1CXaC2eWY+dafseX7HaN73892uUD2vtuXi88JoiToEaQzqqDvHcivtrad
1OXyYlerExET2AWPYE9N7KZsn8yW1Oz99BPHRjzy2FS79LaZjVGtWWcm3IasM2+gWbWCUzjr7Vhe
MzM9PIvCA7tvhmDfepTK2PwQ0YOlOy6hPK5wcduforro1cwLMgJnePFIx9P5ysmEzmkW1EEqNrEB
cEt/U+zWAeZPDAJL4AT7vYjvr+HV1SVZUNOzpZFGDRtqMv5N9P/O2SwTAgIjTtOyoHnpf/49hRtN
TL8OQ/03ZgmaEK1DhLsgnlO14/E6x9Y6Enmj46vcZ3uk8bAWRN2aEre6OgELxMLkREkX69vG/T/M
JsWJr2lRuJLDFiA7TOUwZK/oRt8Cc4b/bOE1FOl5vGEJiIc8zEDYMUnt12uZfxdc9JWvNWl6tRjW
bnTPmBl0fN2/BKY1T6UVXWTj2t7/rU42+Sut1TyQkL8/7hBYzXNMzeeISRHq+uISuQ+G44Bnbkza
0yvdJpxnDx1oDqD2dsim+9DqMecPxujtK1wuhfBD2rYM1btHyjMQgkZ2ZraoQACTixjHzafyUQKV
VLqbe8CrIbPubRWLqDuEEycwMLebJUURo9WTzt2xusBh8QPzNv9r7Tf+RFSGXJBWc8e+/1kfaJoA
1ItGOTafRexTfJNDSIZojc97J53fhE15mRkm+VzpwSAOSHd46cGPYLBPSmkwcOEOHyK74NUQETtW
7mvYr5vws80cC34H1S6H/6Gy8x7pkFHt7M8tpSdj9mva0iW3FX7uHgCpPHhbIgvKROEWJKQYQaDC
nd+TlcOh3bGHPt2OPGQy8THJxPrR9c6HkV90Y0qhFRNrzaHtWWerH4h5+8gwaBmQhGnUZwLtc+VU
9svs7/INijPtZi2+JqYM7hVctDNvH47hZJDGbmKtp3Fqk7k3tSOBu906y0jA2uhTaYCURjqNDjoq
f92eVRwNAiKT5Fzd2QjbvjIBEEab6fdPAM9aTTt2zuLK7QwZHrYeBsRl7QlzFNREjDXUdz3YGX53
VSH6sbT/x+EOYlS/gMwooJqTQU6/z+05sLw8Me1rg3I6v1wHOApoUrW7mQprZXCMeMHOmyhSdppw
kW6tPY0JYUoZRN7MCgjSuy6BLb0vBt8I916dK0kVMYMDspEydfiYSKA/9u9bZONNvqnJRSU0S2dL
CGHIyOwaFy483/nawqURqwH4MhWfk9336/E/LVvddJ1ubnEVokFq75zQcnCxWTHefuL61vq8+0xJ
en/TofHtW7Wo9beKI0APZssELAqht7ZwlJoD9tSgH3wy3CToS7+0PxxMOu5cJRMIkiK9D4x6gEiw
4KGqrxXCtFyZ0VATmA9wNYxapgDndmuFSPPkhj3Ro5snOxIHZd4X+GW4+WCYwNTZjFQNq34Z39zQ
Zrb3Vjk+xbkDGWqvr5eJ4HwxG0EGw71oSeZ/JJYmKuJ4nT6XL/6SOX9qSY63KIKHi8B7JUs/jvFz
MjPO5ogAKwJHgFoaHyyTS+vLq1p5OqpTNqM3oGGEaD+QQ3KijhE80w3nmaasX9Z/0RUL719w3f80
1D3rEqb56CVGskvZnjp1VfJw5mnEnpfOvc8KK/y/hqWXYMkS0ADkBfIBtafRalyJtEfC70451ipH
9EAiQUw+FkrycwsEXmTomGxMBug3CIQiBK0KpDTSnMK4u1M4A8NSzqQljnNXtSg41Y82mZulk1Vz
zTiLnbFl9+z6JsMdXlgOaDjZgd6/7qzpQeeSighgvH2A7rKGBY3S0EE5QzOyyT/8BH/cx1yKsZLi
YLa+EoAXJx3aAg827jN7PsApGBjBSDLuswAhS1iCDdGtYIlLbimSwug7EbYrCmv3ZNoK+/cm8wlZ
ApRqT3h392HHZEq/Hed12NJWIPTctWYsM7AO3fvXwXloZ5oyi/Wo6GQ7G/OqXkzaJ1qOt3x6wRxB
BY6Wc/rzYgtcimcwTO++iRSLW9vOCdEH95ZbA13ROBDNTj6feSo0WUmiUuwG3JVMMPLuc0ov7hkt
SHfD+e6Bb2YemwQC6nfyMatQRfHKOGutaMo86xBh/v43dH9x92K5bf7+sdrhwaPa6cTQv02RbkEV
grnO2/d8r0SREox/rimojPUI+gksG7aYWwyQU59a6UtPsiRNkaLxuKZOwFS+gTIdgVg5N+6YE2AE
RWAxW0yEumLpvIhy2GmrJGindRvLLZPIF2f5H4hjLYLoO0LSP1v0HqzUMrLDhkYLYoroYBO7c3v2
HUNHpTbq46Wv43besu1r18nr5+HSIQb3hy3jp+e/FUbIfKZBt+Vb07x/HS8rgw+G4arShaK+IqLC
T6d1tjGJMw7Zs1JwGwlr8hPod3b821ADHSE43uzgBSgWsPl6k54anEwJtSYja+QYjHBuCn7TXwVS
8bRZA3dSDJjeqYG+F61fUCSG7UUUoUPzZ3uxfq1Gu5sM7UKdIEkeD5xXEf75ztNe1eJxMeW/MXch
0cb2JlSEtVBlwd2tia/AJjtkogFlWQseRFOh2PUcKsCl83greVDPkSoi+lbopxp2dXmwZGjBcUFD
CwCuSRC3Ozadr7Pu78SeUxFkuQMa3g2VT9WKdgteF042yGU4oEVlzwMw/XNYxh/HvP9BlwqM7joR
duLm2X4AEa0JQxcSZkEpsKmTZSKgokZugH7sbrNlRcpDkfRWBipQbwVfnf4j7iVYOuVRx3gsCVvh
gN9g9ewvr/xd2emVhNSKz3WBpx7m6C8ngn/WcBkkjXUHDWZBtZm+pa9Ufkjw1vkuN9fN0ixTBgb1
RML/TG/xHXWb8nJRjA7+MWBSlVURQsy7cowTp+SXiY8lpIR8ZWVbi/xloeWT/Q94jPcH6sYyUG1G
9sBmLgtfQjbrDVN/au4KMBYmzXth80kYgw9AEO3Jh4Resb+I/MAxjwVgix1L6i1qGCrGJw3k/Oj8
MJfDOSUtrKKVhtXczz7Pskl/i4GxYtxo2AwomnZ+1xp6JdTDFqYSfhvI5Kyrtn5NxjlzYNXmyL44
GA4PpZgO6NHTELLsWgUiHL/ofzdyZLNjDXiduBzrHebgvz5iDxCsi6bUuC0/8+Q1OymxSHwgafZa
llVmi8hMo7RcLnYmlQ7aJ4l4qu+QEG71e4ZlijdakMkkoX2MXoYWSAQH/HdwVg+qZdL4EVytBykr
2UxwlD+5hIso8elgX8OtReuwKSgUzowK3PjeFCLt1g4J7zx3Bb4dPGY6xJNK3NSIdih9OTKvosrI
UvIyDxVGzpG8ND2nHPpsHMheuvPPmtOhnWWNt8Qqt8WLpXh1vMPUKesT9Lcz9YjUZl/zskayuUOy
OiZJRLPtJveckPP6oCO09khBB0QkQp6PrXQHKnttuQgZbOtRf7QrhyrAIBdyxQvRD+R5sJT4U23e
OcmuCvHpr+i3asOO3Z5vCL2ycnQyzzTCNjV2lx8L0JUSZsDK/nnvSgw7VlTiEb5tDCu6XROs5V7k
0HVPLhbozGUd8v2T1mYn7zY7CrxWui6teKud8MvIda45iwze2DLwCYsDUU7m/X25eEguS0LxD8sr
80IumniGdx/Jp/zC48WbJdSjn2YJdzGWQ7dQEBtYtSNj5whrMeARkPLKLINUGswTnOE99XGzr3jy
DWN8p0jIYPNoH/WE8iDM21qvoT5pUfSy3FQpWA80aaFTvSXq3ZP0xkxNWUQla1Ap0eQFAfdv+XOv
hEeSfxte53OB3MOV1x6YZJTSWrCuYbqrvVD8+EH1gmumpWFyfMuWEUfqxtB7/LN+H3cTvFqHNEch
iWF6gwxz2rAWtI7ejImS+jPs4Lk6RfAw3fURRPRkP1nAgyvhUZg3vzRPYUMyWmPs3mq8CdJbFIHD
FkalIZNCaMaaCl0wsVb69R7uwCYFZ9to6OYWsfPSo0m5ezYzSZVraks0ng3DDlK3aXyd/dI3xik4
4CzESBeVgX0x9czZEtyc/ZiX4DfVVn7uoFZlnIBJUaiAbd/EXWeGanXem976l2fRvrrWmpc5IhFZ
TCuy/WuwfDdyQNp8NCOfd4UiRXC1HOG1l3blr1FyCgPxr68+rkI5y/BRh5lDF+F7UPTUDxv2qUHH
8IgVRFBgu+SHLxJNmLAwFUqpzmv8vHoS4Q0CzsUiQh0vC3f3/L7CRTjXZZD//QRlsSfleY/VSS+/
i3OB83skYHPQNsUxisHwhOPPkEtaXHrTl48vav9Au4Nr4FXgOR5wrtYUeric06z/ZtZfirMhR1Ms
CFkUPo8SoUCzsrU1HunnBQ1OcSL+bj5jfOvVpNeXEL5SXOv4JMpHjfjLrcV5o7cDk8qfFinRS9+J
Oa50Lha/biCQ6E94XtxxL62Ug9+VYbVjrFjMxymmpEE1/9hMXP7vXmUAsm87+w0JoaH7uUVeYcSX
9I+e0e/26Jrh19jnKY8pARsjPqOQxa5W5UfkkG5nxdnUa01UG9nnh+nxnpJ7Iuj7y8IKj6lRmKcp
oQ9mj5cLFJODavEIqOyUYNk74LJ9+n9AXm9V20Jy9a+TMRj7j14dYDHHxUDSfhW0JDCjbtF6+W7c
qoKyh5qYMjJ5hGRZdO/tVU5vEiv2w4mVg2H6Xmn5YQhANChShR+R9JHYx2VbO2p8mbH57BJO6dS5
+q7rxaN3CLLIOwJXm5ZbkNQ05MlsdSc1qZ+mAf60S+ECqyR0j8cMoUmTbYtVw4s9YhAwFxW/Djw0
jZa9vLbjepIDv0e3KQm4IK7RcWX2gsXXDyPjYh5fLaIrkaktdJDKJ/xAlLL/idyL+1P7mRKzQqpw
EybZQ+smrMLizQ9gXii3zYOnngU8x1aRp+LDwymq75v5fqHyDVO+tGs8moBTvzXPQR6ld4oJPONp
yi7f9jrs4shWmAxU7qOyYRmQDrLxhSi38O1GyIzdPNHPDyi3BtQIy3mtsQg+YqOW3dVI6svWckwh
/IyWFNgV3kOKKhRSqzCHBojBuc7MP11VxWjeDOFqmoY3zIiVMkiQ37kEagLulmQYJpJXOQTGW0Mb
gtWIqBRX6wL3QXCnh/R1FkSvwGsppubmCjauctXTObnTyqrvgsnVTGmVFz4H0UaIYuCR16TF1ijY
j6CR6i+w3FxAg8sEgmPm9AxMKrkoYDIBZhi4u7YEiEAWHw/J3NlylW8X0sUDB38bIn7VMlqAOdqb
dlJT4meAlB+naRMWoMXtD8+j1e+UbQ9etmGkwkb2O2JLAg4r7zG4UBdsWQauq6CUBxDmG90S2UDa
ey7zzsm0I5QlaPptgR+R01To5EZgw0CLDTcccZF6WMSmEpLMUp/xVZSxQEpR5ZIUhLIfICceXXHD
khJKWJonuqkeMyX4ZHvlmK+ZwHWjJuKEy1cijfjRhZtqK59DTdTYmDsLM6qVQHgwyft8cnmV+AXT
HtScdkYx5nWqRq6ONv+fYhKaWIWcmk1D/32kDn/xqgLCTd8pFqKb75M8T8aDlxh42Vqr+gJ+8uy2
4ZuLB4WgYMPkued2aJktHH30fPV9nvnyh8BH/j++YQqWrhhxydI1qMihbTfSMyA1jtrvUtLhAXtM
snMI+Yd4yz6Q8nA1G3NoWUjnVbwJkLZxP5WPkdYCnnY5HWBJxJ5hQFSI22sCkGpnnLhgc63Lr1qi
73Boo70FNSSYPndhGOoHYIKOS6S9Vajzb19Yyy+6pGnxKJUIwXPcCN8W98yplnFDF1+skhddqWYS
cjSZ8WnKENhEaEm8rrCEV7XHTmMHiPSLVSkQdBfKR7XQvJeELpaGyMbxSLNBAPALCpURQZ4EbLL0
KjCd0Xx3O1vrx6bQ+PX7L9Y9SyXrNH9gLXmXsu+K8sLB7SdCMKzh/3LgBcDgncVFQj927l0QUspU
Vr4yUjvFmCCN6jDhs7xjOWl7W6MgJ9+xIDFYs4zbKqmgKhcOCI12MxsIS6r/jnVOKy8y7JS1vhE9
EmUnS9sIe6v4O3lX5zj1b4m1qcvMwVlm/TZnw1Zwfz1cnmvkBJnBlr3k6yr4+BbDoRvRX7vIrDvK
YLofBcC53XugjM2SoJ1nkyNKVV3hVXcMMUV+dBRAMUCj9fUlMCFXPZT4eaxAlAzg66zjAdzR1qUB
Pxv9kSFGXo3TiD65qGbEEtTCY1v8Ghq54zcZDbuQxqiAquNHoVoHtQs02Sv2DGwGhpeWqpTDRs1+
FE6J9Sy66r5/tlBqHDft+awMp1WoXW4APEI//B8JKmfDoutojirzUa6qeVZHb4A2zmCMrARRQAMq
08Bx337IB7I7hIRxgj1Cr+8P+I/rN3r9mEBuPU/sM80ow9DgjmSnK/aJTGlABsoW4Q7kfjOPrKIp
HM7hBSY23IfJchnf/5u7TAtbi79UdjpnMiAuR9MbbWezG7A1ZSX4h7ueN4ijc7N1zcsqza4uz240
wbKsq+Ju+3TGfmPXcuDkZ2zWLxXTv7D0EWzlUsK9Qjur2M7xkBBmZQHQ/AOTP/rR10K1f8Wber9q
1auHwXoe4GFvA9yhqtsXN3RIBREjmU0eD4pn3WtuB38K1fSajzWeHt1bw1v7WJ6rwRAcJuzEhpcK
T4tV3U75PpM5VI6dcqT1hkDKVRCY0PbO6j60ep0y0qzcZBmd8SEPJsG4qyYOeMgLcvIyokDl8OSZ
r9N+mEswHz3/aQv0YW02k8f+f/G6km+ukI3gJNGF+4JlUcS1c8SFgIf38cX11Sb2wpyGP0LPPzKc
MlA4Do7P0gtdzV2lpmQn7KzNEswyxmI+BTKGyc/6tmSK6av7G7Qywat3xWXBeLb5WDVJa8eTYvyM
ooH99UeaDnugpIPjtXTh2fafKfNKeGL+ykS/8c0/yl6UaZVLDi0XZgCjTNYY3F0YvgtxsEvXDabl
uHa3DjvJzgsEs+MO7TBJMpbL94Oa1UlCCrqY1IXMrwLkl5jQvoY9waw5mLza19AZX1OIZhJbQWOv
GftAk6oaPT8CYZndS+XapWMjr2J69Fd0ENU3yrHjCM2DfBABhXbdMoz8TK1bGQ9VI/QfNY10Fn1P
XlH3KLzeqYGuTjIsZWVWSmxlWtykb710YKQWV6REWSDdV+y+PoQLq5Mjtw4ZxrmR6xvUK37ChOQ2
vIXF0AlYXW0q3jUpVDQP3IJd/55D4ZKQuYYFTJvPJ1hoZ3Gwlp7e25Q31YlREZ/6Q916tT+rB2Cb
ASWieUlMHUhti3I14pvq3KVDYn3OOY1q2GQUlzqr28ALRMltpOdg4WMRvfyc1fDyF1ZO4fk2eKJ8
GhR/7JJW53tjov7ZbuQaVJyNxCPdezCVic175Aur3iNqWRlh0ejKUf49xn4iRP+HCuS9aJCsUMcP
JFfJOoaGOeYmjy3l3pfb67FdZPr3Du7Y5YOCo0AHEjb1SD9h+zhF8KqafLgSmQ5JpZWr2ptLjzIu
A7Txs/u5Pb83oRXnGKJyOLcDM4fzhK1KYymscT30bN9D4sC+CAs7TJ7LmEzTUNgB+GZEXUtmQisj
r0+zpFZ87+G9W5whSGvgq85n6O6o4daf2fPeVJBklaIfFD7o+ECkG52sogCekwxKaNyhamj9S5Zt
+8l1/6cRmrqWvihpbd5ISnuleFCVqP8dcGuAFXeOSEtKi7EkFX140HF2Q1mrtyeJz3cts61HapUp
lf7qz/flkMEUCrH45WdLiJV8Ie6Mo7SGt4xiu+9/kAMksLhZ/0W+PhSZEuc3vqgsco22wQErYGaj
lTxNhP9OmH3egtaQaj2gvceISQlcQgpACZbO6acR53N1xer48HLpyzH4MyhKzs73zynZ6h9bHrB5
/vbtSh/LdE4Z67ZhEflVjBo/ObxEFpaIUsFnwT5cPVh/E3EpPkF4YTbVJa513XzbJAWBhYMpkh+N
J9JlZxZnn8ioygYiw4S7Pr24+mHNAKKBZAkRhdybUPJMxJtP4wLNy4n2aADqgc00TpNo8UOxo8ef
Bpcvlc1mm2HQuw/qX+YfWNH1OQcR0kU/P+ObLfDhkav7vsjycYp1udNGbHdy/1FZNlBhigT42pAn
up3x+9GxLiN4iwRNPCrpn03IkTZo7lZB61fPNAj2TOoAs2NU1VOc3OddoKeAPMFAkO0qYhVkY8K4
tc8mdBWEGwz/tOl1ejLaWNWyPfNqyWijAs1vnJLpdxUCEziPHNj1rNrqn1Mt/sc30ZGgj9Ziw9fW
uPihLf1qvrwR3t29h6bfKOOsI5H3NQAvtPHDPrqdlM9TUdRB5Wo+JeurVLx5dngl8cqpj69urE2+
ViF0NbKjMsWQsnlZjwx1yC5rkTuw+RNBjM3qtpFR3TjKbwj8gv96uisjhnGNJZYEEHKhOZl3p/bY
YuoQf5i5eFxzFWyCI4VM06kT+D4sBMzXWI5ne8Qx6Zo85cW9+gubFHgfeSV+cxPITQHXe9OEeyj2
RQTWpEJqIU0+fxaYdFfeDVbnzWhRbZj9C2c1Ng8d7fbxLZmuVnUxq8IkpWu+AGYK5nfblyZU+IhJ
QtoQ/oZ6H88cgd1e0ZA5Es/dlUfiPmkT7fM0KSGQawqaZrLqUCUeIXYwxjBavHr9nLS1/cYvt3LY
rRNlw1PBh/SBUGlW8xxz+ABHkMq49KzPCrmeQQbkfXlfJtq0c2qBTpFDvMBl0Ma/QeEh7K5cDj7M
UXId2CchF9NGZY1BTfVW87LiRzjQhOlpvm0v4qw3mWJ0STxt+/j7gsWqYLIqsx3GPHwKOSU+DfMO
yUo9gbvHS4CFC686HU83H7fG5X2iXTuxe7iFgo7RNQGzMenpbXrp7gPtAqAD+w75Za6cOrOd8sZ2
ffKBI1Kj/ams9cItz2MO3BJ1YcidUmPPsIzGecW21W+KEeeZ/R0TWvhV6uc43En3fdi30skwz7xt
vDgjt/a2hd8AwolGWvGzxTWIZNlwtBGi4QVnCTzlFqY8IWl0P9rjdF4hkiCJIyPi8pb2mTPjIWC3
mv5rwn7x8U2Gls5G7yK1LKaftKPzsAc46en8nuiAxQ6Z/NbgaAqdEqvm6soWFWDCE94t+XFDULHh
3XNe8U14JZKbYkqio6MnFzZl9xz+aFMKh63x8YgEOlNEdGgQI3ketQrtbG8XAYjCvi0571DiCcfC
JJcSBqCQIz0M3Ujyut+a+53SL5kvdN1GzSMLaUVUi7GQy7rVbHDXYdJPpxcU3TiUqtLOwLApuqfq
po9fpN9HzE/90THgVGPN883jxUQDvhmoTVt+B2aCv5/U/BpI3Mkee4iVsFkGWNPgKfQqxFnGBXdn
/ZPPmHIAZpujKQtymqO43C7DH7kTcYyXlOyvNjS9fz4cZzbtKUwrvukbt4/I2k1zubDP880q1IUq
pSC80kVqbX2Rm/ZOMZwTaN7ZN1/5P5lXUTdAskCEzvR0UZ5uKBZj4sp8mwIwGGMwbZqGBC8q40BP
3v57Mnb7ZKB0Bf0Ti6awoR1pG9jYxLgg4njcjP1q6gqE6YtJeMzcSb9vWGUxTIRnOF7xNqx3wb+W
n/kYfc7dMH1weig8lc+hi6HNYycgaNDTD4T0SkQgXXrGfhgutg4j6PdqONTdUk6iAxv4Q8ZefDZM
MCAjWd1CQrKyfpwHQ+c1dB5Pid08smD0IMe9r9Bt8Qix0MI4a0bWMX5SZCoOakpVj9QvwichQPsR
+ZsPssNi3ZILkXABmru833QEqU3ofdao5E3AzRZA1u0kUJrWx/GDDaKct6sThIfSFjt+VYp/3kz7
3boh2Fi9IpwA714OwA4MwgF5mvs+9+XNB+I73niTGg4eZ0Twh5HYH8aAi0op4+MV35G2PLgqP9x6
3WQDhD509iCCUDd/oFJ98sUHzAwLQ5Njopfv7J2Bjif9OGxHXotr2VCMmypwvWovBzZJP72lVk/W
evWK+ZLd9tIMRI58pFX5habAiWKdrIhA6D8l1V/rvrqCqP+31hTXASf1BMB7VwHDC2eyT6c96zet
dt1X3Re3nS9OK8cfAkhoxCBCA5O/kAatfNfdmBz9TfAY8iSwO0cEQ6eilCweKxSkAtI7UC/73H3d
245tyKCDLlDEdZaw+Dsk1k/XGN7HV0LNUEKGIVtagC8qPtSmuFvvWNBwy+Sg4x5eBB2z7bd8RqdV
sN2qEBChsQm6JmoL5AEqx/wQ5yQ4hQJejhB06UzSPq2nF9x5sRFYx9JtOk0lUSd8k2l9nz8T31CJ
K7+pCnEv0vNmpF/uphTxJUotoggGVOeGq7nTdV2lpe0yTsLWS5H8oXx7fmTgnSR944J4z6gkVSgk
RmRfCbJwcf9tbbjQJmphIdJa+xGSAHkVntwETpN8hFd/FLizXm31vstjig33+CRyfsi69mZ3SAJ5
WXca6mR7i1jv6jByrQP0eYaEW+ZxrVUVFubLCHws4gcbPV8OKoLTML0fUMDDuHUEGoJ+a2O/zz6I
3EBOq8I18uWoZjixqhWSNQn4LMQ5bA1S17KF+GY1n2d71ZhrgPb3S8Vd7DtLHRlV4Tq5kU3UZ9xQ
jdh5h3eDiyurdJ4xFSLxZ975l9PmN+KL4oSyr94LeNWy+5r8gcqo1SStcP1lVXQeYh8cz50fUIq7
M5EK4/Svt/Us/FG5w/TaWqgO+P5NsfGhXba1jdZRrjGY5gH0b25RGk7hp0wGuFF3QZYx/LNxdwyz
OlMqBjl1+3iilWu1ahNcmKU0LF5EjKbo67IVemMTz7xPtnZSR+6lLDp3+gfmSnC+/Ov0dTkczSOZ
cCN2TzT0i54HZ0I7sCcw4VbaNXEmL4RVYpxi7NyDRdvTeoVxrzsVNHA+DmnMr/YFhSIEL2AEZ7bK
TE7MRIUmeKQT01aHtDqs68fUZMa1n8tDf/xwC8eLwEC0XeV2LGd3zPlhwiS/FPsapeAtjmw3o7dX
F1av5/f6I8syon2eDX4/qK9sKBQpcdaoa0dYUVcJcMKyzqH8zWVrDAdPDmr6B8Nms6gfCAFnWT9F
MwrqqbcMNtRxqqp2uQSgwQnhBJuG
`protect end_protected
