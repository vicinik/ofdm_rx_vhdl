��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��8&����3xp+���7�����`Yb�H������դ!��B��?ܦ)[� �2�x��*8�i��ZOr�$D��c&x���
D��X�jOn�!_�j�=�&��{#Y�'��ԆB�7���������M8;4�J��>���̓� ʟ�,܈��ڼ	4������R�[�-�Js�OOk8����BT�|w#�3!��1;�M�#s�4:'#O��D\L]����W{{�'D�.-&X�n���
L�5�]!�v��-a��CF�@L3�8"�Bg�$~���������y9~���� �Ԗ�ON��u���B��IdZ)#v��?��.Lx�W��h^�Dp2[Y���}1]V��|������06$��?�X��B�/�߀ynyAzf>ƻ���u1a�.hr��o�ks�IK��D�o�r���q�� ��t~<��f�)g���I�S������I�te���"����y�F�P���1D�*A�o�E�"�E���TN�\�-�M�w��msX����9&����/�sr_3��Ȼ��Ot7���?��s��Ne	����!�P���Lƽ�E�F��}�gʄ}W3gJ:�������3o��*]�Ƶ��m�:,���m2N����e��} �@���Z�*��©��zpD`��j�B�"�Qe�ܢ]�9,Vw��h��1�ߴ�'3K_S�&r]�s��'fEm;H��%�23���q7�p�[Cn���e���Y�^���E,R�g"@�k���kZ6���a�.�I�q=�q�����h�ץL�_3$�H8�ͽ�t�(���>��e��L�N����$滈��V�#�5�|�9�-c��+�`$Y�~��[թ���C,�W ��+M<��rٖqW搟����"�� ]�o�r�DQ��th� ؀ϼgm39E��w�@0�R�bH�),��40����ŷT��:6�bg�q/����&M�c ���f�j*o��]T��װ���Ö������8V�ޯ1��ꓲ��p�#V��s�=qil7��,x�.@�h�Ǎ[���a*�&A��
i��F��w�xJ��a\������	�1�g��a&fb��A�FAHJW=X��gۿZ>{m�p0�/ ���!"Q�?��D��Ӷ���B4��f�o��Uԏ3�Z���e��(�4�����:���&p�8eLbSqq�˗�!c'�4���z©(/�U�O�K��xG�W8%�=E�|���5 ���<(p�,�k��י�ݑ�3�˶1�����vt��fJ�v�|�[O�E��⪻#s��i殲��6�<��%��A'��We�=p7��	0c�xg�㊹�w��2<�^�~#�a�h�h( Jc{Y�=���G:Ӷt�����m	�oI3�t�CPO�xOt�,}"�T�>"ቿ�N�A{c���2x#��a�}j�ul'��~�e��ٱ{��s�O��T�C!g��L���f��8�sR���D��!�ˁ�|M����
�W�꾰�IM�WVH��%L��#?K~@1Isy�{O��_��Z��{���H�|[$�{#�y�FJ��bn��$Xz���J�RFJݡ�}2����u�]�߉�(=աhG�q�z����-���������4;�y�%GTEy��Z]J+Np�_����,�0^�u�k=��FD�(����#K|�K�������`Z�����t�{�����	���`����h�b��Y�!���"����A.jH}S�(��idɓDӓ�"ơ@x�Z���5Z��z�N�,�.v���c�o�-�f�Vܴ��R�z+��x5#��C��A�+7}��%������p��Hl��\�Je�l���!/)��=�������z}GJ����	��4$�����ݺ�@�e�rj;˙�j�FW}��ضM�~)�aC����X9�mU[@�'0u�� o����s%�]Ј�#�J~}$���jf�#���n�J�My��7w�j��P`@5*�3{ڊ%jG!�ШQ������fS@�3�O�:M��$���ڧ8mc���x9G�L�@�ii҃���ci{���q�3*s � ��S�bKɢ{�?� �`��u���@�8{�U.���ﴚj�Z���x�����d��@�E=�s�*�l��Ѻ�q�Ԣ
|�K������E!U[XM��[�ōu}���Y��{�Xbv7x4���>]W|��Y�Wv9i���>ձ�����}����J�����*��.��[���|)%&n	���w�5���3�ψ�k$D÷�H�%�araG+�fL��n�ʵq��D���Z�㖤����K�Z����@��Xnb]�}�C���e/�iH+��z�bA�킽D/@_C�u��;W��S�;/x�/�*���h�r]�K}-�̂���QF�z i�QInΑ�h/��D�u�˺ŘL)�A@Vu�@H��_���!|b=��V�D�9��4�#׷Ġ�����0;��Ymܝ.*J�NF��l��?��ߩ��<�p�~��=e��Wk��'����C� �I(cm��G%��yP�����H�9K��Fkm�gz6�O-�f��K��ޮ�%Hq(��$���\�@e��S�ܢ�Y�I8�b�������TVY<f2��!Y�%R?�@��5k��_���Eƫs���-�ρ'VL����g*�e�Q�J��<�����2)��B"aP��@���G�#�|T���T���o�U��1mh{�b�v�ߢ.W�����������6�/� {���%(=�T��%2Nޚ�ܲ�E��ڈ*��vv_9����S�6�H�@��/o�*���O�g�ʌ��{��
N���{�h���D�ˣ	S��N]u)�&D���dF���"�x�9�N�A�T��i�ڞp�nP���Ө<<��TOd�4�˒�:#����P|��8)���8��N�ګq���~ٞ��'`�/z�� .O�/�)x���+�r;Q�����(���n�Z=���X��Ɲ0�H�\k0�����8��CA��h��+��c?:p��w��3���!�tP��]�-t�Sg��l������5����z�c����5��y����	#}UfoUj,gߙ�1ʻ5����z�l� ��� QbU)�t���4��wo3�l8��!��-�_kǽ��|U�~Er�TZ�%�*���p�i��A���TO��/�����M��N]�k�]�գ�R!wŮP��Ld)���Ã@:�~Pe�I���+_s���۪D�����ю��Bп@dfT����J�����I�%��-?��q��)��^�~5BH��������T��[�e���x�/�n�b7.2�Iz�#mw�D2��]�*�Y�j&{�z�P`�4{��I��L�(�c��q8-�7k��h
a�@�m�G���/uN-i�-���^k�L�ǌt7y'V�z��ڟ+c!�#�C���N%�t��kV�!�=���� �:+Cd��ŕV[R!���]s꣠��֏B�6�"�^�s��0諰1�ew<O9#�$u�LJ+��ehR�^�w��oJ���m�|K0β����w��޿���1�}�1���F��2|2֮В��2�9�l�Q>�`��mg�oĆ�nS	lZ�O��Da6��K�t�rq3����p��v�~�h�ݙ�z]ɒ�r|B�c�nj#O�!��.kMPS��V�af�����?ՂA��"m��e&��uTC�`��g�ֶ-��s;!���T�0ۄss�s�����Eݘσu�����l�<7c�S���/31'y��@�Ťg^Y��9��P@�A/wݭ֪p�~��r��A�Ǟ�RK��0����@-�$M���c�M^|`Jc`U�~�+�o=��C�k�õ�`�"�>e�u;����7ZT>��V��Mx.hfm��.}�C8�2l��:�.%G�� ����VP��O �PUr'O� �+�
h���g�ׂ�.q���h`~Ppz�رy�g\a�vkS�1��M��пE�%�n�>)oЅo3��"��*%t S�c���ܙ?;�i�Җ���\&H+O �9�0>m�L�5���2��%����:G&�e����euk�!����":�=)8z�Ě=��q-��:��O�� cX(���t�|�$GQ�����oJ̮�c	�vu<FR��:�B�:�:������)�i�d�!�T�JE+qiD���a��7(��/^�ϴZ�˞��?�B2Э�I�䷞���h��6��y��#	~��c=9F�Uvkj1��^
FL#o�G����}�o�L�)~E���V�DV���!G��<���� P�1����lyA��b~4;p�ksaA׏�9d��ѽ�ڂ�X�]v\;�/�.���֕�|��@=��?�ޠd����(�.ϻ���2G���4�ADm��ܒ[����M{ؾP#G�;�9r Z?�>��8ޢ����c��v(�ܑ$H��Tuq켣 �ɨ�y��UK�b�֍�Z���d��^-���r��N�x*��Ҵ'�����]�Us���ﷄF�����"�����,�haJ��t� 9���W"+|>C�~Ҽ����<=��c&]m�H1�&XC���������ku�m�f�b�j��8 ��J�(�}���ɝ����#�)#x��_	+�v��}��ӓO�e�GU����
�"W�\�F9KH�(�J�����c�����*�O�ʋ������o�2ȃ��B?f'���1z�͒�ٌ:����R�y[-��q1(��v��("b,G��T�v�?g�3�Z�s�2����q��N�R��ઢ�A�Dd�S�X�! ��� L�8N�:[d��H E/�:Y~/��d	T8��u�s�G��M��̔U*{̳�۹�I-=xܷ��UAM���s�%"�T�a�л��t�n�[��>�s'�ϐ���;.2Mc�X�Fр<�܂�M��9J��E�O�H��~nOB��9$k��5�	��,,75:7��5���!�����D9������
-��qڴ�!����V��	
H�c��o�fC�[�o&�qE�HYx�背���C�&Ca�s��?�Yr�*.��Xpx�
���A��(�H����ĭ�T�i��n�i}�(U��g5ɶ��ԽQ!���o�A;"�>��d��aV�r��a"�@kXnY䯃Uh�
ˆ��O���/$���6��q��س��6��~L,Z�>8#�Zgt���]�5~:�^�w�
R��e�v�	�HxO �&MD#�t}�$-���U+=���@8��F�i���j
�Jf5�>��q؀L��T��B��Ds�}9ߠSN����
�����ψO�nc��92�sX�!֨k��_�m����i����%;s<xϾ� l2�U�W��u<^B�R���]O���(r`Y��� �ھ��1�o��N8'��8���_J�{�f"���	� ^2{㥐kY5�,�%��c'a;9�,�Hp��	���u2�%�|Qɉ��kLz��sZ�G���� $�Ov��J\(��"4@�[P�7�8��%�G
�q��7�+���
(��<�Ƌ�k�Y1�OEI��N#W��%����F���_�" 5��WzZ���f���Ey���G|˃���HOP�'bs17T*�ȋI8� �G;hh�AFn�?I��};|��<�gX_�� �\oT�,�c9��<��K3yd�HS/'}rA�o ��Sq"�S��ɻĚ#��Z����h$�bo�[�'�M�U
N��S��N.K���-Ў�K*o���~yIܮ�
��ʂ���6���p��ag%�,�䄽�Y,w���U�b����o��ɡ��5��f�_G�{��=Z�5�=5L����f�� �h�:�6 	G���=i�/~/~;�8O:��q㖇����l������J_(��&�J^~3�R�?��<7D�œ������<��rF��'Jt�6yR�n!����2�Ű�G�F�z/(�C�-_:U潛Y��j��2ݖe���O2�彩o������2XQ(k�c�^t�%��Q�4��3a������zFe.x>� @G%���g��ϮT���"���T���~�%�<Ѱ�s��7f�,�}�K	�cT��Eb;�WJbu�N��2�}��>�V�d����{Ӷ�#�3��;����-����/<������� fU9O���ݳ4T�0@
��1�U���R��A�_>ڍ�(�S�Qo�h���wmf�Mj�.�"���g�k�2�ӫ?�A�x`�:�����ߎc94D��9�l�N�K�{����JB����K��!���z$jDq��(�p�&��%�.w%뿕���y�f�:G�d���{�jT9i;��\���Yi�H�I�9��`�{m2(�Ւ��DҜ�m��9a��%kݒs���H�v֘�2~V�'�WaE���މ�+nǌH�D�Ǟ�k�&�_��꼗�Ho��GI�\��O�0�C7�{!����g��tu;�-�e�$�
�W[9S����<���v����;J�'�pB�|�,�-QHI�{/�7r��U	��E��|��e��B^ܚ9����z�ߺ[����E�t�m�z���b3G��T��Ij�yTtӏ�paTu�d�5G�7��W�m,V�qr��S��*7+�ÖL�+S	�12r�Z#��0l�JZD̄&��a7K��a,�'�g�A���^�+|�l�R,w[�9�>��Ifb33���
G�FnB��D-�����KԚ��pֽ��Bϛ����x��0�����Rh9{>D;"B��x|[�~�NKf�S��}�M��H�'�E�X9������-3��y�p�(�uFw愔��}���:�e���p��(�d�O{S��jg��U-i1HRܾc{��X�
�/7[b/�"ac0�t�\����|���H	��dJ2���P��v3��S�J�^inK��KF����4%d���:�VI+oil�:L5��j��S�PvsPK�;��\�E���e���:�b3eY$}�;�D�矉�W!5�W���>� ���߬�`�e���y�#�y���+�I� y*~p�Z<U!���/]'��&��~�'ݕ2����]{+1�D2�uؿ������dy�Wץ1��a`��b�3[�O�z�3�>��|f��Y;�󬹈��&�]��nU�͵�U���VSx���<O ׎���Ԭ���sz�Fo�L��/y)���݌17v�/�1��~���4`ou\�8�u��P�2��9�yw�2�j�Oޝq�|N���� 1��l�m���H��ğ�*�g��@����P>A7��Α���S?3�=�p�{Q��R�u��&�&R��4c��J��\>�3�2d,7���}M��7F�����U��aA6K���e�(5�[�+ym��W��턱o�#�]�VU�SI�I�	����c�ѫ��,��O�MQd�1\T�O8t� ]���w,�`������Hc��!f�J�i���(MJ^u=�Ƶ�@'�&p��4����PS��d+;S{袋'pk9V���7�z�e��kR��%��W�D�!/�~Y�zB� 2/�!}П����7�*S�_��j�j1��t�x��┑Xa&Aҕ�Td&
0Y�.b���a�KM������,�I��$#j8��)>��W2�(�����ǟo]J�ܩ��D��� �l�`�>�j,_� ܠT�L����~�	.�*5|�C�~�+�j.�F��(�)�_��Ȗ�Cz�H��g�W �8v�%�N����fn!��-��Q��0��7-�<�B����z��%� ߐ`��?�N��"�Q�]J�� ��8� ��zo��+�M��{���Z�9�IU���V&E�LB�}��Tq H�dL�^�:i(ٔ����rwN��TJ=xeQ�hSrܮv�A�J,ly����*�R�[{�[��m8\zvWv�|�N��Q�M������?�T {/J҅ƹ�j�8 %ĳ�p��3�7i�|q�+ÁY�+;o��V���B�ա�&�1�#�㙶!�c [;ʭ &���Ƭ̢��<��m�-V�ZRIL�֠흅#��Om�?;�{[��Ï�]��*��؍� ���<�jcB5�G�],gw�;O!-=�E^|:�7��ŋ����+1]>���8��[������͐ؑ�����*�VͼQ`�y�%
Y���ҳP�/�n�q�8.�gܡ��J��X)t1\�0Gl���ml��z��uAq�Hp)u�e�E���|���` �Ԯ�e`�P��"9�3���I��x�ʂ�C�:�h|Ӟ9��~kdI�IU߆i������Q�Rva'o^	K��u��m��I�K~�AW�d �[�����E~p��3�FarG�z�s'�n�"��|��}L��I�i���63�IX�j	9S/v�Ym��r2״�&S��X��O����O~H�ɿ	������Z*�3y
��)J��4d��G���؊�_hi�A�vk[_J2�G��.[;+��H��x=��p�Y_����e˛��L�8-�5	��*g8Cψ�F�O
ń�e���bm�5S���	u3��q+r���X��%�vX2mBQj�eh�}����39V!A�WS�s�(\8X�!��C��=��]w1����J�0'�(��Rl�J3"��������ǓR����E,���"���$�c��O�ઑ8R��3�q��ZrE<x��;6�*�G��;-SN��d!����J�7A������2�$�{���q���*
�	�
%8=��NX��~��c���{�"��\��WQ�9s�Ő1�	��=f��SuI���Qd�b�c���pf���
^�_�x#g�'��1f^I�����F�|c���Bo��<�`�F��<��<
�9�-mc�	*ΫD�B�+$��g0��tȽL�g��bW���.�B�tr���(_ܭs2SH:W]bi���ҏB�vM��7�"��9̷�X�&��^RP��ј�D�#���4Q���a*`��(Ӻ>~�YD w�'`BK�Xh}9�t.�!k���V`M2�p[J�;��|��VWS6W��]2ff{7"�a��jꆤǨ.\��wBȮ]D��Æݒ�$�.8#l)R�"Wo���입I;y(.�wxxjG�+��%�����Ц��a�Pvֱ ?���:�K�b���PY8�����]�@���c�d<���O(�Ǻ�,�h�#��L��gYXuc����9�L'Ń��M0�'���������JC�0?��㰂n@-�'�Ť����8W챓�h���r�B@'L����cw�g3��@&ď��sw�U�B�`t9�1����?��ݦ09qa�1ķ��@E��@(q�FU�u������7�$���7�Ώ���J�ǰ�rU���*���nZ��n��s(Ocn�!ve�Z!-`��v�`��0@�R��N���ue���HL����rC�֐��ǃ�*
4+l�|�iF>Qo'�	'��\��i���;��yՐ{{���L�|�C9I[���P��C�\�����a���[ݡ)�u�q�U���j9<�j���4�����|-�c��������Uf�9f�iQNf;���1�� MP���o�n��*b0^<��qy�a�)�E>��V�R�y?�n�"�uQ��=�ށ�0���@U߶a�	��"��iv����]ɿ��K{�W�fH][���ի�۝L�b��{-^��@���xd��'E��n1�܅�
 ���M�������4�
$\���9��>�7>=6�����*��Kon�ď�����7x)����5u�%c�J��7[?� �vzH"�iM.���8�`�Zu�;����t�G��Uw;M�|1 �Xk5[��a64��o���×>\=DC�M���.���=4����'�[���@�었�Y��CT3$�[A�"A�t3���}�9����7���]��)�J?��Kw�/x� ��@��]�P�B)����0����#�Y�8��/���O ���l��z���F�Ez��F�νVC���텈LL�=��|�4!��&ǅb�;��^DQOU4�9Fls���L��,�d�9s'�XI�0�.I�����}�T�5<0Oo�W�y�����m�b���1�_�^�A+�����Gu,��G�6f1R׶iґ�U)"x-��.ɖ��}��P�3���cI��ښ���+�����E������8�$��s�<P�8g��	�<%�,7��\B�v�L+��auȗ��������N������	���1-�
�Y[�Ri�O����%$)�X,]*�]���jc�eC�}�����]���|��K?{�������'��uMze������-����ȥ��IM:��#��l��i���`�$@b�a2�K��3�a�+%>�2��b��\W�r�+Kj�T.�4;.��]�3�F��E���2o3���h��/��*j��y��;y�X��L�K��r#�7�T(@;�=���XNÎGn�嶂�k
��~��- ���)����k���V��D�0<7q}1�.�d|,�*Lˌ�U��^f��od��y^��!�þ�V��H�j.1���̍�ŀ���Mt �����Bsi��7$��y�� ��a;��M�3�i鱆pAZf�/���=Y\����.'���� 95t$�>{AR���9�Y�[�0�sld�(�S�?�X}��X�衿��w�ll�q|���=N0#�#��M���)�| 삭��\�?�<U�(��a�������u��]�ͻ��q����#��_���\�~�|k�wyr�R	��%DO��`��L��zb�N �$�!��F?ܮ��d�v�,����.����R�W�Ev�#�^����@3����T3P�9�` ڶQ�:�ܒ1 �2 "7�aK����:�˔N/���/�M��tY]�ȫ�>S�ClEy��q�^s5)�{j+�Ma�M�}X�jl�y*