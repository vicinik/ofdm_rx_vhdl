-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aKU7b6FA9Ztg6LoevI6YGdYbV3rPAl59sw8p5UFG1IFCdNUip1w2GQJ+0FeFf5OUdcDmwSEXqxUq
DR/rcVcX9ecoH+JFuPTRGZqyhtMZ/D2XTAz2jE/+lDraFPxbtBsmdoHREa1KHU4OCfQozpMx+wlY
6ROrpXuad9ZL6NMaaK/mtIBELHajajFYO1GEDJyMRWDJp7+hwX4CKuoBmywh+Y18+/va9WH9DcpD
1VdJBUGp/T/gpPBtjGVZleXiF1j8rEsUXOtVGnxEHym4AUpESOo46VrcFcYrevrrgRkwfli8Uyfk
g1ufTwuptooFf/B8rwzry1Um/vpN6FdOOQcG6g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 100896)
`protect data_block
lzDS/cxnNhylzMy+vj7tczurdbVNk0cOg9kZ91DoTcyH1aXM2oSc2KYwDWqzUJ8UdY592JcfjaHS
QFirymlCQbfvQBeWHFdpAK1iYs48j3IWq+rZUvVMowyWcbgqJQWtO+abOgnWTL9Ca8t8kVFUF9D/
oAcdHF6UvzzooHTN9VVmoxY2CGWcAKtww/bfbjKhAfFHhrpzHQaaeEfHknXRl+KIDr5/WEsYeUba
DDCsAO0mmWE4FwsaE5unWInevIOHsmEtsu/lJlp1v+evPqaJqh9yQwt5gt381SUkr3HX3H3sY2Sj
2bbMHQVYFaSwSeSBk607z28v+z/8DmkckOZetXm8UqfDd4gCxNJRRTkcCdeSP+CuPL+RUvWqukMz
B4X20WPJvJl/WCIEY0U1LqRExMHDM5xKLMX6UXv17SMw79NZ+dhpnssE3Pu7Aqz/HFRQXO1iPtr4
hl3nCMPceiNCUBtvWUUPc8Y67p8q60AnZipUAgQGrYZtBoFYSqZXTwaEN3RMiH9YwfpFv8WLvWYt
MOsPA4LEy1+6LxlIkSdSo7BH0tZ7OMfHiu0aG7MRTET0iOfIqioNH26lzvvBMm09fZy9ATnXZBxD
CPark9B2SDYuKTz3GHARgdOraTwN8UREmTuw6s4Semql31GKZki422X524haKVLHUCwPMnE9jXpm
QerShn4+MaeBZDDJYQoFKv94cfinu8E8uyRh4OaHXleznPws5MFh1szkHz9S9LMp8qycDzHfq2g3
7v8VWxqwKPSSP0S2GZ0EPVJHdlKk7oksug/NyA8fx+t8Jn45tg3BuTr7koqiSd1rz2nFkAk5v3JY
AXmYyev4C/Yzy0MUoL+xG+gVbG1ly3H62M/BYxBb3shfZgxFJ2mSUd0bFysuXtNVg1xOFjvhUtXQ
YOnfm2+iiHATz3AMsR8VdVvd1NHtQZy1KxGJvq2BieLNygVbZ9LypApYxneRZnhG6AXOdfS+9FMU
HZ73gbWp6+KJ7LAhIEaS/2ObVCN6Io+xKjznvt6kR2ppdldNKTHiWoI0A+G2o9GQoBhefSlexvCm
5g8i6ZhAMTAo9e1xrq17Sv6gAHL17F+/3+NMDwEV4rCIA1Cz8GbVDJyGU8RkC/frBqCTXI6WK290
Hm1lVv1wCYGJRzPOP4y+vtRgPTO4rPhhHo7JCB6HpSuL+oXbbbEaV+c1XAiL6oVnueqUQzltIGby
IsIXNC1yFjgWyS1f1clfYd42oYRjnSzC5KhKarMOR6Vx65fVB/GYmwILzy2VJsjB6pEhEFt9aRLZ
u94ud4HsylVEQnCgLw7tTj3R7DVFlpuB4yCbG1r6XUfgmzC7/RwSj4mZFuc+tzfOgRljYh1jrTZz
f2okobKFLfy/0CprUHAh/PS60xule7yDwoxABSedSafthae3qRWSU9y/uBdqYNcOhh59xzw3FLPd
Qdly88gKZS5edvEGILVDAga2UIge+WMpQsS8PombjYxUqgYsID0CDcs2xVxdB47YXUD/A0N3VP8s
HbMq61wahk4SybaKLiqbYXfdBDgX/saeGJZFGxXB6WSwjXC6l1BSrRB+6yKAo5BFY4YtWuwoC6ZV
ezaFwqRha/awDxwrfr2AIx5L69p4ZrWbRklYjF3dga/9MenG0HpVOv0Xjq1q1g81MdoKslWBqnoV
rohobKxnIH982ePM3aq5kNfnjAwGhdv8SJ11m/xvIL8xAt+/UnoA+AyZf8QfegA6s88BoIAnS0D9
aBXCpWW3NGUr6dXUHbHoebenOAGwhcP8qWwnCXm+d1IV0biae37LZwKgseLYYyPoSnMPkhRSMe2m
WDtnlhrgzQ1K+fMH1DYpcmqZjIxrcEiblA6ItbwyUScLdknZq+OrXiB3pGZS8k7dEhDr4fbp1M+C
O4EpKXfZxNAhnIPoFokujLx24ZBznkGUBq/nB9Hv6F/5qxHUxrXFqxz1UAQ7MS00w+8S35IoaCPs
6K6vckTh/5aIPU0QLQUeZRe3bo0FA7WEbgatkGXp1jMKMhIBJyQHq9aKe6wAQqYr/EFpb0lA5Y/f
ABlfD6PnqMHsq4in7VNxY0K2AItCSg9JcnTl1q+zzwclv1osduHvp4geolUDSb4RwCzTIEHrgJFL
BMFSazDm8Sf15t3YNlU5tHaSxULT5F0fSnLKVPE3ZOWoFC4XpAmYMEZCn34MiZjs8hsdepGODLt/
cCTC20+Xn3yuRo7Xzu7VYVbS2UO2Cn8wU2C/+lRXVLKtPXkpxoSDfH/vkLm/J6LW3fFVbySrG1MJ
qQc+ER+qnxpqyRV6nOZ9+9J5fD/Lkx1bwceNaXBYYBg3I23/ZdskgNnWxuBdbh1PUW27k35TxJwL
dn4y+SBO7zl8xYkR83t5YfpWjlJhejWahGcbTo1NsIeXq8QkPr09YyE6mUde5POztlv6TW5UsWFN
g+oGcTDemo3HsJ/IDCkVL9U68yLszmlGBiXELbOnZyk89Njx1qUrbq0EojwOjLtMzZNZmUjjpZSj
H7rRmzP1ytaO6DhB9wbyvcEIzyRRqfkYCv9PVFYLUKflcvgIikSZzKQK7I3gPiNewrGXJ+5OwSGm
DjnI9jcT3K3rp082nXfPp04bqaUz0Zm78tYHFNJtr0cZ107o9GrbVmhd7x8WsfaNtYhOS/6i7eW8
HkQtA8y++wjJrujpLFLLQ6VbOhh09mbMYIHqJj6h6vy5YMvSsbbQp0U0VLoMioDsaV4t7KJHtdde
wUoQsc5mBxE2/TFVI0p0xagLoII7xbZi6phw6JFlaYUHwIMSAqohuylSU52TPUUVyPF70QHi81vj
RsyYliIAmf75BOkOnffhKC9PCJD2zWM3nRlIraYhYHQCIcxAC6ZZJRDM4e/i0Pd0eckYfmDWr9zr
sZeqBZfulsTBTU7nGMXtI9LulRmMP/mIUSQ+YS1Xe28qOPH30EY/BNNo6K4Knl9DhzrZ0guW6IvR
LM4ARnwtBY8zi3NMlE0S7MQt5oveLYZt6FhV2FF05nmdFVNRe+N/bdXgKeyxVX7Fpx5+g332zM7x
r6dl2CJRPOlP5VQo08QRQHkcZt/NYz4tCCw7hBTohuO2ekMnDHjSy8yywmriBJg9WI/+ZRg7esD5
S+JFko4SZte8taKwzKqxIJDdbmrXA4OEF2JkrtObW0Qsyprwr1VulGILRDiw1om9ho+QMYq3SbcE
65erHKYEPgj1P/i6cil0MweeOD55QQKVbtGiUxCpH+NbNwLm57fGn/5FwRCZvdrrifINjC8U1kNU
KN/3I0QIutHHKFI5ToXjuGc+R1t+TEdXHjmHc5ERPeQ/F6vzNpIMlSlfMZCNikSj9sw6bGgTA9+y
ioSarDCkdGhZH3TsNE4yiKAOWrbhCyi47VUcy9mCly9a8A+AP0bxGgVr+WqfPeojyvKdhUH5RTE1
VkEKSqhjIyWiaHsVUiEvLdNSbclKM3C9wasWXncet0DFS7w+Co0nXWlqbAMehp43mukm8U6jezk/
rUNT2XTDMl/XaTCXHFLL+rTiED10NElnJpynV0w0APe3yhDdyiexvEBpFaToDQ+WCjBqevWeyRJw
Aq0XZNR9bYgpaE8an57IOp+6l1XoZk0Tw8n6YcaOfd5YOhQ2Wj/swcmsa9InBCuw2fhkjZZ1fV4+
DfMH3ajxHP3weK48HYVRjUz56cYjHq/WphKCWcwhEoqhJNPstt2y53EJZJPR1sBU63t5yyS8eYWs
W1YjdggcHaQq75DK162wwAzIGPUx7sswh+u6eAGfGNYUdnmupztZophq4TRhKoKxPO+kdyVTQM6Q
jChblbI4fyodvbMfOdHCEdGmvOpUqblfOduUt9VryKFIAEXt6N7LFg3yvbDL5vyXHenG/9lsuaB4
wjziQfPBy75XfbqMIc8BCpgOk+XGtZ9/TBdwMsP930aXroKc5jum/Z7fTpohU7lIMiZMva1uoupP
vl1CuUnulGeBp5dAf56NNXP0Sq1VSDAruhRioHbsL1bKaqXYYwMJN17jH+huYkQBitJnuY/j30GG
v5MydZYriaUoVTfIsF8iRT/QRgJJrVRsl2SV0voAX9QWt19WkGaOTcLpwSfLxwTvfx22AyXa51C+
fZAdrirZhU+odH01urikyjKP6Kdl2oJVuRsRV5+mzF43RFslgrgguA9KKjFn+RpPg4LdJDKrH1bJ
bR+NEM0rJ2MrAlcXk0pXpRrdaRFBm55audTo9fiIqPGvi2IVeX9Yr7Hk87Oqn0ZnFz7UjuAkAD7B
uKNMLc4hDaHYzWw7+94vxOBrPvePNqlodrpZGJU+6HHE/J0MbPzUOlXbugPI38MhyL0MSa67hsvV
G9AuVhfO9wlDM2Kig0clCCctnKGQqtPcMHDsBOM3DmXlA8zCaNZQ0nw8SwZudcO4SdROj1SSY4LH
HLWlm+TzhJihMH/dmUh66BXOv81XI5PpAFm3geSyChYtRHiiFbiBm3v9QxyqyzTlbivPpLAZmJvl
44PN2UJobDq7+uHwhehYXg4s7iQzdYbTmW8X8nxxiyQN19RpP916sbKeXCmJQY3LqkPXQpqfhp2A
+VBj9ykJa2Pe2dI/QhGrCz6EXkgyunWkEX4L89CHoOqergYPRBC3fO6iA+D9AaXHliuNWIX7gZqv
7l5PrCO321NIeyJd5nOxd3agOL3dWXUYWByoi4QrFomrWw/ybQlIE3ekhTv1I77SLPmly+r3VFDe
zW87TbvL95L07daJEGde3AdOKRJwUkUbWyOH518TcuFkvfy0pW7wKmd7gj3cH84mEQpE/X9whVHP
dtRtSMFuKqBbgeURHe8cxPbXZleA+jZ2Szxk5MAcKj2r/ioWCL+ov25RWGHHGN+Hm1c7dAr/uM8H
nXHsU/Zp/RPax/RmPBrslOWjRoeG6E/u1DdAt2m2NLRoK3yZ1xlBQTTdE+Zh8o729liW4KMRqT+e
C1ThyM3GqIueK8PR0ElXe9i8jMo4H3u/VFtAUzLSSBklXRIPSWKSAjlon+qA6EavkBGwjIsGdmQ+
PbsjuwynQ9ZyAl3nAEjn4fE3eqs5BL42WJVkByQ0ay0AP22JJQ/Pt0rBimfF9K/GzgN3xS8vTbj6
SMdZO4GlMpUIvXflkZ5ehcyVZJrIvo9QN76c1dlLL1Xs2fj6Ejec+nNKqCTJ/OgBxHTEwnIoz8tg
jBD+FOzjRRy99Dag29sTJd4k0oPlM0HalZuIoHhfzXVufpuFeUCE6bF36EvbW510tVpWaZ7rhQyN
BDPIKkFjS494ohzi2NUc6ROC/tGCCYS9Qeh4qn5qJHDJ7PS/jZrji48b+Utgs3QEx9PVXqxokK0N
3MKXzpP3I2lOSTUxCBSp7YupRjntSSx9pjdrKPdJ3uQ7z9wwj1vKqcocjAwomXlMFylurQ3J3czq
nB5uC4GhjPzF+13oTRdCINRcDKPta3G4nyf82qdcoYXGi8tdUjjOWGTiqZbz2xxTlgq5trIkulPc
3sU+Go8cOApXhjudyjs6DIYTElw+mC7vZd5ssw4BD0lwu9w6ww3t0nEqB4sezIIPnvekffC7l+Qr
vR7qbJX2+nVNyw2bJVdkbczMN88Uw2fo6AfDHa/KOvFcMnQEqrlW9yJsIUg4A5d/gmELyLeGB9cm
fjD1RoJxAqU43a54LrelWE8yAehT+rbOHu5DNVvrFYWxG3Pits8JwgaHilHwMcvzSpRfSIJdJyaT
fiH/iRyWBbXFOLOQ0XGSVnno08K/pxXJv+Wfc8EBd1FYtnTMdcGM2wFjsaGczoKz0XUIvSbcdbIK
ZSjF1Gzmkub4tM6QRig1DRK2aTESv8kZ8+TVnGC+b+J5ELz82mMR13NscC2/uh9Z29aNnljNhiHs
YnrGuEpf9lw11uSjNTvvjoHxaK+YAfThpHphJSWFLO0fGOLclbrhmjKvzoovOtTaOlkK53SvMabN
+6CFmggGvAjfvp5xJzzHRSFU3KR9SJKI4I0MNvC3SkAih8QQeULuScz0uRHpvE9lOcZ5ntD2hWXo
Rh2TA7CkdI9H+nVm9t5ScqwFA0GTx+IFeyZ1dHOUAEadF29UdlwOrXR8umPzJmLHDZ4MhMkmjC6V
icFhXo2dwmFucLiRn6GLnOF3l/4fsjHYVzE3nNMwHMuSigJgM1Bcouy4v3Llfn7NI1LtMcRpnobq
Ey6QsvXkq7XDrWwEfNVHMgKaxvjuE/xkiZ8+9wLNjeJGm2wRzzlcW6HmJzhHhiJhExc5e3CZdSGK
jMYCwPeFWbO5UEnjV/1Ms3JW6YbSN/baMyZozL+eTfbnS8xBOqGmxW/w1tAiKIA/BqZTNg11Os7n
LPi8muYjhRo8ml8LG9+ZCXzbFrPYJkeBRePQaxMeggWcf2WNFAdr4Cbd3w7bS25TCZfd7vnVPZzh
TB8VppdsQvWAvBfI3ej5FXQLwsLGQwVBwTJdcfyjosCU7LDSs2jsT0pMv/ulnjjpAX5lLy0AEAou
NZTaBv8E4cGAy1wcXibHfTx5C9xb0g2f5DaUs8s0i3Xkmwh4mFs2AoJ23kU3Ojfe/GxgbrnV6AfD
Pl6NaGPX2prlDKDd2LKsiDfjYFpqJkqEsfDdtmzj5hT2NuX6jHQeTLa5yxNuCt1rg+OGhah3JIMw
l2KaVF6yAyFdJLbDDvEDgPe32C4saceJ2L9q208/CgLvfX1v4/2CAjtrxFXMwWrgf2Mic2Yf9cVu
UNaUlT/QjNdO8orQXheqraCGQnUugBpoTi7jbVdAXLTKF5a5mbdj72mU4KxBv6OyfeMeFm8GI6gs
BGSxDV+4hjngNpOiP733yYpIq5XMXERuDxqK5awSBuPgdQNHlIUe+rc9gUnuV3+iMiDb3Yk6rHYO
K89h9gAE4xmYMVKYOabeHGhkWRv2bJgrpQUS/zT/2Z2BqQR8Rb+pd3uNY1bS1xNdk39fcsFsBbSH
amaoTM0Yb1vIhLyE2VUFQZ9P0IUmQIeEqNcNRrBdpnkcvQjgjd3J79AgCfxputHlmFVH4Mqpg+A2
vBTWufPj6ghik++ogkTFfzefjrOhzEp4sMrz69NJblVuZMssBzSGzatpmUwIl/xyQvkVEFQQZGjr
jND8V8kDB5I6pZWi/4BPhhci8kJgRLvJxohPQxFADCThW6ASOZm0Ez0gr/DhtyHDBHXdDuM0YMnK
UwVSkjWbIBYAdQ2JEZPK7aRHmAKADz3h9STeUy5Tj1daxc5d/tqt2f6WgiGWUDqsc+OJtQh7CMYt
1+BNn7tVNpu+LJB0eIvFwKWEiv8NpKMyXI5KpAbd8koTNV6qPDZk/aId41WuKT06VgUNLJYMxHB0
UZUOlLJ4o7i50tVr9kcQUGpV3QHiMR69St0JJMdvLVvW5LfJ4aUCPA9AeR1zI8OuxwS1Hui/mg6D
Yh/Xqemab6fR/A60JUO9J/oK9RRZOG6yn1Su1finW+4/Bn7Ko7FFJLqET137bmtMCAflVfbQAYmy
H74+iYzRa6RndsIW54V0seoo297tLjfhcq0bTHYAsCMFZaxxs8givSrCW6HaZB+bHo9t3KsFq+Q7
sApmUDu/fvLRyhBiXN+URrCPUIwg+4u/pWyscJLSMa4CIUrVt863j0wnPiEHUO12TyafuGcrTGL+
DOPqzMtsYwLwr1z8GPMt7gfvz3wq5R5Ntnzzgha8BLadBpEYDhMZqr0tuwmMU3loUpKHtk+S8t/l
6jBpUobxFDIMVrwfL2okhJ7Nq6aBHoRs4FTZr0mSU4LziyzFdepgoAvNG6P5W4PGbL/cOHLbysFb
ZWTgJt+tjLlbwe4Li2ae4E9bu8keMxYW9tYcwKRQc5hXF4Tc7WirFVC9l8rPhs6aL16Bnt8GGBQ6
Kbk3C8GONlQCdANcXwsn7rPwu85VxWJgkMk3VFKowt3+xd0KMo0chOfPDGpX5KyEOAhzmqOm5moq
HeM0E6lK9OzL4lVPEWXbN09GhQGQ560lGsMHadeOZvHtlSMD0JjGIIT8GiBhqOkC2nGodqvDdPil
kYnGYIEHT8d/vdaxDWkenkZeX1ULZj+5tYoV5n9cwymnV4wkUwGa9cH5Vi0Bz14O6YUK7PJ+xyqG
ThyemB1G6saj8HyragG0kysXuq1+110DU5dR6NesXzsGsw8SQznKFWp3nrbSwR7yepy1FdpqCqNm
jVmg0CzwhFDIcLmN7n1mNcLdZ1vkEnwVaIHmIQvc84d7sBB9splofVvpfWqgmt2Q8hcoSp1UrHZ4
SK95ea0DpBo+sc72ae30jKqtk5IhKMKLCapYQ2069SwPgrd/137PHgc2rFiiE5vFQ3re/TNaP8+t
BaATBh3/SHNnKRO0SLaUWhR/lMJcvhvcjuNPq0aptJDWwGh9nlHv1RtueCT38iSbEqHOwrctD9Wp
Ramr4WD65pN+LuK2mr/z4Xuoi8ClvTm3BQPRVY9nNqM9k2QJkKyFQe36s7XMmFiT+PUqzzC1OjkU
d6uaK5vkDf4Q6YC39wcM7ElthDH1CfZPz5hH/9cxD4o0NYKHCRudFS60EJP0vX2+38V9avPUGYif
MVPnJwVQz1mCab4532D8+0u3XFwjkl7OG6LXmdZnh34ahcLPRNg7yn6+vLmixxMWO83XZ0nwe4yw
tKIoZzXgyp1vdLBzrPHvPC9f4KW2lJrzKLu/iHvwF9MnOHtqY2urkLWCm+gkuoUSp0UXbrdEEZzt
1GXwr9Q/FdI1XYBp4B58nlhNnx44HslRL+wKTh8uJLrUyrMDprADPq4+fHVpUIMXHegPO+K+Sbxj
swd13hIht9v8pOeguJdzlnzKDe8IaeBycANhiU7TrGsfEUMEMLP2c1yam17HLz1stkAWPrsDv/qw
KDQG3/WsoahZDhQ54vhULDhfgy8PdEawg+aTwTPxADmMrYb3NVN0MbJU1x3fmPIhSZav1Wmv9Tnn
VdvSWyAVsnO/rfmm6E+hBjWzKzGjrmyvOIms68E5br5ZQdfB1UjqnZ3pOFwi9/kZ6SRd86LWxgRg
B0kguuxPf81ECBEDxYcGFRdqdQLQKmwp+Oap7oaoLHBRqfDnF4m+80Ce/EtpDSdSlSn0L9CeApry
IUor6Or/ppyfdR2VYaDRBhFHnMy872pcquwOIbUOlvtYa1+19JjqEuCvhkhFZ48B2ykmsQKuXOB8
moAg5WZqBzlsIkfiNC1Kh01cmAXcwa8nuiS1vbc3GyXPX0dx395RLDE429ocy4Ffj1T2nAOWaKx0
erVL5prIg2Nqfr+JFdkERXpAaUgUglo1ZfTSGWcgIUmAkLFIwUpyBteCkIlUvQMoP6E1T1JpoGuE
8VxQY53xnB1tC+H/+NUsdlaD4oTiSCSJtc4mLp+ldeaLL4EmoJ/kEJwcjtemK0Vn9MvdpLodcXO6
hwMpNApDrsu6wAQluyN4Ohy2cosgU17ma/xUt0nJfvrXoV50O/FN+fm31yIBHeLIMvq7jffyq7x+
0WHHlh1fh1oPo352RpT365z6FAAT1qyRhCi1aDIZdA/LfQp7CMPpYutPfBSrNY3s8CTSIV0oC9Eo
gz9wJkNzWBkJ+h75jFfNpPZ34mnZ3f7b7K8/RBbQ7WdqclM2KbxKBFp8E3pOzXMr6IiT8UBqIRp5
JKQ/Yy3V6Qoxw7x3T08EiRfpWmiQwA0iwGfdrpz1IEgV+B4mxJJa5x9dsUVyBPLuklmYGlut1447
fpoQZ8sA0PPN75TSXmw2F0YvjxGkrM9mWA6awdIIssoXuVMPCs8WFFQ1nQjhkKCpsaKHnZuPZ3Q1
Oojyl0SRLCbW8YVQQPVkpGQIATOgqS611iPWPuxYKG0/931CF/p6vqPSSajnN67dk54ncuDwpqkL
zRYFhd5eDGGOtUvc98NYyTK9FXrlkjm3dNmW1LWGbdkQmg05wGhY1sxuFDacY8kxZSVr8ZLOSX6N
8upXQBkfi3Ukxm/OsA1GPp3FvRx/muCjkNBqPWrcSyV+T1De5WDcJsHiwrNeVHNyhkot4Ag1y3p1
igoTLcDS2qOf5THzmIBS1uXMHZ8tOLfgH1K2pZfxODoKDm+mRm/xgGWkPTizvC/pxZ7jYuwPN66X
Kd6usi/hR6A/6NhnIt8QoLmP5HxsKkNgwmpYchZHZAx3g2JIGstwbMMceQPE/6AcIZJ6CsbKyXu7
OxCUvJGK/aIcu2fj/gBwupkcGOHACtj6vOdqJ8oVhcfaYj1TJYh8DkbqRRBdEgPznlh4AnN46WFk
JXQgFwT6Qyxw6PnP4M9AToAYZkD6Sz3ozaJ4jKxEy95ysyWmZCQD+k/jcxaaNaNiGjMCQgwueo8y
8AgiW9/8WlWGC49YR4SordqLH786IgJt8tJ4ugG3X2+kUtY4ClHyOqWmUy3MLtaFHaJQffZFpQdC
+ju+MM4et7NaQmQkjgI+tUYYT4ez4pRDlUXphIidPDh2bOqzrr9v4Pk4nOeabLhj40Vhf0BW/i+W
+6nNATZzkyITQ7IflM+cS3RlkILvayCF/LZTAvcEYB9NqWan6s3KLLrOrHlaCxxO0/aTdLVShZeC
vXfs4jIFD69FRi5hkDDoamopQGreWQt/2uLRDV30E0/PSXDSWBbv4T6hooeGk6gJHfGwNcKPi77a
KabmliZrw+IxRSNDEsZdAn32sJOEsxHSrqTNZWOZxQ+RTtyIvWbrb7ydGOZgSuhVIsLL70uZBivZ
UZZS67QiYqPHUAMtRy6z6qciS3kuN0+8iSAAcBKrjgDuhIwcPpE/rK7EMkp6tlBkzo6+RY0u0r1N
AxJi+4WkCDgteMhjtCdV8HjWbyphSRBSLgUZgfZN6Q7hI4R/Hq2oyx38uxXj6c2j95uCGxhlckP0
OtT5Uiq0Z7NeVCyBbCRFZxJ/AQgyBKrbz7JlW0NWw0xcVQgG/ULpcFfSsRbRDbsnY5N2kbZ2ts7b
zZbFSkSCD2si3XXQO4cR+GzAKBHPZIzy3t6Xm3fVItBqlGplyqboC7pMljcqr+sreGs6mXLqqiI7
cGnUCdsMs0WJpLkzSZTxDR94gAMGGBS+uB3xNbgjEO9E2bIZRsP1YhlG0gDdHKBFO39+EE+sPdll
oFX7bjiwWSMzunZFWH2LRqK9+GjKt9CQUpkT5Cth5RdOsU52aol8bxHvSVkGw1pKH/3RXEDLQcdL
GWNWRUhRTk08JhvAcALGgEvp8+TeCyDOGcsRJasEUbTm/JuB3Jyvd25wRPsVooZzB2S42uMMbbig
V7Xa6diN42AMHz1Opod7ZxOwMnTdzFmaUZw8MpQtMXzmrAU+Zfqei5KBnarFvUTU0eRGJhe5NJs/
ZYMrwQ+upylkbPGCclfZFyplrSLbMoYSLfVXennn2E4Xnm9KvOrjjG3CkzawxhMTFumb1uPOmEZn
PL2uw+MLJsMiwoPeI/w+OowKCccQ2wuevX+w62eO0lMrCzCxCyMUd+PCOGkCUTimQ7XvHi7ErLHh
MhwXIG1esREhGOyLKhbavnKYenb0OkcE6OgMZk9mzbjTWvQ2DVr6bcNh9OOMM8sz9+Q4O26Sgssu
bwIREjT/7WXdAJVwsRsn3heGn0j3p0H/9Ul55j1Fwjg0oBkPdTxnGg9QQR+ePsjVpyzhLKNEjFHo
XbR+edQccrXqrzlkezXmsXS4FF2Mnns3belSI/t7FBU2eR/wSpGgUfj/bJfp+kpN815zSsoowYok
dXaHKmeOzyoVRp6m/Z3RFydQKXNHPdDM1zcJeIrfASTU+53bl2yNqlB79S0RGom0DK/UTxRWkbuv
8S/gpaQirPEKTvX65B11fAJrtqs7r55tnPIAu7fLXzWQd8pD/2vFeiW7p7Jm3sDvVXnticNMcSdk
voMKJhOEC+upZWM/CtmOOlxtJakp9uByP2/VjBjbPGi1SF9K84GnH8M9rg3A3vnB9WmsI6UxSW+C
OtPrHaWUgXJWJlBz/zAA+3xsk5QdbXIF4cxm12Yn44oDXph8R5GOvMPKKP3AWOeAC151yzm03lF9
irb5/rn2JniBhTyG9WirrXyvYxZmRidT0bEs3V5B169OLDnYRSKR1LEHw58Wo8cybHr0YhGgXj45
nJgDqaHyRRODezKymFPHsu/7HpgQgUFmMk4aR41LDDD4Cq9GbEAAZsL978F4GZ9VHF9RkANN+5yf
DY2Cg5mIGTpuRgZU4FV+nojS5j+8TKmJ2TQytNBwCZHMD5UpGcz4DdOmIDqXXRP2Y0Pd0GXng2Gr
jfHcDLJmW64rAcVEZWiTeTMyl0fyyf2hPOuIOc9kc+fv1ixaF4ss/rmDM18mn8qBAIFWTujPuAfQ
7j8RsciXsuRg5jw3+bigJUPyWCq8qoTMm0LA6C9tnpgEIrQgTjU6sTMhE/b61sclFnnzgbay6L2+
N5Yz/FPD/NqNVEqq12YO2C8P7MM3QMTKZbt936uPgkS9Q5znKda4x5GtqyDDzcEJ5c8+eIrZsNjO
n8M8Yx+r9mN8wI4VUAnowl6Y8ajxVt9NlpLgaYSKt0SSgvVEgZGiHB4PgfPCGSZN0uadnMJbRVUj
3ssfFvF6XJH6NbJVS/EQODVBAVsC8BEXyFdzegDIdsTuaC1CnNCY2aD03oRv7aNS67S6+WtdUki9
5FgPxteMshr964h/fn8Cto1vZ3+3AkBVFI8ni/Ax4eCPO3efbxg4Te6T45MgQInskvOR+WNBkCln
aGR1AdNBPYbSIj+ODAvO/H2vJm9Ffk1F2yAJtmZscrYQB0TF5FoMydJXh/yUQRr/VZU/76ygFter
JaN0yWw5MRtuS/BjEkz+c2CP7LBSy/QrNMrIGr387d+nhl9QCd26GbG5UjNSPTeptCYsRqIfmR02
654bGdYQRUUKEBz6puTPP7tYwTUIkcswAnOmjDbM6XumBctmkYUHcFi1Q0HLOF0NXFD41wZtAuLC
xHCkxG4WPfLqb1GKtleAk4574D3qhcxfwWUfn5L1X+OHoAUtp4Tvi7RyQCRNJn4kEWggADYCLQPy
FtARMFxVpFh3czsfKQa7yFP3BHjNYrSlqx7/4V8xdJxamP6sUMQJne4HIaMkmJv4yYqbEEC4eFA+
or55eevdQSHAPSbo1FVeEHLvdZ7TE+4+DXn+TeovFzxijuqiz6rSwd1Pp6kLqMYRqvs5KyTXJEXn
GtTksXgoBSFIIMG75+uFOxYXFkmTG792giHIYcrKOqaQ0jDkUGN+J3nCDxcnrhNSF9bYjy0QZ9GR
BDIIhum/yeXaWYnHW+Q730N7MQDGt9GRhke0H2sHFmUFxImZcVYtjrB1d7ui1gliFnqIeS1AzR5x
w9N0DurFSp1l5oSNUY+ElnKAmlK/6x2ioaaaJJwufY98/qK6bRW62z/N8mCyCgZJsEEV2xanZ3Xw
dwrRNGaW3ebV8n+VrpmS72KsqWilf4W0RCfrHnAGbDOruNNTR3x3wl1i6d0CYCwUzvhbqfYpmG/8
3x7wgq6H7z2SWlJR8sD0OuCbW2LbPTeG0tAao0s5wBnKYG7MU5dm/RmZjU0JyHp8m5ESf8YR6Lrx
J5tjWYLAsbSCKeUEaUuuMVfmcu+AyOJleMUkzFEe90l4lyvT/MIzWZ582MO1Iz2WKAdMrF88tSDq
ezr9NQDpjGZQPcfrzb45fuASTw8P5H4FTvb1vO+feFUoOe/OrsO/tple6ceO+euFnoYBtL+Ia+mx
5corEMGI0Ix4JwgairNB+Cm+PFQgXh8ElvNSWEEVkSQ1qbc2UWXG51d+krADqVI8rIyK/mRUPecN
XW/+g3NBj4n+nGWz5vbYUWYUke8egNFnjBVjOmcBHqeDczqYeZ78twuzKMu03cnkqtqfzuO08134
Kdy2LsFDG7N0kwbIxxqmYHLHTd7SLEKhPct3ZwKCEqKsWKpDXiQxLm9vwlTi5qY7bAdUqc3X1VZl
I3bN7l9rQ8e8VmN9T4Dsh2tGE8x6PtLymVAi725Obed5joPFeia0uNyQsP+YnJVgTgvMkrzBeUeB
ii57b253BKCkjWHr4vIADvuJ/oX57LLhqNEoY4x6TT8yvrANOUSAQDf4Z66gfnUNvQPbbNfWGv+J
gSgv1LydGlUATVwacdE0yKHt42RawDGaWjuK4QaYhk+NafXACk/GMbgHmXNie1CrzEElstx44NgH
4KMoavBRaM5kH6rAplpZkrvzfeHHTs++dkbgAy+xqTzp4poisOBoA/vefGoL6gfc45jZIv4Fid7T
ygQL8OWoSONPD+a+6rT6ac82pjVWE7BcL3YCDQxM3Mu0gpYKfqGFkyRzSK3vpBHGoHmqY8JqX4C5
lEYa8rHwEvFw3ip3YGq0HUB86vLASpFBZgw6U7/uykD2CQ2LX6hVTRtKZGCHmBMOTO1n4i0+6+PE
QMko2O95zgAlW6RPXTJD3+nZ2QplAFFNKccoUwE4B4Bat7J+Mz7ZW8yWdF8rHSugIfSguAMZDo0z
QIwgC/2mkEEXVmlrZIchJgeKOk3huhDpJdIsP9XG7zda2Lx9mg38QjLHMZuFLVL1QCdTX6YMPD5L
Df3Yj/6yqw7+zd1sQ0ruKbRBMlzDO3h+O/JolJ76FqYiR0b6x09BlJ+JBP+3dDiUWvb+GrMz3trY
ZoibwOKdkc35Qh+yFHLUNyde0qmL8vbxVASyJd9A2DDqgdQMtqOt4W33ludcLkshlROSzya40phX
6X499QViXuqmM9PFXYyfPyGNPcSSpShoed1NyRrl0PNV8+8PP2E5ETEXfwRA//x9V69Q+v7vXHxM
V09BOPAv3o2CqFQWOtIzTGaVmX6Y8sESKaZGIl1jTT4AR/8EJtX3Z6nsrXoMVGIHLcET4qqw8UVi
9VDh1cmZftAagsehhUIQdkbZyz2zuHFB1lXI7FSdg1OGxJctxmK+79zuvGFCSVZowW4ywPB0f7hP
G9jbcCDChe6QiBOPkSG3Wtsb9Zg5yD4QReAyozKgnpBy4kxxF1i9gNr36T5Pqt2XtRxDrCB6J0lI
e6SXSlAgjld52QAmcJId6t1cvgtXaC4rXTDJJV4s/j1vKkxzLRgVwvVJfkhistFXSZKpmNULYSSF
3Ki2OozHmXZRA0hZgqVtC+8kALm0vExCiWagsJYPk0uweay4Y1+Y+DwRfT+Ynr5SFq9RMmPMNqa2
5O6h8Nj1FUulfn6lmx3aquagmbUK6EdY16IiA24QvCQzYDrB8CtbgxkHaZQfcCcczsVCWIR0biEv
cbgpWfBw1SmHYc+/CpttekDAX/ARsM+l2LMoIbIm05i4rg5x8eZg0ahLgOaUGmhJKQ7tf9BdCR5N
kqo/O8CiHNR0TXNKtmrZmULuPfge76RdsFwc/vSkgK2ce5bTFMKspTVDXoYWekIOJNa5UznIjY+m
u4WOdCJICMZjzqUgZzKjnlweVH1jVEFXWxnImMJkaSQnkG23bzzF5zBk9+AbFUP7FmyUKksyWGvC
uMKoT7zQ+c89ueHQTDs2civY3ZSoGDHx59uPuxjF341a+y5MzB7nSBJKX+9p0oPxR9oeQ3J4k90u
3/iwkR0mZ7q7xEuP+uTZDdz9ZoFVwfowgV+mOinH6mZ4T8P0hlXs7tv4CX/YSBjHhoN3IFieqmp1
JBEn9GcAZ8mkJIY2WO6iec0VZdfxMztx7J2o4f99gBxsQVMOFN2KdVcN/Q3vv2j6xw6PkPgqZsVS
849krEXEac41EyFPpEj7BnrAHvVvy2PsRujOBpP3fu5kvBcpGn5PuEMmYy7GzjuQ6fnuaptbteyM
yGWZGq8gHdHcw4NMU9L/Vw9RcsExJLkcUyPX6HuuJVc1Sak9Qrw7Ibz+EU51pQHvwnOSeikOVQ06
VBc+rjzARnjUBeI4VyCSFbKb+jPn0D7d1vmiP11dXa12h6nP+wpPlZ83wOAbUrf2PxWD6OTroEm5
LUb8O4qR3ADVzuV3e6UE6JDTl+Ly7jJl7bn9TkD5JW7qY2mzP7EHeEz8lTnKklnrvhLMoigti2LP
1O1NcqpQjY6iW1UErLRJvb8jlAQc7+IWknLZP22mvyC9TJD/R9LzRXVZ71Ad7qQhvrsc0WTcUYgB
30nwcfgNbkekl9NugSxZz2fRpfJJVeMSRCub6+D8sZf9CWNEdBgAjvNusqssMBGciLmUGRz1lvXC
ksh7aiNeDZaJxGUkKC9Loo7xHR321hcvccfxfq2HDudOji3lgrBWcmIKOGKBy/UHMaxQ6ISRVDEN
IrWhJR53hVTWEn9oQxw3tenBiH/lYuV2Ir9Qm2Yh1rwuRdfQgsJsR6yPNTuiGOV35P8aEl3rlx4s
UI4KQLPsILf/sKdMXssrZUQyU+IqqI46bNVGwUOWwsO2l758rwTGzJqMFeUflfNdQJ1kgQ0nq4/Y
B5+8Srev4yJjgx6JguFI+L072k+os3TDMQQv7CPRVUMBwidSrRrSfeSeu4TsYSiErIuwfwJBRW46
Hl4LwlJEowKvGlBshiizSr756Nevxn3KyhR0s8bW90r3NXd85CEpc5FQeEAoA7vOzdIFDar4Iaf8
xlJefoBmtaQg+etEN3jy+kFK22223bD0PtQRrBSXOuW6ij7SOtC7XLjq8AXP6UyheR2q9nUSbmwq
k+3bWll1AHwEUqOeNyQL5vIkfkPPBAb/iSYuIVI7b/SinpJDC3QtBvv3qGHCOuskUa2maZaqNjrM
fHnUApvelDZS1Fg+qbj2n5e8hJTuw4whj3JQrWV8Nxiq7FwnpFjAH5YiCe1HfvdEtIxlCRdNDpqa
qJcAnSqli7DrkT/agXmItId6bcK/PAx8G3QhzDq8nBa2bfzVX5hg6PzrWDJQ9gdzRQSyzs/4fWgH
1BZtDMmhiaZ5VHX1T8pvU/U6qCkREDtGxlJ3hYllk6OM9P7bjcLUtEDITYBZO/o32C7QrZIYJ0bY
sX+AahQbmwof1Ns6rSNaoZlCJ619wTg6FG9s/pKBqFR2l3pb/woFfpJWHw0UKmQkgAonVpqxIuHK
0Ld7jBtizdeoEcuGjFwbVVSXaN8F3Zv+Buo45svV9GjAzwIKUNO0N8agM+R5c5Zog+lDs5Uj+20k
Jbk8yY0C8UqQkWcNUVYp6YNbZijbEAnpx/BJHsQdRTXmu2fWY4EqMbseU301YM+rcXhPCWstZtaX
toDdpy8IVSPC/Rd+GqgieFLO8YhDiFEUKE7jBPa5yKaq+zIxM48XT2H8AvaHKimB9VVEnIZTiHtI
F9jLmML5Ux/y9KpoKB+I2KgNxa2QLmHPqryEnlox5zty5m2oiYLyIxF6VtyipcD+SxH9nwvBFWqw
p2RNFO2JhLiwqfJ2gKQZbSuciZv2Szk7lt6GObH7Ra4GOBrHefdU8ET06at2GKSS8gcRP8laFwcD
tT7MWTSfjUsgjfIFR9TNfPMJdDwCGMZsbPzXEUf8YPk9TqoDdtS6Vf/uTjEtHVgeApj9HDZCkV3g
676TTPBfPQiCnvYHUaDxQWvDoeQbQlr/AWBy+hhaEV60rNT3k1SQpybKDBI4vhnPMf0PhMokphNn
4qQW9YTByUKJ2L8oQlXGH40iOsA/wZJ2Rki/c5haCwiUbZ16zbWQ2WoUfJs7DSYosrtNR4zS7otR
CQ7heBBVtsZMeW5zFIrcDxxNVrqLBuXsOwsg4SGJBKXHKOISghqUym5npIOHT1xKJmYI4kbzkEE6
G50L88do+gq8x5jqzoLOgflY0Hfn84QEZr5fMErji5KpseL285Qiu0tZ8hxeUGNhtVv4+8wzPJ9z
7ByYa4R1VnZD6i2Q77cQNfbxfQPsbbWmidwnRi7rMlM1pgDw22xcfXpzDjCeAFFaFgYFaJEYW9Bd
G9kV3SoUmCQYivMQN+FNH7aYAvmAqgb3lmRfEUr/Mqtfxt48gKxmzJZj9m7hoKb0mobWu5OcdWQo
A7mAiXfXkXksSyHVJ9zWkA7oAUYKP+/PceM9yFSoWtqiGBcBpwwA6XzuT/yFt3Du5IN2bF5CcFO5
aL76/Y32+rljhXPmGUmlxAiJcwo8tyYv+wwxxXQOQvFZDORNczEsUCqdSni7tBe6lABwB39Yi8OG
ZPhpyjWxWS44t8oJSBFckh44/hGsDlHfz/bV9k0iLLGJr0O+a74t+IP1TZe0FceGqckFVtNFttOC
RzC69HaGr/moVJLy4XbAbZV99DsxCrL5ZHlolSleeXtL0c/ogV4liaT4bOjMXC4T85f8+O+Hgj33
g1vtwxNkw3FqGr5tLXB/dB/gjBHTZV8fO7OPEKz4lncX5DR+1WpnQr07uPtiEb1RakRzp2qs6/UO
ww5QNHCCCGPPu5qXOKNRfdliT+jGGAGrSGu26OWLh9f/CuysfZdjQhA9yd+NEaWsa+VBsGsClGE/
kcRRo2+oVdmC1p62raOUrni64px/FqIjyf9dy0C+h/9KJpSWxVJOb9O+DZU3nXh2vdau3IZdxig2
W7U13uqv3sfxZpyabS7L9dsfhrqtOXFZgcpDEhZ8Pl+VcGLrD8JmvPxhefeDA0i7Bx6oEVjcQL1z
9Hj12/rtVRerh0vNTDyxMd1QDtM2/LUzFEZ8+CYjCFVnrN9Ek2uIE8H/x/ebBaB+YvTLUOZS9Ihm
qXhVezuhacGh4ebCzGjwD4F3oWqAGPQ3PP5WTeJH0LRVN/STSUGGDXolKlbbh0xMbIWnfGrYNLTz
gteKTwgT16+tt8cmhPrhPUes3IoaLunTkco0zctrvsMF8jl4vQeK2Q+z3q0uWkAVK5oP7Mxb2nBc
ZTWUEi2AM4DVgmnQvpZq4vCdXWN7YeaeAcHiwqWNjf8gEzmaeV+DIl5WzDGB1+Gt9FhwVa4VX7vr
EkSvBAg2tjY5vpae5FDaky1n1hvQZLziJiaNNop3Hc/ZHAEeZI+E48NLRRvDhmz3q/fAif/3BFQv
41vFcFUGEMUglhxDtZOY+IDazl/MzGDG7aoSopHU3af9EASQYXtSNCxCfasbMoM+aXaf7Gbho+0N
YYakoRip6/vTxFsORDIWGgRDugGsM6Er5tA0d+7DlgmUq/6/8ajSYML9UIBiZfGwOpMKR/003tYf
1PCUc2hVAN3WjxC5hfndGHfC8zyo4ZxIttm8GmOp+Gq2qjbsFWdA2LfvE7ByPOcERgOvQUWk2OWB
BNrxZcotg8E3W2VJlGKpEVcOA69fqat835/Ns7dl5N3cabZAvLB2vkRnwSfmkL+UDj/Jy1YJ4Glk
eu4OuE307QJBgqp/9ovE24zIKZ+x1YDzxA9FyiFlTGNHy2YEqwR8vIV4a00ljtoia7TutNA1jYoW
GETwQwZM8XbKcrgskBeniE372dxjFf+iDGB2GHVfR4pu1kRZ0NB+y7LsJcMjtulLqqninqaSbFUk
uuzMSrpPFZ7IHpjzpXKGktTpoSW+wZKuekGHp5Snpvc6H6/dMWQFyUILR0g+EUgRhoqTmITHgCQ4
AP9JFI/DeYKnBH4BZd92LFxOf+mfNxwxXui5/umKANv385ESDUVYa4JqfSKjNDULz/6NT4affEnl
bWNd4dRPoEroL2xt6zKJ+bK5XXcBzTXS9H83ZmzXecUtIKsXjws0H3x3Pssy0AIAir8t08D119JE
z9pXsdoz+Bay+pyL2qP38zquyHXeIfiDbzKci0k35XWLKj8xVztHgNSGh+bua5RQjzSlZLf+utwh
F7G9XLselC0Y7q1/HlDoJSvNclEPp+dif8jmLeK6yCtP80nxRzWYiYiRAP5nUCbzbgXAAnk5rVgz
8d1TLACgPCeunQ2XSMSSXppFRwcfPMEnPFi3gqNJTYMg/DZNZc/XuDd7vgfVwXaFm8IpDBm+Coa8
DNSnAftvuNFOOX6e/9+c3mljbqO+LvxHLOdgGZ6KR289DaCwvYE5PMtDnuqGA05l4Zf3k2ms3ZuW
Z45RhJ0ddQdf3tvI8lFjk4MT1/rtY1OhOQEzCJc6DEM/B3fgekYZTsVPS9gnQvWjW7HQFBhbjHEV
ZpIfHBdac2DrGJGjjYLvPrIq+yVgLRUDEk/kYRuBwNmToakyQEoWRTPL6eUibCQ/DGcW2bjkM4+W
3+jyG/h0a11mhx0TlFafxYZ1zmXLrqAIw6/vO3JK98awxZyE4byr5i2MdhcO3bvnvXBDOkBgzaoS
TlMAlOhgRj6j9EfMnt1JI3BRJ+cL8e7QG4SPkKPGSJHBc22lHmYeSTUG2DRTOvrDNaXqTJRvUatd
APTa7isDsSM/bou0KfYiBQYSiWv6nu94Br9W25XgVNPueuT2cEGC9EqDpoEVqMEMcwnoRCjqp5Ok
7XRWn8TpWn2X/NxYmZhps5F6RushHwCnNPrcnLI5IhKjIUkpVolgzgKsmPzvxBJ2FzQYNC8BVbvR
stYz7UyUEP/8NsnW7QDMMUOGYN3YFi+Cn754Hxwc3V0DfE5fZrjCwkLJ7jQe3oEjPQ22BKyxAugv
7MPvnPygE2QpmdI9sQnayLx0U6gXfY02+FScfUkgs15Yay+a31T02hUvRO6NEfSWJxlXpf87p2eK
km7WuOcB4j3w0kIebDNLV3p7mqSdv/vHAVGZyDb/YE+Ncx1vzsUvjnRWVUi2D/GwrYAuZY/s6XHr
QRng9WTKxlA14ZtZoPaw52h1QNZ9e/wO46bJID6uT/rq7dNibP776hhlF6759AM2zbj2skkZ87lT
46SUHEweOeXu/AHx345C1M1EG+mGvnJ2QM47W7/xSRpv/HFdELyvDu6BNnxDE6SQZg342zdYFZuG
ZlykoOKC6vVNIFQyUSRW257VQq/zjZzMnxePZeM9r2sSE8leBe9a42qKu063U0gWrSd6TBCmD7HL
waHU0aaVl8R4F5lpaagQHe7pvU+1Bijj0eA3EgezTxPEvSZDqAaE33W72J0XSD+Ym4/0/TgxcYp+
+3QzsMgl43iQuv8mibiHFHfLEeO+rFGHI8lB3uEtTsNxC6yI4du8G9dDERzpoFM4NUlT/lnQ2iqD
pAAkkhtiIWOPGC78JZPklR2Myod3vZEhtjdZsMzz8ByjqR6QOys+8OHZDK+2v2XzyZfYGj4FFwwl
aC+jVcTwMwhcfOibmfab4rUOxAMAxxarVdhAAkWLPo1Ru216WBMdyT1si6hrAcUqC0VraXLiQvGQ
0S0hp2vYjE8+P6C7WRa36rcDswu+zoP7JX1K5L73uOaJ1wesqEtUGR9R3SUA2msOjcG4iTBxwu9I
NWMFPeNfIhqihB69nxvgeg8DxE1nAP74rbN/K53NwX9zQKe73lHtCB6uIN6jiBIkFiri8iq7C6R5
hpVAhy0fBNeaXPn2TUN3Ui14WA8u5C8Ojyxxbgl5saUVPc4w4ELcXoSNO7KzaA8Nrc5PYnw/18ff
srLaEpKC5Ug0idJ2crBGPh/5YCu/kTS/d2YMKD4M4IJGWbqPnmbap6yeLOB1lJbhJ6rRmE50o8YG
x+bg9LljN8aH794C20VUX6+20qgCDLXDTDomfW7HUiwBnxKsCD0fgh5HTO5ApO5BqWVs8xM4idf0
zysV9T/8CreJk7kuPwIOlYnHvuuXDauQJtozGaH+7kBYU6w3V4r8uetUMKKCYR6dMFkqymOjYvA5
AYj12H2g77UhlCm1VfmJJwf1OrJsQTV+4qSufSXVDGeEpa1IKZZoK+TnooZaRnOSqJ6OZfTA0ovV
ZA3abQRRGzcb79oVm/hJgunJgTFNKQUsEU3rxpmc5HfVL02wfBI9mLxqrrP4e6t9M1A3NXFzxP8P
ZThcJ4qM7sq+DYBPYgpXhMEuPKbYF1XmKwlcBK/bR+U0qj4DBg//IyOZIEsBGIkqnLQZOkm3qGNj
EkHK7qTDJqwjozougvR5TC5eyBpAfRTxtje9Rl/RsA7ckfge3mXmOrJB8zHyptU9FMl28Ss6DZcZ
sg9JYdfFNqqEUFUdU3+DJQ4ICWcOo3/FWbHSYQlSM3bxxqQHN66U8UjhH3O3CT6TjHteMb6Z0F6H
3lCTVpxwWkkjc5jVzBs8QgqMRiuLaiUEg38aR29Pbj9pKyhAg3V9cpdFMZ2eyD4tb9OYIEdlLeGV
fOry3jHewx6OwFMZUDRK3Pzb+bBAp7ECFuSZsuMUy6pKlkCTBvRNFOZdKKeL8vrayN2ebQbJdo0Q
pOgc3p3k8tUdmWKAxtlt/oS4+eRI7bPaZUu9keYCNTCt1noAV9aFMLcOW6rJAhuPlmYwSfAnHIUt
g85njXJM4pDaoVZsTPGFcFTRhjfcOE8WHxsmEqmIJwOaq70lT0nI3NTwTZrYpsV7r5wsMGMSKTiV
vdZZSxQRsmyPm/x+J5r08WMK0OqZ7TL5amzt6+/eBiEy+uhjuJMvDX0tl+jgNjtE7PmuysaFkekC
HVJmk7KjhW1GuIWzz3wjV0UUrP1TjBgOnSZ6snT/3m3GpvF5OPgF1fdckJFW3v518ZeajAdZpMZ1
+TlXJLL0loYafKZcK9JdjdjRcfak+E1bQpIzybrUxjIW5x4qyExejfNPIjo4cD0rrFKSaZWEcevx
cpHqFkxym1yLfCE5EQlllnfrlz+uWtmLM+A7pyL41vxRKABVaFYxirshASNJbBseU2wuDx8pnMRY
C850dsVQ41Czs2unf0n5JkXfzwNUmXtNdGXAEPMV54tx3JC68Xt9KUzgxDzV0pGNswgLkqSmXkWx
82UsvopseTOBQbGu2XxQtLsgu4RGI3DojdG3gQzbx7C0YK24kuolGeccTZGvi8HFIwysh6lYnm/9
E2pL0A5d0BR9sfNNNZNST3XsA69TD6RM3Zmb6tp8GtZqz3h9qObXSCVcKeuvXmJmq24F1XV89YI2
u58VpwsQ8/I9sG4hY4r41Ct1W2yEgkrIlU+aE59XTuG24VCEQnz+C6YW31lG+cV95vBs8n18Rl3B
afmIGDw1ZFaXr7pOudLwhfqs3n5Ouc8ZhvKGi9OgXoMJPa5e9zxa7y3nYuD6WC2eb2y4QK4jYcTf
JaEyNTYVcb0JDnmhepPYwC3AebkbWatPoaIXE0B72eFg7p9gK0qQryriyoQX2DTjuXRL3U2yto52
aAY/NaIXLx0jtxnfE/3nsVBgCNtGfa9mkmSUowhYjsXOxzrQC5goGjeUVeuc4AxVpl2jC6O5nVgw
+YEn4cChO2CGIb8EpDklh1nX3k1Lcx9zwzhkv+ZeM31oW/INv5yjefVzpzmdtOCqHmYpn9Ex/VEt
oaOJlSfVrMeURGzOSc7LDd+ip2CM4VqRK+cpf2G8Z4PxA7EqENWkkedctXzNUpfo5M/gcFYw7mlj
2vIg+iIfIhJ0vYVA49NftjmDcGL7HoU43eVt8sOYOtt0EVOiMRpXJD1pKPnIi9qMNb2TCzPWVGWh
rwV323x5vuK/uMZnek2yE4wuPwkV5u/s06M7AWgj3nLO2yTKrWhXgUday7eR7N72o+stMzgqOica
MDHw4BJaCAzmx072phXUMS7V3jP2VDU9gx2hBB9dTUj35c+6Z/DEK1bWexFph8XENgY02JKBdW9B
8JySMd3c/2X9i1r7xJTdxLJUUwHf3iGqBQh5PS0YAJgIW8MWmB7jVVOeSs3C0iqokzxzie7UUVua
xg3ugqXZZ28owezKGfHA0cYcaIJIBJ1LcM07P4i5pJNDDzgicMLi3oMJgLQm/j4zwB7QQSRl8WXs
iy14Ecw9o2pM1ZGlCOYG7gSdvHM78d513hV2K43n8GRAyogsh6esRMoIU6tAkGgUDNV455iOFk4A
v2AYcnUiQ9oyRN99Dbq9UOZ8bTURmWTg6vIvAOi1/VBKMVsP03iYI1egkOL7o68VOYrL7oUHKfFy
ssc5HNflc4lcWDEzAxDCoUjz0VMCitwgybO5jBZJZYxBlclVzUi1t+7AK8iHaiN714p0GqR/QnLc
kwhpGxCArrPbLyQ1Mm6h8h9tyM+hLin5wnU2OsQwu75B9g/J3RCa2HMeGiqIi2v3QOKRCOeriJCn
POjuFwWfa76yU4FmmXqEXdbSyC40gmPhboNGCjGSs0C2BwjnwWePT624ZA+ds4Ky8AG30zGoS7Su
iJoAU1n7odg9CqS6ZdmzcqwwKr2BNb1TdtpWcnlUzaCmY1mz3OFDDqzB6f0fxblIfxPr6roE9xD6
q20NsTNC5yatruoBsEfwbZew/5Jt3JXxgVxKWEjsOMUEYLtu8yQX2KLh/dPEJC3UCszvy1NiYX2V
5WYptb+ktf13azybmd1COw5z9Y6OdZJtxUSpyjBHZvJpJUH6eTGBBfbsHDNRShUPq349s6Qj+OoY
kOpOrKbM7NsTXWN57ZcjvVajz6OKymPGPnXneeztpGXahVH8KYokMBqRv7zWroDM4lLBLmoJNjYC
rGPxlD1NTgiZhxVxuynKBGExaYcJXNy2l951+tSgHYYminr3cCH6a8LCC0IiRgks7O8G+hb+J/Gf
oTgBEl9nVkGZhjP7ThPPqlPeJ3EZ+Nyq5VVcvB1xZIP0rg6CAn1IDEa0tBhdKQONQhfX4trdAEvi
Hyd7c2mZLefgDuuhy2kMyHWySaFvsupfDDL3yOcwsBTJen8rHOam3KsevGHbrw3bazIbFPKZ/1dk
o3pz/GRZO/SCmRqyLn+EQtmaE2Z/6kST5gsLRUXmhHOGJJFqSFIFohdMWTnlD011qFIX2RBjiEDD
L309Hby5FdANEeim+GB7UqQBTiuO/T0/AodnQ2wl6aqT636W1JVGYZZWSEARAVFp0bbIZM+2C2yM
wb4kq9zUTZlAL64sXeWXuWCoeOnQkef1oOnNuxWixco+fIsMMRwUkDuJTyNFbAFYTAia57tMXVlz
emkIcwQ+z18eGNBF+6iXMLwg6482CLTz1NVzVKuzNN6g/yIoAHq5a/aWq9fBmWPk9hNMZITyKneB
y2PS8h35IvVI5AjeAjPLctAHFUr3YJkcIMKbh1tEnYe0AJutezpK02nq3/6XD+JVcS40LCLlBE7W
f5bD2boG2RwpD8Bw6DnxgeZcxPXaV58HqP4/Y5EPypU8lgb122jmXMr3ztFTMVJ+dMqx+5z6apD0
AtMr6yjarpxG77KM1mwi+tN88nATgH3z+EkEuKRK3OAt3OLF86avtjWn2tHiKUAFH5UyqfDIezpm
PyvEW6kzet08Oa/zV/wx8bLS/b6VHWfraB5kp9kftyM+FqL0wigJt/Zne5XaW4yDqZZvcBeoWxdY
DYAhWYyaTqzr44q5jyhFuSSUb/CfPQEahkODIYunX1xSnVkxQovKZgIxiAWbMeyipFkMMxX+v8an
6LA7qww+fqnE4E7S0lLbVfn/LF9/idfEUy1j5li362JHS5RUwALemqFcZFtlIlyAGMiZGZpQz5xY
b8VYddYkUC5SaHbEJ30dz9gGaqd19qowtPGpMUj0ahCSfrdEDK72viWzxU56PzUD5ddjhedBTqGy
rB1HiNx6of7y9Qw7jpzKduRYRBgo+Btc1UZZfbCxh5gfW0ukmQaamvFdHr/iw/NLpPgZcg5YCswE
Q/xgs73WbqqesPvR7YgpjtO/92hbucIxl1aV8FPrpgxDCMDliZ99wMforuNNKweAaVh0f/oDKFwj
vEjS8JfBht+DCF8I+nwQ7/4c9qpqCLTpxZbgTWF+FjSd5tQkQeKoqJM0VdCQ2lYEz7a04kw90hqb
1z1xgj1w+UnMWErcbZv+6FWCK2CSPQRPUbiXBIjbevRsC0JL+TGgc982HKeSEc2LKgRMATnIoMQM
uH+zMx9SYnmwTUwHVG6MQfGhiLJ6zMw0nd35APCL9s86LqEN/PgL9NX/segqine+ZTV2EtB4ahUm
EfWKBJHfDgxRQovjwRGVSJeD6CCZ/D7RycmvIC5ZqaIfT6C2FLEJTK/ogEciL+/pZYp38DG5PwNO
MZTWYGctZWxldFtdUvtc+Q2wMmohR+Ar7OgmT09ONOTPqHipvFtWFxiTSU+iUBM8J8+0tDurC/8f
HERPVxRSUfBU90mOYs74K8G3ABke6yExLeAb1Qj2Ld3LRvAwxV+YvFbf26awAWhTJu6uNWo3Z4e/
fgxqtGooNvqcQE8N9gl6V2//H9Ri1RVB4iuRvw71DE1U83Ns6vM45glvZgdPsBnZXMQMREfGhnWP
ToFQiRYurk9cHGyCrLtGaCnS2DmswS4sxLVRAT0WcDnTWs5opYt8A2MoqnNuahzq/nz1C5phA/M8
A3I99U5mfUT+dBxsOxtF98BCHB3FicFf1kWMfHX2ul9HKoCPVBjsNAHEi5+B5KpJAKMBsa2D6sHJ
86TvYBgp98vdGIykVzgGFmOlDPLYKaElVMMvXFCoHqoz65CfSjNlng+fPvSQuonGzTe5Pfem2SD+
2m0l+NwvfMlPkUHOjdKVFGVB294bN+/Fz3ftg1OiFp914W/O/6D9gI8WWpdsdlnpdNORoO1swtNZ
RE0NdGCXFVpqwIfQYbWGLyFP9wJvpyL7G0dxXkzRRSPCuLxQe/e3PDYHbt0ihr+g5slh9BHgWcq5
rkjBIdoJ/QHG9m2OPfKllSZZkegzdz26xVHrANDK9LI8oFBEviJ6F5t+1ewn5aSrrFET5661XyUK
l+SM6ZXRPBi8cQdXhSOLhEhfwobWTrEbjFSJn18kU0JVRE41Cou0j0jmHkeU8MlwKA4K0uociGgi
zk1l5OUEILKd5KAore5R5FO3nCGEhP1jTHXfnx4wbZTVjgTDi3FKj/Ruyz8FGUQy7gXeMxT9jONf
PG36HAXvps8lCuo+ouBOcY/eb79B9q0qgBKtyp47I4B3Yn/3l6zabQqrVbTnDHai24eP2E+EBCOM
kBvSIDI6k7RYgjsbFSikg0hAEL8i7FQIXK6o53t8YhPV8JhhwXCLtalmFKy/2oCzKBfe4cqqzZ1V
Vw0PwWaDBZcuS4ELPmudZZqBylfJuVMAeVv/mPOe0fWzq6MX+rfwwejl7Wwho1nRnBx6c11z0Fc3
MFYK5TJrHuhrTm1vts5gtYfHuEhJU7jx9gGRGDfMH2iqbZAblGNsbFwYXby6zQ02FPLAntwmp7S1
qHabUqGkqFSuxL+VioL7D94fTDZIJe94indHcSyX9v9abZ0IASWY4BLAW+S97NzEwH/QEyHfZFSv
CCD7wxEM+GXQPYTqwXIvlITAtg/RVqOAqV0EtPalUOacs/jfJJUMt3OMnQ8vHi0z5Nw7iVEQdTpa
0f511OwGupU+k3bbHwYKiqeAurL7W0eguJY+nzDi4bxWwmWj8GJwVJzEhOJNnCwjOC8l0sCHF+9G
ziLFP4O0FTbVs1u4GyBVQvhFF1xwfIPpXi5e4X/1VjECOWD2KOFSDim4j4PRl6FruXfO8Jp41XHo
8UbuYmV2YEQ+NmKDPO6fRoX7JsmExDPRsO38WCr0mUr8WdLSIPpaWVrMeoHuZqfq/GyvaI0CT7za
s394M2u+ovHCWTC1d2BOjdu/nu46sBCkBnhJiC70Ul9+VzcRukOQiRAXAnfF0uOBZsC3qvD6/s+5
VYxAbTptIWe1tu//jE8aRV8+iaIJuDtIQE5AWBCs3hf3U687nogjVkhEK+nU4+d56bZ3i9clsVEf
Qza5TK9kkU8k53+AUb0c0GcU6EplTlriZMsf4PeiHHKMzbj++vJGb0LNisy9/vXNmLTMvrUE9seG
goR3PVTLfW4FXqe0vIitvJ6xEf0JYu+9ag92zG5Gz5n4ZfTibCwGSyqjBRPw6zBG9HnES3N2A8Vo
4BnIuT8mdBA8ypMjLxiLnT6n2rLCq+GKgrylolFNzLIUQg3SdTSdOIpxmKxyCecQh5m3/q5ma1N0
zlgofEXxytjGfZxMED047ehKlsfZnL9McTUWME/IaH6I7F+lGA/CIR9O979qccMJ/VwlUA9/hOXW
5hKOkQ4V90qEgaB5xETy1NnK/CUSgYDkAgiAilNNvAL7ZilgOtVWyNK5Aom1K5xuPl3L91zJKc9B
cGZirygh67zyPhM5cHOvb9QjGFBGvxOIqkfUAUUXw8euekxzCUpHFp6qPMPwcirhsuZaYpZTWXbi
PYDF1NagNvv3vb48J22ErDZRevRvcbr8D9jCQkj/Qn49coVKCnNjlyMUUmha2w9ZiAvfpRBVkZ5A
1VzY2//65jbZQXoI54WRne+2QKKXw5F7wJsaHgXy4FXbNhXUl+Ql/v8kToW3Ae6gAx0ab0rwvbGx
8M46eq8ttWFqz/K+xhr3Z8l7O0BocRmoKJ5QIxdrqxYeMk+/TGJmjw5nh0g1ul9r+xNJg5kGBZCg
ZyjtspfhK0lgZAPfOnIZxYL7yDVkNqHK/7rQfWQ4mbPG2YXC2YLsw5qJ0r2bpor0sel0dpyTL6sn
mVGbXl9+8hHZlHDhiWbELKrdUb8+ptE/As7dRqmOqj8CuTy2HqQ2LtU0eJVbc23sBSEuTw/RJcGC
uE3YeY/2de2szqQ/WiDXIyJDYOSmmgnpPq7mhNJ155QNmk6Eaz1pfQ4bMufWQLD0514qPvCZLuEv
PEiIenVO4DTB5M80qTiJ25VOdseBHhyOTSeyHsDx9m97aG863RV3O3FeVnpShcFnFzoNjKC6SBAe
KcifkYLbQggP9i8b3I5Li2m63z+ErOUClCOcDBeOBHodCEpqr/zo2Trrc0HcYuIXkn1OYLvmn3dR
Tf4kAdMU19hBaPIFxqnrcccwNkYbo5ecPt3+8+8c831glkpnjSsExa6GyyFWoyiMdE3UbcAGTw9G
5iMiR9gYcohzaZ1pBqoovDtR78hcnubVbtvCGCHer2iEdeYrzdHEyBXjJXxrCaaMDsOSUpYLdIzo
h+urjUn5j+VG6+BGAlH2uRM84Z8fd+cDFCl+Db82mW6VTqRVJfOM7Pe4/r6GL0yJPijAJWs9MrcD
uTPuvvwmuhDQTKJ/8PW1/ztjCp8JUMsZsi7ybPp/XAfo2mWhX9vjPYgtDVzhZqjiufazpfyzmOSa
+tQtGY47sOUkzO/scTW5J4QgQk97GkkZr2Y33Vi4Flw0H+8sRDtZkzE0AVveV8nGNJzhkX8ohDFp
D4Q2SIgSNSNzdbXAIpPmUKzxEthJKu/WuC1WnVumxQ5x9RkuZrgEjs2BTdxBC8loVmLUnF/Z3mCC
gBJyNCMMlHxyJHeJeURqvSLm/G4fGPy+/pIuGOt9S1baxs/t8f8yicBVRJrIJ6ncaLNYkIo4j0SZ
yh0ZCJNU9tYT+cjrj7D+8LpoSIamwwBbKMBCR8QrMmrC40yz5J5kNcp5UYk2RPGuZTypEC++rlr6
h6u+Jmke4o6rM0PvjMtuZluVA8Uh6SLut70D1UMmuz2He8al5KsjsHSTLOE4ZxEhT8bk5rWTb1TJ
fYeWNUQtbM8geqp84eLO/OVpUMPYNBKrqMyx7ifqHERKiG5W0ekJg2vP1A/DTPpCnf846XQgmO1K
UK6K18/HRZV6oqnqMolBBA369JaM7J6WXDJ9mxvF9dQCs2ptyXY63Ey/m9An+J8CofMnWyZ1ZqCt
krO8dQlUyqtOrsRQg/0GHOFkzVFMLUtUC8xxvraCHFVuj7v+60i3V3F/fSatrG4SZ/iI1fqRrKRK
ToLi5caQbLoRMRItU4ot9PqkjlAFpg4dPZc6+K0gI0H958fshZ4XycEnZfKiJSiB9lHvAXB4nHYO
WOLhUGwHacBL1sWRGo/JokjZioF4o1E4QyM9E3+EJuK6nNSdr0HnudoYDuXxmEnCmdh0X41KQHVU
MJyT6qB1KU0X17PUOs0QXYByxh2Zh6BqEUxUZ3zt1qZnU0HbTs7ppPUbaOYbJBH53idPW03x1Xs3
USJy3A8k3OZG6047RSWcmVQT10Moj/PR/li8CjH+jXts6v9rgl4bbCl02DWP7OKNuQUKwknkzroz
XBwD3R6UQPbOalil2Aznf7CfhdRCOHsNi7Umx2YGFeOmpBgvOGjPMIwGHZRgiHRi6aKK5KSmjwtU
6Xim93FxHW0ZetpKLNttroyP6E353dd2x5DMkqvlaooLOtoHtwzkhHPIJ9qe31TqyseCx71Tar24
qHegASTkMgKkLLXHCFQACsFAGoFd5w3uqR4vm00oheurWepr/s3tEMI+PRprDBt14624g71eOmGs
0YtuNTT3mRHdDq+/VNmABqY0KBDx80iIDe63EgdnTb0UO5qL2zGizitI9OrXY1S5AW8ucySxn7Hp
/l8nbrEkekyNJdI6xn+XQav9zGDt2NBfLfJmhvEfULYWhJCm+7X+BopPj70KSSbFfYC8AOKDRivr
47hM7iHvO0R7+U+QNAhtvzq7c+bzrztew/LnBWfhneyWgFQmy5tJ9AqdFVtzVNrZnqH/PJ9AoK5H
zZFOf1chT6nmfECFGCvDsP/RlaZGf/w7TAF2tnoqNtY9xYCdZmRL34osZEN+d4zbT8/Ao01AQNk6
OYDEZVcnANzY7regRN+TMAu0bUtvLb+WT5QVlfPoHqeEwLsG08TNKbd8RuILs+cIekAwAvb8qDI1
FPZJL0+zxXXrYXysNuz8itcUNZhR+W5OcBmupPl8q3EgQ4j9RooToiwbkI0ea/Jv0Qdl7xuM/pT4
JcOBR1SUB35xcSs0OiF6+eeKtSgIFrZ5ttdr5rHesqy8Ndk3GCS1dWeZQfro0hKVSGZFq3vxGow2
YdtbHxN+Xws1YxexB6Wh5TVGR01lVUh68JJbnnUTyZT0gdG6RRRnF8/r7imEFFqM+Qg915hTNs8G
Md5iMIlM/ZRkwAzLV1ySOa2kH37KnoKmR90BgpuZ2eJ6YM3eJEBfTcC+P69rEK7PrfJeWZ+Mz8eN
5vaa4IXVHlpZhiQec4WEdIifl6llvkijlyKytIHdGykkdG9mdRJXN9CC7ujNMqGwrSe4VInWcLdB
1WjD1JM+IF75SXHbVe6Tlf7t9bZa3SCeo2AUYvcfp9lBsRNIbD4O0CI4u/V/1Li2JlGAneEmIge9
MMKcPdFXj8Zy7soMhL3QX+wjKGyEC7X6hDC0lxQjz3ahfU1HWHg4iDr4KIT1hfQaOhg41ZPtix3g
J8OchgaOinmAcxk/S3z1IsscUr5NRNqmwPYQJ7YnU50RHtPjWRHW0ErYZyPGQrM0tpPuc2E6d2NQ
TIov7Be90u5JqTr7ywtvKqrO8pR3XLhxdveO7fDBBVKZngzSN1mBCYKSmCMNuoql4sUl5udxBlQ3
gohDmdu1K3E11oa3cLGQsJwa69F5qpo6PKLQusQg2pyWwZf9EUgFOh06aDZy8nf6mujMEpRoA3nG
5eBKI9+p9ESP2/tO6+9zDDWF/rujyJIDgaRMVfrpD2BRblNNh1BhX5umkJv4mdQJQmaEwRxXZuSF
lmPYDW9q0XeJBAzep2u3OUAOSSjjzoNMiTq94mOlynKYmb1/xLZxY/XEHrB+nqJBlxyeaurVGkkt
ZSs6TQ7dglO+uC6V6lR9vO/RJSAcCh4DxjsemIuQBYrCKwMbhnls82G9hdkm6fBWU8IQq6dtL391
Xks4HvoKN3jF8sweu1taLhL7whveSqUHuICLaIAtbW2zsUCBtNcRXEqWEURBIDtOdU4wRPCORd6G
ID+5KnJGjorjI8ECwn1xI2TAbwPLDyUGXw78JHlLKUYSnfoGiWb3BzDA26PCdxI0lPTR2eSiIono
zomDqTBi50JgU2asY8wpRT4vWIcLaoAoAs+8eoblXCV1jDdCtZM3eG6Pd7giLlzPk1Ir3MK4wtzZ
GX+SLSXf7A/XjqqeQHZrM2KUzBX+7SLHaJnYqAxNkCHhrdbKJxKHLTa1LaDq7+2rbUwsGNE3eiUe
YQroHqwJrgmaHZSLewloWjED9VP+MFCfD2QfHaZXAqjlKR6CnAJM651jdTPUVP9ZwF4mg5WglRDv
5SnTHozOxWx6nKqQTeD/+6xvP36uJn8c3ftHzHwulBTfgIwAAjihUPPRFu9KLO5Uoz4uFdBKOjof
n5bZ46wgeYiy5z5JcidjO9tTw5MAOAi2y+jmwxWzIGjku+ZQ3IgWnQDw3WdHTcVeVb329E5acNA3
GFQ+oPKwqSTlItAW4krdoM+NStYBc6MPsowm+uhmyu6m4LCWQfUbe/H5RV398ichnHWTP9uOphHY
ydBdCVbw1uNUQk1tZ0WyNIGusbgxytWaslBcq+ny9WxZclhp+skjJzTSaeRfBO2bqiXYGWy3182c
zL0OaFprqg3vaasqeEP40lp9JWiXPVoQHVFS0OabssurdcNYKW0wBt9CNw9EmJCSDSlWN+ku4SG/
eCilQ0qZLENH/SHmmS+tuUVOkrAXQ/wDCpESkd2TtvvxevgWoDzjFMrjLYK9+0aOpETNbcm/pjgA
9VARgH89ktBRixO9kyYFaw87WC5ihIawOYVBpiPm9bsVhJnPpoJe8NFbIzcoZd+ODqFurqL9PKGX
yqBW4RX60EBWy8uVvubo1eoYMxkw9EazGpZ4mcQtKEGDC0Fd87/K1pInzHZ5Z9mc2XepcAzFjkTn
cDMiaUwUijbTG8hKzPZYBb0RbwPi2eAingaG7QZ3H49zBfr+0nFHOsChSjWg1FtwmZrnOzmcZD2g
UpQL9//KSliVMI6WfUpsNN4WkWh5A5YRqwu3y0GoZBQIFzS1XbnHTbaxd1fl4oi8H/zHr2WPgvyf
xAY9zvebVargmyfKfNGCUM4MePW59GSvOBzax9rKNB+xXMC8dyQoORpRYR4FecBlsQNsBLdVtfes
+X2/LOodG20DYQBfDEEPKjBBLnK0cgShctREQ+bWYpZJGPiQiWHcNCj6B6q2WSffSqnH4MiBRy4E
7tT9KvmcrwxGoiiqB1ANIJI3FcOFaWoOlTQl2iviN2xnWlKM742+LN4rfoXJx4zBxzmi5RyA+/qi
fi2rMlJ/CAtKhLmNfJFaIB/PMEcZwow0sdyhyC63bqeBdpmTbuh+lq5TiaSJFdIaKfYwia54yEuk
2Z0hdmdKLzwDJ1atXoTE+Whxi4PE0JcMSjOyJ+ncYNhxtds7E/G/Hi4pt3fub+D2q5xHpOSDQZWA
/JuN31LsCxI8mhFb3QNoAX/mi4+9b4UpLgmO0lCICFvVAgi2J5TaMFG91yvhhGYI02Q+1YP5CJHC
HCcqXcFAXbazYb4jMWRKHz/nqrOM+HabiGlwekx1KRFe6eO1NbvuboZQ5rXPc25SiEe7zY9kaBM9
6wYyafZixx/7XCVpZxXdcmwi9zb74XlRETT7h6kQ/GJOTcgkjwFqFzKkfPXL/sMyf6jcL3ARGdVu
Jl9WphVRxv+DvBfiVtab1/kxfWsGsn7Cf0brADEzV/bT1rJATSKkZiZZ02zfpoXbXQ9DqMGCisX5
A/yMnM4bkaAEzey5ipsuWzFNXp15Vk4ylv9ekmADJ6JYIZnwQNzvh8wggAylvBs42sVFevrSGl+S
zFBeg0/n33kqSYOXzlwoLgALjPIJkwCRPK8H6MtKrpP7CRozfUwfA0AqzbBlNLNKEYj1EgDof2Ow
+WzV4Ot1rRg6M8dRriYvln+zMaVQTTMeNZnMt8Kbe7GwyrmF6RBrXCgsORfAF6DZe9O/pi3ejlhF
JUNSRIEK8K+hqVh73sp+BDCCujIXgvzgr5B6hh1ErFIOWaK3c6wXRC19c2Vkrfr5lBNcnbL7EJd4
OlZJgZw3RY3fH+/THh1bHPsCnZpkKEzwCxuppgFuHGDo7zqIH70/AJuBH6UgO2znkS3eO4ieQ7eM
2sEXtxy/QqPEdHO/OSnMmKgyMBG8eMV2Ymzk9yZhfkqw5bIxhPD1M9UySZeIdKak09vByG01s9Ad
WiAME3OySnJ/5+e2A80iLmfiof2eeYXxIjrqeXKbmuxEkeowso4bLYbPwcQdRfrz4QkuZm8BRlRM
GUyuN755sBvqCmHk9mQq1x+5prhlzsoc7Lz2smpVog9aAdc7RDKU33rECAUGm6zTsRL9qbaa14w8
HLh2xlp/Ck6AmKJXzcEah5Pg3LlHJtGmdu7bUMbO5146FHs8vvgXxH6mo2HZTi1SCIUzIfgPJNCc
9TBx5Pi+Y4qJNRK+u/fjfb3MT0WdyuOIGNSolrpmn7vZN4JT2gsjPrkGmKRLJwdttqWZQJVeZ9XH
rlPVYKyiwrB8G6pwpJqfnKIeQLKjCoyCCQ+raR1TW1Mfk5nyahkK3JGPaCBJVi+mz4tzdA6hIuPB
YiicQlQcqdPo8HF6wYPI3mUD0k4wHE6dHxSawKiVYRQegX9sWNYK6ZG9Vvoz67qNKHU/EEjVFHSs
WxqhlHn+bcaDsR7GR6JLTTBJ7TfOJwkgRbfBfuKH3DbrSCyehIBLlEJ8+st1kpQizWsmk8bOrfzZ
6x3KhQSMGDCEePtLqTkLABCr+j7N9xQ8Yv1yvfrXOS+X5kiAKl0etbMYjouG7nVl+5A01naD7M/j
EHIKfRIhYPPbgxNG76tbFeymmPiRRnJqg2yMRhQmijdL9Q2mLGrP/pP3mrixu0xPAAdPCFDiw1CG
MpRVPpyvYX8hZ3BmGcrYTR7f46hASU/CIA4WocwAnC4Lu6WBOMspIJchEtnfDidzODnp25gLmqJR
OMWP7k5bK1UD7Jtp5o7Mcj0VZ0R+Eb1UCUwm1Qm6M+EMxvE5ZrqWE4v3+6a9yg/Uz/bbarED2Sr1
9Wt3h8AkO8Bc4DfOeGiedsys0NVw4hKeSp54Y2iIJ+gxlBEJ3RInfz/Bt2xxr9nWMPcvdFU84G5P
YymIPYqdvmw47i8DROh8272V9+KTqUtibk9rrpp03WYLdcdkCrrp1PA5bRDuSLcUQC5eP9ofaXs5
oYk5WxJO5UciceuSDpiOwO4tesuUBAPSYo8XqPZYlFdqrb5uVJq5DTwQs7h691C2TfUOqNR2mvps
PxbzNRQfDOUmaB0uhQbpR9VLjGxZh+dv+h7/9Bnik3yBnIjFdSaaDvayzZwPiv7khvvdTNKpVwKC
+P0oa8kzAGtQiT8sIpR2p2GM+V28MferJhrJT1rR1jlTIinntjypcEqdyWxfY0tQIaV9TRcw69kA
CyiAQn6pcoxQlGyJe/p2eeeuE7J6T1CpEf3ktTsnlk9faTz7D0g/QtJRLK5cP2nv8KZlp8PZVLby
Xfuus1PGW4BpijMj7ZgNy6rfxzq5izsjWtsVEbK6Bo0c5pxmNHfdb9RjDeNbvSfLGtxqSjbDOSoF
5vCKKFdwBleK1Bj5ay0kxBuyQdUlt7kwuEBiNginUkqglWajAnGr8gkW3VY12tj8BOzN9hrd1ojR
OmA145nfM5p9w/wTkT1yOrPUDmKfncSw+UFFbWjBiY116PAKdHMu4JK7UF7Gay7zXapJgesVnfHF
dGBCPC1MKGuZICPLxM5CUlmjYGPuSGs5DkQnzb3BUEWIvKY0sdKCSe6u+NHlU8Q2aBBR1s+d0eo3
LfM8rzpiDCUx/DXvc15b3FJ855WzL0HYj4sgTlZhDXSKLZ5DXwfIfOG17TmDuBBtGx5zLuy9rU5D
tAI6KVzVPvQ633+vdySWVHG31GMg402eO9xDBmzmTmIwxBsL864ejri1G3zhtn67592DY/mUedil
awVk+iZkq+kQRgcK5ArE2GLWZLr7YSfhecGSqY3XMSFNj0nTIRQsb0kB8vGgiwgNZX/JbUKs1D7+
vdDlVOc62B2cbaopkPB2dQjOyn0/gpbb3vPSr6AGmvywTHhZBU4noEhOrhryYZMEPlnP0WQ/CIlt
veOTF0sLBl5Ns8UeZTE0W0OJJWFCeVXV/HcJbJWd+CCjqCAhYAzTub3S5ORAXppkUpZ5iVs9E71+
oYjvw5E3AsV2mITCUwTH/n0btaLqQpEjwImtNSZ9ZsrkoDrxFPWFXGjyieI8qP9X8jzGfACt/x3T
/25ZiVqoPkRvi+2wCq/RfPWKOkFIyBGhqU+ak4gQdiA32xMIZLYeR7/FPhOz4ejeu2qQh590c6Eo
oLpdp2CHcChSD+n+CJ+DIMk7I0qwnSZn5YTYuKttdvcKTDQFcFL7AjNlmgjLGCZMnMUqieP3lVL2
sHXffjvWQx7p+j6doiQaA+7CHiAZnsDfoxsgUIibDpIWVVQ39+oZsaBazc4lGmAqD21J6nJIqx3+
ZcTC5a6BCfeShHzfOGMQWb8y7nFIrXGlXzT3zvZtfFUICJ1dHl67JS4qJIDHoClZE+9r6fUQ3Mj3
a8IIEdKk/uQtZ8cHseluicJi3W9n0OOKQrlZErD4sPovdqrrhxa4q++oLW5CDKTBZVRVYgMuW7cs
mAS1wBg4hFwZ1c2HAhCsHaZGuxa4LhctN/lfl8qBgEJzFBjgzlQE+OcHR9TC11IBxIUZRiduBHYR
kbr33rkuq/u24XwAZymBiLJloE1Ush50hynh/MBkp3iF1FvdEuWRwX29QBkOajg+VZjM3Emx9l7E
pIxLpWwOINp8aiscaNSZRghRuS1CwZ/X1P6ae/T7g3Fl0ncHDxoLcStWjElfnqBn2m6qjZlmALNF
SZ0yUnWpLYZjzwKh+lNYhfT/zZ3PKu+E7JMZdpwCfx1H+ByPXgPjvav879anGcxc6Usx0muVe3x0
XoCEdmOzmn8GR2Jzv21ZSzH8PQ2BI+PQPVQVgBIh4g52g4//7BL0a2bkjVfyg0o069APclGHJdiy
nCF0ukxYahOqgjhMdtOE/6OYV5Ov6a8MYVoBnMvpwKlPMyEqnFVvjD0TukXJr3qGlJJgTwSXdzFs
VCocmNsvmGrVOm4MakCl5GvMoKgNF13P6uZjYGJxIhyQCvo6UIA5yVqGJ8gI0ltyEPRs4bzyKZ7c
PfS4V0lXKGTAmn0nw665A8X21g1CIx3dz5RzOBkUufBKvmE2HZ6ZPXvy/BDWlz1+tcpxiTSfAU6q
O8PmX37C6Wf0Ha88VTQg52fPjC3RHN5LDrc56Euibabw+zMZMHDCGr/YNDBF6CRpcy9SxukrJIvC
KNPTHkdmNyal0KMzp6IFT5i6FOToOOE3jW7/c0604L0HbhSQe9ky+6nnl/Z0uDXleFEDhWI1EhQ6
VRdHAb4/Dp2wjwZgwOk/QNgUZ2RfV/vvPZD5mUIqPEZUueEWaY0B+TvlTIvuXSazR8+UYMmAreN6
/vnbJ0f4rn8l/yjWT6YHZJ4NnEb4lSW9iNyjBYSCepbki2nrOO6HO6nhBjNIwLZ16DBfWNplpeA/
g6VEKK7p9aFGmwvKxW/GB0rfra4rkuF8w1uF8FkNzcYMDTo3VYTRuI2FO2k1gH055CIC2iO8vlsQ
JrizxJouraU62/NZynfIB+lxweZhuUZaTaKOMHvE9N7GEBVn3veehfrk3ndfavtc8BBaGCyfVRSj
V9KHqaMlfA8GqLeiGA/5iu+g6c6uy7jkCJtAxKwDlppLc1gVlGLXDiNm+80QnSRtc3pp+c+tah0r
GT46Y5ocIc185qbgOMGnSYqaMALHPgXh153xrYDZijgpDa+EKcjHC3RgcxEuKkMF+Zd1aOp/kM3O
WC9i6+W5wpyP07BViGXS01CjdpQQbjwuuAsEr1932MHpYGg//dYIZtZJIvmwJc0jcEFpY4PkVo5u
AjrA5olmx2idqEauogpochtkxN9opK+9Ho6IsSgHfW4lRdLq21UrTvd8hmha19GdqAmEM6ozlaYD
S3Q24iKI9YQkG579SEHiqfikCKj/mr7hv/IzXsLVORzhJ3mMSkW7x6i3tbun/cGkLM5hgwVVSW8D
/B7PxE9BddH1XqueXhl6ERdd9CrHGubAMYtdngRVXG702nJBpo3SYaMGj4ceTEMrW13wCM9uc2ga
mbxIjMw5IburjMXvnbDbQltxSFp3iTQHVbMvUaaw9PwNHktMYaxeOA4WOu++k2CCfani0Qe9rggY
RkKCMkSbs7JczsIEMuCHvfzhQl1/R/Bd7X5V+ZR/wnHDkYamwLVtBKDGzdl0FnoyYZCDNrKc1eTf
z2BntLe35WKNn+YHqCKxqPvQTCzJD1iI/yI9kA9hTK8268MLAUsgjzSzhQXSCe8rWapnE26z64FP
ibvLNnW0nBDQ3CHTNSh/TaaZhJjai5WVdjY5SAo2wrfLt/x/ebIDSf+C38dCemCDUmljIStHkDn+
0aDtT9mgV6xaHEdmgcvm97i7rpU3o0qwWCU4GrGxsDLheNubh7MRc2ft1d1qDEVSygbYZb1nqYrY
w702Z7EpuBOQE1NbXM5Sa5bxUPiRuBeeS3vrQYbozak3YKXNa/3iMyYEaTVEfxE8rZ96c9YbYkRK
tqSWpGho4rV2lgsxEQ60stvaRfEmLSS6zskGXONriRKwGdNJK/gLP6hLn+KIRxtwXr22M5ZOQVGR
R4d7Z95y08Jj4RO9imEGmuyZA06tXb4YeYHiOR//eARasVu8Vti1Xl1T+IsZBYimp3JEp+IKQVlt
ZJ3HPieq2Sl+o5TTb+4/CUafnPCZmaeW+cxEL2iSpG/eq1BYbv8YW2zw6Up+pG4fNVP9GT75L9Eu
5/0ebFSPI8flCDlKHIYwVVP5QPk/lg0gW3+VIgTR7vmS7uOwhgejNSa8tWK289TsP/O/7MqjTuFw
wxBh1Q3wN5d06F9hRW6sNU15o2VxJp3fF2fbH3ONVnII+g2v9X6O+ltopGipLjNcdg1to2ffDQki
V/ALFGDJ8eaB/dRo1YtGnpdDyZ4EXKGYAqFfTc/mEJxYbOrc4H96cl3Bg5ITWaGCYYXZp30eEbfp
QGpI99MPcwCzqpIohZETw5rHta8Hi9hDJG00UcCh2kT2UceEGnLLZu4x+pibiuDMxFUkakELrtzK
iOM/wCJbOH3pJYBpLNX1+1N7LMQ9AL1j+TbdHxuBHz34+g1HR02Mk1NGBiESsxoPHRDGXGXby3dI
RVhKlieBE0yIo94pJfOKt0QpiQ5OKT6uPK1GXqersTo3lO0HVjCr10nj1hu0qmkwQPA6DA+4Njer
YxHTvaanFFrTz/MeRTpGx118YJ2RAmqoCkKsA6glTuFYCniewZiAVjIVOtZ3/cjMCXEHms74yvjK
DvAllWYeeeI6K4LPCuVtH5Eucvo2kEClHyeo0mDUK+bXTQpCRXUglUu598Zr4z0GSL6ih+83K+45
MJUS6Xdb08Y4L0kw7pFk8kkLAc1egg16GL5JnrrW8KuCGHIhanMb1UfI+/SJTRq/ywc4FQUV/Ojb
cZMk62DT3n7cNJHr1ddoaQjGBhvGDzW0nQ+viYZ+hz3vs6n5MCNDIZENAmt91nICKsCzBBvkaRiF
DsrnhA0dhLitTg1TZXmrBeY8h3hGRvp2QhP9Db3Cc1rrhTyqoS/ZsY7maDzkvpQTUgvs3/TX82o4
E+6Lgl31ALgxFf18fW7bfO7afmtN8vksHQjLT+PGQmdDKbv79rPPvzWq6eCchtcxkxSS6dLKokDz
mQHHyTKajz0t7x/XyZBjUetDdR1vK3Le32jBTtskl39IMO6Ga6fIds1fGKBvhHT5MYOA9gBiHwi7
ylCG9rRxGDUf6YetOb/KUcWFu4UR0CIJPJPNMP4djra0aLUuYu2mnBEs5+nKifJqhsEZk8faQWho
vCla9BmJHhZL0Q9IOtYYr8EtBXjLcLxG1gmOaMqnYKqdNy4je8QsIIZpX15zVf3HWkbNe07fITpz
2hsCkTUS9IisFIGJzcIXXngNjRJNyXrlEJyoA6z82y7aXzcZydWVdjmyHHUIg6ubBBijnPwvvJA6
9G8BBYuV7KpHgHNku707WcJuQPFqleq7yU6VG5NYfn2oY6jy0LXv2FjOy33EuAl9DRUBKM0kyl6H
4UQVGJIRrhGLUU4zH3x/x2maW4Zq7/frFHRSTkhuH8YyXsEj+v2M0QGYSNFEGSGcDBJaCBsK2NFS
JLSOjkglYvWw28gv643ESMuS7zbBEI6LdoCDXnJMzHxXPNKkI7kfF9OdWBeMrxKUXFrRVgDIe3Oz
XWzY7q/quYqc6c9/A8pI+5mf6ENDVifYFaU9wZnP2Ddfelpqfbpwa6pwxTwc3L2xPDlWXz7QZNWC
Uh7egEjQjsIAknwYBFw4dBvbUEyAhu4I5hhgKyJVSaj9bDnsd7oDK/s/bGpxooAvsw3rEjAWq0iM
ZN3vYG9eF3vXXdFn8E/r+fzx5wd40KOeHD9MNs7jQz1k9ovjjbngnrDeT0A15jhBnq+s62sIjTnB
xP1Med+hVH/eg9oCatmPCk3PTcOu3BZhayAkVD15Jv5nV+MkAzOpf46XNh7VCAmF+mmueMAG8VJ/
KOiC9lmueZrAK7axRf6KOJ9fSBxEXFFZ7FM4CdJptKfbkxJvNrIyGd8YhjIQOfDCA7+gsQO8uT3w
q3sHEMeKrmENqAxTQzl/gMk+lbKNGujHNk/HW9RHnx3KIQAjThaFuAn4oRnGWeQcaLvWxYZhgPNm
LKLay2zJvlvtYGOtJnhI+B+ccNKg4OL9pTm/udcagOhUMOIe8OABCShqNmGw5FBypRDfD5ZYcsDE
EBuXNWa1VuDqo/aKL33iCkOpdSwKRMbgUBAXf++ojNkkHCBP0+OSGnq926YDn1DUMzaJeVZpvqxG
Z6JiIzTRYfvW59zFf6YzNwSBwCss4VpLFdAB2BGfgyfTe21c0bpbXxmST+1757rhh5Q0lUotBzxG
bsgOa1C+/zvFj8xczmDdH6+1x0C5uF2EqtThRM9DvN7jDuDE6k71BUX+XLh0jRWufECMxGXBYCKv
5MpjsoFD/J1DMtC/eAHHhGWfuw+/8XxXZhRYdMhCA+ySYHN/KXwORRQXsOaPhKgNg8q6TPU4gbSO
E4JDwIGac56rzcrFtjdNKVbatlb6w0u62efTEFggz9F/VU3BjslsePlzIR3int7t8QvNT7zs9y3s
nCU0cdZ9P4T5DlDCb8AMnMMEkJHNVlyxGMWfqKHDYQS+cBk79Mr91unQyJnTFMufa7LOqUkc1iT9
f5AxqTnH8/NdlXfua3E42gaocQZ39Eh5BLhRGa/9iTfVVK/wrw0nkNRo0a6IhlBq+l5kolFfRqop
raXj1B9v6rKz7FxpMjCoQByTQ2p1mmJEmK4V/HSlIoMhqk/AJ65POSTnVpZyu2vvYZcPn6u5NnW4
ryLBGzc0JKqygTsLH3f6/7tj7vTieFHt1gpYbwtgjc8n4zcJ9wmqd/TunMkKhRNe1VZZm9zCPrdj
UkWUZG1gzLSwtP+vs8v6paZROabTktBvkmBh/hGwPospTfIXtyw7g3x01dknnwvSTOAU5sVqv5eL
WYLNZZ/Lj4EjcJ2oUXBE02zFl/CZUtjmDxWsqpqxgctoS5LwW6IJ/sivFjVzXjO5+mtoSFI6HrLL
urzIhSVsFS3Y1u5mU3VoxAa+kWCv2dajFdpX57g9KmAijl4Wa4Uo+1AIN+1OZSuzQUeSwwfHHzSz
UJahh1rRFYDpVmCpyHYtAYdX6y3fIOJIlPlJw+4qCFqr/UgBCZS73fhUF/2CRU7/Ik/NW9TeXBL/
KJdkug4BA5rQ8nEooV3AubbESsyhHCsH1/MxOOQ9xPcTtyIXlXPppEMfTSOo/V1Bm1nIW99pCwuW
SdS3s70NWmcq1r3MvOV1Logt3J+foEqKtQaVrLDh9HTFIKPmNp4Gzu2M5fmung159AHrpi613gYP
fxP7rJ2IjteU87t+3RmIWgurTEb16J0xHQRwT1XLKBq7VhTbRDh4bd6IaACvpfRIDyiuEaEa33q/
yYgwa+AI2q8qUGSDBCS2pTg387634w07GFglZ68VVTIp8RdL9rcWLEgyOIz6U1OmZQP7N7MYpNuI
/Z30DkCINQNMifc/6KZKk9XSIrPnvlyuXvF1DPB12DvmX7OkXQGr8Dca7jzMwOnuAYm3B21/lVyF
yUEnjVA5IjCitTXUJDjIQdjjpwSd6fQ3Ms2vQknmMLlzY+VL9RND+M7WfIg70wztECEX1foVLLM4
QS3qieXNWwPhVFNYBfGOCG9gJK0oBbGRTd5Gk3qI8M6qa4wvswyKBj8cidqzFXg+SC6jPxXy/KsZ
VWyiC/XWrVu5n2gUWjuGo6FwjIpbWTaffTYiw8hPx0RIKFLYK23vElYc9AcKyb2eRx5iX54QpXLj
mkDzMcTDybwz1szZHI2NreGpz8HAwONVKtkyv8DO0FXhhDhVZs6e5I3F/0NClq3NdR5EEzS0DlM4
elYW5fyCBh8K19ATmeKcwPR4if+QyE0H85MGQSpnUV9cb/mKbAqDRvzj9WgFHJnD1TYLnVe0+0uQ
3DS5ATfNp86VHoeRVAAwNAezZiBBXA+JdmytEzavBLUc3vKvKTW78gF4pe+rpXfPmh+R3q3FVzNE
UqPp1QFRgVxJqTVG+Y0zhtzy3JISMVBSBB277AbhWHYXZ+2/93/xr3Th01nJ001CxUvDA4VGg3Al
VK8DOgNOsm8biibv5GNXcoQBC01D3CMqlkxlsKUVzXT0UxX3HFiTltnErwy4ACsuGzlLcNKlvzPJ
ofYKlyOCt30ur8VjSas6eeWrWQ4CwPHF0pnZLwJZl2zKBHitWmvDEe6bwDhoMN9rllLGKdw3E4Wl
dmc5GU2QOVGpY4q321uKh/CPcVkR9OzvGtAlWh2Zj/tV37dUfhhZjGOZgG81wpGtHdsbpcU9yfbC
wm2XnSTajzPGe4Wmx/vZirFQKBR9vA6rznB1Pd8LKohnNZxAauC3ZNXREYWzhjucEeQce557IqSW
k88fcMBv8t0Bh1A21Uq0om4eH7Rauhn3gUIDuagyZeTQveL3rhlh3ojPycYznhmEo5VN9yMfJ/yN
e5eRaN/05IubnGsmSkL19WDgv74nfPVLS/MQwLhj5eaPoicbAVl+BjxMEVoQcQ/0MzOapPxwhdx/
V5PJCZmV/FaR7RLBO1Z0+KsihtRzqGaA2C7IQGrDd/4UNracVhFcITxg7nDSSxIqofRCgV8SJ7Jy
REtsuMjawWh7g7Zlt9jZCRtZdQPkNu6f0w03Rp4tp/69s6Ygndoi/kksXsN+rET4Rc9ORWOmHBGA
vipd69R2BsC6ZXKjhOjZx1VvaigA+OIq+ypgSW+ItRfzW8gN17BE6SunSXJE76fgqPDNkN384V+R
NQF92OM0dzzcWBKtfr8pITSTEHrpdaUIZ2qUZGZb7L0Ss1g03pUZdE9AENfaTIRDvjjnhj0I7l06
Aqi8tmaEXeZ8MVTSYTyKa2DAU5LC0VVqSP5PTVkhyac6r/R1Up07DV5D94H54sOVg7hicufGzr5M
PH6anRf7tgll+7/xS+YBvqv7juRu5zOpxFGXSFhktUNGQ7y8KWJSeZmsc+b3iCWbrRCTnSeD9pyG
ACCtKzid6e5U6p1Up8SNuXGDbn8+a9iMGFRA7+s9LiSgxDCw8e6uptQL+QXoqmCjvBVxVa7TiEOX
x09WVs/+grw4jxDGpFeHUFZDTS12bBds2J92GaJ8vtIeYd40tpgVfVkNuVTFIv4hwcxW+9SJ2wds
GnsFKixqx5tyl37RVtPlIFsYjql5tbyeSu3Z7iTQsUrVYvTaDUHHZxDmznSyumXZmz4RJ8lLgzxw
Gt14fUnw/QUYcUyq5SuEU25zPthXOxy9HQgQW9jWivZdI8UbRM2vRUU0Wm/zZL5gBzUZvzSvlEuL
dsSlb86dGfKFwZAwpIhO8pmpaXrIgpPErMVTmxnQLybN2LMrkZYEPSBPsg0sOM+rDL5sn/7q01NJ
qm6RrpYeYOdx61YlEXDVDgZm58LX8eEYnB9cROkrcIJE1qjn4jyNAIvTYyv2izc6tBX/MlDa+tcY
7HYqPsE49+rc2Ndpa3nWpYc8PbMO2thprecEIRwbrumRZ3t+cMu8Ma//5wVu+NdXxK2iAm6YGDzE
XqOTGe4JJDVbmXcb6lfFhcwx3kZgm7MPrFYmbTRUMCDO1ovYse07Es1C7SvN5aW2NXUK00vm8SXg
5SG2YKvwNsyJX/GImFKPaWmKuF500XhMNZSJFoCLXIradWEPG8s0ySEYLimEFKnOacW1k0gPzhcB
4zZzIYRBKnSGYDn8EXsx88AGwodEWxzZdDhqZEPvEbJbaibSW7VWch2Nl+VUWZ/Pnz45xZa0n3vB
4ASp8ns+wnc9nBqMrBIPb3d72O/5TtLwJ538onmpXS97Ud0kT7Do7NUvsDCsNH16NegwhbCwMa96
VMEyJ0h4qCNe6sZ37dNpHNfr1WesXPa5aXCEO44gMZ2ssO8P+Y9XEaE7TOEL2TFEbUL699XP1foV
B/8HpR1xfTAEBBPj/X+ntdrN5xevN8Fg1GJUQsZEkX+FYtT930pswzHBEPTGO/S8Y756iD6/T2uN
o8q5/DBdFcjLijJoC+zJZEmgOeKodlIrPPqBlpR7hgadAfTCxUH0492luyzfHJ4b1+ZSC8zubIm/
p6j/Q0zbgbWwZLlXvR4VeXz7VT+RzfdJ0EdtO2YOHPbld4ei9wt+z2ZVyloyFGaTFqP410xPosh9
zn6G0foJH3izA/eEmU6VDZCoDH3ZaJFL8MVXhFuhzIYEpAwVkiVkTIslofp9mfKZfTWxVkkbHQh7
NokD5qOVax3ORYO8Cscrjm0NoHAl/vu6fDKclp7Jv2M2HG0d4rXyNmHxtUxr+gMGsNGPDoaVwxUb
63OOb8FhbWt4SO5AUKEf3whDjfN6RauEzOGX4CB9tVAGDQCGMjx3Ptp2r29g+k+jjcnnKMFhOA+A
V1tnBuwfjaxp66/Z7xgm59y3gECrB9PbNTnwJUZsb2EGZiYfbDRHFOZlqDlmj77Ts3fWxygZgFIK
i2LHYslotJ/ex0OlIE2HnTq/uCT9BT6OyyiZ5RjgTPBM1/+7MaT5yqaArERW58yi3KSVD6lUj3xF
RpIK6GNIAmte4yTIVXc55IxTNq60gxz69sJKdObw5iI7P4x8o+X7tF7jerp8Q6ZKnl5Qe/j2eCZS
dnW2F8DLMyzN0HbUHaLSJ5VS0lxcqAEjNTsFOXQgWaLjmOpDrp4k/T+wyZICrRuve/zgXK1BIdNr
KpLIH26Fmf0N/TlRwcDjjOtqDpwWJoZgH8e8gfX/0Tie2x2LgNxKtFXlyNaMnnmbzwuvCl1irHkH
rsLFjkHzvdxl0cHjIMMpqLH0hnsIym2AuBkHLuX0vxTfmnry0q7bdl3lo15N63FThDcrAgFnNqsW
ySPXZOLivjGuzjb0UFGVmzEB/xlg9fmxNbsM7tQzY4WNcxEY0IB141x75BIiXXHUs8XMO1Oi3DYZ
hbjrKlgHwOHEy9Nzc+VClozjNPVDrxmGrYbyDjk3jk+LDj78jXlKaGPCN3gw47IPR309lwXfwP3m
fpaWvj1kDO0v5PNeMOuvYEuR5Pb2lbn6bw7LmX+LRNyGq5XQjDj3RKlEYjAO6aoS4M30GYDqyF+t
4n5sTYbCn95LGYlWBYXmLOEvk11KzGAgpXu4zYEUktmskxQtuLhS5mKTDptxvVotstHTeeii/0B5
f0XgtJtz7t8o8wHLETARjJDnW0pS4i0Eh3Y5VcOvg9BNzFcwR9hT3pq4V9D/wRMIfHBloWXzeHMP
IKwaorPGP4FALts4mjHBbjbZoOdWQ3U21QOvxwZVOz60NWYGy/sYD5CCsb9VCXf5vkWnwi7Ge71Z
HaRrtEBkhawrN9tRro4deMmmTS/urQ+ecIJajCqGHH1fRIgInQjyyOVQgtBsPVqOMcAV3TPE+Cbs
7CO7n2FDtx9tOpjThde5PhCpCW8sIRAwxJuyhdiz0Vf0R48Q0OC9vMsGOXCGEgijgjPsrxG2LPsR
uAyZugDWuaPL2dXAHy1Oat/Waj0YGCnIVum+4dsKfXMRrrFlRc4h5YPG0Gfs9TCIPbeMgtZeOxZg
YNHUnAXMSYqw69GBwhjOU/f3TkEqIytqTTgts8mm9Kg65b9MIEci0uMbtWNWtY7t9PGBvWHhYuVZ
dwZ1jt8/SKCbtcR21G79bM1Jacmq12plOb4iF6N0Tbo0Fn9PwQSnQqx+Be6fCxt0jf2qkWGiE8PQ
FdHgvZMYq5HaXzpJUl5JilV89+gvIVoMBKhSw4/wcCWtYeU08jcr2qGcYHFQ/zZusvVvOhfmnmEl
psIy+HUe0JYxtIiQnI123+jZPjN0FRZnopbWhk4wa/HOU4PXhEeOCYUq0fInB0K1OqYWNSPn8Z0j
uGjtqwd1C9ktr67OUhsfWpHMl7HQIi1BnUX4c+cuLGPql3PBGJsww6cmShJ5RDhN0fpH9IQfzCBe
17ibsChpsXCFPjOiTbCSU3Iot9bOau+lM9Ua+G/7CIaeYJksynYq5wnR6F70Hiz3VKgOQ7OxrSrw
H8VKLnjYFu38zFi0ZnuMlOi09czlKXxImNTLHaFVYxiCGnizVvWaAKW/wvRPCwZrPFVBQFnJklnM
XmC8yJe7yre/fBt3bPPdw11ou2YvKXQjcXDyUk4wnuZqUxFvQTdU07auzNNFKgAvabbalZk9cGIu
43FXEJQvoYqIyEdBukw+Alq4JVWf81LshenL1gFW1pAoeb3BktrnVuislMXLwpdC1UG+M0XJgLF7
od2Mkyvhf0ZfR/9U210LxzYhWhymM3gYjpYI7yOYpJGAmnCV5RVIDUpifPpA52vCR4Ue8RtPQfzs
eyHsGaxh5UO6EASGDO/RZrlSY5qf6KYoxDItHeWkYlTpilRGePSU34Ce14x0hdq36x/+6K7/eOmX
QjLFX45pSiQRCQW7LbYmL19DtG2FFnvpFXZFoYUeg/uOk4V5Vnj57BI+y+8QmG/26m/XLwHjiCaP
J74H0+aJDOld9TSV/NZZBO3dLwLPGaR2cPBHBHHwcm1S1YGMC7FEI+i4RslvpSUFbIWSGiasSHGb
YTxMcOIVrReOYJ9BPNxYfIcqrjffpoeHSiR0LORxH8ZBWt3dIfAb31VzagxMe5riY4sP5d3X2DVj
UP/wrDZDY78JXalDWKtNHlGWnX6zH/vyI/GaLznmhkfl1/PvySeKA8vg8Ufgzx1Gmb6iR/3udrbp
GOQOiag98ncQN+zRcru/hsTGx0y8IPW0XTI4Gi6e2EsCSlHZkISLfRPZ5ipdYEvHuO/tRgsJ74tj
eG7ALgoxTT8tmfiYhQPuXGVapXAPUUwzbXYBTp1GVMvNgyB0hM4i/Wj6qwdI/pPrVVdD1rBJt69c
teRfZwcjRBxiOWUSKWiljtnK9snKlaOA6YAVDLAWXF1/gNjWb3M4WC4wvaCHnyhSwPyGWc7Yxok/
fApmnB3hNvwkZaSve3l+DG9kUKEwmrsJf8bbwyviijBvXKrGWxJ8xGozTf8ljEhFfEIHjAEML74p
43RytvYhEbvwVrnnhNhhqCIojgQe3TSrnTRWwcHbdU3pnuyJnuZ8Ig1vRnJb6Arkpv/7+PhEwqBy
6sfrbp+dPLKmYNuXmGReM8GVciiFcT9YQT2rOFlpcZuK800aV8FufwzwO6AGOY7LXfnB+FPQOxas
VFQgiNRq7nCtPZ0JWMfw2738wNYTteBC38S5/RTADh6pMMj8IZx7Z342cDtFspS63+A5Em07DJL6
LWv+AmNGFeOqX66VsBlSy1Y5Ce/9O9DKPN8D8LBVnJaZChbghg5HSTlnupvzOwduJlr46xLBI+7z
TpKoAlpQ9CSDyHbxhMS/18dLUw9/7/+SoCgqvtJZ3vBKhWJ+B4mdeQFiaKxxg+qBx+6ylJDkIXyt
SDHMu1hUitKFTeo/KRk7T0ODqgdUXHYbjcaVyOgasoLMxeRcCd1jeBctNUxzNHLEFsTKBFO3XQsB
0J+422pLIqu0KSSOsBMHNn2YxwAjnI6wcSn8SHfyNBWoQW0CkNLe54j3qPvbOKfrOREf8PENR9C/
v/u3zn4Edc94HMGWAUgt+ey5Ta1SnS+B0FBzyTI83DTlVyQCTbVQhvnE4cArTVnXiqq/mX9B1/xX
77dcFfL4DuNirSlID0P7e083GTCwem36shKeWaMKkBpjEBwSAuPlH3AT29khbeNWsrHsQBw3tnIl
RW/kjLZO370VPSTmoSlSnAS1dMMxWs4d39ZYxBWsRjqQubasu6XKQtPpC1B94dT8Uqvb2aaaIIaq
HGDNAkBGjbcHZPzHcW4CbwQ8vTDprvTd2VOgVgaXoGQB0soxDJxG3gS5zl5e7iiL9ILlXcnbV5w6
Iuqta9VzT/Tb9D4ENrrOoqdQTNk9cxNvCWCi0iRnisHDflBrlx6DTVTFyKeIIlXFbQI++m2W8h33
EwZYpoVW0zhjPfj+uOYkiSsTHfjulo7hjNuJs5QiFcHdwHpQ6YwieiUKZUdn9tFFBAPI4PLC5w9Z
EJkbctPL9Bu+QkDkUbw8yLHT/a3a02izmndObPl10/5E2aMm4PEqRG/oS/nCCG+A5wH0cz7e0XGs
FuhUKRi0qOPN7cZJQBSlzambmHiw09KAAOOn48F/0JhU6NRDBoJx8j0g8AJd3sDzQdVCZlhZspyz
ppr7C7zGVhXVK9mbU3UFrjt5rrmz/S6u6Frh3h/ADehFMHRZpfqCOr543+5Zuqe0x78eYQ3Xh/fK
kf3NxhMUVamG1j5WSbGGXYSEfZTGqhjT0+SKYpSv+uAQYiMKC/UYWydOSxNGkubA5txPgAIJV1Ki
P4P74PtWafw6JT+xYe9ArhcT3s22vi4C/q1RQnL/FE8DHMYwC3RhjmSDvqO+7rEv0z3AHWunXx9T
8mMpwm8L3AzI6+78xsAoGrMgjepkR2U6TGxBik3CXwhO+JFrzMbZM1Dp+2hLGWya0LX+G1G1YWHN
bwcnlnXbz4n3zuvoQaYQFeur00bjLCcDL5+jbIONegew0K50LVYYHhYLW0SSeStXMqp8N+30w+ZO
C3r9Z9CKz5uq7nCpnj8JsppD3jObXQmqUej4ojLqUcaB/GV0NuU6lsxTfgiTDIHQzMHVPK2qfHbU
T+u6Q65QI+zTW7ktBqyhFUZX5UCLvdmipF8FnMha93PGqraQeo0BeBTZZgq0iOAKfnQ9JEtByvWp
m0ssdbbN03WGX4aTXYoAvBgnHXedxUm3fS/3aojDMZtJ0nYAfcqzlokukmWLi1V35JBUTkcpCfcz
7+hqEwz8bxDr31AAxlFmzmlRg+K/C/RdvOT1UHIJ9I5ULHsqnwT9bqK3aGPlbNmz7wveXDWSMts4
hV7UdtppEJhtn4rS2VHvcyU/gtmPmRkGWoAZaRYWmPK3fkdXUVhsDawMLHgWTI2+676xJMK/ARDm
avpd/UiE0hI5QptnUEqniP/qxg2c2H8KB0YlBohB3DbtVBdcMY4XPyFPAO6UwcZpngZfas0FIAYN
kSuDHRWnN1vn8GwOSIi5B80xn/NR3z+rYatDEYcdvApws+g6pnjT3f1QqXnsIPkWA+EJ2hjUGAgv
w7JBVSZF3uXeGOo4qU5X+fNN2f9ZPWIS2WNniSfnjGKy9oiCHCtXg36cAea6fcJGeY2Achy8KkO/
/CKpxnEat0Tg78H+NS5HegOJeCvy8eUwwc+SY4lsmbEugrwmUyrJ22PpuyHS5/OeV2nC4NimKUHT
KUs3IeJJ4EjTcBt1AW5GbCuKL2YR3Hg7Irvg1NnCUbPo1qgKokG1ACdCv7mbn7uo4GiFQAOPTHHC
dM7/Th8LR/0uTPilF4jxg73yJi205H/FyFAQeCj2ZD56ZUNEJJHqaKIblA3ZJuXoz/NibEqEeuM8
F0uBjRojxgfmMOP+3RmaoRiZR+W19HjMdgJWdTm5QGrpl8OtSNz5zxYN52ZedoMZcaSM3Gf1ZtKi
H8akzscdZk3nN/uF0f1PpBnl60XuTLpAdLcJTvCR596R0u1bgcy07YRMI1sUyyAW0Qtv67qHbfa7
4KZntYJB396df4hDwO33x12LAd3uR8ofgFEGyi0UtozIcgrjhwJUM1Yrr5b46z+aDzUhp+cCJ1FS
+s+QO8O9otyc2vIgm1YWDDz4G6Ti0VRlvY9vdLov4Qd0svHoBSYVHDPie1N5NtfAfKl/yfQWHgoW
ZrK+1Z8cSmDyHbj4OlXqmQf4dpFYMrN25XFS4QUh6WL4BDNNKXZSLwPHq4KtfKUuYUk4I3p+Q2W0
Un8/9tdwUnaOvuCbNjrOObgsfCq12ksn8/7N9cK3aHzRBhVBKC0rXxyQaMCZtGhnWepBwl+kI7jx
TmQBo/fjixuOABweR1XhaxI4Jf/nRSLT+L4mwXNhUQqnlzxxqNUigTMcU0NlBGsgemo3jy7UCFFz
hGqpnLczNqj8zrv6GY3A977NysDw5mqq/PDYfGXwRHtzM67MXoVleGMgt5ys9z+1qp05UKiCZ4W5
cDMWprYUc8CBHrulWd/Ws5kifhFSmrIQvURJDxj0fuzlurUzOVtdtRf3UJco68So/cUa1C7v7JmP
ATpkHf6ksxSx0x9CWg/uE03m1CANFI0xTU07Ayb1Hyjl1SubnpLArvT18WyvD8jRywKNfj9hK7QJ
ow0ArygvBQS/DGl7SIYAHka50FesFmPks42rEhjRP077HvO0+UHqV94oOHlOsusRzeULodQIVU7v
uhBgPTM6my1WrbXJbkWwOWbYx4D7JsDbGiqJGoNa8qCgONXzwyC7Q4swKUWwhAji5IHTeibmdORF
rsoNTaJCAGDHKgKcSRtJiLrcMQnUEcFDqcj2eQiXxkcr5Ah7zLb4Vh0ImmBlhF+vnc+Sp5LP2BO0
xqcFS6C/d+rGJsUZSb0kp0EEnEI7K5cqUISU9yUtaLMNmuU6wZ2W9dvah+LR+oOcpsyzUm0nXWp+
C17+fwh2TAEONjBObeA6QglRzBDdcBLXClVgv9EVEjfg6Fooy8Xi9bEPN7v03eLp370/vGxDii4k
dOBBaine6IzJvTo26qQH3RRdt5ZGid+1uRYlMZ4uwb0WHr3hGeEbqmmhcwZV3cw2xUFOD6993RIr
GleeKXioLNwo7y/aqZcYSwcpBTXsd7kfXSRh8+QQzO3TxCCwbWO7LJQKxuSGIWlcUhnCVKZKX96n
mDZWUXdQizCCQn7BeNd8+9QW9n7IT16Q8jcCJc+7NAbupLwXEi0p4m4iT3ZmpY3IU0t41Yifj3ZY
CizXBfdd5sRDDPiYAkITq6qnTkjEYmkH99oozNXn1trJknr2VK2LUPTNveUEiNXLMTg1MP+45Xt2
lreZfgzlYJktAN+X0AJ4FfM1jZC8AfQuS7B5yJcf3MRAcdCuhAhaCaPkl/13Iuwts8y24UURxjZy
qq+cAE8OHfcIuTmvq5jRPXap+6/1nGH7wv9XD4HR8wU8GxGaKmSeC2XSDRT+xoyseFdVuZIPy7As
ryBPZyNZ+XxeCPs3LMZngg7mcKrfGeurUXJ3+F+noWxfRwkyDinwJJSf3ymiAdv7S+ytKJSBp3wm
cl+SzfEk35vEQ/qlkNEt+CnoqNd37CDd7o9w5YCmPGAOn8VB8Z/Z/kWMlceir6JoDw6q1glHjLm9
2yqyO+Zw+Nl+V6kefEefLlrhq8E+gmXQDzNp6ve9G2uJFI0o4ux9ggGKXF5eWOSHBj1zVwB6YMK1
YWZm7tR/4u10Mxg4wVJ3kUZGEDQDNn6Y59S7RKhuLw/oK4cCkREa/02wvjKKvyT/TXuuObLph0qz
ddeZBwkqvJ0fSq5S36JSoMiu7oee9zEnmKsujIlvtB+mm//+/CauZRYo20wMvkZ1siqH0ROyE2IT
P7196DJ7Imwl101yX8NUcq81PkGm2bjlYINrknp+rluds7pOkyxKlmQvsP7CfDzcRPN6E5KEBu/O
tE4WdVCFbWw9XqPPFG8cemrkIX3QTA0d1FIvUNKoMOAcvgKjscpBK+9kfpsgL8qnRut9YtdsHPZI
2ahxStWOAQerC+POEwEiA0qJ03WzDfzuMFEPWjaON1IOrsBNXlxzy+nEwJ8pMBz+eJ/OMYnzBFVj
aNXUT6f4Q5YlNWc0k1ZxgG/PSs1Z+YcyVAnbjxmHGWbeOn7IRAUqlyeZRZbwo97vZQZXkF/YEh1n
IpAERqx5g4fLsoNiIyiNMnwrQW7cjuIvdnKItcFTPP7NI8Qlj+6TGK5iK2V3+g2pDO8qiQVe+tSG
97M6b/mt56HsZF/sj/WNetfbNN+OVPc6ypLO1+3dvxRJMim0SY+1WM0hZXgkuHfNbbsj9cnErZZE
T1gJytpbt+W96UGikf2rBK9vIvuJXqNWeJG643qAm3E6F5Sp4QS8KgFz2HiRvPJfZlxrldAhOPqk
up/5wKx5DCJDhxCccLNlRasfqsWnpdA04/Incdy4gPYOssmFE+lW2IPHsMXsMPwoI5P8dkjxVUMg
iLd/Xnv18naKJb8EczcTsFU5tlUbI7H6TM3lYyd0oQqdR1XQ8nCM6KneyXwgJFemXUBWZ3gG+sMK
kXzkut6jr+VsH7boWoCIOzp3wcOb7ew8mOpOsvS/ufgQWMSK4l8S37G/+4JyozjoZiqqCSMXpIMm
k7x9jXgznw6fYU74f+sL2b9ff/wEyqUprNrJfMQZNZ/3FP503QhIkD5gHOn+onE92zCXTPF1f9e1
3/TA0JgA7Lg2Mde9NvXFeB00L+jLwhmAqu9sVrgVlxUYPPBIuQ31FtltwIoL4UcZc3Rw9sBLQw5Y
QY91V2O4o+HdpJeIT0ObYDVSR0pumJGEJWMQL9xTkVI+L6gXGphN0P93ZoSzPQcW6WEotzsbdKuG
Hq6inpyqMoSxMktjIOhrBiQqlH7p4EfOGqcjhYmhfeWUuShLv2mR+XAVrO/DqX0CxrlkbUahmmVB
/ER4bRaE2c8ZVTG3gjs7a+YZOIx/Zu3XwfhWMDjbzFSmME/49wdPPwW4rQOZoEZ6paNtVJvxX4Rg
IR2on0+j8x7qQXuUmfjwaYvAAiX0zZ0feUUD2mnFIgaHBKbFEN+5V5qfF08OGOogif0tz5EzXIs7
KGKFcYM2nwFvZqaanrn29Ke1IpHQKDCSwAGADY+Q6SqJcnVdGc6R6zrArvSy9L0+VHeoPpbtvjJh
cGPXTGVfxyqjAfupeyWIdSjSFPJcYc0E4R78MvP/7/XUNPynMGtcb/djWn7oxiYN+AlQ8+P6YB8M
4ANsVecxiiJ+0oQkCNx3yv8mLYv4UXC6zHRX1T8YC3FBhp4841GeD9V9dH6YQ50pf0xkqc04Ke0z
EeF5bjSGcIhkt/aoaEXJ3NHWFEDBCOyPbBXx1s9cVL3qMT9NmfDE/3f6B6LxOpwsVcnUxodgG9Ps
j5z5kg5LX8EYiQUAJrZOVwGHVl/f7t9pgQAsO1CTcmiIBOuAbu63SmypFVc0eiPExZK8pi4KJ5q+
njNK4dq0vWXMRT3Dm5QGi6Ny6l/VsOzZtvFmgv0tLXNcD/m5D0ogzRo6SpWaFfkn25YdBIvAoA4R
M5nPZwnDpNWu/zTD0c20+E52WafVNXub4XcFDqwp1gqNBCeBWbsYhvxkanwOJZaQzLzcl9V0+tT0
YsxvXa3nAi5L3thasjzo/XqpEQ3VTMbjuak9vWkN7dsjHQGpZiWL4ENefM+H+/o13T22cnc1UkZO
33WaRgB4Y2BWfzuRV3qskIftNPT3cDC645QfuXM8RVMHPnsN48ht27g07G2HZKEDHhoXL2RaP4vv
GxyVxj7acVmbvDQWzkjwiBbx7Rwc0iHEuJEG2RnvbtPBLBCvlre71nRGHtMePtun2xcwHqlfd1LX
lMCg352vHt0/s1tVMmHTJrGPDlfjZJmr02Rz/zDX13QfbNOTsXb5LW1yMunc21WIY1cb0Hmgi/TP
5NKKOk8Ur1H8bkoKkH0049S5KiQqLfI7DE9TXZ0OwDOG2vCVkjEjFvlr5MX5vlL7YZah4LIuaWuJ
7bOU4I5E4D4XxAUVwW7FsBh+SWYsi97lFluNKaXUb6dGdeqKqwh4SFBlFBMbVQSRjM1D4XE0/bwF
ecwSEnhKC/Sy2X9EY2BjLZdfAcqG9B1MPJNASxmrvtwiEOg/MZWMV+uHApEJkvj2yZh9v/RPM9oO
VweOcpDgD8Oz56m0122dDXtPZ8TXAlwzacQFxE4QnQubFOgDriZH3CIpbESwftZsWdOvy2JIG+8E
W8eNumD72x/VknSXc1wabqi4DtgtngnoYD8sD7UGh7CmKiRkv2+sfN+uV4am6z87dYjACBK/S+FI
Bf5LFwo8fkly22Ms9CkeJbDn8VGENS4SNMbCsdQn3yxXIPCShiunUuCSbG7t2McLyfoU4i2bUEzr
ag8QaGUJsticjvYpfno/xJOINi4mHWGhV+uybvcT8Gza8+nNFUcH7gG1Sm4XBcGsoRu68eewRSw3
0LEuW4wzdVYLY3dU25fj0YDj/DSPLYdELg/2wfNPaa9Vq+qv1QWd3unr59ZQrKlbGPl9ntmXscJd
jyQTEeJeMShvGlYOzK6PBKrLjGqwav6oiaA8PRo6cACJ1l+SieFzvUtfpNq/2XJ2xD8HFe0/k+64
/leqDZA0dUvEpPApObwEBGWO8bZJs+NZaEvHWeo/7uzAQb1p9LgwJC4sQBx++7K9/hy5PA/SIfzg
g91XHzL6UILiGWlx5JSrB9PHogQLnk9CTuS8dj94myhKnR2QdNOlklxIYFJHwxduTluMVxktz2ta
vOkARJayRTFvJ+YT0IUE6oci3ks9P/ssOvjcP9OE/tmbbXlXfJUkaNpwR0L+eEc8yibghy4fN2/8
NlbHFqLcDYW4jysEvLw7FBAtMOBRXVl2/GHskKtimE0VjEvkT/w61ALT6yu8oRqjvNzcytjieP2S
I1lDYTVSBK2DnhcGPn+yo9VFDp5tBqDAU5kc5jEAIshlx3kv0jybjaDoOigOjBIBT5xYaLHMg5xd
HWQvaV8qIOMTjsKKNyoS1+mUxdf6Cbmsx81UjjBiaYSeSLTzShziKJaWjuH8HRAb+E4P5w6tBX2j
XleNEmWv8Lt9IcLL6JqoyXC1ZSfof0+EyB5FiUKzP1oBKS2Qz2TrRFJSAg0SEKFxkRujbJpd3rhL
+SIMgLBhnHmlIbAAQLtJSWu8tbg8yXOTO2lDzZyuz4LzVzyg90dxRfcGxDMthVIkVBxr+STWiaj/
uDuqXhCI6QVmEN3U8q0HgdnLkshk5Ptl7retyIJVRLEe2i/6//8U7n89LMqc2Qo22slAKKzL98WQ
j7GfGc9sZdqHG8AmzlVI5bIfOC/hq6GtSN2HBl93P7AzdLkfoNvR1u7lxTbLxOk5IDUxeNZ5bqpS
Ni/M1NHHJd2SbYnCsuDBxflmRm3uRY5eVTuErom/K9ulCKqBrsV4dLQr0MzHMo1d1jOhYadMIzWH
srSeI0qRkOzV27RDKqBla2HCDObOtBCsdgni2cN8BmPSV6JuK/LysB2PE4112mLqkSP/IEJMW4Cz
NMeYAczAzFwjIdlRWPXcdbrNyvYtFENE5HY2DPMwWnWW1KYqeor/YLX6rWwm17ZGAbP6WM/8OLpw
4Q2qp0grVpnO9Py5WFOqq4DWggkWpqy6mnFomNbErJ/MHq0eyyX+gFFNMD87KKGzQ1vw67jRvwbv
NVVBox80KW7ZnkY9fgO9qq33bRGNa/rJUDFrMoB6pFuIyyuTb8RZ+CHLYkbF929vpDUVXn412auf
uiLJl5XFrgAYhip8E1I12/ODT/89G/6m/u1NOHE9DPuDUu4GfRoW4kDh2nk1216gpT+rYjzdnTpi
UvYo0fLilE9MFFFTkBqh2BQVnb8kuE40z3HG+ozFVhCq8IP9gz0RelUuDzT4Zw2h0/zcie0oFK2k
2PkJOv4/K355BSjUwfTDXBJnw5+fXsJOIqNybdPfnB6LpyP+DrwvSChtPRrlLELgCtBdbUvTtnT7
VIxAuPzk2J9t+cUse0GKVVOBiFmsW/BdnZ3to0k9Lwwfd3sgUm25ieqFQI0dskVaqMubkiEiVWi8
f69Hgevy6Ho+9eWy9Putm0DtV4loOWEjQj4RzNjwOlhEj3c6j3r+KPbHoEWrweO4bRFwQx/KbYOv
FDqsF504BYUIoo7+P2yfMuMkF7sG65W3pAS3hYQeuP3YOuTcdscWAXyN2DAeAEk/61KuRNmT2bee
1M7db51AeNZw9rhMUsyW1rUJQZs7Boylu5i81pHAzHM5b2PHAJrL6c4EmzyYNhMP2BePuiGxssl8
vuKsJ4t/ybhkR6wXW4hN3amHATLQexVmRZMpbqOuh7+54Y58+wnyFHdz42Z8WL2Sp05Ffi9nmIZh
o7b62cARSqnP8vtcyYUh1UfBe4bQ4P+7bAUoL4xmOfMTmyeg2ae0tkD4Z2UJMOGOs6yu6EelRxre
Axqd69Bo1h5iGbGDfl1bcdCCfwp8AXFixf4KtAC8tKbwJfe4hSSrh9gk6Igvk+WChOsSwJsSoCDa
BylFMkyZV42oa2RLrjAjnQwCoqwTfmUsx+tRpqeXYDoFPsLDJkMIJ3qqeUlnbNPkJBQssRp//DBD
PVOCUKla7zce0n9+scif6zDpg53jTlTc1TZuhSlSaF38mX6ZnqAoWAmt0xkYZje7pV+aBE/gtYWd
4Is0IQ4jOM6mp8/89Omru7t7DibnP7nCvSdZpczWiytxoo0we00l9FmOf77syQKjZ3IuwzpZw81P
IYUfKB5TV9+XI075koLJcOBkwchGzp9Vy88kG5LmEqAXqMgxSrQJAQdndN0z9wp/yQUywrxUnfVc
i2xLyRCFquqa4kx9/gek+QSTYQjNZtryDjaw8O6sywspeS3BpmZQ6GOhITSBNEIxgkvO/awS4RKo
CQW1jClnkfKeRdhF5C05atSMDEvy/+c1RmCL0ktSwQtVuMU6wKgC7jjt+QKc9Xnq2Hx2sVM/G8rq
q4/BCZ2WspwzHW2XZAd8oTp7ngRmyVoSKtATAiCfR8HOKu8rCc0yJxoq/tMwNdbJtD8EasgpNsSd
h/LP6aL4PlkY4d7wa7+IXZjE9LKa9DN/EzL7xsA0tcmj1fSCM+1p8CItjB6cNto/DaJBao+09/oU
d9hBHEbSpzN64UROwXDeA0FqNtvcoMoJO6oO4C0J+dhYISwl6lqrxJZT0WTvkP0nxZkCpdZy3YZp
ZfQEcHeyCVpQ8AaszDuAe/cK4DAZIbJOybQsfQJaB/e3ydRlOdK0aRx1h7c5yuVmChQ3Kh3OxCNZ
B9CJQ2v9dXda3dB78ysX74HpBlvxUffm+l06QRqZNO+PvDh3KIInHPakkKH5rhqa6llFpdmh77Gq
RW7QvFxybYvMfMej4K1CECMYb9eo89FjuTSGnzfAxR3y1Mjt6EitzxkRfIN0Oe4no+epzY0M3m89
5Q354SKmg++MnCuy57yezjDBL++XbwWfCDaxd6V0Bxg10502DeYqLpr4xWjiNxxvLUWJ7MBh0fco
Kpz78/ICb4PzA+uj0UOc9CRLd7eO2eT7h0OpGaFA0TI3+Lc8/NQLWcrcsqzgfrutRXOnkk2C1467
mzJpAso70UcoP7asFC9kD9ZRiOz9uEsAs5NpHgNIPwlHHOb8zURMaHYtRJ45YlXnBBF609DNuQ7a
ln2XnlPIFXwoLGEKBbJ//X9ARgTgy+FsttizHGnzqZb5ywl/gBow7KDRkbAeLrkG8zWWy0fOoo7i
F6kg3IuEUUa6OmbQuDMAhvANvsSaDe+ew8OQogbdSZzOppbmMi1HLWId/VcW6Ayw0hv/vU7yjR/q
oiQ1ZCmr4nU4ALiPMM/837rP98r9DE4AnjDJuUM4nNcSR9jpb/xaFHhefd/zjUV/QunHJlm9bduP
Xnv+xayg6TKOyC1/vA+SUxDeuqn8Jdb+OnlzRCldAWTiiEzEwEXM6bqtAVA/BaBnbCA8TbkIAOsi
L3BicC/qBcJcF+6D0x1rmb20KBLaIQ4QG812iIHK69w/cZQPsBrfQc2zQtKyejpfy1EPMEGw4bEK
AcfoR9sJGqCbNxd4IeB0F8X77XR1AwNqcAY7cAM1bsaLAiiTU525UcFH7UB1bMBoFUgJjS7Q7xgB
yWoM/QffXCNhmNLMCPMk7tGRAVX8RZmwEE5BJkKqRaqLdYigPbuK+6Mw1AGPkqfIFt7GGS3jnDEi
hMzVedRBGP7YmvflbQQ3x270sqOHqME5p0GwWT1Dtu2lN0RgJrxTCkZHWAAbgR7qWinQ/wGaUWdq
ik1UJ+pzWfe27qHdR0wsZT8krHWQpy9yodUgafTo3LGH6MOeN+Iqt62nRRAdHtx2b8GtB7ToiKGu
9GxlNkMK0f7nIU7Bd5H1zo9w2M/oSq3hijdkKOv5DNGiNBcGMqXCotaA0PXlCJqqEGdn4XFZ8wrt
PRMmX+tbIvvQk+H9OId2hBugGCG7mhw35TcVWlbaG9LN0ilHgtj8Ys9yaLV/Aaz7ohPc8xzt6NeE
57TMtiBIOEzl1zih+eBBLgrxfbsGq81R+duatTh01jtpFy3VCkynnUPxdY4gQfQDDH0FwjmAPuiU
AVOw0BE+jeWCKVx7/ftSQC4+CB3s0vyPJwuW0uOhqhboO8+3nY1rg/w+N5Kv6gBBzvD0D55l/dAh
SCfeTmJtHicJnHOCDcht6396k2QcFn7/uuxdEdYdyacd+e7yoHu1Xh4L2K63uq5rKykfqgmjX44Q
76JU2hQJ1VbI+O07ZPOAqLslP7mL/0nyxtBtwssYLkthBPX9/fO/k8QLhRs+yIhfVlHIZT0J3a5Y
00DGJiZZfOQbUKxd5GxXyXQJTyU2PVWyS79/5jvvir+9KxBSu9DlzN0pk7IOt7pKmtwiKuq07INH
otSFFJe8JiFKL3tVVdTuEfDbDOrLTy5eG7M6oHmIkrwwU7wGy3Iyf6zd292AEa2OA7iF2aSsXc9G
AVEhOzIilvlEMPiBdF5F3vKn2KkFp6S0QU61Ad/VW+Evl0XqsC9faqnqfCl5JCfVZ1mxych8ChN+
REzPqBELLUxJZJxMvv39Onx8tqmbm1YoPDSVgwqsNcZNKjdAhU8BUNGRPmk3SC87x0oMXK3D1AQB
6eR02H7YXoFZ/ih65HjTBiQalb2afmHf0t80BSqT5simzKvCghx+K1ZBwO+x69wBwhirXAEr4V/u
PqJ7g4gy0ofmMQf9fjsQ7uaKs4U8Nlz6xhCybibYvDwScJ7Pvdy5dQR7mY+U4an2u4PDjn3Bvulx
hV3+PAtw0V1DP26R5wgCuEkXYgf38YWs11PcHDhJNxpV3SwSb1bG49SkVC1GN6nZ/ZFbOu+eHY6n
9w1r1UH1/TEuwN3Y2o8D08qV0k+QBdfzGlS2TJ6jHtYvy2+wwoewxf3jEl2Fc/aVNbykIYmhy2f7
s5oEvtgFUWEa2i3f0PplAGYAwr5kiXxHG24It3ExcFVej9i6tk9MTKY2p/Z1J9DM44tyQQUdnbUK
M4x5pd708VfbLmPPpPQFs98pl0J4RPxh6pIAILLMvGkvP1eTDxepMtQ60WqmL04s9c8JILEKmmTD
D3vj5HarlrEuQ3LkfD0TBdkDNl/XnPdrYj+N1iKIlqaZHUI16bbwOZ9iqylBhsS4w1E8JyAfscGa
gEdT6XpcPBuDL8s7E+nc6o8sEst5uYujpLqvL+c1cprF1Up8UKjjb/ZAMLH1twrkNIbBuc7If8sy
DvLCu6R9MgHJWGXpR1HtzwB2AmyZeyXo8NjlyqHA3iusZLyGP/lNbDoHmOMDgIhqfiIzYcTCuB9S
cBKEB6sToYHaXPAWGfOLBOPIFXtiXTWUe5p+ftniHYGddB55ytSTE+kP4n0MSPzVHJfDOZhAtYBI
JFb3KPetR7CFhh34p1BiLB2CO1spAFviMOVVz8zn3J8YjIHdcau8f1Na7gqjptxi0UHSV5E9OUui
ElAUv7Eky14xoVqfN8NJnCV9V0Zmrs3gfy65j8JQRd36sonOEfg2Bger1VnbTbFTuRDW5FKa6t5l
q64vxDbWwki7WVpSOx2YCyzDTPgKZwqiqZIfspm9T89N9YIou/ISYXxS0iKTFdPBJjivfTEsYXIy
ncH6bmiSWS2PXKd5xbLwWoO7QfxEwofTRne4Y4E0PmZCh/+8V3XOvOd3P3ipQRhPMFV1niWmrYiE
u6x2/kJXUGTiEQZnooAHg6XHHPFdojAMhSLTHVJH1t8WOoOP5M4IRsBtpeQ7EDWIn3RKJrB4f9oe
BEjlAFT/nzRbETjAM9ekWCftf5BfxpEa8qqZkPO/JbcctseFv6dhyrRQHqUcdDv9AFAI/f8UCnL9
tm7NZIYMrNFk7UDzS7ulUAiqcqINZ8ymk4M6oP1kB/WfIsU1qYXeUMpoRlnY03dSVoSIhgZArqrI
YEJQtD9Ofyr4BrvezQmA6W3/JWkylF0m7D3cv10WYln7/PXMeyqsQIJcS2/VBvSnUKMZk631lto9
3DauU144tNpMUpR9ZqorS7Hb0tVkTMqn+d+Afjx2kHO02Ii+qiwVEipARzuYIbXmPFMW8EOqLtc/
hUA/kUHeyj6VBHDjIvTzDPeM49H4ACc2686O2uLH7q1PPBASpDEzXMJtfE5MCG+mVCYTp9dnfhki
QvRRTjTOXrtjBuLAimwKhWf6ANq03uYpvoUQXVMOTWbepP1pFLlUM+OEFr9Cy9oH/QLPleI3CON8
4CwGh76AAPjCHYx23pGhkA+hr57E23v5RvVEu1Uwyv2Y4nXO9DikME31hsYF35+AQIT6J/W9O/r0
2plHN7kBwB9lWwHGyiJ2OMQwFHNL6DLniGBgcMDgLw3wJuPcW/RJZLYSKbQOqLz/XLhyfki8JKHm
WthGfRfFXv/t4iAIkgv5lCLCcF2+Of0e9S/T48tvwEWmq+3e3GGdzVcEpjgfC+MosYA3ECT6hKq3
0VW2Vcd6qWn/wEPB1FP0TEDBVMBQ30mkhJKYZ+5io2NkglwjLk5ItTMdSDm8wee8oRpiD2u85jWD
C8njmvb+lbFvYH80siWstPkUOj6b3rBl2Hu+jvN9VotR4zlP4GOs7O3FFr4N/t6VOHiPz9aC8rrh
AnuifLsneTN3gbZhWQtgUHInPSQekVRmoMXpXFbHbnodqeDViVC6SlSltJsZKxfOLH0bRI+JnNzO
ejd16cECvWc/V58SCq1IFU/cUfuDeyF2iCm6QNrPaCR/jqAcmG9MST1lA1Cp22yBCjlJvMEYomhR
ZOITFW2bFPvxIEsV7aX63RIAhv6xOH0N7OL9UNoYwq3sdq6BPqtLGzCs6EJ8kaYm3Gew0CyYGg4Y
YWYEyH/8g08W0Vq582syPFABZ83wkApBecZssKuX9pL9QkWZ1o2REuqDIu3FQ56KDfqkRvdn58zk
21pFCRILoXrwP6GEj47Ef3Tgni23ZDGsZI4xNc8P8KeBSYZiEnLMyu3EopDLy7KYWKj/HecKPOfj
gzI+GxGGM20XDizGrCIeWYTQI7d/kA4DOXyvpN6vdfamO6Vp7tOPAjMQ8CWi/RprVTlPH4NqDdwP
fKzeWFE+gRQQfnz5Hh8NkJB5pBxevm2oxnAKVYKjVxeJB7/NQSzIhI87bZ9DYlILcwCtrc/Wd93N
UnArqefg7lNe4pAZM3kdaiFPuWsRQ2apv5ufZ7/BslAuUiGoCYZJdmMye+QYalTAsrrxz6ImyTMZ
36u7Z7Qf+Z8I6JWH3BMuC82mMjwAu6ldOTrKwSvII2Uf02kVrouTJ4o8YtVccYrDGc9gs09cxGko
Kwlm2A7HHdOY+RJ82BVq4dWipqsHxR/rpqIwyjz9uY6fyE6TUqGE3/id8m8fqbbOnrx1vXi6t4NL
D3nLDo7zc19Pib2MW+Wkm2Bfb/EVzUcIKxskiDxPB7+u5VU/UKDZWHJL3/bIgP115U2IJnWUfqyd
b7er/3jZsHbB3wIKHgZpEkEPsJUIZzitrbcip7rb1STYzfm4jVi+tAEj4MnDbGon5rCAdATPL9/W
imB24djR7Ho70qI31Fxn2u5sd+thgSAKnnU8E3VZq9hRrclcuoReHLHJWUCtG0sTutcPhWBEFST6
LMa5lSFWtNIB8pJnYiBetjQhA553KVfHWle+zWuiu090+4WHcXBwFdKMtB1rmG2hyrDt7Q2DL0Wj
0tnCuZRKRhGR5+kDt/Hv4k3X5zF1ftHpVdzxUEl4ssZFFI6533x3nY40MPISJ3HndQs/HogHpsxJ
ebenpt3PRgbfsrKHqpDpepFG8SnfxgqTayKLaCpz+ys3Bc0hPVBIRt/s/+mwC1o8PKQlrE0skDSt
7ay6LMJRC+RY5eDI8KCXFWRaZicO0lQE/DmnxGxiDQSjnQ49Ctl0pwcdmPyvDGFEnGdGi6oY/vfC
mFN6lW7si6oHlPtRB51qzT1u3UEXjMMoIEQDbydOncPHBon+vBdil8DP61LsT9CbmEnuBpbFbkm0
27knM3J6w95M9MjtE4urvMKxIRnmgKp6CAV4PEfBZEEAqi63doUJn4EKnvTLnYglQ2M+kmtm22zL
Ag90DWdT/O3A9a2oF3DD4zQEVCEKGhWKYqpNtyHhJcUySlA4LlU6NNDFRGW97kcSikV6MWaFS1oT
CAG7OJfzuUvBelwAiZovF11M0nXyDcRkrzRD/ivLHQLwzqWlyiplGF7/SiNkIsuNtPQI1RkvA+en
AhXUEWGz2mrh37aLYzVmhVI28GkmZ4iCiJgdR9XfqTYV3P7xv1UZsDVXO+ffbhkxIgR5y9hgyTBP
4rj0mgvIcUb/CbWezkcvyu8jmwC7LpBRfM5uem7FNI4ZkoE+p13/OR+wlNlNhQjovKrhm9QBknBF
UTvO8Js2pMEDMBO5f6+TcDRxyjJnSzgXw2VQ4uEfzVdarF9ya8uqsEw262xIcJ208X1+0YC2/rxH
eoul8tR7t9W0y5TcnEIotwJKX9mf+We/bmvmAog5m/UxqSJ3uA4P54cuusA57sEIh0excD7aINfE
NvhHNrK99V+mQTqm31rUPHTIjkpsvAs31TyrwwmosPZrvn3lsYas5otaIxAR9FNec0p9Zl647UZA
tpCh1kq7Ll4b5Y2Zj1umsQuLUsMuAmiTCX7pt7z7Du32V+NDZdK49+8zd3p4L3KTKAYUpiVUsCkM
JGN/HfLpyqgoKDv4whPrbppR0t/zzFbz2PqA58E0ChxcElSCX5+7agE5js2uKGQHuUm1du5BsBL6
Wm9fKSRuV9ZUu4y3CIQj16/HJ1+KNsos6rFz/jjrGeeokHjzvT1XOKKAD7JU9lG5/JwPOYqjonrA
f3nD+p9qhyjCXS2z0Ihjq83Prxr6rgCNGMXU6R1cPzRWtmt6pOG3HrKMoFu73g7Ggw33PH2eCiAY
6M/yZRx+WsGL/hZsIrryCkriZFC2qIfhChGeuBxC8Gp6vbMBys5uHrQMH1xRUrkj/1YEZkfL/qHC
KLuEXby3swEVdkG4BC9sdxk2QdFzSXQ9Eu/97tQhuPmAurHYszGcuGq61Z1EB0sJJJqygazfzup+
RdbKWtEbxcTv8ix4yswe2js5ru9UuuMTrNR1wwM0v4K+dGNXMPAKUbLvR2Dd0/bJnoQX+7eZs91X
WUuSSDkUEjzXanknNmNoNkCOuvZ0PUWC2Erq+EC+AVrjcjcRMtijq7uK5aGpZOB4okbJTjbDwBC+
B/3pgMN/nTMEUnxjK2MAVtCQLbAqeHnLrDRFZZjb9uMOQksXa1reu++oCYDoOF4RFNzJ8gfc1B6X
HRxwWnrpH9rXGRo5hnQVApfh2ynV9KBZgeChCckiKeRbKeJ8hYGAqkzyiVDHTmdrm373GbO4vPV4
dsg0crNKocG43T/x+Ez5Mj0YA5mMEn5kNXsDD+3usYcK2b25H7Y0GmcMLufw9Pko8m1RDdifjRBy
0+MmAkxPqdthk7dparGAVpUWA0C8/gF9Y8gbHw42KZWrCDnnjvGNBrEivQdw5g/4yf8kKunjkpxa
QVflpurZh9YWCYgajNsZlCgj1BZhkqeKsfuA3TgsUP0/t6e7mdDQX5cmpWlpeHd1aBJJBPAcDsAv
VKC2y1H3KtBMqy35hTdNYp2HcaRwNnHcCydUKTOriMplPwE3q55a67OT4jDeZYMvEmTz9QoaTOCo
WL7ZBXaHehwFP9/Zt61fM/PfGuUFPjyarkq2dePKHjzZBqnYbQElToNCC74+26HwxGHDEF/JsEZf
R+HLCCyIQYsalCgBe5wqKF4XmKMY0i3tGE90WVjfZ38qMXqqYnoF6ubuSxI5DWMMMZ+RNKtm5kgc
3nD+c9HrPUk/Jc45LL3LOu+5TBrg7zrib6HljCUt9FthYm8xLO5C8uzIQ/mqiYgJXI+PTdq4W/yp
NTZLhPYNZ9QGnXFvHY0gK2RTtd5v0Qao5UI3zJGdEDpNn/Tqmf7CEAfd/hSLLB3DQAySOVWIythP
dSbi6yN+SbIZYotHw+UvFq2l6lp/31ttuaoUcycFszhy6WnH8Jg+cYMC2R2eTLN6oxvZEXMCfkoK
NdNcE3SmjsaOyEcWHeXtYQxmPz7os4CNaImYT8siJAnsLCJNOq1f9GjKbTkn5UO3pPvQWzKsbNE9
U7kDcJiRUmjCOof58/jRUNvMIQAOj40C1LqmxCPw3BQjC/ImNq4hwVF/EBqskUqHsAU4DRewJEqV
GywKr4RjLfbEh5w2vYupweXiFjd44QeY5m+Ocuk6i0lrh9kRZy1+vJkJbzsAFDMOHFEHbS1s1uB9
Y5/GAshAef1Rix1tezHcLaSW/nK7KQ8Wc9UHDWqs9QS+r7bb9rY13Ro0Y6sXR1T1k8TMYb2BJMyz
9P1oT1UJ/IwSVuryJWCU6cUkIC4ass86jYem8kzGy6q8Oxhdaqqgcss0Al7u3lFo07ggjuUEpwUN
ONnr1EkDw44j4DP0RkC8LIKhYDjGblebZARt8b9xdyCFVZ2SQR8c84ktEP0YJez0e1IMu7d7tqg+
SPZUMnzvQCqwozDpavRY5u7Jp9VxSaW9iBOCgiMZ6XG/jidbVM/L7nSH0lcPyZwei8RpaznjJmWd
h0k7HcACiG4eIN4yzAbXNz4PFPIwQI+jHfEMyiCNjoZjRdVF85cuYT0PVaVXiZM1c4cbsgOfJd3q
E64oyizoMXMlSjycdARvKe4qUUNZrY7BD0jIJvIRSwd+RixADUFwkcFjdJZmLw/6lCVnQP2HW4jx
wu/p+r9LYS1RqWWrbALlihtQ1BwHqJ0U3F1sB7k8KEIuzLppBVTMau1zWicTHv/j9bcspSrlPStR
4BKD0yiASPPjaLqc2karXj7JBTJyUY0xLw1B4Gmv5j59mFh7mQlB6sqt0uJzpmEdUsESIYrlm9TQ
/Rc460Ik0u4xNhWKeMeXXx7OqEtDg6KYwiZzqcFOznW713XlzCTvJZijkXu6Uy5abWGaFK/qM8uH
Xx9kMKJL65WAZ9aVigYfoPPUYMlTn9TXH68AwCNPJPzqkx8+jwzFVlvAb9JjZStyB5z+8nUVCuDX
5dZqmVLTVFRby94q81iSv/4fn2sHWnYutrgkejeloVJSPgQShLPfdMJmM9DOh7No9mzCHTRebQkp
O13BY+tiGRJc3Ir9MWzRBaCSk1IKCmhdAmo100B7eBBEZR20itdOKRUFUqaHEPoUSwgtqfriX10c
KAqELsMXDruv5fA52Ljgeyu0jxx/aimpEDpExiokjnaPHgbyq7OIS/h9YtKWaf13zqMROxQor8lU
UUv5ubl3JO1FrCjhU0Ls8AwPx5wtUa2hosWwlRkfN+dWoK5+YzcQBKO/45GP/hMD7ERaQZubBJ5Z
Q9D3tDEi5qIvOKd+ZVRjF5DbG9iFejTXj9hN+ltE9Fw2w+gFrwKt645iLNxYGZoBmB44Ml1BfF/m
kQKrop8xIwScG5pvZInzDF+IemjC+vchdzLDMkL2DJe5eMTbyanR215teW8PrykFv/ljOXHbhjQ2
SlYzcp0DmG7KKDs7+zf5p/jZuKoK5v3dAEWmomxi72d2E4VVlBHosT52iNBASAVHq40YjX5hNoCm
W0bC79Es2fQL9yRqlFbftJUxQzBD5Vo4JX5c20rqEzQP+4DlbLWI/8y3G06sILF//luqc2j1O8t8
qletoOsaUZvERd4MHMjYyCg7z5Z8tbWhkZF8Uey1v03WNO6KqAtRddLOAq4uIH2DLKWGOQDM/ccq
xvZIS+X5+s0eJ3Mh6FG01oxaH1qiZHT8wD+2CSnTq25X4nibiCjJG+cHYZijzCBiWuys7nkcx9Nw
qd+hhTCkhqdj2274w6nhpwd6gtIf3LIazs7j8zTuxlcG139R334Ztkgzy4eeAHQbK9+EcG3wrBxy
d6ml2pR2tNT9rKaiPM+lr+aG+JsCYYb6AQrBUuC+8An7SWnqV08a6CX8E/6Vra6Z7/8LS9YBfenl
93kY4iM0VWhtGpwFyI3Frp8P3BWfPpHIs7ig6Q08mo3Zk6JGvVKcmIqCLiNNfLnYegeo7Li1sqKe
wlVbUW8tUdkZiUJttq/S5Tdh1Jg7wYTwHN/I4g4/BKb6rHaJgg/Ux4jqNyy7IuhfgdOY490BQDKy
I2MCq3VRJJUG4KbWHLbcqcPnIthptAom2Fmlnmzpf+t3LnF16mfLjlifVxRa9NdEpT+mQ9xIJjSo
hgiSIrbIeHcZctFmrpFNLobYMPCOlHBW9BkEJDIXNEsJ67qTaNOVaZ4xKxjlbZICLKwgJUuI1k4n
Z+IzG7AzLErdC/dmHloTvrf+Y1G9bIqREby5mvF6tdd9v2N2/VGXH1CMRkArVqtk4F92EMsceM3T
8oECCDOycmOJrT/TlGr7wSkiV4hfAL/MODuVl/WObC/qN3l9iAPz9sQxNHmV2MP4YfsmdO3LZKPa
19GncEH85lvxlmg6EVJcqZ2sK7mnIGJVI8ZwKI69G4vetrtQ8Kw975iU/rZSF8636cqlFd50pE6X
oUsofW1iyJMVALvnOO5gkZD/xJ44sdyPklHnOwduTLYMOyffDOjHrvefg4Nb30F28gIO2V4D6VgN
eyQvlwPy9/vP4wffKF8hCYpznE0kRgjJEU1EC6bJUzPK99COz2f3t3Ux7EEQcn0sYzSOnX5yKN5F
HA1jLJG8fO5LBB3dXgLg4r/g38DeS1FYM5KtOY4XizsKsOZ2V4u39ZvkljwghGkhbfEK9ZunE6IR
C8lUZ/9INrCQs3+Ap01N9qVhmFznFelTNV192OegTk2TUx/8hbSwyHVFa9m0N1vnq3ExRz0DUMUu
R3eWq0rk9PLBjciVDW926DHNEVk3fbP8GRpj9MFrMZbrSzCLyjzMe5VnNWeXmc5pE+UTarHisPBy
ac4RUkDQsLvKY8bTID1m9NGEgF5p1BG6ptRDAJKHBPDj8lLGIyzKF9djA0FGQ8meh47f998WNc5T
9UEAoAfovwSn/vvE+MQFzOs4VfD8fChtfwuUiIWrc01WL6AFuQVf0W2XFNdjWpdM49ZLhONW4N/8
E/RUJhmGpIBkw1V3THdDQLCnAnrwTC2NLmsWUIHYr8+31MzJrne1+PtbIYQgjerYIIWfu4vZRqxl
Dy4GL36X68N5V7Xqmbfeua0iYjLfr2Y7pTcO5lxLEFPgTt9z2yT46QNZvhqYcWwIi9euP3U4qyIv
OrSjUO7Pw06cbQGFk6ikYX5CBlW7hzCNd1rF15KT5uFDiBDMIGzyMINvZSevEP8u4w8DAb2cTnl6
bA2rB8jkdKHQVIKlKsdCSOJF47peJJl4sQfoNtf+JxDUeXxq4ZmljfBnsezw0iOV08QsrlV3FOQQ
rkyw4A/Plv5NAAnVypHN3XQkdUMwp+WGYZ2owI0kuCodHzy4aQaFeOpL/nwDsne9D70mkmKYk6L8
OlIoQuNHWzfat0D7idV2Q9di5uiQmWFrxGocBzJyZyBS+frlOcU8QKUQgGaA47seYeXop5+rvegI
jh4Vx633EZtYumDhDvCIxBwMuCDPzkn3J1dxayo4wCf9+tkOXVYqJfwDnLsK1WahPFEonlYjO7HQ
OlsC5SOS1Os9j3E+WDLwuZy+wD8axMCP6CaQ+9K8hBeF6i2JdC2pMXKSlRn/8XeIspeSnvIkDr4E
v2q8DyqoNTa0xlBAKYrWEpy0GvAaB1AOREOesTNXvUnSweptbMYreDols32xcnvRHHLI7ch5F4ag
ZTRqa6JlUq6MD4AvjNim+kSR6Lb+Ixi50F91pWOCb2oAUqrjD6gEX05B+BaHzs8TjYI7nulBdYys
yb8A2573YVsK2ciWmYJnyIs2QCLpr3lOBkOxG23wB/DAmR+VyF8NS0eHRIGbLpW+XsRcMOSabopz
jNTkbojT6mLQD2z69H/axr33RzDOXK9D9Q9iAQmz9AN2MzJ632+MBTqP8pvp3eTjm1Ubx0T6NR5s
0IFmr53Zc3dNTNi+LXVCGJJ1RHqKRI2DYFPI/XbrcYnghcS/r3U7WE8ZbsQKd4kZ/1TG0j13I4QZ
VXCDF5kCdFQUS9eiVVYlrJwgqu2bLzmPWyzgNrw6ZqfB7oKdK4Q/8yNbuLdln29MCrimdassRzF2
aYzGQO7hJ1KGJxQudiWsZXfNlsZ5de0uI/gcDNLE28BoW+6VpsIfeXztt9zkXqTmTfUVfnkSEHZF
7+vq9d1om7ytUU/VN4X4Jh/e8MaKBhZYl8qNW372RANY6vwIsvx7CQ+h6fHKsJZ7MITNMpHnePjd
C5fB/iqOgFc7MrhwXAJ6V63WzdO0SnZfQs7TGWI3BtLg5bu0wY18wikmtO7E3HJuXu7Jn+sSWBP5
YT0OYwXoznpgHUfg+0C2tl95rMi1MxZM4QV2Ynf7K48brCHyKnFXPNUTISTjgwM+D+ME8qoI/T7f
XpWJ6A+hna085CEFpmPkuBpXwO8sBixUbYjhsj7VQ7YNW+ay9G4dQXY4Tx94oaepQgTKtiHSZo3w
KYbDcUlxqtD8/0JUG9g6e6MgBaIbtZmXsD1BwjB6+eq32WJxse+iVtLekeLJshM3mAeAkCFyNCPy
wZk2Cqde/BmCGb9zlZ1YYpzTvsgdg7AchnGFgxOy9ug4QLUW/73hwqY/39OPU/q9tHkHvE1Iswbb
lDKYx4quAMnYyORvlUxwkqtK5hojt6S+o5ZWCMPwn1ZurbmhM2204iO0Xme8GYryUbFCE7IY2Pvw
B1hzacH8/+PfvJOUemGZn5HWIxfVE7wUgzF8FK7t9k1dN7SNgM1gV30tKKwZ7dGkEbxLae1weJRY
YCE5KjkaVew1bhetbgFts+ky25da1WysQk2g8cS+xsrTOMaLrwBw2bhjog3ExLekSeWOILJL++as
NxxgdzwHRW52SPzHwNc4kLpw9l9OS3qpqpvQrDhyMdGpvOPIVWniBmbPBGk8gdxDPB3laHSW4lsT
/u31tnzFDJ8uLXb/xQamnW7nQPqttsQBFg/HX+Dv7A5arb7Pu67XmLjIzu5z6r59wuW2ZaPYCTE1
V2mc6XYotsh7cGOUGgWpZb9O4cC5FcK5/ivVgtQDnW7CFIHTE38EVFz3zBJZNr5axphV0yxI4iCl
e3CXPOKB3o6ragflCVaHpv1ffrJ3SjNChjgCfY91hNNCps7+IC4M9vPTwJLt0GxmggBE/kstHEH+
88aekVrdSwWIlR2+CgeT4K/MuvuBh8i9CKJiAJLe8LzAZ4Cgo8DRX0s6VCm/N7HIezApo++/AScH
mXSCVRSVIwejWDplmSm+4szorU3TH9+VV8lTxoNhQ7ziHtWgXoOrDsuFG1xNTs1WpzNq/Pnlnaiq
Z43VxjxCj/hZOPr5mncnhd8Dz0KkZPODKN1XUwrJS5jZxLKAOQOztxcHE3RXfKUzc1PQTpwwVFS+
Ur3Gcnd/J9ZJJwEpVXfMydFq7kMgVYER6IXZSuS7pQfNJSu5pt5WIdGXcvhEJTh46Ncz92mKX3zZ
t4Jz/SDZP9RbKaUX5ERlMIxiqlqCwrMjjHQDRuZOJDv+SWcs9l99THu8mx16TKpnGujiMLda21OU
SkNirqz9FdSB1Rfk0B8nb8RUL38fQiugPZhR2YLkQlsNixmx2Kjm1jlgHO1OR92N1GuGN1eUYM6C
vwc7Hd+5Cq473fEqHrXFewaIKRMbFh5Q5TL1ZgSu1wuOHoGvinWToHgAXbiBE74H/juaFqM0VXQh
QCFK27CCn0PFMrmLkNHyXi+8MyYjDWBJBkzfHnPqJVb7lgvoJBFcIpne/mSxNyzt9fBbT6QK5yg0
fElxraFgiRPl18cfOlj5veaDWUC6fEoaQ+qyzbFrv82OJarNnx0biE8ezqkS9kEC0Fh4JBhCJOHP
qYIe/Gr2V+6ZQ+69rfwULGjOSCzQVNIedg4+bzGSjr3aH5bRr8YBoztaFC24GAzLuBcLdCDVBEXZ
epDEgtnc0j5IBAYg2g55hGLBqd8XcUpaedcL9Lbs1lzHgsKgu5uhR024DV2A8gHqNiD1BJI6MVJX
2O6C4T6q9e+MmgS1Y/UZHlr/mW6hIOYUh0GKsb/c+iBaw1EMDvLNpKU+Ysef/jPeknwb7vy1Wp5X
HlI7oYBhZFwPVKW2QIBQPNjzFCxuqlKDx/XWX+JzglFX/k8LFn6Fnnk03g+2TcN0xw8XP6rMqys9
EBp0l+k8N3AarTGkm0NQnpSS3DipFYw79hzYDdGwCR8lv4ZRf4nQrwTiO4951wgsD4WdAE+dJ/kz
/9GI9bEOeVMCDpR0FvGk5hczG20hZQplDpVfHwLCRNVKUcsaWGeC/qbYH69o3gssO7MMsNneH/1O
4TQVWL1lONHuxUbJiZTeQXSncuU7x+AFwBK89rxtvEsDc55A59eOoEoz0eLEEBoDZxA71OKuyXGE
pKqhbSTpBfJqXKDagABIns2HHrPQHBI5iTxYIhsCGq6UXSZ9zJ8aK+QnjDKJHn36eedHYKmzGgPm
+4+24KdnEkl1K3Cy6e5vFORiUqp25j7XGwlTSlHJsuNqRODa+rC1xUYm83Tq5rpFxmOBnoTgkTp5
csxfUioS3M3rgV5otDENJIY2eRYHx4Jy02U5S7xhTQS96nL2Udc90LwsBXKm9AxiADKhR2L/ZKT5
CEGpOOttlmNoc/8S77p69Ci6Xt9uBFZ9tpLaO1mBXNn+2NT+XSAHlq9LSTblzTp5lMfUYNgGgWn8
+4aCS3RjOi3YhHTpvP0dNiT51qlom8GusfWZNBcbf0Keft+1g+iSf93IroLkkoz2JEZvQMPJrhWl
irFGrg5ahJw8M69Fu+zRVCaq+l/xA5UclfyJjEdFK/SFaaHCPUzwe+NKWaeictpdkBQrLIWSkqEt
Zb7kduK/ox0rKKJeqYxOZsI0QggMRK+3FihTNH+bgvtlcSr7CqcsiXYG/ezZTB0jLnMgIACCugq1
35JvogluJXanG4A1gzUKYcj2cyGC8fNmvV/91bYxANm6WTUPp6X6/6eYhaaKz0WgJKTZ6tLyYAxN
qGqlCbu5zbsBbiyQkFymlyVVwKQaFLtcEycMOwsOMQoJyLGkpGEpn0hP+ChObitraiMSnD93+Dxq
I1gNyUUgKqDx0tS2+NpH+66WdOrwsE7+kwRqr8YLI7HP36W7pgzx4672txGlAG9FBOTNYISBEuMZ
GXRfo/6woI/sqhiKJQfZSI4ABXqC/o+V1N549jh62R0JZPPu4RRbiEpY0gnKkTSJE+n4COvcAJQg
oQZGiPvSzU6BAs/koUx39AkSMA6+eLs2Y6ypOFcmMT1v3xWJG4csi+fq/rS+cSfoOI8SILwUwNZl
ZVNS0Jn0rUfe+90kTXc1lEPx/IOrlpWbHP6lqGlW9/9rNC5T7VlvA6L3coF+4R6WM/dY6tiqt8Xd
39DbZmE/jSiucez5cSwfAhtCQLKT4MqiV0gvyepvQ4GbNuRxQ0id2qBBUmHA5nO0W5tRXLO2oZMu
+GYanRAH9H39yMhclhE4PlXTRtdCgHSmbVZgp8IfLyrjKnmjrZ6zs+KKMQF1QqySpZbZnMVJypFF
SevhmXKwjdlbtmPdPsxP4iKs6FriyGiV8nyLQrt+9cVWJzADru4vzNNwuiAOQldnACSBewLx6xGd
uP4p9DpsuOb35Ih4zO0K9VbfRPN3Jkl5WH30izvYzpx4qmXoQErf4F+9SACmzHi4YB6MVrV38fYJ
42bdorj+R/VmNIbZa7v+XHGukyhxCgc92Z6QRcJFGR3zyYhea+HHLdpQcTu1vBSde98YFP2xr8Dd
NxbUr66Z/imM8Vy1zL1kuQ4vlpx5qdNTAVOfSRQdptod1BxP3UQAKEqAx29FMXL8+YEdn7OCNk5n
9NMo2jKhP1luYacQ+3+zZNCiKYSSadB1ihaVRd6BuFe6eBt3x7K+wHUuEZqU0Dkv8KU4h9zbyHgo
nJGrSqtrLs465B6emXcL3H1ZSm/z5K1hLT7YBdgAS6esN2uPkV8i+JLitdYHHCtkP2gW/hiJBLaR
+/Wbgi7hqPJyR9Q+AYV08VW1mTT4nhVvubn7xbflpRmWTU+gAeZAc1V7bzZ1EliUviTVu3jWQctr
S3f3KpFT73jsXIRE2CmYYjWEe1qD10UJtGnh+BX1VRP4f10akBR+VJ8VY19SUg2R3cyxKWmwL+Vd
NmZhfMX5kieKYnlPNFlvDN2VJQ8Y1jaQh8Gwr3YDLbJqp5NSwBiuGnFJrlnCMiJmPCXWR1IXNU0J
7tPYv9YX5Wk+uTdG5O+dZdx3gG9XkHkhBWOT9JWdjdDfBuqcHLIM5mCDjEXWQg8gKSjAvlYrVMUD
1fIYU9YnbsSXnPlReG9fIG1LL3FsEH2BMOaPcuLOH/dBW2RWJzlGtF5J4bpN+QBr/Psf9eUmqbkr
AtSq6a+Lp7qCSJx6BX3GUBtfC5DNxsNatGtVmyfA2JGUNfYDYEDKLCpe1KHv9eva5uXvGmw+AmWn
TlgeHCPExSHqz53qIvzKaaMZ9Fs4k8uBebUNi5ITNEzOihFzRdaEs950k08xGGXZLEc+Fis54nUN
TX+mUgesHkXYdgfxWe6hb/3U2r2lRJh35L56pHEO5qaozXzYwGzZAikrfMhvkeDN0Z6W1Dq33rMh
oaQsZbRSy15taHgwuJeWWyh6GVzirRMVDEg41nVPNrrU54tsuu7rL7xnUQ07CQwbPhe8WwPgVNl1
E/JWHk7Uek1i6KVrO4znzg9w2L+WVXzOsAdGnJcDXs9cvFCPzLoqIIpOLpClQGJK9+CUtpaXxN0r
pXY+OcfiVEp9pGtfr6wn8VJA9a2vq1ITod6JwNrwtBpOgEN6hNyQ19awh7BMQD6ciAHR84tGkhpg
b9S+80U5kDHjYdB1Xoo8EVvFmmjnkmR+UDfIcEIIPSsQEomroCpsvU7zQD/Fy2vXTzgWgN18qH8S
ilAyxeZdjpFpCMIziF4gWMNWagg/98RQ/kYSTR4EfhxBktaDwnn3rdfqrMzPJVnZuPJlDdmrzjBz
Gr2NbdnvqiUrN7Dq47ewATzWoocmJ8AsFlTWY/IO9s4qj+rghyQW45WJxavxUZOsYxeZ0YePSTWk
YSBYBj7f0L5fEOBf9rXrbpo2D1OMUoZMKACHXgWUE9gpRWTlxSWiVECEFddyI1MF2wMsXXz4nkkF
pVSaiprMRaOUoQ03X5/QuaZ6Xs7prdPFw92b7Fgdgj7Yys9kmoDBq07z+sG8LCYUpvJZbVk7sc/G
zUosD1I5LcU84lnHgZUQ3Hpw/YSP12lVMeXZZMsErTE6xDZf3OCfBcbjYyoYTZsj7YDyCftVXIY9
ngPKrks2l3ZkMlMviUgmrRYViVknJOznW3BkPJ2nFVt0A2iUjBESHpLD7r+iFfmBl4PROCTWsFdO
luSU9Z7q8x0/y3raojs5JWo0oWT2D7nZL8lCyvzP4KDzvpdtYBolbYUHq5cUIdknhcTCaj1vS1FV
3yJlhVO5N+AS2sDTMTIHl40rToKN7ghd+eNxbfEU97LISegQYBMg0o3dSMv5VNCF9jyMD+sErmwA
4uKOxXuoArvZX+0ICEY22X4V2QZUxAnTuzbskpvIkVHNZSi97v/ohPG8Keo3RUivdnGOvUXUV1rQ
csHQy3i4HJM3lubeWsIzDtJ9UPsBh9K3EVKaMWy1obDkl8Quq+dTsgjkRcvNQgV9Hgqrm0zWxcMF
qyPfo3YqAn7puVsrVWrcIR3m4bfoPOdiJCyUvN44Fh0xY2OSk098W2vD69IgCIe1Qn2abvvAX6V+
043tgUntYfc1JQPCHtRq8h3S7bh14rLR1TwE9Lyq/G6TUXrZmKBEnGj/hYkpsOkt2asIZFBObZlb
hZy0ROotVWhKmcHvILc+M+i/TsSXoHssW2yz/NHwA630jmS3feik7asYvU0iWQHly5gt+9rQwPpT
ExbjiBvhtWcyq+I4SHM7HhZ7rxvauEqJzq/naHeBSpc/A1Yp2fhWdaVawkoE/JQ1tsepm9Ihh7br
U19snKkvn985zFakIMBxpIAKHGdW3VPbkb22RDjB+CcMyPtxLSEpfHfhcTMxwdgHLt5nz8eZcLlq
7tzkIqjgJ79UL7o7GV7EZCrrSFTEBXinhsyZt5BbKjo3oknxqvmkgF8k8wdv6GIf0qImnKGlwapL
rA/LtuWSHhJSQAsV75bPQBZ/UPg6SseWlBpGcPftN/5gD63eRrI+p4ZBJdUnOX9AZRXQfsNKia3r
hnfPfGghypNxw2lQDDLSKoMPxRcIUuOYSVtY1AmprnjrPj6/QVWhpYAJYXo7d2DstMHroHR6x250
uHuLitxuJDr4y2HJ3020sRzkpu6YlCzoeq9xm0ai8tp8nT7rDF5vFmtT+bMonD0EPswbBL6IMOR3
ej49hrXbSR26GEKUFsEyAFpEywfK9VHBPqqoixbi6WFS8Un1CRLs9rcO1/ORYask8xasZBB9x7ll
SKTp0DQTE5oOulZyW0xMI2UC6A0RO/Jr5zBgeGRdEEtLlGMwwJBYD/d+SC7tL4+rlZj8w+2RRw7m
dSVQ5cMLkmD33TQoZ9+qpaS7lVTWmckfMwUF+qZUvpv3cyb0LVA4D6XCm5T6IAcixMVoRuLoVrYo
Iz0p9TPFM0QNyIeu/dRYsD4U3iMSuMiFLY0RsY6evQX3xyUOn1PcYkkdS2UqRcNlRu22EJcyQA7p
wDAmngUmgv9q9FhNOCr0NAt5pTXm05+vS++R8reaVdHgFNEfI9tFQNLvmHO3tf1lVF3qdYe2GObw
E0KOHnnGtq1xXmsLGksOepcH3TVljyzEN2W7PCutR1Hnax0LjbvBRLwPbEf/PHzgzIz9M9ThmiaW
oUr58U4T3qD6KbRi/diI8iK0MzlZYOtRAAvjxpezYn8mCWiNQu+ymB63rcE+xTy9bbFqODUw/ZPX
nVTrWBzoWlpxfinHdKOleVTpHPaURO5meAzHj3QmvO6klQE7fbBwGY620ume9KgB/1hdjohOSGc5
vPvYk77LdVp8XL51j7c+Y2TzpokZcGROMsglDvPBB1a2qNE8rdDkaX7YW2DTq7FInDWK6vC3ohKg
9qJNFP1xMJ3Leg+00V/nARA+ODpmseysmKSFSICxNZcgtaLzeW7NYwaCZBKA7bg9Usjavz3zhPXd
OTvszYF4M2xnK4opvmRJRGjueh1Y3u1FT7NpW6dO8zMUbpmLnTW3WCtmJNBWz2f6klpftjTlL9Jp
MnmMVCq+LmZEWuqjeUd37VrFKAVYRWjVZHE6uHYRioRz4HzsWnQXehp21fFbKSS9lQhrjLOivPwU
L9UxInDzkn31b+sIKPDdnTOxcZV6aOP3f9abIAWN3ez/zkzQBQH+JJ7CVQf+XzcvuI/Xjp+3jqfN
fKyL9oUU5IbrIijJxBqufo3nBLtMnK8xYBGlqYBOY7ZjqSf0ZdrxHfjYlrGEZfFn+T+BBTEhGZxO
FzDwkmAYbqtc2SGLBRDCkafpEeG7fnIrD7DvBDVX8IFhuFWsWvmKyx288QuX2lvXgXvjd6S8pXgJ
vBlBHYWu+qdtRKP0uzfN0WxmDBowSUlTlBtj2eOP6dt2kyPjIc8zsKze7qnbNBtS6n0pMP3SSm4k
XLqpUAn8inlQyw4wLU1pegMGrYeB2GaWMe+qPuEAu7pMH1xc5TLpusaVn/U6KUJGb5wu9VYfWd1/
ESGUEgtR137iFs2pAW/sjQlHrIQmWqy93/Pk3Pn/IVNZ+NbuYyefntE1omR+aP6HQyBrL3Co3gEO
eXRxXFo5TSgywTlqasczv3P6Ssy0wLLS8GpmVB7lK1KzARCRBb83BHMTA5bycx0EbiJgd1MU9WIX
PpQrrXo0w856T1UCAXqpv1nlRZ7ywkIJzRKfyt12pFAfAxtvMprwm4lAV2JStfzYLN8nLClu/glu
IcrDLedQOvMY285iN8jLEgYOslXr90TlhrhdLXmFK4bl617gSpEeGWxsBCrRxi/gCV7DQ1P3epHb
JBJKNwQolv5Vsk9ex0MAX8ail+sg9V/DcT10tdp7xwRpeX+HzQGIArgovVyZb4lOoJWNHNWKxSGI
KG9O6K00v77gn9leo7CfZjaQdA133zGgOKLm5bzSlXZxIMRRvA2w8szaZIJGwQ8mun2MW4JGPieh
zOXPKYmINXZ5JA1YK7EnKJqEHlj2/C/NqTM/IjhC3xuO4jrRl0HOHA3Fgz7H25xWIsdfXJ6h3Ggi
bxukU2rrxW5uH+LpfFquBZAvpZU4L5NT7baIiRovF/iKu9zjtu22ZBjRiV85RrNtdXgStJaApmc+
OZ/MQ3q+zk+TBL6r+VrXUfxqkgHbXSQBCkJ+12xenx3UlvPrmBCKEx9a0lyXgz7FFMeBG+SaFI84
XSF9kQ72+UO8J7g3T6J5eUEHn3hGR4XjdXmBVioo4Kk4trhVRIaufDkUs1rDjxGjt+1f3Tf0w70E
Cw11r8BirCvyPweNPYcQvJP1czUPIf3JW4C2hPUStl1+cU/XHPtOR/TfoQb3z/McmNm5XATGscfJ
NDv0dJq9wL9GlZXsqTbX4rhwRwZs0e1b6KVWg5T6fFDoMLdfhHn35FPCPl8J5v77Z6AEtkraYkRS
t5VdNzaoslWJGOjhl2BAahnb7Igq8IwNXYmKrTRgL9ZjQ86J1PsNXurm3K1jc7y840MVztKdnGTx
P3c5cpavTk84UkdxG/zHxk0lrwuEcVGNIMo8S2cIdyTYpAVI1fe89+ihBun5pVWjWNytibOH1Pf0
OCa9MKD9t4+AdvnQ0f+yj9MYJYlPCACamE2xLzUoC+GsGbJe1V1i46heBYGMawFjiufMID3TAlz+
7cr7/neW778JG2HzL41TzRjFNNQzknP7mgEWcmvxy7J5Dw9jRKXqIxnsAkTJz1Xr3KEkshqvyWKI
HbWk43qOAfk3ajaRmp7sMKEMElx1rf8qe9C2n0537cbB4QO7lTsb0jfk568e9BQuA0R9ks7F7Jxy
bycgsRcj6cAbdRy0ADNHL+YDLfT1gGAJTonVSf7yU15AwMR1Wtf26VwneoRWo1ZNeVKeWjBIGlsB
pEsz+Oky6nhkNZvXf73o3KHvD0eC1rx7oHExUqwudmXBsRxQpdph3JtQTvhhcbufTzbVh5o0D3cO
pHNaDeHQ0PLdpJTZ0mv36id9AWlgtVpzMN2TVcN1A8FKpcvc0AcsT1SrWm7iB9tGOiBt+wyYq4ic
6tWnUuJAaas8ZIwNJJeI3Qihchmt0cne0p7FQYl1tKnyfheozBs1H9lplS/nfvJ+jLZhDbcyhNGW
PEP1IPl04E+GmLcRWvbo099zsqYq4u7nBEOqZ8V23iB+TwUOFSz5gJ47Peo4Hpq9+ghUGbXdu5qI
USMb+RsUIIz2+zSK3hhZHZXvUmV6U5+REQlspjDcI3ZvuyNLkQip125CUhhwHI0tCoXFNAOaYKF4
LUwx6Ju35iwtkyXSShNoN9gRBppSY1gC1W1bKjKhIvt/HW9foMVgJeYE5EPJU+LDvZtm8varNg6T
DQjEE1Q/EVJShIalRAfdIqkEW8JGOC0Q9oe1azB7IIHnip/lGHsGlUb/F38DRfJ3LODmt+TvAWAG
5Ppj95xadHWaWoNeR2sWk2mKYG/DgeURsa0ttkWH2uyFyAwLicROuXv/gtTvYbpipomehDkDJoaj
7LJsmOGlTFeOVYvJhWdueSWnuLX2auN0gViDTr/oO2YfwuzNqqMPQF+nxW1kLBsJ7Xp0z2u3X18N
+cxDNMWDUK9CqfHSWPXHZlIg/1xKHE3pAoENHlt6wdMlU08WxYUaNcJ0tSj/evsPBwAtdNwAynRh
E2zhH8Sqma1zYvuK+XTmb96MjL92YbNQFmgOzkt+zqzClW69b8kMZJVM+iaXJgEwbmlhjiWh2UBs
OP70vTw5O34Bslx/a1v+MEQkMHffpxfQl8GyjCHdjmoNo5tEZVtmeA16flPgjvccQULGj7i1LjKm
sibcDLzJOFGX/FidRqtzhPFkXyTqrfle4TXI8r7ybnfWRxXu/zLC7epyd2MXTaUk0T8QtHpXWMIE
hDvk3JtkvpSVvsDTqoNhemSkp/UJ+S7DUZBPEaCTGhcLuiAskPW62iEd6Ylw85sBgGOHJ55TwUat
iulvzxOaP78ZZxfQiux5srzCfRGzpUg1GWon+V4ahL9gqWIPzisku+BvR5WvrlNitnjKysjTW1SN
OagQkqWLGb5Mem+/ls977HCylbbkFppTlYdiiT2dYpeHgko1z2vLKShY+u5SrNSdlEVgVZFDgvto
+P8AxO8iEnoRbv5jMtUMSe/d/8oR2T+cf0zfTF8u5NhIzJjrtQg2l8Lq4w7FD6PYAUyv6Kn7Mi6V
gXLlhxRgyTHGQJJJYWUYFGZqCWQZXfWr/lt77K4dMyQgEwPe3QY7coYlCoj3Y3FyKBBqLj71/Hzm
f+LgKLRCgHQNUoq/wjAGlDLb8UONrZxjPCdv/owETZ3tGYLvP8aYft5C/cwpDgCb1kKyG4DD8jYv
YPWvFC5/mfPK+Zhr0rTpZFe3lAc364EfT/IXvzs9cGMLmRo/bVu9dWkG72LZvmLr84UFcCoA12ji
/4dgS95TCJk1k1s1cwEplUEYhRasAnN5phTe+p5p7YPf1Ze8jWpBgCjM/6EoenQVa6sdl1EkVAPR
mZ0SH1wMW6bIopvtzEuDvL9RW7M7dGaw9tEMGTp/Oblh8Tpajgaw/mR8KehiC49IF8Z2fx+YluXV
lwXfVpW+6xs0RFzhRui+xPFXUc1pNbIzJ+7Z92OfVEe9VwCO/iUDIgcbUJ5EIzrA2j2mknyxlkCf
KYfce/anVsJo8YNC+1uUmEMTL7e7Z8b8iUHQBil5ToUlCDDD6LT+d6MCg5ygV3AYP+4t3NN1v3Yl
jWPRCGjlVmFPWt5/N0tIsgstUh9U1JLSwn1UuNQ+PNCsbTV/vo58GFMjESWc4Csf+zmjlwpWrryf
/KE/FvyJQSOo4rJlq9vWO8qBsZiZ/dQADX8jByaq7IhHwpr8/TAotPh1exFK88h+scjAdxzulTeN
HNOdcxN5P/cBGDJuuivClw5x8jIGBeqUEhPtrYKXtEyVGhvS9pore3W5xq8ngocoqIGPIF9vOlo9
jhDQV7y+XGqErJbXU0Ptz2c1Md2qyqlgX4IqBDdh9h2EOEtM8fgg3lAbQYL3weRGR72eBSkTemNR
G+xR9KrfSJfft9i/Ov/TBS65NVF/+3ciBowgpe0Iy2tYQx/pT/AzKiFTGsScWsBs/GJkKREXr1aM
Rd+hwdaRGvl2ajifSbJkPx3s8BtCaaOowQjq4KjtS6hmsN0RUn5BDmhKTYbs1pQegtVquI7T73sg
VR4lH1lOHyNQhFhK3AMegESIov1pf/NumqyHFu0z9m6kNCEo7e3IyhAxnDdP+AkEHtVFoRsn20+p
fO9gBVGkuha5oDuOeWQqr2qiXpqJJ80BsoS23ddoCXGnpWi4Eb6wHI0V7n1kI02vlJxzqGONJmPo
MtA9QUWnUVqNp3VYYeW75/z+e7c9xQiWfzS/AeA9DP8j79GAmhamllydcitI/7LBnbybzoKp3/Wr
xnheWoMamoBrpvzI7M3XIdqL7jrffjmAc0Yj7uBA+B/mnv6uITPMK/kCBPeCUep6stUTyFu//m7v
G8xadqK80FlhWqijjcCb/rEJWaQ23/FNtZb6fefpLWRgJ8ptdDmCrLMUzKBoyAcHTE9dou/U0pNq
ts6ouz08ljDpKyqglQTW2qFOot1ByM6VKd9oeoLO/eF+dGItZUHz6aUsIkGw+LIFdO9jF+xFRreN
QCI38DujhDEyBKnKBN2OSAcIvd2CZJwJpldJ4GQe+RXRaTC7WDRj/Lzs5Xvr1ooiVDPBIZ6DQjbm
5HHzU7Tv88rTuYD8v4++P/Qzq3jJOwrFZx/TDCnh3sIuyE/6jX0Bn6lczcB0odwy3ujiukMXPbu9
NBS9gCisVvm+tmpr/eWQkKMTMw0R8CQs+tT1u0vL1ibsCiPR2NQGtfPgo0Quwu5EJmlBKbeZGiN+
Hkzkwe/uc+JEblPWlbPQ5VATog9fPjfjBCNrkJO0ANtZIbdRo1VZt9HJa4rmmmWnGzI4+Dck6hzY
ZU+bTNTWlN0iAFZCvWeP/kdKmo7o81c7BK4FCIruuneKGiYB9HFD0R4XzCvlWcKCTRd5DN8sxywY
MOe2V+GmWsiGkuuR9x9xPX3XfFp3dirxZ0n4rWAmse2bIUZqYqLKxFoPZFJCcSe1mP4zEe9D44ww
HHwsAj7ghYWWAkMs8giCr4UhOZPFo46UudurfEC1f0qSFVXWhr1bRD82WIwStLkBhWULBWKoonVE
aM0RawBf5uLrAE/jxypfkcHbXQZZXG6D+gqEjjVgJdQTeHUjV0RKYpsKFDAhEIuDF4YmfeO4HfBI
qntLuMkJAT8s6DKkNcCYzyV2vW1Ghbdfu9/xoX95GcKBaVYD+2vrZOyXGx1zrjN6bXJKPyh/8BEu
Ed0ZovyC0HjC8PY31pk3vxf4TcMQREM/H5yM+QmbAa0d7nL7dM++1Ocl+Ri3ODyZ2rqw5lOy3YY9
6We8aa2qog6xCRHjke31Gdtax0HhGbMgH9vDgiFsksynKQkgjl4TEcRhaOVnYSI/TOuBqwxTx5Lh
6/tGxYpK9c+WbWzlNdQLpCi36oGrJzTWj8p4PO/JiT012YU4UXCZZddaCmINGzQpSS6rbF5T8zbd
m1H6Na1R8B/UM24bl94zjzFAbxENviT95v1eyfYKgweqUMT8iCwuI4sUm5q2F8JJx/t/fug14LJj
VTxd9PlAAC9RQ8pMf/24txFAl7xaLbVdDwZ6eq7xre2m8mlUveLbH/JT85eABV7i0tAs50z2rnas
6ugwRZoBjTmxaRimf98G6sAaLi5B74XOI458fRqj0d7myLx8tlt2CZrl5vjczH75ou3VprBLkQ0i
paDveMglnoA5UpFxZIzR4xIwWTvEWq3dG0N44NuvUQ7nNFmi14DTUoMM2nnfALxX4cNFQ3H2nWt1
0ibLNLhMJeNs3XqWjCd1aZDavSVS55dqZxMqrdt7GzsgaExS3YHFZHB+DAo5MHmz0+REcl9RIXhc
QJkXC8l2j+03B+6bSBragiRJuJKspdMT/l2MgjTxWK8FFlb33TolD4aHe3BU2A0X9uEUfpKbddpd
R/Yh5CH1GctWk46t7H4rjEKO4ReL5RLWOpeeaplz6svgnynYUjeDw0ktuSGaRn01NikShhonQSuC
a8hnt9IasJuJhUiNYvH6i++vgP4gttXEWViY02SH7h2WfmjDoSZ2PM/rjz4XNdSQ9g7IxuS4KQF5
WO/kKr1OOnYZc+jumd9AZwlxHWVJNVVrP58+qSTFZhJkiJXb1F48GM2gENEwHYdXSPXlvrfeiaDk
cQ469W5IbvgvOThSbcnopnOQgPNYzz7nwP/zpyxJ2hZc/kb8kfJzrq+WsuWgZQW0JP0J47owxN9Y
ETIrIintIUOuEjzgokrhF9QALOwRjZLVEloVCXSYIO/riPq5EDhNq7nSVhEpFxuxmYKANFyZuFuH
QBbAEzPLFwXrEv2LZejkIcsfdiU27aAFkBKqLEC8BwbQBGsLeMuD1+seAUTFGwHl883xVomQuryW
f1jg6nrWulcdeatn3I1Id5e3n12doNIU47rGl0n7b2kkGHz4Ixj1D5lwIr1QFYRavsbjeTzrg/4/
I5CPFhm0Jc3Ta4psPnrY1TKN0lHvZeYSqqlYCRz2DWOFBy2LtZtZpERZS2AzNS5IRFmcAyBCQ/yX
1M3LeUoZ6N+lbxKCwjN5gBZYrEHc7fm1V8DFKCahx+30hvylMfIOxsUY+jH8TgRZlwCrDY2QRWAp
pNCDG2nGO/oToxOPyc9/w1zOhwsXVOXSAhpjUw6vaXmCGukfIGKucwuAJpO+9Vlf0MN9Ws825C7P
8AgZFP+iRBjnz+fe5Nm9TFyuQceQpfqxnbDQTsw9ZB6seC6L4iQDzb2ttaW/24ZIbzPHpBsLDk2w
z1Mrq3UgQ/A6F+M1YPNSzFEn8I/4vUVO86ywa9mPOEzXDjqtTfimKuklJWhdFIy1UblPxpfJxb6n
q1hkdY0pwe6fC8+tr8X5gPq/sIhOILGqylH+rz5qBSdwy1LTkSecQCg18qwolQiO3+PUBHfVqwVx
HBNHc2/ZApSH+QeqPpWmszWCnUIW9JuO1nWRlVzkEpIDnWUaiJlGWD6ih6AGzT5SZWt6EmFsXU8Q
1MInlfdTWnfggz2r8H1zhufktSc9dWLTAAklD40RBfGwluwnXQzn3qfUc1V19N+Z6LpngTM0s5et
q9F+A3S23dk38KQRlkHggWvmpgtqto0Pzyugueh30XP8c8CeLhn9z1NsXjwTb/3LIiKJYh1bB5z8
R5dkkbTDq5nWoEnobDwCyO7tINtXTgREwyymfYkcwtzbbOnqAMwjKr4xNjxAXw/5y7iLkm0jQJVs
GpLpblnZAXM/pI+KXjXk7Ub5ScxFamGBA1L2yaVeazzmSU7UZFDfc9b642YgNu1REp//xHhGJvey
2+HFsu+6iMbOaUJVWHNZVh7DqKIBZsbJRM0b0k7zBObdIjljSmuLW/pONBz7FniDEzdtG948+r9A
K5qHruaX9d/RT9Op8CAOo8OygIo5ZnEPZ4/qqwxqsmAinFh9D6coboVuE8AyCy28LwBlIOABVdbV
xXZ4QPMnnNRFUe6NP3AP2ddOgkld29vsCXgHyaEDPxzFg7DBzJOhUJxZC+45vfUApSBdiSmM7sHe
fgzMxf7ssoboLKAf6QUmb3hTpNeTR/Bn3wej9bGeNloCCAaRQociL0VZ7WDb2RdZiWW1VE65eKF9
klVlOSPyIylCsOumetu+UDEkbZ5BfTVLV31o/lodPLMV2Dxldg/dt2h2yQj5jBN3kPmFmBuCAdsj
Ek8N/90vP5AqyFQfVu5477v6EWLpYM8rQ+GUDVk/x8DOJbk1Ic4/z7rBXxkURw2n/8QHSwMz4dwI
Wh5s/16ERaG/LkYR1UBKHDTd7yrge21kVrlm+Aw/mOCQTyT20rKer7BtSoEqklhGWtVv+G7OyWYh
i63LaFfQOc/LwpYNpNIbQZ1HN8F/Gt7KPVLrNhqzq+h5Y2dhm9Vxb+hOg7NJMdpV+OkCx7Aq+79Y
CmoeGG7MM99S16lMBiG/ibz4XGi/gB0gWgwxg9y2aeSCQv+5+wWSGrqroYAqfFQtDrCY1siqqFdm
rsvS1KeTuqXCvTREyExsSSfyEF9BoTn5FFjxC5ePm53HY4VTwKmIpMWjrYcZh9SaLh5KpGHQbUzt
kYb7Wh0uQ9iQEzle5Ze58KNaRsHWprYXTxz1ZbY6D+Fv3Wyka+G5/OGP7n3I9FzqpunGLUt7Oeea
EbDY0RKPI2K+JsyPJ/trLxea7Vxyr8nSEpo2MUfbTzVsQu/S9aseIBz6Jioh6eX5sMYCuE6TiG0c
m6ISGzuTeWAE1/Ww+SQlMB3LgwgN0FsU/x4u+BAG4KGjxwu6ooonlbdkv7w+lLnsHPVfWGo+wF7q
F6ve/PmECw0NNJgJqcKMpbGrqhSwJW61slwSsvCsFKa6UZUSSHqa5LVcUD8W/BuqzQEciYigcxrT
78mU8pL/QLSPEzfYCOfrSUkhGWvFw9j6cPI6VrQwwQ72Kdgc70NjweXdHcFaCewQDI0vDhUrfbbw
TJOmWPvbQR/N5y0mJdE5huz4HbLAmq/IJ5JV216oUCntOletnl5Dee9YNcCPq8kkaydPqiDnT8V3
s1zJAEBnqFSRhv61zOylaStM2VNjKyvDPv23MO6o0zopy7B5RsBglSq3KJ7ZxOXEW7wF4atNi7A8
EsC0MZM4V3GQtRZmlbnUiad3bxucAT0yCvkGAnfU5VtBT9BsacYoscppoQ6CBnevwjE3164lyfa+
eHbZJLLvFb3okf508BEJ8/hvUc7YFKI/t4Cf87rHmporw74fyL+JUtNYEoCiRLI3hed2QFb66tcV
xK3t/ez3zzqT1hZscMv5FC5rbh/CMZtENv31f5XkW+VyNTuamPJacZxY4VKgKKj5N2MVITZ56Q5/
kcga5lRuiRNeODlk0CwpQg0L5LCoa43+Epim87uiI+sEObEnXlIk1CE+8M0qrp/MZR3eqZQ6EvEJ
+NGblAqPShxCj5bKGTcLQsgkEnpX7+0lGenXbgHxkF4sRzsJStz8ZXPYczHk3IRqiDdOoz08dhIp
RVSANhMdEU0T92EsZtC+MvzJH1t70ak+fFaGOstBk3DUFwDVbYp9EzqHJLTEO5eYzXUGnvickMWu
n3gPiwqSYxskYyUD1QeU1xeSAK3jXS/igrSv7nj6dQhooNeeHM3MT5VLyf2bnkplT/zrPk0ymXT4
5hmi5uQoT/xvpn5Fpa+hDubEkz6ZcSUaHkttzgClaXZK2hDOmZF1BaLYi+O/eAXVNWIALLkJflnx
aUAvQVYDXbtgOL3v8vA9EsnxttfffA1qsMmH2Qkprw0VX6yoAjnERS0u20J9lBv5vtcW1Sa7M9jc
brMKI3ReEGYnJ08eSwepYnW46rx4rKj3oYHpFIDsWBeqnkDtNlN84/Q/2kOHz/i1h/9bzQ0QKHsW
psrik9B4xpjhJj7JgA/Kvh41U2jXJKMRl/D7cctacHoO+uI5I4ag4BaulKJKC70bIW+PhFYTIdpg
PxbKA2FSOHil+5xBA3R1HECXHblqDmVvozG2hNJzNA3ZhXYNsvCp91e4DvsBPjLVnkUpkyYiGaMz
O9MoA6Uc3IabpZLuzYZCjLc6ZJgFrqV9HjxbN/0D+dtSZzo0Hk9/nofv4So8fgXRZ22t0evB6hEa
T7d6e5VmlKuFXcbeHka8cy91JPfVtxLFIdJt4KaNsjmru5PGwwfANnFd53m94xnxn9r0siiDyWER
m0XukBWEAZPohbNT6TfkqU2Oiw2+n6fzSSvzBXnlY+SvLLnkwVkO0Dk7of7CkbYzJCLYWGzRPrg8
T0in+Lkl0ArNgBTzIlQAW1EEdTVznmCg3nwwnw1sPYEZCw7em6P1dgO+Uf6QEr/WcgrBI3pYFC5k
KX8U8Y9PDx3vMnuy0u8hr1+LLdF7W3lHxF8FEeOo/Q9HCMmf0CMGnqMgxeuF99QnYKbgMHu24Elw
RNapvnIXE+SobuE59+fIP9iMib5R+esywPLwSlQUwR+k1ieoDmoNwZlQgtfdWem64x+HpWJl8OnA
RVXf9BEWbH7t4zuIna5kqJv0hyjWe00jA9uyY+Q3dL76IHzJPMG75d2H4PzjKbiljkQE5koJ43ZL
oYd2GVDtRK3TudPaOlQzhsuJnh1yDpPWXj0vWtK67zNde0YzNQ3fs4q3wMGVrJRChwEqKu3tT2DI
XzHe5NYnLEzva8nCJboMRTuOPfqoC2mrRHEaJkKLzXVakkbH8sXJzBekRglCKy67LEKV3ueyJ5l9
fFGii6D4EEMreaNM0b9+irkx3YuZDZIx4OuC6St14ul1J7yV2r/1BOo2R/yDOHPraaCQ0kPCU+ka
szoieozZlMfsyaqzSDNzMhPmLbZsIZN/kfhM77yIfhs/iv+oUI0sE3gMWZX+1JTzybZJ1v53YTGM
GbRKbEM9NaEy+wE5v2TorvavfApiFg+R6tjfCgumtV8EsJ9lw1KTfOta6Kx/dghty4MsOeKFcJID
njsT542ama5Dm9fEO1kH+wpJBaEoXglpwhFpiYKD8JG9vVZ4P/S6MR3+lv6+F8eDJOil7zuzxi9d
CIEIHEXq72RYCUlgHKyUPzQbuurn6wFNqsEcUAmywMPjyuT+QREjuzMKNGJadrg08u7Mpf8kMQb+
glvfbDDpLRURgSuY7QCbzoCYRoS3ps3q4YC+bMlcICDnuiSJyDFmf5EWNupiZnh7o+9swX1zoV4R
TmUXDJaplNYDx7JH2QzVNNgsxCzItdNzgas8JFyMGbPoGZb4MMH9ORnYhFsB34R03lhD+9OZGUWc
eKMa62/1vey4qY9IMq5ZMsY33n/1xgFy/b1f9H6og6bTVdpznkKXRQlYFe4rIzmGaTeR4+wHNL3j
XKZhat13cJVw+WT10PZ1EF3mYGHkXkeJggnvBj4ukocJTKlKf37AmuhtHKtNrAAoicw3V8lelWbW
Vp1KyhR3LSvdPi68RZT8IBUvT1xsoLL5+fZNyVoy86ntNyGceLi7B8k3xQ4HFY+qsZUCQLQz7mE4
BiSUZnhKaw6C+l4Nj2Ii6fnti/BIPmbbOjQWbzDofa/oEKzq+4rOo+ydr8orIdIaOtXl8Kauj2Zj
npZTgodGS336q/8qDLpjH6qMOaBHv0Q8zoaNV9YIxpIvQPRmEnEIAre0ktT7VxiyIuc8brrsT4Uf
x+dS9oTUVI+Z33baT6AvUIVyUq3vYIlw0E6AFlD/H9jt8wMAYnzHR6JeWiUlF/hYQt+QGYClnB+A
Iz5aOp0dEANTavgvd669s0yhdH4aSY04N2R8CRwCC0em/tZuCUsvEHH9f7J1icMwvK20Vg7y+97z
0Mw/aakm04EG/Bu42uqVS+VtskqM6QE4oXKokiv4mIZrK6B8LXiLXIL5KAAGAPuAEokG/9TSUGqS
TKrPKHUDtj0i5MYie8EBKyyF59MK9plfYsRO2uaPoBa8/n3drpaemCza7LipE1JV1BtgkQjz+3Sy
gmikPunZrIX1vcYDOfuhKjtcDhVla3Z/rieJ+7abFrJ12eLKzFOEpsexhaFBBqc82f4+EpxnUn6p
XCOIcCH2XSbP+zQFfs6VdgOz3zcARruq3NZgHGPtdKqePPzK19Ekpp4RDfF+vSkIf68Y6EbmC6Lr
S/Y4wKRcfJYZFOBnTOnriRX9m8/wWltFdsBHRvQ0no0TVxga0FhfLxvbN5rImpnrlu2jHONNkup+
oc/jpcq+kvtrorcKlE7fIp4xHpxa0shNHsvZNQM56FWKWENkks3H+yekiRrzBqz2a5BmCH9o67qz
shmhjj8u0/7UtRExou+TJ9RT2LDOGGYPgratCSd/6JfQTmj2umkyK3Y5cLpWXZJ7bOwfiGVbN0+N
79BAMFS2i/ynqNC2JBWL5JURx2pJTjMF2AppIC4qDs00jn5HU8fXckEItyoq9ki9wWjrWXJ1gIh0
ZbgB3mosVoLcgJtSMoAq0Qy6lF3kalezVUyES5nDMsNUhOPzLRdrsOddt0H/rsZ8AmqnbWpjrxri
3x1SjbuEPzTQTTQLMHMjy/VYhKCZXBT7Y7A6CZCrJGL3ZkdP2TJH+XIlgQkz89GWWzsYRw724wGV
QVRCW4Ejp8osPnthISxIZUCRmZqx3glvBgvl0yTJzHjujs+UkbiD1tLsGMj2I8Dcg8WK1Vm2g4Et
wPRrBzh++jy80PrAby0DGeSEEurLMZe1kfDjM/YD8TSyqmTVjjgOv/w8ws9C3W/r5tah7vGaKZem
IZ3eurNXA8F3nSK2zjhCmN8ZEcLCaKWUGaoegleI0AG/EyXKCr+QJjqZmy7d49uD5TKojxZTxoDP
mLuTOJtiAiFl992uF8EzFjZ+IDbiTGL1PwuRHbtaiH5MMLWBS4AiyaEb1BVCl/uA4UubUU71rUfG
/3qg7XGZrVZc1cD7EfIflMbMdTZ1RpISgFORFDPzl4/9PDn4KrftfEcRY3QV6M51Bb1fKUyVs5Yo
Iim9vKy/HFioNwx9otu/JdpaP+VGA10G1S5HHOITcT+3Q307c9OYjMzNotyELTmkYLIfwI78wpN2
jyW7sK9Z0vorb8fQIm+nImRVuSGHh9hnNvoAOqp/yHg4SIH3vRh7dNqqZ+G/nEZfF23GUIY2BBeY
YzD+FTj4QhreLr7DO19EuX3jztHL58bx5zaaxZOEraJEbi2wYOnhOGhNiwz9Qwo9fEBi8lM0j1SM
oC5eX27JzHROYjB3h8e4MDFREH8lsAc7Z1YZa9O6Nlkkl39f57DnQwjOT6LB1dDy3jvNImc6yizo
lyiamBut+BWN8EXFTrEnNOsvLFodU8aSq4cj2R7j+2tH2pUf+e0STmKXUnyrKA8XxK4qUwEq39bb
NJNZ77t3YbMMhLb2X3qQ83DOsumiJ/7f6hbTs2McDcCukJmMHYT1iTMJmUtiISra6A3XV3brBZLI
4kw6ZC9rI0A2hq74fVRUW3GJxZsUorj3TsnoOAvQULrreOUOFvFooHWOtCaaOm9r/utGLn5TZEfw
/Z+cD/N7oXc50E5D3MTNssycg/WA0MnWsG/K2xHqYieAreXm0am8wq8IYC3qc1y2kO7g3VuQ1x4I
ig93sRAI2bU20MFHhg3uFAA98LRI3P0ksvkbWCcjtr0wIM+8Bx0YR9REYdcU1juIJHHXUkq4dnJZ
2AghXyVpU2+E+eVFy64u61p7mWdtY+vlCF1Y+IJJsuZy+61SCeNxJzsNIRmRSkNWnmy2eLjECxxx
QfkQpTKLZVF1+2jumHMl79wVTTHmP5ncxX9o25Ov3l65iKy152sPgfOKE/6wEyPKU7y5TgHlbVWu
38CQD2ieVGONsaAsSHh+k5Y2uXrtTUJ6YjauU8RVJxT3M7q2q4vTdaS/qOWHHhgBaBqluUW5sU9f
oe+QkrrO1p1/7lHx1iu9ZWhJ054zyGXcPF33yVf7EfWXOYC7epsUSMgRSaeZYW9Q2utTBd3Pv1Lm
5sc1W8NedWEplzj3fI8oC0QPtCQhw3gaoSFVE9NxoaCSMXPN5c1S5NdR8u8elTdkGlji/u9zjWW2
0aBd5gkMBGut9Wpcm1c9wdMGZvtrS3brAaQw8yNSVzwURFf+rE1w0BVjJKt1XTPBRtaxGhiABWA1
YJYr6af0+3Y6abTPgaPhfYmBeNyLeT5GdUP7D2XxWJnLGnl2JdtW20IIk1hN0rxdfCIiBUX3QnAK
Fg63KVuiX2MRnHo+6wrkaQv9tOTKtb37HP0saoygW5pW+WCjAYO7MqMs5JxqWseJBqnmcO5r0pir
4u8S9E/aFF26+3vXtvAHgoWlCXvw2sk5XosQAOYEtI2cvNL2ymfGdhRqvuAeWyVKmy5/s98KIdt7
AUfF/y6L513DDdpwIfJEWSJLFNm8C7UcUY0k+QHZLEVZSKijdvw22JbB23fUpMlIZJIXNsSdRkWI
WudAFNsLSFuHmDe8ymSXRr1kraoAJXEzWUxJdP/WwzwLOIKSI+i8uUt2e7oD0GTibQ14IHe2oGPy
99yhA3z4AVIKE1Fan/sd+Aihwa0n1Bzo0x3jQsPjDFsQad+rmAVNaMHuzAF+ckHc3PvCGwhCal88
FgWHdHDbHwAFTt46ecKTECX+1XRhmdXHq+/2fLxJOoK8Mo7yG/8JDEXBdq8DRO8AYAQYs8R/nEzm
lT9uqXJz8huERrB7xesROK/w/5eMNg+1Pt7ux1/vm5N/TAzqzgjvCMxIxc2M0/H9Z0sTvSU0fiou
NaO008Su0W3S4X2QrRdiM16VzIPwOAuX5PHXigS3v4zfRM3R2eg/Twzy0pAmzqsmqSUVZky1yu8W
GmDCvAKXuse36AzjnKi67HuHcaTfd7VhDVmQCDwAhf2DaQIsgmd2crc561lM8BHa/i0zUxcmGkT3
HziJg6s+CUCMHgcna3zT+CI9PqVhhXW1h0YSbNU6VQIuPD0MuYm0dFtLYX/PSgUfgWV/F4UtUCYe
RBQMnlgEjtn33ZMxOxQOtE4zu81sZhO49qgtSLbzklJlfmqVQMfqZ5rGD5pgOuQMDEh0HcftxaqE
aewOxX3jVFcY3O9kzdM1mE+3bHtZpvVzgxZTOx70yZRF2mqgAHiBzH9P5THQjI7DiqvpAVSenfka
oGDFx59IjI6KesSSvdULRRV8iVMPIWzmnl0lK66MtGPwovfgP/K6Xp/vlXhBIvRg3kOFdBQADPEt
Y/puV9H6rzFqwHHoyUfpP/ZkPUIILGPDz7ND+jk22P7SpNl0lkFg7GCLCVqUf3Riel3YNxhy7E2M
AqwRy/N6PyYGHB9SGkalqt/mYoV3gJNVYVKwTYHU06q/xAOAp9Bugodkct5lZLk1hS+01CWq8B5U
dUwGBJTjYQBtgyUhAlmHhxzJIQcmVOipPZ4cW03Qzb7DGb2h1VsMuqLt6q/OaOSEXxKO5My4wpoz
wMtQVPxvuRIMwNz8C/wAJQLYg/XpLdGb3vowHLyv90BPxDwS6FobPg3bgMKllc1Z8yhB+F8yZ1Kh
20CTxayAD3pUnJGBRcVCvSDsAEfYhdEM2qRF1FGDF1bRBlLx/GjzNXL32tVZy37XShK8EJgVWQKx
5wTFLJmTxtNzKID8ztYfJPD29SE45jN+BHVRBW8DbsjomU/34Fdvhq9at2k/f6TCNLw+3Sg77+KB
WFngx5CUPuIFY1rZ3NKnlxw8qaN1Ehq1NWre68sNk9u5gmCMl+BlAy9SXehlV2QsQQXXq8TIX8IV
ZehVhw51OcDEtUJAC3nFWutkBUObgfQvXDpTrpxOIfDA8QpKnOtWnQgg8j8xyfBz0LtTEBUjWqZj
7McOKJn9CEIGQwxFLELYB5VKdAKOyUUlwrp5AnuaQsG2NbmUC10SrWirWpf6Oe43iFiXQuwtRm9b
xlWO/JQ5Tka4v7IhCxuIKRitGmsaErPkzpQuruAtVpqSSQrE5/F3gDXvGC211pYSoS0x+0OnV4dK
nA78IYXx3YAUyiAk1Ehc+e8ArikRgvo6qwRxZb+AGnn+Na2y4dOym5lGQAuFAZYHaMhN08XbxbZa
zwUUY6tt3C+julbOh2EGg5nDmhez7weXFHL2u/9oMuQmR4ecQW1krfQ3AtIFgrXQcmmZyylmC0za
I2D8HUht/HrIJHwrQKQahecQ5+4ybcUeQGS10w0X2ujdTRQIlI8nHTe5kOJz8NWXSHtz9DQS9XGM
EtaMtBGQx+gNkxUludKkzcyBKE1o6+rZVWAEwrQoQ2wdRY8Aydwykr80R4JLSQzjesSWPOmo6zn1
HgbTmw1KiIjVa2rpi5c+Owp98d+WLzkBzY1HGLBrYN1vh7PjjQiRGcazESvM2/s7Bw4EFa+gywdv
hyiz95WUHMIpCLvV/ieD6riCB31BULvXV7/ursVgp0q/6wN0UrcaaZClc6/mho38lzz+uxV2bN1u
V5HnoM8Pi7uD1VYQs5pNV9bxUjRiCosDK3GrcG+lEX9kxvtxVyJ4osy6dV2fZ2Ue2mXQrX2tldhl
4087I0HBj5ZCTdRKXjx7qblDM/7qLZys9RjnWZjG4ZfT9gLbCuhAxEoVgja2G9Arr7w1hJlVJPAP
7CNyrvbUcu0uKPHOsNJO8w1AptslTnTEizrlZW1tsrM+4HmErK0qN/MfqNrtzsf3lVplhjlRRWSc
SvEIyJZxvoiUeMxYOAfHrVHqUDID+BJQUOKBofapytXWvs+NcV1/n3xya0QWhYgnm6nOJ0IreIkP
f3x6Swcewvkcjuaup9G0qG0oEntcMpzadmuBBBpAAR0crkeR/0oy7GeS5o/4nhtgAoydVs14Mc9Y
PR1/cqFnzWoo13BAPPiNoXYb6oTIXoPzoJhOg9kAVzQGFUkPEQWVh0IAt7xIpotYz4hejqfNxq1j
G8ZrW6S2nb3lEUlESMG6UBZtgrnsVX0wOj/Twl8l7pLvJf300gGPViowfVwscDhAQSLJEhGCJ6W2
vpwquGr5WQ0GPagkjyOkdQgQt3NYDXAT7DngUfNY65QpiyX7LlxJOttjU46pSI8TLssCL25ofrNn
+kXMk6ozsHLftCvyOAv3C9KqHz/5y730um83PdEA++1HOyq0B9uYAgRRW9fpqgxDHycX983fjujX
UKWqOUyJBc0rH3/pzLX9Sut3At0p/kF72EOaHQPqyI4QCecjf6yoOeFhN1pFrNAPtwA+RiTnQT8b
Far4UznAqnDnaGl+fMe6dUUr6VC2GQ+0J4LarNCXmq8FG3zE+LzLLMKHqJ6d7mF/9NiGKFnmKrzv
Jm8JmpckFuq/T+WJD7vyWGJgemio7b0EAMR2s9vVOGzNxvabxq4A6dZ9qUpAFqjeToJi/rFsWcTW
sjZGsCWH3Mub3wDgPOAXBVkmt7AA20YVi6KPsfTXtGnqg8sTt3xFOBjC+/11/GPdKgk+75IpsJe/
2LUvPfKyeuRmSkF9TlbBoPIVD/3y4+gdnS5uWbDe94ZHtcYm5CZiGuCHMmRn8nOOW9OkpSyNpES8
s7aOFigCJi6dgrDJc8dINdV8q6jQJ6K54YzjykyHLCU0j8c4SUch93pen5ccRIl8u846Kjd7kXST
gA7+QArqoIs8YYEGYnMutJ7chnP9FfmH3h83QdoHFnhJ6HbrPWEq0YmXKfbcQ80nRDDtIr8Jg0DV
mK0W6vOC7YFWA62fIAVVN9UJ4UwYMK7CHj//u5hzQ2VNQQ3fpIA7WhnkMowLeAz0PLBsYcZrMeX8
pg2/CzJ68Ox6cn3nrt8IeknCY3a8oxNPmfF4xj+l3j3KbDktSA4oV9+ufO3eCBJKLXxNkGvC5nsx
RP+x3gjbgp7sM959R40/KBZJKDieO2nGR/6BZxetd2H+NFscTE/WJULWctwRdIdVilyNtQVBoT8M
+mWiwXpH5C0LwgIIGueDP3O788GdlAmv7zpfwbgu49+g1SLSJhdPnxXAmndUtPMHFwS/khOCfHeb
2xwqgSS2447S5O90tBrWGjW3lBHijwrVT+3G7UOUMDialWC5GGyckr7SH4un902H9ouTCD2ZLunY
TU7FH6HDnHlmZ2+O+oXwFsEHqK+Os8pJOqnWKdwVeVCSQzvXj6J5Eyxv0O1nUVe0hO5e9/p2uSBX
ztsbKjFbDVjHTMsm1wqrts5Zhr/vgsedRUAziby0a8goGGBtB75TT25S10Yjj/cTJTR7Ac7JngyU
+TWdGxDv4TvmI/fog/wwpLNYtLUnkssP9gixIj+GDrrYlICIRZAlvG1a2JyW8VkMNAF9EWFUvarc
9p0mMxPSUjCcJO3+vszEHXw2rirx6K6c0A26SnynqBqVWH+HAgo9zfnYAwMOeHTjqDWL/SqNx/o0
r5yBOV0jBCzobrJ/qaU3PJlaqyZh3OG0KfmFNRhRI4oYiPjW9DMZm5LFivknBfVS9d7oJBIAJnht
sfwoXUtrd+Mq73cx6rCTZxHPwe/qdKZTOjGs9c1F/VH3tGNW0yT0S65jcTKousfHmYZKsJRJKnNF
jGz/qMyFC67mXEsWN8dkxFP/gvVYaxaiA2Aegdg6nd9JbWpQfhRHuhw/aQmmXg5SrHYlHbatPo8X
TIUKM9pUwbGG+zLyZukoRbOg9ndHm5D7sBEo/hXsQy9N9Hgeuen4VEZZ4UzBSdGCgsdPDRYtp4As
4viQRK/a3xXxPKXGV35yU1/bn/jMuCAEI1v/ew37DW0MgL7OiZUFcQ0l+bo0SXa81WwadkHWfSYf
rq0lr72eC03vcneqVmgLqeg0MphuH7Go15e+I+TqUOYDMSb57kAghg8kvxa0Z+YDLx4uj5H4Sok8
lmMFOm/S4WCYKDhzVZ4PFeB2s5RaU2gb5zpW2WPXJIq/PoWzFLYMiNaYdU3v5xB/JOVXnWf+H3py
9+hrW70UrBDv8waTA4JWzycGME8dshz6RM/+rZJqEDR1RnQUIhcjLzktdv2jslJimM5qPfXWvP+8
VOO8Tf7zpA1z1TMxB8TCNtOA+aiuNeYAd3f5ptsUIf3/qWhR1krP92nvaFL0ynnEWgTvwWEKuCwd
TX3VIvTaxl0qw6w7E5I9S1bi/l8p9PRQ2UUJIeyWKbZCGmm/WSErvhsf/mPGHGL9tNcJNAdTVpKW
qh2dU2CS8vcMV1pv7+oUwdOyCcpgXkscCaFYgotMipnSTvGYSCNpZyIxu3gy+v52IUNGD9Vh5Hxt
5DH8J+6ZVB/nDTCm+hg/1fNyV28RffmrbSv1aUaB/jGhSgHAJhWhaMTWg/YMUmsLwf8cno3gThYH
bFXuJlAMrkRjps2sMqx6EWWecbSyvE3l4rlRVQrXkMLOfFq8h7II03hbkFdtSDYGthH8y40uizUC
0pJowKxn5flDo/G5+uLVGhGCNEZ4KfAqnwlOVyGFTir1aYs8RJo2iNLO2omgD5lXi+5UNNQ45MBT
Qgcx9oAMbgFKPivPUO1ldTjS84/YmVJFW4DecpRNTWen4u5zxWqGIh3UnHoG7z0guFG4Hga/curz
Tymcw6WMcchfVvZinKEvrp0iqd0h3sjIkz8wdwloepuz9jjVvaaWQVoGWVPcYZzoNKxEgX67/sNK
KyM0A/3/YJ0N81MZXgPy74Pkag66EIcR0wesoZH3AU8HxGpe9XUI91OtsZdmJpcs4IPC2pFrehQO
3/JCLmCAgEBykMKX9ia45u9tF2wgR6su+we9B7X+8Z8jGqL5TPqeMO06zZ9s3ibi4cMVt/0BRlHT
zxixnEyVTAP9by9rz167hnmVxwIVTv/WsX5d3Txe9KWz/msAUh7x3561dQetc6elFkUn/WUMdjU9
T5JvQnC8YX8AwT6h2IsHvfhEId2fCXBEbhuZ+CnYSfz1l5juoSSTV50bzGEOQfzbvi1KElX+Ogmq
mLVcMSzuz/SNfIaeqU0WzxKG29QVhQ7TptrRG4gsigmzCdoUk1Nt4WwzwGqCAi93rUSuLp6Cz7Hn
eGFNOw/0P+aA649iOr4FCeM9S58VAuFbYDxVtNkGuGChLDo571jEZqT5jpdMYZ5W3/DEZPDAFKmY
zYWz33AwiHgjFkAa5yiiyPyx+S6TmYqxFiZpwgR3x+CP9kgajKj7ub98WoUV+HmbMewk0u57WJ+O
e/3YUpvw0h39/ra5w8zOsOE9apYwGGchodozssBm3bR4xdbWNgchDrH60TYEBxQ7Fo5lEglE64oi
7rsrQu/GQWyLl0FQf/KuOTvODQUymBPUMwvz/jbvQyVZg2/nvk7T5FqwNCGFICieu63MCoVPXWBG
zsuBGGEXLNCynzPJ2uhGUgKgqqbpiFL8u5mm1cAFOGOuKI8Nh7IpIT2lskZ5Wewe8Utvxga8T1BA
PCkLsU2eU8wZpcVViK6+CFMZ2gaduIwd0QVdzARwUir/fAFZlA6YCCCo7Fa8rkgk7yvj6WX9kgBo
3iyzHpfcN3VHVt9tzP6t0stWjkV4wmRq2Ximh50XphphhYY8YcHLLQHdAxAyuMqaA6qvO71L3FGq
ThMZd22ifGrKVy37dZonTSqvsVZb6bu+otgw4kOjGr49XSLJk5AZokAADmRQjW7ryDraabvo+821
ik1vx4LClFR72Hjyigwb/VQO9MWfcn/MIteNixYwqF0fubzkOHd+OXf0XUvClOBMwZTHvpJu4z9o
cmeaboJnWgRxGJUCu73WEtS7PUbhCEj8n27NOJgfiw7hzeo7emKoPLGWWvlux5RUhIZwkBInTNxI
9J6SXACcnR7Lq+TBLozCCb6wupvQNTSNL/JQBPFX4fX47GSSCudb45HmGUOdgxnEY8XgzP4Ibgug
pg/2WBpQoZpDFwdDoQKAue0wyfbYILoAzNfI0arS/b4MZR7ZaFu19fGqRniZa6gXZYPPOSqg0Ico
/+UgrXbXLmaMp9Ot3QRZ/dkjSWvhPwZQ/7BVUvcL8+wQUZpPI2axBs2OWaleNffXpWbUVrShKvC5
jSAihDIPYu273Bl7LcOEIS2gx6YukZJg2mQbKTQPBu3CDwFcakx4fJalG+18VZ0xi0mzyt8Jy91O
pQ9j0EoxvF7xEo68WDzT8gA3WVIUNaZTEjdKet0mTG4RediBQTuPhq/VCdU3SdD9pUvHakZaP7cp
mSr4GOxE1s+W8yi9U/FJaq1mwnujaYojTcyqvxUyVhX6yGHY/BeGeEgmHpD/zhYiUKE9fMeindzj
XEnKezJ1MNbmx2/HIbvsCWkRBrsgJMZR/J4LEiD9FquByiHIBypfUhE3uDR5voEGrTcOzuDn/QFQ
6VedhF/9dvNNz25vd7HnJ1wK6cWiRPoj34jDZFfNb3NWql1IYffPoR/dVzwJuY5Ex/a58b5S7dqE
OlCBnKcqyZPwWsPS5VFBTe1uOZtmL1AnNHCSt0/y/9MPr+D0x8a5n/PKcIKHmZOFrPJcR/LlHqgH
xwkyYh6UFgcp8fXPYwwUZ+s8UbhzQll+cKytZCQtZoUIvbUnQcDNQlIFwMi7wZHhAANuEo/wHm6w
sfFwn6YAx03RRpW6/Zfy93CuQkgR2mvKB7iJ12T1fhKYj2GTe0BGTOfZUtDCqID7Z/fwUl/yWoQP
FNa3J0G0KiugzjiuwELZsZOirvUpIqY/VETGm6l7gw9Ad0xjNyMQvQ2wVBjILXY+4hrOt16+Y7fN
U4+UXFGJ9/9QZtZXy6jtrC2Fjd22BVvo44YC6pCp8mpuLUDsrqfGLs46PCKIn6jUaNLUtCUzc2mL
orvgnifJzbCLTI1Ob/nCbKN3DD3sLeM8/zMae6FMVHq8EBfncUCQQhGv5CeQ4T8m8cZrfHrbQPLJ
x9kmm+Ht2nAHBf1WX1UtIz5i4OtEaJKG0NN5XnHd/6OqiNNhqtkPE/aky+q6W7+z1L7/CdQDIzDu
7uWgqr8io9YprDpJW9Z6KiJ0tHxQEuoPcOFWkrBxATiSvTqGwvb5y2NCiiu3kbklpnyOFv4ron81
3dMWoXP8yIWmlaItfS+9syCXwdEr28z17DOzDyBSWQjbWNtm6xAN7zkwhH7b+F16UlcbTgM7vKSB
zXDMTzrkdz7uVALUANuY45Hc4tu7qpZHE4/XfMfEpkeRNBZNIxa14Ljky5xxNP/guH9vbwyWY6FV
tn5hjxB2iO2Uo6s38cXtnIN5L/6p/njS4m6ANrESta00MIBaur21JgnD25CKYwe8/Bdiu0Au2lUd
eIa+wCSvRc1bxE7mSDN7LrXMT6rXojD1zKeJKmftB0ztFp1AUhdnKElsdSju9+Gssk72hzOeCLcG
Pb3fpS64R1/ijV8r9TdzkLUhSNrR2g4oyxn/Bjd4zERawg6ecp7/jk+NyfBX4FN/9LW4vA9desXT
i3CXUdi4UFxxDhC2WeYY0m5UTgVlRm1P3eKck5KxHnYfCL4ZNKDY0S6fz5pRhhecY/kNHYQZQky5
hwFfig1MaF9alxKu2eMDifKzaoJLAS/gl4WHnoystajZm5KtGqIRyfDr7QVw/8luNNVCb6/eezfe
8ibVDHxnDzWPBwej2V0HhZbAVgNMAirhxeAzCb32mdu69te8zkdCJqzKNgQn/5vg+M9TeaLivDHf
Pcw83q9k7FempwSeeMcPC3b2uC/7dX4v+JsIflkySXJxIFryfX9++RrBkIAweG74MLl0ekkg+/0H
dUn/9p/mgpjuUP0yPAFSKyM47qyRoTLCfQzDzlt4dC794YovXqbN7PHjDbXmxgLWuhq8gXe0Se82
+97ilLsPSV5sYZd6cbjSQwsmcKIRw7Js1zazxJZCXIHa2daOGNtnfnZ4gjyhvo/aSWemT8YlmNuA
e4mWMhDwipS1GpMEBjhLMJbqJbbsRoAqpYxwEuhf/Kf8oA9phlZBWPp+vxlzbdMdOKAAtQCcNTTh
CYi5tn9L9auxLkmhqEkTSt3D/wjbvZTpEhwA3KEsM0/t6IsR7VRi3wwRsTQadRLF1mN0S6rmeaiA
WhBclb3pmJjLwoGJ6IntS8NQu5XCmaBKwdo3V7MRqb1vGkSDjuH3NETCw2CebTxJ94LBsMneVf5j
NdZ2jt5J+M2w+By6nJPWlr8WuQpP1bhaiwtDaYlx9rIV8eh+XAMZYG4Bqe+m2xOk3pAcXg/F4YHl
FslsgaeOLRZsvYa0YndHOad2D1s9NRcIVszBb0Dz7wCtkQjEUQbE7F4GqMVAdle/uwUU+NaEBFbG
GqzDsdQLN3id8RsfUeLl5fTKR7AHQrvjgToH+869mco0MGc6KqsyTVed/w5nR5v+It76cPEsgHY+
XvKpffO44V/WQoaai2rlMFy5yK3xggYWSDQFNFbO1cNRu6kkuTeZs/++GmidrMxC2daH4bQqdDS6
M21nyimIb22mIVHaxRYEyszASVNgKu+QjUPjfCpsBfiiNGCo2ZFJpPPQK+mOI41kX5MNG8YP11Eo
K3Xo+4GSLe8MGoOqQVSMjRhk1xtuVcQMwevyQvpvJ0Hwe70kPN0ZuBU9Ax+pcM+pbql5pIXMd+3B
sVaHmFiejDZMB84U7POQiFGgdjAisIjXBbtk+oHsZ3TfJDuKg8/DIVa1f6jHfUhnfUSLqO66MxD5
NVJCzzOdOGH1oxM/LNtD5knErh6IXo2an8IQD+BdRgeQWYCT3r2pSncrYCVmnBumKxA/s3o2MfnB
YjK8d0DNQNNGtb4sTidIjJhmG3neEgv6J7VaYSoq51mVUCPdz9LmyXj6kXmq6qHiFf101xxO8I5j
rvQupngCeL1DqvmTwV2sEJWn1innrpT67Ojgjr5p3L1wNtOwAyljTYCNhpjFsxy39rj62ac9ZuK1
GejTaGDZIcCozPX/m4iwWV3BEbV4ebCcfeoSbOY0shiNyXDeqz/M23vX/WafbzunHvZ+samqU012
FBwuT/aGg1qZOi7dlkA/dIwJQrO42Nfr2j/NfgFzv8c/xrKSqQIXY1KXQYTtR3d7KTliI0VgWetQ
l5+kvliowqHDEi8iFEmxoLeM1RViblfQmqTWwexbZiV4xPsChuLkLzlSe+KgkeToNzFRmjBdzh9W
ZmjBaa1dAtfB82+ypnlvBektfZTRPs20ReCaKcjRvzJhD+4Cc/e2u2uRiCmrxbrWnXHJzx3q0YTZ
cnKegNlJY4ntGLIPCmiRPQsvRlOIknoRSPGGtRMwndok+zFPquTu0AkSZidRM8WZscH2VdeJeG75
H5UGg3PZIkiy9o90b3x/PN262nlgKxElknI92u6q0aHiZucIqBMu2HlEr60SPGar+gNUS04jnEKf
AXjg6nTVdG6ww7RdCet6E6RpZdzv7QKdn5vbqVQ0g0S9R3mHQVr3tNhQuJ04hqCB/a6Gb6L72qiq
ME/2Q+5RzvTFDyw1BNnC+ZDgBikcPbGUQzT7uBJPaab1IeNQo8kamtmZ6OjesU27ngNCLjV/LxFT
ad30WoJIaZTThVeqWuEJEep5xbrYVF5PNHL9Zy6O/CFHQ/8rruaCMNCnDM2oMJkoT3RHDB6Xar7e
nNvfqS0tGM16Zv5VqrSKyShBhAcQ48RnY7Mv/W63UHUa6o6NT/+HAgkRZPUQkDryX6OIgpn18fej
vR0O1TXtRe/V/CMh8AktMwoRbl4HL1ksLyVjexpK1FmExzPvrrRalWSiYC7mei/YqdeQ2P5175TS
BiJyTpoewhodq4BcPyiRKGWxhlTc0awNXBSh8pp0pv3xa4k9Fcrp8bmRqa+F2GZtVcZw9IL9CAPg
oG+EZLSgqI6t3T5ScTQIsGtKN+lyIQ+H5X36UmMKtn6ynMS7Z0arYIqLoThBkPHd5bDlEJAbK12c
nCohqgShkrFi0Cs/hVeTJq7GuEYaIO29IU5sPnafRkQjI0XIKvVRSeFAxNbx+0WLgKC+JnxF68Pa
FWKBC0ffiJTqNvUQjYGCyNvAf78x9pvYISGV+qPJIEU4yNduAsVJoi6xPYygghZxIYoW5czxlpGE
z5eq587OcrHJsJtgIDzSpL8Rw2p5RUTEIZ3v9jw5+3oEHzrDyy2mh5dO1GdIe/CTnnQVbtl/V6VW
0OZzdTX9ic79RrERrROnkwylrHLzQh8gLAFK+pUKIwKTaYSObQVdBmhADP5K/8Ddju28MYJI1uFG
HYDO43kd/HJclj8gLTeLby0Vf1+39uppSRCW/Xr4qEfrm6g5FpfneQhwt9+ZSJ73cPe7N4aXpwZa
9r7pl3wUAfH0Rq+G7nc/5mQOJMHGkV+dOCKH11Btbt+Iru4yejjdSj6w1zN1I1taJ9/iSN7AK5Xe
ZqwhXlQkw2iVauS0oj3QKZQnG2ktgupsozZdja3hJWCQ39uuDhvqMIyyg3T5e8xMoR99VvxQMMix
v1W1TlMAClfOHs/lG7zLppjlFCZezQFVgPGqb+J0jy9wgBuErboL77fn6biHUsRIjn8pbWywW0+I
4rYNs0rPqMQeKbO/P0Qcobu1KgjOHPMwBIdPriD9ZBp0vr3/R+ufK3x5E4l/GbzDWfhm/3oDO981
GdpwFDfmwbFgu8CZEY8YJHomOXgwnhaussU120TLlU//yJmx548ys8MsLNScmPKFSwzOSZIh9VY5
THRmhw0Lr+0KyYVw2DhMTSWl9FCFvIFAIZlhHOr1AysCPe1rgIevYRbj97usrhFVELaMxemu+QZm
ZoLCsfaQ59HXLQDJWLqx1KsK/JZ8D3ttQVnd1QmOfoNDlzagr8/pB8Kjhk+TY2pW/rDbHiVGp3p1
ENomjumoCo6sMHmE5sJNPaQV7AgKBLiwJHH4IR4TcSdCCKev5wKUYt4W9GnOTQrOCheRAY4V+3ix
xlylPvoqEkHrN9iPpZhRrRAxQKUxMuUmNuxdeRr3AhfEp6MlR8SeJqAHo+aON74hofJI2xnPRe9L
pHxn/2MzbHJgCS+DhPrWYBoKiVAXF07qt1dNDPNKaW74YUJ/SoUHO1kGowLbvvmsRwdnPHQ+gOfR
8H3x97IeXZUnBcZzG5HjxlvEuNsjdagIIWBfNpihoVPtq1KNNM04mi/rw9YimDbalxpu1UttruWb
V6IdgXUO/mb+RGD9GduqGRr3t/WNXfG7p4U2BwVE8IiemgrWs7hEyWyxTwc3EOQDasuuwOAhLCWh
W4fnV8rEBKKAEG5mcaY2cqQ1SycRkCxdzTaJsECYM0sXjYlJjljk/0c7CrlI3HSBn8CFuYOnqxS6
rKlTsrLN8IWPlrJBNTbnhLHZaMUfG6i1ZNPV3cNXQ5hNJcyLfpEYLaIyQaNARVc96tCCiMuG7oVc
zUC5Tbg1fYhG7j3Lcf+gWQojD1+XPmhRP9Xwaa9+hRTyZrXJZuqY5/wH8SYv8ECD/UVCqYjVb+P5
hF1QU9+/uiStSUYdHnI+1YfW8CcA1A+JT6w2WVL4f9v2Nq6vOTYB+YNTe81NpRH/Sxfv6tWO3ylc
RRhIro1IM/B4Gsk7DRYVd7DKkklf0YR78DAJgVChkht3mcJ7qmpXrImD694p21GFpYZJb5TpaD+S
bqQNzGq5zB2GvLp9A45hInUWAcOsCk83GnqufVHIvP1sSYNBISAgWDjNMTh5IMmXTl+cBqQlmCz/
czWDCKfHj9aWwJqYHCH4S0XD4YS/Dbs/f1341/uGc7WWFck5YD2eEQUi95b2CNFUCnd5P3K39q1t
ZvfMKJ3RIymwq7Tjt+FxNbh+DrkwmQREzwIVJ+w8CrTjg9E8pML2dqPCXSudvaQJzMP+g3/rPCGO
1nFr2g5UizkoQE3RPoIMT+j7eUpXmwSdTxvbcUtDBulB71lQqNHrqHF9+6O7vhDIQ77LPgmZOplx
Ifk6SJDNgr2H58NtfEYQR7euwwAKRudW8ExbWgTr6m57HVaIctiLaER1YDcel+lmUylMvLILswFJ
HH7eFRPsrQ/sjHT64ntqSk+XqEBDoTVaAOKuS/LpQ0U9Y8DNuo9Oi8a+L9KM7+Hl5yGObjEiLOOh
foSGBLBf18tjh0fCW5NRuj0pA6lYQOCYfq76Td7rrVZhAMyJmp5pcn0sS0prB7mPSMDufb5b1pXe
EnTfsBVA/V8aroRk1SvFwLKxe083hemH+og0kG/4sy6kxuDk3PSHPJiED675JcoZB+N6XsvDtfVX
PiZcdV/OscOrAE+pkwlJUeOqo1LqluqdbLqjSjC9/s+feGkfGo/1FhvameV/6KCkLMdjfGQZCPjH
zAd9Urje0zu4joVogFb/SsCaYmMXAs09L0MMsmTGv0mYp/I5PgZoIwkpCb+GYevG/pGrK/UZ5rw9
Z3Y/qQo3+aMiUABWHD0pp5bMw4OrAY3XLCdNe7u6nE2FkRcYIBEnEY/NuqZ6/pDLl5QIAYpydkCM
4QX9qXIK3CpfvwPFSN/MxQQ4B3uQhT3z7wWmStPKtwRv2likfW4cgnnpvmBbS3pLyWr/DEUxZ8m+
nmocozVx9m6EIRrftNtYt05I43D6MKtnmIgFd2P0cZGt1UHifLzxet1vb1YEpgFh6VbdGFJbi3lI
f/kPK/bYmBCBmX+6GF/cnh0tVUuy123/c1oDjp4hFdjQ3RGjlKeBDQS4WauXXfs0NoWIatslUihs
ZMpgTNIGvPIRkKYx9lG9gQIym/a9LeosAVdGmyg3Iw+NkSEVrqquUm0ikL1tPxV1IUja93RGnTCh
vDJAlrSxA+WGzqBpLU5WcjfShOfYaSUs2SiNZw9PCk8S/PfHBZ4aBp4HuPvaGwGx2z6/cAbHKeFi
4TVqJcanDYv+9jS8u2i9GcfLTiPVy6A92PBlXS47VOjjjQiVJ1PsNPoMHA+18GekGRGhTmfbqilq
EcMwf9yW9zXDc7QBpVDb90HSexwcNqU7YEz/MRDhnhb6f5w48LbvKyxF7Sp5jOXEd6Z5n57vR1QR
lyNpcAIZoj0b/49c8+ZxUGwoniAUMUNKB273il7DSFb6G0reqC8WrXgjxBE0xrD8fffx4Bn1IdHw
YnvdlE0Z9SbxeokY6O5mhvcFtB0JMtoouMhnWSC1pPK1nFEj6EkL98PaLyoygxjfVQqUmClrXkID
USM0LE+jo8wG4BDXfunn2+dG9eJSXVHRf2/4HspcW29PU8d+3pbK9LmySsZTq335mjgQgIukPkdA
iFYleVz+EA0mdnMPPinOVTTQPS0Q/ruHKvhDGpo60lPPTSyjwKOAOJRF06y9HD6/XhBBL/OmNXtR
3UD15h37hKBogmYLOBeKiUKfvsvGtCI7j+t0Rr4x4oab/YKFlZnO9EziwhipMF4/6AIx33SXmwub
DJSefFFlKtX8CmC7bCt/6T8xR4aTRaxWsRCVGKelQbayl8TLFV0F387IfgswHRQhBF0MXelHfsMy
yvvZsWzrkpEftRfX3JhUPTnN4aQ1Pv0t66yb6MQmkt8eiZgN8f1iFjDG9l7VRTUdIDlB04/Uy5CR
83q3/ikAGt5gZoYn4D3yyNBQI9uh9WUYDYcjmupacg3QfN0VeVzmfIn9lzKVEDRPpztJKuyMHKU7
Vlj48osF3BoNzwWESZAZiqLGYOBc9jnyXzjKnv++a47Zppd9p7lt8V55F+cZeRAyB/w7v85rJMmr
HomxIw2+fmk6kRoq1kThyHeNZXVWNyErFjw1CHi/zqAxsSxnBN6bieSRYK+p6R9mAfdOb13paYi+
NxTPrltan3yRTcXLHnNIPWYEqqcvUQahXr/4eX3uzF88qfajzFsrSHG/LN8rygRRNnk8GBatVasm
LAA7pR2z0Tjl34oybsb2RxrfbbW80agAUrbYDBDBh6gBF1EjHinFWY0xac+8tZ3csJbuK+/tHX6q
n2uteWxMrEguq1TTNWTwJ5+LQDfkmoIIf02TScvxdsOSLuF3ny7kmqg+3iOFym4ZqyQs1IU2IZe6
snC5RsklH1YmHE1gnKoy7RdoKKfAubdbMszxNRKk2DVWXVqe1J83SXk18wpvzyPAIFzWSQQX60HR
XRKhsmx+x2+h5EF0E6ajGTgPoZ2PFgu4QDnpaPoofgWhVVGARONhkHT81sDtRhEAKQ+j1lWu7f5D
jjvxGzg2NLeGpQGN+EE0bB0UBdMruLsO3phEKLGgKI95JJtFUIP52Rx3ZWA1XiK9K+V5yK+me5G5
MnHcCTblTYpDUgz4ViINmhEmtcWSQS2HGI8ephgsboV4B84dGVbkPyeLjGXlLE8bU+aJiLGkX4iE
gRIHrdSnZg5R+2ob4hfZuk/7Kn8T1+953YaPpgIAq5M1iJ6SzacsYl32b7vxARvNgj+iOy2xQksI
4dywKezR/2xSf40ijE604l45/wZIxlMGdayc4er1noS0q2db+0ndXdrcgOQhmgsdPL/JxejAGwp7
QrcOGtQn0+/WJFgDqzStjr2SmxHTyvZUgixgH7CWhbUJgbwlcCrGVGqcUXuJIvo4AabldS8h+pf/
gUwuQOpIoogvZj/YNY//02wLnpDEeiYgFQF90uehfUsHs0FfeAvxLUpv09DIOSMLcb9HFEgmWM1O
/t8MdD9qNZLNNKbjsFALnL9LAcNuXZ7kn2VehdYVilksN7WzwFlqiLkZotm1cTZU/GjRGEAYw5Eq
D9wob+8TedjwlL2FXp6Ua0aShYz6linb/xtShMZ9/ol9tBlSg48IzidLalQkCVhoB0ox8MnEvN9b
iOE2IITOq05DfNJ3QPzoXVcdAHTd3HgwVY63Y9DuSokweaODeiJZ9En41uQtOQDN+D04f4E8AyEA
rEmgw5XJjm4dJLOYNOTgauk0usfnwu6ptDh1mGM6Q5ygKoZesVpby3HWX3O5r0HZS8QOFfUkk8Z/
JyVfwbqStnuTc7ygAS9onSpTCmIywWcqStorut/AQATHeX7y8GuA2COqwGxubeg7ZA1TAiLKj1LK
hRgjmiYua5FM5wdBUdkI4Von8THwhFnHo+6vnGYvPOy0N1iR8Rittwi8eqaPjs9GIbG4iOFwDSUk
BnUTjwUJfErFkHhtUD2Q0iuq+S3qvHl9xcbLPxYsK49KpPRL/Ctzf8fH+07E67C2AhXIPryFlLWv
hPH226FlIWkqCMDGN602neH1ktiueWcHhYnS0AdM2jGdC7T3DEdbBLktg6V1H+3A7yyWv5XvtAEO
l+3+TVeWCBxp+13Cb3XYQ8YtBQI74HpLKSV3kfdL9zst0VSIWKG8JBforX+38+AUU8kU0g7KAHzz
MKU1ZSNJhCxgUMn/XIz979x/BddDmU+Ucb6sKg/WJixoWrv1+Q+b52kx18+P+fDq9GwQz4ymMS6F
0O/ZZ29yTGvEN165N6b0k1w8myuXtOeXeiMCu286lCtM9XZ6VGtoAj5XCYuELvWOVL9YutIJK9/e
J5yGmNNsd9zgeAbhmQtj92p1vdUZMf2fQiK80tdOI827RA8LU55FJiA6Y5qNe8aSa5PqIfmpKCDh
rE/fR+dZ5AtUKkMKh07bdjKNq2Q7bFPMbFh9c2VvtNHetJhzRo9SC0h5JwUEVX9cIG0BWyy99Aqs
NiKRm+WZrmX5oStVK+Dsm/30h1wkYXbDnVuO7LVQaHXwFzn4uGKkkC/Xz67KWC2V026csavTqnq0
BKvdhY8O9+q7a8RJlpK35aKZYxrxUrpq9RRC1t/2gj89jtaXL0kKMsPcWZd8aJzYySEg3MmsuIJj
WgAMNsCkQBs8BWJ58E8BclVit9zaVtTD7USk5IiQXLDHMtGxp9eo7rS15cbZwTpZPUmJKDTohJ8I
orDV214rlcGMEWuuA1X7TcRNoJwFpDCVKaqdyhDbk40q7LqSIaf5QfITG+VYv/Z7AgZ1UmsE7p6b
FOdaA6Mq9P8j4P0O+/RNtN5iL8WBpl4nAkhVnFr7ssxb8swM3nGs01nOLvszM19AbWO2VYKLhQ/0
LjmczsEenEuhdbH9X1e4hN3K+rRxtSJlqXFJ8xRF5iFFjNYVFOtF+cVvAutcVPOVWgLUCWJGg48k
0P5nebfzMZhrDtrat3m6YLmYDm7VQB0yRZKQXG10SWzRY1xLjZ2NvlKgcMqVKiJOgP6a8H80rHtA
naMp1lT7ahFm7TnbThoesACpKlo0nZLBRyPX31zmGsEH/ZI/syn6khd6TwNC5MzoMRvZDymMCruB
+df4DYgdTonMSSkdW1KQ5AEXezsrI6YIRIfq7gIBrOo02xCmrT3A2d0G8uDjrU4rtJFTWgfm5PUU
0BDBR2e6EF5ZF+XzTY91Ii7AIqFYSXhwKdDIb/6CDzljz6/Pke67/0oLxwFkz7AuoQ1nCRDjoN5m
meUT3EsrRK7H4KuTV15sgprnAnEgq2YoYVz6sFX/venfA4OflX1VRSty2h10vdnElnDbGGc8Or2P
xAGEoDP9qwB2nrFPJZnn9RIeMqmSgP0+xRYc8JFvFjmTjz/GN/7laJvai7/ZrL87bdYf62OOb2rh
BJFrDMOsSbNEp1fEMn47qtKr5p0SSkU/L9aLwPBe2XKC1e2z4YqssqDEWuMw9Tk23t5Xr4TIJDRz
Ek9TVsvvoo+6da9YTbkAgVz5BQlqq0rhhiyzTJdxKklaYpIPYX9P6wm6uGMyDSVkLIcMt2OjAYyJ
D5pJXx3CvfL1pulfJMQzhYUZMqcjFGl88qXnF96Yfj8Mfo4ia81IL4b9LAwSFfbNgik0Ech96kv9
cmblgOAwRmemVW0V0grp4y0Ze17Nk/KZRLNQKBM7YGgRB3xe7DXL2Gc7uMH5YhMYZmxBs9I/lpm7
Db+HSDaiH+qH0bH/hlhdwwsnfkM59RPHcLSC/8h+JGJr4l2FSLotUfmQgxj/vMuOMpSNDNR9OvLP
MYHqzWFVzdLiQizGdBN9s2ubYUmI9kKh5JVeb1/yjZUusyJPMaMHTklBxhZXOSBysgUCgd2FM5Y1
pkXFk+4aFbQDREHiG7pdI0nYfd1cws4MuXhIx8SRLmw5SbifgD0ddWMLuiqH6FeA5KfTkZ8G2dMB
wWg8b0kWrVLAhdwvEay4THv2Z4cNmcWolVBkLsAMbw9HaeX2uJUGSXLIauWeOqy9dT4k+9AEzBeU
/2azPhbyUqiMvNabgdTwmBXMIdIEFgfCvFoh4/qUptakDHwIE/A8TvQF1+OvvJCp/cKZsMlDrLVa
0djKn2cAHLPqCP+8kE8+CZeIOR02gwVXn1bP8GVAoYBQIOAG37rjg3NVWv7nlc/grDwLOV1c2Q0o
Lk0VqCCBhgZOnMWVDcml7Uqmbie4ecm1IIehYx4ZUX5rLOgV+fZsPyk0Tpu3tVzDcJVTRFhCFVfo
/K/aABFmbJ7TKFt1y1c5iSqutasbQad8xuvOdUSJ8LNeOUBbhrwkoRYe53EXCzO0BiMHlJDI4bOX
ESmHi42mRY6Tdq+6vvt/t+V4W7EGZyw7hDpggmvdGx+wcU8IcqzKU66Z4Z1G469QUBPwUHr/JxTp
5Cv9UKBejbfIDDqV8o1lCjoaHL3gX/PQK1JHWD7qwYkx9OR4ONo97672u+l1ACYKwnLFa8SJNk95
VwXoumF/NvMAnjVCEpRKKbHMIC4zvADHTN5PsTXh/p6WeHir+z3HbS0wgvbH3kdtfI/3Hy9zqDIn
yIn+uftDRdQb7XR9sGPoaBD7KHNCqk6fumM/Jziou+rMwbGSB38TZqSD8HnJy69KXAvKkUAwPkJQ
qcwsd0I7chthsfM31y63JJuI7WCJRehuAOVQ+U9SY5cx8i4eYNKBV6uhiEGnk3TJ874xmQXD7ZXZ
D+R3Le38jXHFta877APf+aVYisCa+xywHF2Xw9u7eCha98IxFpccgDdOc/ZHQ0PbPmXYOr3PPxf4
j8LQhapEXB4Gqrnm9mjmG8eiBm+V/k9ILI4ZIX03IbghgeGTpOgSTPXKlcilGTpRIipECsnjpevH
c+KVfPiV0XN/FfAoOyfq9iwUGtaTImy0n5C4IZisqv4IZfRD+RMx2EIoyY6MA+hTesuor5IbVh4m
Koe7oYqxC1EyY1Wm4fbCufeoNOXYR9R4DhfLbqviIkUyECgcimRfMUigs3hU2mIS545SXjIRA9md
dZxA8/PxtZd+yqe5vYpIzwk3Whb6Y7By0Jg1aIvdwE8m76YwLEtJfrxaXUnVsDnvdH/qBg4AKWlL
Qk7NKLBbdTVYTdHzD40lbprSm6Cz10rO8FzD7yBwehlPw+E6WsvCLLLbh7P0F2vyGlBIwoM7q1i2
kUQkaZWPZ4A6O8vTrKY7XS0xN3zaQ62O9lfNo8tkap4n2Nw1lnjKTzK4BopubmvSL2u0Vsl8IeHI
c2ntH8d4CyTVijDuR9NF0Qm/9zCAZPrSRJYJmNW5IN+b+TLkKVU0WtvBQR1g2pDTSNJ/ebwfoBkl
WYLVfuUBFoQXSiXoBjYUK2Ro5B5fuiqMMpaGdhpI9krC07xMuaF8XKaCq/+/1nd1ANvwkIJxLCdJ
rqQiNR/HTkU6SHbRTURcjcFhF5ylrQrmqpUEEyK8ocgiE+xFFL85KRonBEax0AZZ2eWdqxtLFmOH
x8FWW0LNkRk2rJ2nq9i0P+mlbuoQ65kNMReUF1+Zx9rXwHAhjn43c+DP/gQyJr8g24fzfMFK+6jo
H2Ku8vYbscnpd3pA+0SANflUsn4VF4GA5NULHMxiPfq84sd3W6DCmtKGCKKwX1IHtlKhqoAzEO/6
HWjXfybU1avk1N3j410YyD2vqWUVWAvwSun99FyphpLImyNaHvrizZstRrhm8+d4hAMB1e04/Rfe
CsXTXd0WxM4vxy0c8hB4MXXQ0NfjL2GJ73ZHVlKerx/TP7rPXBJu2Mjmp4UltPqaJaTksyYXtbco
RrrS2tXdJHynKbPMaxZQwG5bXTX88aWfOAzJ9kvoy5uYb9YyIDRCkP6PrfRCVSdqAKaPcDSD8kUw
qE1XSp0S7OZVMKr0rf4GFKqKP85U7IXaFp2t6YS7v97u3GhM1Xk6Z46nz2RRmEEt5xZYh5g4Bbzd
jy9Ba03/Mq8USLjFtm79t2l9Zwgy5rIMonZ0fMUmYIfZ93kiwQmeq5nBMnNHHjuJor3lCzPZoJEX
vTVUcfQ/fjAV1GKVQTiYqZJq9YX2daNXCsTxMbmfvv8dG5zStte9Ml9R/1+5TvTRJA0BK40qLkR0
KfFLDWxVcd/bpr/wT1F5Ytajf/L0bsDfRNGDf5GHaV49Bx5XAPCylrR4xnqyniSipsWny/QguT+3
r+40iGorC7uzj/54EP7spco3NxAg9aW5CdNyq1i2RAOx7cvmva4DPutQ34DLYluV/hmtbyrKciAT
+y5b0gYhY55e66oJsa7omAw7n46HOm9CEF13DWPeZvrmhsJ+ixKiKHXFnYXa63kEHoLcGyU+G6Ma
d+lgQq6JoAHG9/sojuMQX7UEAz5AoxJlmQwcOp65OB6x7djBv6JHF4kq7zI2GrkgntOxXwGh8jND
98bao4PMD+H2uilWwCIk0jWJdKq0+tpzQKp5mExXd3MhaEAhTakLlU4q8sFLzdA4YtDFsRZ1IQ0Y
9N1FdQFf13nHpYar37ErGD5eT6+3qZpSsgkDvLkERI6ePdET0cFK+xYWdfp3u2+IQHnMgMs8EMaF
BVlLhNRpKZmzj+T4bNF9G1t5+3gw0wVOvqSLO7qUjH2icpm9KvSq7yXmEmVSj+JWQVQOKbZeupIf
MmEqAqik08X6r2T+5a+wFZM8XFGOmWeg1nQkr3Pl7rU9DP6+ku774zRiB+oCBWoJfJgbYlLZfOkz
ppWQJQz3wzlouNLnLHPopHefobg3t59GWkoyokDeDxCaYr2/hOGoZYSCmSfuxP1MNMQcBPOILZwq
kDoe0hov4yrDezI1s2ldmUxfo3FcksrfRlc9hiFzyd3Bt1q2Xmw6lOWDW545PsaP/+RoU+bGI/uk
VHsJ8WcNQGyb+mjxiqrIzLpZ9rhrywdYx7PaUvmFMzPys8ltvnHeouuY7L3Webn4C0OdTX3PBiqP
eTQQuLQ5aB0jMCCPDuS1243CPysrmpVtVgUcCcJ8Kj03jZnRsSUkQjCTPrfYY5wxrDD2Bf7k1YoG
acHqK+G0eBrbw3TxzngVzrbEmt0M/Atnj7FcY0ymWasYg9sdIWluOU9yT8RyK5Lpbie+C9rgeGID
5vcKwFlpOhMJ4uuTPMtH2323bw9+jA/pzGgqHQjC0srR1rp62xMfx1FU3pp0dNZQGaqrpO1J/Q42
gyA0Bb2GSTZ2AskeKp0duto0XwXjzJTXcUpPDr+Oak+KB1B32sz4aNtNycmgb8S4Z0pSI+nJ9IxZ
0zRexjF8Kdw58m/uUPwS9QAiVLxupJwMxwMifjfvZkg5zsmJ+2JIlwHEhTfCe9vmbCbgJbpGFgSw
+5j3mBsc+nDte8xb3Yo7wDrEEwoCzyNWJ5do9F17jp2uanHi8pFmezJl+xDWOT41RG5hJzuVEApk
7qLkmq30GPFX78XYTrSewoHW14UsYxk/hTsczhk4nCCtGycVTdtLLCV28/FrMdbc+we36l4KRSbG
dK01QCpup9WIf1GEr1n2fUo7Qd5RuXOkfJuQ3Ky44pR3wOvU14mhfJQk4m+TzcQalznqv087+by0
D41nWZA+uYvEZJwy6t+eY4sqFoPbyN+NAE+ERJiIignGnq8TAoucq7TFZ5PZ1f0XWNfMABOY0dx4
P6w4EKpTZe1eRyVlm9qcheo6u/wpjeiwR65t8tWDNj7RCF6xMdfcvRyrB5fQ/HeIGejI4sbPn9e/
nNw6AgrzMR7g+xuUsCd89dQctZOscq+VBJ28rP+6l5QeijWwU0aevfcgGrU3onIYWdBEzcS9+oBG
STnhIl2mDpJIUVnL9DdETNDzsKPVZE46iugJ5uoLRoOAsWCN56/MsZdnL51eCvTZgTkg9JhVGzv0
WP6zE2CaYD/CGdbhKdRRpRKP18hRc4/dRZ+UmztKWCTRthHxTZ1w52Gt9mKETNSCmWPYlFC80d4V
kvcCtQqZVQlsC1Xdmd2GMd2l0C5zMy9zbi909VrWKCK98aBhkEFuXtREk7LeWkszH/LwbVJIWIS5
eZrEtWNml3KEAntcltA2Szzb90Z5SQGI7ZiiDOrpPsuqoAWsGO0suV+R/wyOMii6NPgyWt6rMpQd
AnE+mpl/e14Um69qPraBjMyaeu2p/nwKgxf3SM1pbphhrmyAAo5ys7wlTSV3bXNdadQhW4IsUavO
lBN6HnK6EP8nKlZNxsOykXC7pVDB6hlUzXc2Bm2NtMmNvsJksZOnQLLfxnwb5RQHUflBTxQFFSVJ
Gf4FHwBRPKEr2F95RjVHg3wvDD/kmPmp8uvSDJZBOlswtltIio/CnYtW3n8b+fGlS9paPaYgjKTV
NOTIenp1UtsBlZzD9SNvqViQYV7i3EFJ14Qb2dUdiWsjdye3+gfqOMw4e8Dg4jev78NQCM007Rl9
BA2jU6CM1weUxhKReT28vRDl/223rIjH+CV+2GzFwKKUQuWMvAiTVqL1+lDwTUnX3uJKE8HeNxW5
zSNWfJljE8vSAwTmzsqJlQ+qBoaohk4XWmNLvze3jm1vXBO8U+TlYS1nWwyuJqQlR3QG652seTRY
iGt3wfj2iy0fZurNJvVg/9AlzPm9c9yZljiUHA5BjZWvZVdJ2Iqr/bjKj7wZQPOT6YUqhtyKSv5U
jPQtiaAD1KvYUwIr7q9sHLqwXAXNS3GbDZ+elp6O94DSJAEEaQvfMH9Lsbl2PGH43DB3Qlwy5Dig
aVSJlsIWsxMO0WRDBOPDFl91Bp99tM8DPjvrqrZd5fPf42iNTsL+t//awcM9mwDLNUxrfM/UnkJQ
PDPNEbvEw0vs0emkiDrhHBe/FlPlCX7GcTpwh/qvGuiuDJmQj88yL64w7vlhYb08diOgJdIVKnWv
1rXiPtF+KaQs0zdB4wn1+CNGeTEeE+hS1obXK3PqFMkzlEw3zFyyCvzJb7XazUrLzAaQozhvP3aH
C0Vl/YE62nTz/PQ8D0ujvinIYXuIYDNR09NPwuAHm/+NVeFrY1cZl+wmsNdMBAfyGTQFyx9jVpHj
NcNDWx4DwBpJ4yfnoqS3tARbflJkPSUNsjuKHjXkcV2BWVgsZm+Qq4u3pHZyTx3pL12pLP4QMuq2
lqEbNFWzXTMr8MWlagQYAYjNjqCyCjKUVvxgwXlZrdWlHbIkjWfkD3DAQix3atSjsbPALvA2a7hn
QbCDpPy8qJ0w1SDfk6Kgs52R+xhV1MNQSF/6pwRPhdkkVsEQI6VJbU/NrE6BmD7M1BXwVQA5cemI
W2Jda4C4hzUMea3dDkRTx5CfrnNoJgpU211so0twyDdBysiQIKka9BirpTSyAUA9rSrSh/Mm/ntk
1+yy39b/7xIqQk4Bx3KIf686yd5l5zglx1zFzHr6tCp5tnfbc2RsogIJ7qlUf1OkoNlY0GXF+NBR
sI0Da+WYHuiSauzP6jTA2x1q+z1W+Lz6CSUdlyQFiktMjeg7nFk9dDE5gxchFj3+pukb2eVTIub8
1HFyuoXAvjPOkJAfQN703r0rnSGSHIcoHyoQEDWkn4hcOXiD0LUp4eF280OIMcDAhD0eA7WjtURY
sPw5f5+e8vwDIZXJsHoAiMYDe1ZQbOlEbtCARWAl4g5CL3Djd6uXnzOyEr54oevL14fz3yOVv6rH
B9Tlb/ad1D/hdZy7gaMu4i2bhDNSMBRE2J061t1Yuv0hUG88Ka2cTBhXafzVLmFjYtMR41llsdEh
YUleBH6yt7MgwTZStVPOSaloCiFZZKg+OIMqrdNDTVsP1clXrZ8WGrun2Fgrm9gddgwOGAok3D5b
m3xbDOO1AqX4L5AVC1uCfWmYDb56hlPSic+II+cftPc/9qeqj8TMxDjXoeaW3+IOvC1dFvCSeGgN
QdsOAKurvNyLu6AHvWoF9/BgK7gGMbMcz0PTNWhg9W9oRFf6KPlO9oYS+c4sGzvwMuiwP2+Tlh+F
9aCSneBVNGuZo7mNFZ/WB93SuMyATUWACM79aOg3eodvalf5Oivv0tnfvdb99xI9Ik499WbVBIqs
EVBjcvqQAMC3qXPFftZ+WXkGX42SQie4yqg72ymSd4hza9+cZl+3pVQ01P09tp08eQ+jj4SNq1i2
VjDZPJT/n10NXkqySMlE1gKGqxg51OKbmhAJvwRCRP+9a/rc+fsEtl5YKPe81XSU+yJkhOHxx2hq
dFKT93XGCY/Z+S7vR62QEcIug7Y9l0ftYvgcyBM8/sVE0qtom5wZvAmCppODhB+BsYbckVdizjT4
hbufmE6I798ci6AI0wMX77VaAewmgVXUpkkbfWab4ijBJSidLsJvOVIi8pXBRWpIHbwPm8UPqD8P
lGCQ0lVFLgrr2/Ew0ouIZJADV7OmawKiU061sPZyDpm7/eRPTqVlgAbyRPUnIh3VdKUYTV42QH8S
9sZ+oCZFve7MmDhZXKlZqKGjTZucWaL9HCWIjuNBicKMK7d+WC8cSK80dEh2x3/zxTdUPXrVTmIy
+2NCGrnY8BzNQcJlF5KgWv8Wp1iv4s8KSqlzT1ZBC4vicbJfVNjn8+bL1qpxm+Mp7XinVmFx7mr7
HocsAB+hwhg8fuJSSudcIQh7BAXDPucRrAjzL6uD4Dl8I+QOHzZfhQDMngDDijg/oPuxPljEPb+F
hn2FdEU6rEq08FMkNJNvXIjfc+9LAQ/i00Dnvew/GrBbCvilhPz9/uLB9dD8czQrB4nwKUmMEgnI
ndxxmPbFE6Gc4vPb4iAR3fdoKgrBCD02HmmYXoTOBxDSwCfq0W7Y8irxJqwVF8YYeZbxLUfx2zku
WjP7KcEQ7zk/h0UTS63er8L0un/OGPw+Y7UimcgKqhBZEvio+LKZhyNw7VRnPAwcSU8J1k6aIOfD
5JdauKxPUbq1wgrVPU86IlN5NTMgE1CWzShsFtoREmJeOrOURtW1V+Wfs+Ho3FuTHFYK6a0PJ/sK
oac6PiDB+8k0jnF5nNw5ZgSuri4m0tm9hjPGCHSeQgrJ3mIAzsLOWmPT8inyPPf1IRN1YVw/qHnI
PuUVKOL5ltAKPVWIPzHEFe5z5kfw+XyX0ySPSmrQgI8QW7evqmsw/QsfhD3cHbAu5RSQNX6l/CkM
xnn3/RXa5j0xgfSZilDMFZJWmnQYV2X4xP3ekNoLiiQ7XOCWn/o+VV4GF0413JbfkWprr0ufFof0
a4+vQme84F/3QC793r3S4s+34az9c7yI6uVSaJ9BWwDuh1lN4b1iXb8J5v8ZOoKzhOZoK0R8g3Xn
77KMUCmU7rmvzDMBr001nM2jN0nAlnx1JEe6JqRsZCKXwT8G3JAE5vAoLE+mMCqeDtC1hG22QotX
IFfR83lKIi1mHhG/qVibgXbbp7R7W1fIV1XryLzRoKQBXpwmzDIR2652CdCdyryKGe+M95Mm33LJ
0TUEdPeFOOevWp03SGaIbR8YAck6pwPluFPYARx2ezsS2pS3yj8UQr4VGOjLdy1emr0A5+1Z0JdP
H8dKHKsdgPniH7uhAM6+xUUkQXS+jRlTZaQs7fDy1BwFVwH5uAdgxmnqd9NFOVha+Abb5o10e2Zs
P29GRVPkd3mhBxpBilwvGEgnPxm9zS1snxOjn7qm3Fdd6UkFsqhql17N7IRmmb8J+z5du6PLZbz5
Oy8sU5yeHONjWMbROD8TcsOqYnvSmYOtgHxeCPxA2aFEs607h1eYirKQF4mAlx/vsP3IgsUZycFy
L5wbaSahXXUVJ2qU2a6s/KEKFu1FVcLMizNO0xJJgxWghQBskqxqY/NcpCBFPPl5i9xHCvojx3sb
A9XQ6VSap09YbH0YCdhchpORggJbtzRx4ZLhcXRhrJr6Bx0fGsexk86PoRJWlYLp9wjgFLtYqBVW
O1yNOtobqlA/jWpTTJd8aZ5duAvOjPegRLXU3N+cizj/Nzj5g5bPmWwil53QLPE24HCqGPZRuk3C
h7lCOsF2h85rOaD2e5Ouj6JGmCx73RXW4QTs1HF1e8A63ZRj5rNFzhpNsJLW+DIw4HdTbZM07MwS
qHc7DrHbYdXErdYuEflsYOA/1hMRRCW80u1jDUIDRLRv35IrWXUhF8DIHCVfust2tDZBVaVaTngA
9kkcq8YJdPWNjcksmun1kYPb1tsK15qqQU4UveUCZD0qkfketKlaGP68RUFyoXvSdlLxd9cPCwIC
H52zf3oBUPceA66u1vU/9eRR7KD1tR5hCsvduXLRmnFUNKJWIxDSPhtgZ7/8EfrEIa+dRpV2yuZQ
Kd72NmMroHSRCYkiDvsTLupy7AViCeIKmvZQsp46XUCqW1WqVLy2L2fMq9R+u3EmXonv5z4LVG9n
75/lhiSqaS06Ug6pFyarCLWZVTlEqsGst+pZ99olVSJ+DPODeJpH/GzXd73MrjPQ1HA5koeZx2yk
lMkSI3HGDaScKNZH0ZxMWq/g9SXrLFBIQ9EL6Sbt7Wt5YRzwSd3xNy+tlJshJ39tEsP34eadmbOP
OfjuRFK9pAXA3Ac7GYF/hc+0JPW8kgZDg+LEhwclUEcONV9Tc5Ba22Oqf4Xo2ScF+mgSr9J3IrSf
w4udPhQ6e+7p/Yno+v+bCFnVYG6AntYA0m+Er8tIOWU0L9eDShUWFU5BiBA32aj76yoGYWFgQB+g
CKEuCaaVM/0IMnmJ+NrbNV3m6bbvTyJp92PW0bng/UVF5iirnK/nIzRwIl6bi8Nhxwev1wtnJxFP
vtNm1GUA8EkqPFbCEYH5BM3tTjKW/6b+Knyte4h3UNidC6pDOgwg7GR+1vWVALhIfPUIfl4/FyA9
yOvfDu6DDCYp8NKU0wIAjQuQRAg1qMxvQXRgi/sEjFCSVFc0d8tPx6zoMVD7ttVzM7QSZQW/DZJf
teekjxB/C4ybR/wcJWIDFUr0ChCk/eVJ8RDVv5XaqNhb+db85u0VL9jxIcMs2hosRypb0hH/MXRw
encqyGZDF/kHldEeY0PLC8WX6kJx18tibmcWkDfM4P/76UVsxYqtgb9ZznLiHS8rwXwwzjVygo1V
oLml1sk9pvtAIaSVjeCQToDettRlZxAoKdToGy5ME4NvllA9zZljcCAXdf0N7mAHC5QlbgsV1dC2
/ceqsYLmS78Y5tdmzr0zGCTXiie0cVLSVrfcXLJDZRQEz8O1MOpVQ93AtvyPAYbUJsuQC9UN72zb
LEAUSPl19h+hFXRytz3ExFEdKSq8TJB86HMnIXM0Ah9+PDplUYR7UAlZhYNZbbVyPZorOe2PNgs7
TFkbLZ6PR3kfjHo4VAoFYswk/xN/HsBdhuX78UZQ2fkCTz1m7KlI8qyFOOctRY60D8o+uw8ipwNA
+CoBdbmHFUdsy/IozLl9EqI9ZorUbrcA5KwYyPLphgL9aVrxhCe+opfFA38wpCFlN2vk7nrUAhpP
+YAc6EnTPXuJKi//+joIWXd+4pGvYo5CW6OYjFCkVrG19yytPkHqgtlMrHihYaqyTQD4/VjuEpnu
zsBlMCxfzE9XKYif+WPj6e3Han1TdkvH5JiDGs4RIy3HyuIw9nnKeopAVaQJxe9lFcZdaeunZktz
jByOkTJEqEUUu1fOU8Ye8sWeT7WoCvoCgQ+fHJN+uqvfWxiQYwH9YJpxCNp4l2UxZ/2SjAf1poD+
JpuEUZUZt2ODdcboPvy4+Vs1AYJ4XWzz7JbbT/WUVvYrFv1aKfI9A4y+poj6oYVOjeepAbNDuMmp
AjTKQMdP+8fQ9Uv1bCbS4o0i64ZYfi5VWFGQZ8Ewr3jYHtc/YK7rObbWvPo+MX8Z+OJn2tXoWaMY
RZfWCozmvRYt7sTtyPtvFwg9oKojeXPvgomCesf5qSqDnMiyJqyZJ1sO024oqQJDy6plvcnLStE4
ZkN1Q/LJRC1K8mydeBGHWSmt44tjPfsW3LOa6CUS01RP+24Fb7jheJsjJJTIr7pNWnhk7SOM+Njr
fi8/2Fhb+f+5jkOb4Iw0oaEVRwrh8zjCL/C2kBbToUgxO/QX+XsM6kRLXtekmLrxKURUy5kPpCOr
/tjYwBonLab291ro88h0h/Dp2derCsGcf5CE3nclRujQ8MJylwsZ2uRsiIHBZ0o2TOUs2yI/93ld
RTaFiSBHZu7yR/Ezc//JDuqCWnS/z4Yd6ETx4kU7NLo5PJjhrd67w++d3GDzR3msiAlGk9XLjXsk
EIz1ByCvgEpPKxzqwL4cL03Yihcr8Re8HA17b2OzojE4QGZMbpQcqqzSadEFSxX1Hed0UOedY9W7
Lbl5ePsGG0Vep80mFHo8o7gW1hIs20cQQTJSZyUoU6edncJGFt6xJVcREilq9twrYbikBZToR4f6
vJtXfHsxIFsGlVB2qCZh10DKzEAGv+ZgAmi7fOYkNwL0vUaIcxyR8o8B3LeVOpvQZxM6sqQItWGB
arVcm6IBAQeytQweb12HzDefCMPwUx1pEBARSmYZkNfUIuDJc2ApBtto2CVbFUwjq7ANX0c0rfoz
Q1UPDVzmYtZQlWrKox2oMLrAeG/I1btSYQY3TtEhaOeGOzhJxPzL25Ic0t8wjSmKPTCVgb1qafZa
I7xk4HdAVZECb3Cpnv4SwymBm0/mklS/VJL40yLzP+gEWC+Y6W2ZzV2a0zFIIiljkncirhxeChs5
9z8zPU/UBpW0BMt6aUt2J/hHfk2VAKGDEM0FnuMuvzcdlI39XKpuqJBbwKqce63zysOX5XsiZQvC
FTnGUCFEyi3dtXxn4/FklCrVNr8tBajfsmean+rQg7Im0rWzM15Y+SVXQlPgVBu+MINyb84nJqjc
9vbr2paAqozVEOHRAIJ4BFVWF8yEIVHBl64UKjkwyEBafWx8JIlkydfKjUOZTkxjR2euckNWJHTh
WIxD5Ngs1w4QJVFZjynrXua5gC7Lq4vSS4VQ7ZYQJve13dlRpNqVrnWi+HS0opyB4cWdQp2gUcNV
sq63A4choM6IQVNuZcHU9kMilo3AB6+Lj+46bDxWy1u2g/4s1zQC2wDKP0TJn5SrwZf3YIl8vjlh
pfJOCf3Hi5bfcW+sVzSQq4Z9mzH8L6va7lch26XMXWFWbNCGv8P0jDmbhjstkttKGnVvvI68vhIs
nH/m7nAqtc9siecwUABsY7s03GcnXopiL9if7DcjyCVGOR8uxHeJiURGtczogi+uNNeft3JBeLkd
yvGF5cftNFBtJB7HqntCXWHk8oisqxVCMuh8DYDXV0gN1FuP8l3omFedItPc9ipm6DfOEFnAkRgY
gX212k/ohLDjlHE1KYYGR57CXIm32uJjtzs10C4szMfIeDadPhq6gtuMA60MfyLovIwnObA1EULw
Ek3lqDMwfSVoP1Eh13OgRaQk5Y8os/4Z93dBFqj8xBHbky6qfswEMDiJTI+G1R1rXZcwAj8gd+Ix
HXVdFEQCx9zX3usx5F9zHWrKLq1ETWV+21Fyvr2uNB0GzOaRQpBaYEUk3sZ3SG5ogqpyMzSfG/IK
4Rf6ZTKGCR59goYrbOPexztwE9GKibAUR6/IhJ53yqryFPoe861xofGQs2Wqr32zIUI03aM/vFal
46VRDXc8divFrp339DMBZCov4efFTK7shXf/EgE+lcCtkwtHIVt7Bp7+/Jnbh1duBFeAOBpCxd9L
GnP/7K0e1GqviVveeyWZSRLWMKNHsikwjhSmt+Dy1jP8K+6r92oOSIVJrxNBZQe8XkY3xMjv7aPT
8ar+C41CeE39kQL0aOBlVq9rfLiR3erD8jmBRcTgCjCyqnbKFiX/j9ejZ2PV38A2BdpgqjgO8faq
05yE8CxPG3CTZe1U0pK2GYXTqjrl8icWdqLihOMz0iNJCDkq0xrVKLhJ5SZhz9Ss+b3nXhxozyB1
adKNwhoWs2ksJdow4EjxtMvI1WvFdKyfKR9Qq+R0lrrkjp8z1nZc+aEm8RaZdRTaxe1VAnvaavui
jquegPuHJytjYmDR/Mo/N0xnz5bNNOlFJc9Yaqe7RfIaTkS77wYtJ8yh7jOe1rQX/U1WGjQa3Ag6
ndv7eF5smDk4OQAQEnTFzsau1xVrBphS2w3B5YDH+N93DJOHkOmOgp2lIPTYT7G8NaB7LWDUTMwx
D+KYhOrNxDJFHLeRycMFhbpKlHy863DG2Z1OHxlZG4dvzAbW+7c/uYFy3DbEnMC7hB7DYMATr/Xk
hbJ2AiksEKgMxnSKjRjISbpmiRtT0/FuyjZuieeKfVWbQuds4gkwrVKna7iUaLWn3vWgkbG3hT/q
ytUFX/aO7M+9/zA4JwvgpUmRCi0HKU02jkqBt+zVxmvQfd5Zvog6wBIp9oaaHl8E4vypg8UoJcU7
cf2xhCzlVDLM6Yq19Mg3Ecq3UNB9gGo5vr6JbpvEduwxxQ7LuoxSG0CFJXMmI0eYElD6pH7OUEN+
/D5aaDiio3c5tvlRRNtkGTafmnXbRflZZQ90IkjwVyLTY6uXuC45YdjV9j1NBcvRh8fuNsC2yiTs
awR5XFucgXuDa1MN+As7d/yy+0ds58YjxttWooCQsqYLBLe/CJP51c1IqOFqB2EjnF6aMvewgOXn
qxamC9xmOwr8IdyoWLVmoZa+E3cpecJeivnBnVHgc7iuNdBzVxQUSCs5YeQgia02kOvvmYoZhPgB
TzVXC3TzNlmmDU5PV32h6MBYmNrhv8m0+Lo9TesjKhY4X8atjGhHc30R5Lw+XUwcVKxUa/z7Hknu
aNIei7uTDAfUWV2O17SGdv6Ipba2UMUNjEpI6rwWg4KNPAP3VqKIvZdmhZ9vZSCQQ0VgRhGaNv1G
npq44CKFvt6gKk8sw2Qf4bv7/ksY55duP3eI0ZzU1wTH3H0obKT7T9l2uNIaeUM7qeXClMdMV8Xb
ZWj4JlwqFqpsNmlv2jqW2oeE+HVgHg1npHL6WRMKk22PwvfhjiT20eDJEhMVPRnUKVUNG+pvMzry
V9ZJl2l03Z2wE0ffll5CZLbsPr6zn/Wlp2+7rdcqmf9XeAi9b+0RM8S5AipifEs0+AmU6GOaFAO7
ktPBTIUrM6cgt1FHQ27ZWN0cY7PZ67mWbYoBmwqULlex4WyccpzyroZiKWSXdVmX8DeG9evUxC0D
3DjdnZ48oD5Urtw39s6W25PQuLIbxZ6dIz9WOtMebRLFN53fDPdu0I37mAupGLlh4uutyGnaNjeS
TFKC+cl3IX9KhBgvBRwHd/pD6//6Yjc1DO7bgVKN6l1nHubVpH/2BAEJTUEQTheHvwiwE1pmjF3E
pl2hdlmBmrrHYm0hrzcoC32hKgCtpeu19ep1WfIXKz5E6Y3TabFtvSNF+Iqno9DWd6N0NNcC4UVF
Gzdd0Sut517WbIi4BMYsaapFp+8+aJO3EhO+aDxCnmNpUCJsmKxZlG0DUqfex0tTbfTfhY1IWce8
002QuoYGAbESjGAWmIRPWJNBHvSzfmb5quyJPJGMZeuYD3fx25qVvY0Yecai/wKbop5MRmF3CT8c
ke/TYMtkUGJjDaV4RhrJox3hCHOG8FhHQ195pcJHkXOTafYojluVgEngfWePD2u4p1vFmvqUTtm9
Crfo/nueMQsd05zhPyUFx2KeW6wSkRODhwgc+nV+otFecwQO7hridq/0WIdON44OV0Z+hZgISwvE
rCMgZcVJU4dT8dQ9NfSZKIcaIN7Dl/VUCbs3iQHPkO06y6cUxiQoPW+pxSrkECl6ROgCxG0fIPCL
bysN4FQ6zHNbVxhivQ7S4hE5IR4Niv/Tl08Ksrs/P3Id82jQR/s7RUeJQUiO+3WodXKeJPcsRBoF
+fjzKrjK8KBN5PHsLPzjtp/GdpG//y20jxm495tscdI2pipwBOScLvwqXQNqVt450p3MIfx5CtD0
6FDC3Sd9/crFp5dya/LPOyy9J5nZ13nnHp2/QiDx72OCYFQYI8grjWUU17baNr4iWCQdBEwJnGCw
BDvnZqwmnRxZyBdYR/nXaxpwlbriNh3hxHvlybpAZZfc0LxvKCEz5ZVYRLIGELz0ONw0gnxAZcQF
MWwzhL/Prnb/LpoQrrppZcpf6G0oLVAq4dhbEtsp0htQOf92vjn+RXsWcAPp2Hk6ZfIk1AXw+41b
zfSnKncgrgxweldgDDZvTM+0NX2m/T77+J3xbP+RyzQKJU5XerHMn3cEQCHsrSz7RVUl4nT8KiQn
K6LRSebPtN48m/iPTys7qUee8dwqA4I+xHMswrVQ4wJxhHqT+4fYMgfP4IUpUPDHTWG3vAZdexRl
0/eB3T7atbkiEIGCnBxcDJL/KvpgzNSPfq/5nssGpYP0F2Jx8tye905D+WEy9DdNu0Ix7Wz3qKLm
4GDn2k+EmUMJbrHUyKLoMoKU+ZtmIoSpNaL5QbdMZTbcAtpgDhQp9zzwAy6ktzMm4AkDY8sCNbs8
EycLx6K5dbZ3x1UUcpMJVTTXq7lieYTBY5zcv8SrCUoSRw6ny2tpmaeORCvSPRzkZbmKkC+Tl25X
HhFUGyT5SLr6KkigOpEG65MRdTYp/PGGOssLQwnwxnAEgonP9ej+Zw8GdZVORYC523E8urPKQ1Pz
LjXzsAF3/yMEqDkhffWdvtXAyPS4+Dh0HRSCIjPWWKNRY80idQ1NoLDLeGDfl/Ka3RGYKzgIQlLf
M2un66bkSNGk+aVad4UtU/xWixDSjuFQrMUSKzL+L7s4yVLdv8GWmow6m2KIGxrKJCYPW4bwKR3D
SqOmur5Wl4HuGdqLP7W5gs3lDQKo0uc+Vmfj85qs/nsCoErKA3jXqMniD71t3JC4qQUjRv3/Fk8W
4GfiD5Jx5Q1DH3UN9xWSXZt6TQ4A3q2q2B5M70vRy6TyLaIzLZoxYQcQAZN6oucydbFX8x6Wjxmu
NVdrGtRbEU/Ad3w9e4UXcwhMFeylKxlToLsU24/0YpGWzgFfSFlotqV9uekS+KRLZusO3myYSE4w
V+1hXNG8fHbhCN4iHHArm21WhA3SYx7GEh9pmhS1Q5JgSDvMTmPmX3a9irL2iDY18M4+xiCTJEPB
3ZnyNlp0KbMjYVuZ7bCGW6Ot3nDg2jDsZQ9Mu7+d1sGDENT4wLtAr13c6u5+MYeBnjYghKWMSbE9
2V8ERK2Ovpezz6mH9MQWVTT9tPRr3jn7se6fmDVF7WMKEne3zMsqJyMrfSfJU3LJo1nOCiUn5j5Q
cqAgj6az3NhKEZEty+lVxD0TZKGxSLHa7cJRLHJTQqp4d4ewWsgwtaoQPUCcuaQUSP5axoNc5UUV
AtE449+XZuw7q2dnpgBYIvY6xkSShnvqcPH3gKa8qJk/2oNHRJ5gzxZ/NxpRCmU6IrQjY8Z1IUCU
aFx2lTsK6M7ld3pv8y1OK9YxDSGWkgm/jS0GnNYZ7JtC2eDuhfKvBOp7xjC4WUYbKCFbHSPdP91v
tDuPUaZpneojStbbrrmjtIRWsPW3L9lBem8LHkpZ5p8wwVhcQzc9ow93W+NrlbjN8BKV6a7DH8Eo
7zChpj74n95d+LvpR/c1A3fyWDynt0+3aKKxCPn/JyIIh7vfYY1JBjhFr3IyF5HQ5GPdFecp9A8y
Y9680HfW3lRZu/hKAk4YXFuSRtgHiavLO8RP4FO+lWJ7R+CL13GzLRHRUQ4nCKkg7iWaoHz3OFRP
5IQZsRUewo1S5UegfxE+gjQwztjHcYJgoHEbf4ZRHnzUERW26Q5MZtoXXzA5K1xlUbsxPstbXlyH
RvC3RI8q09F5uF6powoNWRJ1MMdSl+kMRjBYuQNAyi4GCAv0T64yfgCCy0l9KaP65QXCao1LWAI5
sEpXdbXQaeeBTr+e0Mq6ACyoFcqqqIZosGQUR4NXJ+NjgwVtZX+8LCWrJiAmLTzh4SMGXxg6fgVO
oXU9+dWV2IRA2w2mFR3IfRVeUsmiDQHQRru9n25VCvpOtKHNcRXnflUQSI5lUJ1fdtKLDvy9+bNM
zW9CmxNWzYbKaWemY0gns3eD4ihEPyjogNJXlM2lRQsCJXTn+f/JUfKZRYzXn/bOBwXvetkVUAGs
mV4mGt/x3w3SBagtebmrIKNzV03d1GVHcd+3EsFZYGDsED0X4cyBGNXY4ApyuE8JvL8u4aGbGY+G
H8xEiuVjpzH2H4hI8RFNR+3571cvt3aUaQFmwD7+74y3W+O+XBy49Tqz7CdtAyrAb45px4aNLl4O
qFn8t5zObTu2DpNlkdT1x1W8I5t2sSyC1IdbokL11ES7JQbw0P7BVJrHYvRJnNkkU8NcnkxQDRKO
VIuetAGv62WtKWoCspRicedM64KnIW5KjCzNOkB4V9COvzGHU/pheG7sBDNDevzi/QVyFnvS8Dgv
hCOswSqFfyT2hJAS1o71j99err74kjUwxKE2T7k9e9aFiODkEZ/dqP7M2/Gbyp35Mi3meeURPKTQ
eotSzBOZQm0hw1mPesUfnNERCacYhmmQJVyCCIJYjJLUrfs1Vsw5pbskUHFNYPaG4OGrbPLiuDx9
UfEXHSIhPyxM/vkn0FthEVJYoLqGtGrlvzspkSsJKSEQ+L+6Ay+fuqmrvXT6zqbnTGmr0BeJpZcU
Dl+uBbb/Lhdw7J81fX+4stFUQzOhkj4XOrTMS+1vXc2vxFU1C3ho+UaUCtizl94nrj1x2Tpizcb4
lQif5BOQIJl0TTa+9ca+zj18G7uEAil4ZryFuYOvP1t1UEpTCFpVuMu8YYtbkfuzBw6wnF9v4etI
U7C6Gv/QXf4vdhycSdxnrB/2y7pr4Y7peDUQFDJwsjsohxEfg0n9I21cl7TeYM7jUmdjlxXSii7j
xbhCCPgHm0MD4pMAJJ05IxyEg5imJmiXdqP3USXPxlOLXFZGY3N5mn0SJzzTn551t6YoJ3IhfIif
MG39DvQMvVrMLYIzxha3JrIBBUqrOcSXCfEKBcWp0ylEinMdfsWJrgeb+fAkbbY/2b2UjvivzHDr
1Ej/P/+4ycy5BRr2SqI1dmEeLYsiAOW3NyMMb09XcyfutZamIkbCIeHKONZEo3arViE7ZPzoVsZH
qEBbW0FYrTpYExjR/wOzC2G9EMxnODpmg2esn6iS8f+ob86yFmusBRq8V5SB2R87Dt/3YC0TdW9w
Nn6/RkuB+DX3exdarergOsSnfmr5zM0wYiQtjLHeM7xfMpKedVSmDsbNIFMp0CG6I4hnqKkvO1Zy
eH+h7t0YZmzV/1MDCYTrrV7Bn842q16jaSBdQaZhUOcdqje2rHCbKXihTU89J84bTOts3n1P35Zn
a0Ow8KhmcIYcOTOpaK7nqHRZmE5RfGLQChe+ckCOrmB3Af3z1m7Fe2OOaUpaGjFIDAemRDTzq5w+
mHKej4seg1/ooMHhC8zrPx3Q3X9y8+x4fs0lVXFArYWUNXeqiGHlBDfK4rc/kjd2UJOMtp3aCcjT
AOYnkGA95jslodF1p4QMekJjaufAXDAhRj1i4MwOymF8aDN6ySOD0RgRuBqZI6UNx7R2Wiysum8y
GxSH+dYl0QAwXlFMP3TumALJ/mfKvyG80zLgz369XY4BAvsUbq2VKmPNtAYx36xhI3dSLBSaEuwn
Uz7y7Shlh94yDEkyYqJ89i53SJv5yZIynXQudReMe58RfbISeDo9R59TuMIhA7F51HN6z42cF9nt
Orp6GBjtgAdKYH47Aejshj1inY/JpirBxdoe4mAY0Zk+n2v0G91OAUvd6Zyz9qrG9n3nw4VA7b8C
m6elPiRcPZhydIXr2APjLf7gIczcRCtromYnAHTdWVwgI9w3GDnzWNSnoSNdVjpS0f3yogY0yDUG
sLJFsnvxRd1gcq+5u9PxvS5omh/cu7U8z0xuEwzki+BcuxiKPLyrG+tbL+f/piR+2AXXxXzjL2QW
mLDcgKjXeExJ5AS/YVnKPqi2L9F/cjmiF8b7JjPOXSxf6DIj6MihgILcHpviy/9f0vNQAKl+tkBC
/OM5d0NwGm9upcj8NKhOTx90G8VluUZcQxYH91a6pouh5HeZPkMFh6yNBjp6tYjNTtmSNUzFhMGJ
DjASyBAtmw8p4MCQzaZ+TNRKXzB21wn3KAZygTNBI0hTzuSjUYPR1PMsHBrbzR4xFf59BvftNEh2
htjzzbpkL/eGx5rs3hkrZM07ees0tVFMAUxBsAxhzyEzfpBDoyYoZVycZCt8U0Vay+t8GHLtlpkz
7bunze/w6VgIKcQZN0psDoANUNw0QTKGzdxdgTvxNg2dDxTbqScoKZUcuQ5esOTiyQDVHCZ4WH/E
ETBgIEDrNqfTU6zQJz1QyHF2Dtu5eT3XzE7TVF7Dsf9CYEKQFVmkY4FfGgOR++U+r5NwcWEBbpdQ
SfOxNG6/PnXh0gCYR4lN1McBmrihkIsiIH1VTPapGtunu+rrsPS+8ip31c+UNDminVdvnE9RwFZQ
uWBKN6slj0V/KTpCddeDCKqKp0Jyy2qRsoSqBqiFiKZcBz/36IbdMmHipwZb4ngyXdaanW9kbCAq
8jDy550Q9nCtZ76SgpbNooiSP03oahyl9KqZxyFzDkN8wCzZsvlG6J2TrNpZ14xEM836gijocngW
BbwioqA7KrQhrEbUkx9lPDyGj3aFa5RwXlZi5VCiuAEBRDp8889z6W4gsoC0q+mz22x7qYDYfW2E
/JrxLFMu6/kaqgDJiNIwIl149HjptwWkFSQHbdnmyqNfcfNuk3MYmLepVvHbB6aNV60Po6hFBlmc
wpwdIh0C9T61SW+yUIeI8wq5uthCtDJgA4AVyp659VGx8M9F5DgH27FwYn77x9QEmV6gUnBrXUob
GneH988k5P9T2aGqutGNY0KMpyZGI/6SnENhG4LDIzjFaYCLg89xvmnOoK1ljuBH7mmdwIj6EVuH
3xLBuHG4LAq0ZeymKd39NiVF6I8KiekabXzCum1mpEX9ICNqhk2iBAn3ip0B9ItFgm+AYruPL61+
dgTy3Y/ogqjM1Q5D1gIMo9crx92oRYP0xqKXTYP01cy0JOgT2g7BaK/JCNNl5aHoTi3JHEF7/z7Y
YZ23dx1RmBPZ+wjksCD1p9R7j7cOl7Y6Rp9A7QKWPiB3OASYB10Jq8jxdMXpeuKJBp67zKSXCjNp
i3DYiTj57XUPYaI0Y4zgwT0IU/JEm0J01FndXXOChE6diAiZRflo8N9G4W5lT44a0SW306nu0eiV
klfD+kfFtxykIEmcf15mVNs5h9qKb3Cet4BEKTjTliBXgBQfxVkFKiXHiRFbPZdUkeG9CX2R9JgK
knDnf93uNcpDAxg8v2Rv7PEol1//jtuXH22MWx+1J3Ff8tLRuE9A82aYaPM+gKpHL+CMX5RR/Feo
uzemGrVDs/ubja4Kd995mt6yLJfpZihrwFT3QtGkA8oSvvLoWBpjItDzEE6rmxVFXsXCKLAvi6ME
yDbncAKVjazAii/6glR1tPDkyCsMPeIAijUvqnyPgZ1lh/lEGOpe7JVkSQ1n6fI9+qjQQTD36R+q
Eqnjc8Yepbn3ct05xDFyEOXG3eGyQUtHeqrmRw2MbqC2avP6WM9fhmYFI/Qw9lWJMhXuIIRM31Wk
QyPc2u0UQTbhgF3gXQLEjLtpQGxg75Y8rvdWSz/oH9oy3oqeeFw3Oo0zgsHLOsdPihJvzoPZYZM0
ulQuQ4rwlP4nRaXQUsamTWHzTFqgCLt0mcRRj/afSycAlDFsG5lmiL9a8/xIvhYzSqn11OA5wbsG
58CnWwviIDh6/qpsz8/pgniKY5jGgYZe2jOLk82Oh2tzvSXyN+G6gnn4ARgTyMNeeB4tL6T6opUb
OP4DZJCgCNKOy3q4VqnsBhe4i3ese7iguNgYdn5hWBP0owrjgbKKSYs+zlI0lOTlxN7t8nT7yAhi
+aGnLjAx4kxXs0y1zbryqtaIBaA4vAwB0CcMtTc1I1f0jhdIsWbH3i0tGV+VSXsPdOrJEdSm5tLd
B4UH4T0+kAsqaSiOE3eYuXZ4iaMPXoPxdD+PLlNIF5BZHa2YlmN+DZJ4CS8Daml8aRKH+E9v7TLv
hYxDvMgA/Fh195Pd6bBzNKV4owUGCxZwwXn9oF5enc0DKEJRjmUhZMBFYRKWPdRsE1qM7GKqsBeV
N72djzn5jLbiANDa7bdGZyryWeIrn+/QmRhnVKj9XivfuTU86cUwvqjvJX9Mq0gTrHEriJSV5CnW
CVAL95KUQNgcjZmSIOqSwhi0AKyYrLCFzItVtOU5AptVNVyXJpXQU0cwBs2KqcHsjcn4G0kgTgzZ
MSIXbxYKTinIJyCU//4Nud3aHUJFWFhNI72Lne+jka4WAl/vJeWRrP3naL8gf4Vwgyvm9yatm+Kv
3lAIsn+iOVFL7gT9abKxKiuCEk5dOEw/hIi7u64zAB4YsUtTFaGvF+yIbjfyLxUmVYzX8tOIe4Pr
ZJ09ewPsf/Xt2fQamtIusAdNQE9sUJGnm/Ox3LrKQiZ7bhSwGRXiE9Ro+AFLRahJBMjq1/zbCdP3
XYtKYD/zSm7OU/itzm9+8Tv5GW1RyGBke6cj9RkcTUpx5By/02PAoZLGyDWpuRNk0TOoH8tLR88c
Ln+aDz8T+ULvhzdBuF1ZCWmHqzZR/rngC1v4hvl+mAToHQ9/lvr0rsttZrq1VKmoig3uZUgL753n
czSyW1lxuDazBsyma/1RamR/uBpnF3CSktt681pjz+HueEJonxm17748+dDQOC1Po4x8pPYAYvt5
KY0I4eUb7lqzJQBrh14rM82oT+hcwOnpoa17G/eQJxWrOLEw2KtgvXmuMpxeDUgNXPe4N4fr3QmO
eabD4ZQLQTfminRzPPevRM6sxsAE0sdcPGxlnaF1WSf2CyaXkQ8DDuo1cPyhNEgvmBhotFn1UvGF
AV23hcYrICi3fS5djICHbEOWtHjGj6utFZ56WVAHB94l0jz3ZLh+ZzgBX9+fPjr/mpbZUUQntL5t
6yVPZwk/CLQgi6UEqso7VlSDml7vEM96/6m8pBxel6bFPI5KNmOQNNH7rUuSWxZgFc13/kIBnzw/
QexTdXZ1Ep/w8jkf4UspnQ2Axqs20CWN7sq+ncLEjKLRm1mJIhkd7f0wNXkQJARMvh69pkJMrjHJ
06yWO5HwCp1M9PZbdwkwnkJlco/XDQikGB1S2a0I9aoK4n30sjiuDMJO7rKx9O4oUb6ZJ9FAqeCV
8xF4Z2f1q13kxTrk8pJu+5D2dof3kXDsfFUnqhCf1Qtny4v4TvQuwWPRvRCBJByBOE0JsOJPvF/C
chaR2yX63afKZF48F4K15LaJ788DwQAOhh2jtTo/DtxFXCFhW5ByNCAJHAiGXsooQo/eRFfq7kwd
q6AWXuQYwNpR5pg68RbUrzI4gU6OpXk0KujbyYBMA0ivLjdigDYScz11sk1h4EFVySF/kROy6Jdi
j6YB2jiHvIUGQ+PBbgs54M1wQZI39d1f9P8ozARmsaV/jVllvtNNC/fVJSsHZ5IGSg9XRRrXt3KD
pOOdSmpwZiU6nN3zH4iBYcAu0Dg9uXg/2YWGzOOF1oU+4DFJZaKc+/X2+iUzsGkn+t6sj0kQliqk
KQG1NH8m4n7EKnVC89DXf8ygdF6J9jREY3lZC0MWh7IdErCkJp7F2NFhkMc6Fu55FsUgrifRYEsc
W3tz5wHt4AQznmKsy4pPdNzRrbUckqKBWqgV3+0/N1YV6CQmHhT+iMy6Hotxdx6BgBs+KlWB5+xN
ds4CrEj9qaUMBgGXsuEqgO8tYm4xh2QeOpizzzv8lu/Ey/pgqOj9d06g5DDa3fZp2bx9kDxJZnnt
mbV8PNRX27s+XZmGih4WQXDYOgQpwXjHYmm5hyVmfo8L+QcifEXLZ05Z9V0It82T10WUkiXixBQg
bVoj7qBSnB7SHw8uVn5L6AhE40LwrXyHHhD5G2lCmlK6XrjglcainPM7jyxX5RIe2UfEHYmLLKmB
lnTepjCeFh0rwDYctBM7cwy7gzOBR9QZCTaT6HHJFl3GCAs2iRhsYpc0nVR+0s71ynG70f/kD5MV
F78SBeytmuml5GKRKViUCRyF/SOb2x3TGt3U+9yHMQ0Te5PbkqhgxVP8mzvwLURdsL7+jLsPvw2q
lW4xTEn5nuHJfDdJdvOvlL4/LGsl8jdZ6E58AdyeafGr5FTjEf9jZ/nUFE7Iar8pIpBVWWo2+pwH
T+SWdedYGGPhFNO5yK6/12dJlWoCn3ORNltpHo5U7BoeLcgtIZ2mbvE72KXn5sd9M9SxpxB69L+g
e30/yG/ngIx4Q4y7HWv/thgemVX+7YjLoUnHQFarYKgCKlI13a1XcNdSfry2EM3V6ZyRs0GjynPK
IVfw+o4hGkss8l6Lbas/CSrYYLsJdNm5pF8vaJ4whOofxHnF4Q5z7sXbJ8sbUBMg2ZQPOGotbjj+
5a7BvF0YwMgSV8QX02ft8ETnOaJNRzKZFjEPRqcs9A5Lj/5ZLg+3PufvhxpE7AB158pWt+slssG1
ENuf7J8CQdwekdUbtkzoRCcGosbx7ssVjUbdSADYRle3xang3TqoobtLib9xLptrv0WqNDa9TtAh
t3nm9RIz9+WesiCgjHzdFAufCrJo/UCMIYZaD3dcTzdt7sEqIsbop5lVXMZwNLVv8PoX0vytN2JD
O5hPAGpEQSe6kBef8H+oC5s7PAZHggdVbO4Lhad3sFsOmOeATlN1NCPB8x6mPU6K35W3D+qZWAlz
10SbL/dk15VA8d0R+jvHAHSN/ZxByUFfZy1rIvNR5lL9C0xRNWkS9WlBncbEZB03UOGUP/up0dLz
C4r+wc43YQV2kTwHJq37eAgJy2YSEYfBDNXf+5xTGGL26qU9vd+31z5hBg0BNvtHNb8fhaMEwjTs
cMWwMbwD4b8YKzwq3E7Z8+aNrEHMlm9ia+VZa2mHpKh1aXHAnAQnTOkwvTvIot91Vb59WZzs8ymu
PwTzvjuxHbxYMj/sKuQtjaX31X47JWJiqUhUFAt55YADlqkoIdr1NMdWTXQBrPsXKOGY0MLMz4mg
+KfFAMRfUo6xowQqzDAo4qiWt5vKXP6FGM7Vt0ugLdu1c4S71c32+9nclTl7y8vqqcmDNTOCbRvM
5+V5qXj3qRoQmThZDFlYBJqomVM8DT8roFZH+7BW516cWDKrYNe6wTtOQoKuEHCSQgbowZ6CYp4R
QMI0MMxQKA6w3tAcf1tJ0Ou0NUHfCKGggXRwjx3iH0SLB87EP0ZbEoqnRnshZr57+bNa3g3RIwLC
Rpg/cGQ1OcMVc86nMxCZz/eDiH0alWaOiFxcjI8/7IJSUe3/L/kMtKFMtmq6rfqdUrK3dOZ34aSQ
vbmg99wKrdJ/BWs0va4wvL6j2VNGu445FIVXR6O3jq9tLY+v9D/h3Q4SUGP+WqnOwmTglADU3opo
ev2v1gxLaKq7HMGijc/VwWwU+0GEiXqgZ4PTUzuM7lZDqEwsgOt+d3nqHR4oEBAFG2AYMkYS3Xw2
7TSat1e4uD/mi1bvHN3BpD4uRZDnnLQapc9KtUo/bxGleMlwEm3z/1r9O1b0yZdeJacQPerFJBn8
aGpC5AnCK/TCblsIov7xWxmdtuOaJTifVh0+yEx17agw3IWcZFKl+lLnn/tJLdBI6KZ6k9tGChaM
6UtCaxwpMdqVZsPMWq+5fdnfKQPvf1I06VYcEWAvDHV1nvYIQXUViAX40WZwjAVIR8bYRYJoCwEI
gn/Uf8ceRNoQPyk4HncU5KaPV4s6ldNKHpYWAh5w6nwuhBPhMTs+46E2f6I3g7+6FXNovCOdyekx
YLRpikslITdPQL7Euon5kzS3a2D+mqdpkOWfTkGBs41sF+m4jeux4AYyEeOj00QwuIq88I/LOf1g
8oywvzyBnXOj+pFAxAuqK7wO+H13E6OcMwkp8K1FaIXzqSzjYI563MFnFro8Z/4Jlm31KSGCIl4v
Keekd6/+LO8hzG9UdbDOmxegyFzbN8aa70HluzSQ8H+W7hE0Be/jgx1mKaVH0IlP57Xe8uyvXVn3
dN3p/5elohN0JK51lJuRfTgWDJ50dYY8WDcje/tveJYOt6zhRJnNGASOt6XjobYADkfKHg+ZE63p
htJc7+qxK+kZpAr9yIfgbDBqnP+qkBfSjqU0NbZn957c0Ekyrev3cdH967//qSEltlLwuKomfvZ3
D3azTsV7bCDM1fXValUpsI8wg0Xer7uIhumlJQFPvaUsLaDrjbnkZVw14io7cBNty+eQ6mz1Bd5z
gum263nu6vSBl4L/ELohFoFgJdzrh5KPPREMCv4hBLBsU2EFs50ISik4Zb068i6ZFp+XQFLZ2YH2
iA3n+ZXW+zXyr++JYV8h5/+6IvHd1xZY9xmnN4sOEFACqURrHklB1L5C6QexC4ch8Ly9NNnlQYLq
mvjf6WmrLIntYuPqf6nAngS4w6pCUHQUu7/dDfnb21GGaBSnDp1OV0keMBxvmGPJHfDBVkC7174P
fMmwElRCNobeIa/0nhXDHCzEQKX9yJOKUYDnF5xcahZnAzuBEyXB8G9LKHPzfOHMZAEMN27zuEFQ
8TfRbDuUdY94k91CCOPKFsnz0LP91qeI8Ie+nyU3/DhLJITeGQxjpcVWSwgj5eorE6HmrFfKU5WN
jIID/sn+VFwbh59DVgApxbs18gYEb2ZWjaGq9q91QPYZ15f3iKWHGpjXdJaz0Wuco8LXw90M0+kE
Z7q6eb6VvBZRMPEdxKpqY6pgwsrwN+rKAqlhhT4/fYV/aG3Okng0hyWZ1EoHtuOpI6Zzb0hiuc8r
SKNML+4aUQcDEQ92V59yS4+VLGF+ZBJDw7teYmH7ccX6xVrWLlR7JXbztjoNEtfmz7rHQe5GhtwI
fd32ZXthcDVugV0tGjrzb+qSCmyrpOVAb3T9aHlVxdFJGftxvy30fkhzLRhVf3eYFFIp6QHxe5V1
myIihkpPQ6pi1SKg7eg6y+NyP4YCHDaRTm4F1JzRY0efDdrcOja5rOaUOUCP8IRyYgKBjtJn5fMd
5ZjO4kz6jzkllRcpL8KPVWN89uagCUugmj2ITnYtX3tWqlgWE9CX/fpSOY8DJa/k8IFAvJbh+BGB
Uac7vwsvmpykUOhGuE7SMsOf8Wfzz+M8myukYAlY1fb6R0bR/Q3z4/02A0pxNlU/3lARht+eP40F
ZR6BHeMacC4/hsYF8nsvxV90fplkgl0Q6tga0hiy7dwkgxbPV0bdQpoiRfVektEYziJdPYrpuPLJ
PJMTEoA707/PBRQbga9nNmJuwatvpxUfxysmqHVwMQysc0CN3CTKyXTsaiSeRaWkozO10uoy6Igu
lBsNLW+F6YXhvL6cbV94jMKyx04s3pe8HKYyF0RmDV7ESvIThptNNPvVYaTJ6HqE1Y9UxJMDmYt1
WbiFSJ7nlgNWdUNarPB0gYpvTREZXylepTYta566KwYzjn3wJp4RJhZMQXgueXsM7jIAo36ZpTgt
OkMfmkZ+fM/DWD0zgskgNaO+3VvwtpfndrOpKXoZoFfxLJrr8DaijKrPRy3UXfsRpIUvK7oRmILv
jzOCkZKJAkTb5DRy09qXHSrHw57kOHKZRAuXhyIIS98kNJQangldWLe/jskXKoOzZMX6/r/74Pn5
wsFbsZorO2qV45YPG0IxBh9yTh5cL1VhS6fbSDkPZdlQl7yUtq/GG2PdxsraAS8+OBv92pWBooqD
L3jem5Tbd0n6oi7wcfBWr4SA2X16u0VY8EekR4D56LXXENPVk6+Pzyrlv6462fHSzW92ue3o2qeT
QtdEq0EOV2DR2vEB8+w8rzC6aFPEVhzMALi0QLD1oMU2I95NE4A4y4mbcPNB4nYTz+M0T5tRmlRY
2OFDv99ADHnuZzYp9wmnuNaBUiLIP2QYuMNdpZU6D6hBQ75bhOltKcxY1nO9eNeX/cM5VvhoEYV/
t/G3k2FZJzH91aXc6t6swb8mmQMyVD9tMkRYwAlr++npqcE1PZdPUo89SoWPrgznkyDRxuKIvhzL
AD28l04Jr1isR12hFh7zVJRlI4XrjXQl5IzCfXItGk8DLlJcz3xAKNmO8IWb76+8K0iOZV11ZRtF
L+U+jiF6GDjl5jcwTbE9nhV1K2+okHEeOSWwIM3FYRwPu6WxkDW3KmS7JyBtEzWZeGVOPCAlNhfs
UL0mg2AdHly28f/I30K/KwvX9XDnJVyeUIYHyou0y/58ZQnb9SWivPx2kkqmvFZhp1kU4SyEwLmz
lga+7+SpLlOqfZ6t6PPY+0TA4N+IoJwq93iU5JLZ2ouXLsXo7hJm1lfnk7XyDL+RUPZNzPxDZ674
B+biTStzNWX9nkutwWNfnxWrZhwXmwLLT3skqErPFeqxsCgNE9w5dOCSOwvfZWCH4VjIZUR9Rs/b
VYoxB+8r00F3/dwrZYlgfX/nzGksanWtHHFO4rfcxzud0fqEeAXwXcB55EEs2X/XK6erfr4Y7GhG
i6RitMGoysDhmoPvuiRAd5KbSR8TEU8cDvSqooQlF9EeC5JJmw8uRiGU9v+51TTszrGc1uIEcqm6
xIJa7Jo2JWWXdIxhKxsuR4RmLl4rNVq4QjiKe34se0iVsiKwtPKSK4U1IRbaCYpBoSap5qK20cUN
SRqt0XamGvpEJPEFWOIjQjwlkSiyURsokflt1Pfr/36HnViyfzz7eQV0ckr49NNSzMs+JaOMWopc
DjrUuxYfqXhllalVrPcRs5HgVazCu2haN6VbUuXTH1GIOG8OPBctF7JD7wfdWwP+8hButPsab0mk
Nc3KdKnFriZRhIIpe/4wKlDn/52iyr7RRX3r9aKQLNGd2RfLLSq981bD0OYeNlQBxfF1FIdGPc7K
WjZw5uiVuQ6eLMfPvrihaT5WHLawIURyp5OkPpAO77/isF7ruTOGlJym3Dawy4mJ+AUwRxfh8KoO
vTrpyXdkyaJ4GLC1KoN/KYXIu6czGKJN4tCNdmpNLl0SU51P6hLMgSYgugSd8J7/ZR1lQ0gg76mk
DdGX3HRBzz93eAbUW2R2gC4ivJfgNqC+0XUExOsf/uNCdEnXvT3qJNXRxBuUSypu/+Vbkt09hEjL
P1fR76gEYblEu9f4Ts2c2l9o6ttsdjHSy+5ZKdpO4q4FASjJrjqAcC/uc90FmXVDA8qGSEdHxy0N
AYNWoCx4i8Zt60PeKvFNLu+WnA+OON6qrfRNYuwuk7eL10sC5rTS8vjU2XmFXHTOWvzyo8kNANwx
tZC6fzaaigHlsrZyvB+3dK0QKNnuH1BWg9/JGuKGm/FPmsTfbgpf5TfBFCxucam3Lv5t9ek4+4gd
1QwGGcp5DEbG4jlxO6i4vhR8H1eSPbXmkEn8hkkPwXA8eNHaAaEjXIjTL77bW/r8HtBs3WG2mnJY
la9XZMDaRlNVQWs47IVnBg6vjTcnuOVBvnFnfDinc2hKXis0e8cn7T/fbzrEIG3N34IcKjBbCpfX
GKElnDsXQDDBMGuKwIeQge0qV6wo6uyhEip1fGcxEQADoCHjOjSJIYyLQowg6A8gh8cxMwWnhh0O
x02oYfG6ejkwnl9Jem5W0JqnO2NXNlc6DdYUJCLUGNUj99vkiVwGUAGHg/6Wp1rcRin3uXjHNUZj
MkO7Dk4rHJ0KV/LXnDz1JszF7QPmaZxoesnp3Khl0r62NhLjOUXIpB2+F0WU3fjCN1F/FXaIImV5
MQs7tm0+N6+TLQFWynbfb4UjAUpO1dsa9kNCZUxmd71tjMg3wtz9yo+Q3HDaKmc0WHqi00EcwzdN
tABbq2MtmVasdAz5I+VDzqcZOwZMLFTOXGRhbUdueKfUc9QLW4gjwr9T4J8fQmPmX1YAFoxdx0OR
dVirfnDeN9ozsudq5d4/ZdxMyYj/DV8E6a8KVQoGH9grnhvLqQTKSQ/y+8PhHCcq/Hn1sjIs6BM2
1AFiZN+e34NOsVKJhc7olgIcAJbRUFdhisEcBVTAJjzdVuQvMAUcVbFWA9UtE3eBFKaDsHJLAOgh
jDnU9NpfmL7CpiG1wbTDa9X81TvvvmVPxEGGI2bi5aGxaZJuzM6YOHiPQaXWpeXkiiMFTdecjdzC
7keB57ttoY4EA+H/YEzgRkCJsFbPWPxr6EZH3UU2cfl0lX8KLjowvx2YsbQ6ViUK3NAp+PJKiJXN
AUrwciFUAtVkOQ6jtwL66x/1mMb8gOXhFd8hqkfLj9+8NmIeV+Byn3jnpUuKZOBiad40lEys6FpZ
6i7aJgKv56Mr1SYgkBYKmZ5vv8L4b4oFuE30qFJcMiySxVb2KZ8Gp5Aj6GarYQbGdAEUeIoZtPTj
mCajSOCOOY19sglv20ABR1BMiQuT1drJgeWxydmc+mdLdm2a2jr3KfAe/fGfSjpLqlB6gHWHgHvC
BgvPKxgFBHOwABli2e3DUY/R4Voqi3sNspP//qWe8GwkzYK6qRQ4t1S4piwjaYzeXEwIJ3dcO9sE
BKUJGvP7gbYa/xDuKbTrC/SRm7AaCpmBaQi9OhyqeVFxMf+Uzz5x2n1fnFmiFURWE0ta/HMcNHOT
xBd1l2X6l4rI0QfW0v9K0v5cQJkc9HwBCcpvgXLvcVZN3JWDhvj/qyp8rfyk0XnC3AigFooS2pQ+
KPWzhz7Z8Bcx3K80W4I6nFlFIDqrz1d+Bve4AkNKFDa01N/ySMmGvN1GwJ20qk2cVmN5RY6SJF/L
tnl1gg+W
`protect end_protected
