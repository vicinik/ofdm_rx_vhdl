��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`�����T;�x��Zg���)U�b����\C�]ȧ�n�ig���uWg����Gb��i>������o"V�SdsR����r�x�����5�%[x�
�e`J��:������D��%�֯qd�����D}`��н6a�_�	�ͯ�m�B�jpG�zy��b:�1v�cn��H���G�#T���n��-:��L�L�;Ha͆{���{~F���pJNG���&�P�>ҿ7�Hefv��po�ڐ1��R����J�䬝|�-�|���/���'O���l/��Tp�i��7Z��Zx-~�P\`J�{*c]��RȾ����%�T��I���՛�BK��W�1A� 	g�ڸ�ISGgEg�؀q��sn�A
��k[۲��4��IN�A��_���-{���9+��,5$���X*ч)l�򦆖�=�
⫒�?������~o��5Sd��[���m�Ȣ����/?����ݨѐ����d�<a�¡/QE��N9K�(VD�0D��]�pDY����U~���y�\io�����`Z�.RZj��+�N^B ��H1Ws`K'��6/�Y��P_�O���Q�Ru�VIy�I6y�I�1������ݺo�n9,*��cvt9�X$�x&+1F�]�|��wE!�[�0�YP��4��6���1'G2 ���Kw�_�
���'�ޘOn�q/��y��Yi%�q�\$p�*��uc�����\�4���J_U{R$�c;�O���[� �Q�}�#�ρX�����+��X/A����� �UgAqw�"��b4Y5��*�����]�9Ez\W �~1F6�\{�pf�����G��YGN48皖|�B�)�v��P���y��Wmw0	r��P��\� Ta��܈���{J�a���yQ��讵Fox�kE�]�Ҳ�S1�0Xg�
��O�����G��2g�؀�0ڰb����T|99�&�V�ǧ��O��_K��s�mΗ<�ҭ����Â2@���|Va�tqا���ݺ;�?X��#db��b3�3I%����e����h+��;��6p��,�E�"c��:�7`4�}q���6�B����	��큚�t��`#t��b₍���B3�4 �R�>��NS��H�@�v�
0���N�z�:ҥ]��"s`�8���t4p�M��1��v5����Uy!bJ�l�&��)���e�h������(\�̎��Μ�u��װ!̏��4��y䆪A�� F aٜ��u��;/�>OvR*,1�-Gf$���A1�_�A�Z���8��e^W]q���*�n�Y��G_�x�
��a��/S�^` I�{A�5☩�s�I�^3�p�͂[/�A]��w�^\�w���vU�ܩ���; ��>/C��}�P�3�Y���y��0	��p��8��������tW`h 變�nȒ���v����!6�Fѓ�/��=�L�`���6��}Re磲Ø��k�[ӎ�Z�.�q�]k��D&��7�_������W6�Į�RK(�12��1�4��"3�^�*����߯Q���G�[�L�M��������>m_f�ϵL�	r�ڙP^��'QKT�5D~d/sM;�w��qOH�'}wll^DOM����W���[Ğ1��Z�r�n2���+�sVu����qX�.{��3t�%���g���-��V
x��c|�(��;�[���׆m��:�m�}����{�z��x��%XJ�U���MRq´%�Wi�����E	�o ���h��,�i�~��z�&��9o?4)�����!��KD����x�'���JIeu�F��)��S���T��_����I̾���G)\YN>B�SJz�vռ=zz�d�"*׻�T��m>}NȢ@\��C%�F^\FJ��	����5+0ޯ��j�42��R��0��닣�2�Yn��,���xl]����W(�O�K��ܯ�"
O��mZ�l=�p%�Y2<��5����I7֧��ϼ���Pb�i$�IQ������,�t��=4=CN���(�#C��A���G�M���y���Zχ�p���Hi�ؒZ�O���k�r�����KnܔE=��`�Be�B�]������M��ܺ߯V�����zD�LK�v�Ȇ�2�y�ybɄ��K��IA_s]�a=I�2��~�m�����;����wM��N�^��y��^��0!�$����r���i lK������R�g�/x�������C��2w	;e����r�i����G{"\��>^��n�]�=������;@�~	�uW޶ƶ@R;W�N��t�oKpݵ�pTZ��k�+����!@��8�Ea���Q�ͪ)4ԍ��s�#����N��[$ӍuvZ�A��lw���R���-TGP�q�͏��W�a��+@���B�<[Ps��7�|k|���Sg,inb	�������[�/qc�R���:h��Wy���lV����n��#LZ���A��-u�� ���*P�g�?4�}�,Y�����.&zyG{4sm%/�BAYY���ÃcI�(��G��z��eri���S�i�Fk�̱x�I����U�ܠl�����m���T�H����|�,����Sⴋ�u��"�.U�Q���5�J��Lv��6܃^��T.�ѧ5�{��V4�,3D������������4"��-}䔏&-�ir��H���^��>����6+A@/F��~ڮ�>��zs�t�~��(��OU�ǸU��+�R&$#t��%D��T����]�ba�-j /��+m�����+���uwmꉱ�x�	�DS�w�˞�si�'�|5q3 o�$Իd���f�45���[f6]�[�݉�B1\��3�)
����Wc[6����ޜ'x76(Q[�����ngR���x�ʠ'�7�R%2�I�O�/�q/+�ͮe
�f<�g>� ���P�y��p�z�9X&#�����|��5<�Jnqᮽ�:��m����a|F�:m ,��١m�E�i��O%eh,S;���-ɨ��G�`��c�Xba�a拵F"i� >��UV�Y���>)�i�4~�C(�k '��.��s����Ef��	�<�{K�j�q�R�}]u�g �3.X�e���]��1����u��������!qJT)�:xP�B��!uJg��"�FR�;*V�8lZ*Ǣj�8ɀ�suVpJ�띹�_v	'4U0^+(�ؿ�Z���0M��x��I�K1]�,\L���c�k�(���o"x��x	�ɛ���_f��[9���α����%���w)e�SH
Ry���]W���"y�9��w��!�+az��Đ|_0��c�����(Ә���j	6���A�W�C��D����cP��kX����~�c9DG���v� ���!��3��w�ؗ�<*.��L.�>W��[kW��T��a��r��ޔ}�*L��ξ�D��u�yf?]����p�r)I�H{=��>������ȜM>��`;?�jN��,3�Y�9��C� �]�D˪�NO�b��_�'ȟ&���p�P+�^�C��۩h<���2jU,�OͶQ<�����z:���G-�d��p��c_�V�}"<�h�T����u��� g��	�1��0��8]��%�á������
�zH�C�HO�a�����9t�o3pVD%ߠ�Ï��cp*7_Yc��m�b J�^�ĳ�ԇ��:����ޭl���Wa՟��"�곀-�![Q�Og8���Oڍ�uS����ə�x�;����[�	D�d�,�X�%2(��31l#�G���*kOr�z�Sͪ�̎�V���aJ�\$B��$ĤH��֨�U�K0O�O�LCH�_*Nm��_4���E0��A����e���R����}1�����ё���������:2o�@�}Un�:���su��$�g!��Sa3b���~0��d�=?$À��`���*Q$�?�XZ��wJ�ڔ����l�͢B~��$�L�U%P�	}����@�3�WW~�F�̼��맬�E$�iH�5L���7w��S�ha�,�e��([���Yt��}P��2���s��8����2Vk�g��)���q�~���5�&�Z�q����a|J�P����9vZ�ĺ3ʻ7����#MF ]Ϣ��d�(7)
��z��:=V�-��)t`��n'oVPĭ����IFW�*�t)���B|�t���^T{,ܻ�hM<���2S��^R��.h��2��1[V ���6�e%�޸e�%�*!��}���f ����һ��ɡ��S&��H�bv�"�:k��
�Ȭ_��������7
�f;����W*�7��ܕ��K"��_���x�u�j�ک�0��:̄��Y؋Q����A5"*3� VhLY�t��B�?t��J�`�C@-��| �7�4�i�1��{��S�a�7������;^#dd�6
TPRf�|oa��L��O���Xb�as$ӠI���
�r'�;]�Nj*9;���G���y�B�Fd����3[O*/�Vd��m���k���|)�Ӌӷv��^�m��|aq�S�w��g4h80����/���#"P�Ϩ��8���P�
t�T��	�ܳ
	V'h6H(�{Ѻl���+�_��f]��^Z��Z�U����$k�d�>D�E�Yr��f��=fQ;&�߰l헚f1#��U'����rdk��!-���R�G��5��x�j+Y~�-���h�T�/Vg�D��p��D��2�iȠ�6$��E�q������{���q��J���D�p��o�����9�1wc"f��E,m�m���x���~G'b�.=d�x�tQwr����TWO�p+Xj�|;�!�/�!*z:d��J~��R"�C��*�5?���:Wf���Jml��RӉw)�)aW���^��G0*��\aiF�i+�<����BwC�횞�<Z��	;�̸���C�B���
I
���6�k��I��@]_���HIY��!mh��A ���Ĵ��jW�a��V����ot�-�O�C���%��i��� jwxg����XdEtLJT�l9�~تK�
?��=N��p���^S��e�F�k����(�nC)��~k��{g�y6��`<X`B��o��V%�h,���	�P옩OʹuG���� ��h{
�y�_ ~����d2�rwuQ�!~�G���{��8����c-<�n(�y���	:�� �0W�ۈ�(� ��k�.Ѣ��j��Yo;��t���m�D)a$O��df�ܷ��E� ��6S�CZ+<F�{�O�9�0��n'��]�>Qjކ�Y�`�$ţ,k*�J���t	�]knJ�����paI�2��4ۊ����(��ň@�9��pC�������W�,��w��Fh�}���7oD1}�	?�m3@K��G�a�i���ɥ�Fd��%���`67�E��cj+~} �vl}��f�+z��t�D�b����c=�S���nB!-X��=g��{��H��[R��C�#�x�s�E��,�,sb+Yn�K�W���EA1�ʙF�ɻJ�&�YB+�Q�)�XÈ���	�gпGEZ���ZSz��ٳA۲K�+p�H�#�A&��D����,&9�x���״ݰ��?�{(�o>��Zui�3�JݝɃB�����]��%F��z��)%:��  �a�&�S�n��vߕ�-o��l)>��d�S}�4�+B����@Dڪ��8�'�N�E��
��{�4�㪕�d�����ӾAޜ�~��)�mG��hM��b�g�?�ŬmN����O�?P����MF{t�>F��쒦����?UɥXϚ�&+�;��{��a *P�܄ y_B��q�[�6O%W�쓢���y틍XT�04(�V�U��YJ'r�=N����S��ꁈb��m.�f�f'j�����3��=���°�����Ʉ(tkE$*�R]�N��S�#(9���?=��H���>i�5��^ٟ�������[��!����Ѹ�=�Kb.t�l[oX�۞Yc�j���:2[I2��h�dY��{}�61�JT�b{J��4
���C+PN熫�*^?�#� �wo�v�ޗ�%�0�K�mr�8��1a1H����=ru��IÍ�$i�CI�,{��XR�N��W�x���<q�8��M.�\}U/3����0[��ډ�)�qe�)�>Aȝ1���_��gy�,z2���l&�fp�nf9��,����W�����6�TyNпu>�0�Ûpk��-L*�X$��z=@$��c�?������[�a�Z��\���&�`����2���3(gWFຈ�Hm����Rm�m/%R��,�����K($5�I��=ɛ#��A��k52Ql���y�o�+cr�<�s�Ze�e@�c"Nj��v4�E��lM���$D�?��N��̑��K�˹ƗX�	�Q���<p��)cb�E��K�S
�mxe���4�X˾�Ӡ�~�P���&��ȝ����2x!�e��ptXaDA�C���Y������NVbTcC.�z��� ^��M�G��>A�T;��CW�\�������qḜ��oӑ���c�\��;>T�Q�H�wzq�#���J����?u����E5��<�75o)ѩ�?�u��m=\E`��R�	f�����5"���r[�a��Σm?y�,j���������H&B�讦�ۘ���eDZE L���N��g|�B��x^J�g�p:<*���;���ɉ�:A��M��h:n�m���ԃ���Cz������u�Ebm*��#˧ �O�u/g`�Yc�ZC�H�!c*w@p�g�E���	V�*r�iѫ��ßWͼ���Jȣ�i����S%�ڟ�~r��X%yҘ��)9=��l��fO7O3N�"?�a!�}=�\���K�kj�+��5��b��Tz�C Ґ��d ���&��6M;���J2A�� �s�ș��|�E�.E�hd�d8�g3~0���ٶDdȏvފ�t�:N�=¤T�M$IC�x)�D�c��pJ�1{�ٶ�%�������H�Ę����o�[�u!;��*B�qGM.��U��*�LT�>?�]y��◩�qZt�W�z����uS��S�,��֏[��t�X��ef�D���j]L�#\%@� �^T����3�lݟ�I �c"5�Ix`�uۃ��r�)�m�|���	�*h�������譋@6|l� �z�$ю�I��	����d����މR�7��&�/8��cꧺ���-W�5)-�.�/̩��@�C���wٞ�d#��ɂ�]�M�)^#���o����Zʮɑ���'}d[Qق�݁�{/��ی1&���=ǜX{�e��6e�������t�A��#8%����X(,�Uˢ�$3�Cu����X$`�^O��v������,w�/� ���M�c��z$�65W?�����[���x�:'n���C>!�v���YPe�sq���&h)����}�P�����M%����"4 �v�T����l����ؓ�qf���5���3'�w�o�*�������g�'#�nԋM�$��4)F��ex�T~'���n{�}�A ��z4�u@���A��Ʉ9bT� V��'��n��)�+�9��=5%���_ o`� ��V(��)YK24;>�-��������$�׃f�*��[ ��(��릻T�����(2{���W�����B2C /v����Eǔ�ν�_�z�R2 ��V��k�["5H���}y�G���ׁ��k�ܭ�4tk:�Ǜ5��� $7��4�f#����ԇ�����EgO/V)&{B�'���-{>����P�ЉTAQ�N�5P�p$��*�,$���x争�{��訳�tT$�w[S�WZ�Ϥ�/�Oo<��t
(B�O2s'vzSdٜԤ�,1�m�>�[]Ѹ��L<:Q��$��{��K�7?��V"T�1���'ŝ#s����@�$Zӌؒ�gs�s�;_�1�O��'�6�I��y�L�X�!e��g�wJ�Q׵-4�0`��gg�w���z�`���^sg�!p 稡a<��F`���&�s{��k��`tS����g}����}�~{���! 7͔qL8IW�z2��VN
pr{ө=�sz8�5E�F�\v�.5G�@j;ժ�A�e֔�=�k� ;��ő����"2�"�U������s%Z3;��h�8M�%:���j�]��Ҿ�M^�>n�:�M��M����ߌ�Bp(����M|�%cs�T��{�u܌�L݇����6�9ښ�d�*��:�*}] $R>�[לn�0�ǂڰI�a��ʊ��b�e(��s=�G���s�vO��P��X�ܰg�m~��Yj��k�N!g��߆Q|�!1��p?p�}D_�e����|Q� @f��T�f�YW*��Fo�=Pǽ�#F����,�����0�?_U���B��.�Y-�kU������ m�mq�8V�r�Jb��E�"TVI�/Zzoؒ��#W�OL`�r���`���!N�`���k~�Y�U|]���
��x-�����%<â�b䫷������r�;<����J�R������,�Y��T�I��c���U�^L���Yu!Ö��|I�j�@pLcg��<�������y�R��`��@8�B�Td�����e��9η%I�I
�մ	o�*9�ht
��z,h�VG��[Zw�'�'+jӮ�^��R�=��+nAsz>����r�ْ^b�(fY�j>��ً#���^Q�wYnN�0=��$_2s_��$#:�D];˖�k�Y�6�N#)7}	���f�䃝�>�R�Z� �H�a�[����WF�������h6�&x��ɵzޔ�N���5�T�5����(�1�4}x�
��8�l�l1T>���#�x[�GU��^@�p�e�� ��������`~�YtO3m?w.��H7�1צ�V�S0Tg��_��\ϒ���.yl|j������Ǆ�o�nZ�JE|��2Է�~���Jq�{�pU�t�1l�$��R����Ꟙ�6�h�K����w&�_HI	����3���7�+#ֿ��ӎ�QGŉ�(�#{�R���3E����T��(���B6|^Ic�.do�W��y��B�6��c!d_�s���~��S,�'��l��P[�-���.���WFb��߫b �{��A-�>��������:�n�@y����;���|�Ӎ�\p �Hǧ�Xa��E��S�o��B��i������M����+%�v]�7CT�W�//��m�W\������R�l+��Pz�.�Yu$6� J��`R�C��)yB94b�Db�e����\!���Ϻ:�7?���L�/{-6ϟ��i��P���T����+s�[<�̋��:+�
�]��v*�$Q~��)E�%^�S��`����"�����/��S/7��+N	�K�i�5/2T��'<ADH�OIj���en���
`b�!��/���#�����zp�R?@S{��$�|�(�cې�������%}g�rt���"�bz�f��L?e��n�)飰P�1f�6�0���)*^;m�*uQ�c��e�Ո���ުҦx@����;��xJ�U�'�:� �.R+q?F�$���3��&�s�z����ه������Q���Z�X�Y{��Ԑa�~CF{��zP(�7z���*�YM!㷙A����ˋa�~�d)St�/�w��w�������D]}r��,b�(�:C�4��36��i�q&�'��6���z�N$)(��e�e?�!v�.�#d��&���Q��� �:�"v�9=���Z��C ��{�CP�YK���%��d'�6�-���0ih�a�ژ����o �{]�kt�}4;r>�]~n%�ls��'�����FdL�ܼ�W ���i^:~rok���m;��4�;
L͘�E��jJ|���/�\"�Ǒ�йtdw+ʥ��#5��A-����p7�V, v���{��I8z� ��v�"�Rg)ߟk���K���
\���Ϩ��E����Һ�OAu�-�R9p�R�Ȳ�6ެtH����д�Z3���H�J��q�������VY�n�`}�{�y�u����	���D�
`�Q)?6c("m�$9�׃�y�kA֪�D��-YS6��uu@���*c����eZ90�
A�4M{�U�_k�J}X/�)�~��f����&A)�+����ߺ���2%(�Ԕ��.�C�r'��F�׉n����F'r����I���Qz)�������YU�K���lQO�lYKT!��bznx�-�菿�~G���`�4�k1�ht�b�}F�E����$�P�_��ފ̍��P�(��7�/�&��X-D/�6Zr����V����t-=�����J{��^κnP�������e!Nڏ��j�u8����y��N�[�{�N�y� :|h+}`Q��iN(�]0�����f{�.�3 E��Z}�5ƥ*I_b'�dܿ��K��.a���(�S�� A��nv��$���n /8c�W\�3���fc�9�:��V��&�.NĶ������1�r�1xRӌ���s���^"_��7dL���Ie�Gw��K��
u�,��:4R�D��y��$�֮/��!#��[|��T���I'g��&J?��6*��'�?��/rX��?Ol����g����@���+�趌U�,|k��s�W�0g��>p`���R6j�>��MUMH��P]7V�-�h@�|p#l	�ӫ�I��G���dC����-������R��u��aK+y���?y������27ix,	�����V&�G��5}���@j�1#����9��>��Vwǰ�0\�k&������z�	���kk[���<����(�[=ok�hg��X%+g�׹u�� ��� �~G�j @�b�Nb�{C���/�+���3y�����k7*]�X�:��*�(�cٺ����� �ъa�-�k� v�ߡ$]���sl�d��Qýo�b�#Ю�=��?5w���	�kA�����+�$���Uð�ԙK^-�"�K��'��h�[I�"m��a��^s�<8���7o��K�w��Q9�uFR$���l��H�������e�~�ϒ(V�RbØ�|��§�T��FN��Ĥ��W��N�������uw^_}w�i#L�����P�8������������j�E����w����-A��Tl�h-��>�����]T5��Pk���f�.�:e�#�z�C6�B�Qwq��y�&l��Ӭ�u^�>4"j���'-�Ϯs���싈z����mRc�nK����cY8�-e֝F7ՈLغ f�~�'����ԇ����C
���=O���~n� �Q᝻��WB��q��&��$���!�*�:���G�g���D�숐Z�S#(�t5�U$�����ì�NW��u<0��)����-J���T_ki]�矑�匊|v�ζ� �|kYJ��P%E&R(��F,/v�'D���
�ۿy�ڇKW<����IC����!~C��Q
��o���)o��:�q�Uō��o�!}�ql8S�n9N�Ȕ+�o�=��>E����(uO�n���r�ç_b2�`%k~H��� C�_�\5�̽s,�ƚ�U��bR͎��-��68>�z�G�����d+�K6c�+�[���'N�S��jB�{�	U���ϳn6+����j�։&d�������/�/l�[V�\�,m<�E�k�X�\��|��;Fa����5K`]��^Ⴍ������ŭ2�r�MY���s�1�N�7���N��۠fM�B�兙ak[����)u�GΪd
g����e�;�?�HW���~�Ƀ��/�U4iy��H�kﯻ?gi�(v¶|� ��N#�����-��-0��I=� ��S�|�nUt�#��C
��֢�����7 &/�h��*c/e�}�o�]�h���Go#����Z{'��<FH�ʯ:�7�/�^w��g�L�Mp�i�����ek;�U��w<6���x���W����iU?Q���=;:&��y�Q�����8��n2Tj8"4[��|S��.�����mUV�_ ?*�Z�#��Eq�m�jIA����L��v�A_��(3�x���7��:G��d"��p�O^H3 �&����z�Y:�A��P�lR�D2ѶQ�T�/��Ơ�Hr��f����I9�>�X0�
Q�֦�B 0������a�?V���+r.�s��xժ��_�t{�x���s�80�gj���O�^�hl{�\mV;=�#�l���.�c�4`��kȹ��˹��}�V�X�6x��;b��{�$�!���{��5�=sGHwY9�>�_�� ߎ~�9Ώ��M�f���}hp����>����7�E.;� .�:�B�5�s��Fx�>\�A�!���Q���������xq�j�nt��j�o
J��:6@�	h�Z@��;�8�����SK�*=u�cz13/���xW�*�,���oӔ��.�_Mm /�]��O0�J��W:��Ž(���L��v酤 ����炠lNl{��{�f::�ҋe�Bk��.�_c��fB�MS��s�C}/�;ð;��K�-ʥ\�>[�{T�=�u�E�/k����5�߱��� N+�دk�ۏ5o�M.��T��mI:��r���ˀF���q�e��E)9�>���r��8͔�g�� \�c��I�ѕb��|�D�Al�%	�yb������?-�����'����4��P��qxQ߭!_��iH�g�`����c/�pQ+��D���Nh��De䚆�{�aOM㪴HO����%��2	�sQ�)��A,0c���!d-�(�h��s�}vReš�;d?�3s�'B芿��T�:��Uz�K"��B6�����(�,P���oq|)GH'�A������ ����X��a�Y3�ڿ���A�c{(Z,�H���3�D��K��3�*����aJ:�K�"64�8x!�>��a�������n��ۙ
��)���a�?��t�xD���of��aJ§�?S�6�blOS��}.����'�/�)-n2�"��>�!����Ǆ�k��h�u]�%�)�WV�Fv9��,�x�kX汧4�Z�86B��c�^�-k<�;������p!*�b�w[����u��F�p�8
1�ҁ*!�����(�����`��I�C��:�����b�w����V�W��f܈?�R�W��t�,L�����&x���-���$�`�4�к�@1:�}hqI8*����5��]>�	�˺@�R����A����0!]$q0D�iS.O�Y�}>(�B�P2ȁ�f�W���;��i���Ӯ�ӾΗ��|U\2��m1����8�wF�YX�j}���ʴ"�aO��&,�W�y[{��D��1H����H5����a��j�I��(n�����JL�T��3�P�^�nɭ�X?q��T몷0���b�N��hf�k��k�U2�H��X;�=�@�:��Z�Uc��B�k<�	-Z��=,T5q��S�WJA�v{d������=j�4�<�%|K�#�
zkx/#�P����S���7e?�W��"��z��0����=s��֍�L2B��������2gc������2g��>�8��H�� 2���W"I�!�D��M���6 ���2r�x�	iOߢ���v�ƼEy8G/��p/��TI,8t�,4�V��Gpa`�^}�>h�(�PN,�Q.D�T�-��Ԫ�D��C�[�{YCY[����%���LQDQ���n�Z2K:�a��^�. l�u��k�'U���2h�N��!7m�4)�����;��77d%y��vHm:ӥ,1i�h�k{�����KBZ������2Ԁ�u38>?W��U����r9�B�U�g��i�J�[8��Qft�
���d�ܔ�29��=��
�y��9���z#`]y�wⅻ53�l�V0��C[�����s3V�[l*��x��`�X
��1u:R���L� �EP�Y����1�G���u��䆢{�\�&�3~�T�p���1�9%���f�O�#L��)1�%��%1�0�}���酞J~Q��UC:���=j���^����0v����b�i�U���/CA��Dk����3z4�����1y�|pI��V�nĆ	����C�h�R)+��ԑ�t�}ȬL�m�jn4Ox����j�0�XE���F���b����ųa��ț���_J�� LH��ˋ��Ƀʉ�u3�;ݓ�f�jr����y�����[&�d��d�v����*ә�L:Vu;�=�<�Z�Ql��⵿�l�Fk�W1���N�B��ex�.߄�5����e)V��8��B�p����Ό_��S����Ʀ���P�|�<�!�>�~��&�7��d\%I����6��{|Ӧ���3��8Һ��H',v�_f���=����(�ܛ�[D��ȱp*�Ecz�4&mv(Tu���b�1b�$�4�qd"�w%�2�z�Qw��q��{�w�h��LO�K�8c?�bq��%"���`��F~����ð���]�F����N��L��3��$���YS�dGnE�G���u��Tp�氁[�Q=dzo����Ce{��	���l�R�ʱ��x"찂�x[F{���C�i@�>�q��ʥ�]q���Fp�@���{J6^�F�~\�LxMU�.d�Ȱ�!��r'p�Kq��Z��G�u�^���RE�ʚ��6�?[��� H��AR�� RٖgY�lQ���@&�����g*ek0ǜ�H��B@�J�1��䁝�Cw������O~����ҍ�԰�� l2u6~Ya+7��Ϟl[�L-!Ш$�R7z�)�����rϥ.���>�(놗J3�?�;�A��4��J���������X5�n}���� q�t��4�"X�����^�a�н۷�z����x鈒�x�U���IL5�� ��ڮ���S��y�tWv:���u���-ws�]�6˱�mt0~�N����J�E�+ճ/���8����h��;,�"q��� �v�d���t�.��:њz*��Z=k!B��L4������X�#Q�C0GtZ)�v�v�`y���l�q�j%2��_���_�&J,�!we�fT��Y��;����h�Fk�u}�����i	w��V�0���J���;�Mf�ўh�����4�1�E5�T�x�������T,�������Q�qu�2�w�q6u����,���ǀg��&9���h_EG�ъ+�)��}���=)b:����	�HA9=���u�xqO\�(��h�P�V@�kWD�}���V�˾a^D\��h�t���w�6��ye��thS`6�M`�e����Z���!l�ٽm[�d�����j��G��r���ZO�Ե�t6M��
�����:AU�_i1��az�HAd5�e9�D�2���e�&ϱ��މ,�0U2,#)�U�S��6H�@��-�dq��܈5�%�G�(/'��؊k�C.���O����GR�E�,�,,���S�1�ܲ���:"���긕����^؄���$�XHA�{(`z��Ş�o�M!2����8Tm������;�@zR��j��}N
��������G�#��fA���+_<R��)��0]��_/6i1�o���KE��:8�bյ�R�Q@�}y:π`k������F����N�b�ON�K���=u�B���q�b�
���#w�-kz# �򎊗YK���FQ�w��d�F���& ���,��)�ܟ^��Xs~��r�
E����j�ZG ��s$X�{�k�0i$;	�����)�-�!�;���ŋ4PX�C�<�)Z��Y������o偅�DU[]k��rT_1��z�G]�Q�R�7бɽUIf��ͮ��� L���Ӆ�@�>�h��lߑ}-�X(0'�X�uK]<L��.~�u��9ފ�P݃<F����1!4�f�ZA��j�*o]�5w�M���$�Ya{�8�ԟm�k{�\����4dӉ��ZυtQ���J��P$e���X:g���@/��ȏɏi|hT6������ڌ(�F������Kb�ȲD���m����J\��|l�z1�/a&�H$����)�[cwA�L�� �SH!��d�[���J/2X:��N�Ճ�H �̑T��qe�����lA&�W@{kqIL%��h�!�c�O��j�D��@��
P��Vp�-��iV�X�(�T�;�:�3��Y����h
��z������+�X�s���o������92k[/엽 �N]��!����Q���\�J.��⊧R����Z;Y�� �u��\!Ⱦ{$����ۖ����F(��y�l���z��j0��D�� 蜎�]00H	�<պ����ndɕ�^��L�����X�i�)��Y\�濂�,.]�5�@���+���hF�{�s��}"끘�J���Z+�{��������+ސ����?>0���Q�1�D���?�m
9Z	��N��k@Hi��D��;mu� �Y�w��Ռ�MR� g�~j����W�(jh"���|X�aȥS	I�?���@����Ew���L��V�e���7v������.�Q����͌V#��`l*$	��C!g|v��=Jv
�y�V�fQ��\����,��˻6r�"W�B�f���~��`Q�Դ�5�����p ֈ�ve';@�X4��W�|\��b%�v"�D�7��&��t�	p.`S�'`�b�a+D��`���5�>�砙5܉��~LC���������Z��/��UXx��摞SD��3J��� �#�g�T���~�O�!8�\7D��2*�K׋IFPU�/�מ2��q
�<Q;ې{^9����EM�E1���Z
4L�����y�<W>�F6JG�U��ހfBd�2�NB�9I�����c*i��.�m�����j^�jt�g;�0۴m��H�	�#��H��
gߒ�7{(�s=M���������E�0�uO�p��P#%ƃ�(�I��.���*�F��ȍ�+x��M��G�9��'�8<r�l��Io��#��]�{�1(w������L���e	�5��j�O�^k�]�thCӰWv�>��K<�{�D�y���X�`�a��_H�y�;��T�2��$1!�t�������`��N���7��x������F&:Y=P�R�l���%�O̥���M�^��`��s���}�BÌV��������E� �N����<rpW�ze�;�xU[��1��>�B�(�9�dMU����p��J~e��3��lr���(�ދD׾�Y8����svOR�&� o�#rRs�ph���O����Q�֊���q�co�P�*��|���*�L�l, }��C�����!Mz��M�������3<�^����
	7�ӗ������LZ%���m�!D�Ÿ��-$����Iۏ�*y��z='�q_����������n)-:W,�/�tF�ˤ�p I�B�j]�r����!�hH��Q7bLJ���c���c��,x?�"#�.^y�A�kJ�x�)S.m�Vf�`-v�.���4:��/�)MEn{9������tf�D�'��
��h�n�������-���D ��gׂ�Ƭ�(�,�����Di�<�Kew'ʙ)�n��a��G��m�����}(�.x����}��!�=l� ��A���c4���P��O���2+��}������>S i����zhdK6T7����(�zy��
��V��Ny�G�h�CE�Wm)�1����֣>�Y���D"���U�`�r[��ε"�5��y2�nv�q��� �P5��e��V��2O��i����Z���}��[����Q] �Ufs��,��q�[��	d�#��S�ɥ���q�����}m5�D��J7�\�=P8���sy+:�/%1!<<O_S�RVt�GJ1^��dLh����U�@xa�nz�b���e��Bu� �M�a�~�И�4��)��uuV�!��i݄*���o�)�j����}+X�8�EȳR8$�i����Hr�G�?)p�y ֿu:�\�2�V�Q����E\�	���X��4D�ǃ�r;��6I�͜��Q]�ir�� �p���-�'�C7v��a�	K��w�7v���F(`�������������g�[�"�T�`�[p��tBŵ��=e�� H�@�A�m��wb�%�)b�)�����z<z[�"�H��2 Yh�(~YPr_�tp&�%b��^�A�"K�6k�E׎�C���s���477��sc�����H_;L.���q^�/	�3\��qp��TӨ;��.Q� ��%ޔ��}J�I"t��kTG����$-��5wR�ʆ-����i��:. ˺*� -�LZ�E'��x��r�gԤ�2�Z�BF��L�WAD������~#�.��b��R�Nak��V�"�����F��X�_9��}�ʽ*MP(�E�%�)��<�o����h9N2�6����0O��C`W#�)�MQ�' ��F�9{�@Z��lT��m	og�{���d�PA��Y��Z�a�/��c�wc���٭ǒ�Ě���+�	U�H�t�XO��[�m4NI#"b�@�{�����g�6�<L�X" �o�U9/����KPFjv��in��BȜ6��ϳG5h"-��3��-$EEF�.�L���K��XϠ��L������N\�;)mD�v���H��eQ����A���z�r1���.���Q��}����@�J%���eжR��|7C��#�p�.Xg��Ĉ���1��ҹ�p����\P0��!�4���Ӹ%���r荑��	�ʀ&Q�XY�i�z�1td��W���ᱚ$�Y�-j�����L��7�����H`�tݒ�`�oI�F��7@e�~y�������~.y�b��rx�
ONsr3�U<Uh(���Ro���='��T�V�r��y3�+�ڟD}��,Fi��!v1偅)����G�㥹�C[� [���d�b:4��d�9H���&���Uir��S9�6�N}�TaeKᆺt�2Ma�r��_\�Q���1ņE휶�oq����{@�Q�����Iy�-����s����c��=̚L�怶�I�i�虧�K�2a@ T?���IT���'�Q�XS;f�Z�Fõ�U��E�HкN1��?��P�8~�AO������.i�}�3���K����[*�ys��սx+7� ��/ٕ@E�-{��N����_n�����R�{]Q��G\����#�#�r��s�'q��0B�J�j�Ss�Q���Wk��EdU�a�)�ޢέ��ew0�����"���mTRK��mp#���Y��ǰ�nrH���F�K>3�g��p�ρſ�{��ߙ����K�j���[�9���EG�ipɁ襻撹aE)*��+AX���n��]g"�^��P���;�����)u�M���:����+O�岢$ s4�s[�#W��c���)�-��\��%�!��\}��]�Pf9��J��������w�H��=���^��]Ŀ�G�6�q��'��WO���t&��+���5��/V�w������9k���`�Z��}��f6$�\��Ve3�����S�s��VoQhm+�U�ű��v�S����sE&��)��@�=:b_l�f1RC�:��������l8����C�⸈�YZ�@��ٞ��&����۲��NI��c|� ���8��ڎ�c�c[�"5��9���iY��30��<]��yɀ�	i|ߪ��ո�����x8��e����p�3A�/#�O���+���u�b밖�F"RYN����Kb$�P^cGN=�<g� ��^�(�B�J�|�[F^�c9���^q�`�5�����o}�7�b/-}~=������#����/᝔J����c@�n>/E�]XWqv�y|{���E[�Eyi��������:G�}��q�V+������-y�v&��qmkB�\��b����rĊCUq0q�9�5��Q���*�{]�0��b �[��=��-o,�Wk��_�|S���k? FA@����LF�HK����9���wYNӵ�Q.t@5�V��9�9t�Y䧢v�+��FY����%Ć�wG�rf=���V�-]V��Tؔ�p�bo� *T��x"(�����@[�2l⻐�S�	F�@jČ�k!�%����'��B/9L���{��8�3�EpL��0�~���ps����	va�$��(j/�����в�t��HE�96�u_��댟�{�}2%C�!��g7SIyBO����^��2z=�o5��y��p_�vT�&�jR-;̪��:�����J��Q�S��p���ݦ}�-$E�>?x��s��\��傆`����n�h>j}��ۈW�N�N �%BCǙ�حزXW��_RkJˊa��
���'R<G"^�X%"m/vI͘;�OW��_>"�<��B�\IE��>[�Dn�´��-��
���w�XO�PHg	=8�;��gx�����Ŋ��l;茁&�U'DP7>��Ս�v#u��Y�>Q�����$|�d��=�:� ɯ1��vK���ʙ�"
�j�k�� 򵣅�ԉm��V�4g��|	/'�|��G[4`
&���sы���V���H�V�0�|ҩ���^'�	�Ef�۝;O�/�E�	�@�eh��@��x7�G^{��؁�!�w*�H:�{����ݕf��1��1��f��]�#�����,��΀��~�-H�l�īoi=$K��@�z'��M�(�9�^�S����hw�!����n�>@��QIE�X�{�}<�ʽ��A�ZMA�O�$���GgS�l��>�fJ���u���ˑ���5���$uel�����3�	��;wd�p���|���
%?u�lQ� �&��b�zp���3"�4�o�C3���r�o�]�����S0#Z�ްӼ�g3���H�%�j����)�H�.p	xk��f��7���re�]漝V�O/j{|n��ỄN��>�?�)0�R+5�mF��Zˈ'���A�m<��2*�tzj�)���3aKN��adjf���rl���3i�BvհCe��1Z7҃{)*^�%��i*|4i��:��4p���k˶S�~�O��7�bM��6����^~�_�!���d�P�4[d�ގ��k|ťC�a͌�Kx�N�b�W<1������dGʙ��E�5?�ov�`dvlT��	F�4�����|_є�΅ֈa�)�⥍'R��h��Ap%������I�0���\�bB>N
J�U��I���Я�G��V���.�j�T�u��7'f�(�v��5n��wV˚zsV_���I�:�
l}n�T�� ��8ż���R��x���(���a�
�#��(��B/@�¶�[[!��U�T���t��Po��m�\j�G׆
���O����y�sj̐Ʀ���ir%�	nL�H��=�-J�7�U���Ґȏ�*O����v�G_�{���T�s#P�с�v��*g;�����@��{��
�o����f<\V)*v�~�cc��ZK�)G�7]�[PM���;i��^oq�+��[��#��(�ۙ#>@l���y��`)�[���-l��{���6>�ǡ	��nY�x�H�w'E�t裥_t�R��m�E~��-E��W?��#R#S���AH����<.����k+T�*�l�]�MB��o�w����sΔ�o�<�ď�o;c��D�P���M�֟��Y�Z#���J΂W�TR.��%o���J��ɳ�FpG�!����Z�6�`�Ed=�mO�ա�Ap�'���|W��`���xT��{���ӷ5,e�,g1%o�W@�ܹ�.׏>������h�)h�<�h�X�<<W�c�^b!����]P���p�_���Z5��:7�o�㔔P�G�h��M�)�V:8.8��$�P�o�aԨ�����z��Xk��2]�}���X��.'?�h��YI���%1F bǺW�Ы��K����t��
���U}�e���l�~@��ET��o���l̸�^��s�$�=A������E�O@ply�;��sG����
�a������dmS5�����jծ�Ȱ��Ԕ4�Q7�
* ��5�$�[�i�m�յr�����1ب� <=����^*��7Vtu�y�����^O�CrmLr�h�gyD�����x�]"�qmo�,��ݦ�͘����-D~�,�T���^��eZ��jD��D��:����B��9c�d�KW�4�P������)�%IZ����$3&G����_r	��:C�71f�w�)�_��*��+͡�/�/�n�a!.�*1P�H%�O���e@`��l��Zȳ¢#�����UGg�$��^�k���$�!
�	S��؆�y�c�"T�ѹV� s��|����M�T�0��ui�;T�3wj�\y>�j�/�m�����s�}��*iE���F�5?�lA1d5DZ�,5�����K��2?.�1.��r��U��n@[�k�� �~=�fnh�u1�Or�si�0z�լGh�(p�q�j9�ݮrd���~�Pd��ڜ�ר.�]�"�Ȥ��{��w �%�%���5vq��>|٨'��Hɛo��c���LsӉ�^;|�ͧ�G;���(�Ңu�GMaSw���mcý�OM�y!n�_s{�?�L�ȃڱL'�$�*Q?�ϴ̮K'�)'�\�?��)��rNbz��>�U����;3t�^:��cNhݔ���,��Y��\�߯�ζ�"�y��8�&���&ll�盲*�rZD@��Q�:��"�U��*'��u�n�����ז�l<�Q�?h<i����,�"4�#��x�셓L0�&*�����o	��|DD�����BuE0	6K��~�bO$$V���mܣ �-�|? x{��+\B��5x���o�������h��{䃔*N�}�?�
2j�S�Y�$�T��ͻy�B��g`7��m�9 m���!�&�O�˃�굌�4�qn-bڻ+u;���=O�yu���f5�����Td�y8����v�sc=�����-�;�x0��×�0�1�T���^2��xH�h{��V��Z�<��&ѸpZW~�o�.J���)��Y�O]fiY����\�%)�w蛾K��V;�_����Հ���Y� ?r�����q�m��5�Hq�h�J���-9f�1ꕲc�/5:��9&wP�b6ȦD{!KE���B�;��������C���P�1� B�y)h��K���g��W�.ǒ�������7�ԫ�*�P*St7�����`�j7J����c�)[1��`l������a�;j*-p�D����.t
Fij��0yH:@?�M	��f��:s�L?������	Y��u( F�??���7U�d�l,`}h�+(���dY�Ld�����C�,s�޾4��&rf�s�ᓙ�@Ѐ,�}�,�����[u7,%u����SI@��3�:cEzA�������nZ\[��X��+�Kc�>�D2琏'.�c�>q����9]����4`4��j7��tC���PV0�m ;_rǲ`���&��� eo=�� 9�o2=NZ�~�^I�/Ѷ)" �sj��9m���n{��h�%Ut(�&#I�~��B^��T>OD�^C|�7�H�s�	��boP%��#��Q�P������w�&�+��z���V�<���Ye���ghI���������6=M���}�Ptt3���"�h�_h�u��D�}XE�i�JE p�T��Ws�(��u��=V���Q�;��&�0�}�s���9JJ�u3��Q9��%��)��e>��GE��	J������x�cNL]R`���ډ�蔖�@��R�H��>W���j�<\IS:9p3���ə�7C�7�~�1�)4ӷ�{��} �W��F�wP�y�&�w30�#BG�u�	e��m��W]�H�31N��`�=+w��r����e���b���	�٤�e���W��8��ْ;c��m�'k����d�!
���[����-����Z�����,lW�L�!j����I)��킇7��4ťB!SO�������6f��6ʾK�P;�]�=������[R~��g#�-��z�m��#�^:��&�$�F4Yǥ�9y�����[OO=�d��vH�����?�p'����`y�wh?â��*aԚ�okR�%��?�^����e5W���d��;���K�gh���%ab?H��=����9��Qj���XZx�4y;G�3�g����u<�N����rp�A@��j�k_H7A	���5�YU8�Ԙ�]}�?nᖿ�T�����n��:�5�YW�¦R��~��r32'��Wm�bz���I~�ݹaE.��B%��1G}����!�|P��GVL�(�3�h���G����bCy|;UЭV́TO}�a	>�=�G�pM�d8�$� �Ӯ��-.:�L�s��B�q��O��:�F��^�j�rvޔL�q�7�J6��?{��5�O��) ]��*���*����}����C�z�.�y5�����"t��Q�x�C��۽z)��!%�!`���d	`�e�����̱\������i�<�;����6���7�4G{k�~y�0w�rR���&�L����uۃY��#Ō���'/�Mz!y>y<���q/ŀB��v�w��)���2�7�r�Q��U�9m�(�z��)���,��|∨���z4W���H�U�@7��{���o���UP*\t��T71:�V}���I����u�r�o����˸��yzv�ox�f�_�eR�ݿt��J��ny*.�YC�������?��x�?LM��Xf�X�	 fG� k,d��-�J*"8�����	���}1Γ6�ۨ^�J!9�A�\4+_Q��dݡ�fD���^ ���-
[v�o�S�@�A��G�jYƎ0��V�e���{M��Ϊ�m�tOғ�:� Q�o-x3>����TK��FE�;����Bs(��Y)M?�I�څ;K} �Rn�f�>0L�Oԯ�"�}��U����[�S��)��Y�T�7R1ޮ���X6|г�6�wڰ��R�0J�>�'ZJ>)�Qr�k��{	~H	��'(�|���h:��׋��Ui+�Y�����&tĀ[����MiaQ�WI�x�E���z�l�?�Nǵ{��я`�2<5�F��e%��͛L���Dv?���g�Ub|����獄ilFBſ�!�،H"n���x��v[�mX����������?ϝ���|WX�Gp=O���v��H�	��F
�j��l��9BZQ�uj	X[ڂ�7�	�,;��>��M�R�]��@�>
(�S�� �
B)��8�~�ǆ��m�2�ܣi"�%��b箻!��?1�\HΫ�Ϟ�c�ά9xUp �
��gXo�M����h�xY`,x�'�9��+���wF���r��������3�*�t໒�I[���0������:�+�AɏC�t�C7�7*���Nߟ�P�]^Q���.)��ݛ��Xu7ʅ7X��͋)ڝd C�U�̢U{L��r�@P=q;R����LlMXN�QV����}C�u���j=��h�b��T�Q��6<�FsJ/��c�\Sn�V1�X����J<K
H�b��͢A�)Ra,�po�aV�m�m�����+��� /���ݨKל��]lr�G��ϧ�%�@�Hj=ĒۆJ @6 K�^��,pIx��'��P)�12���j[`6P��3�MXM�c�׫�p�� ���l��A�V�KhEM�
U�}R\�'��,�P[`��R�s�	�qճ���z&����}��(��	1_���џjd&��T_�P�˔J8��i��f(�=8Ȗ�d#:{���jnE�]��s�t!I:����f�}}�p����r�݌-���q���t��#��P����^�!���(���=��bOdf����)礚B�09$t]t6����1V+�ZF��	z��֔R�<3�5���o&����	���
r�,�>vI���p�������/wRܸ��*6�X�P@|ly��8�nc���cX�eQy% �`�γRW]^�hSq��}d砝J�@4<����eF&��'��9u���S-+e�#d �i��e�5}O��_fj���`���S����}Ә�:Q�.Dj��:d���ӯ��\(��je�w�L����"�f$� g��W��ϤIq|����+��� D�,H@�����oL�k��6���x
��"m>�M 'ڠ��`�\���=|��S��`*�6��Cv(���2�����[�	9�1��u��Ϛ�є�!X�0��,��4�9L��0��'�9�W�t�E�$1��ek��}��٭����$�8K�Ή"��J�T�^!aZ&~��U?�M@���ts!)��e#e�jgNԼ� ��4颾��7��+EM����/U>��
���q�,1��hw?`��v����m�f:j��^}�҆�gO��~(p��)�.[��Hʆ�k<0�`�!��d)���p�PG�ի�
��D���o���	Y*�I뼏/���X�f��c��s�uI_cmgO�V��w3.�#P�<!A�"�[	yU`�v���X�r^9���l��8�9�i�3� ���N	��)^
p�l����.X�����{�Ә&:Ӳ���W��Q�o��H��c�������tul,�^�	�İ�r�n�&`p�uk��8۰�$ԵY`q�EN5���4�y!�\�F22�$��J�]Cân
����5�~��z�e]9
�J�K���K�̼��������L�'��#Oj#6\�����Auq��_N��I4F���$ʯ�3Ջ���NV��5@�=A3w�bD@��%���ރ�y��Q�"r:6d���w�gH��-�Lt~�lT�^RA��L9Io�0��i>��r���T�e~FC�A��*�^�����[y�g������`��5%�&�P�@m�J����~(��3 3�S�-�i���l�[�Mp�F����N�.S�ȉZ*�w��<��u��w1��s	���ց�MͤG�'���O�������X�!��k�2<G=ʢ��]~�Z�U�[�T�	)$2��/�DZ��g�{�� <�1`;+�A/����yu���(\��k��!Il���Q�[��z�>CN�w6*�*�*R��Ry�
�/Q���Dd�N1~x�T Fy�+��軟��W�G����A��92%���yq��$-: 	C���fu�����yС0⯕5ۨ˅�C9
܇ֲ�y�V���������[�9�ȉ�]䦼����[��M��]��]��~�q�b���d�s:mt��a8��74���m�$Dyx�'��B��Mj��^%���{�6SD�������1�pylIw�	�3`Fz)�.g���|�[D0S.���b.8�㨑!�z�!�n�p3��ߖ�&�	7E,$����V�"�N���3���;1��7.����*���S�V����!S"�f��7ަu��>�U3ɂW�HQ�d�����|�T�0.Bt+�gq��#���m�ÏH�g������W�@{�y��;/'Goj��6"Fv�U%�(J��gףg��e	p��O��C�Ի�c5!B+��a�<5�����ٰ@�H`�9o_�G<`w �*ؔ5���آ��{@'C��>�'H�x�a�
� +�{u�����������lO�/h�]l�k7����Q��ē���f�c��qP���z[	�����]�~�hrV5�g)��1C&�m	�E��˃��m�����A�@��5ޯ����.�d��f,CQٮ���͜��8�Dي<"OB��'o�hO)f^�|:��w�^ͥv�w��}�����d���Ȍls�)x�� ��i -��My�ha|�@[�=E(@��&�b���6z�����U���w"�����hx�]����[ qv����,OX2�W��J��X��ڪ��23������o!�sq�^��h3�pK�UW�k�+=${��c�S�G�Gͻ*`�v���2�.��!6�[i��q,۟BU�4d9�;y�Cv@��9������h{%�G�=4LMdL8������d�%�
I�5���B����s&��P��ʅ) 4���
���g��a`��t���nN�8aπwC�~ۊ4<�	R��ǡA�n|�iE���q���Pc��z&�g�%Z�����\�Sɭ�4@�$E��E��[�Zt�;��ZXSh��*�,MW~��?�"��#����(W/~d���>�`�b��m�y�`�榿�f1:���V}R����aK�d�h��&�@�o<.!ˡփ�`���ζso�3�����仯���5&��;S��L�)�J�x�j��d=���U��z4o�%��d��N��dk�x,�����F��o�C��$���T���{ṲR#�*�nW�6��ŗk4� ӷD��| eF�qQ�D��R��P����9���	��7��O��5|�������<@�G�z�$��Y��J�*���d;�2�'t$�F�1[�t�U������q%kķ&:)U�t��=LB��B�A;	o;�̊E�
��*p���)�R+ג�-5��P�)z��a'����VŘ�y�n�9Dg���ledyȱC�b�����2&aqƱh	��#t�u[! �^�-E��{�X�:����* #5(��,nK#ݪ����a�芐�&	Ȋ�B�I�(�U���)!O9���x��-���F�V�ϥą4 l[��Tf	�)v��7�D�⸀��7���1��5�:����^~����̼q�U*d��!^��%&>�9�����N�d�$�b_��o]���RF���9<�R�*z�-"r�tOeK�oڇ�K���k�Wpj����̷��8yYP��6�W�7�/Ƚ 2���T=�R��9'��:6e$�p��0v�"� ;���AiZ?�q@�G�c������/ݥ�_���bQ�g��" {�ձ��x	�B�r���|aN�d�v�q�!Ƀ�{�1:ȥ/�y䘎�p���W]L���Т��(ʌ&Xǘp�Ȼ�9m��#w�8T�F ��)VQT�y`,�/5��oY�J�����D.�	BkT%$����*���w:�ʦZ��d��N�G���>{&�
{�aX�5�-3ov�cUc��HC�Y,��pj�v+��i��k�F߹��GmIAA���>ꧏ6�|�ߗb̜�ml�[뚃0�j_������cڿp��Z�.�'P��U`?�^ǡ�a��#����)����~*�!�t�B����� ��H��=�S����4Jp�f�b�
?�z�L�`�-����ë�#�0����u8bs�f ��[�if�9��ꄹ�&O�:�a��H��-;�J�!z�svZO��6��N�ȗ���1r^Y׈��
��Rۤ`�e3+�S4<Y��u�m�nP�O�����X[�9-��A�z�Uh���_�>��hq��]J	�����b�Ǟ��y�]��:��,hoX~M�"�f��N�_g��dL��*�
�ց��V[��"�"m�sѧ�j�W#�R2 P��0z8�zx�9C�9��E&�ب�|ӲV��^�`�^(s)�����s���1�B�q�N�Kh� K��~�Gԥ�HJN{_��#*���,^ok�aH�ִg���s�L�+&��X *�f�����^K�UEx�J�3������2�U[�G��5���?���X����H�����%��J8<�$ъI�z.������ؼ����5Fk��`Y���E����A�p��v�M�@f��i�eۑ�ldCEyuU6��1�_O6�M�J���}�\�i�"�����tm��pb�b���~Nj`mD�:�FK�P&2��Ha���_?�;���w"��
B����k~���aW+�6�P�&�u��^/e׸W6������>��UjG��W/aOD"7�8*`Wi���~B�=��U�]��/C��%2(�+_���B3�yu�O���ԱW���u�9����=�od��:�A���f��5͏-IK����?�#��5V�R�=����KBq9P#u��$q2="��[&�*�&�p�����5�����xe�=<�cU��*�'�die�t��#l\�����'�zb�UY���F�*�]j��A�K�� &TN���ю�v�㟬\`?�;����be�^>�Ɉ��3_Ѩu�|�+�u�'  `&��`�v�%�e���ΒV]T~dQ��f}�	�kg��S��|*p�^��t����z�s�E� 66�KƲ��̈�Vm4yf��	�ǰM���v�q�T
E7������=�<9���P:���m^J��rV����)�Hm����Bh�����y���oB��~ ���K�	Ig���s*}�#8���j���~wHd'�>�αr;��qy��?\�HN,̗ᚦ�/�i�}A��������dm����O��p;��F��@i�
���6��m�gr��t�2q�z�]jq��4+;���ң5��eP�������h�>i]���R��#N�x�F��C�i ��������2�T�)�5�-D�l$/���[��h1i:{+-��P�ӯ6��Z[ˬ��7��� ����&1�k�'ׁyU8�	�Q�4ʚ1�˽�3�y��i�'��s�O7��;���2D\�6���&?���B�R/��O9��h)s5�Y��P�_{q-h+��d6,Kf=mՒ�;�q���J ���>�;��u�ے�O�✇�b_�&��9 e
fQ8�:��F��%�O�0�?����m�/�h�e��f>�Q/n!��TY|ޑ�Fz��~�ظg�G�g�ڊ�����tE��q�����
��)�2�|�e�pC�����21�����
�1�Ds~��tL���8 �=P�$����H��?�
$2��]�#��A!�a�Ǆ��&�z,w} �h��NG��}ו<�`,*X���1��-S�U��� DV	�5$f��<E`��UA	���W₅��2~��Oy�5��XųsUN�xg�U�1���,��W�ˢ}�35h����@[��i|(����HD[4�WŔ�B��/�@Q�;��Ynhp6`���:����.��-ͭ0?HH�m�CS]1Ex]�$E�9��q�d"���jԹm-��m`�s#+%a�2@�����ؗ�	}k�Z��\g���6�w���9)�*��B)�0n+M� ?m�/�AF&��5H�?B�z(��X��皥Z�o�foB�XCiHҧ��t�oUA1�/���S�"�Ty�b�݅�Fߒ[e��r(���~|�.�`��8��ͬ�\��܎�탖���^�w��M��xl��8�� �q8H3� ��2X��/#�Ƅ][�w���~/����������U����V�=q���j�R*�՗V�F�2rʕ�����؞Q�x��y�����H$U\�=*NoEJ��IO���B�S1�2�S�1S$%|M�:��y�x��c��7��XUx���9ol6�dCM5��=���A�k�EN6��@I�\5�t������ ����� o�',P�9z��������Ǌ�,�C:`h�\k+���yᕱ�B����m������6��_#poU�ajF)��.��E�Q���#�YL�{�AI�����&J�K�2�{ �Mln��<�X0��HP^��L̵8WB&T���~K��j+e�o���Kz��k��x��w��֬jaM3���c0��|�_��҄����q��v�0�����x�S������'�~�FL2�(T�0����4��2/�����v���~G��0��� ��=����o��� ��VL�e�8����%m��,Zb�$�4�y{ġ��s%��]@�¤v@�Z�M�|�*��T�pӽ;<p�$�Q;��!���-�g(ɺ,o�3;ă����g��qw�G�1y�kOP��R��et�1EA�T��D���k�W�P��4W�����3SNb�F�VHI�}4p�t�]l;y�4����GR��^�P�6��J�%�A�9VoYb��N����ux�Y�4�m�ڃ��Q��<��S�h��xC̭���(RN����T�]1A1�Ґ���
�6g�a�f��d
�֕��uy�qp$�m�$�?u>a^֤
�R�&$X5��oA�'���T�4ATͦ�U��H��i�R|X�'���t}Bc���;���w�A���)����z���N6����@x}��J�N* /ӭN ˿	�b��}{�tV��"��w�(����r�(_��
l���i6�b�d3VA$`�,b.s��͖֐S�d�Y�{qؗ`MG�q. �8�C�mR����Ϛ|$-������P�g��ޯLJ@���a-��r־��ٺ��>X$�8�6;�F*�;k��À�5mBj j�'�K�@�����)�ŵ�:j	�k�\EY]�Ll&��gt#��i�5��@�H��"7�k���<��#c�B�q��f�>�PO��ؕ�/��l��/�):n39���/�]�h�Ʋ����kAi�]�ၴ�d�^ڱզDf<�E���?�Fya��
_`%�e�s@?���3�Dc�IC㙬���w����ڎT�a1O���>�P��Y+:����Q�@��(�t��9Q�/����h�,X#�0�8`��Ls��J.\�7c�)�|��@�T��_;�m�q������3a�=|;�I�gϜX��VP,�j��IX�<&a�9@�"0��!���~�
p@�Y����}K,��
��7`�G��ʠz�<�pT�|�|�BI��G�$�ׯ��M->#�"S��8�/�����"J*}f�7��� P>�_��q8��H�7�仃�@V��vP��m��=)Ή�E�1�򂁤�kw.T���z}]?�W(�,�~Li?{c+r�і��-�yu��v��S�=X�+�����l���Y���X^I� �֕	���\8�#<������T�5 �����{���x{�	�9��d��<+��#w�j���d�Ɗ�)�3y�M��������˪�Q���0�7j9��B*[�M���[�[�k�ޣ�A��|�Pz��5^�L�<�H�+��q�s��>F(�:�&�͐j�S��*��$��7������H���Ӹ�B^G����_�����u��
�T������1�'ȗhu�a�K�V$8!�^Y��������)ȍ��=�>���\/M���'mq`�r�	_�C��u1�9� =mX[�Cr����av��;�����1�d�bH��g �/��G�O參RԴD��1Ou��'uP����}� ��q���[O7�Ҹ?�<�|��4�ϸ+A����ϑB�VB"��Tw�
Uۦ"���i��x%�C��~Ļw����S�C�w�g�ڻ��(�����gz��,����Ų����Y������6)��sF#����O�¿���rtЋ�Ԣ�5�u�
3��o�rܤt* Y��@��y����~��8�]�NC)��:m�%�����&�6�^J���\�̭��ƭ,D{�$aG����z��<ἅ	�Y�<	j�M��N^��纉i��I�n��7�A4f����p�}L|Ͼ�#?P�V�l��ؼ����h� �o ճ�����Zq�|l^)m�	�*v xJ�lJ�������y��[���a��Y����Iܰ���VX9��'d�L�-d�؉h$-�0�-�>6ZnY�"!&�y�sA��1W�O�|��=ҹK��rf�x�+��B%$b{<ʉ��ٻh�$Ct��c�k�+�=��u��VBX}Ǡ�տ�����zͰ����M������������HkV
 ���Vأ���k?��9���'L�ޮ"��������2(��HdI���^��̯Ĺ�d�Y�f"�$�[�b,4�o�)ʄ4�Qv��c_4��֗�[�:��f�ޫ���y6��=��`�cV]o�y�m9�R�r3��\�I�L���F�`r��V�az�x����P_�~�����8u�����}�9�{IrY�L$��t_����[�w�S��?g���%`�_�lb�=��c��?Ʃuh�#�w�����۲JP%�r˼��L���c:�N<v����(��4�t�2eW�?B��s �F��'W2�R&=|�$bU��Ȳ�"�,:Y�j�?�1��j�ȓ�ǅ���-��3��\�h�J�A5@$*�v�;@�ɷ�r�v�/<=��S�̢qhm5>��|悉Eʗ�`e�jW:���_o�v�c�2-l�ʧ�k�򒩕��8{�xs�>K������&l+q��ǉ� _�|j3���枢��,IЩ��BR��p��\�`o|zx�f�A����v�>>��.(|�����-N/[�����	�,�ƃ ��b�c�p/Z�����n�}�k���b��i`�Şk��*�=����q/(}�PXd��[g'gS�q������� ĝ��>����Zˀ��(x���O���㴲�A�٪���p�8���w2��&�jm��ՖQR�������sèݨ���[�c���ڳI��������	����Q2CT��HS���KV�sM�9-�V�x&W��f����^0�Y#c��8��p���>+KPX*tQ|�]>*�
V�ޒ��-x�K㏣n�H�˹�|DI��h3�6O�h��	2�gpH���ANǷ1z�Q�g�����s�5��biE��H������ө�~��:=�l5�ׂY(�Ǔ�u�\:������ťp!U]1�C�_ކ���l�\]�`Q!�d���~�Fe$:vO��̃�V������hpx��츷�@�l	�Yz Ӹ�d���5گ}��~���+����>_�eW�e=��
[����߽jR�Ҝdm�g{y�a�)	�(g&���mjS����N�z��7:�q���f���X<��\qw<�rX�0�EsNT����;�X�z�av���hJ�Afɀ�py����Nޏ A���WΔu���RA��P�R��%|����(���m�����)�nkR��v���ב%C�3��H䓳W�5�M-B��'��ʚ���i�����BE��
J�޹�(7ĩ��Gʇ�_0�R�ŨU2��͞P�e�Q���}��
,��]�,s���I���a�p��P3���R�����6E����1�+�T�R��l��v��H�J�ܰD��I�O\r�R]��k�-�H�X~�yP]-�(r�wh�έ�"�l�R�]�ȣ{$����q���H�+��G���;�"�����)WT����/N��44,FX��S��]�(9�M���3��q��v��u~l�6�P��n�-'�Rl�Zi
/�W��_&m[vO����*�̎y�b$��.�s*C���/{k�|�^3sg�'�
E�ƽ7��'T��I�.��X�����K�Ku�c��:�z.Ei\�uk�1M���za�D1�!��c���"76v�ﶦ�5�r�z2s��[��*���mh��{��i��>�[���YEb��и�]���/|��я���]�Y�E������/,8�9����^gI.�F�Z�.�nՇ=-\�'C(C��yp������8��]ٝ��0E_{ه�T�T��_�0�o�ld�a�ų
��{<�N7j��wa��b7��'�����9�V����6_�؝���p��v�;a���i�E�� �9�Eu 9��7 "���>��|^I� :��R��tI;$<�$B���w�_�ȩ5�
����N3�~^���nA�����g~"��O�s�zV)�,Dz%��2�'��ݓ���LQ뺫\{��S]AtQVv�s�F1�b6�-/��os�� �th:�����~c�������ݘْU`������m���'*=��h� ��*0�}���~�N��l*m���Z��R��1^,�i�9�������b��������Ŋ�^�s�;�;n9�'�{p�	�9\x��#��1�'>2���SE�)J�~\����׈u�C=�Ǳ��,� �#{peZ�OY�%�J��p�xЇ��MS������h.�1�Sd�z�K�G&��h1S\�Qq�p��
�N�~bi��ݳ�j�@|D�ޭ���G2�e@\���_�kQ�z��q��P�ܑ&��495�;n�4_�C�6:��i?=�lV���$�B�=��qP'����
��]� I��I�VtI�N���$.�M
��8����!.a�D�B��텁rS�d�򤤮�2�Z�?S�L. �b���Ko� [](��y��W5�u�+N� ���%�2w�ʠGi�sC���.���V�v�rcا�:%`����Ja�ɻ'���/DNM��ozGnc�Oc��s
ed�>;���*�:���r�=$Ad�P��RU�n�[��P}�!C~K�Q�Q����>|�d\	�:v����6��O��x���;bd�K���<��cn��`�q�y.ss�q�i.��� �}ri:��O�<AyB�� �
�` ?�B�TS����T��2�0�ʼ�ܵL������ u�f��n���_:[��ZZC�g%!j'I5����D2�J��SZaŦk�'��9t�*�H����e����l��S2�y����W�r׆W�I��@�,Z=��AF��+��	�� �����s����pD͖nls�4Nϲ�(��3*�r�\k$��v��B�0����y�\_>N�o�朕2؎j��.��AV��s��YA��ĠY�8{	�Qek��h���T����D�ϣ!K����tYXD�x����#�Gs���hʓ��%�Y<kN�����v�9�b��76�&f|�b9�<�qc �J�q�zf!��j>�c��=��4ބ�=��m�����0���6sEy�	j���i!�4����:�JF���^�0e�d��:8γVE�Jث\�ؐ��k�B���c�_���4�#-,C����ܸ����Cc����7]�-zCC����!�B{�˯�~R[����-49�� ���׫A~#'�`�֗��G�΀��P<�5���ȪzK`���ub����T+N	pd�Bi�JM�����A�}a�T@�Ή�z���7����ב�IlQ��oiR�#�������L����!��tO�v0�n;Yn 6:�h�N���ei��$��Λ�.��ǃ��<Z��3�쏛D�z�;X��ˢX��h�"$�������䣶ͨwѨ����,R��g�z�<�hX7�����^�MB�yl�G�rK�m0:$	��\�d�����Q�`�Q���sK�3Wy�k�-���;��\����� �kLt�e;�Y�%�E��̣�;5)����pM�$}�dkCK!~.�"<�w��w�6�F���y�2�E[5�H3� ��<�WQ�_x�t��T:�d�V���Rb��M���,��#�����c,M��ڸ�E	�Zk�!�t5�~<�qۢ(�9��vj/�K��e/$��x�[u!�&� C����ͼ��^zFK�^�����,9�T���3S����H���ܬL�@T7jY)/�p\]�s� �����Y����튩I�#�>����0~ԉ/��S	��u~�;]�q�D��}+ώ�h�0�]��%;���7��x�o;�\>�`X�U/��~՟�GpV���-H����1�|j=�oG����\Ɂ��ӯ9�F׀,I���2��I^�lR�M���3�KQCw;E�������P��#.�fB*����'O���B������QT��������k��������^1��n?�V/Kג:�j������0[�9������J��z��$��+�'ш3�8��~���B����n�Y��� �.�?�J�m̀�u���?��P+���)���ܡA�����c�U�z(� ��(O�ȶ��:;�Y,�mw�jĀ�P}�)�b�f�_SO�lG��-f�>�K�{w�!�6�F��/��j���:���|R�58��@���£9�r�̾Ɍ�r�� �}�ɕ$��`Re�\�!���m��T�:�B�C3��,k�Nl��Y&k���u䲳���v��ng5� ��$	����0��k�����x�d��)U�T�m1EH�K5"50�ܑ�o<A�9XX�O�b�(���T��}r��P������2,h�KpS��4g�gs��A��M�,��6-��s�] n�\
CR'Z���Gn�d�C�Xw��,R�񝖆���0S�A�<�v
'ȒNiŷ2��ȏ[9cC�Kz��N?X��W�!�����E2�Ҡ�Yz7q�<�`bWE|�|5p~���ό����⚔Nh� @&��I��/��V�!��+��l/�¯7lT�$�0�mi��z���6S�zb�+�]�wR�-SH��2� �kq����տFp���j�����<�=M��b�Y(N��(@�Y��[��	&hq�"d��
`��|2���@�aR�6�/����q�"4����N�����͓Z�TG��'0r%"46�
�1kl�	��O��?����a��qF
�y\ߙ���k�6@��E�j1쟝?��H^Z���\�O7�uѵ{8��%#ͧ�`,F�[��o&�p|yZ:��{RiS-���~�[�* v�V��t��恱Q.���	�ǐU�H�[�l0��\4���cy; �&�H_Q�j�[Zm�YY��Aȅ����K'q�3_c�2���L��]
��9��kڳ������Q^��6ۓo��C�9�N,?7f�ځ.��?	1�(
�p�<l�t�-���QG<���ڟ'�&"�!j����9�"A�8W�Dt.�G�	�.5�Ne�}� )t���$�d*�e�le�w�*y�pk�ma�ѱP����_{5O}�65Z	�z��/�'@j�����<w�У���� ���Oѽ�&�x�|�d��d���SΎ���K�w˴;K����E�-xs��`üƼ�!�P�-y'{�,��p��9����;�x���@@V:ND�E�3,��Ug3�A���>�^:�X�s�5Zsq �'�!Ƙy}����כּ�&n����u|lEo�_Z7i�+�1�j���)��p�ke�B�^�����\�kw3?��504��6���G���2ړ�[A��H�5��ù���c涠����|{�X5��=LO`�3+��P+S����|e��X�A�?h�GM~����$R��o--�{eƂh"��#\�Z4����s�F`a�H}�,�����!�l`�FyX����qڕ�+;�^���'N�����ʞ�s�MU��q)9%2|����� ����$=C��9���\pnϕe�%q6 �.�ν&8ɧ��\MRFEu�獚�%��n�|���`�,6�p 3t��?���K�S�ߜ��H��˼������C���6������J�
A�M��(�n�N�Y
s�<���Ǝߋ��o�K�9��,�EW_�a�:�hW|{��^A�����Rza���ߏ��F<�nb�R�����Z"0���SA����-���6k/
F\�b(��'
�Q�s`��9!ʘR����\8f��4$�y���Ƹ����.T_���dܥ7s�9��b�V]H#��M	������8�y���34���P��">�3y��a�zQ-�}�D���ܩ�C1+�jg��
��l;=tivz��fg��YT�U]br���qw�!�	F`��W9!��>Jڃ ��1���Qo�rq�S.����S^�����Ík ���[%�L�q�0h�uU.��ԣ&8��Y*�f�X�x�ࣲ ��{Ξ��H֧�7ɑ����'͠�T�������v�b�d`�<r��a
��t���%����u�6K�s*�����M�)]���Ac|��6+���.a�����=��|%0���VJ��<�gS�<X8�ɰ 	�veH�Z�I��+h�.�UJjv����:�'��^�ݒ�:U�0�e{��������t�|��-���_d�Ebg�TP)m�9@[`���w\�&,m���ђ��x�L�D���p��o4g�HVH8Oy����,��?��q�D�7}u?ݣ�>� l��ӡ�P A`3FHfQ�q�c�C�x?���ŕm��-ߌ��#��j&i���:���1��c� s��y���/i��n���ֲ6�C�~X�)dP;���9Ξo��?��o��m"��9ۘ���G΀����P�8S��R�WDY���ql �g��!�F!��P�#G����?����:��źu]�4�G��TK�>MqGj�}��3��9��G��l��uǡ��pd-O<���ހ�h���o���:9���\�.���cs��l�$/����N[ՄtmD��U���َ��M��s��VnJ	�Զ��2�6��.v�V'�VY1u�r�<2�c���G�AXC�LG����g��b�fZ���-�.BX����,�4�9���A�
�q7���5��$�;1gm��f����]L$L�!���W��\�0�E��(���·��KU]i�=G�hy�p��D�������J�Ǐ]�D�a�YFW"w��A�{�����nRCL| h~	/뚙��/˃�Տ@�:&da�CP9_�9��6��5�*Ck�O\�-#GNkt�C���V�q���sC5���EHbZ�$�9����
���0�
���}��~/*,�\*�I����׸u�A��/_!���7Z���~py���_"|3\����Oݏz3����F􄳤-@)mα�cC6&
�"}:�cd�,0�I�3.V��T�a�g���a����fTz��b�q�B��5Q˧gU`n���f˒�!���S<����o�����.ԛsa�p��\�{��[6n��B���e��)�}�Y4t!���j�*�k6��><�`�`WNm�;��1o
�{�1B/��PX,t�<�����6�1hk�G�`��/����-�j-�z�����5>b����m�E"��e���b`�ZU"Uls�1~Z{X�=���fI6�'¤���ӏr���.1��vF�L����4�논/.��}�] ���h�kCW����C�&�ܙ��l���n����|�SrԲ��/@*��XД8_B���GcW�{�V���ړ$�} 8ccEV.��:=���Z�FHr X@�<vBrU���:v�A�(�/ �+�7v�CV#/�5A|�Z��ɦ�nx��'W���$�\T���A'�*���~�tG�IyYe�.<���}�;1z<�������@�tz� �b��V�!�Z�26낛Nn��������Nˆ	A���Ǭ���K���Lc2�0��:�$>�2�ptBۑ9�L��RI�<��)|�������eV�}3��T�:wj[��D��.�b�{clM� �b�c��4�4�R4.aס}����k?dgh]Ia�1넗������iM�o�s��<�۹l��`
��g�)v!ۚG��mƳ,��m���[��hɕP����<U�I�%'�����?H�/��3P*K��WG���7�wi?��᥇Ђ�-�v�s�3vT~����~���SH��S��眢c�T��
s��l���%����l�fcU/�}�GjqaU������V��%�?}��iݦ��یq�nb�Ԫd3�~�\R8�f}fw�?|���fy��),�g{�h5��'��M0�����r�[���{+��� �
S���4���I��EWf�G�H7^��RM�ERm�_�&M:C�c$�$�׉3�}�N'i$h,���Kfn����a�iŧ|թ��,9��zy*�"�h��6r�Pe�
�l���f�W��4���N��?ꓦ�j�f�D�ި��kО�x�0��@1ra�/I�uy?Ǘ�o7����cX����!��@��c-�q0w��s���x��Y�:��s^*�2!���@X��$6�����2G�n���(W�l�/Z�#�H�1�8�ݸ˖��l���k���� 1���8[&�Z��gg��8��C�Y Ɲ0��������z�1��ch�Δm�*���2��"GГ'��[�������\�͇s����J�䧨o��k{S�q���|U��}���Vkae}����]���M�eH�'Px4o��c��s	Q��,��V.���k�1d����H���R�W�?`�G�6��ؽ��-ua���HJ�+�Y��U 1`���*�v���k�r"�0��M�f̢u���r�!x�l��=
���a��)�>�I��6�:�\"�j���j��F�a ݃�4���Z�R���}wE E�h-n��\q6�b�ݯAȷ�G�jOV�K�!�]5���Tf��XI�Z+~ja��������������~�'Ez���6��b��;qaQe\�?'�����-�������?FP]G΋�t�f�d��&Ŋ�!S,�F��ܐ�ؠ	�ĉ�L�x�c���@�c�v)<S� ��r�+��`�p��-��E��*CU���^{D�*�o��JwN�����JɆ�2��{�O�_��u���*�>�D�i�X��SSD�S�stE�z�gA�$G�e'�5[�h ڹ<��`��eR���@<�X�"H}���)�V<�5Z�G4���{�ak�WQz��Q%1^cA �t�A��S{�SA`�KM��BBVs?�`	&�
�������kxS3"��^�^��f,���M*��~�~�({SNu�f��f�$�����V������E�Jl�oj�S�[g�����=����N(ͬXh���8���F_�?���(�.����iv,<�hQ���&8JN���pC�8�˄�p�=�E���"X��q��:��O�=�~yFVRu��$�x�s�|4��\l�'�K[�;��T��I����_����	Op<����#V�$���m#���!�S��V�/]x�A�F�����ʍj�7��)�p��2���\YRZW�9�b�\-�dd���2�$zMi����r�� �>�D�����PD)���z��a�:�a~�bM�a胘�˴.��L��Zs��k*�R�?�GQ@�:��L:�RC3�4��Kk�'��AF0!<k�l��40��Z���Fsv=a�{�Zu�h�e%�9bڈ�V��������D��"��G 5��ux'���FM���m ����솠����tr�Xcc?4'��:�a�=s����jB�,odF)1(�Þ(HN��ٚ��18h�X5���K�6�Q�i�����)�!.�	,(*�<�R¦�m�d@eҙ�:�v�B��#=�lI �i�g8�;W��J�6r��_��4d2�('�t����<!o���ѭv�@gN����\����Dv<;~@��d�~|ʟo	��Yo�T���q��u�`� ?$�0�X�44�ty_��/����{��E��Vm�s'�F/做�bl��J5�s�͠v�Vy���w��_i�	� '�5nugP~�� ���ŵ��� $66q=�4آ
���H��� �
��%f^����Ü6�&E��
 /,��=�<C_�N)�RE����I�j�aF��6n�j�&���o�)��tz�2Qw�sP����e�Nt����+I���فך�����K!������s��������d-�y��<��~�z����v�T`���&:��J����8РE��S��1�t}�ڠ!�����ށ�Q��3K��"=:}n$��w�ځ���.��u���)^qk��Y�bfg�+�&Ė�+74��N�����,E,��g�3�����&td &i�+�*TF����[�#l� ��8�
� ���-��	�D���PpR��^�Aʱn�S��%z�r���	�~��z/��w����~tT�5I��Ws�'��� �7�U&�=����HO�f����&Zg��CE��*��e��[�:�i^�0u��}�q_��
(Uz������LS��洌�l��r �1M�������l�g�"mo��O�hګ\���AJ�����i��2C9�����	��^�����mޟ�L� ���<�#�%��`&e���6|-PS���ǢnjF��
D�SFɏz�����k��l�������)�z�O1HD`S�H������w�?%��m�M4=g��"�S�^$nQ���@�9�AH�a}Arŕ4��w�d�����M��~	�e�ӟ�D(c��^�n���
9c�âw�x�F0�/�h�����|�Mj����O��=|:$�+I%%*�#��8ǘ{��}���P���|��8olm���`8cQ�)-�(�dY_����B�M�@��q���#'��(V��1_��OZ{����eE�x�#nq����s�o@�3M���RC��L}�p�Fp�UP���Z c��5|J���,�k= ��i��Bqz�s�鵴.A��NGތ�11��u��s�> :������!�
����J�t�E��q
NB2r�,<9����L@��f&I�jAa��kSQ���Y�^m&�SY37<T���a.�"=.�h睢�����B�����H�\��G-�@dE��.�.o�`Î���5���m�3}KY�ؠT|�p�����z��?U��@��	������Pp�#��Hzci�
�T�p�����͝4{���NY��>�� N#���	��#�C �U�%Ʋ:ϳ����c�T�ڳ:�bxG�Z������Ənd��Y��=o{�2K�<E_%fL��� Ẍ�8w�ye˃�> ����]R �\��������G':��ǳ:#���f�Z	)-��Y��u�)�[��T��i��
��">7>�k�n����HA8���x�Ii��f��Q���UE!Οr����_�w�	0Վ��2嵓Ds�e������z��l�(i22��&��;7�)���k��rD:�<�Kd�t��=ρ",1���(&�眒����T-�j"�����>ݽ�"?v�� �Y=6�m˂���|g��.o�����ì�$����������h� 8�:��u0�׌�9���V�R�!��rC:�HmK�';���yɔV�e���ˠ�|w��|�a��)�������cV�J�pفPl¡�
|��8�~��W���m9�-�;��K��c�\+~// �IB��R-_��}�i�0@�����jIHP�dX�]�)&�$�����l4��l-�+���d(Uªl�@�:���"��э��OQ�VY�5XJ {�UH
矆)T3�����5>�� �%
+N��y��y�JE�_f
z^p=�1H��K��-���ґ��LŸ�;����������"�*�4:,�s�@���xڨ��	��7�u�EUx{f'D�����=x��C�P�� _��0�&�gf��bg�q_+>k�%���඙� ��Ӕ�L��#�3p~��+���^1@�� ��p��Of�����Q&�Da�ʫb-f&�òF˃	欆�j��
�p��2�3�Q����
�/�5���r^��ltϰ9�qԾwޱ��</W���@����?��b��U����ƻ_���Px4�H�k7���Ix$؍�#�];E��q"�jBIi�c�h��Mpa��M�����#<�
E�7�r~[��	ň�=�s�_�����4"�o"mjr��ܷ}F6p��մ���YzV_��j��v���p�B�G�<*XȾ��Y�ywrْ�5��Z���m;����X�Բj���g羆�}�7�N�M���[;9�cњ����v�g�l��8m��jn!M.���s��gdדxav�|���8mn��Y�{^�T��W`-1^%����]�p�z���- V,�C��aݖ����#5��E !e��d�gHW"���=rC��\��l�X��}4�.ĨSd*���(������U�w��xz@se�<�������V��ׯ��Ҵ�mW��ή&�m�+�(K� ~�Vz�W����bP�9_E�3b<�]�ә_x�W�/��{R#�J2�bHPGυ
�fp�?:?Չ�r�j��9�2-9����I~�=A�-c޾�	�S��y0��g>��r��UR��`CĹ�у���g��(JmiP�f��!�8)�D��J�'7H�����]�Y��3)��?*֦�P�z�DM\�h����������4�|b;CW�{Ġ��BC����ƪN$ۃ�5��j��ެ��"�y�U@�����Z�~��Z�Y����]�����J�L���]�)䉧?����>|�\��� �O���p}�Z��?9��d�]����D��IXd���ݦ��̾�{�;ds�\\OW3���-)���ɚr�/6���҃Pр�gQe���5'����#���Ƴ�Uo,v^(�G9V�f�p��i8Z�Y1W��+`�L�������s�[���_߿��b/���*�pi���VI����2�~/`��zHO��oU^*����\�Z���Ύp�Yv�j��܊Ð�/T��~f��!�^[Vk5O�h�c�ň��E(�+��9�O;�'�u^ٮi��Z��0�Cw�/'�|�L8����H�$�+I�O,㦢|�J$u8%蹮��?���������٥�;�y�2STg�	�Z��7�i��2
Som�Sm%�i-��A 	d�G��٢h?���e�/��öC���������^�|6C"('��l9> �I7�O�h�
d�W⓷����l���,!j��X��3��A�ʋ�=��Mw<O*�̣l3=}hd�<y����Y��r��k��
��Y$j2����~.��_��@���g6����D��q�\�M��\�	b��{��ԡ5d��_��� �|�I1S�j��T#�}�"p�sG��rs:0)����T�@?ġ�ʱ�F���岡B��c�.���᫊� �e�α-�^9���5�9��wOv�Ojk!	��e=�[+�BDBu�g	@�Qߺ�2�iQu���1���ӗ��s��-�$s0e�"fS��ވ�d8��J�6Ma]��S^�����ub�3l/X�`~��* 푳��9߮j.�W�/�[�3E������,�d#��?
��r>�����QoO�"��K2��ɕY��t��mu��K ;A�+�K�ْ��]k�L��-/�^���
� X�?[9�6k�����	&�;�+b*�7��m�v"�~tD�瞈C�a�ߦ�!���A���h���?��"m�^B���3�)��y�=2�z���TE",� �� ���6�4	��hﱱ߈ ߗ�����C�^�-l�,�#O�X�̉�U�"-�;�~��
;鮥�[�`�%��,�S|�ڙ��̍[n?��0!�MQܩ0�	�tͺ��O���ز$��n$n�D�84�+���A�Gd�� #����