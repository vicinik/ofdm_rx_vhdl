��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�e:�G��P1��\�jHiV�PQ ���dh}H�Ɯ���I���v���5:Y��K���� ^ԫ<�Tɓ�kVb�V��2T8�5��}F���}h����˵���t<+5(H�#Sv�#N�O��R���n�d� �K#�_��Ȥ�c�{d`��|���L���Pm&�
"ef)����\�@��gb������P������	z/��JA��Upc\Jx@H9ڳ��+K��1�þ��W�	ί�IY�H�<�>�<�HOhn�T�Q�A���A�<�<����������?��W� �@������p�o�� �O�����F����|��+$�jAͰ�V�ў�67�����_��-ET[Y�t_�^�^@��L2�,��>tsWxf�yB-�f'Y_9�I#��.���
T=�/l}��/�G���)�\�Щ�y��u�#t�t�m/{&5�1 ��jH�5�^pc(4����H����O��9������AY7���s��<hMP��w��L5��](�v
@v��qJ���8\�6�9e��w�E?�1��wَ�}{=��bҐ��*��exM�V�	����E��c0+�K����f����J$�{6c��B��� ?�D����
���Q��T����gT���?Ѳ�V�1�6�g|�^����K&������ǃ�yޟ���q��+[ݰ`))_:�,y!�אIE`�7���Dr�{A���ٿ����nG3����q�������� ���8�P�e�g���nZ�N�M�9y�er�!:�����Đ��|�x�e�&Z(�`��ۗ����!�K?S��Q�Z�M���J}ckk �(�;�:6?�4��:${f����	�#s|	���k	�.Zz���gX�J;n�g^t��xq�E�l;��p�sh�Q�4F�g�V��j<���qlA����&���0��m<;��\T���K;�%�O@ʓ�B`2/��N#���w+��w��a�R���q/�c� �έex,��j��v�Y��<>�|�8@U���D�$�᳍�P���!_��|~�2u^枽����:´$&6.�y��f��O��CD
*N֊ ثR�j�.q�M5FP~4>߮��JN���j� w��VD5��K�A8���@r���Q��X��k�<�!-aw?!��[A����-��(�����I`j� ޱ���E�@qc2"���ŷN[Y	GI����E���8N�de��͹�$<�iDeu��&���bm�Ņ՚�67�h@��"B��3����[�����FD�A�A3?W�1J�n"J���{�-	����	([r���|��0��c���u�`A)�4󴑃	��o��N�������2��+/�cpnX���#���&-A�� �e�M�j�$ ��cO~n�:ip��[J�q�3wW�""kÂ&�=�g�U�`r���x�x�"��_Q�.��Sb�p�ز-��}z�u�͇�zz"�x��I�#�8/_2�u�v�$�9 �\ה�h��'oF�J��������1b)�jq ��ښ��C���CU�l&�z��S����d|`�Y�
7B�@6���ƕ�.G�vFD�T
��j���Y�0S�)j��˾�(��b�m���,��!/�o٤3�=ķ1�D��	���A�82�\�,�-f��H����/!��A����|�K��̲����2�����%.r��	��
��ԵC7�d��3ÒU�0�՛7��V�#/��k��>E�%��y��s�H�Wź������ޛ.� O3���1$�K��K�tr���>T�_� Զ��^8�c�耩	���}���S�LI�G��M��r�����xϹS���_Ų���@
ү"yy��,�q	J�w:���'��#�KS!tw��b�t�J_��}uOP���~6W����v�j��hФd��3-�W��⼻A���t�2 ��#_|�[3&�Y�-�V����p�l��,���=t�A��>�={E��@5n��yg��ۈ��mN0�B���������
����(�X���4Z����e�?z	U3�͓�
�s.l�n��i������w�(�w���2�ʜ��	���W�H��	=�.�{��/���&�߇�dE9�$)[�R>6�ޓ�j΁�ĲEF��G[Hl��P�0�Ƭ��.�
��Tp�\8c��h#X��R���zS�#|�x����ք]n�%?��僂#/�G7U�e�vr��Ѷ"�g;�)�z�ѭ��ll�qM�ͼj�����T���eT������ѿ�ڮꅰI���<Y-�S߸u����k���2�!�cw$�f�5N���k��?~4{�y��N�R���ş��Eu�x�y4O�����|u$.���T|Ye*�9n%�e�;���u]�g�V��~�,�!+�DUi�������6o�m[���J����Ҏ��P��ue�"�BPb%�+v���!1��M��9J_$���Փ�����(�����k�T0�,�`��C�ch]y�ao6�t|�E�k�z�P�j�ƻ��.0gE#+�Qk����|�?wU�$u1�$zF8!BJ��H%���Ԥj�$�;t>[�3�Fx� 4�x��6�R/�ÿi#*������ʻ򇴲{�B}�%�@Z�ӟcaA�!����PƷ&g�*��'`4X��ͷ�c���(��n��[�r�=Śm�j|�E�iী���]o£KO�5���b�Q�ɂ��t�-�Ư��ؼ�q%�W����Bٿ�G���`8�۞�A؄n{&��`*��Oy�J��jjƤ�210	]o+��*���o6õ���(�&�|��RF��XC$QC3R]�	�(2H�K^�m�����D}h�џb�V�Q���ޜH/��2�c�Z�Y��)�wT�^B�*�έu���C�J�B=� '�{<�D�k��V�_��Te}P>�غu@�T�MK�ռ�毽}����S
;@;=H?XVD7>pX3��(u����KA\J�-��X/�ā�c�6M6��kd{P�U��u�yaK��P�~�C'���N 
C�o��S���
2��I�1:���yQ�P�ɫ����x
0?c�P�;5�8��t<�}F�//v(�%�V�S�L�?:�O+հ+=��!�vwiΰ��?i���K��Z��d�����
�-�r�X�����Wd?6���m��s�!e9H�>�l��W�X�&h��Q�B(e��[��N^a�|��[սHT������c��l�(�Y�ْ�N��?��ދ�<�QKXXvC�Y��)��xF��{��)���:�ɡ���S�as�&CE��&L9EP�����Wp��n n�+Z;�T1O�ob�SoO�YӐT�!�|$Y ��N�#$�Y#��t^���.V�B����i���V��A\D[5���Ԭr�Y�L{�ق�w	�&o#wM�H~$�z�k�����'T!�����B�+<Ӭ"t�Y	ps�Au2u0Xc)��������7ȏ2ڞ������6�q��,�W-�j���3G��0�g~� ǖ����֐�%���~M��R�� ��%���T�/��b<v���������fa¼�|����A��r\����<�pK|{��4�e��
ǽ\��)�C�8����$����H�:�m<2���:I�$J��a�0���4��5ePd��Lj��|�
�sǐ�W�A���UO�� �7>�Y?�-�����;�=?0T
�}�+2�:	rB��p�3oY��I �z奁���)#�"[O��R��s�/��.x0i����X����1mD}
�l�.��U:���3�I�!���MQ5.%�)�8�� ���&d)+��8]%=���K�HՆ�Mhj��>X?�ɟ�-*~;���U��8��1�S&
��G�z<�$�7��8�����O�C-6��m��ü�͑>4&���*+�G���|֙�@3�f��τ��w�������`�#�L_��/2Tx��c�oi��3�m��RK�Hʷ��=�Zp�o}2�$	#�EpX��A�=�i�m�P��H8��Դ@�83��QK��8o�0��%Ȼ�ǒ�;s�Dm���1@CVI��&8���"Rs/�k!��U58�\߮��"��8��o��Z��H�J��R̦%�mT-���l�!�(8HD42�]�4��I��T/l�Bp�� ����*��49�|q)����g9�R6	�x�� D�̞hJy�ڑ����l��qz#��0�?�X��b�-���^��?K�#-&����i���������#��Z3��5��J:j|�[j�n����������� �Vx\@O������nuw��

�U&f��X��wK��� ���E��"�c�G�
���H�!(z��i�<S���U�*jPukk*xZb���g�^�6�{��T�,�6�s�{��@=v��L����_A�
��o}*��pQ=8W*w<�[�/�_;
+V��?<Oxߒ�:�3�?�ׇ�t���WH�̄�Z\�ߑ�=�2Y�*89����`�����MV�Q��U�$�=��<Շ��L��j��4H��}?haViô/Y�v�J�)��L�잋^��l�*����	l�|�%���|��!�zZ&�)1�`No��aXSX�'��1�V��97i��3�%�ě�ybw�c��Z;s|��~9�À��/#Rߩ
]'��3�t)�gd	>z3���O(��a]N�-�a���u)Z�|}j�o�� �
��)B�%2����mQR�.��%��ʼ����z�e��<����8n����Q����X�k��,-o��{1_���!��%�V7�`}�u�]}]\�y9���t�U���{���]�D�Gn��?���uk�vQ��.K�q�$C��S�&�Fƿ��M3ͬ|ع0�6�V2��:s�6��zT�m,��K`��̿G�B	���~�v�2F�Q3�L�vvyкr��~�_o�Z�k{��j�j����ܪ�lܺ�����Ω��n��Q���ط��O1/w�3�G^ ������+Q�����-��T�����v1$�~�%���OΛWgy�?h�WCQ�!�|����$���$k�(��jô��;�q�ih��I/b�e}	\����۽#�߯�{�?��
�=87��o7��cܑ]>�U�Zv�,v'�)!s�'	��b1��m�֖
�0�-�N���4�=����מMM�6Q=�[b�`��� �<E*�O�×_{鑢\��#t�����*$��5�au�ٓ����O����]���$�h�=����mv������b�ŖMJ+�
WQ�g�+c�.8�$��D�e$=m�]e=k��_�֛���CJ	!QS���n�W�vi��0O-���I�~(
�c�r��V�>�u��_�6�NF�����:�iՑL,aU���ڇW��ZG|�SKγFz�RV����ł.�;�M0���k9Fݴ� ����n�ܝ���hf�������w85Z%�@h��<��"&�A�IW ]�8���חN5On3sE�>�����X���V��Y7��V9۾�k���Όhq�&\	�D�����y����{�3(C�6�e�!!W�R]&�T��
��s	5�p�J`[O��˃/&,�<bM�����Վ�^�-���%��$���!MZ�
��yS&J��=�һj�|z�pkW���} ���t����:�x�;l��n�PO��+�{F͵�eae�nڃ��&�Tm��s������&nUD51��)���SsҞ���jF�xI��+��/���U��L�����N-��������r��{ �)D�p�kݠY�������`�����ΪlI7|�߰�Ti���$��!�sI�I ]��^ķ�EZh~)�r��
�r�$p���QM��5���T�lm�xU���E5�tx�N���~^�ͫ�P�y�q�\c0�H�&��G������=����YZ@�v���#b�Xݖs�xg>��΃�i�Z����gP>��͜0�@�O�3�3:��x��,+���.H���+b���C��V+\ܤ�ݥ�%UޚM��8��&A�9N�;�{��[����^�h7��޻�M.���F>�0 ��U���VP��w�����S����Ht!�V�W�H3�����h@$�����oe�Վ��e�b�}�aP=n�u睭=�M	�1�ؒ�a:��n���sm�ɸ��KN��$��c4r��hb��<������)�ڑhֻ�fL8��:9�},������7�V�V�&&��]b��Dc�`T(-~��/�L�ł�G7�*ڤ��T����R��� _�!t��~/z{K,��utvb6%������n^�\FR��U#8���a��G�c}�(ߓ�+;#����$�����X�TK�t���=R_����H�E]`l��OT� pD�|�C��y�80���w��r�
r:wM�.m��-�K�*8+LL��@�H��4��<_\������������S�E��EE)f2��SLA��g�Fw�)S:(.�`�l�(��v[��y�E��vDN��e���TP����D@x���4w�Hb�]���Z~�V���A�`{����:�E ������ʹ�?����O">�~>`Kyg��q�j���z�,8q��s9����%�!��&���Q]���a=���Ҷ%��Ǔ5!/�?n3K�<3�#���G)_��o!E�TNŐAa-��C@������b�N�� �vA�ط���5&%��%�z��|�G��z$~&�M�� �EeMq���)W�47�F(6�+�(+ӵ�o:�mtm�A/9.vU$ ������N����[��ޜ���5��Q��$�()��1�o�2P���޵b��r�Rқ�.��_�N2����,UQ8빗�
gD$��ϒ�(R5�˂��  ��5�t���M��#��K��N3���+�m:��Mq��A0��߷tBsd*�];�R D�͑��x�X�B[S-���|;�q�D���1�[�ѳ�vW"�Q]ї��y����~X���%-��=� �Nݿ�
A-<�4�>1���gT�����������.�D�ܰ��-�IbJ��Ƭ󅸆@e���eQ��9h�JnM����};�l(�r3��� �܁oAqi���Qg�N��&L��O�@[��F]� Ϳ�&7zWyl�}�����x�FS� !u�w)γ�@h�&SjS=�7�K>2�����a��ډ����x�������L�cD����٭�q�������NiZ�K���~o|o�j��`�S���R��f(%��4O��B�'�%S�K��t���=���P޺0�B5����|�
¾��i�ݳ85h�Z��c���y}ݳ���|��;ov=˽�b�*�X�_ra-��a�	(k��p�o���H���4��ѻ�$���N=tȂ�n1�h|��Cǣ
͕��tkf;���̎�o���2Rg���!.��?����E�M�ɽ� :��gp$:ו�k�@��u��G���#j��ҕܙ���;���K��/��H����>�ZrM��h ��h�����v�V�k�r��B;��h��_2�!t
�v/�P���}p2�?�P)��;�1>ـ�B]��V@EU�Ϡ�x-37��������1E�ʍ�8J�H�k�#�98�]�_�u/�[=p\�t����u��^6%
'3}�p�� z�6H�=�= @c�q5�U]��Q��b�4��L/W������m�p�ge�kT�uԙ^>Lȋ� ��D�����>A�=J�7/M����N�~�2h݁����{��H���I���S*Mg(�n��M����Z�U���y9Q��F+�8|v��&�®ʉ�}:��%G�+���Z��_����T�����U�������0}�F�C-Z�7CN���j����0C��9����Q���ಈ�UB��W�p��$`�W_(�˻�Ґ�@��pmݦ��-h��%�Zm#
?�9�3cz�t�S��N�G��ʝ�-Yd7�?�- X�b���,��B�'�af#>��i�!����Y�s
�kj
g#�����_˺[�͒V���q��i<��m����4&�.��k�q��ف�~>�[錎��� �廣I�F��0��&��yS�W��8�bor�{(?ֶM_g�����h�Bf��+0��Z��N�'��L�G���fjz��[�
����eX��5c�J���Li�.+�K�`X]i�s��� l�������Dr�n�%�8,�%���oH29���w�N���Y1�?%�O�_q���`�B��p��(����AV6N�mKiُZ2Š':����= �`
Xۖ`�ӏ���c�װ�lgPWl'92�8h�z��)���,�,3 ��?`ʮoHR�{���T�~'��������Ų���9���6TN��]��	?#�k���JH�r�
!�=�AN���i�qP<f��}��/�,i�� [H��p���Z2�*fԳa}8���:�.GA�qZpp_���4~{z;Ѫ�țgʐ0?g�� ���.��6��y�!�����m3ca%������H[�<��eu���ꜯ�!���v��?�����$?u�ם>J�л8Y�41| _j�� ^s� ��Ml7�����jpc&YܳkZ^g��<�l�Ҁ�%!��E	�}�O�%0p�+�T7�]�T�M+<D��y��8�p�Y�׏[�DE����/{%�#��!_Ȣ>��֭hųP����N�3�bE�L�����zZ�'�P����N�p�r�b��!�{R�7�]쩪����/���!޶�9ފ1�
SF���*�I_�P/̹��l�y����^���� [T��2[�_	�����(�a��΋ܰ_њ�q�a��8}�����UϠL�%�I];��_�}����Ś����D>��?��C|�ʆ�@u��CE��<$E];�X���1�!<��5�A���"���ō`�����6q�$2� �������?�(~2T� �5�mghxO�hR.E���K.�wI>�A>�`�6I� )8 ģՅR��|ܽ&��*f����ަ%Z��
�d�\ϡU>wuQ�U(kӼ�sW��4�E6/4a��l�W�G�3�+M��CGY��<은ۤ�Y�M��O���W��61H}���ǻ�E�6���c1<��29t[$���w�<�yT���s3��yBׇ���<?��5Ҵ�N7u�,O;(��b�r႔�x��h�ӓ!�q^���F�Jb���'�8����8P�7�N'���V5���3w[Pjq�|��퓹���w���F2
2�.�ƕN@blH���C 4���h�B�M'��e��Y���'�\���S�K��A�n+V�o�-����b'�"����J}������	ܲ'�e�]�r�d��A
�P�U������>�S�n;�U�}��G}������h��*l�a
=���`tҚjj����8�{}��Io�ό�Ί-���*3kG��z�!O!_R����1��0x�M����n!��ҧ��5�6f��,�A��]�Yk]�˿��|���s�`g���j��d'��p'.#��x�#��R�g�l$�+��_�%.�?������)�5�N�uT�ҝ���ŔO��3����_������ĕ����o;�7`1p%�ܫ1��{qo;Ѻ�=D?Lo�b?�8e<���xʽr�h���V��^�?�ET���$vp����:������_c�e^>=��XO^�m�����L��n����v��b|�/�]	�p���1-���<�ڐvtU��������Eg�?�8q��W�j�.�-�������|4E�l%[��D��h��42�24g�t*�sRb`OR_��AP�!�z�KE����o�^X;�79_v��
�[�2.�\��q^�ʼN��Eɬ;d����A��m�cwo��횮����JP"�aFYJ$t��v�ô̴Y2��H���qi�����e���42��n�i�����f�&�#nߠ�n���֫l��C.Kr�rK���6�dpޏCy�]��C��r �,����J��CUS�F��R������se���B|b��>�Y������R���n������%
��4�iz�x��k��GV�qA(�)XX��O�Wl����4��W0�"T#vx��J$�u�����V<�L1ďE�g�����W��� ���"%�Ɵ�6��g���fJ�w)vleB��ď�9���Ľ2>��|>�w��7�$��.�#��6�v=�$R��[q3m6TCu=��t2����VJ��!�^������.K�a�/fH����;7��� ��*g<���C��
��P�]�Ɓ#��"g}��f�C�_+��1��@�d羅�w=�Jm�"���艹bli�H��2O�J��r.�s"�O�+���onI_6�����R��=t� ��a�c�t���"�
Ed���@�ꊹޯ��gSN�.D!_��S��W��vL5 �>	5k�ɹM������	~�ƤW������C�~EI�Z@QKtdjQ:@ac� ��09�A�~ ���,�C�7���i��:o�ED��`�.����cB��CO��:*�%�2�9@���+�*�C��( ;>�p�f�&jq�~,ự=t��dKh�͏=ĭ/�~/E�t/hc>L׭}DB�(�(�64���b�Z�
.�#�e�XZ��t�6��8��K�^�.#�����lɅ���2�����Z�L�\|0���<�E��?m�r@ZTZ�Y
D��%%�WlXsiLv�U�d�[Sm�h����2���B���N�B7�Y�Fi��3j�V_S�n
F"��ZD2%Sati0F�N�Hs�j1���r���D��ۿw���!#�M׉��r��-�Ny��B�7�}0���{�\p���O�]��`�eaXH��{pzSU?�q�` A`m~�ԧ�[���=S-��@�/6)c�p�4���&��@ ���`�x/2Cտ ���&�?1:�L�X�P����R���2�yE騬6�K�R������MJ3c[����(�)	���V���:l�3C@@xCjֲs�n�c��'�?E��E�n���|� �F%l�#�3�O籬�82��3DZKi�m�V������nB�r����*��\M�A���,`�*"�o k�ֲ>j��o���O
���$lClg_��p/?v��Qǻ�GU��8v�.�m��ZM��D�|�v�0����������[��S���0��rA�4����ݤ����]<�"ź���߹��ȉ�+<����:�u~v�<��o.�Kk�p��O�dZ'�ϥ��ʎ���v-�3�`�z�ʕ3�/�MZ>2�a�.N3�p�}�b�}w��Aw�����nC}��9b5p��E��R �e�SA���Fz(l��`�3�К���9[����5[$�I������N���_4���.FR"��4�I����!}l�E��w�X�9�.OD=���F���{R�щ}�j�i�j�yw��ל\(>�|wZ�BvY���Wl�&u>/��1��ir�l��)o34;h7�:�Р�_�h��V7x9"�}��}��$V�Q��Mi���t��a�2 /�e��S0䗽�#�ܲ�H����4�q�~i�(5mǇG�b*i|����w�@���bE�ǜ��7s���A��?&w��	6+�)���D&�L��+T��	�c8�m���(�8ɂ��M$G��`O�������#����<ݼ�E���@a��دY�4��Xa��6U5��x'���Uҙ�kC�N�����=�3���H|�4���Y��Z�սc��M<�������6�����&r^�ˇ�M�~�p�
��ƙ,��!���i��<tԗX;*����Y��p.��éO��N�h�4j��X�98�#�鮼(o� �^�vv�j��s^��)��J���Y�eZ����-�;t���WH���@���[�'p���#~{�ڤ3�}�P4�q�2�T
5�\�ɯe�JT�<WC63*k���L�!A��IBޏ��A����w��}��L�c�Y1�`�@��G�;F�I�y��}u��ˋp3�`��/!�ͧ�áGp[f�ͼ�ѧ��j��-fs�g���h�b�%�ʞ�F��3d�G���('�Y�b�]��yB}MOw�P[rM6����a�A9;�8M��z�d7i�Tͧ�GfB�\=�oi/���"Z�0<�f"F/t��`~���f{�q+�{��]S>o��yd��E}H<������UM�!��Ĵq�*,G�LBp��W~#Fi:o=�����S��']Ƣ��H�5����f7)�X+��-�~���N��w��w�}��z���ci,Rk�cQ�rr4�F�h�=�;P+��*�5u`� �^�C����t����@q����ˢ��V����W���>_��Y�A"_���3Q`�g�=��GK3Twϗ�z�ݳq�&���e�t��	�?w����4�~F��k6�F��D��-}���H,ύ,��*o2�����%��?l��G�}�o0�0�䆕<&�&+��e+�w������̆HU��Ê��꫹����=��O�6� 5ʀ�4
1c9ڇy�k�$�0Fh�E^+<�^{��ܨ��f�7�c��0�5r����O�\�г�!�sL�(6�Ƈ��>0 $�.��8<�KH�|�2E��Ӂ�/��F˔H]ཉ�O�l�E�b������Q��ACR)?��fJ\!��&��D��h����΁���a��8"u�O�di$��_=v�x���<�'�w�#��B���_�z���u�Χ�~*���Z sf�1��p�S	����0\V�@A�(@r�LãeMiZ�s����?7��ު��k���Ά*���e(��	'ΫZGyҹrs�Y&<��x�\:�D���-�<r��ؘG�R)txN֢����\�-��B[�V�u%wU�h,��I���-��u���}V_�O�M%m��)��a�?_Y�3�J�h�遥��9�����P���u����_8t���OIU�!��Zr��	��Eb�bӴ��e��sU^K(�>E��Q���x��Kϴ����r[V�{jh���B��K�����&M9Z�u�e1nZ�Y$��2�6���ߢ�ĕw��g9���r�K�e9�x�O+H���1˷�a��h����!�$���ʅ�_��жB#r������������X�2��j�9�?s�%�4�:��kQ��+�U��nĦ)��N��-)].l,7҅��w6P���΄j$0D�[jlam�&>6��E�'����}��V%�p!%�֤���`j����}�4����<=V�#d��?�=9��2��/oR
��Rw��+ٹA���[�0��2Ύ��Q��(Ņ��a�#�/$�<���@���:{����;�R႕W�d4��3 �C�ݦ��_��+~��=�l� FC��f*ݧK���D�gr���8�wdX@l9'� �_�[ⶫ�3s��F�����ߦ㶘�Lx�&�7Jţ���FŨ?M��i+m �]h-��Oh���$���2�1Ŋ���}ߦ�0@���2�A0�ɽNy�z2�id�������I����y9a����{R�GI�-VC
-9�i�����h�=`�l����/�CFҾ;'�I��j!�xAA�d��=��x���� l]y�l"۰N���Rd@X]zS�d�OG^�sd��?�=���,~�`[�z��c}��������O�L��qN�d�Bu��\�D� 6�
.�ռ{{�"X�[��O�
Y(��4rE#ž����u{���$'Uq.���`&�����ì�y/Ov�qU(�ش��� 7{�9����ڈ�U0>moۀ��%S~C7LRp�(*�	�w���
i��-�}D�뢧�1��@�b�="�"��U�h������8W�.�*��Z�ݘ�tb�[�b��&G����`����y�F��M�!U4	��Y��s��Pw~�J�&��]��&2�:�ς4'�.��M��`5�G�4�-G�6Ӯ�x�P�cx'�x$�ޒ=f�=�]��"MX�!���qb][b���~3� M$g�D�il�t�7���:%0���e�&�u����JDd��!Ȅ
:�[��Ѝ� {����/I�|yW��PI�g�j[���C�ݜ��`�*��MXPzC��y$&ϣ"W,hQ�U�	��t���5�,�tT�5q}�/����p��m}`^m���0�2�alL��N5-@<�N�hD��%8"VXS���iD�?�K�ƚ_�-��;�KG�����.p=��DxA���S�$XV�WV��l��Y!��<jj*� u�Y)`��s0�͓��tJ��wuBIMJ[`C�`�&)�>L�+/N�)VW��U�9�7�U0E:M���'�E685��`��9��_��A9(z ��$5۔c�QU0y�c7���F����	��\���:�/��`��y�{��^.D�^���k��L�����Am�b���N\̖v2�N_��aڨ�C^U�i�bo��m�YS����'������rN[�_���_�2����\Ύ����l��o���V��j��`��/� f9p�g�
�u���}�9 �_�������,f�ME-/X Ò�U���A����0͌kCi�iZ$����W�O�_��WW&N.���(���f>���3�`���!v��f�lr^�G�).a�7a�qI���+�$�V~��aP�ڈ�W��c̟�]�PKX�*�z�`��ג�`#�/QU���P�T�8�DY� �G�B�q�}"a���ɱ��e?����*��:��K�Im�y�.Ii�P6s�g�
�Z3?u�WKy�D��D)�����g����n��\�k˻ߕ��\�Δqm��p�v�ia��v��e��g�ͦ�f�g�8 O�L�.��s��aDMtn��y[��^���ۜӘ��x�]��iˌջuKxP�����P��T��)]�Vԁ]��;��16�~���q�y�`$�^#�v�奈��o�� ������yveE�J�eeʕWk� �mCu6Z��⳴�ՔF�#i���$�Pf���
f�Tu��й���k&�t �O�T+��z|r7�{��Z!dvd���J���.k�Kpp�Ԡ�wζk�ԝ5naVjv��z�{�]�M�z�t97=���+���*=�}�wp~��i8���C�|{��䲌]!���$4�_eM�ű�Sް� %hɶC�U��d���$�c�s��]���Ř�$b&̮yz����l��'д��F,$��Ѻ��,�iS@d�M��ُa��wi���W���j��O\��ͭ��;dSR,�r�=�A�]�ot�LRJd(�r&��p4~8J�"2���_���ɏ���.�%��'���ﴚ��ꑾ�*���.�c���y�Gh��/Ok?�%��I�'e��\3�%�Ëh��Q�(f留\ �X��f*��B)/��ҙ{T�"�[x�:��0y�$�ձ�|�Y�ujS���c�~��	�	pV�9�sdU����fk��p(��跊䑬�ɠ��������*c��*r��D������{Nd/��}�]q�"�Bu�Q��T	ɺCK_kKon��' D@T'I���-��bt;HS�y�����۰:�����io���iA�U+`�(���SM�oc)��'�O��J��7C���������/%���!���y�?z��(�
F4C����A�E�`=/�O!I��lo���TC6�-��z���zNҭ[�*FhBpGtt��O�3~:[��AP��ܫ'	5�ԉ�5__�yHǨox��p�� �����_���b�E��5��{�[��f�.c�#	�ű��k���rv4���,�woԤ���<�T��7�����g��۽5�6���^̩�[9�`����MR������a��}m(���%�;���m���m�︲�8���Ü ��A�>�q��PV�(i����c��������>qVΧT�+��[o�Ȑ�����i"��
��ܣގr}():�l��#�(o��_�Uǯߔ��7'v�i����:<�����A���x@�u�[�h�K��g?�Xt���3�[��z1���22GNW�lx�R�VA&b��Jg`�g���d��K�"��r��6�(�η���v�2��M���IB�̒� �Mv�&��OO�0ӛ�(7�_%�H�����ث
![Cm��x����0���idJ��#�Q1��|\�g�c:}�.��Mw�g�$ǁ&�u5�5a.S�,��~#�u�*8ΧUtm��F���C��1վ��_�3X>;Y�ӻ��f ������V�s6֬kQz#�~/��(��ழm��!X��G࢙�F�W0�zj% �=t�7+kHK�ݶ?dG�@9�5���Jv�i���_��)�hbh�l/���C�.�\1ϕ��(��sA�N���š��^3�R�'���6�Ⱥd�3�Gf�1����k��Y���2I�����y�p@w��a�Ua�>��ΡP�M����|u|��8���5�z��x�}_��AB��v�[�c��:%cC�<���7v���>*��� Og�O��tX����]�V�I��,L���5�tǀsyQ���986�c�.3�� ��2���J*Ii|)L7���Jd�.�5JCF��]D�m<X�+���рy�� p��B�ͦ
"�p7Z�m��x�I�a�ӥ�����0��O�&�q�i����"����?�M�^��@���kVjo2;h�L����AAI�}"3=�O����?x[��D����0_e >L��)O�7��e�2z���o�O֥�$�l�^>7ӽ�(2z�u���o�D�O�h�J@�Z}}`�+}��ԥ& �I4�|��ho�~w����6U�Ή����<���sl�����f�ÿ���e��#@b�{��M�����V�������KH�>��P�a���F=�)u��~���Q)���[�k7�m4H#o���C����~�X7kLV�%���l΂�֪��;/_ԒעU��!�Y��,
�ڸ���I@%/�p�ѳ�sd��t/D�E]��.Ѭ�b{�K�bw�$Y,������/�p���p0e�D Ս��5���1/�`G䧧���b�^���fq|=4mL6:���X9���_cW����Vx���E������t�'.���\hYe�ߦ���=���Qg��Öe
,�5�v�Gu4=y��,3f���¨">��_�k*mQJ*�,��Y��t�Wf���&����פ=��]��'�?���D���A!�:%�H�6N�T���%*���bm��埛vpP-d�fg�E��.I�_�K�d��&�I��R���*�]�/��Ms>��Ω/�A* 
�/ҎWy8�Gr����J��,:�ք.@�3���
ZО+6�G�G׺��J��,�KP�'p��$���7�k�fvx#q)J�Hc��HJ�'�b�ծ�wyW/4ژ��m2@���[�h�L̫-k��2�
j�>P�u�3��W��mvQ�����ہ���F aV�W������7��nN��磖��G�O©4�[4�]�������̋� H�b=��m-:�{��� ��ݡ��Y��xx8��5l/\Ks^|p�eӌ��)ʡ��␪���ObU�UQ9���'�����/A�R�f�7��u������|I�	k�vWTz�Y�>�����B�?I'c$�6��ɶe84+�ٛ���&c(��� �xy)-���(#��%'rE�[ ��e~�:1$��qgw����A1�;ċ�� �w��;؂�d��,�&7"j� N��y�4���� �#ϯ��8� ��t��Omr��N�	6��x��ex<Yv �CТN׾�~���"�+.�jzBr�L�R�%I�7=:~��%r+Pp�(pI����V^4��E,1
��n�##�g���k��aN�_3�f"�pk����瘭}��-3���C|W��v|S�g�z_�_�)��D��B&���*����$;��y+&k�ڶ/� ǂ3/\�N8_Z��}!�P����x=D�y�kx�v��>��������Xb�5v��󓌶�����AO�ZeD��[`HBd\�%��tt}j~$'�B[�_!5���4��4`p0Q�Z5�ucٝ�q��)�Cܾ�5�E�mN�� ߬<N��)U�̼Ҋ/*`��0X��"۾_Kx�6�@�h��1��-�mBp�jq͑]w��^����G*����:}�\x�W��쾅$m��g['jٓ�Q)ԍbL�ٖ!QI�E|�o|�`������#C ?DX�K��T/3��YJ��g�XC�y��:j�9��1���"�:.�xfg�?������H;p�S���5q��8X�(��Q��{���_ۏ97�`0]Xx������(mfxE��1a����!ji�<uj�'-H����߹E�]w�DX�Cu�� aL/�<���_�I��Q�eU[���AR'��;�4�_a���?o�x[^�"z�{:]���ր_Y�Α�<���w�7t|`���5����H�����>��,�N� ΃t،�LYs��0Ib��Bp81�U�|�K�s{K�ş�G��4b��ڜ3����p4-v�]���f�����(Ȅ��hn�����ssEj}���	�Ǿa7�90E�i2��"+s�c����%��������5�=�o^�Q2Gj��|?�?�p'��fE7���=v��P2eܡ��1�Y.Pa�f��h6�4��ʡv$H���]��FK2��w��o{��RC�¦��S��,m�0\H�?K�V��|T��[!��XCp4�\�N�.�i�٦
��=a��q�@YNg�Y1�)%�MD�:A���\�:�Wb����zKi8�����u��{�c8e��;���Dj,Hͱe���s��H�j��U����@��Ġ	"ո_{�7��<-S�T~61�|�4��I��[������BE��G�䊴��9��)JB_�2�+ㄥ��$�ޛoT�I͇y�!8 J�TO�I��+6���֞����H� ��2��HK7��]*n���>�i%d�#j������ܭ�����CR�&���v�A�]q�e�/��hz�P���!X�t�w�
��M2��q��`nŴ�R�_�Ԑh6^˯9�Ɛ0�`����C�E�qra��G���2�.^`E����b����'S9����pL�G���`sN	�Y1�Ye� 󄊲Ujs+��H
��DkZsq���ǹ��@�O�1o�U���$2Zd-� �p�޾6���_���7��V�\��(c�N`_e�hk�ސ�w�I-��c�p�F�ua��~p�ƴ��N�W�K~2��=6SM�~DM� I���F��4��i�*H�{Ԥ������9h��6�nus����Q���IV�@�Pt�co����[�5ɥ��2�v�yܤ�!d��L��Eѷ۬�@�$b��E@'S��]�}.xg�N����!��(�~U��i�͖�U4U�ۆ�����.��'�J�rA���Q�� z��c�'�>�}sLaf̘�7�����U�";���}�h0O�p�0�_�
`��p�d�8�3C������f.�̉,�l��Ѩ�u6<� �C��4w���P�t��m���Z�$ �p�����l�������ltI�r	V�x�-Q��k� ���+�x��Φ+y_��o���ᣜk�pI�W�{ǀ�W���<2.~H�ٌ�3��
W�b���X �"��E��d���_h���C3+`n� ��Ìȿ����<z��!b`�
)�I������띱f�2U|�LW�S島�{�lW���ٔ�<y����:�(o�[��� �:��BZ@͡yg����g��ډ�.�dh�P����ˆ�bXtʥag���s���
�dVҩ�{�]4�/�q�ߔT)r��d?�N��L��B{jC3���UE5 ���מx�Rn�F�]���#T���e�5\ڑ�Q/�&��aR�u��:{�}�ݾ��"ȁs��AO=񕨙n���H}P�'�0��ID�����<�bv�mC�n=?L$OB��U�/�ۏ�����~;�"�5p�xX�:�v�d�h�PA��B|��ȩ�ķ�n��(U���ґ�&��ܬ��m[6�Lx�F�LV������N�T%��19�(0��X��_�����N����LN��"&�ۥV���I��	Y��N|�h;9���=x�>U�e�%��5���P3 ��7C�a@�c9S��k���oa���r杝��'���N�@��G���ՠ�gr�(q��a~G��͢�����[��+&%N�������{�KZf<s�%��.X��^D5h諔��}�xa+�z��}?�v��6׍dx,�,�K�%1x�Q랸��F88_0���߰�1-UF��S�X��r�Em����'��:���*������9�-s��5�2RB�`7
);�/.ea^�[NZ1a�9�������F�a����A��h��3N�'��3�Ԍ=uR^��4����xl� ����߃��p:Ԇ��h4� f�0eU�J��ec�o�����	K͸�Y!h҇�M�x��w�V���g*���j���J��d�>�k&r���Q�b���HP�I��J��ڡ���-�������B˲/|U3�`]p��$��]��D:����a�/��_���}�9�?���1]p�w�|=*�K��L�@����g*�>�@E<�RcF��U�D0Z����:���Vؼ͡��b�WM_C岵�9�Nv�� G-.R:q}�1�+!���a��������
|En��s����:E.)��S6wb}�U��?o�+5�s��[Y�v�oL��
�q7��y$�gA��!j�s�F�J�J��B���`\��g�;�ȧD�B�X�k��-quh�ڹ�>��4��7���dxD���B  {;@�d<�A����o�9��Ȑ�����s�󯁾6�z����l=�i�1���x�K�w@��*��GOl6 a����~��f�ۑ�����O�8~,Y͹�И*���rP�����<�M)�9�Vo�>��G��o@����N���/��(��D��E:�F�����\��W�'���1���u�����J�ײ�T*����s�Uo*�cC9���u��[,�V���abg�&a���� �_��N[$G\N��B�p�(DC��)�w'�s;�&h��UZ�G�+��L�|�˛�>�$$ħ��e�������#�Qo���`��m>X��W-%��gm��vq]ʩ!{t�"c�[��Z>��|0��&� ��@_"a>�����p��e������#��X����1���S����]�Ώ���qA�����].z%2y�F��yp��u��:=!9|��;��63�S�����z�G����ĉ�%?�;���GeD!؏*1~��޻ڱ�4K��խ�ؐ�v����7c}���00t��[�c.���Нu���o[����}��Az�9N����"��8W4o���y����Bv߮���5�,;g6i^�VF�~$���\�9����e{sx�sC�Ј�~g\a�2A@8��V^��Aa"kTE�'_Ej���-�n���j��Ү*�Q:v��E1t3���e��L�P+�rG ��b�7��+uz��۠��C�+I�w!�U�P
̑j˳2�����Q�T�w�8��D���S�,_��N�����?Fu��7<���L���׾Y�	`-�����l]�O����ΰ�l2(����T԰�)�I��H"�E$ �(?��õMk�5��B�Z>{�%�g��r;�of:>�����#���A��I�Q�h�ޗ�F��>u��
���D?��SӰو�:�� E��Y�˝Z�t�ߥkt���1�
'��6�f��6h1]:ovW�n1���|���g���^�����i�Y��tK�j��i%���uN��<@X�w"��wb���E�$���7��DDʞ��2W���J�G��1{�OI���c^�\Ul"<���T�;�V��1f��h�B*������E�G�:��ᮯ��<��ZR����������\���.�����b]��=Rl�'�e�Q��Ę	�L���׋9\>Л��4d��l_��Jqmz
\���n&�!� `�_�G#{cR�S"��e�"Fu����E��/�@�I�"D��HBC�Z1>�9��L�h^b�A2�Ĉ۝�U@!ԑ��v�Jc��y��W;�a�jt�󧂢\�6&C����X�_��#�?n��S��q��g���~����X	ͷc�*ߪ�!�O�����0�u}��*��QA [
����Y���5S�]��j�M7�C'0�(%��.�L�]�xS��~(�@M+�Jt*��O�����*�I���%�a�l��F$4c���4����rw\��Ծ5ٰ�Qҽ���L��E<��OZIը�e9��s�<_3�c����έFeܸ��,�#A�O�� �&�� �qC򬇲=$l:o�����eBueG�f�YG��в� ~���@��$�l ��׆� z�?#n�rB�;��W}16��&�`��S��-	�L�Z�'F?K�R:�^.����5	�I��k����GOlᏛ�d=���%�eھ��1��Ϝ���ϖE���a�g��D�i��Dz��c���-qy>	O�h՗9�_aW��2�f�p������S��h5f�����uYOis�m�%�e����/P�Q/~��;;�x^]uZn�� ��v!�l�!�Z��k�U!K�I�"�h���qd(Tj���UM 5�EE��mqez}Q������ɝΖ��/1w_�K �V������e�՛�pk-3J;Y�}~Ӫ�ڤ�I��l�~G�I O��{m��g�9}�`A��,Ʋa�Lm���nxM���=*�L�I'�o�M"!{p�ŏK^��cNy��V��9<�A/v�ݎ&�������k��8Y�0Q����c�qj���딐�H` ѷ����͸uC�]�!0�0���L��u������4�;ψ��n���$Ĺ��A��{g��������Y�W��DY��<	�����m�Hڥ�T��OjCD�i�Y�L�A:�}y<7ZA�:׀	�!��q��aJ����&Y�m�d��3�gaF��ͫk�>H����#󄕒8��O�����/>��D��n� �
 I���h-���j8RV�`���w�����?f���T�'�4�D��i�a4;�T� �2il_��(%2S�X��0QA"�n�nˢ�
K��-M�:��&p��C�u>���N?N|�YhlCl�C&KtB���y����^�0P�b��v�Ei�4���,7�=z&�?{]�J0������+,�<(�^�^g=��;��R�qd�b{:Xٿ������P��v��ML+v��Cs�Ȍ�w�y�/Q�gz��I�����.�Q����m%G�[���
%�0�a8J4�9�p�3Q3-	}�z��0��X���
`�m���檕$���)M|qha�Û� ��,Cԭ���6�/�Q'����<D�|\d%�[ds����n٧����鳚^��-xղ��:�����AJƔ��"�Ү���ɡ�.��I��@�Tf�}:@d!
��5���?C��p&a�KO4�..�&��4�TLii*�)��i�б<��.3�P�ϡ �v?`1L �g[��w��c K/�bE�%� _�`�@ʍ��BəXT��ۃ B4o�ERt���:��t��%~4���1+���Z?������:,x��U�!���ӘT|{��H�Oh
˘�U� p_'� ������,sgma8[�CuG�Š��,%��w.37�^e�g�:�X3҉�BͿXV����W��3�X����1lLV�V/���3�d>*����v�\O��Eb��:6�4v}�(z�o�C����:�0"D!NJ��B昍���f�9���nb�!a�w�R�U䅯��:�s��� v�<[%��1,����g�η�ft�^<��#�2kk��|��5���֔иX�M�(nv�����n"���T�����U�19r�D���z��WB��v�l�B��!��������ҙ�i���/m�l]�os���������.M�W�QqO^M�y�eYg�g�<��͹�W�����#p1UQ+v���[}D��>��Eq��������V�F�t�@�R2��T��  Χ)5be n?�V��H^��L�:%�a��|}�YN!��)�$�0靹��5�26�+X�����}U�!h�Y� }�����7�A-gf��~Gn09��)$mqU�[>9)#M��-�99�bR�{qV���N_�X��}ٖ�+C�V�>�	��R#[b��U(�h6��xAӢ���2����V�&ҭ^�������s�#O^�q�A�+{Bv0u���r���^�*x}���l����cO����RF����sǯm��Vbt�fC� ����A�� |��b�I��77�Mل�{a��s)�F!�p��z�Y�����]��˨Yؙ�xi���oɳ��M�	��L\�0�� �$�tb)��B��^*^�P<_C[������,�yx}n��&3�U�g�*���3q�w�x�������̷�[�_h��Uφ�~u�\=C'}����I8ｅ�m�M��r�"}��7���Vc}���!0�	x��B>���({���.��{�t���)����D��X 緊��������[��oz�c���/�IB2h�B�<��QQO��Ì��p��t9�1;^
����OKЮl��HUX������N��XG���K�j���c���'��Mp����P�H���`��P�Or ��5X�п��c{9z�QG�'�6�,%Zg�lr������$�3|���|c���&/��_C�ٜ�k��ئO�@T������T_$vk�i݆ I+������_wEGnM�&�1��|T:���qb{4��0�?��^z}��*t�����ծ�L`U �@����_���a`�Z�� �[�֥�#&�`�WtrX��N�9�X�N�9Ko�R��KK�/E��f���QȔ��5�����Ew"��$���F�	�射��A��h##�5:��M�3�1'�˲�t�Vt��@�{:���2eV��� �y@��5x�k/���	C���@�Xj�O���Y{%6���j���9Ͻ���������'��5�^ܡx��{M��ۦ��7��)I[��ubP�^Ǣ���s'���`eޝ��9U�8����į��naO#^��f�`#եL����I��	g�.
���K�d�?�b.��S��[-�֜��i���H�3��a���Y�i�еΌc�&�Pحz����6-;�٩>�17:b_������F�ƶH:�'
Z!���;}y	G�O�rM 0 ��/�A	B��ԗ�����N����I@L���3��i~�>���0�s&��4�v�p.���%X�L^w��
����¦��C� ��?�Gx3n��q��lh�.����%��ԫ�Wb�K�e!��S�jF�� 8��������nѕj�����U�
s{���� �����M�l�2a���w��"/��7��_����;�J��8W���7����׾�6 �f�h|��BlNx���?F@��Q9" ㅕo~�=2֝��M�F������;�R�S���t��I�Hy#�����e���G�W���XböikM�'@Vm�h���w��������O�aW��C���% =C�������߁�C�K�p����0�7*�2<d_�� ���?È���xe��}��4����p>����^Ȱ���~u�}�i;'����m��P�Jlޤ'S��Y"�q�<?��E�B�m�s��S1��o�]CvY���P4�����xY�)��r�z)�8��=��Wrm��m19I��;�h<k�b���e�|�C�ηw,M�].��Øܟ#��*٫�6�[�9��#T�㾔_[������L��vx"y�b6h���1��yd��ډIk+YyD�zM(-O�*[4���QG���hW���[�תL��"�(-��r����,��S��G��A����!�T���ժ#�������%*���p�~�YpHeh�hZ%�~WQ�?+����)&�Cĥ���@�e�J�%�� ��4�D1ݤ��^y�⌆���J�s�����E�'��eG�l�vn�F�w��z�a7�.���dÿ�#��������I�Ԗ�F�owb�K��Pxc�l�fo���R��~f�.�>i�ӬUU4�
�E0�	RFm�c!1VïmS�	���A�:��M����ذaΊHYY�H4���a^�hl��@v��a�����v2,�u7�f�� LhMa�lA*�@��������@jS�>px�a��-U�K��{�=N�Z����p��5y�>�<�]y�<�ؖ@�S���>��� \�zy��1;�������5�b���çI^��� �D���t��������������r��x*��a��)b�f�v]��m���*�Tu�?(Q�	�9y	��K�Z���.��|��;A�Q�"A�?r;�C�*QZ�5�p)�d�2ᜨ��H�ۡS�w�+O��Q�-լ����Ѭ*h�a��<�j�!�ch+�o�6��<����!HĆy����7��J}WQ��y��ţ���D|z�� �����D� �y�<��W��m�s!�@2E�i		��}M�H����mi�1�V	��tÎ�Bi�h�P�MO�2�&;�|+#԰tL�t/r��Ă&��L��g�bU����9FyuQ��$|*$���Ä*��l��Zo���3C��>�mm��,�ȉP瑃e�9�YT\�FKH��9��*�N�e���;J�kA�h��Ǥ��D��f���J�ä�C����$�Q��	�<�pո��7�]���o�Q4���3�A't������]���(H�!+޶�r�=n:0R0��{M��:�4�*yz�������%X��N{�s�K[ǒɋ�H��.��6z�}�B}�:I���4(��J���Ε��noX�U8���S�&�w���(�?nz��}���8�n>��͕���>8��H� �zGq�M卤��n�^F�s�Sk^~�̫MDcE���t�<�\��x�rz:�[XJc2j:�6�L/	
�h;���\�c�#�-ߚ9S�B
�{���y9 ~�>�W�r��h���E[|�Wn�ÈY)�ӌ�6�¥��%���'0̂0��IC�D�M�����J����@�8x�H`t,L�0�S�θ�9���ڌ�g����[t������f�����Fz�__�) � ������hd��.��'(��қ�;UQ+�J4��ۉ)e�M��Lj�J%BO8ׯ���������U}Z7�8�=�Ss÷�[¥�@���	�W��q�ו,��E ^ˠ���=�t'/��4�pv(e�jF��E���������At۷�=�?FS�/�CnU���%����l2��{�\��mW�s�0��f71�-�ZW����3k}��C�~6��q���o,Q
�f�S.z��8��K	n8�B��zGϨ��a�3��,RN���S�k�G��r���j�9��A@��t�4w��m��>�;�����{��S�]HӤ�n���pU�^i��!oT-޺�Mԏ䍺�(7y�k*s�5د�����~�J)i�i����E#���܋�QB�z;�r�A��-R�g6�&��~�ٮ��lo��
��E^j验I9����,&�/�y[h9fkE�Z!YW�[�уIb����M����Ó3�^�n>�5���@i��]$�;K�i��m�O=�&�-W�����+���8�ő_�qƂov �v0�}B�p�0b��ȍ���?�z��3��jW¸<����TŢ��Q ޱ5�/��g`�{5���s8�*�Sa�
�*��F>�By��-�vUy�� @�Q��xZ�qC}e.dE����l$�>�t��n�3l'vO�*�i����5U5f�ͺ��K>�Qw��Z��b�n|[�����'��G:�1��/wU"���%���g�,�~��Z~���z큀����w�K���e nȢ7&��l�6�q�g�ls�q��`h/�0�Z ��-�ݻ�h�g��@�JwPp���1������D�d�>Hk~	���L�_?�Ph9l�[�x`�cG닣Mβb43-���h]�0�&D���Y�r?H���n�ѐ��ьJ��*��6��"��j"p����vq�v���|<g��0b��M�F��C9�#mbp�a_����� N�r�ZE�ΩjO�P�J���;�
��A��	���ӮV+ːh�vx��٦Â�&em���cR9�J� Qu���Y�"4'8gY�i5͊�l�����^o�������{և��+�a"�c��`wr��wy�����A�n������­R�;����������q�+�b�x�A5V�4�S~��F��7,����6+��J�h���'hB��Zn�z��c����t��|`NL;W���Pt6_�ҭ���N���U��� 7��KrL�?'��6{i�hwR吜�X�Scrm�j�ĺ��|�D��q]�al��0�W�)|G����
��G�� �pH}���^�fVQ�#���OIq�
�ȓyC��i��,��ks
y�BՍ9kly��N&�3@/)J�<�G�j�:��a�
��i��Ѽ�D������?i�l�*����q.���Q�2T(G�Ȅ�ڃ6�7�JE�f��J�Qx��c���.nG�8��!�7�@��;�Ύ�Sqtۯ�r�����>��Av�"�`�cR�p %׬}ߛ>b�t�Q�(Ae�E�*<0�~�Kߚ�uk�Y���W��~�3��������.M� ݻh����d15�Ǉ�S��[������ЈwH7h8ͫ�� {%���P����ǝ.��NbD������4�b��)����7���z�+m�$�J	�Bh�)��/����N���t8���(�Rx0�A 0m)����}%?�g*�겲:z�̑Aw 9�%;!�7$��(�s+��s���o5׆��e($
Uo#%d�t�9�T�mK�3�e;H�[w*�ì�(75�l��[����0۴����5>H��Շ%lF�S_$ޜln6!��y�&��-���p��~Ouo���w�-L����F:6M��ei�u�0V].���%̺z"3�Ss��ѼT�7����=^��C"���:9������7	m�%T����ʪb�!?+��Y�b[��ɾ�
��~�-�ړw�m3 ���R�q�p�ѠIg|�q�PI��a�7:��pË<������\��J����z�J��I�1�u�j��UHUUG�
~�9�{�L���:��D,ѵ�v$ڰ��Z���?���`ۋ���xL���ږ�q����H��W�y��AR@�=[%i�K���HE� �2���`�m�zDȤZ/)$�^��lI��a��R�����vA�Y�����٥:���|)|�cY�B�c|����H�q]C�����gA��hU���0�b�C8� ���eT�5�"Rm��u5�v�\=�lB,�������^�Oi��v��9N��q�ׄ� ��$A�Y��J�t&j��!��Џ�k�ŘՒ��e�g���R�<�N5T�͉���:���:b��]e.h�!&��@ظ���Լe��S�mZ0����>ڿ���2�i�\3W�#��h��5t����{[�uJ��
J�+S@�f�K�F���R�:L�G[��}��D��yv jPJ��u����[2X�a�����R�p^7���x���jl5�����Q���0�$H�?�$A�md7��,j��d͊S�?�".�����%��׬�K�b�xִ����&s����_�$���)����V:�LP�s�~%�������KC}V�P3M%��Ƙ7=GJܛ�\t�� �aU7�����˂1CS{Y�Vȭ�V��.{�w}�����RO��Er�f�_?�o����3�*ka�.cr�F�.�*Hy�y�]�'�w�u�z�rŢ4ApȔ��q�gc�fo,�)�3nUR����t,�w�#9Z��(B�>��N77~����3I�NBϨ�Q��E���������+�=�p�\W�۴�w����^ńп�{�
�2D9�b��r��G����M��tk*t5�Y����G�'9�Ʀ�C��ů���(n��a	�S_8 x�6�
�2�NpM'%��4J��ӥ�EΖbR��3�[%����g֐u�=r�_�����h�=��8��W##���x�7����	�� 9Zg��T9�E��a[ˤ#����&�䏝�2�K��f´�>��'��U�+����I c��s|m%�o�}A�v,�vd��@�L�{�L����0h]�|�����t��$ÿ[:�S��ˇ<�?�pxUZ�Y̗��z��VM��4TU�&����U�_��1]lp^��7|ب;�8.Aq���f�ok��M!��e7H�(�K"_H��U�T	����EI��s�����9+K���S�t��BU�{Y�pί�Q{?�>a	���v�sTg���S�G"S��C�[�����il�k�%`���%�5�H��k�pԜ<����T�WD�2��;�b�NY���6�4�l�i�
���7�h�!b�V�]x�q�1�D}�;�������}7�*�_I�y^@�k�u���e� �
0��؅y����q>Y��˕���)�����U�'�-%?��z�tP��Ǟ�������E=��?�2�h���Xʾ�L�Jl�nO_�az�0��o���}M&5 ���3.��H}�����E׫7�DPTv1�Rl�)��V�n��&�Lh�dN/B�Au�)�����j�oɽ�&������q;�g���$�����&�)�T��⡝����[L���iw��lJg���Y�˘��ͫ���ܱ*{�%���U~@��g�d�ſJ[��\{��n������70�3�n/��YU-ۀ2쨾�ELv渳���}:]$����,N	8��=�M|�2����O`7��/�t�� `!]D�)�:��0�:!�עj;�d%��f�����9�hi19����r�@��D\;�� �'�����hْ�a�a�s|������g��=�Ը�������M8G��~ �p�W)zr�G(쏜��n��0ZX��u2`�2�Ա.�Iz��w�+�Sd(��"� lj�k�0�J2^��|	H�D�7S7*���L�I1�hN�7H��̰S<�C��[kb˅�-zXr	�q�q�a�?�'���I�I�l����H��8X+�Ga�/���� ���[A�E{\�zX���;���,!��Y"п0�p@�}���\����9�eΤv�,�����~�bM��r�B�q�bv��Ѐlx�����I,ɂ9��[]9<�RM�kU�:������:\_�ƞ�"���-#:�qCcJ'��q+�C�=�K��(��:=čd��)l�>"�d��k?�)f��S�vU��立���ٌ�Դ*iv�mۂO���k��-�c�c�XZ<������DQh%�2�
.���bJ������J��S�f'�h�pښ���X&��ܝ���]U3Ic�	_b��k�����9=�W�`�]��|*���0%�i����f[� �3~����{,+��A���;������u+��O4W�H�>��p�ߢ�76P�Q��G�6�{-��D�l���й���~UѸ�ی�	��wT�%�"/�;��}�lA��O�ʾ���T�Pj.�L�UG�,l�ߌC��7I�;��~w����y��<z�S�C�<�3��R���/D�
�m"��֙Q��S���wKΆ6V���P'F�
�����f̞�X�|bIs=�-�W���+��?�#;���rTfk�m�x�:���ij��31iB���y 	��/^C�I�n�*}�p$mQ@ӽ�yh~�X9}�����x!��a%�

\��+c�d%a�77�����N�ȗ?�M  �����Mp�
'��3��py ��j
��j_�q������n�`4^Y0CP�nHh�J4X�0��s�V܌��Q���(]��6R5F������yYY������{���=t%_؎��v	>���NX�w)+uɗdqP��QC�3��W�8���-���LK�*�ཛFt����|>��'w��=�"�f"�<J+w:�ۡ�˜Ơ������:�0&����.J�]��#�Ŋ��s_�K�-��ܓa�) ƪ#X�г$�����ˣ�RX���
�������9�)û�Ix����	����_�џ��StVi��mg���)z;[t�H`2�^�cf���|n�S֍*���C�ix��N����(��'��RH7�uc�V�5F��P=�]�����,x9�c/���K>�E/��Q`P�b�R��{�HIs�����~�6��ي���%����g`$o6�p&�F��J���a/.��լ�e��>���Ȱ:b�����㣐�:v��[���idU\�����ܷk��Q�/���E[�u�����XZ�l���2�h��Smee�(Oq�Qk��(~ 8~�Y��k6��ޣ�*������Zi"�a�/i�P�ou�;���8vCs�rwI+�cQ�u�Uc$ܴm���G�nN���/J���Q��,3of8�Y�ʁ\a�v0�/����qK=��V�����ʄ�>�����}�� 1c53`k���%$U-Y�H����pt-�P�����7�P`�)���/
���	3��bK�x����1�!�)��-)Zӂf���b�6���[�ꆆ>PY�d�3��v|�o �^�>Bg�z��ƶ��a�D��⡕K5`"���0�\t���O�t�{!�o����pg��!2}$|�a�s;�%�),�YN7rD>R�i+�&�Ap ����ʋ��v�����3�$�%'6b�$��O3y�r�K�9�~�ur�H5��Th^���T�q?�Y\�B�z �@�e����:�U�=���0j��e�P\��R� &.�Z�y����f�~d�ĀBXHU	+m�i����^��agEQ��)�K��{T�|)��a4�ٮ�+�rq=�i)�A�ͼa-}H^86��k�`�m�6�rT�yma�-g���4»3g/R���N&ҶC��oQ����F��M1i-�c{�{ ed2�o����翌&0��v�{џr�$�;�f�.�����bI��BSB�B�9֢�"��6j9ќ����ؿ���ςt]���/atG"�_����j�.�J��E���QH�����A̩��r��H�B���X?���ʾ�?i��yw#OQ����o�m�&�q|9�Q ����{��}r%̅G�J���\(urX � >&� :�4z��{��;���s��Y�pub;���1,l�44N���54�����<���,�UDm+��q�¼�F�ߩK[pHl qx�L��D?g%��Ϫ����]f����S����C���4�Yi�zi
G/�*����
��9�����Nu�S�Y����*B���Xq�oY���̽ Ma�'O�,��y]��h�~������U�,U��5�|� \*��4����ysK���Q����ۍF�F��Eo���<)�"�)���V:s@��VE�=bm���@*�M����G�rXO1j֏����-�Y��ՠ�� �{�0�ٹ������S<�SbU`��`[
h���<�C�d��0�(sG�A9�4��s��3��04x9|�m'vr��U�B-���N��x����;F��h�]C%m�&�[���M琴G�܊e���F�5���+�ҍ	������z�'�����i脈&D�x��?B��\��2pͨ,�O���g�`�����j���1'��I ���{1lM\��9���8�d���^_(�$��'���y�e�S�)��bN�53%�^jf����a���2��l�k��P��2LZb,�]�k��
�U��J,�>��+��sT�E~����F����,5��y3��5N�O��&�m���j]|ա%u�%���%��&AО���|v�*0iѪwt-S/N�{��I9��e��4n�T�������9�i'u����eIN�'u�D�a�E$�ѽ��aSYY�Q��P�Uv����oe,z��pU�1��5�iR�F���^�7�)af�1�m�ѕ���^'G�t:��������YT��C3F)�?^��RJDo�D���!��ϛ��F�o9�<sGCތE�^K͡	�BD-�PCC�{ٺ萊��fN�p m3��c5��"J���þ��X��L��X��)��X5{w/q��ߛ�¥31�e\NN���y̰���u)i�J��E�B������n�GӬȝ:�h����£� -`�s8�t�\�~\��Ԫ��1	f�E�?��4Te.���D�TH�V�$�|1F/�
�7:%�?hCDD�a�	��\��z:,b/}�Ai^�I��E��&B�>��ٌa�2�����\<��'W�AA%��%�Bq�@��0�~�(����[���*�d���g�ꆉ�p���EG����~���y�$�N���h���얦SA��I.�Y��6<��V8��&��x���b� ���f���wvgK�Eɳ)�Gg;�^hr�L�Q��Q&}<O1u;)�݉��~��dt7��er(5�<J��2�#����  rn��}:)=�P��A+�S:�U�S�1���"F��,<e	a�A�q���]͟���������X-c�䐤��(B��I�{�rgP��ꜹA*�h"7�ʭ��q�0��a4Z��M��E�t�_�i���t\�K(s)N<�W�?"1�����xD�z�"D��Bf���ʎ��R���I�
�4�&�)�k_©�j�����<glj����-�`~+H��W1=��eڟ�e*H+x��}�r4����r���_M(]����1�~_D'�wn76ɩ�`�M�F$��h��T��]��u�ә8y��n�f֔Gn�����g�Ikn8Y
�C:�ь�=�1Lj��9�A�r�4R/�-f�JJ���	�o����/8R���b���4����ho�+��k��D�����
��wV�`J��aV��!�gԫ��i����|���Yqӽ�f���Eā�f�w�zڝ���	(x��ْ'/T��݌B�j���wO5��~�-��$�����ݿҲ/�`�A"pg�cr��!Ȍ+��.i!�g�oEăRVF���h��g9�0ڡ�����G|ݬe!#d�z����-����#i��sݗSr���V�³�B��X�d�s�}�1&�Y�lW��7Z�0����%_�r�T�� ���E>o�����p%T�n�Q��̇D,n�$��~|x��t��md���Ժ�1�pd�3�HD
�,�d9*�a���֣9]I_�ʬ1����W�"�dQ"���!-�u�1���rm]N��d�*���g��x>�w��A��K$����2nM���3l��֢Jp "�Y����~MO�c���a�a�ۅ$���r�W� ,I�%�6G���ۘEq���?iѝK��y�٭P����$�WC�ޡ�2�PZ�7���@*�ʡY�&���P8��y�m��;ouA(hW������'�(���lȪ�+k�sM���Ej�:�q����h�o�,M��J=qRD��v&���U�ڧU�Rj�E1˻�4t����@f8��d�O�&>:��� �eeA���A��u���I�:�������av8	��2������xv�<����8�ǥn�ĳdi�:�l��@�,Y���}�g�����v��U89�
jo��eI;��z����(������d���*�=VB�	%�C%o�?qn6�&��g��U��`� ��pSǀ�������"�[cxA�r�]�ݶ�����՛G=�<.��=(7�E����T�ab�ϩ�~���+��@���3�� �N�@s����L�w:M�RZ����4��Ɇ��fVw�!��O�0��Y��w �,3G#2���P�=��w�W�L��� ��TD��}Ɗ�Gt�D!:�+*��6���������d����̂b�$�����[�UM��b�T-���x��!7�"	���P�p�0ot���w�^ �_��;���?�ެu�s�Y����uh�p�C_�˸ܝ��ћ�R^�.U �VH0���<RDJc�C�m�O+�D�7O\by����k���ĩ˗�bz�蠺��-�o�&O���Ap�"w4V�lD�#/�t��|=J M����$����Zs;8!ܨ�y�>�L��[��03�M~V���h�wV�S�s;���'�@��	��%�-����	�A���H�#�T��k��<��ûY5�P/n��_��@�j�֗M6;�������l:}앲%mU�$X�G3U�˳"/-5�m2v4/Ė�5�1���U��V.յe�"|-T��օ$��ɥ��x�${�(I�\͌~�=ĺ�]��q1��E��H�?-���0P��j��`_�e�o⎬�7����p8o��E��x�!/�t��n�T�p�0��ڹHYv��a>ap���zhW��=��c��\s.Ecφ���A��7n�cD�t���PYs�t|-��l� s'�'YBy\������;.��.e�������j����L�:�~���#��6�G����s7�D�j����Ɨ��tG6��* Q��f��y�����|�t��S0���W��y��ʳ\ ��'���}1(�/!��𳮥6� #��z�����IڡJ>�tj���Z�m���j	^{_����}��%�������`�|��A:�7��#����O^v���@�w���Yԍ�~��߽��̂SȪ��������ķl'�i��CQg���|�g�`"�X�j�앓j_��oc\`���Br�ͻ��5���L�S��Py�ӃS�6�NC�Al���X�t�@���	��i��6���8�����:��Q�FE+p�`�z����m��p��1&(�l��S',�6�?\:��V�