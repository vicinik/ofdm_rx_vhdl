��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��8&����
/BZ W�� z��L���]�9[Pk��kO�c�W{BH��^"l�J���߲�GM�b��IL�����g$��@����c�E��J������Is�@j�z��^�����p8�ɵ�FDqLT7�'Q�)�D��xX!SD�f��W��v�=� ?���1Gj����|7�t���r{����C�<��L*�W*﩮9x�Z��ǡ���~���zl9	)T��|�I� B�)��??�Ǚ�sZ���u.��4=�y��CÅ��R��	L[�3n�ƵNjK�_����7qc}����a�e[�Lu����Ad�9l�q�+Ǚ��'ʝ7bjl���Ŷ1`t�'%��k6���.E��K��T�tO�N��˷r�p{��YF��J�7��_>OT4��(��S�@$<�N��+uW�&�"��JM�`x�{��}�� ��6��n�hj��}���'��f��ń�\I�:��^������z瘔�]���c�ry/�|�=EFM_�$U�+l�WP�o����³gw�x�5*�z4F��W�rڧ��xH��ݡ��"�lGT�A�sct+7���^'�g���9ַ���":y�ܣ�E�a<<N���9Ln�3��(4���Ǉ�s����eP����3��YNxL�^{9"�� �Sz�i���\�0���7����[��ɴ'ӣ�&���K>Fm��C�� i�zr�<�d�
å��tV�k���ZR�H�2� zM�c��Y��:�w��`���}C<�JىF�� �ݨ7��\V�i�7�_9��+��?�*��1k<�i�c
�ҡQ����ٟ��n)�7��|r3�# �C���!�߾U:ڛG�C�~&����[��dQ��(��A�5�
�z�����)t���⸿��zOɄHKx�N���*__FH��a��q�-�Ļ T�,��
��x�UoOk�
�h2
�1~d�na� IMgUn��طf?;S��Z�Oz�5b΢YP��j�G�{�.�O�[�k0Rk�F-ZQcjbا����@T�7`�UE4D�˟e��_���А�
���zP�8��U��R>����^�e�P�NXL�86��Z�~]��G��nE���ɽ0���{��"���	Is�pP�}T�0�����}L�cܒ��ȆCV�o�y.��o=ˣ���_����Lh�IJ��P��Ww�݄�����:�<C����p;�[ޫކnB��>��.L�o��2�ocO#£�Gu%ؐ7ŉ:%i��1��+�{sߎ����t�F��doP�W��s�e`: ��m�P�֜�����Ɋ�90�gh��1��W�+�ǘB���d����zNŚ.�a�K�����Ȟgl|4���
�Eˈ_�z�t ��r�0�{M3��/帇��e��Ž`��*ک:bm�	�PP��X�K�1R��3S�� aB-���}�3�4�4��h���I�GaxF0vNB#��?��I롮b)������|��W�3�
,/D�|.��s�nZ2�#突jKR�34��N���AF�/�S���˽�����O�ō^q����^d��5�vq¯w�zX�&�4� Q_�)hs[7�fN̻�*�}-�A�jr�Ŧ�CB�����Go���c�c�\ĵs�Si	B�>08�*s�R��ٞWy��;��uO�3q���
Y��`����Z��η�SAb�`�����
kY�*�1
����}>H�ku߈���I�b�VL��>�}T�n����ƺV";�/��k��DS�����!��5C
�$�\U2�� ?�� �7�t�"	�Ͱ(�6��U��W�XFf���pQe@	����]-;��]җ�\O�x��Ɣ^�ݟ�"���v�bs+�J����N9DI�Q7_�?8Ȍ3JU��cV��#MsHO%�G8y��;;���B�V�i,↵��H^c(�&$�5��LZ�@�H��b�i~LnN^ꥥ���e�� ���6x�o���T��=��o�FM���=����v��i�upRN���ĝ�~K,���0��a��U?%i���N�5j��t��W���x"+�[L�S���a�D�,k$mo�R=��r�h�hȑ��2[�W�(��k�U�����^� _J"�9�Ȭ�]������؏i��5��}�u���5;�J��Z�_��BF���&�z���Ae3�;�ؕ�����-�v���=$�QuW���y���+r/{�pq���uI[젌�.91��4`&�/'��Ǯ�F�a�M%�N��1x��L`{�
s9�\��{�g"��$�α�� ��?�1��
P7o̾��3�cڵ��/3]�iޣ��j^]��O��:��3U[�M�}��xn���uqd���6�Vk�nv�����Ylu�������"6pZ!��@�N4�r"p��\ukШ��,�g��A��MX���3��B������ێ�R!�Z*^GT�)P"C��ф�]�9Nui�5 �v����8(ox����&}�D��P�V��fLB���9�$���(���3`����s�*B��O���k�%��0���/wJ5��;`�7�4��|Ƥ�V�ؽNޙ-\l D�~��d1�����'P��� �@�=��Z�A�����Kc��fc�w+1x��n�b����׷�7�d��T;s�l&�O�I��C��%��Pe�ZK|�,؈4��� �L���Q3:fzMv&e~<�/U��Bd2��F��`Z�xp{χ*�M? �Td�$c'�����>nd'������2G)��O�F�h�f3�3�`V�8p�W�γ��,�#��!�K���p����X���]��t�!���ջ�J�pL�3�U3�٨|��6Έ4�4'������U0
��҄�~���=�u�[L�%�~Xr�,���Ro����P*%yv_��II���$��Y��&���c�a����kP&����j��C߯�q3�-yq<	�ة��.���3�Īۭh{�z�mR,f��h�YNV�P KW�"�:{V��2����Ĵ��ڦ:A�F;2R�[�4��%[*A��83�����O��2�_�����q�,��mh#'����M+���db��T��{)�S���#�4����*e�]�EWk�
��e�W��M ��`sB�Ge*+��Kl�<U�����+]7j�Ә(��ת1[�0�6)KoN�k�8{���G���$s�����ڡu�6x��k���/Q�_��u��̍�O�p�+G�����paH̋�g�q�u�����D;��o�?�F�sJu;��K��̠�T�ȑ��%	��p�bF��}N)�#���,.o�|�v��/(_L����P��5�=�8����ӎ}Ў%ۣ$UU��T�Ju�(�t.\�h�7O�Iz��Ǳ �P�	���h\���3���/�w!9��`�bt#
1�
��e)�lm�{���B��㪣fC��ߋs�Mh�Uo��$�aJ��.K��"��>t��$+�;G 1��.�+�,@׍,��M�0����:L� ����C��+;6�y�o��m+Mh��F�N&0�cGw�%��}E��Z�r~�k�� ��K�k1���և6�(��2O�r-Ty��^��w��� �����h�(م�����n@��r-�b"��c�Y�/s#~��b�
-@�\k��죕�ey�:8DR�9��>^��_!��V��5&Ǩ�K؂���_��ء��fS�Z.��7"�J��េ8>�r�����6v�F�6.-�?-�P�o�$�Ǌ&�0x�7�Z����իpu��L�q˔��M h8<�H�}���KW��D�l��^���F@�m(äR��ݍ��Ij�~/³�G`$cT^�3(�3K,�&I��0e�:{g�o��)=�	o��K�4Ɇ���B�M��(��m���W�]
�\d�i�6R�?dLK��<�h��Kʧ���H�#���f�Y
D�����O\�Y"�^��>K�ﱥ
� X$���f�����[��K���� �%�ơ\�8ݲ��=�<P�0
���,#U�v �s��U	�n
>]���G�熹d�1����������&�����Zzsx�:aH��~˲C���X#��坛Q=���|�Q<�?z1m� 6��e�Fl��l8m�z�*���ޢL4V~�k��$^��̻Ϧf81qoT�W��Z��2L5q�,B^�t���K#��a�.ІE���C��	AnPu�؞ ��U]���	u�+<�<^x����A��+��
�������,X��|_�,?�X'���*�YU�+��eM�l����|a�©*�Bgo�U#�Eu�{dn�)�"��ٲ����[�-Ѹ�Y���Gj |�G�Ď�$k��>��˫yq�s Ϩ��� �K���O���b+��A�՗�1��+����3��|��X��p
�#oC�6
#!���������R�T���3>�Yv��\Nzs|�B��m�1�έW=\GF<�3�/��
�]"�W�E��<���>Nj����+�yh�2�_�j���7��1'>G!(����D�] Cx|���W�w�T�
��k�ll�ѧ?Ls��E�X)�G�9S,F����4o�u6��� X�pO�<�<_,�ad��o�5���@7y�3�v#pH�ӲQ%O3�Cm�H�Q[2g�$a�̡%� ��E
W:���TL~>�K��|&�-Z��(�Tr�v�v����;�1����&n><ʯ���ʲ����3=.���>`L�535�=B���^�Q�Wb�.��x�:��C����kXe��e£y�3N��.���>I�,ˉ6��N��3~!΍��1�*�{�+w¥t�\��� �*�ʫA�᱔��k��D�_�@������'�����7�Q!O
�[�L*mVBp�w%�a����9��J�rw$���בIh����B/��߿86�rOiH���V�ԥ8$@��k�R�R������^AS3ڱkG3�Z����u�����MXׂmL���- �>_�U�5q-�!��fpY��_G�	�+	@��M	����5��]� �A_���X qAk�#���_G�L����O�9�"~9B��܉���oY<��]��8��md���jܷl��:���J��B\�m~��إ�ҷ̝���?��)�-˭�����z9zXֶ}x����`�5��A�(YZ�	�&��x�\(�E����c�J.{��Bm��4۸���{'��y0��5����i�����㍎f�5|��� H�BMU���7�ê�@���Cs���#Z�y5�w<"#��\�';w�@	��꠆qz�j��ϼ��(�P�qM��I�f��Q��g0�5����8ҙC��3G���ݟ%�a.OX$����Y�V}�'iR�0]&�$���z��f�v�ūs5�l
TVtïV4
y���
�+z�0gkΔ(QFm����-��4}e�{��dKTw\
o�w��FC'{[q�Rh�2H�]h�a�=��g�_���mN������hak��Q\�H����t����k�Ѐʐ�Z��`!fY���������6����x��ʴ������o�=�Un �)�e7]�&�l_��X/[%�D�Kb�L��B���,��;��smH��X�<�ZF`�x|�E::^� �	]w�q�̻�g�1��&��T	����,'}�+��W��K�KmF�ө6��և�vt�K	x�=&U�|�}߭����cA����0�m�S~O�a�&�/ 2�7[��O�Dl�� F+6�]��M���ܿW���+:���&���h���/x�A1B(��nQl[2!6��*�s�p�Z�f��F�����BE��+M��UU[�s�G�Q��3	6ϙ�J�=I:�یl�	����:���?�����a�z(Y>~���D��9:֛���b\�4�"�i�2���Dv{��Q<A�xK:��Dha�$��66���l�	�`Ե6���x�ÏL��r~�ޢ�~���*ȗB�ێ��x���̻��euM6\HbVa$s����{�G�{���s�ۻ�VC=Pm"R[�mI8ϡ=R��ZD�,W�ן�K��k �j�~�o�0Ra��Y�Ǩ�Z�5D�����K4H���(#�<��g�������J�@������V������ʥY�����j��;X!�rw���H`�ks*/z�����枩Cݦ_;n0��>�Z����M�dr�;�J�<(_�����X�1�k� ���</�Ǳ>)j�7�!�b>�L��-�bZ*�ւC4êx
��E�b}�3����yH�9��Qٌ(5��Ÿ�gJ��ZFh�Y�5X� � �o:��u�������8>���⍣ �_�N�Dy'?:w:h���.�(����M&�}�/�p��?J&8�8��-��T.{x��R=-�F*��cV�`"�sM�I�ъp3M�\��\�G�r�;�rV�؈ʳ֥�(���K�h�����y�v"�.�����Z0�>��i8a%�wU;��$|�����9��������f���i��G�]�(_v`�a�3�����8��,kx��~,�H�Y{��f�tش�U	�h�ͳ�^�=��.X��`�L�T�����JI7i�\��U������0��4��t��9`�}��i��C����\Ի��Ĥ尢�ˀ��
���ũ�
������>�=��*�a�X�~����~>!��o��8�X��'5?.B2~��X���z����/�82�m��_�j������~���ǉ�f����Ǿ9p�3�zl;b�X�Y��Ӭ�4��_���JE�`�W��f�&����XgC����#��Ɋ����Ma�,��}�t̀�М�T�4t1�ל�X@���`w{��^BIn�1"5|N�2B��H������!�y���v������\���^�A��8���W@��S�È��nf=קɚ8�fz�Q��� �{C�|�R���M���4<Bp3��1yk������a�h�q$[�d�M
fN�S]��ё<\a����)M�eCD���g+�K������sa\�LH��U4*�=��" �*��F����W�9Gj_��eG8H�)֤:�]��p"��"�	��M�[Zp �J�!ڇ���NC1i:IfC��1>�
�#��`�vƪ�,��p}ն�O&��4xxa)<��(GtR��k������a�p4�a�4�бĐ	��i$�t�|��Hڮ���8	��gr����I�o��O��f�����Z�5APFr���So>̈#Q��as��L��M'и��6��/�P������-n�R���ރ^�_ 8��V�xSu���*o��m��� ��l8k��~�!�V:��l�7tC_�i���J���2�j�,c�Ŗ�#�n�^�@��z��$�����q"�n!��|A,)[�lGZG�mjeF��&O�&�oa}8/�����w4*5��F���xuH�+v��-E\g��Ά�cv�����/�nM�ݞ�ƚ����#T�T�g��gÙ���b<HÒ⳧w�x�o��I*R�yd�F2zw�I�cF����ؙ�� {;~�=��p��ڋ�"�Z����h�i9�:��s+�k���;��W厠;�~�A�},�7028x#$ ?O� ���U�,�`Z|M> x�Gv��-�5� >�!'JI����1����F�X����}�R�}QwK��T^��}Ov���_�R
{���O�0�q����()�x�Os��B�����e�Gk�d�,��3�����jbq;C�#1u�[���[#F�g��]�WX��5�\1D��`���U6
NX��6ƼL�A�v���Jq�?��X�O���T���� t���t�a"L�h�+�.�P�L�
��k�W��t\��:����|"���tU�� ��-�^����|U�m$�Z�JY=��G^pJ_�"��b�I�v��M@�{�?}�p���?��G����Y%� �$���%<�iorJ��;�x�N�;�W������t��A|Bd�1��ad�c �I�Z�$U� �m}N���:���J*��G�����n�1���g�(��3��V�b1Z�5
�"�D�����J�����6�m��laV���L!���]���N.��ho:"Ob�K�z�a<��g���(�v��'�%��)x��V��z036��xѾ�T��v֋��/V���4����tz�������\����ag��L�j�e�S;�����[�ǋ��{���y��nvV�[y%eOb2��@j�'+��0�S�QP�b��2������ě��Wy���Wm��?����0�Ke��}�M�������C��O�<�00z�M�4T-S�~ׇ���	��{���C�(���0ή)K�ĺW:('�yE�0�.�<���mQ�1l�JeY|���.�K���w�rt;"5�Է���S^k!�Ab�7�����j˖:'��N�+¶6�,�,>�A�p��<q�MvBICDq�Z��ڱ��7ۑ�u�G��1�*\���Б��JO�!p;\.����:PK�B�yZ�Ǚ��yB�z3%6+����/<q5йq"y)���r{T��͡�H��~�'���G�^���lA.9�M�8VΗ�|Y`)�5�X��X��&��l�*�B7r�p�M��N��'n�B����}G�]��w����D�:3²����24ʄk��.E�CޔĂ�7F3��^'G�� �]�+Pa���+`ߎ�E�v�O��>�I�0G̞w�'5������E�6�*.�hZ����y�'�8ݐw8R�L�H�V�����9���1-���I���X��S��+C?;9(K�.V�
F���F�5�9R�w�"Elll+�1����*�u�`2gnm��Mt�'t��/ձf@n�[���#W��u9
'�ohD� s.-h}g^Y�)�a���>銭����{��~�����ˠ���`4���� S��,��๜�嚘,��Jh"�уo4��&˂�N\�Ѷ��ʝ��R�ss>�/�H�¢c�F2I����!���a���ǌ������5�#�K���Ȕ���B��qAD��Ȋ!L�µ\��_�R�"\(���8��]��h�S7��P����'�i�/���9M�D�gL���u~����N%�sнc<ؾ�M)��"�il�j�J�r�)Zl�K1�i��bOd0n[���7MQ���	�N@���uׅ7��n��?'��"n��uq��[
��-�+�G��xM/Q#��W�d�+���t��l [.}:����Ƥ@��2"�m���W��_�d��F��IE�Sp6G#;�)�Ц�c�*{4Eq�ύ���Zmz)X%2�.�\���w��%X�y����]��DF�ċXXp�M� �w�W�ù�woY(,�Nxr�2}A'��	�rf3���yef,ZQs�+��� ����f�z�bork�z6~v�C�6�[�#�X
�fD)�Y�jbp����l05*�j�e�@a$ M��s9lEC|�O䐧Z!�;Wڎh��Éu�q��z�ָi�����I��ڹ��z�3M[��-�Ǣta�=�ux�"�SMW��<wg8�ǂ�w��A��l��t�^�X�9~K6�:��>��b2�Ǽ��c�|�Lr�����8�$"f�\�D�U���֬2�򀡱<c�B�H������G0����`H}+�h��/��'Ī�$�=���b�ڱS��,��%"��>S	Z��|x�.��D����,߰�|�g�My���g���f�Ҳ��ۼ�E����5��wA����u���;ȅ%��8����_�����X���e����խ�E���Ժz�6!+��;Az�H��a�ȯ�����\���֩~4�+&t���� w��raL��y�qs�0AHO#������Y�J=k���)`81��e��+�G#�v��޶���z��%��>����j�&�n��6QH.�q*��G�|���=����4\�R�����'�y��
pa,}�ؿ/&�q�Y��M�U��\<C�$�A���W	c�.��q&��7L$���������V�h�!�i���l|��gO0�l��T��v"<�� ��r�m�)�w&�r�")Mv�+�@W����@LD��1�K����K�ʡ�n%sPìg`�����=E�ɢ�J�r
��^h�~�_;��^�3mD���V��^�x󳏁0{�Ҿ`�;Vn)d��{��c3�� 2}y�Lؖ,R����]������=2�1�r>��$ҙ���-�s~T��c��ALD*�l'�X�0�(5��Ԯ+owAc�ؿ�l�B�灐N(m���:�Z�;��@]QP��������-Krݐ�w)�[�@����_P�!?GG<����o����Ņ
���@�i��Kt�sS�8 !�M�"��s�O�m�e�����Æ�}�ѓ�a��=
ӓ��VC3�#�ԋN#wPrr�00� �s��,�]�o烶�fX�Ŏd��CgĥXxgM�>�G�}vK��6E�R���9FNp�\uvv1�!`��V�8��)P�7ԩ���}����ZuGBph�2g������sd��a'Gɒ�2����89�i[�¯�nu�Z�2����t!o���o�!����H*��@?%k~sU�
�:�a��4�����45)���k���v24 �Y��ĔsZ�h')�+ƞ�H���6�x� [��s6��"�84#�K�q�k>yDޜHo�����>��[�Eܕ��x�|遶(�w��mm��Y�i�|�p���m��1�m���)�"�VAS�k�)~�ww'��ªf���d.���R�>#�ãiva�U�U�6(�L�Jc��h���ӿJa���G�ud^������MrTV�k��$���o�ߒz}8���q��Ht¤�+e��:\G�5An�N�=�v�$�1\X���"�|� �q��1�/߭�-�D�P&0�s�UX�4�l	�?��"Pa��2��uG"���Kr��{��92O�ɇְ�wXW�?��i D�p>������<U���(GM�6yy5��Ug�`���ͣrq֎x�,�U%Ym��NxJ���<M��� �02�;�qH��U;��� #
�:&(��`k�1�{����iis����N���n��Ν>R*��a'�y��1,XY�!���u��=Y4��/Y,p���3l�	� O�ӵoS� 9�#���Bjr���
�hͦ?������XX¦��U�\&>N���UQ�u�*�RxLw2^q���הVOnfF����=&-��|4���
�X��ԕ��(��/&��Nn����m5uY���E��Ȑb*	��o�� ��gZ�,P?�M�L䍿���µ�[�e!�[=gM,��%L�cX��]iQ_J��(��3��
�7t�k{�����P� y��o�����9��[�>\*��7�cn�����L%�A�3b���>v�0O@f���C�N�_�e�+�uH"�}�Ec��6/��2N�e��b�z*�2�e�1��Z�����g�_�4ו�K�번�tp���u�X�e8e$Bɶ~mI}e7E��i�Pa?�m�ڡ!&���ե�tO��7�Ȟ+_�O߰Dܳ��w(�]�7�R���C�OP��
S��XK�>��͜3�MP�6�B�9�Mv�
i;�;fG&Z��t���֡���C�o�h����6>�%r�>rΟ v���P��u:=�����4��MU��{��Z�
&�f��~	�qM?2#��-]�z� v����81��f��C��Ue���Y��9�$qu��h���`�px�z]�/?�|�;O��z(S"���񜑫���^y^�Ds�F /<x����B�}���S�":��9����m��:l_�`�Q��m��.\)GV�0o~o(u�6�o�߳�t�^�s��S��DY[uS8µZq�Ƭ�7]���I��x]��J� m����G�?�4f�	���Z�
>qRE����4{��+�g�s�����d>����g`bQ�A5�
M�>��b`GY7����r��%d$m};05�4,�۱`�C+���U�� 5�մ1/�j(c��d×�l>(yHz���L�܁�(�Z�Jj�T.{f�ULUZ;�Ȥ������;>R����;�az͸:˨��]��paJu�_����KgI���Eq����N�8%T�! �,��rGJ � �ug��ŜP��o�]���"�Y�a7�@u���O�:��&]�x4�m2v;��{pm�F��RI,<�z�ط@�^�ń��S��*�J5| �zY���m�5pp!�֯rg$6X��Ru9�g��&���N�:iʱ����x���q���Ė4��μ�w�@K53��9�h����J�G��]�n��Rr��BWhU�9���ޙe0/ާG�����L{O��-	���TM<@��q������f��ZP<)��Ɩz��b4=!q8��`���8&c�:Q��i���-�� *�f�z���^�Y!��0SH6i�2@Ik�����Y0z��6�QJT�k"�	�ӌ�O ��x�v���8M����D�[�e,��_�\Kǈ�˸Wp����A�&"���*��$c��ui�؉�n� 4޿n�����K�"�E�����7`08R4E����V���R
�Y�kdT}J���#x�>�dģ9Q� $1q_sh7x�h�䜲�u�j2т"2뙆/�g*��/��Um��-��w�g{r4Cp��"�+�+�m�
id��"1)R����`��^���"�q������ի+�Pa	���(��6�ɫ}�����at����3�S�8��dC�vNh�6��`-b��ޚ��OH3c�����:�{4=ڲ	�o�ޣ캸�M�� �@P=h�x��zy�,�MI��¡�߈Yx��݁\Ѻ�ʊ{�%|�?b�ٟYp�ʪ%q7�w��Y7<f�M����ث�IaL��*��.Q��/�*�d�<,�8-v2螁�4��7������7U/��k�'�R�:Z���td�f2j��h���bƔ�$�����g�;ͽ�r���9�|Z�g�r�=u�G�
H��ة����rYNV�b����Q/=�dƀD������ ��
mfc\�e�]V�5}+ �s��[s����a���Jd��c�����EĒ2�ԭ���
�M3ꁖ��t�����;��,ѱ���h'�9sRU�/�D�%��3��?���H�[�.Od������������6Ӏ�L܏��wܖ�n�*����R(y�+n'��H��9�h�U��y��c����� �����/�I4�h�6�IV��z��`F���+�Q��oS^~\����v��&>!.8���n����"돜GJҦؑ+����;1�|�,)�M5t4��Gj��o�Y8K�	C������>����H*�<]��	H�sċ?��4Y8����8Z$�Z�~�g�<��-�&t���`���`�)�)��#׎��HC[�&d)D�S��\�@f�D����2��qlg1E�Vu�tFj�u�n(�B��y�J=�@����T?\�����x��e���X<Rut�x�%�$�'�S���g���n�V���S�����we�1g�K�7�tA3���#�LF�Ӎ�ۤ���F�pgX�zpK>�k[j��qW��2���u��'0�O�;~h6�
�s��K�N��F���C�o��(s ��v�H����
�����������s3+����C����~}�l��[��\���ۖ�	��h��\j\7m�	Q�#d����y�S�^����?�ӡ��	���$����3��QH��h*�Вa/~z+�L��U� ^����N�������&i�e4tW��w_^�b� i��<�0�
M�5�!��RU��~Xd)�^V�b>������������2;EFESb-ؤp ����?6���?���L~����!<�#�~��A8��ɲ$M��>2�+X���T�%����2G��~��h�A�fv*W�H�qF�v#Iܧg����M�u.�P���a�6�[yɚMx�4�0}��.���GJ����;�T.�@�8�eh43߯�{hl4i�i����XP�XsѸ����|���{�0ԑ�@x-��7՛�e?p�}�(ns��cD9�`[���^՞��` �'@(T��@65�ACb.�L74�+��b��?+�=��9���΢a��K���$8� ���[��Yv��=۱�������~�����[>;��j
��z��	�ox�E$d{8
To#��Ag3���_C��Z�^/٫�)UW��@F�r����1 =-;O�^?���r�p�T#g8" P�[�x���>EB@1�p��[��q�]SHZ���ztZ������,�Jf�����3����5_��B�!)�5V�$�a���?��~�
DI!S�� ����Y��.���'��,U�A<ؖ)�m*��{C[���*	.g(^}�?�{��?k(Wx[;������ٹ[�_�!��Mo���! H��Qf�SDӞ��N+�X9m����}�G��	��5�sѡo]f�m� ��d�P���ti����
h�$��Njy#< r���g�'�¿����2��i���dl|�u�x�{���=������N����|&�K�E5��؄'t �*
u}�$b�	�g�'��}9z�INg�$���.��cS����Tle��̅/\?WoW�2w���^�}j�G�����3���xO�y�O�{�=�]��`o�B���8E��~HQ��H���L���I�7��Z�<����_OPuv^í�Ru5&�N=)jq���a�h,cES_{qC4��!�[��A���]��[QV�����/���S�@1;��LB���H���=���+�����6ػ��$���S�&�"(^�|�h�����.�H���d�Ak)��	+�W�y�p��Y�ْ�?0<g�9�uS�庳�\�2�2��X;H�KR���.
��8������d���w�m��;�B 8·�.��G�^���!h
2zr��:�3�2��>G+,*�,���םV�O�j�\�Y���m��9w��{|����r���p�T|c	@���*3����
"-�^|���F�!��#�(���l@��Q��8�a~	Q�b�O�ZcN�nՈ��S�{���q�rPNS�ˎ�h�=�%�����HAl/<� t{�ԩ���wq�#��V��4���Ƿ��Ğ�:f���ty�D%@Y�f�£�����bF�Ā~�^���Ѧ��Z%H1்ڟ�x�1�z��뛽L��/����J9'�dl�9-�T��i4�h/�.�/|c�����p鶠#~L��]h�����=k@��ƫ�.��pߧ�Wnh�Ӱ���vd�=��$|������R	��Se�O�r�q�7	� ���8�w���8~��U�,DqX�"ֻ���3��.�
.��d~��%w��&��8ʎ���1C>�&�^b�S�=��U&�3!��r�b����@�d��'h3����QEkh��!��[�"*m��"S��[�������������?� !CdON��`?)�a��]-��I_A��_f_����2K�Tg6+�=�9�����ż��Q�ͦ�	�q���u6���ge񛤉��Y����P��'�W��rۛ�M�2��MskFc#Q�}��̧塱�qߓXr��u�k05?��9���I�m4��ez���e�O�� σ� �v�z�1	W.tC㧌�_�㣺�'d���|rW��0\]
�q^>@C[�"�-ε��@�Z���s|F�ꑵ
�K�J���H=��_�7�-2�{Y��=V��+0Յp�E�e;c���&,
��℁q- �ᗙ:r���6��_�cQ�N=�j�[�Qf�dFu!�@����:�7�z������!b����ce�\����mX��YN>�♋/ v��p.��r(�铅��o��rf�������`�r[*(�̕A=i�4�W�������l3������6�<��3�o=��Fd^��7�4����^��_���fd�t�?���[�;���4�)����~��܆2�j�R�c�!�g"t�%Y��HڕO�H�w��uh]]��Ij�����C;��jBs�qD�:.�f"�A�μ��!�;��m��Cm���Z8E<�c�7�+^Y<U6�`�1N��UuY)��'<	�yr�i��ţ�V1L���y4Q��Ft�&���@S�j�ݜ�C�i܆��������zCW������\�٘�1�;W^a�k�Y��|'�����bR�y	�)�hL��޶����ҡx&G5a�zS0\}�4K65�\4(/
��7�.G�5(�
�%Pg�*�h�h�,j��T�VI$���_O���^�t"���/���ɩ�TV����͞߾�Y$�wX����`<��d����#����Ș����O*b���J	�o�>*���$�*;ϟ|�J�xr�%ƍq��j�������[��U)	�Sd�=�=��g����0we)��K_A�d���e��@(#_�װ��knj���"Lqm���]�[
��[�W�d��&���2�����������n����CC�h ?��/0'9y|���j�y�(ݬ���mӃ�/��_�D9>�V@_��x�G�$��[G��^Γ$&$��"�X�G&�4�c��uN���?���@�B9a�l�L���-�Z\�3s6��3���$=.VrS����C��_e߼/�ütc+���"�yVs�&�~h��9��%�
���,��~a	Э�DK)j1?a{�|��^0�^@�E�"K܌f�#GB��uq&E��M�p���$�I>	��_#8�GI�[;A7ZIl6ٜ#�;��H��5/�	��f7(�)�O��%�2&�뛋n�2��v��J��o#+�Wѧ!��=��G0+K��%ژ�:�1��
���.Vȗ�e`��u�����0��!�N;��(�J���N�����km� �S1-���?dJ[�u6�'��D+�X�1<��%���rѮ+'��RX,@`�dEV2E��߫_��s��i�����/��[��.r)� :�K|�1+`�y�
�Vֻ�b�TA
�KD�=�`fn���!v������m:�^�)�U�l��n�w�d�?��n���Hv�L[!ئbR��5����%dUn	�ɂA�T!8���^e�*p���A�r*A�7,
��]c��X���a��<!�}��~������xvYa@��ι0�����9/�s���"ݗ�ar�>mv��O`-���I�7�#�]ӿ
�o�/e���u�DeI��!�Ҵ�P4�����-g}�1,Υ��(���Ў~'�����_8(c#�&;q���z�b�	�ӎ@���0���oXj#MWyϥ��>!K�d�Xr#9�ia���w�pTT]C������^���'d��uQ��w��"W@�@9��!�h���^kV3�b�=�y�������4p�8�����4\��K�~D�i��y���w���s;C�U9�pv+�8a�������4B�"�ݟ��ێC^�Z,��b��k�c�Շ�=fx�
�;�7j3�d�Q�Q'�eij�Ԉ��TJa똭���Ըm]�򯽟���V8,p�����qG9��R�;M�8�R�Hz5ч��[�qEv�����+�DC��7i��,�c@��alUgɮmte�]��j�M�)s���v�B������� �&��ՑrA�!�f�ӵ���df�%��R0QOY�s��&|��Ci�� ��X#И�/M�PR���T*$<J�����4�谞�a�=!k?�
����&��Z��,����x�Y���.8�U2�?��HT:(3B�˵}��[t��M��ܥ�u�0���W ~,'˾j�Y�0�7UMG�~�5���|Vk.?r�kv��ݶ`�R-�ߓ��Q�I�t�{,�UO��Y�&�����Flx);� �W��>�ΊA�܏�}��Lq�p8�en������;�?l�$	�uq%�	��(����Ok�n��"_-iDt������c��>�
�&?u�I+֑��9d4-�>�e1�Zn:e�N~�^U�q�j���G�Ř?-���B�T���߈���"��V3*��3K3#�]O`l(�������#f�D5��tU\�l�h���z��l��̒4��c: y{v�l^��T6���I�[T�hȵ8��ϻW�uMZ�\^u?|\�ig3�	�;\N4d�����/�Q�6���S8�E��'�w�Q&���]!��W>I6�m����^.:�J�V��9iZ���N�]i[_����S�L三���1���$r~9FԺ��gY�%C���P�����f
Y�V�����p�R��󀐠�<$re�s��C���1'h_��M-_�#\�:=�u��L`��l��aA�?�X�*9A��p��e�h��L!��C�Z�AWj�z�O�q�>�8��|��v�a������{(>6�&�R���+һ8յE�hr���,�{�����s��E����r�.�ݭW�/�b��Tvz�W��&��ddw*�y�4�S��O��F#]g�4Q����n;��ڍ�o(e��I|��v�$�tB<�u�u���eYq�ż�PpRY�X#�ro���.�l��ҳ����U��林��>7`=���`��Ԁ�������_R�kN��5��-Zl�f�r"��0��0N^;yvq	���	*R�=��\X��x��c�U�^@�>F��&�K߲:��ىZ~�zʒBE�YW11��!�,
�o�u7����7\~3zL��8��n���o�5}A�G�SX�m#*���7�}��}(��$�+4#�X��m��E $�<��CiƢ��A���R����@;�q�Q="��@rL
J{�Xm��\1a��~��K�I�R2?�`%�H�*��1=#�j	�+���p�jxF\C���4eo��ڧ-��@�yJ�+۽!�������(ؽ �+W�Q~Nt.�?ܞ��/��7�l��|h�:��a����I�SSHB+��4%>u� �n��É�~a!Im�]���l�t�-���b�
bnt�[��Y�ֱ"%m�:�p�[��/b���2Π0�0-��mrmY��\�l��?+'xX3Ic����Ԃ���m�4`]H�6�v5S���i���"�~a� �;ͯ��"� R�,�E3�<�����ϕ8�{ ��4�u��͹[��u����e�ٖfbcVDK����Y52�d3�JD��`�#�`Xi=x'���'�j܆�s9T1a��
ez�����d��J�7=���̀k�J���icc��u1as��|�D�~�[�?��^߂wOt���H���8����"���g`(��y_�ډ^(2uvݢ=o(��EO��H�^�d��B�(dHpg{D��V!�Dc�O�k#H�=d���7��;��������`]Ĺ�L�6q�@)�B�}V�R���M4/ܳ�*��p�Z���o��"�1�T�=���X�E��+�
��(Ǌ�$¿�q7H ���k�)�B�N�%�`�H����!v���ܧ��:֭^J*y3��a������C$��.�ȯ Qe���J����_����)���"�i*}����������
� �uW��4�%�	��1:ze�^zΜ"ch�7�\��I�O��(G;o���Q��T��31�%L��X`߬��˔Gx?�̈Ԓw�dI}�+�A�*�v��N� ���u�}B�B��4����R�H�����߮i�k~1���^���Ww���K]�]�V\������\-�x��x
7HW4�P��u G��J�jY���F<�|J���Xܲi�a�9b@���G��d����F���0�t��k����15PXb�3��ON��Q'�;k�i�gy՝����]�MNF���ď؟����O~�6����ʀ01Ȅ�$_���[��^��~��w�
+5l
�FȄ���p}0/�P�3�y���
������ى�@ȳd#��ߠ����S�A5'�љ��cJ���$ c�t$/J����#$�z�W�x�C��0u����a��4S��r�$�w@�;/QrR'ԸB��)��<S�\��N���0c�p`�
L���l�`.;o�R��B?4���2�LWov63�$����˔��j$o\d&�Jq~�%"T�G���}��C��a&�	1�c�3�V<^�O+�`0a<
+EAPay���̑��W���q���7����,�d��_�����M���Da���=�C,yr��(�������$J����8qR�Z�T,5뉆+7ɟ~���r,x:`Z]y��=���+O��yL���"���3�-�5Z&��~�6�egB����v�A=Q��}b�w$��@�(D��],� 
�l�?	���yo��T�z�n�p�5���)k^�_�~5�#թ1�ñL���Q4G���&5�&�5 븊wu#�,��� ��AA�/��UV//�Nc�sM �XW�vxe���	��l�t�Ț���9Ͳ<BTٙ4��ٺ��Ğa�����W�I1��:�
���&�l�S��@����&L�:2L�F�nOT�����Gֆ���ͦ�-����B�AE����c�9L(oP�������tXF����X��U�.���΄H8���~ ��g��)�3z�ר��{���+s-�O;S
mf�?Y��u��4g�A�{�]��*^	i,�E�^�R9��V���-�-c|M�� %fPվ��ء�18$�i�m5�ՙ/ݵT>�燖n�̗h~�?E.&��lC����>�dh����E���ޓBP��������A���f��&��P��kqCqz�� ��)���cAB�2�eD�15�56L4�0C�{�gP��`˵w���RPz�I�5��C��$����(yԃ$�݂��<8�py�#�矾��e���ȥ0| �(�����-�2z�2���{�Q���t?��Q۟MmI���
);z<r��A�$�K�.���
����s���R�.d{G����G��*}�����U}x��K���_�T��o��B�W�����w�J'6Z��}�� �M���9�Tĭg�5Dpw�h��[ؽ�ېAQ�z-�Q˯��t�>{�������Eq�,�A��i����fR����2x���$�Q��By�Y��8n
=����El���Յ�-�V���!&)5��m �֫Չ|j7e�RN۞a
�H�܎;�����Ѕ�tPG'KIpz�:��a����`3�HF��P�ؑ?M��P��}W=���B�w��_ ���w�NG�l��t*K/A�^ 3 t&����,/��mҷ��uuJ���c*qô�i���j�[">4A�u�Hݛ����o�8�Q?����?��9O�O���0ˡ;o��ٯג���XwX�`�CK8hd#N���J�t���6�Kc�E�S�Ώ9Q�aHw�֎��,Kj�[��SO7�g��*}�QYHo��+XCH�����0Ⱦ��<�����`w��3Lt�J�[~��]/���^�|"�29��D��ɥ��+�+�����V��@�Ϙt�M�b��	�
.ח��� 8R��q^d�S�l"7��3�;�37J��\�Zb!��4��`P�\��E	��?�� �_)!����J�>S�&Ӕ�)j�!̶-W�<[��V%���A����֚m�l��F���4��38D0
�ra���5˼#Y٥�~!%�$��hS����A�Lƅ �!��iJM�� !8,��n^�t3\�״,���Й�&p~�T��(`[j��?��K�˥� �h�u�֝�C� xc�]J��q���7���H�VY��I)ܥBq�@����J�W/x�?��'�y0�c6�R\T�=?�i���M�^C��l:5y`r7/Ă}�;�]��~%�0Ҏ:{��g�Z��N�I&V���ԴH��'��������^*����P��媿[}����gʥ��ּ�A՝�(���Z^@����V7���9����6 ɏCP*��Ib�>�)1"�mFpL����͐>��R�ē��8�	�A:'.]A�^�U�B��TK�3������.>H�W�֩�g��sWA�x.C=�Xx]��?%�xJp�}5�����3'�U&=��-�%�&��z�!�$]t�܊�� cR��V�-B���&��^��`H�{�A��o�F�pB%˅+o���W%-�4{�U/<���ʔl�vQ�s
ڛ���v������Ez�Pb&�9~���b���fg�6��)�12�7k0	u%3S�����o�!���Sӡ>ʲ����9�7(�S*�o�xQmI���*k5�,�A�UFjG�|����.o60Rq�о9h��oͶ��`��_w���kq�剮#�ь�Γ��L���/�)��D�������s��?�3�L��緲�筨�Ȼ�/
%/ZɶY���X� ��W܅̋Qo>i�@�����>���5�Y�0��U����JH���}���gM�}a�ݘX�Q�i9��v��/�>����C��������V�~T��n`{x^f�=�r��b�P�GA�&�(����`�pSв�w��Ͳא$E7�$=����2+-���1T���Ƕ�4m7,$C�U��m�OpĜ�A6�� Cs��1z�E�ʾ�=+��7&{�{
�^�ݶW����\�YX:�jB�C��2ߴ�k�+��q=�2'� ?	�\Y͓�L��R�� �� Pe�RIӊNB���#(�u:��C���z~�C-4:�[c�Y�;S9��(��a����a����L�n��c"ם�O0����A��i��!�w�q�o��^uH�N9����&��xH�_�A��4���{a��b.��o�H����!�fVe ��|A."�vR3b�v���D=�YY�_$S�G�A���Q�K���{\C�![i�߯�=��vb�=XwG��R�r��G�+��JY{A��.�e��X�D
��+����BO8/��E�R�Q����*'U��+����%p��;�Փ�w�� ��x���֕@Ca�,�5�"W˧�S̹;ր 3���8����tM׆7�\�50�6+-O�1E3OZ�O�����&«T�HZ�{�T���A��fCE�rf?�2]I'���Hb>�:S����p�������`�n+(�+d�eVb �dKJ��%���G;�ei���Z:M�
�W����_��'X>��V�.�7���/3���D�a�Lc ��J-AS�p a�e��m)�΅�G�,gY���f��Q��#E=CL*���6E�9����X_ŲN"�5���X?�ss�җ^�,�]*LN~J=56����ㅩϛ�S���q�ۣLX�1�,.ߵ�;�u��4�Zg�p3��΁�A�v� �
��(���X>���a��p����^?|J#�&�"kk�Zi�M�6��Q���e��h"}у���;>_A7��ᴿ��e�a�r�4�E6ɕ��·{�U:&Pр�R�!��<��$9\R#�KRz��t����z���$�E����-m��qX��C�S �}��U���Ho��� (q���;��G�@�=W�N�2�ؒF�����O��2[��/= 81ł���3>pG:F���4�B"�MkԜ3Cp�zxO��
H�,p�}�G]!����d%�j�s���C�����KX|Ճ_����c�6���Dޣ���`�@�b_�7��|�9�[���<�*�E�[��ZG�o��7��F�C�` A��,�q��Q�7��B�*�Y���L�Ⱥ];F>ha�],:�`H���?�(*��6|��"�ڬB<�AY�<Wj�2��s��\3�����撮����9�y����o��GU�� 	��7�bb����oG>j�c9]���glT����cx0��	�u(1 K�4=�v�m�vS��`*�C�vv�};K��`���l<'�I'��s.iwN)�z�!�S!�a����tm:�-�x�.�]���Qk:��"q���7ڕa�����	�Jk����c/�+
�f��Z����_b�� a���VP3��K�>�cC%��S���A��p)y=�:2��[-�L �����R�^a�_n2�����������!k|�G��'�Q�Y��5u��O����*{��,�k:�a[V}F�ő8}%ա�.�������-㊋�v�O�Q*q��\sS"
E�ʶ�7<�B�*߯XP�n��
X��}���gs�;7@f<2�f3��+^cӝ�nȯF'&!�Qf x��zC�mT3M�g4�k͕H]=�'��3)�d�SA(��p��d�o�b���t����>�D�+L�C1!�;N��4G�sl�i@�<5wZ<���N��\S%*�2����x�@����1��"�Q=_�-��}�&��.���+���p��k@ y����<|,�q@(��G��X��:幬��-�d����.�C��c�Ur`�Y��a�^О0�T�CY�3�9�॒/w���ƹ�cz�_F$�v8-�ꆘ�%
u\+0�8*F���f��T3鰇u���]tN�����X�n�Q�[�xo�B�=���b�`.�{c�����KS� �i�;�gvh9�Qr��P2��[V)5n��[��Ek�(����я�}�.���~�G�g ��f��_m��;T���Z	e��2G�@�p�H��ư��
���Ka�&���Ӯ�_���י��U��]�ɟ�E� �ȚUJs�8�ltA�|I(��!R~<X�������+�K3 vW}E��+"`H���j�>�W����\�o�
d !�ᄱ��٥)��k�ۭ��%�����.����ڧpҿ��<Y#�Q���ç�c� H:ke�m�~��"ʿQ�iP��K\�>�jD����
�#������g̒�L�Ut����*�:{o���3I�N@8h�>�-ԇ�M(a|��(`19j�6��L��ٗ4D3դ�LP��o6T.�:�SM6��R�՗��O�	��� ��p�ʽ-���� Ց��Z���%ނ��̬��]y���Z�I8%�ɩk[|��\mJ�0C��X�}U�Bj�6-?фjx�:k��f��H�C�+��0���ϯ�~���̈́x��Z�6��V>�[d�v��L�n�c��h"L~�=Q���?	-%老�>��7�����H�"�����qD^��%��j���e�A
��7qvs��o��3z�ٸ&[�e�䋤�e��G����w�/#*q/P]*������R�&pH'Ix�>���)�.��C����*��� Gjɱ�
9�Z���)��y��W���"<AF�A��
��&�%7d�Sԏ`2��ݯ�i��@Za�G>�;�������&�[d�X�Q�w܃�`D�^�O?��0n���Rѯ��8:b_�C��  �A��ቂ���2����*w,��hrc5�O�+�19��%�&���H��j�_�R���oÔĊ�@��̈6�uy(P�a�������K���	�{��ϯƴ[�1X�*ȰN�y���@�~���}��c~a�4pS�V:�ܭi?� `�]E�V*�A�u��x��� 1fY��<tz���rx��8 �7��9���Tum�1%�V|r��`��9ma�"��E%huq��Lfc<C ޠ�^�+e_&E�W��4{�F<��\�P0���x_�"J�#k��Z��{���;7���O:����?M:��ؤM֑/��#������;G{�i�e�#�_tL��◲X���n�f�_����qDU�2�~��z��\{�C��I�J�)O���\��Wl�H3f�@��!�s�/��Z� !X��tY�͞$m촓n��Z��̗��D9�����Xǥ��쬻�bJ�� oj�Ia��Rx�k`I���5|���YM�C%��3]��
6���:[�*������=a#ʠR=�Rl�""��Š�ض�沞�>������M"��=��Ԅk ]Z���O�<���#�@�.n9&l��=m�y��+��J��������_��:]�X��z�����/��_&�aͭ����(�y7L<M�j���r�) �ttR&��.��rz?�o�:ɢ�d��;5?wJ&󛢼Xv,M9|��G��tw����`~!ܦ�j+��5�t�_��T{��*��.�/����Gj������K��mA,�4H��>}OPO�!9�P��3�C���38�8��5���I�P\���-y^�4����q��޲�����nf�6���Z�5c������$�^*���G�����S�{b �k`�if�W��",}z���,�q���?�����g��r�5�<��y徙"k@�����^�9۠Ӹ29��ҩ�HY&>�H!	��P0Hiʗ#�0�n�� ,1�f��)�<x�Z�^�^�Uxv����gJ�w$ t!�S~^Rqc~��ۓ,�"��_������z�̙����Ru�A>{%���΋��!�@঑?;:�gP�0�z���+��%�0��,�{<}�{X���D`[�C2��	g���p��W��a����H�ס�l#.�n�� �_��-~ӭ���Y�����4欂���d^ �_�Q�V�h
��)�A��%�o�_L�/�7mo�Ǻ�;��� ��D�"���\w�ؾ^h�	�s]�����^��k9m����GsU��-�s0���+�> sk�X��
�o`v�d��z�)��q�ܦ�W�B��h��^��i��$���K�k���xq�V�"3?� ̭C~ѕ�1��.��� �;���N�F�2�CCI�J���T�pkU{9z�ѳ4]c�Gx��D���N��,�ێ�{��zR�Р�դzM�Q����NCr��h:�( ,b�+�#]�0�ܑ��F�j�d�#e��G��q?	ք�p�r�C�v�h�kE#�kɐ&ʱ���B�B�`����u��N� ��l��=��SU�D�w��b'�C	j�������|���}�3Ov�Š�2+�]�����)��}�A�Ȏd��"x�~�S��r���g��k2�/$�i���E@ZQ���7�}��A��/���Y�(LS��w�㸐{ץe@��D��O)>��Ѝ��)��"�.B	Z�},�(f�����E6�뮚�5RR��聞L���>}E]x2�Y�N%��}�>p�� �0K�����N{66z�d��"�,��G%�p	��Ȗ�B��*_�_@Qa�kr�P���5J��>0N�Z�����a�9�Ӕ	�[n�m��<U�-�M�Ĩ2�"��Nڙ�ZXϽ�[��H\�}�3�HK�5����COk[4W����rqZ��߈��0p�Ѐ���VA��+C��cO�1]� y���W�C��K�����M�ġr��;����O�˰xӊ<{�mǷ;���p��f[��F��!�E��5e��Wa�	�"[ �ܖj�S���o�C���y��-u+��r2?گw�l�ܜb��TE�Gn�?�nS(}Q�2�0�}�ݦ�+N0k��1d6�+����u�͢Ѱ8�^����؈��0���1���z Fq����[�>kp���%iMi���9=��*�;�-���ƴF�2�;6z�tD�F��nuذ"N�_��џ�n�8��C0��$e�t��"T�:�}���k��x�'�e�2'f
�ӠN[v����M:ZJ�2���