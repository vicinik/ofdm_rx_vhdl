-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0Lce7Jz9r4HspifQjkLqUz69dbqdH7Ap+jasz+DHaFTXBK9N5EArxrigR4YreN3f9W5IHIIgfiQJ
gVQICimxOT40AwLlnli5LddNeFQnGhwuhGGfnxb8q6SrGzauqqv1+l/sUahHO1aCEwcsz/2/6C+5
LPxIaKrDcX5gYoKETxZ8Sdta7BrNNz1CGsWoOPilyYq5FElNDbFQ1Jz+CY4OF+vhAoirDWZuLapM
XuyXwsZDlHlA3fndMPXcLPURQ1dUG+ZzbmsYa48mdU4l/VGxmyNj33p9balH4mXEsw6bsZn+Gx77
hDg3KPmDHKbAaUcdf+d6WA1z8ngc5lyjFksvew==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
xPXaQWNkszN+67oPkYSS365VYmekzZGdpASnnsEnoIvsZfdC/bsudQ/IYco4dK8Rbu7Rf5/8C1cT
7mr6qCKRkXprlUs2zqLrboKnNYi/mqCYhtPyhw8JkOOxhH7asp+LbnK5N6AQXyAPc+bKNCH8QaWN
2vwKj1En69z/NrDIw2JmnCUcgbUKvPJOEuNCjyw4PM7yCeXBwsQIipaS2XTg9UqopV3aAgm8fZXc
Hq3gJfG560+CG3qkuvI5FRAjMHxacJ86RdQDJ4YAoN+ZQ+zh8a4Q7Xadp4rsBVgoDv2kYx10rxOc
ynM2MMQltDfJVfaybNrBSHrnCUVxm/kkxseCIWLXaIn2f5oZAzzZ+aS8li7NYFqn0+Eg9DoBu4Wf
s5EhKr7S8uQbejZAFK5ubz91OXmNQxwzjHzCOiSBYmvfjBHj30sfQXKniZV5xC9tJo12auH32FBO
W6260/0zoMtPrVU1J47vo2FI3+axLPKc/6ICvaFb/Bs7fXIcnCAEAs4dsiidv6TOUSqb7vl/6H1c
f8NuoCHcAY7lrjb5mD5/3hcdeBBiopQjYHnuTfdkBtHETk54Kz6oj/weDnQTTu6XVujRz2vIOmEI
Hc6TkSPLxB6KvKzStZzxOvN3Wh3k7M4irecf1SwgDhLCAf8bDXgC8VAkL8FDDOEYhmQ1/0ltaa6j
PzRuW54Yr/mI0oOyYAb5GEcEFuQ3T6+YLtKrag/DhQfp19AmKoTbpMUyVDhUZeLv9ROuwJnY7TKu
l48ab160ws9Rbp5fUgVKfrXeXDBiJZam/Mt+WMvA87vCrN3Vy7MxeaUW9LwnvFDHTIPPa0HWmLoM
Jo+D3i9avhoMDhmMdvk5id1LCJZHM49hi2JKPoXTu5XpDmrxxp2zAIuugyDe2xibYfYpFk4rf0HQ
mwrdR32Bl/OOzFOrGLEFu6j6jdKGNg3iufwyJsg7U8QDk54nrYexqRPVNQ1tfHkmIrjTPme29ecj
dtLKGphYAZbYxJ3+f7Ez/GyAXE/EsBBnHgou5je3Gh2dgHTBywEsbS3HlVdq/ElK/7IKbIhwywPy
ihByMAZzlER7VFHq/T6WChipFCSbcIXqVBnxDft56dRq0WB+5/Ymtq5MKzpha21iURP2zLUUa6Yc
3eesitwoQsj++KkUkYUQLr7aB9nVnArbiUAqc70VckfcOGyFcZhwAP8nZZLV/TrNkWsEohXt/o10
K5dXtwHajpWOv23xD9giFeDa21qH/h/5KcOHoQx1Hf2WpXdNSsI58umfnvIerVEy+pB0sLFTOkce
sfcmq2JbOlk+3S+T4YEmpfDOHo3k/9uJzwJ/h0dJ8glF29hNnl9ntUVKz80HJlBQPHcjTI1sdQ4c
1ztKksexW9x08r6kVdywGgtzBMc1NCF4XWDbp9cdSXRvQE0LAJyoLjjT72m5nsI1a4Kz2I7nCu1T
XEhbaWZAaD7s2rfF9jzuz9OuJufaQ1LxEyxH9BLakLmBZP7/IUZhldU1IVS3G7iVIiv7mSXYpZPr
RqnJGnlK6Tq52VwUt7tS/EGS1KGn0yk1uQl3Fxw0HFVotEKScWrpohRK+unwSCz9G6Co0OKhlo13
ayful2+fpzh/HiePCY3VaagEDFgh2cNUTMPT+n5JwJdyjHan3u1uvg4ybMBhmAMO4ZaNdqEKrt0+
/6+ELNAyU4svVZq0h1P0kVoYSg5FjWihXWd7s7oJ390kJV0HQ4+vFu+UOKnRTl2HjRKbcGhJ2ZY3
Ddq8taXpEvsEiMNuf5phswSM4lQDVSG4lxeEnkE595p0zLjh5EXgCgQgme4ugDoMjKVa0vXtH+Gs
PuT4eEgZ9syJM4TrU0EAyWoarEaLgOAIdBxrz2XW9Z+zM4Coc278ybEgXNxA3B1jPzx2NF+c/Zgn
37g+4tA3XnUc5iyDEyXYNBbLrTJSXMrEkm0qwCxTXvBMv5AifxTDK237psSQApALqveBgTYxlcWx
+hfGwvF8TlqE23U7M3LZiE8dNfZGxPuV0zABrV+AVKufeEliYugPbMcAL5PeN4tE4+RX7kungZjI
bSBY9pOUQn8484adObLn8bXnDUtdV2eKvQLEw/IpGM6bSN1oDNbJuZCc254tob4jxzjglA5Ce63a
p6dA00fQLoxBqN8KNC74s+wtUPgVV+UOfk4KyrdEusuMEqnI6RhDpMZAnTZoY0P+odj+Yx+6KIMG
eNLHm5yw4VooemIG5l20CAJUDGIB+4gAhfd6NM9mjC9QQPF1CTD3c7OmwT7ohiAAadfldoX1bHtA
Eye7ecFpSih0KJJHFvBhOejWIl2LWt/QtpxJIbMMaXQPKNOQ2rAvIOvw3B5CIauDS/DEEuffVXW3
dNiEGQbzYKA+Xfi3tIm/juhKfU6YxF9VJdSwEb35mSNvDPdd7Yl9pCZ/ykllwJSJXp+E9C9qVjcc
WiQ++kj8Od3JiBvUVxSCMY9zmXwNTAr1AsfdhXAPHCKFGbkdN/sDBvQaMEny30fWe4VWvrhjNcAS
1pTwu/L+aQCYWmQFD+gzeX0uCYc7lm5b9wNmnIALWgI+Ut10x4lzlPjBBCEwi05yc7bEjtQI6noS
yhqC2+9x7B8336DBAkqx1QNJlLxq05QyyXhJQSZg/z6GFwONkpNP7VHgoytHht54AiKZPgtRyWlp
3wflAjo1rozVhj0JEHhKNjx0PS0k6j0k308YAx7pMDTvy0jOu0je8JLU69gDYBaGsCFwSMGyoqU1
x4CRmby07ZvjKyrjcrW65AkuqPKLqVScWXaGIqyXjaqq42k+welolWzcSbosKFraJbenSSKpaMCh
XO2RqM5Et68N2kiV3J1bpOv9jOEPCnpeSoP/H3P8/jsMx+kWcfmVI9ue442UckDj8sybqKwq1Xh6
k1qIf/i/c/BVkgvMgUO3TsAz5P70YwA9gd/Nu/fI/L5OR/DP5aaxhcYgaPfG7SM3BKEWKGqoKrs0
0EgDNqMTWW5yidfZkktdPEVC9VyZqAiQte+ncFpYxNn5v+8ZPRzyMlmhG1+71GiMJrJcluFqJujd
Wn+e2pFjR5CwA5s7Gc+7bHyCzMI1MFIDU3Py1tjrU8D4dIIVv3mPkSQm0eonei2xCdjxRJUzR0Le
8CiRU+CKNF8TrXc6w4osaBZQ1YbjrNVDn9GXs/YpjkwNPM/Wb3svBL5A8kF6+UNwpT0SodUmFhTX
Q/MnP3M2ZQBVY2bXDTtoKKbfWoDnsjLaejKT9y9OzTd/11377fJBoM+oN50BBw4tOcyLoPLPS11j
M64K318G2WXEy0DZKCHmp3UtsMbnMjzaeL60cN8BMM+JYjGYcDQNkpMuER2iymKDVfp8304h8v+8
PMxzGyZg2AreLHscn13jCFce6iIsJmYpHxCbpoDrYcIXuKXeGf9FahALiWHszHpq5pSSowRWkHBg
qsgl5uNyUNy8wDo82G3G5VQ6SgAHY6XE3WVNHr8JfSt/Ou3I7XEkEwIwcxPZj5pNyZhQqbvEtDFS
2PElJeMBO8t9dz3SykWrdNe0P+vxEyKXyYiEVo1jidvyumfIQii4RJf+yfaq3X8GqkFxmKULZnf6
8SXyKe7AvFI8MLqklggdP3ZQW+qLg0Vf3I0chcWXfu7kTjypA4LT+uOydwRX9XVUJM5JK265MinT
pchjxnHP8d9PnHiLMkbpRpZWpiYmf1gUHnAKmTsZYrtrUF6FBn3isu2+Dy0/nyKr8rX+ZASb+thw
DIMc4JEjHjp5iI0lgmZWLtloa7yDBBHaVVUuVQm3D3iP2kDpJEsv1tzmOMzDTkA6TfpO1eZmGsC/
If8yaLTUmYSxNuWVMuPNzwe6oGp19E8UXfivV7/VPcp5Q5IfZHlyf2dEZp1GhqNPDlijm4KX42xl
+aWiw3NswyDhLNZjlHY9/4HODnDaoRemHfDv+xVHB97ri4V+zo19ctrrDDs5ukJd8croYAecr1o7
ckVVrxPJc92IjVg9lkbhNkJRQusA/yVHXtBUptEu9s2Ayamp0tuApg94cgy5NUBobHVOCkJLTzUT
di6cIr4DOd62u9lGBwn0lA8Y/WqBbEpQ/VQLK6AVYObOjM10EEt01DcXUngEdc7BCLQU5aOCaP8P
8P1t+Ck7k56rRq1Gsf/Hsvj/Hd14gS2KLQEuAZgcVS66KZsTx2iP8IssexuOfKGBjB2VkZuEECbK
dtzJscKPQFozad3fXtTsX3jh2sD2hXzIPKpbQ7G0ZMHz5bAgwkCqlhgwnxZO/F0xaQA3s0YwKVmB
tzCy4oAcBJpmvlgVDkcGsRhbc9Nm6F9NgltR43X20wiSLtR11INACxfit5M7CLmYk9NmQsgzBjPn
HBCU4H3zTcyh259f+Q7U3DL8+jUuzU/WYdp9JJV0td0rFIOtTNm7YZergE2CGa7MQtgkXV8Jo/tz
uU3V4eGznlM06KqfeQwWDAvj8SwNEPJQSIlUGu66CVeDDl3nSuZ6yRT7+pXuBRasNuF00znVx7uo
/eSMFRlM0N0Qfo+FaRkDA1SRPHFIXSxxL5eHCHZhPbbWTsAmLC4SW35zicG0YNyGGTCp0iTqRXkn
UU/zhr8GnVxm3jMETjVw29KOspW+gZw2DcpEPWs5qsVahBqbD3IUd4Z1eP0TaziUmy6mbESwHG3/
TdaFGeAzkYcSDTH2/Xfp3fLrgP/+5v5pTCExs1tz3Ng2yCBVIXvhR/rhSOM6vb7mOS6fsN+CxJcn
J9ktBMnJQg2qGyBaNsObg9hJJ4b84WUQhHGxe0xBvTFQOsWjog+fEkf5dzYZiixXKslXvZIEdLQ7
JCbjfr+R4I6pnP0td8KWUuEZW1y+TYVvoe2xB5r5dJOJvDZ8EYUbedg7DFnLntIE/k32Z6QvGZj4
C6gzZu5/T/B0Lg1KZeCriKOLVbvS1FOrX2jT5+sD2axMX8yM/EIi/zYjfbzt9txi3j7Bofi6PGwi
FRQJPlXe7dkt8VIBVXZgxAQDB2q9J753L1yUWU1bA/eGtdYRqChHHWQ4YIW74BjRxCDcJG0vo87n
GFRA5X60kPpT8Kjo36j0LdOz9mq4nLhK4N+CmfLW/uNdEPLUgTVIuZYKDJNdpGzBdEgv3m335mRK
AGUlhrzkQoU6csjGCVvEP2iOMuWuUidleSxxYxWr6DjiSBPCc5QpLV+ppDHEpxePiAojojcxJjMh
kFh3EQgRpaeBwThADLMsOWNBqG7D9ykg4Qj3Xz83L3rmy1kDQWPO7a6FZx3WtjjMm0qnbLpQlmtC
5+W/GRLPt8pirwSJC5mn5BBL8OFgTytyrcyFH/RFrLzeKly99hQTFE7yaMkniwPyoEusVFFLt+0m
ziJDi4GH7bVftkqx69KgJlXJ0eJkM/RknWq1dwCZsbu9sCMUJxad7HmrdYXu87bYg3en5JNg08y4
gbPu83NFTMe/6sMNmCHKwFuIQHtWVj519D0zk4L+sX0ONYgXbHpobQRvgU6ZKBoJd6PvW82HKTSj
HvfazhcSjlHpsYrpVLL9U3ETrBWBOHmxcuMoqE3S1V36eC8A6kaas1e5dTYLAdVTMmPfWgU4DrOt
5Xt5hUlj1XMeGZC8jy9H1KHiyHJnKDLZ/26KEot9KXZjTC2Z6Ne8Cf4p6n9GRvycKbNRu/vXVqFh
71xJ9NuUWYcNlxy0/g8H+gWQJ8ZOwpRI1aOYV3xB9nGWUR1Vy5f3FESR9K9mdxJk8mrU57CReg+m
tiJGTSVLN2/imTGQ/Ba7fiafWCp2eOQ2SORT9dW5rV4WBzNWVdm4JntWoB8aw7phQ1nqib6a92Sa
IZzYTAb8/H8tkgcCYvoRwa6HzHWOFatXhlIpF5YcgbgVKf1J3YVgEkBWdhp6qXJaYzdTLFuzHjXv
kx8xqTvih0u74LRBDe1neHAJ8glHPjrQkNkX948yAXwmEh7hHni5TIFHOM4+2BBSORGgnEN40Pxm
OoiWOU+LKECb6CJuX+erl9Je3+Ozdd+Ro9h0n4hnwbuTYMGRPxx2KwK7iOJztwSzAEYF176hsbw/
Vm/t1Uj/W0VLkZZucGjhMrKuLP8HMO8Xsp1KQY8xMb+9g+sawvxzY8ikiDz3/jhZZBkMVSlorcDr
CYmCv/hH1/qZubtQCXWmBy4AfAFebOasIC9Zbs0zLgITzyod0GBDJy08CDejkFShLyZiydqLZFYM
R1OvPJMstS6GE6hKWAoCyzu2VmjKgj0Syqpb+DK6Szdhuk9fwv3psscC9J3nK0dyamLlkYD4KhzD
IxoQV29pREfb0j4OCtjehpZ/akRuZAWvt1f76Jt+vN0DelT6qBgCsscHQVixcn6LXhi3z0K2EYGF
RLrkNo2fogjCC5ZSo/ZA4tQsF8fM312I4Zl/YJ6c+jMgeeUXmydzIpF7nOPWRV+T1HM1wHrmE9FO
NYlLgVLmnyjRP76i7cjd5BsOdImSjNJs4e7f/Xu49baul824n3apuUIp/pBPCxkBPTTjdsqTs99L
0rMcH0Yez8YT4pC3fey4AlBA7al5mfiPvgqvMUc+z8JOzV8mHH0HMBI5zH0CsDswn0eH7g8XSpFr
tgP0umS++ctV1Bxm+ODZbmoT1qiqB9Pk8fNHiE4ltr7Psf7xvxB4jnoS7kxeuH0a8a+FyR7tn1Qu
Ut76/T8BX5/5QNXt6wPADYu6mEA68WXYCioVKCzHER90WG8FmhrnigWBMRfOYO666OaWKO+8X9Qk
a1SBDrXRlvf0xR98Cb0MMQiXX/5soVapZTjL3DsO2iHVh/MD9yhFF0PhaDiCZsGxuT/5Ae/r+Z2Y
YfIteNRWc4afrnf9E0pcq8C9IJQwYAi6SHBf4gg+d6BJbNuXwfy4te37MFVJmNjekUj74Yn2Dw6M
NLU5oT6fCNBvAM0FvEiBW/UozUIit53ytMUbtP4FTGKj5N1J2QOGdSHGTNBUm0aRBROla7aQRL2Y
rVJw7srzvI5LYNTheJyBBHjbdjD3+8y/FLBwOT3qRqS1HCDjx54g+B3Br3Nq60ec9QDNacQ+9jOT
ku6u7mUGzMLjl05j0AF2Lip1ZWDhlssmDXnpBKl4RH3ezjmxKrNYAKACNwDsJGdmlHMJrF8roY6l
u6RFQV/d59SnCuwYqIa0eXxXAoViVF32tQBTDi3iGi53pRF+zhLSim5Uyd1RVyRr1+DswdWtirMz
SzD0cFwnQDCVLj4KEIhggy7zGO9nT4dBrzcl4pQbiJ43xVhMFhfhpX3d5RN8KlfAlln5KaZlS/RZ
hGzRLBRhXPXT1m5up979M6f0zkyVLHAEwlW404PZ4tC0nTMSIGeGlpcKpXlc0hiejr07T/MQNT2U
h2qQLVsaiwZ/YQ9jZjwYtUwNuKPKHyDB9FJemi61+YeCJYKa3Os559SAeixixTU+s+yjGDMJLiZW
5qzIGIo3pJsYKRaT6nx13nob9vN1X+YNTy8vujKRVDWnSp1IAve4FTTkfXjSkz6UN0ccqy9h2ME/
VjZry3FeaFL4sXMgGvGv+w9aOTTMMvIPVtPYqLnFt3rsRVIgTsuWohy7fH7iTTh3T8mWowIJ6Nvo
Bmo1gjHl6wsZEfyZeWIQkQ/TSsyZKlg3fN9gO4ekpwAmr21z5xDawddjwb7ACYuxM88UZniAG7I9
az509Ndju3ekWzcQWsxHkbe4XefPruCaaPV3lIyB6d0cQt7O/ptJiLBPsHI3GEWiubCyVgDhRkGg
8dZJSKv2w3CJuFsk8SWHMa5ODS5w0taC5hvc758p1ibs3iIrtwnScY+/gI6QERYMOESZi8K//fm7
Jc7fxHcjkS0ZxszJh32RuJNeWHsTdG35vWtmWvCdjW9bGbNZC/rzz14LhRiThXw7pq5OoU/YvwDE
3SrptlmBF1j4YQUUoTWNNtlOUDBgAeuX2912jsuONo2cqd27BxJEaqjiZN2gp7MUAyh9LLdFzUyP
YDIUtMxSHua7G1S0IZ6HGGSEGRGPAkwC2ukfsTA/xJXF3xniOV1MNsB1CQ+Cr9qY92kBRZ8OLJjp
ojZ/q00nHL8dBkxmbWlkjeCpLlQj6OoszgvyJ7STB90ll+rk2cjc7MdHrDXmofNdgP4+QSScJWbD
9HEIc5AS4RYh9TtsvFV0cRetDZGPCWKdicqCt2e12er511puVxsBwKxhVHGgydAyWHyA95o/RBo9
5oizOwLAfcl+YQShLDaOKVy4jNCpMK6ORHjIy736IqgBRWhGZeL0AlgIJe+zmiZT6pXJyxy05Z+w
JSGZOJRnTmPZ49ZeHu6tZhHFsxfFYy/2e7v79w2wnwI0sllr4YPbH3BUQ5c93XZGFK0KDGDiAmEj
pb0lTOCBoCorPJrgpzMFOcCqlUc4ZRqFDELMoo6Rfuc/Q0k0ZKwQ091c/8NwfcH7Mt8nY8Hl0Le+
0dpk3c7iO448eH22wllNMCuA7jo5vWxY6A/FcXueLT98YN5jNNiPPQHv1iMfm9ChxjG+gt21J62w
uuaOYfi2NvgNDM7aoASwP2eaY5kdVHi94AkVpO1LaIdJWC0gXH6HGr/SO9EnD8Zz2jbvrpNigNXG
KE5HTTOTQOe8p4hUN80od+wTUqD6swFTzLWxfiFwx//nZZv+EFITWIONkgE8rmLjalm31K3Wr/Hg
MUQRPzB1CYq1Fssg2jRGbLpLEm2FL46iB/eSCD2OZcpp+Sl///MDnRIrV31lUtq4Xb+VsrtlmsX0
5lXCk5IPFXRoKfsovqBOdk+2JAVRrW07TrJ2jDQU9kGU/nybolj9htCjeM8BE6WK8PhPF0ctBNqB
/vxATxd17k8qK3e5Ub2783jhT14dSBBeeQW9rgwCXr6bISXTTpQG/+Y3rYbZmf3CaQ9I93Z0yaSg
hh3BAENBhQuKvga6ojskWXCtNBlYmv0F1GWcAwS1aYWy9XsZ3Yg2KnJg1b4YsFZ6fXUFlQhXTPh3
R3rUPbQ+wXhbVq4HPTTqCuTjmrnkOTWtaTylgmDQReRJKfjZ+EOmjSDvPiY4C206BsU7dt8p3r19
gvX3onByMoJB8la8roiVBsDnljKmL8V8d5ewpEKDuB0DxDudGovi50h8Qqchnt0wXPCeYjcF3go+
yTqhsQgrSmEycFMKDatxV7p21Ps2Fp/j61ehp/wTkyfaiMrK2wtqiBlnRzBHgVRRzlUM/qpVItUZ
aVGDAb9lDdSWBgULa/tHoXyjNq3yQ+EivsSxzMmcgdRiVFFG6V2zByRFeEEnIW1cWj1G+2IJHCqQ
gC1MEHY8jmo5OCtkJ2eXEa+WFZ7CoFU/lCAcmIrzhJCEBOJPOT+qgkFPkCp1DUKSJcOMbfKzvcF2
3L8pb++ECUE519JDUhkc6DKc6Gef7LmuRu+USiHb/jLDinliNqBXYFNIxOto2f4m8VLXIqINVSLd
Bc3dTkpfYtxOvi9GYQEmHUo8v1aGousMbdYLbsfqq3xUxpOhgfZV044HLfSS9rMGcg0abMW2hsll
TDFxHh04xTTsnRrNga7I/qjyq3rsMrWf/GZ8V+tEQM6iQ1Q2fSirIP7aJml9if99LvdAG6kIfnL0
bloZuXDe0Or7O71DXfLJsD/dGA8568YAv7q9xhaOr73kmXWiQe80rOtndpxQ+fRpj8tiIYkNKDwy
DnD7GYmzieTjTSAE9HRNTduadOKRkOi4sIsIrm6R8SELgTqux3kts3PkfpjyXL2D/wAod9LoOZlt
xYki8K2PtF34eOxHUnOJaXxFBPINkAhXM0T/DJd/3GWsy8nI0WlQOa5Zxx7cjz8qkq3CyZ+srPGk
b9gf2RlzRmwK6UQaw27fMWWwBfQlf9CyFp1wRyAsSAd+dZAziK38eYSzaE4P56JRtDUOHQ5CckdF
HZKjtQsnudi9ve1pfkBJXgZxdgZqkMG11JGa0gBRVxgkJiBwP5SXLoh7+ZcKCrrKb1vCCq0yvgeb
g+si+heWchpjdXfwfLTmLljG8KsI6MhlPZxPxycZmy0z9tb9WQxJ6wTHupk9RZf3Qf8+sVr0HX+w
9AIeaJnGBj0dEzxshLYvSdmrYXu1wnPJP9oXdczwJfDC2L4sqzWyPeFCgwIWIp6Xf81WySuYHlt4
/Yyajlk0iM0N/EDfleSccgqN1pqsoRV/aBTRjkRmtdvZ3s4+2U9O6jBCebaUGhY1FusNKQq8oXde
i5cKn2TuYnO9J1IVAIo9Vy21I4AEnm+iE9gU0dQcwuzt83TcpaQdeEmB8Ej7yv+gQKzNfYwxBBHp
dY55TQwVFHbnFSd7bOj9l2koR4YDZJFhtSy+U1sZbfDDZLpxpCothbGwEmNzqLrZcrTHsNjv0O6x
GWvwXyfDuENg8BTYHTjzrSvjQcVxZwIKl3ZGXXiUXL3GtwEgDvORgGjXhsK/hvJM1Q09lTfZ7Pdt
N1BqiJNBZALCH5JfPAduJcwVE63ZMpPYuYnGLG7GrAF5zqNIjheI6eKGH0ZAqh+xP95rFa1+lJRJ
Z/MZiuUEUnb/U9sC10/hHrDnd2FoDyNTYw/dMN1Z1iWq2ivc70rSbPMwpDOdct8cyx2rfafJ2TJG
lZI1PWM05Pqhr3GpBAIGvj2PPObBBqz6G+B/8KIYNr0NOzBeCMgQHv17HoS2C9Ms2yZCima4n6m5
vSIkmgmev6amF0Ihqg==
`protect end_protected
