��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`�����T;�x��Zg���)U�b����\C�]ȧ�n�ig���uWg����Gb��i>������o"V�SdsR����r�x�����5�%[x�
�e`J��:������D��%�֯qd�����D}`��н6a�_�	�ͯ�m�B�jpG�zy��b:�1v�cn��H���G�#T���n��-:��L�L�;Ha͆{���{~F���pJNG���&�P�>ҿ7�Hefv��po�ڐ1��R����J�䬝|�-�|���/���'O���l/��Tp�i��7Z��Zx-~�P\`J�{*c]��RȾ����%�T��I���՛�BK��W�1A� 	g�ڸ�ISGgEg�؀q��sn�A
��k[۲��4��IN�A��_�~o����Ž�Űy�z���z���\JJ&[Cic�H;ԱɰDT|8��z9���w�,��ݪ�����*X��j�th�ǐ�w����Z���%�6�������(�ف�X�\�Js�"�;4���j��{C	��z��7���p�s��k���U\N��Po���1է���uQRB �19S$h{�-��kH�/�;�7��!7)��Uq5����%A��C���U��y{JH.�s4i�����)�p:rj~Փ/�N�}E�^P&t��i���[�80iG0��:��f�\>��p^�K�%��#ՠS�&�k:�Q��q�4`�7�X=e:N���-�����_F�K}
�Ta�qvM�7�iU��-���ЯF2�H��,�~~������P��A��򏔄vW[���f�a'%�V}��3�e��:��˖�b^u>O��e��=��Nt�@��4��7G:d�Uy �N��!.]����?WC*�@�6�D��xB�|9A˓��+q"���{����}w(�Ԥ�ȍ�]��(���z.���Xt=Q�;��"g�A����-k4�u����cΔ�36���j�2M�wU�R@��zy@��� P�0Q�6: xr���Hm������eF���S����>�<�Co"��P.I=�8�ٽPY<�%�o��Ҥ��	J7���13�K����x(pE����{��q���|Oa��Ul����C��h ���3�/��nRPB��֡8t<�ɓ�Tj�u�������T7y�)���D��htHXE�SU`%�(w��h18(_��eȑ����$O��1�P��b*�������7(�wA�]޲s�Z��8�Z��� 迫��]NސҨ�*'wO�����-{%�\"A:��þ-�^K��7|�H9�w�xi�nK[q�vB�ih�F�%-�4a�F;PT�����P�>jC��}�[��c��	0v�;5��i$���Y��O�W�P�v��Sy&��Z\�0�!p��i�2��^���nlиಀ�����MA�5�y���\98�i@o5�^���tA�N�4:,�^�Q�"��^�Y�6|l� }=7�;!;���u���4�
|�гl�ؐ2'l2Y��o�����Fd��dZ����t|��h\�y� ����1�+%�";���#�ć��6��:��բs��\Z�{�A!�J�I�UAĨ.k���e{f�F��ڵ�Bf�B���.>�X��#�p��K���d��p|2�#q�	��3�QO�k�1�����VlBjto���mM�YJ�G��dc�.Բ��-��)�C"J���Z M��J�d�����}Xx�Ço+i����s���:�{z��;"�Z�6�lv�b]�i#��y^����.,���,���9�2b�W�Dw��c8�O���Z\f7���J]*����9��<�`�_UVk�O�5�N�;테����r=��L�8��h���� K>9�"��l���'���	qv��а����?��;a?�k��UD��G�6��F�����x��|��$�p;��)^���g�<��)!A9��@m鴘��U�ѣ\c]pB�l�D)m���^Iq<u'���·���/��v����9k����O<URL�7w�'?��qhR�3�e�=ٓ�>��)��'��\'e`;� fһi�p*Ԋ��Ӊv�R��Kzf �:�1���X���]�,`&ڍ�}sa��$�"8�D�B] U�M_�
*�WA2
G��m|�����d���wj��fl�g����W�V��� ��z�������?mŠ<A����b�Z��~��[ۃ��Sq�%[8��|Y��c�x]�'da��y-@��3J�m/ ��D�N(t/M�������o;m�+'j��I�K�������rɳ5[��ճ��;�������=ꠠ�`��h����>���V�[x���0�����9ږ��C+z>7NJ�a�٪dW�p��{�$c�2c���F/�,�$~a]gvy{�!�j��u%d?� p!wmB�Z�EG� �"�7n�R>��5
�mcƄbu��Ż���ƣCX�J�i�z���nt#�S�����g�y�ǌ�C��|��i=��#�_��)���oCB�c�9J#�f���rs�^Y��|�2��S���D��}���#nY��M�O�������3A��3�#p˳���^[�IVe�{�!òi�&h����R�Fepͣ|b��HPw�9��
�ۆy7@�У�66I�ƻ"
�*�H$P&jF��u����H㲳68β�]���+Mh��}�s)����v�������Ā_�)�T�������+�s����""������l�L�-X:���[}x��Cf2{�O��NX i�ۆ4aS:��#���� ���@&��A�a�^Ɔ�<{�$�����^���O�4�2X��^�{�;sr� �8��-a�~(W�.6[�}��q�$y�o�yaS�þ�9	���&�5�ù��}0�ݛ�|��ڡŖ�&�V��p2()�C<T�+����q-"ὒ����j§���S$S������뒐)S]�%t��'��_{kG}��իoO��eVb�Z�x��E�$Te_���4�0��O�Վ��C�V�W�,c+�ڵnD=A���i�n�IPq�;������D� ɶ�;dj�d��f��}���?@nX�6�D��x���/�m���E,G��Z��I]#�o�M�
aX���/�����3�t�G5�'�]\���H�_�JTVQR/���z���lK&&�����Y|�B�u�rdToD�6��c���^�e��e�[���Xr��S�h�Zj��Jݑ8^�e��A�U��ca�8}n"��e� w ~�^�5^7��������쿅^(tz�As��h���[QE�Ѐb]9�BT��6>9P�y�P�4K
Z�d ��z ���:!zq�y�3(����[�r1�5��ߗ��ܖ��������p��r�r���������' ��Fl6l�}<$Q�U��r����{͡�[Цg��%3z��!�X�)6�qx�+Q1�b�&��I	2�֢iz�2Na_p�d#�P�x���m��s,Lŀ�|�L��'�Q�쟖���3 �xud���+6;1̼/7�R٭��#Ap�"�L�ǲ\%�}�bҀ,��f-'���g.'����@lj��J�o2�f٣S�e��{��r���IC���¨��
3Fhݒڲ�»8�Ï�\˄��i]?�Z�����9�σ�����<{RA�t�Ow@�N��!�t">u�L{��he�E|��/��p���#�3L8։s�C��^1�h��OWj�b~n�(��0�n�8{�9�z6���gg�j�c��~�~ш�w"<�waBx�V�0��1јbz�t��5���9���������IMM�>S�9�M�CY��u�ױ{n�Q���C���bm0Dǩ���[������豲������f*�:����;�I����A�*ĉqz�&����e"�px���;JU����q;6�3w��K� ~�|��{t��#1Y��?�N O܃<ONL���Խ)��_���$(��-���f��&�͒���vB��!�Y$e4�_НCb+\l���6�[&b������h���k���+W\x�"������$�\w�W��k�8�)��e���n)"%�����̗j�k݀��q���̒ԨD�CN3d���BvR�3W�۬��7���*l����}v�!k�Lj6mWG�GէgR�;z�pn)y�F�[��@�i�մ` I��T�%K~!����D+�����1��1���B��p��u��C=��G*0�c�R�P$!���a���%������޺�)q�"�lދ� ��C�һ:őj�c�40��2�i��LB�1����Ȫ;�c5�{L,�����R�K�D>��}�6���Z�@���@<ӓW���ɂ�lҔ���m\x	�':�ܘ�;�X6y��L-�9px�@+��>���|�n�	O�$��F;A`b~P�>�}(,��x��?�����/2��VB}T̉�ph�&$}-<M7ͩ&ߔS�GY�19:��Cu���v�/��QOi��s�����	�������=���4fH���E�����9��Y�G�]Xc
Ts��̂m�R���\G�j4�~�`\_c���y~��VmV�\�^���|�O�Xfbs���j-��2��yȫ�?�������G���S\��f��D[a��+* 8?�O!Ev��g�_��~�<��6�Z��U��T�%_��%���:�$�x7��9GC�J�E���๩�����$T\��*j���7��O�e���}�>�+lw[z���X�cR��普�Rn�sC���	���mi7�h�<|��zY���:�-
;]�Ac��vJUsx�rO���Q����~�j�eTL>3bh���`H�bvk �D@�:������$!��BE�K��M�M}|���k��a�h_y~��N��Pr�9._���$T���J��xLm<Gg�I�:F��pW���,��u��>�I^F�a��pC�SM��9d:��3[`\T��#�c� �5������c+l��1���AK.��@Z���!�,����I�E~��[Y�7�2M�ͬ�5v��c�u����sU���'���=���O�~��m�;�T}��A\�{��cSG������M�zjD��闾@�c{�E:�����M�_Z �i�<��PΗ��ʕ�9ϯʨ�)�R�z0?��a��U��o�mbO�3�A�.k������T������[O2rh�� $H��T՝�� �6�f6'��)��҇8Q��d#���`(����*+�b�I�w��!gSj�><j��yV��&��+Ũ�4"yHF�|��oF�e�Q$� `�ߊ�6g=9Q��/˷IN�E�&�R���H� }�E7��ːq�a��E]ed�^���<P?rW�.��6��ř���Q�9����8��grj1�cjA�6"�d�$*K_*,d�\.�� p���͊�F��ce��Qx��]��E�BTl5�ܙ�H].��姗ߣ�7�:�Hm�Ϫ��p���"��Շ�7������/�+�W��x��G�Jc����Ke�z�wQ�M6:�s��E���\P�E)��TΟ[d�֩(�򢠲$��H��ph"Wl���1�UcZ�oh�>A�	��է�"0�ʑZF��؆|q���B�)l�{���g��8Ɠ��G�#磭�Z�w45�C�>�;[�:;A8�3���po����/�K���n��:l��b\�1�V�L#���^+|�������2�t��� %�"T�E�n��^R�ڿџ��T�\��@%7W������Q�C)v�`��K��t��U��|���6�?��1�ʔ�TS�γ�6QW̢בI1w9>������H5n?9g�@YV�9 ���Io&�L+BY��qӄ#G����t�P��:�U�a~����-Ė�#W��AHI� �y��w��ԇ�ʓ�ڂ�đ]p�9а4�H�*�4��:���;{��:��_��4�I~]]ȥ��C4EIxzj�W�`�OĖ:���Cm��Kqw�{
� �f�:�{�0���Jj�[M>24E�Ɩ�K�v���t���է8�moŝ��ff��w�^�;z�W"?�u2�6�Ny�0D��!�����@,��{���F�*��!m8��G���r	>
(T{�Ҡ"C]7(b���h�~<�*�=��v�K�&͹��[����`�b`ҧxX9�v����U��w�٭��ԃ<f��_��p��O|/=������2�Ca<B}��Cg��8����"��en�掙o�X�S7〓�J�]^g�4��쐨@� /�Y�Qx�g��I�
	- �z&u�cM�_���}���y������\��B�/�fGv�&��g�_A�0�9�����ZZ&��vͦџB������V���E���J
J�OJH=�WK|�:�b��J<e�- *�ú�j7�/���zȝ�~�R:I2<N�����f��W3P�����ۖE�G�(��Z]v��M�'Qh�JCn�e�d�;�:�I�P�����d״G��������������� E�S�VK��0X,�4ӻ�M9�(k��ɩ���Oq�,J�NJks���^�[�-��+���x�R���!_)�OF̑~�Fκ��L�X�Tv���J�D|�5h��0�|�ّF�ڮ,�_�vR�0)=�G�vM�-�3��%���h�BW�����b��Q���N��FڇE�s��'��s�}����{�E<�,�ƕ��O��7w_C@FO���� ��:����?����'�F2�,�Fn�"Ar��ҥ����jJ k�kX1`c�����4×���z�j��a��B�-N�C�}[��	�b5*:�S���!���gL�B*ک^�O�'O��t~W����д��Q>�ˮ�s�2�M�a'�2>vΐ=�>�W_�@]|%�?~��f�� �����>�$���|X��U�r�l�`���	_�	�Gd2_u�sSdo����Q���(��{�@�f��.�c�V��j}���3��ѝ��x���A����橄�f��W$�j�������"���8�^b��&�*S�� .�1���s���C����� ò�����[���F�H�ަ�E�J�N�c8�ux��q�e��o5ޏG���̺�\���h�/V��I���m�L�����m(m������O�Ct���}VΪ*(���A%"z�����'^�� 琅�u��>btՉA�?W^k�v.���~Ve��Pr�a��RqXVX�D���PŲ8�|����T	|��2��s����{)vEq��u�4Х��Z$���Y����*_`� ��$���[)H�%%��bBt��0�[K��B9۞#J���y,�앢��KeT��n�I���[�\����eL��s�O�L /��x�U�r�O�0���h5N{���M�M��Eu\�9���r�P�9��R-����i9��Iz���r BY��M| Qy�:�6e}�E��HF�;֭�蒱�tt���4�K���}�lg���7x1OZ��3�2����`�{{�����i��h��-�C����b ��wď��8y\���b%�ӕ�l����5�͡�:θ��|�V�Q��}�z�dF��%Z�����T�]C��垎�(�WV���{�Z��vƄ-�ͷ5J��,1�b�*�"}���7�� �����C�.»
5'�\NW��j���'�LOj��w7���pQ�X�f���8u�6�.xSt���~L�<$�e���Q�`6IMB~|0�������?�2�%3�[�jh����tZb��K,c���<�-=E�ڗ��g���l��A�נ�ZʝE�0K��@ϗpf�b\7���}�{�~m��2�%�ξ+|��'<���6����o��"z��3]��(CSn�_W��ͬZ]W@7�ّ���Z8V�o*���p��|+}R ��9��t�*�^ӵ2�o1X�tL&p�뀣�Q�r���;>/^���ã�����d�Pـ8�nQ��FP)K�ӥI0�t��b���9L1?��79�㺝��Yg٦�?�+~	����z�}��scc��ƚ'-�r���@ �J�k�Eo�E��y$��o y%��Ÿƴvp�!	�F0_���P�롎-$�B����a�q@Z��(��|]��ː_�E|��ڪ�����m:�$����0���)�kh�w2/�2v<�+�7��V�G�K�of/>��
:@K�K5}H�V�R3�(�OB_Ap�m��6p�E[��"�v (�=~��PCTTh�ӳd3����G�Q_��er�~r�Ͼ��*��-��Ǚ��)��L�sTWH�/�bt*������>�X@̃Xg@���2����2c�vmN��^�)�|�>���r��)%d%w��Eٽ�%�>]�����,f5��[)�|²z�p;�`�(\���|�N-'#�`�Mĳ]|��+�ge2u^(��w�ϑ��/���;�_��06GD<�4]�@`˝���55���C�
�%�Xh���P�7M�ց �'âu=��(pt3��j1��1 ����i��8{o]a�?jJtqM�O�:�7�ՙ����(�FN�>j����9=a΁�#�������N�,�#�b�W�	̠y��G>��Y�r�E�)�<j����$X3N8+���CV��@��d��B�S�f�kf\�go�����KU�c@S �U�Y�A�g渮�L�yZv�����Sm��e[��)�e���C,�����Q�/�I�c#�h���A�kiXS�{�/k6Ӎ7��'���ls1����N��kv�r�^��.�d���5�&r`��;(��5]m����Ej� .��1��p9�{;f/�t���� ��w�����IXo�A�W`����tR�~G�k>6��-Ά%b6ڄ���[�5�n`$A} �\2(�x��05;��Oz���|Y������c�
�Lg��Q�R)o�:|��z��ۭis��
-�����2�k�W�[.Q�k�[uG��:��T�6xd��+!O��L�m��˸K(/�����@�Dts���`�}7�y���7+#��60;�V2����|f�Q�Λ\ی�͗P1A������w'���qFFBW�J�6#��"�Lk���5q~���� ���@W� ;��}��#�M۳{�ҝ{\Q�y�v\�/�A9��IL'e��bJ?Nٸ�9�J����U�m(�Q%5�����5E~�;x��I��Ԛ�q���ʈ2��������0�U��g�J��ml�*L}���qȳ�h��8K`�Gu�@���L����z�xc6ҵ��@U�����_8J��m�>s� ��7�������dw��;��k.�3m1Ԁ�4]�c9OR�\�}y�vv�b�,-h6ΏS��z��Ey�hQvF��G�(�ϕ# �T��^��,���ـϻ��+D�p�3��"���P]�1�|6Q�0��� ��82����<g�8�����)/aQ���6[�&����-}=_ց`��}$���Az�,�^jN�t����G#����	�o�(NH��X�9����)
"
g�=;%}&�F��ZVpR�	�\���\O{c#��iu:���dk4��=t����٘v�z�.BV�����^�-o�!cOA�����h�����Puk�v�4m�\���$��KCSD:s���^(�;Aa��I�oZ�O��u�+�w����F\O�@J����H �(1F�z�C�@��3���ӂ��-���0�T9��5
']�����/jh�|��E-ޑ�绳�u��_2O�J���m�4�?b:RX~�D��?6��|�4�����u��Nb&�4��$a2ugQGC1���J�}��&'0&z��QA�[�.li��Tz����G�[�b)Funq� ^߰NØ�^�C3���D��)ի��B��Fz��d�N��9a��;������Vz6;����~��V�I8�msܞ��϶9�c _��Hs��X���a���ިϪ���EQ�7p�K�#A��]-�B9Ϩ�(<�����I���hx������8}*���AG@t��X�����S�B43 m�M&�=����Epb���6_�㴓}��]�(�^�3BvX(y��n	b�	��=#l+�dQ7��#�P�䉩�j���bW@����_��`�P�pu���l`�8��e"xH"_4����ԫ�=���e�2-���(�B7� @#d)2xT����s�`05���A&��V�Fe����wR��N�l��c�y�Rn�fqk`G|�FD�6I�E�(ƨ�dx�$eQg���H�;����N�Np�ʙp�I8lq�P����xR��@n�h(�AT�����.�yё#)TܜC�g��+2��Ђn�(CP@���?	����'v��嗯Q�����=������F�$Ô�F`F��k���ax���t9�ź� u�[ΐ{a��P>���ٱ�ꆧXڷJQ�y�Y��/�\���"�gFĝW��X ���EN�����G�c�I���	�?E���/H�8�=w��O���5QȕHN�A���%�>1�;U�*�=��ڳ6�1\��g�d��q#��
"����� ��B�[��4#p;�K���&�n5a�E�����̡���aS��Y���c('T��)�Vϕw�鴢�;,\dD\Z��g�z�.�-_��>�U��5�T�D� �L䅂	�1'�R�-�����:D ���r�sBF�ث������o����
��):��>�&��nF%� Զ�qs7�;���}
�ss��]pa8W�$
����S��Y��wbB�Sjp՗¤Ulӿ�  !^�Z�Z�*��i�R�4J�����[����O@�4J/�x�����kp�ݵ[��XĹ�q���0U���ث�Q����[L's�$B=�c�
 4�LC����c�N�hX���A�I�\�%��Y
EC��E@rř��Q	��Fd��bA��2��S��v��&�y�������c�cl���v�:Yy%-/}�:����,��d�W��~�<*�W��_pKڡ��j���zj'�&��:�)� ���B�����\��&r���\�&�q��_� HPv��_�$��l6m������>׭�%y1]�`��A��2t ��9�����5��|U����E����@�sy'զZYo8ɳ"������d��Xc����X��Uc�x��?���!�pϞptCur���H�h�m�="S�Zk�ww���>�M�����ϣNטf!��ݔ�T�ow?�	����T���т��n+r��@�pH�!��u.>V���;m����*5@X����Drl��d����:�Z�h9�2(l�����I�1�0�A��8>:i�/�]���9��@�饭��Ѩ�{mps��E$8G~�-|ex�e ���Bo��f��a��˜���g;-�0� �vg� ��#ޢϗ��nx�O���A�32oV�m�$���#��M���?di�h�t��%(@�%� �� ���'����=%ٳ��c_�ͫB�\�ک���ܱ�|�N�f�E8�@���OP�S�&��z�xC�Rϻ�R��Kc�.�y��q{�D����c�}'�#���y	Ie�J�Z�Y��P�eW���GO������yv4��3���r*,���&��X����F��y�+��<�Y�2�R�c�>�:��A�������d-c���2�b5C��s�t4��6���'`�m�n@Z��>{:���M/�D�_I�b���E�
� oَu���-6T:L!�Hc�q"���K-OH�/��>.�z��b�H!��l�Hׂ�]gyma�J�(H��R�:.?T�Fո�Ǹ����W�&w�w"H��i����l=�����QTP��������P<M
�Ud-��}���c�Y$�t�ecc�63�8���ܭ�1��i�8Pm@t&9-=�h9�8�H�FV���9�����Q�]��XL�ѩ�"ۺ���G��2\���oǶ���:-���e:������ЕJ�*�[PgH�yn���\�7
d ���;D���K.���ZL��u5�܍�9�:s&{��y�6�W[�9��`)�<�Z:p	�����-�� �wu�'f�B@����X$��'%]��1�;�d}�2H�����$2#C�d��C~��Q�}tBw]Ne�9�X��c��eK �9^6`�o�$:��U�R�P��H!^�8������a��eHGq;�O���y���{0����/tX�@��ID�]z��a
{�[�j��d&� �`�
�@%��B���^�4[��M�}1
�(R�����J/bdE|��H+��=��8�}��$�W�(��� N	��r�Q<�厰�.vBҹC7	���H�u_�0GL��_��. F5�0�M���^(��4����^6��P)R���:���?�Kv��e�2�I�'�B����%.\a᝵(r�@8��������q��ԭ(i�I2���:�4g�ɔ(T��頰��̮�6�/��Ś�`�i�hZ�2dS,����]d��CuV՗ىB�J��ҥv+����|�î�0���rbxeo��t���Y� �5�L���w�[׺]5G�x1��v�{�o#���饹��Ջ^�1i�	�j�|���{" �}��'�\������'����ؕ�Q�,-�.+�ZpnQW�ipM;��:�&o}?����>$�����g�"��q�� Vt���m;��B��5q�����Qaf�~).�����̗����F�<Fn��.(�S��������d��Uo�3�|��f��7��S�6��5������g��p����"%2{ߦ��_�j~�<�O�6�nD{��l��~'�u9���N�ג�^�� �j��|��\=�X�4K���R#��`��D�WZ�����wW���d0���{Vڮh?�Bs�};)�Ƞ���ѭ>�,�{���K���C\ۺJ��6v!�R������� ����Zk�k~q�g��#��qE��x>"���w�����N6#��R�&��~����Vo�Cj�gX$������yxf���?��R'��a5<��rC:J�C-���td�yi������[�0:_�\8+�I��?-�Pp�϶��U{�;J��_r-�z��cW�'�b��I[���^��@,���\<���M-�l�y�]Z��QC�Z�E�_�`�T ���?����"�dǷ��rО��o���)fdl�do�ɁW���?��6T+@VimVpl�]��mo�����93�[o��e����P������Iq8��L�=�e��"�������!�/:�K�^+��s�yX�?�B�۬a�t��P�,yj��-d��.xo�^�S�6����g��)�ߵϴ^�F�=B$p5سnt�1Rʵ���N�c.\�̪]!�����,h���c-��>�Yߓ��yR'
�gRth��z@�j*c�X�~)A�\�7�V�H$�#[�\��s�W	2���v����FF^k%�v@aET��,GR��1�2���ʒ[�͜.��$��V����=�ZK�I�*�g����`��4��C�E���2���C��{T{N��f�G(9IF�uny��`yPȲ���(����w��4vVL�o�_$��B�Ae@�}�y�?h�� u����h�h\��r9�y0"�H��Wp5d�0R �V��M)8U�(Z�ᝯ���U'�ƈ�<�tCz��!S5~�.��Oe����5��7���77[��t$�bֿ�Jchw�o�#d�b�9�S$����[�{^K�н8xd�xVcWkU�_ˍǫA�i�Y����~��dl�¸E��8�u���H�\��.����&�?^枟�	v�_�__��ݽ>��ˤ�d��z]�p��{�m��yg�*��g]ؼ�me�V��%.�Wt�L� THNBlJ��>�:�;�y�xU8��V6�O����>���V�˖ޟ�Xr�Cǎ����T]h;V�t$��0�:�Y��ï	��y�o��Opy�r��~�9ȴn���Ep������j�W��=�Ub��v#m����~Q�I�W(��Z�D�ɱ����>�ʼ[]�em��ICk-��U�V�*�o�c{��p>L漡)��)C�����L�Lt��I�B"��c�܃w�R"7����+l��	�'Ys19` ���G�I�;�u<q�Dݥ������;���n�V:��M�I�y�AL��߈YQ�YTCs�ΰ`ᦱȔSRa#��*��fK�;P�Z�gF�
?w��^��hnb�OT����J�3Z��XS�#W[�ek����\��U㛹�����q
�a�Ux�����!��>N6w8�<gT*���\�;"�p�����u���O`���(�ڨ�+���P4ul�p-l"������a��[� �j��'�0�x;���d�Af���_��o�Ѥ�5��0�0����NUʽ�#��TŒ��a�k����O��Um�����1��N&�>���=�G�bmÕ�$&T��ę��h2�u�73ǘ�dC,u��>Y��M�r9���-"��5 �o��^~�o"}�L����zG#���Mo��X�~�6z�f#{#�T�NU0y �	�S��0�h\�kZ�x94�{��F��s@�'2��P�Aؚ�*hcx fK:=XA��.���fG�rJ��K�,�����S�̼	{rypd��*�c�s[�~�i��ٟZ>sL��A�~�=W`�.8�5Я�Jn�3c��܃��pP.��e���wq��9�+�bcq�������L�����D����X�D����fko'��f�Q��]4h �.�+�'>�7�\H�@�:����Y.T����o���ІO�M�o��>[O���	K�SD��~�Q7�^�:���L^�Nu�-]���.�렭߷F�6�����ϩVƧA�K�`��1���_��W,��8=�v��dO�#��䊅��_�,X�%��z���^��둥 7lux�i�v4q���_���W�g0���rM���W���� ��:�l�� :��˘ 0����>��L<n�IJ%%�X1{��V�쪅~LN��,�g��rR���&�+ª�^;L��k��3���M�d��|.F�i�
�
Ǯ|q��I/]�hK�$����~�!��>oC�W�O{�M����m�Y�H�g��������T�<�����;N2��"[M�=y�M��2n$�5S�	�"2/ʾ�y���{Չ���ֹa����)1,	<,S�#x��ʮ���-;�[�?�g�����#��V�%����{O��V0�)����6�Y���������i�m +*�q!(^{2��K8����n�������2����3;����i�(�����p6�>)j�(e��a��:`��+��|^2��],���%<���Z��B]�����@��;[��V��������[0Q�'$���r�yA+�g|��%�N,
�h賢��^����)����?e�P.E-���'�T8�9��[.7#i��rǜ>Lt��UK~��#��eB�ǹ�����g�F̵�x��߻}��q4x�/;��v+G������oi��]#+�����S���&��9`�]�hK�^�O�Fd����K��Q������Gz�%�7P�GfuB�ٰ��M u`���6��$<���U��D=����-o׹T��u����K���^��A������i�������=��������w��>�R�9��4�2-�X���2_���B���(���$/���b*�8�'�tr�E)�\1����ǡe�a	�I�[ ����+����V������8P'4B���3`{�Ǥ�� ' ?�c3���,������U1�F�=>�f��HP��A c���%%nZ����",=[{���`�e`�'�p�q1u�KČ��dĚ����P�|6��ŧ��}RE��|��ldjx&>���G0"�^�Ώ�NrR�L�,�@�u[��!D�pErD	Dּ,����7 ������R"AK��ģ�C2���vW���]do�zFp�=8d�}W)��.ض��~��+�T�w��x�����Cö�Ҙ�o����X�j@�(i��W{�冼5p��/h������Y�6i���e�@.~e��c�O
I����֞i&�=�[\���>�(b��j`�qS ��ik<����<��y:�霸1�fI�%+���#�<'Bf�Ã5�v*R��ׯm���Eŧ���I�`�
��\sW4�����ł
X��ϣGD0[��F�M�C�0�`Hb<��;�HN�ۭ�e��f�L��
i�<]�9��T�7�[!��y��d���3��/YDzyt���v��9kF�@��H�d-R�=R����5�\b�uu�-��M=��a���� 7U�S�p�Y���F�_�T����3Sw�]�z���Mdσr�>!�V�}��P�)���$_]��]�� ��J��e���kiQ2XR�F�!||�io�epU�E�D1�4QT~��q�7��~�ѐ��Ƣe�!���v7�F/*tN�j|��6�Aɿ�t�G��	�{^�-��oO��ٴV���MY #���%c�O��v�#��e�kr��MZ�5R�:�Rl*�/�m�!#���sĒ�89;���w\���7>"62Iu� �֟�\v~�(�������}�,��nJj�Q������
����-2nPH�V���?�ϩ��I_� X,�`���e��RI��!Mԥ�6ӑ��8à�����y ?c�0����m(y�C��,���k�݃Ƙ�2��J���Y�|�����ƤA� i���6H�<���x�}W&���-�w���������Ǣ>��9⴩�$�h�P�	��c���r�CcS��?�����zi$�:L�Q��)0��&�o�+���`}�4q�$��a`��{I��ܣ58��?�Xgr�"����zc<��"�v1_�@N�̜8
GeQ��F�?'��Qwik�ir(�����I^_�?G_�م������0F�yF.bH��Rw�-��f�nl*�4f����d��8�>[�2�B����M��(����0sy��t�V#U{p�K��B�^-�Μ��r����J�iK�{����t�,�MX�tl����szv�uw-fU�o�!�!���W��-��ß�@���}���&�nJ���U�6��I]�|�0wH�����eI��c@g�{���gD$�W����*��}���� *C�Q�ț�LY� D��O3�� ��o��7�������Z�0�k�>8��L��;�b��D؞��l�r�|�� Φ#�ZR�\8�:W��8@*4n�Z1��� s������-�A��=��LzO/N�z�sG;��ԭ2�C���ƛ�2p}�Rb�#M��̀����$�pU��2Ծ��th)t�R�x�VH�k���t-I���+�� ����^v��<��O�%9��v�E@�����_	]xp��s�
VwԜH���`��ћ�L�'Eok�?s�k�h:xw�]A�v�0��]�*�.�tZ1��FG�j�#������]��AS�H�K�Hj��1£
]P6��_�=�
g����p�i�z n0h���b$�WD�,}Qr�W�`���p[;���-	�/�>b�b5�����B���n.^SV70�X8�XS�+�A��VE�,g��<t՝�y�9�!�>/�GE�-�p���S���:��w�沙]�����|#@����
F���,���!��~S��Z����qɡu(��/-U\��Ǡ �b�P�
���oLӁ��~Z����n��b	`���m�?*��0��hI	�<�]!ԅ������n��d�l���o�� ������!w�����T�ls �e��-n~�CxJ	�'+p����QE�<PzW���>]��c�و�+K;�������.w>��Tx_H�C����.�yҪƬ.�>av�������L�6T�peV2�8#׾�0�����3��!۵/����q�V��\�~�]���5"w�|��b5��!����?*s�����[��:�w=o&���0���|���fpEQ�ME�x&6,�+���bF��F��qR���OO��Z��7%���}+�hn�\�~kЃj�� �1�x"�>τ����FV�����B%bV�l�1�fb,7�Un��cFhں�'�q���*��9h�<�1E�f%�G֜���=�f�y�H��'�@� ��F�U��SIw� �^9����hv�>V���yf��,}��du/J��A����j�7E\|w6� �_M'$�B�K5[��D��6q��¿���j0L*�v��Ԭ 5{ԧSA�+����@��-yn��2�$�T4T����'���7x�Λ3��E�7������iw�f�����&p0�!����R<Bҫr�2nՂ��2ϢS�4Eʴh���^���Zˆ��Q�cGF�B�us��bYw���A�T�-t�d� ��w ��S�;�Ï�[?��w�99!�D�?/�i�wq�:<W8�P��mq>AEb��_g���w3-��F3��ȑ�#.��������`.�!|��_ӛ�`8]���.'s�"@�̼6^����R��p����0�����O0�K�> '�:c��w��� ?��t�p�n5h):��f�
<!���}v�Jo����7ú�z>��R[[���6��T���A �s��ϋ��66��H�?�QnL�z�����*���
'����pe���P�*��D�{{LJ�Z��Ѕ��9�$(���#������+x�A�y_��d3V�d��Ck�~���h�K�4�se�w�r.*���̡�L.���ј[��,^f�,�L7����N⌷L�$(}k:��E��7g"A�΀��7�c,
lD�Ň��f������8~D�V��L]b6mt@��<�%ǟFN2�� ���2 ����%�N�d3���f̪�lD��J����UTZ��ׁ��F<�3S���?ҿ����{����\�z̩<y�
3��߰~Qv��h����woc�ʷbG������4�<xЛ"n෾��� G��2$RQFMi��rٕي�d']�7������Z9p�����i�Ut����{;��1�%~s���z�K�0r���>��&qb�I��.��Gݛ������~�]�(����uS�&���vmo���f�_aB�UW�]����H������{��9:�82U�ߙ��Y�DdY�ǳ��b��S�[rJ_���gGUy�&����#t�����t����p�R��#}�*ߞ�ۚ�M0�vO��>���c�I��H�M-{b��[d��99����0�b�W ��%�-s�S�)g�� Td�$6|��e��|�Rw M�
��X�mxo��#o�L�ʣ\a�f������0���tT��JВ��q�z,5,5�`�^6Ň��/����yӄ�g(�˒T�h���_].oh�K�">0��
���U+��ܨS�4rj@8���{���IV��S�h^3���ftRdg���J븵�7,`��g��d��buMm��I���?���Ң�<�݄�Is/��T��TjOFx�2�
���(���F8ACkE��׎ƞ:����@6��C���*���i>BQ�x���>H�^�>���LP�������Om�%���<�6W���i�Ccju�u�9O��92���H٠5���h.0������(��f�/����g�����!�S�[���y������l�/��f�š��Sc���K�^����s��#M=�p�A���@���6ǌ�D<~NC`4�]_���+Մ�8
y�O��$�j���}�/�/.�N�q��T���׺h/h<���h���n��{���I�=hS�]K������0T@�s��a�@�~ ��';k�3tc�=�B	Y��gMh@/�A+��ߩ`���yQ�w�Y�m(�	�{xO��t����ȭ��(~��d����A �]Jxk���V�PBu;꼊Gm+,Jz/t�7!C�p��,V@g�R:��<
m�"6x/���g���o���e>E�]I�2�����u�q�aԟ��F	�	ƹ�p4�<2�>vgY��ٶ�!3mx�-JĨ�={�rd2!�L�P���Uo���W��QJ"�np���|����|��������b�!�� y4s칀�KuH6u���J��!��t0�Z�S���t��!���蘃"�b� ,�>���-��	Tj�X2�)l-�d�m[H�_e��ܣ^�ඩo�Q�p@e.�#�X����Ǟ��_���b����uB��V6�ц���!m�gFF�Ȇ���ڱ����6�E����M� ]!br�!?g	���x�&��t]�F�E޸+�7���7Q�<��N޵�h���6�k˭X#�%����T*h�|�������5TgF��?�Z�#	�]���Abk�cx���{z@��њA��O�Nvބ'!��xq����,�vy ���a!}l*��0�'@�l,�q!�D�����Ó�J�ӥJ+,��s���R�!44n� ~*[g �	�7ݞC[����R�GY��A���\o�;���vw��4��HXd��J[�^�ɡղؼ-Lhݎ�>� R_0h.�&��ѽU�{��@(0�t?+A�c��ֽ����-�M܉-_�n����o�8Z@k�������#�ݵI�a����7bU����Dr�p�1�D��΃��p31�f;B�n�����{�^D�[�C���	c���:��y^D� ,\8���V�i��h�UѶޒ(ly�rm���Y�C?��0J���$�*_�Mi�O�� �[;]9�m�+��z�@5�kW�0���Fa IE1�^��S��U��F$����7ʰ�M�Hk��5�M�X ��	�UI�K��rrb�?`QJ�u��r���8����j�� �Y]q����̓"�GfP�&�����N~A��'Y�a$56�j�6�و%�~��}�tR�!G34���)20���"���*�vܳ��"�1#%�����%���,��h�{Xu�1��/�u�v�*/�6%�_�x����z�JY�L���g�2[oƿ���`�~����(�k|T�x�0�d嫶w��y����!����;�骧 ��v���øE�E�*.S] ɒ�S1�`�C�;����s��X(] ��ΠqƯU��~��r��ßS�ۂ���hR雒�̞��x��1�pe\2O'n>
�G����U�z*Z� N_��:�~�	+�xŭp�YQ D{jҥ��O��;�VQ�Jk�v�]�����b:��22jV�a:: ��J���pk��lyŕ˗X"�{�Qc����"���f��0��PF�4�n�	Q�w�����b��!!�0�d��f���>.8�,QZؓ�	�#|�J��BHB&;�Q�2�^�Uؙ�%X�M��H{�.��F��o��n�,�,�wY�{U�f~�Q˳i����ɶ-�:ȼ�w5��/����'�z;8�J�CK�ki'j��ä�C�p�&��!�T���M=�r<j�k# >o����oЪ�[p��Sݢ FW5Ө���sڟ���е/H����M[g|nM�� E$^���p�+��9��]�Gk����I�/�Fş'��i�բ��q�w;��݀�&�Y<�6Ɨ�G|x�n:�ȈM}w]��^��-.��?dr���R�=�Z$�cE#@=�mD5ў���>&|-n5*Ա6&&�����������0�y�]rV�(-�`��K-J|$I��������~" pE�j�=ND6.���%}��o-�2���O�O�?���W�D"dngNr�fDel,K��/�c`����j�38[|(x��2	�i$�e��� a(! �*��y�/Ψ������k��\l�3�����&d�g=�d�0�9��7��b�?���yD���wc=���&�+�	?$��P�|U���!��U��VG�����] O+�0�:�4����D/���|����,��Y�"��.oi�:�������D畒�i*Fʿ9K��W1�z���[qNYK��a{�������Ex�s⎳�s����U��{�B2�D���������+�~aj����vZ�,gwg`B�2�
��a��k�G���t0&��tF��@"���	�cA	*##��4d��M�m<n´��̐�X4=�Ku�WA��j�����|�5=��IP���%�%q�,�?���<�z�"�ݓ�g��l�M��}g���X(�2�C�����?<7��3fΧT�q�^�K�F�8��B���@��pp��}K吓�N�9XO8���t+9uk�=k��}���Β����_���\h�l�I�o sa�����tR ��0R7���x���1��:�A�d42��#�$v���V_�=�.u��3���*�Y�]�bq��	��/S���$���������02�b$���XwN�Vi��C9m�M�"e����ӑ��ʼ'�֠ӵ����Ĩ,9��Ywk��n��?F!.YK�'�tʘ=)6֕������(U_�c�����`'�Z�}��S��i�Ɣ��y�>3��ܪ��*���[k��<�)ghJK����-�wt��$t�=�t���
��y���_�rU�fU��[� b���PW�W��:�~�~a�(Wn�#&���9��\^-ɺ���cb^�����^��>'U/�|�b�)�C�U�P��0��'�m	��Oa�o�ã؇��/��Q�߱`��	��j�7�_�E��&0SW)w+[k'��3x^\S�o�؄뒣�����ߎ٤�mp�?��`@��g�������\Y�ZrC�bğmYciw.ǡ�BC�zll��H��Z�R�F�
f��`��=��j/���e�E�(���𴕞z�
��G�d���i#�6����4#�8W-$
�r-���,�~}���X^C����ȷh>Zr��B|]@����X�0�n�L\`�$ �sǏv�
đ�גN��Q$�i�meڨ�zU��Z��+�ۑ~ �w���2���e/��3����)١:�ը��x�T�i�bu�N쾂C�G6����9\�gcfָ�N�\ɯF��eL����+����ܓ�宇�揓L��B�)c	��c�C`��5��}8@�d�Q�3(!H�=���9 ;��:}B�sߑR5��E��C�R#K*�.�ʽ~�&*�"�����bp�SwTC���7��袡�"���K�Ӕuv��y���A�
֛0�#\���G�&m:3��Z��p�s��U�;�P�0�#�0���MG�+0�S5`�	r�-l���.�ĮM�=D#"��0�p�rɁ�ⲓU	��cYH��/eR�xǖx�Z6��Ɋ)�em�!�moW��"R��E�����D%R���a�9�fL�}���b�c[�(���{��8�ݼ��%ڰ���r��[�VG[�����VU{@VJz1(89U���H9 ��c��WX���V]Y�F�:���0����y�~,c~$o5���Y��ᅉǵ����Ul��=Me}a13�P�5�~U��<[~��;*�%uj��eS�]��_�	���`����7���ǜ:�p$�{��=1�E�����¨����
Տh�h���-���Pw%�^���1��JU���8�P$���ס�<^��� y��z������(OXX�=��������nZ�³F��|��i롥�Y���ﬗN�I��5�ix�n��x �w`/8���{�܎XU-�p�����T$��'_�[�������k�ָ�t���U��S8��Zw%U�������H�:bS˩�?��l�!�~��f���g��-G���b"��=���b��e#�D�qģ�������m��g �s1)_E��{�h`���8N~�����pM9���1����❫��^H�<��f��6EB�mz��(�����,��`W��b�Ʒ*wE�m���	�E1���E�1q�р�;���<~��#xH~�}����6cFяwC�n��&Y0R��� :�2�^&��y���a~��py��l%�����+�5�2����ᴽ��di������>;��U��hP$8J@ࣁÛ���sGo�x�b��Mm��~�k�Ͽ�����iճ�O��::�r�1���a��t�q$ <'�)�X�v�U1q�M]_�F��N�I�^(=���*��v#qQ�|ɒPUO��j7$�AI)s�k@ሬ:`��l:&I�7���A�;������Z�F��%��Nܸ��1M���J=_Ώ�+���[�양�f>)�̧�oޟ:ܬד�&�\���%��$����6����|(L��c�[]4F�2C��X,��X V"�b;�}yr�/u�_��T�&��G��C#79u�pR�TY�M��"�˯ڮӡ�� �&�-���F>�0�Q϶��Y$ f�CC��?�K��%�5�Ȝ>�a��YGZ�x������\L����oڗ̆n'������
��~� BGo����Ʈ��'���Ev�����$Eϓ�X�������p/�6��^��+�u	i�Ǉj)Ž_�4�H�:g���l?E$��T�n�K_'���Q����G����v�� Vs��j�"x���јz�2-;�9���xu $�*�?q�hׂ�?�;�2�Q�34�Ÿ�6v��/�׈Ip�К�>���?����.���ݎHD��������K�o�b�L.6֮���0����Y�{B��!����К����8w� �܍�,�q~R�H7�e�<�*p�hhٌ��$n������9�)�s4���H9�� (�����L��Ӯ�gn�~���H�ʷٌ���/|n��{���h��D��Z)g}�\M y����n�p4�o@�;8��%�)��)�\��Խ��-���d�s�Ң�E�,�~ے��8��"kIb��Ae���ee���p�|�� C�}�<�O���ˆs��$+����`iN����H�:X��f쭝�f=9Л�8�)8lH����fyΆ�bdB�L?l�K�NR�0#�!���8c�1�xK{!� C�:�Q�;ؤa�`6��iqRlB��cɨ�;};�&F௒;�;�vn�c��N�;����M��g�˵@P�|�?:i(���dF4|y#l�&�h� SN�R(CA���B��ݳhk��0�Gá��d0�1s$�j��rQR�����u��Wԣ��i��S���_��Mt�>����=��mi�n�08��:;e�I�ir�����Ǵlԑ�-=�61{\� N�ԫ���qt�@CҐ��B��t�W�B�����O�O�Ud󉈲�4�hc��t�+�����U�
�jW"�؝vE�ܙ��7�P<���YT�����	�� ߱��B�^�I��t��~ �[��P���;x�ƃ2�?x��P_k�� �3�s/�D���#$c�"���^�6�D�p�BjxM��@�a�S�W�:r�_!��X������񳙷`�B:�!��qD�5�?��Fe����GHT�o�i����i��˨���C]"�:�4kD}ख़�V�\��+{�J@�CJ�P��<*���X/"�����ЍN�f���b�@/Q±�R�~,߉��q���~��S�*6�v:	"��m���rŒ���E��Џ�}�� w���l�3چ�:T�|���%ɲ�oK������F�]XiJ��,&T��t��E��I<5*F*rP��<
"�Q2=�劅S!���$�����i��!�SN����Ü��M�ew����`���-Vo{�1�NdsM��=$��QX��J��T���ơ��EN���� ��nI_)���_!x��@d���+���|����O2�j��S�o.3)W	�R� ��"!���iP��G(=�@2Ԁ.2�_Ϫ�2���+}�2�Zhݪ,����{�����tZ�^!��0�ܖ��qġ{�U�Rf��J_1�E��i�y��Xc�c�tu�ߓr�|ڷ;��}�^�9�83�5�a-�z�?9����<y<44�	�����A:�� >2. F#d���)q��L��N�&����P���P��C�}N�QW�����-q���,t�������ec��I� %����)�3�*z(OD?�rϫ��Y�jcC�q���U�����m�8y5��7�U51�t���H)@8[� ?:��W�����eD8�{�7�J |�Մ��ײߦ��GFZ>ӳe�����c9���>��Ll��m�eD�뽛��m�_� ����_�ûWc$L^_��p�X06B��$�܈�0���
��vbڹuM0���?���B���	J�#oVq������߶�zݘ�Zw��	O�iQ�;�Fz�0^ı��C����t�Q���f�#(n��oK�#�Q�SDB�j�K��ZF�;��r���_1�_\������WO�Ro����ç�S9M&����R�P�_��ԽE`�3r�T�=x��	�J��\Et����bW�Il��I�FN|����(r�6v�/$�QPU��d����FI6���x9�uҚD܆\D<��ј�7�8��e[�$`0į���&�-1�O6[ҭ�(�v4?kG��wu˭��G�N���w����C��*C�ǧ�C�����v*����G8�h�oe��Ye������X��Ei��Q����\Cp���a�����?E���*"��_���x����;�0�T���ԏ@�TCR����X�l-~��=��>B���u9��8�:�\�ڛ��bx��n���#�1�D):��~l��|RǢ�ؘ���ifN�N��w���&ǖg^b�����3�J5��"E��S`MU�YF|W n�����e3!��o�Wo[�=�C>-���:۝ �u-#
���Y�pI�u�Dν��[
tz��R��[���/���g�k��Vt�L�*z�ފc��y���C�Rb!4�n��wp�@w����(�@�)���VZHZ��"+���� �}�PQozF$��ޝ�f���JS�:�k��08-pM0�|Tc	1���P��[]�����ǣl����r� �����]p΅���Rv��e�{U��ƻ�5�O�c
$^@�/L��ޏб�I8^��H��1�A�fz�����F����l��fٗ悽$+J?"bR]l��T6����9��osZ<*��A��skEHDuޢ9>Ƣ��K[���Xy��9ފj�^�f-��L�Fi �!�"v�6^E?m����]r��6[τ(F� ��z�J�b�1Qc`�u;���Ԛ�S��ˋ$d\Q�6S�)3�?o�Ѱ`BbϦ�+� `��v�BS�%�*�s�m��,�t���{8. � ��[lp:l���^���� ~f"p��*�#Yŉ}�U/�:ʡ��jQ�.�lخQ�K�|�,�MWH�����<+�S�cl��Ʉ������+�� Y3~�嗼���0�лRt�-�w'�_�C���fs�
BtSh����Oߪ���j0f�g�&�YQ�3�
ˈ��;��.��-����x"�Y_ߚ#7;OQ�a��w[)��o����w�cl
7��2%����M�jd�N`o�J���|��w1m�h���o��?b�A� 
�_���V.yB �l�Q+��M�rey�^3x���\�F+��H�gx�K|�U_nF'�.����!�������W?���cB3�s�����HP@*�D�&���2�Pb�iq��� �Z����/rm��J�XY:�yǰ�ţ,ۇO�u�����O$*�Ĥޡr�	P�#Z{�D�H3�L7�K��@96���Lo�J��̒BVz�{�F���?&1�����h5dr2��T�q9�k-���"[u*h3�[��=�&M�袋�r���_���i>���e�5��h�����^&�� .3_>�h�S>�=	gյ���%���|*K����G�������Y*]j={�L7%���~��沪#Z�'�:�ܘ����b��/�r��9���Qڊ����˟����V�'�#^�9)q��U��=��w�d֒8�ƛ�;b~��T)a����3��t�9�,�&��E��b�-���xRL�ǯ�?&}�}b�0�)9�A̲{�3roaǍa��<��hC�%rcoT�A���}�s(jp�8���1C,�|�.���hd;���6&�ItL���D��\V�TA��d����)�#?Lu�e��f�}�bkxtr�mdF%4H�y�1�n��v ��wYY.�^ ����o���:�h�Z�,%X�� �|���k��A@��ǅ�Wl0ƽb�l�'���*|�9�6�i���
Kb�a633�r���p����9�:�N�5"���)m�Н��uꂖ�U�f��ߘ\�H��1��P�Bi:4��"��C�=��:��j�{?��b�N0H4 �__�3#�ګ�R�����52P5s&Iu�<�gnP��RDxc(r��/έ���Ry�ü��t�O>W(h }���[v�������߷OG״�� ����be[�|��[�q����
B�LG����@�K#<�)��^�2���V_S���;$-"��GE��l�p��ZA�������X���*��]���@A0�C�:�3�@00��@�y����*�6}�"�#O�-�~,D�%_%�vH�z����'�;f؎�~F6p�R�g�C��'v���0��J��\�bg���lИ��Oq#о��ƚ����~_���DV�|���� ��i�j�פ'���%�1�
x��֌��q� 1i��"�*���!7=pv|�p��#(1���i��g-�qi��E\��ש����$��8H�2:�s��O�
yy��/��E���s#��.�.�U�i�G'k2��&F[�"�S+@�>��U�dj�`;�D��n��� 1��B�,I���ENH�Q,O�1Ⱦ�"�:��Ks G����p������!���m�K>�Ի���~ˇk���
T�Y�y����/��<߃_O�V���ד��=��J���(�j�A�x���HY�����}��]f�s�8;׊�'��Q�V��R4��E��t�S��*��s�i��}J�l��e��ۀu����%g����'3�#�!�g�����p~'~l�9]�1�:�@*b�3������ Q��|߳OfI�4��>.�G,9T3<@�)���3�8�~@T�	!��Ek^`"�;�����f�d�, =�A}0U�I���ˉ����R��/���V�ò-y���֡�L�F�1t�Ӧ�3��l��� =GN�����N�=��,oD�� �Z>��+�P��(���	�0�C������X����B�5cn�;'D,���B롕���S�Ю����+���#�Z a�uX�\�fJ-��n,���U�֣:��siV��j
��"a��@SI� �t_lŜ�.�s(\<֠떢�fAXxA�}�}P�=��<������H�O�)���L��ik���2���Լf�k���w�p��zni�5<���p2�ٛ�G�Ql96���U:�Ӫ�TcI�R�_/0ra�,Q�.�JL�/�H�ǋ�0��Za^�_�i��!���ߓRˋ4�JjI7Z1<�F��I���������iM�N�f�E)e���*�S2 V��_����z8�@;���pI���A~����z���%qYe17�������q>���z:�:����	x���&�*-��Ή��;�%^+�L�]~ѢB� #.�P��(�9���sѓX4�EPWI�1[/�SD��u����%#��2�ڔ�Q�����ﭓG��@�㬏��� yyX�>L�	�v�B�R��l�+H��L����tc3���q�������/@����ٖ9|5� �H��"^��c�{����֏Q��i���z��A��/PBB\
����Ԍ�~;J5��f� &�{�����	�\��`��@|N���SbP��z4��=W�#_����_�D;�ؘ]�L�Ƈr���y+X���\D����\�w���Q����F�[�K��^o2Ub��'��6#������ȼө�0��xA8��?�����Y
1'�h2��Q���5��cd�	�P&�7�^y��0��q��`�/������ #�W'EԴ"�.����ft�!h�z:n���8�f00l�X�TҸ�ΩK�9�Zo��W��,�m�s��p�m�̿������[TA�GA����U�`�j����|��v�~*��y-»�� ����w\by�ɣ˻C�*�{R"�Ynd 1I�����w
�TTP���x�02����H� �3*�C��F�lqr��t�
�5qw�ㄠ�^� oD�hbq(�Y}�l��N���4�V*�,�A�Q�anv^���7?�_��GJ�Iq��>+������q�N���bw��9�$'�ի���yt�͙�ĩ�����ew}���A��6H=T]*��,O�Ӷ�u �0�
~�e/T��m[�m�`�%k��������=��K�
�:EɄ�ਂ/�& ǥb4M}����~�:��S,P�ev׍
���B�Ƥ���#]$;�����%�_�(�W^��.����g��-�<�l�5�д����H5p�iG�1����:�E��>Z��(��5j$��3�:C
����'�����n��T��� Y�{�I[K�y|��O����*h%�kۻ���|��m+!c�X���ǒ�N�ؓx���s��Jm}�P��G_���e�)D.q�����"1W���X�I͂F#�Y�&ʥ���q���y��J���ϲ�'���L���!v<8>��Ƨ�=*�śP�殑��B1ɉ �z6'��C�
Vj\33��N�Fae�2�����t�Je��[%7�Z�Ԅ�7�9�%#������׏yz�Y\{"ў������f,�t]���#a�уPN9�mI�J�co��J�6=�z7�htC)��m��o�Ӛ��e�'�����Z0�J�q���>Q7���h�T�9������$1bG�?;:�c������!�9�>{����l��ǡ�"I�,j�l7DaR&���U-w���#k(� jo-�����Mۈ�߲�Q�Y�����#��Z�ۺ�����R�����Tm��B�M���@�w_�á�ah��{p<�)���2~XD�n߹:���wTŜk�]�h|�w�:��Q}=`��܅��-)��U�n����Ɯg�i��Yՠ�s
�-���`�m΍�f@1��Nt�{6%�U�|?�7x�"�LӺ���;���w�4�
���i�ę��Q����T���X��M	�GF�q�k�(#�Je4��U��{����H�h�lόt	U��@���ys�/�+�*�J8�Y�O2��O�eϼt"2Vo�Y�J��Z��שqq/l��:��A2��]�`����k�_���Ei�1���q��].��a�g��o��E6)�4��Z�}4i
q���T�j���$�Xl�K�@���l�o)�<#Ǒ�p�jc�'�r���r�B���1�(��]��Pt�+�6�Յx�%�����1�����T0R�����v�Yy����Zmg���z��t��_x�qS`u9����[��I�׸٨ܱ�<f�����kY8xFM[�E/�̙8�}����q�\!��o6��r�$y�I�5ps�s�7�ǘ�៬�o�>���X�����-�x�Vj������ԐPu����b��ty��p��=���X��kw��*E���jQfI2�:eJ�l�_E�Nц����z��$�s$�e��_�DꗵP�m(��HlJ#�k�T���[\�2*i-'���;]���]`��f�#�����,�X ,P�c��[,�Y5_yz�v�16�9=I�H)�:�dn�c���OuGS��e	H�`��T�S���oM���KɈRx�M��Y:l��_u}Z��8���=�Te=E�Y�6bwj����Nx�t��|-B�_�A��|�*C���E=σ��P���U�������g@�d����� ����E Y����%�4�.�1Ҋq��~L�X���*Q�)��f���
�n�Y$���+�湈���]ǚO��&��|���8�ݟw�7"�l5J��ލ׬d>�'��К���ޢL0�9e�T���nMD����F�$�S�w��-Ҝ�/]�۵P�<�n�+��G*���06t�D��Qb�ZW_����w �����p����*�G�n�%u���^���;"	~�Ui!���O�V�=��8B��w����%�D`W�=��0	�I�Hjs��rW��o\�w����*��� C�q)��
fb���kH��r�Q�f�Əc�����Nb�k^^�>�"�`Se���0Et8?=/~��ԓ���N�7�p�6�BT�.��Hg"�?��b,�%/��(�����L�tܷ|MOh�s�h��U<?;��h�Nږ�{B:4>�,�����o}��4cA!�^ܴ�����ےB�n����\+�s���V�Ϳ4�5�KE%���Hgt&���!���|�������Hi�b��1$Mo��U����w���j��������(	�wA1�Y�-i��]���}�"�avkt����l��4d <*n�b�M,K&��gDbQ�O�(V��2�V�X�Ɠ�45:T,*Ԭ��r��Wb{�4����F+�<!�3�y�Zibfk.��*�S��.R���C�ñ� ���{���>�Y.c&�%���ʁ.X5�ܦ�@�<��Le����CT�b7([P�@{e�~ECrq�j��w����<-!QS�p�<���_����|*�?ǖ�U���)���eqWd�ǢG����I��i�'p�ոq5q.��V�����d6̇�~F�J�v�:??yxF����z	�0�^8�D���q��g�V�I�E:X9OwzO�}�N
Rݬ�?����#��L|��ˀ�XnNW���r��ු?Hf9`-{�=�\�x�9�z�t.f坙8O�b��`�k8�(�zR���{QF�(\���),7g�/��C9��.�DB��ܹ2�C:��κC:����0�H�ꋹ���Ҩz�>�B(���4E��B�8l�H��k�\���=���85�dX۷�x׳��g�x�܉}��I4��-�k��-�W���Yц��e����[�U1�Df�+=��,�Jk���m�V���?<�i��ZD�B��Ct׃��J��!,B,9���Q��V�2:s�Ã�_����y!�� �����U�珷���ac|�����~<"PP�(!�>ۅ�~=�SNey躷�n�7Pf=��	q��v� "��C�,[~�N�h�"�)^D��6҅��;���X��Ս�Yb�d6h�m�T$pY�@�ן�9{>�2�^T%�q.��kZ�R�¸7�/���,���F�`g)>��F����-��� iU��s���^L���2��-P<�'6���C?^��+}����5X��~���s�dn��h[��/vN�:̠,���C�5;v��9<V�˲��������5��C�BM7+��Y0��S�'j�N�ժ�PA��T[ Q�`��ư�u��CK�u�5B����ޭ�<ߵ :nguE$Ga߹�8)���Hd�"~s���L��T7lAT䈀3��3�Jɛ3d���NM����Fxqx6��d(`w���.$c;�1���I+c.ԯE�� ��}y��c��W��>���A/]uy�G�?!}$KG�� ~����{�3������qκ���t��!goljV/W��`���y��j�w���0��/dRo�o׻�8����-��#��B�7���1I��ך����p*C�4�O�*��8��������H�i�x|�\D~�,u�GY�>��иwAd����X��V)�k��H�Oy�+$$N'�t��dj�q�>�i)xBn)����m�~Zx ���Qߵ��j�wǎ'����2l�cY�`��uW'{& po����Q��}԰n��z�2�k?��-Q��[2t�߅Z�ŗ.=���r�e�jG(���#~T�2#�l���Օ�FM<:i!h`���
�i����=/�E��L�1���B~́���(��ew����a̭�]�����6�к�j��l���b���8�ێ{ �X�)��}�C���<��D������?sBk���w��ˀ��V�3���%-�{�n��4i�sz�Zn��)�sY�x�
�`h6�[��L�׬2#U����sc1�%�y����8�y7_tOU��H���/*��7��� �*�3n!"���"���'��b:��� 5����"�,=�r�Q�k�n$T�W��r�k�J�f���>� `�!5[<	�o��oe�J�Q	��}�܇'��U.�DM�[��L�shG��F���7zLl�CS���n�	Fq)�GAd\?n���
4ٛ}�A]p�lą܈���q%Q��3�n�!��&�����������g���.�Q�p���q�+%1��~�.�,��C��Φ?0�U��	U$|����F�M�9��~o�����ZJ�g%m���C�f�xOO�zf���EN#������kL1\D�+%�1�I��p���ט�h�}n$���ݓ�����Rq'�����&Xz�[?U�Yw�pr݋ʎ�S6�Y���2k��l�wں�kh��v�H5`�͂�PH=-��+�v�a?:6�D�.�B=�(ha�L1����Ez�܍�d�K}��4!������,=Tu߅R�pLn�T��V�U|��Rt� �T�y@�;7rd������ī�q�@����ưW�� ��nD��T�j���i��U�/+(��[�Z�9�</����0���z�2[�L�1����`�00	�T��Z��/a�8�9�7^�9���k�-��+%9���y������i��ϱ���Q��f�h�o���q�9e��Dk;	ʵ0�E����R���;�S̾�-�r�E�0��6~PFz�	����]�1��0��
�/�u!���8��Pj�����ÍN*q����6���x�և0U�־�J�ܼ\ @^�#l�w�O$|�Ui�������s���W>pxF����Ȅ�Rڀ�����=��� ��I��؇l���w]���+~�9�;R8ވ�*�u���� -Ҡ�n�D�EPnv��S-�w(�UU� +�%=�������o3k��Ӿ�T�-x%�����wd.K�c���K���)k�5/�Մ���y_`�[�s��b����Za����ǥ���7>x�E����ی������[n(�"p@�獐Σs�\�9Mj�s] h�ऑ�NLN%/P�{���F�� �Q{8\�$�8f��q�������"
O��Q�GW��2A���=0��Ä�#�ω@�����"i8[��뼪����g�Js��8�נ������s\qT[l�<�?�+�x������i�_��0]�oI�)��m� �`ky���w�HvAo$���&׷&nWc�SV�ez�{O�ܫ���_ޥ?���YT~�q���l���л�gD]����Q:M��a���ɠ�I��	2N�(aI�0��Uم0q�����ƾ�0M�����Uh^L���㈺����@��ƶAZg��$�rO �XA'}�z��Ä$js�KѰ����@�����9���;b�6]+l��x��J%>Ê �c��;'ը��m=�TY܀��]�|�V��� ����S|�6I�9�3O��]/nd]��x�E@�3+�0Wp򧪭5gX�/������R��&���m���4�����:�@ ��Ga��|D�'�Y�8����B�f�%3�&1��l��@�2������0�N	.2!���K#t�2�HEQw�c�[W��YA���������󒩑ȓ?�K�}�1�Yn��	1���S�(��Gn<��!:#`�z޼S��ř�!nI�� ^��A=���lU(Ց�"�2O休,Sg�����������U%_#9ؕ�U���@]�R���sȥ�5��V+KΉij��--e��j��ϚWo����7�E"a(�2�b*7Ol�½�8�}�>3�h��-�������G��Ǜ\�_Cj�ݐ��1�D��Ԡ�΄NP.�C$� 6�:�A��P)z]��zh��Ѽ�}Py�F�����H.��9ճt�o�Z[��~G��'}�b�ўP�-���x~�B�z!6˱�j�][�3 ����$�;�E+d`(�6���'�*Yg��I�S�khsen����9��]�n�A�[b�Q�{�?�2^����/���E��+L��L�g�8�;Ý��L�*(��;ʕ�	j7�kȁ�NG��V�9�)�u7�0�}� �S�&������aRI�S�~e��Yfc��ɔuL��'D�@��>�m0#�w/om\��e��*��^X�}��!�F��&XAd�Qt���}���/v���R&�Ε2�gA��m�U��QzR��6 
D��`����xf"��QK�NӃ" ̬��>G�Ȧj�42�G�����n6)w@l��7�yͣln�����AS����*� 7�����*5=�vŸ���T3��������ؤ��IՇ�F���,b�N��-�'{����]��ft�����qz+����c�M+p=����z�ē{!G���S,�N��k"��a��v�L@���9E%�]��Y0^�$�j�*7���}ڕ��)~e���V)O��C�[�k Sb�;��}���8�E��֪Q�D��@�yX��iL?ɉ��34=�{�(��,9!�Z�eE�I��~��N���iR�&��@���u-?�G��HWSh�og�~���h@`�m����R���馓�hG�U��\_�6�Ⴊ|<껤�*;p��u>^��/.����,x�OC2BcJbꥠK��9�LR9l���=��NN砈�=T�ґ�=�J	��������~�]m{;7Nh	�#�p�T(]������<-�S+��ǅ��,�Cs7�,Yv���%����ea�S1*�I�-�����=�hP��͇�~@d�ɯ�E����Wr�H2�P�2��č��o��|�N<�[*���~��PԵc�К�;g�V��P��]��9�Ze+gov�R�\%`��Ԛ>ˡ���v���un��������ʼrr�w��fRx�w�N>������'0�y�LϽB�sM�[X�z�W_+��>�深�Y!��y3�>�$7���-]'ӷ&}�N���r�&g7W!NR�V�NCzW:���I�F°h�����ᑎ��6�k�_��i�P÷�{^e��+�f3�(�y� +���?�����`T�!޵�b�K�t
�� �-��m������o��U���Ku��ޛx�'@�L�q����u������t�-����D���=�{N�E��n덌4$�l�4	f�T'�k�dpA��A��: ��X�tZ�;&�`�ں��l�q����M�����՘���se���6�M�l�C�H���)�LaW\�����E�s�8��WT�H�&(��6���\+���$}6���M)���ܱ�,m`���'�JF���x9��3�:�ڈ󈚰X�;>>ϥzj��jb��R�
*Jgn��o(p2�0}`�"y�];r�90ǡ��8����CU�� 7Oפ^,�?΍�I�
{�W�����d�_�XQF�Z2y>��v[m�׈� ��B�[����Ctr�U�"�����0l�ғ���֢�2��`iMʊC��x)���U�����R�>B7��8!���B�ܵd
��D�F͎�SR<v���Q��L�[����.��s��-����-�"�R����H�ɤuuȑ���b�@'~r��K�j�2q-gl�l6�$��S/�~�:[u���\Lq�k��@s����F�� #��I��#���3�����x��Q5v�X��d�!Մ"��5;`le/9]	c����
W\0�J9U���	��\n܎lن�P��(X�X���H���>>/G\�E��	[�\����%��Ƣ�b���m$�%�I�YXPr���_I�]�f��XH��H���>eX���ˈ2��r��:y.�B�v��I�Ӆ�M�c���a�Nv.��V���C/�>G1��:"ը�m%��/�C��_{�y<�6�?|xh�+�~��w��΁]��\&%��M�o�*��O���U���!����&���Q�0(�ZW�����H���r�2���;�z\��eF1�T�<X��|��l������6���8�2ޛ�$lS������_1��w
���5���Z����T1��v΋2�H-Hց��Ѝ-������/0� �g{ F��H	нv�%��*o��J��!T���H��04�u���<?GV�۟�܋A��=���1�����_�VSG��:\rB�iO����6f�'#�8x\s����%�w��y�(jA2t�Y��f���C �c�T��3հ��9�̬F7s`ҿ��^r_>���k��'/Y:�@��5aj*�u���Ʉ��~ZqdMZKG̶�.�{S~I|-6՜�F�P�1vG��xı��+n����2�{7K%O��)x�A�������q^�N��{���Gq\�d��g���l����@�nă���'V.��I��w��+�����QA�~c���~>NuQI����-�i�����q���KXJ|M����i�����|����U��8ՓR�\߶xXA͋���2�W �ă�!卝��z'��������3�+s���w�'g"�*�=���U�W��	���˯��}+��mhN�ZH-��g]}ƶ(���;�ޖݓ6q1����]�!�l�4հ���X�O߽3����ZD��ʲ4����l�9��,D�"v�	�����x������z���#�Ƙ�K)�B�ڔ�e��,�M��`���?L.�Z�=��Ɉ;���Gh�KALK}�oD{���7<�ԫ�oj5��ĘJ�6�P/E�R�����C,*PK-�j�Fi*��7���)z±̺d���i�잉T4�p���^�|�޲EZ�+A�:���F�f��q�kS��N�́�����]R����l|o��;"sP��s:C��Rg��vk���rS����Z4$pr�v] �M����щ����Ӣ�){
ȋ�E3��-�}��%"`~�y8~���y�K�q�v<�8�@zݣ�� ��S���muqs�/efsSk���&	������S�ؓEr/!�bI�%eFk���H��7�:��g6#~�թ�sg�w�&)����sF�Ý�lÛD�܆h���1?���;)��][��i'F�F*T8��}���0���`kr�4���ʮ�ڦ�0�CH,Z���]ww���"3�u�eP`�C�(���G��R9�XF�:�C��2g�2@�����r	@"}
ǲx�ث��/��W�`����ˡl)��5�߃���w/�`?V�N�*������Ⱥ0�&����	�������������7� �uH��}�O�����)&��?Z�Bl�} ��滷�a|ݞ˾�\cs���j�' ��8���,��z��h.X�I�k�Ek_g^k� �͛JǓ1���˜�rѬ��Zk�� �-O`���-���8t�o����8���E���5�=�k1�5HK0hsG18w���N�ڇl��!KVZ��Z�".�2�r�o4�0�y��T�#���K���B�_Tt�:_�ؗ���������ޏkD�T�`���Ɣ�g��{U��ҽu�T2lꇆ�����+dԙV�-���޷>@ݲw��Q�r�uh��r DĦ�TX�����/���1�LZ����WG���aE_*���#�KFj�ra^v����ыe'�Nq��kL�͗S�Oǡ*]c
�%?�}��O��qxg���ը�A��[SZ8��ޑ�ƓՉ95{1�k�W�q�7H����̰s95�J�t�'�e[T���:'z�+y3�&25^�~pH�o�J=���Pt�I9��\�J~����1���� C ~r��
Z��ƌ��\&���v5*����Ӯ�i��	J����r+�9� 6���P�������8��\JA�(/���z{V	�C� =��iAR�ԥ
j��ح����u�׊t��"���|���]�NT[/Jk�S��UU�\���B$a�5�A�](�ت/ƔPVa-ӂR���V�)��P�vJ ��Z|:�%Y֘��?�-l5�5�JJ��WG�=�	�ʾ�A�#NB՝T��P :�:f%�z卄~M��D�w�Ǝڌ?gG�V�[Ө�	*2�	ݰ���m���[(��o!��+��O5�ۭZ�f̃�`�0��ό�y�r�<����� �����C��{{��@�O���]�US��� �S!����B��u9���ᰍ�l�B��3�m��"�kQ�s��x2�{����-�6��T�m���n� ��)3y��_YMM�{��"�L��s3	�lc�e~{�5e�8�Huc�y%�x½�_Ԟu��	��>f���1V��m���%�	_��`�
=�R#���ZIS�iL��tp�1�G?�GƵ�xf��^hP�h�?�ؔ����f�+��-b�>�~ �@w��ăj��~�<�GZ�Ǥ\����s�L��bi͒�y�8��P��K@]�������zE'�r�*��t*)��QB{z�+S�z��y��
�X�47r=3��7�b���t�Bo|��5]�}�wD]���cL���Jr�gԼ1�����D�ה�<����zJ��v�5�\�5�.�����`��숮?<� ��տv0�Rzh^P|�:��������}�)����A�z�x�b�wtUО9g*�^�yP�1�M�=�Aj)i0�r/�'%��\6��Q�;*���At�=Ŧ��t~��6�� ��� �YǠ�Q �^Y��Ms�DcM*�������B��ĉe����Zt�, �#�!w�D����q�;�cy�*�t9�N�b��[�;x�:Z|�D]�g��Q3[D��^����|�O�� J~_2-�����FZO����S�J���R��'(ļ��z?K@>t��%��K�6����7`4.��|�4�:/��l Oo�p֝:���� �7͞Mr����i6�w��;�m�1bܝc���%�s�E��L�\�_Y�?�s��ZW�A�1���(Q�������5b��&]�>3��o��������1�yY�n��=��*�P�]�v�5�
�p��ICd	��[e�߷p�t��9s%.{:msR�| �SE�Gg�W������y�>��Lψ�{�]5���:���` ����\i��ۑ_��Z�ĕ2��t�Y���pU�gUz9xt��M�q^�܎?�[�K}=�;4��?��PuG�Ѵ
,av�Z>?�n?%�ׄtfb��UXv���͘4Q��u�ٖu�G3�_�UA�P�B�˹_���Oͤ�� ߫~�"�ܐ�;��Ď�� �|��7��R]����Ho٪�ԖTJGʜ���T���o��)�겁�:�XU_;���������`�2 ���sN���:Y����1�@��������y9�h��־}e����6<��ǿ��Z�%���^�OuH��a�� -x'���^?t!�+)��^���\r�P}��З5P��Z��$�a�d-��հ%��!��ğ�ݟ�������%*�D"v��HD�	юw�p�p�F$�ZZ٢�O@��t!d����׊�\�4
���Wh���%��W:��d,��p g� ��r0����߆�����܉�B<sP6��4�IL��z�ջ�^��tOq��)iȔ�w)�`-���W.<TV8��Į�:�f�C�2�|��XϜ�V��_�u���<�}bݦ���a4�ӧ*�7�T.���6|O���c��M�|�%��W*)L�"<��ѿ�5�L�) �K[�3�Z�����B��o�&,���+9��3F�L9?�o�&!�Zb�`wz��kPr2$|��]�C".p����%$�OWfշ���c8P��t�	�j����J����w�&�`�}R����/�7�m�fOKPyV����j��a-O������m<F3���b4N��6�JE1�Mkt�(�A��Jy�XahH�ÄM����䣵�lW߭Օ_.^�WFt�0�	�&/��
��S|�i{��C���֝��u\r����s%kh�|\ ��gJ��ǖ�d���������WO�J�t�����ӫK��u����i��b>��5.����N�5�@�`n����*��݄d��Ҭ�Q/(�Xos2%t{Vd@��J��j����D��6�ߤg&�t8�g���z_u���9����H%Ic�8,�����(kK^�Lp=��&�GQ}�M���oT�q�PA�v�
��p~��8�1�ry�����~�%�Dv����E��5�S�'���@����>іd���(́�AW�'�pA�w0`d�x������1���ۊ�"�򯰱�x�����q�cU�o�,Zu���Ƞ��w:Wvm������X�i>t�P�Uأ����������o�bRgz��y,D�1z����(ڕ�	�-`g�a��Lɨti��,)������6�D�}�񳹋4�kRyBc�IV:�A+���ʝ)��C���Kg?=��毫�d���U�	�bQ3���m,�ea����]�����yI����c�-��ߔy�FȳM�B-�����<~E��g���W�;�L�jA���ə|J^��*�dT��� �[���.p>��ے'��ڒ�j���C#l#tL�d���PV�
��Y5��H<5����U������l�����I+�G���Y�[~���=��I$<���k�Q0mhj�Wfe���HC���ݯP{�{�Ŏ��R�:�o��NR�\�px�O_���g�[?	2�p�ٟ1Τ�s�������A��u�#6i���\(TtE޴�_�l�v�
a�C*�5���A��(?�Z�K����y`�"ٍ������(�y����N�Zd��o���n�I���(5�=^Djl��ޔ�G%W�G�%	T9�ɈK���-�h�bKg6u�I��{���:7'l�Y��i�/-G�-��K�5�?Z��lsGa ���죿(A��JX	3�q�������K	� \~�t��y��M��iYW�EM�C�J�4���B����r�����dSE9=cՖ�s2��+};7�D�F H�GF�jJ7�d��&���Ilʉ��������	U�0i��z�x��ۮ;�g֐��XJd�i� zz�Kw[ �Y����k�����yoLd�`�͚�|�7����,�+N�j���w]�.bxQ7��I���O���#�
S"[���s��PY��Y����q�K�a�j5!�{�6
!��T�?�,� ��m5��&���N�O�>�� �0k��\��/�V^qA�}�g��Ji��LOtb"������h���ƚ��5�UϿG���uH��Ӧ�ͱu0Th�u��������>�i��[�H���y:MA��Ϫh�i���ܪe�=��ʥ��KI^��!�,&g�~��c,�ny�請���13c� �`��L�밒��>�E5�3Y.q�	:F$+��M�(��z�d���V]���i'��\ '����vPb�1�����
-Y:8E��hf�o�����2�旋j��[|���\^!a��Q+�vҕ�X�[ I
�Tͤ�ol���Z�vqL;��<n=.�<�W5��(�,����C��/��i==zt�d�bә�!OQÛ�3���Mi��4����9S{���I��ҩ�w�CK��u �Ց63@pRO�g�uo;Y��6c4 ���
�:�(P���v%b�1�G߲����8�GP��c�qUH�L_�����p8�� ���gR4���
0���>$�n&<I0R��!4֒r�F�6�z���
����	��b&~}[��k �:XB���`�s�2��X����e�:�ld0l���E:]�cԚ*�>t^��d��(Q��mL�0�T���I/؄@4�ً=��%5�%������l���sܑ�֙XV�QT�l����Y0 :��0���"a|'q�����=�R>���I�KB�G��-5G��_����* ��괅k����m�