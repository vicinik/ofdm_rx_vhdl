-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
D5nKrEGsP59apL/iab1wlWKoiTxh8ULtZo3P/jr4dvbI+8WM3PiuGZgbWYSYIG41L4c+SwxAmxXk
hIrCAslfA1g1Gn1vDrO5Z+7UuzT2XnRwZ6nPmNTs/yoIYp4sh7S2tObSGztJ6kt8LnD6SxzWo25M
ia5aBZyvgJIZOrhd9GgX7wSdeG16v5S1OCehA0tdc/+WMTTsOCQrlx2qyjatMm0sasx4HbMhVUtF
QeHRJn8TwyrW8SZ9AI6UKz40Bc2S+Hmog3a1tOLNQp7JYAUxV/yAXfETK0F9yJ5ffbJb9X07Njg+
1PDFJ6uAhxJ5EBWjzS6r50Gtbf29rgWMEAR92w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35728)
`protect data_block
VrG0lubRmW05lIwtGp/fuhb1W29XmcyLCjgdjkGcJ92XaCQLlfVNQB79+SSWu5Vl8qnRSlXdNbaq
MeeabkZ7trhP5YztIqdwNA1WG7B1oA+WBMCB16IZ7XxDf/4cyyC7W5l4SowUy0JCs36Mmzdakz2W
WsNaI9TOjXAGOqwzmtW98FBYGvzb1tp5IMcYRIMZXtvYr+7q5QzHZ4JvjEcTASPf8csPSFU7HPfE
Y/a24cy/pK+dVprLFe1PQdx9167tfaB3oORPaJ9oWnZ7hnbZ+j2Q5U8rDKXkJZtTfdob416JipkN
/B1GaWWvqVUpu4fNjy8GKLi1UbkCr1Z6U5M0xv2NvS6nfI76wqyRtB9cxPTR4aEhCIqJzBE+P0z0
/Egs50TFGh4XHkXKpMTirU7NdnLrHdpqTG+yhv5bk/e1+muGiN05f55jonCl7z833MR4pNg7f1s9
tC10uz/EMs18yBtGTKhqwOi1XiZh2/oV04eeVKAVQ5qRjIMMdLsSddiKpZonhD9HerZcHyxn08t7
/BEMepT55ioW+jRs/xXO7OYYr6q/q+5ZNKFcYbamwrhu7H9QI+dS+RYXvwAQS914nqmb1cqmVI4e
/WbhSuP4Qs01QeeIACTkEACir/WYrFnb/Q31kVDV+ZSrzNMp2XWPKHdeAP7Aydnuoxb9xEbrUvJ9
L4l5Tv5YKfXeGawQTqBxsXESm0tyOepcjUDRlOGuOJqZaOhxGT/bH1Ja0IqgIY/RqWWGMuFBKTj7
yqOMgYZBwH5SjZcfwPJha3ghdGOlRT2pdS/gpaNqKzQNwA8z86CTJi+jRKC2LOmV7HUJTfMQkreU
yIWRonPvYVSQEBwBghJ8oMMWpfOhs5zglSc0DU0jxMJQif+QwwdN0beDvtgvOGDl03AuvwW7qPej
p0xprDXHO0wXujD9a0DH61JDO3+5zRhfBPz0e5C9e+/lSb2xBJibyBUkU5d+iPZsooaiHMku5m3n
TRUi8E1m+0aFBhuvJam7nhYyh+ugjabW4wVP7C5H5OEGF4EetzPj+6U4g/1RzCeAgMnMe0+xvTmL
6SCkOrNuz2BD8GLcZAYKiIsgmUZ43yAx1u6zqJfS37rDUKQiuaR46ux1wHg5aMQyoAhpEnvZwMci
50WNKxVHdpfC/289hzLr9S6UZrMGYTbYipT3f+GHpDZQ1jByFz46dyVosDsSJgxD1DjIEXXeZOOV
VP8D0WK/rqju7yUsxOCMCQV2mtq/V6c641m5GdiVnJ2ZUD3KCg5G3fLJZ9V7oq9HVe807/+WZeDu
DagyWscQ76nW1amVqADQySsZ5ITSTu0m3ibJMmJDr8qtp79HxdePbspheklEC1a3RL7QCzucnZEj
RP3r0QqGA5OUPuXBciKEMZVaZjqzQpItwohbe6o4+SwsvXqPRewpftZ8ZLTNSFqjKQWDuhoxQlsc
K9i/YJ5CTIa+zblTz4BYTGqoFez8VTafiP1wy+O6H/tCwvg7nFF1n1BLK2xb3l3MBJsQfen0v+H0
qF6gQ+em1wvDMAsjZWKXspkG9tkxLZ/EOxYYSfvH7F9fgVuEgnbYKhJBrMARU87+AJAHEOUlB/8B
thH/uS6FD49+TtG2Ayux5xqYz5Ef/HDb1C4ThZDK8yqCWL8cZQC7en1z0R6nFw6pc9CnNgQMF8jB
5pVuwC2Cka8WeLUgF0rKRu5uJyuw62HnLFlNX6vrwSLryCYzvf2DkX6sh0D0u1RAzNBMlm+dwBZq
ECaMPb0k2iTvqO/O65IhQuA+ot7IrbkcqjGJOIAhivdoN7b3GqR47uaJoHrHkQ7w53eL7qDUc/gn
ZZAXbpfdaBC3jyKAqEyR00crXH5zKQN//F0TNBEIHLOmjp8BNrW1N20iPZi8FouCx6jktW1kO5Fy
kPpl2FUScbnLVPo2x516l46+IMtet5WF6Z67Z2wmemr1TwcaESY3bTARbdp8hHWKXv+xXkB2Qdn+
m7Y5J/8ZdOio2OqnsLxp4zBBc4cRhhUVQ+d75SSeVIhk2a/S3/WQ5T7xU473lAu5D1rtR7Io0ooM
Quao5+evuTJlY8zIYOvNiOD0QWdtZtlFW9FZm32qxx8P75K5WZu3gWpOwU7zlK+hU3xmmxdvk+0O
LXJr9x5KmjKWWkTvmg4HTIXefpQEX+1DBkGfb5PhiYN+MDBySLW9K9LXzVXYhrrN7DVL5HUJz87z
Oe2VgPYX3zx4dTByn1RpQrjV1hoIKV+zlQL3l/T1qVz/PQvgV7zGlQyEXKPQniLT6BHucMTyZMiw
NtAjaKY0reAkUDk33HyHVhnuOLtVi6PSYJ7hnfqzqOT4nFnJeZdYuM9Ny4edus1qs1Q3Ld3B9PIj
S0e+qV9R2nd02Trd0cXfsXVH+/1/S5+GEslJxcPn8ukQ9rbX9+QLsm4nL2uS00WdCiQ2cpV9okBU
9btATpvvocG3n9alxg1QGO0p5Ow9vSFPC66RswvHVb6o/wh9Za8RqHw5Rnf/O0/GNU2zQaxXmbyd
L7HYpM4z3H2+nPWjxbTbRC4fX6Kmu0C6cQTpOnrfJ7n8upV9T/w1BbrzMlH5mwWyKmePzSAzrffY
QmzNAUtDAR9hR/UKtcZ21Pji8TzDHeyaK/uV59ST2p7iyUAKP4yWXbpdXmbcFa/wXt1uBKZPjuyh
8dFKYfrwwPhNv6pstYFl5Pm2+7j4wUZYztqryRcxoqWnoWv13FL4WgGQlaVqzDzSoHQT8JNYSsiD
zmUfR5fE/cYt1t6P6hhTgy65ssOvFzC9mk+oXdcXVEoYVLSaFIeIYCQ0K82HMgpXES/PRMMQgGND
zmadG3O9qF1/Q3+clxlHYB9u/SdInkAKl+XMKxrbMYG9AXV4ZWP/5JoHLwicNzTXgdM/QN45pGER
wNdMd+QQQrf7MJ5Xom2U/KPbyu1US1uCSYNToykiHPpzmogR/9j2863B1ad6u2ABp7EMKHgBicCD
lRV16V2LYw9NJ+4R2ZlOROlrp1opBygOsNzdQ7T9kpnhSqGcnPACM0/t+JchYglp6jU3b09nOcI6
oHbQmteb9HPVo5ilzwjtGqP5qYKY4xi/aP6uJLMT1gQF+EzgIYSMVymFhQBlt7fHZqsOwIROx1fR
2BDMzhFZnUxGE8aF3qs8IJpeAZjBzDbTmM3x4Z3mLg/D2nHP+PJKMNvjxeF1lHrCfyWQhRRYqk26
DiNHWT6Z4ygzjkpYN/jlMnDdX5zVKqwh4P3BX+JSRv1lPtWtexvXVztopsAtH+fb4/OExPRmQOsx
4voyMjHTQdNZZ9XUbDK8cBUYkB8SDd+eJvHgga24oN+zA8vB2uATSNrLPTTnt3uH46TxKpBNm6Np
mU1O8YBeOHphQj+FXQ865M51mlcNYhDwxr8m9ejgzLJDdslGP371R8D4BpnhskpqCIIiw8fUWhY3
ORUONrdiVN32gK+N2Tl59ivMdCxAF3BeaBwq/cdvb8dOXeMJKLDkgpyKYmj/pBZhC8+pl1+FvDlg
ry+C3gJrLkAw6NAVgljvI71+TVomiY2u/ZHion1RhXcHhtoDDihxbBRhKNUaVWEt2X/8Cp8nA1Ut
2sXNUz4gkmQpC/7c4NpWyWyWg2+nTklAJMRFik5MEgpQE52VQS3trNXLf9fjKzGXnklN2vECn09l
ccT9rLUbu7PaRz3gDzw6KHihIg0hmRK7nskYMXj/rlU2WYZYXpmo3uyuIM+amtECY2Te8U3CJoyq
vicSDsiNcwAMDxJFbIv+RyMXuXLYdr1NLZq5qSAd5t5FqPcdaQBgvSC+NQIwquzvf4wo2rVxgjKQ
DEp5SURHtyXzzNv1NR0j4gObwQyzkyK+Sh/WHX+Z6k3hTOdCQwdXyOPoKVPrxRIn1tKmUSb3MYp4
8G8oHAsZ50yVO+H+FnPyMCZ7L+vrzhPakCScJ1LRNgrzoYCQclq6Kl2Dtfxqf7cFoqvFzoRRBfhI
lLBd/uo8/O+zzPW88daSce5qVYocTn899QGO6lZoBNvHlFTzOQwzHsKcNqZcfX/jPhg2Ht+h/5LX
4TVhveRd1Etnb4c6YNV5d2rgZAx3knD2fcJrEA4SkOKMVVtaX4xt1JafR5GFz3vRdMOFzFHVTsXs
rwnseNWquTHsrS/FN4GItyxpYAWZyXyqe5gL3I3qhxYqE7zpFpwX0hmxv3+ovbg8ish0mGuhnjfh
oRocQi+SBwOMaCfwx+RBxI29suRI6I8lJBES3mB1CN6dMJzKgo31L3ChjZrt7uwI74Hf+MGVVdyT
qAGH/c9BOTNxrKdKhUnFE3egJGfMa0xgCsxjxA8lSvNKA21taZ9aSHf2aOhMLqOkSZrv8wAqXtAi
dWm5c0xoIkagNLXD/K6iFGxgJu5DHnyKEj9gCjNkLixW6pxS+m+2+iJ/yOW/QuGnXdQo1L+gBru0
nP1pSJ+tkAF3fXdvvTQ5smVNeCg9vxEwfvxJaGGW4tTGK/YkwbvA6ZSbAWxH6q8GeKj6/HzvTeO9
e2kgITLEIb40lWYAXCqr4G6auRvlyZ0xhJ8yg1CtYkmzvye6n0g6K+B6xGIHAIJ2YqyxmH8E7KOX
rMWhjNfEZC9jPHid2j1aEdYDPe0ZiUoo7dlqJv8secRjVGAWIe9zWXxRU5KdEPcfPeVLbVQE99xB
l3Q/kss7ADhvjd0Hff69zjBpiSbgfSztTmsxDR8UXxOXMLKKgGv078RGm5yOo6MnyU/+VgLingn2
vnIUsTM1R+KuzhFXAz5Rfg4s3mWi6iFkgBA7kLJpAuoJXW3cC4zcgiBr4BThDeX8p0yljfmOdYvn
c4B+aroirWLia2BcLVuSGh/aKgqreO8EgNZm5HHfgxo2wYTjEUU0b/7FWcgfkR8UqCuiu5eil7NT
ozelGvOUok+Dkyf698OUeEKdjmEjBjsxAQ0uXFPBh5wtgZ+ZRjus3QkYpMsj/4Zcs4SQcMpXkcZf
mez3fIfkGCT9Lq3OMfqTLQmJaCeQLSNODCBEmZbWiNVi3HJFTF/3sEYOnEF66SVnKntHjBWWPC95
IMyuJO/R8DcfGzD8LqeNTXBZGCiMvIZ/yH+BorgYMiv/6SHE6KPCyETq7KBxNEU/oHjmnwPCa3nJ
2WzvrQAbXRIXf15Qb+a9MVGHIEygXaJ3S6H9nYrRqZ8yrwr306+ysJllKeFQUhIU6I19dkxJSgLE
Aqhfj9rdYxG+/JbR2bh4G4FIptI+Vajkio9U+WT7qrcmRKPUzHwmie5QdtGlFbn+ENH9Aqx7cI35
WLb8IlMGFsOpNqFiophoSxrZTmdnaSxJOKvL9e+pHFbItHw7fs6qZIBwpoVdQ2O1IPn+KW8QbVMA
9eMKNFgC7HKQP03ti1GVVxDDaur2UB0xULHU39Mg4m9oufSA6dYPXKqOPC4yvfUy1SCzBxtYkXj3
E2nNof7p8dP67lEXYmYcVPKkdZDsfkddupaIFiRPKuNGvW7iOaSghqMWxyXXxwgcNIFzatxB4ejv
PX7z2mgcE0O3Kp4XCDIk0TYgq2p040l7BDKB//fsndfDK4pi29uFuLNy9GAAG4lgm7tIi8nRKLsK
jkmnyfRqeeaZxKkwgIg5vgj9Mt7yLueWvARQEuCacYGBCgRxqULcHmByoGfdmiR/CAySsyddet5i
tsFuchLKS/3e62lxo4RtXo+bD2YiiPMgbYrRtgr/EGuCfzLlPCkdSqJ45a1U6pLr2I2UrJ3WxeWG
acUr7qvhQZU3TR8KpWi9SS+XvmJv6Qwx184BB1X5WBwkKqQ0RzC/ysWaFv+53byfOv/ePqHnUjTX
O4TMazj0TxgaCUb2eDTJ8vwIzLZKWOLOPcEh4bQauNcnIdp+Php1Zh/yRJYTZWEZ1RzJssr7GfSd
Xk8NnlAJV4suaU1Vi7suYHPNevPSne2JhI1unt8Yfr/nbd+gjO6ZPy8sSBRaoECoGRt58s7ODRUr
i7y+Lgm9H2xgO+4KbpLe8WX7nUOa7tIogYqvHZEc9OW3wvPBGXA/iHcBLrRy1obdVzV3NvmdJgJS
fMRooVhWdAht2KUjIhcyAGFX9R8h7CJozZ0lcyFc2jhNUFaXsLwe+2KJFnkW+nenUywLFlxt4r+E
AVDqrGgaxRe4uVSh7D5E95FXTv9zuQ/sG7KxWXPothhOWwGb5AXrykWAU7V6Bwz6yGKY22TeTw+B
013i4xZk/t/JCrDxHXpMPcmlxGDzGofAlPzd0kp/eBg86vHmC3cPejuFVBNjHuxAmryZnd2WNn4S
hDEU7vA2EEWIQgzA+UMk8IB0R7UHR9qKRAYyGjqTmmW5mheqaUFmqwKixpelHEfI2iUqeSfFk00D
ExzvyzvFXMrVgRPNCEkPbWRmyvgdjVLllwbS0jriIvfarhD6aNyymPZt9EU/i8uSf61f1SUq21hm
P9hQ/ezxmjpx/viVS1I2steHyudIp7UYz5fDLnSpOtUGQqCfi1dv0TgK2e9EaP2oNGozCAFXtErC
BaxH77Ghg7vJ1D691aohXmigL8uUS/daJeNZiX2pUVDdtwo6rdDuVnQKTXG9CCrUd/RCzicH0Qz4
30BdiANn3gRwXsvEVt2oiTGMSTW/PN8nmTJLjoM7Q6AwYxu4LzMZpwQFsePKbilv6qSYFYESpx72
t1tlL7bKVP27+vn+16kJBG1PUGiM8Kwj/sWP6r3WTmANavShemqBxCvDlCl24ZOSkpcKqzJs+Jf5
IopqneDfGGyWhtkUwCNBBdyPDGf6NwFabuEF81mtOWmCkzSLYGPQEDbcKE2JNbIrLY2hCC4DA4mS
0uLszCxfH+hL5nFoOWMTywlNb7o4JLj21vYFhPp+GC0VZDav0pCv3KYlHeSoYVp26+SU6/CfKk3J
D/Cl8FlaonYcdLAQCzxperjf3FvRNEzFiSKLARNpAJ278+f7Xz2i/euS+Digd/H/YxKDlwlKnaBM
d1Pbm+gT/QrRyK8b1B1Qc6rTtt3K9rQ5zaJT2KKdW1wAx2/M6X40Cw+myVQb24IDoIjkAjG5g4rD
whOW43EjPa9LY+Op9MnAmRWr1T7Wa7mhwHk5eVJ7RJeWm13zIVjcJZVDPEIAjF7D9+OSpN3au6eK
5rgc0ahzynGdyD6VAloupkbnV4tno5OELpVQv87n99KStTKuXlmMol46TdFgmNvD6i00mFp18RvK
ZEwIFgDjt6zhQbkd8Ead6VtMCBRPLjy60TuenY4QVKmSBeUkaGf4n8yNzLd27E+PfIBmE9fA8Q/a
Uz+FFauBI6LZDzCsDD6hKeKu5yQ11kq24DbDjn4/PRpcXdeGjf5TjHsIlgwD5PXkAEKCKwtM15pH
nQ+6jEhVcNhvrlKiKwcBP0NRzkhAJtAtNtfEI7FLPFzI5fCyct+Mzx9lUW+6QIbhmoSVWvT1w3PE
cxt3YH9k9PYozm1XhGITHHnY79fbG46PgNWAkhXWMf4qyDlaaPilciCdnxnQt4j9/E58AbNqbr/v
L4Nhjs4XCRjnztruqfFw1gq+RCt6iZS03nuOcECJxwc/3t8wFKKxjPcRv23yhyOVF3c6H3sSx2aM
u2ea8DMKZLtIvSMRHvxA94pf6tUuBXASbFMZkCRMxBlw2rffFfden9H4dCx+UZkh0nA7BakH5U+O
ohZ9TjLzC0SjZv1EvAVMFwXHnOg+LnEzZe1naI++kmQsz4bycdi8R0kNBBHi8ubClgxKpIZOEtvG
GGyIH/Ck3m6t0QLBArYYTLoNoUEY6S22/KnDFEQDdp97hmC6wfYiStP+A996HPbA7q7ykmduVBB1
9Xb1csMhCBNiUP2QOFnzMM33VrlC+L0J3Wnv2ioy6RrWP+wJfvdjMqULZJrSb74EwYq5Um2fMw0k
qFzOax8HAApKUd4YqwfrLNyTIF8n9b396V8Ayiz15YW11u/JG8A0zyj6lAJkIHvRro7JQWIoveXV
Oa1jhwWmI2MB4v2yDlg1zO1UHFVQn6F7yFnq3WMZKAPvncSYZKs3GwfdMLaOl40bpHf1xBokVm9J
gYfjTN5F0zTISzu3O91O2Y/tKBO2JyvnMlT5fTs4ZI3sm5oyCayC9W8ShJeSAB65jr7Y1HyHPnsg
jqg4sOrAuSxgyq8KalTbZG4D+6tr3NRYgSgYuMjXs2y99XaZzKNeNbHuCbRwN7deTpKaeGILk8oP
DGp5Z0mg2QEy0eUj+kTD8QTzVilbvTyH3Jqzl+fvLuOHT4RuJ7oK5l23FX+iNgBCjRv8JZeL2FHT
DmWeFdxealbRY5iv2JQWmcvYgP0wOTrebfwe7mbFYLIzeCmgfVapg2BSM2dwEAFosXMhg1FTj2kY
R7CpX9TfnupltII1b2kBf03UPEMQPyqAROWPv6DwtlLEtt1p0Il/FRZ37X0AYNveEXMq3iQ9yXdb
jMqZNf0286PwYstayPfpfkloinTkPF0GArdu/daZSwAPBo9Z9+sVz2BsxPeWrrEb7Sl5JXOm3Rdm
2Tr3SQsZOaaDfhDU7PZWuRCdluVZwm9+C9n5kigYFKbDIfJ2NBY4lQQBUbLKOiWalkzQj6LqnWun
bIFT+lTPBZs04iHroMHfx5M5eHAt3xShtQ8PBwqxOoHW7zRzzgLTtZthOZwRoIzl18Eq/l2rHh9B
byzxSKdZO1zhseNU61yf6mHaS7FICpEl7IY7tmvYoXWDqaPut7+LrPvIP7D30fqvw+6xsSNZonZp
PZKKfxSyeVYbWSBPlvAR5BT0CZw+PBbgbto1U0JTnOWFQ24fUGgee0NQrpuG8rq/6UI1sbialu91
Obox8tZYKvbKIdIDFlAziQpe5qaLkyHLDKjnei7NSq6gGDMLRqMXv8gGFl2uVwmL51gu7p44v1wT
B8mQurXnIrRhnUh2H4o1FQCUKhKaWrZ4kNH9Vx+T5MAYozUMDvP4JZ9lxeCyAjVPqE0M2LCwvIqO
wNVrk2g+S1fqaAp7F8PcZttr28qvAXvzgTrRkSg4LnwC2yJxHO4Gun07CRX0aDeSbp8uzwbd3QlV
L9ejrTM6QP1IoRFig7GuvnoVIwgZPKrgXnby9lINRwTuHVBHNJJyUngmEWoNDvB3sciibBmphEd0
FIBbG74n6FTsRYTVY644ZnUPbxsRPYO/1z1ZF3sT3TFn3//xZKzzxZX5LT0iZAHv4Q1QZNki477r
z4NXAo/8DwJVuotRprdSAoqAFGThEwKXqMK5O2zK3OPBOLZjQ4en2PRhSQs4t2Bue7eYV79BWyuk
1yy9kVXrWC1wXwdr/4oWqvwgqwb2UMbwPzH3QfRK2iE6w0nKHmPkXxNUYg5kKjCB29WbpMeB2emd
qtISQLMtH0T7eCUFajyWR+xk2AFry0c69TVcEgDM/L8sb8tM0nVM3vzzLRyNxWNj/r5+eRb1y72u
oQN2yFXO07yTPqANjUO/1WCx1hmsb28Sut+5k94+3r2e783icFa4QYKmSnK7NWbYhfvWkkKO1Bwq
kx3TKsIYtyg36da2nfeZalQAbgHoxmx3GH0s7nJOWnn6alBxbEFU7Uq3iWq89qPa052HZjz8r9jC
iqiM5nofhBcTE+uPXVZz767ypaahfojt26RYF2sYExhZxTekehSPkiBS+DXZGOo2ImIM07bU0Exz
L0DfbnVWEE0zYUz3dcSr1UUuccbpg/Ppvlvsf1IEDxhuGl6YylZZZvUjiyFgFmzkUnuwr1GeAXuR
0HEY2/Tm/nXlIN0prgo/tyvspmLBtNx/0Vrux6zwwlYP+CF4U3o7qfYupmf6N/QgdkHPl1q/jWmR
I3NUZbSIzkh7nxyhcYohASAb3jk+VwxUKTQ6ZKqra5MtfmP121b9xsg9bHRAu+ayubcKmyDSgNKE
w6ssXdPOxLSpKNXgwKcL7DROvnAQzKiltjeFYD6L54p1kFCckt/sJhUDjLIaPneLDB2sit6iG9V7
VHYzBKt99z+1h62rP9Cj4OzNBkymHihCRwz24sOVrw9SoIkm611sMb/Xmpaugm2wfvvt/0OhAv66
IpldxPVaoruGlKqAaS2th4BInOQd10wZDQ9BRexl1VvFVGZ9dSOpD2vfDFy8XLDB6g7JtimtLKV6
egA6u+TGb+ZDNrfojZHfaaClts5/gO3CntP3zOYF82cOsYL7OPwNyxsstkkAhzIn6JSLwemFMpbv
1pBLM34SoKc/YKQYf5CYk/RmOrJ0ry3ikxfbRrVk9NtcXMQu0NOun5rBzmpcBtI1KFUTdR6G5Sb1
wkugQ2z1vMMfEg2oWipYXuzEo4tnh6B5Th13SISIg/mqM6f2zUGV7Ep5z3ew6XS98wBqy8cmQFO+
x9aq+dhMdoOlKhRu/Bd00vKqLbXqsgtA8HKorQElnNb0/7TN3ujCBwpnW3cAGbff4gNwrbqbFSME
yc5AcauVyfB91WZUUoA61/mx8uxh1H4cBJYyV8KtJvK1umHva7kQ702uSEUAySoV9b7ZBluJII4b
Xm7QpEq8SAexxaAJJNLujBXAebhMfqmEHz3GfdoF/HR1VCgXbbkXK86KETJiB7XXCnjYu3XSim03
yveQ5KrbzsUkh71wGzOkvd/w3l7t48ulr0S8oFWTyrX5KJoLgqr35sxH5xHYuM2WfO6Ued0tmfNR
0lLqaxNe4+pmv1CCDN96V5G4cGIq/mEfszckPpPqIP4Ewj8veKLASCbLZrm4gRKpRrCj/kNFMvEP
pcxqIl41Z65IH8wYKsrJi+tiKRbc6Zh1MQLTSgNUcH3lk+qx5zymyyo89Xo36eSLb3pveAr2tSq0
fXdZvmnzTHn+CyMtyZI58s0fIeQKQvaZ+LOX0cOYfbiLURKLchApmUwxqdTG3l+1uhtMMp2pcC0q
z8yLpWB+5YDnJ9DDTZWIM5V3oJfE/UNG3h1d/BmZfL95HbkrDXlIzxR3mhjV4TJVN6hKsX0gyBfG
AzCv1BjWXgstOBRswN7F10VETou0tMqf4O7CWkRhqyX6AoJQ/IbAVKGm41SHsjbvrQv/P6aPpniG
WTtBTHo66b0g26sU//xQztGrf9+egAWNNQcTlOlQ/qTpretmIMitI6WGQAjO8YYScQa4/B1wuL+v
exF61cBVdvWjgcNvta1aR1qIqhQ4XxhUeTdL3MJvpf9b5V1DPC20nHvR+sT8mARedDZ97u4PxszG
M5FhLSOEOiOqj60OIqG2aMWhOw5S6aEZraVpeGwZ/QpGiBhQMAC9iw5wGgFgawbBpPT+Txd5Ox9C
zU+0ZAzW/N3NYzZQcATAQhcQ8mWAu6np7QuCix7RPIC1M0eJZmL/Qruiz3pX+YkaaEgy24JFYSS9
yrD5ZOXiEs7Xaa8Sjvz4Gf5MBJIttw5Chuu87ne3Vx81kw66LtXqJo3d14U6xkqjs5KTuqThGBBz
vBdxhWRPWBadSkWA/BhrzbPYCqWWQa0Unal3yy3UdgyYi6NmU+9WGOlc0cOqC+Ckl3NjzLvUKIXc
T4cLEWJpGUJ2B4o5ti5Odzz+vPrD2zce7vJGMoMzv+EtDF0eX0X/eXk7iyoYvGLmLfOfURqH+XgT
FruHSTZLb1C9nIvSVIRTqcVKsml0nFdBzQjUicZtNkyh5RpJc6xbHUitUWYDdG+6j3/2i6ulrzyP
2/7jj5Ibqwyu6Oi0RpLaEDPTIFg0JbA1z2tL4TH5Z1n7Esg895B1z+rSU+9eflMbV8gpwsz2K1ap
RAKZYUkQE6AFdZSnIfdafko9l8Wv9rcwBuVCV4tu7kMUxqXYqAV46bSwnnOuzZKc8lZGTc46w6sX
9kF+d3E/wVpeAEEThkYcxI8f+gC1ukFhsNVR8ZjxKoVUgvgqjnh8FNBSO0tMTuo5sYgGfZado5AP
hUFuRylrP+qsBN5aptnUMImuvwGxZam8yDJ1G6dLwG8k8C8tozvRxm8c9L+WEl8/PlVGjH2LSTtS
4hm72UZfBB6Pf2jqv2uJwHy9YtmABtrKQd7fS1A0yajeGhJQ3jMXTYIgXoO4cw3rkJtKCFzdOEg0
KMXIhAoT2GHAdZ8XsUMeAJPVL5K14RBQ+W7PX6QWmVn6QtonGFrnDhOkNZHhybXQvXCcD6G5ojDN
l0bHh2FSl4Nk1JGahKIhAMhkwysux2enjvXi39qAKhY2q/lAAtLD5vy9pyN/XdUtxq9SO6kqahDb
RhnWj4/QqFZb1Nx13I/FrqUwRQgfaJEkNAcPiyB1TVVR0rCUKswHwcJsyQn11/B0GKLWPecjKfTZ
QVxu8YSpcG6xDIFdhK6hRQDcZ/pNuI8J0z8+u/xDVKO4orrCRQo9WwNhscU7cxlV5txeKQS8l2HY
E/wjZaYTSNqIXx6JeWeeRN5AjLRs5DMWige1y1nqek4JYmdNSjqvcOt3SinltZsBn8Ypq53EuHY/
1jJJl8Mu3xo3ugLZTFYZlxwoo07BP0o5f5O4c3/Zw0S4fyuUF4YlvpqC56hmMBSlinfVkdIQqQ+x
BkQHrmJU2EfKFt8jfT6M3Dt2aXKjbvGsoQl7xO4Tz2dOV9XTiRpBtn0lVna645Z/YHDctzuHgEEh
vAm38IhDTKvLQz95o32rw26av4wryRBWtto1aefIYHR+iB+qnXPnXuomERfyw7EETv6i+j831xBm
PZMbZwT9J5Z06SBPxl4nvevS6fkEsNZjR5KAHSBAFCa0kuus82TjhhqvayJBMCp2XgNgEsQIbVWo
bXVHcd5tx3c0MlX4/xVkLf+Af5YYAnSlVXnBuadFIIwG4QNwERZ9UxW6JFfbganniYNTb1AMW7BL
JbdXoEk/dFqslKD3cDlMqnfP8yuK547R4DNNI8Bd4gz2UmxrDKUgC+10Oyh52X5LPPPfcEVfDzoz
5suR5EvWgf4VhnOqjZ+LTJ7/JIMXWz/CG+hjEnspoui8cP5tiOJs8HXbjSNFKr2XjkAbesifCY50
0+zeWqo2rf7Ec8QneB3u7Yymoddt0Vd/BunVLxi9KqZ2sGN9QfdVjA3x7OaXhKwPzWGvUsfwNjPL
gbOMI0CS7Xj5vaYWC7ypusv47YF916LxoDUeDVYHkQynhaW5Qbk2/9nden1HsZAvUB5YJK0wMGf3
8JtqCha90ttZvDLcKVqx5l0zCgb9HZhhcnnKbZj2HBMWyr76AkVH8C7aDN9sETHBNmb8ChiR+pUN
fWC4KVVD4h+Tr/htOW5jz4I/SQDqwS+EA4CH7SteOQX5iwZilAa5MJhQv8ssDf6ZwiCW+BMlJ6fo
Sk/rgwcVvkn0W29ByCxBGf9NAdCi7T1JFZCfrnPS+0Vw1vEhBT5P9o9OCeYMnwqauQM4ogwRxMyU
fbxS84uNohlh6mFTIBRdCr6gInaKkEsXSiv6WNd0P3Y6/KMlIgl/cXq20VjisrwH448xXpvmvkvb
2DJWE8gR8BOEWp5+HtDQ13Hw8oUYmPWInojaIDNum554NGmkZ66Rk9pKxyKg76+RvzAUyqg6hQM+
FNp/Cv9P5YyRKE4xT1D+bwdDOBn9RklWOrPKoq+LpLODApGEPFiQZEdUt0xws/W+kR2S0yk9j2Qb
OZI/kwEKQg0GwLeCq4alglwzpNmOYlknVLM28a4rSSqru7jlj0F9R0MjqKXnk/hojXuTueo0Xy22
zU/zRMte/gUfxIxxXoPJefq9Mpg2dx2eD/HnswgR7jSgn5RxzLXGbZ6Jc4vBtBJmW+PN6ceCGIC+
MtN5/vXvhMihOSOi7xYwBLg30eeEvNPw6fSq/XtnklljV46ON27WSrcRfzQBcxpRX7xvO//v03Bl
MK4NrujEZQXVR68skkKmMsCnCBhH6WqZ7EvdgLBeddewoQnj+w/w9Ng6rBhuZF2nzlaDVpqlniFL
rcCF9mbg5fl5NJTF8kBOjP69zVemCjXHqCoki+JXGaaVuvutBd4kdG5dk2RXtPWKvnsMHyx62Frw
bHUYj0u2jg8+afP6sgWXhv/diI52QBGy+i44E5VgwgnCt6S8hVsbun6d/pqQkVzvMHfiRWOFEAwE
BovGKPPAIWvUloSWqRS+6WHYvroBzeAi0anWeuhFKy1XCv8URYVaoKUploJA2u7IaLTrbURoSERB
A/xr+rVviCxho66PGKT/u1RDYkzQtGPo+r3WK0n7kiBE/GXJdFGn0sqxh/OhE7c8pEIqYM0QdErY
IiMl+SkPZ2Mkm5gfC4an5pFfxjWoWiRYPBAiYW0mgtvxB/vs7aUCQt5bVXkAcKubtOxPSLd6CuRN
3sIoJ/VECG1ODoNm0MyxyoHoRaGpTtpTY8RylrLzwGLNAr2YUTasW0n611CV76tI6RPUvq3ose06
p+uptv2F1TY2+S1qNURB2gnse9dmgCPD5mYgrsE/jIE75H2oiBk7rz/U5tft0aciHXmpi6uxQqq3
MWuu5JoZLP/CI8XrW1hy1h/CfPhqR/CL5ApqhhDQIxf4wRQed9AGQNvzvyzbI48o2F/yAbnzr9mf
ZncmgYfKvaUy3FLpCu54IhjpNuXVUoQ2g02slY9RHFKUKfuv8xZMoFAxD+lr49dze0rNS29dmmuJ
P2ZIgnt9RVyfbsPLWIJT9WKxJWf6eGVesg27NzSiK8HVQggv8TYRbmWUWWEicfP1lzwqmcgQ/pLd
4oJ5eBa+tbpjYCG57kzo/54y/LhqZAOjxPyNbuHow4sqHq1upOPzmd7yJPVLKX7TOKIlRtztWj5f
KQyiWuY4FhjzY4wlZyrXo5OBTx3e2jKHR+ez62T7DdqCnn67Y/C55XKxh532fdKEi5W6IfL957wD
TStMq4BHPRQXmNuBhfFiielPStirXU3pLLivm7+xJTW5bdwzN0nNs4/1MkxlR4oyTj3MY0ky1FC8
JYn+B5ZoVEH2zZZyVf2Tfu/lLShdxGKSk4EFM/YXwfTOBaAXZbsvtmtNjUdwKuE4BPL722j8zGEZ
5Xy8wg9ckoEklJcYMhbKpF5VpXGpCo2avhj2JWv7ZMsYUR4JM81O7rGEsDtDsC47qM9aK/tVdJCT
ovGlq4lP1Xk3S9x/bEp/I+ys7x8VeHBaqX8ash0m7yyJHGiar/s9gha1qyE3hCGGpRUoj1f4iSeX
f+J01xxilIUk+EE8A48rP9nnGL2E2mOAZZpKiJFPTncDjzeh094Qt/PqMAcpTp8md79VjMVFpyRF
M1GW+bh9dxFyTtHeeonKcgjbwrSxsUw5iPzLJH2gEqdPGGBeDNHhOU0hIfUFF2p3yAyhUjVmy0Oc
T5G6R044+kh8iJuPOQJaul1Chvy+G3QExyQnepH6ZrwSgDq3fEUhxoGK5Are0YAb4J+NRcpJMZtb
/RhY1tXq/qmMA6vzJNiReNtw/OYHyjkGUxNujGHTSlSGxAn5nL/vyB47goAMCNi+UhKGAlp2GfWK
PHqBCsWoknxiINvmWdtwgRWdWlHo5ARdMq39nsn6ajYcpuPbjzrFIo322JB+0TVHKfxW2j6j6WaT
IQ9Hz5lFgmfxVOiAaf69qXzMaHQNcPiRs/qiuP35lfVWA6N+SfI0sgDikD9VSNMOgJ8uWYzkPF3X
xuzi8S+cH2Wpo0BMuAuEtV7jS3WIMSPtUUVfesJxoLBnXjuAijFMYfMpkzuhyidLmh20uD1kXXIZ
RkGp6C3WVO2ljoy2AwYiB3URvqeBuMcvK/ieOwSHO3w57caDhMNl/WGL9s60f+UGuaZFQ/GsCM57
+uPQIjsrgUhed4tTv0S3Mzd0Hs8klEilEO9umsVRSD8WmZUBu/bucxwsSN3Z2KcCRtd7kVoWv3H7
XFrVOfsFQfX/j5JqKYBkNqX9afYjT3M/BSaGoOW3lRkN1y0RmGvwAOBLFgqknciT6hC3J97NxyNw
i/BhyzQPrphFIFuEiTJs9h3HgeYp0Z9afahkMti4nxOHgkq0K2JRETRniRlV2YRtVqUcp2mXMqB7
Lu3KvtTmD2gZtGmlla7fsGw00/dgBh3IqA8ZR99fHFz6hbHR1Ng27BoqBlDwQNflBEl4P8r/+763
LS9sxQYpEpgaW5ZwBJlFe9g6WNjoQkx6jzjZ1Jv+kHGZgxyONgA18O96vrScit5sa39J79lC437S
LSp+aajXZwQHMC8xbZF4/cLT4XxxJ5VavDKRyAZysazh49Yj1FYIQ9a+VEQZi2POjs3AYltNKR8A
SOoyGpr7G6NzWfZZ8RZt0fmzzr9M8NG/oQbxWF2YouxkOweLx0JCTZ4c2ZVuQfeR4hLrB4xjvHX6
spyrMUwA+y8goieZK+5cuhI1GDpmHubQGL2kOGjs2X4X/XOZ6NDGQxp0r8SfnONW1DF7WYSj9ZEb
95rfPiVJGnGdoOP9eztcsmTJJzEbDryCUSf+tu5tjyDJppyitgCdDEIYMTh7nlNV2COpoliV7TQw
GlGfUFLvPlssl9SuDEt1v6597TkMUMDXI65JrkfpM8u2CIGklQ9KEWC32tREEH5K/uokg+WCVXIV
eOzPp3ebCE/gOrcNR8hZJNL0sv8rxFahm5Oeiiu8vBKYwoC9iaQI50iJ0i2jAk1CRtbDUgyqx+xd
Kj6UzTc2XPrKBBNfJfn7cQt+ECpNbSGQUq2bcODw9djZxNxlcu6SKdghgpoSwtQYWjjvz2et51B4
UHdCi1Tw3BJNV+/3S7pyHDdv6baRFxtG0qR3LIqhizfCG7IXirq0elkDwyOzNstHZxJnisTsTCGq
Q62FGkNYiRbdegfEROmxLsbmrI5+uTygDaFhYB2ArDQFZib/rC4UlrtyEwcArp0D2iqcNqvC/rBb
mrH/VIZT4oOljnOwt0VCE88P3srA5S5pPd6kp6d7N1m/ydDXdrDN51BYon9DfXYIyiqCRfWBny04
9c1Wy9vtjteKVIwVD6F0dmGUbg9KiwX6WCDDxhzl0xROOX+SORTMd77DGBaYYvKhcCKzZ1qtvVUx
heJSXxRlC2zbnkt+19JZnBlpNHaMasOQ+NtglHm9Fo2fzPUsKDTkHFhCsFoXETqrbqeKh/D5zZJp
zxieqmLIRXH1yFParcsVOex7+roCwUe7vxUxLL9oiJLp9u8NA+yodhRu23xZEsyxc9l5+o2GAqjS
S927buI7cY2Al8sBusDhVQWSGKScOd9WN4bp/EeRijPrtFB6ziQnh5wS3kjtOnOeBCDace2uWmOt
0Wex00MoRgwInzxrQ923cB2jaIrLb/WbT7XheO8B2iBghM3XNhqBuZgNR0Gwnh889dbukXkXyKLa
CXZjLcfuPD5ZS01aLLMNzx05XgCN7I3EN2MsOUsDHvjlW9Q2IB2rEbSUGi3vB7XuV3WM1GqyAnRB
EudiSXwTlMGy75og4Mgx0X/tDU3LQw1KthasYGyEYLk73SmrEkmn7kG8L+dhld6yBf0MAuUp3+0d
F5VHTjE0rUEuAUV7OzXTNyM85d2eqnVryfYzHb7PJI9LdZtMa1/Fz0M+SfIG6nn2CFE9mCJxQAre
8IBiInuPKYA1Ub152qPgNeY3Uj7Af+5+bOPhyXLDjEarhF5FXJWFUviO6uUoPmxMir2k6z9oICZC
zXsChm7NqvhA9z0p11IZ8SIPhXNpykYkN27X6i9LpWla3UNe1LOQtd+TmRPax+BR1PaAawpdqO48
wwGTpvmmLQihpncbL37XUEAUipwRYR2E0CD2uMn3Ji8XdM7guwkW9mQmimmf6soDdfpv0uRgfRFv
6i2maGEnkvNFwDdcVFje7KEHLgACfzzuK1RIBANknQ527QERURSKT4McfJ9TxIM8f7kvLwHxjU2g
RPCx4/PSAUEFOcYHPu1c1NWe8ZyRwXBqZC0C2Bldkx55coWZIkppNph2Wr40J+totAEFjmEU3GJd
7q0HuttHWub+8wY5umN5e5y0/4DDc566Lk2PZaMTTJNHLF39xGb+hPcrvrByCwk4nr5uLMmw8KuM
wTLXVxkFicLQQt7sGhCxtSzQNZhHemxaJzDO8bQ4svOBgDhaWfinFvsLb1Z2G94w5Y/pR2lhlFzO
UKn4oKgQYRutstK49FThgm6DQhUORu6feAHemxccYZci3RzQCPdLo7GACOd11B4qBMYyORUccKp1
D65dxDLQJB04dixUW5I6QbEbN7ggej1+eqcbs4/wraQ0jwQIBl/OcQ+/qQsBYtAN04aoi1iSq5R1
p7bRkbq46mdLNJCUoW/nIZSc8DQRN1AfMvL8OZbA3jH4xOgSr7SKceNnOloNIoWc9rTXJgZlc2F/
tx1grZ1zt/UseQzfLzDgk9DwtT4memqLAEzIvniSowt5vSmqkNvqnfw4phITx6j0JiGRvhEsKdDN
PPg3f78YWVh85p6aePG5Ro+f53/tm1Q32vpBGa9c2fDxogyerszWFrXj1+wMmKDN+Bl3sE8xywQi
KZRnBp1phVks+Z07HYfrSVFsKCoU0EsaPq9K6G+l7cmHsgqOUqPkpYILjWW5F0ffDZ5PIWAdx3uJ
6+DlUFC6+AW+1JV+i7DQhDp89f/JobYvbKAi5Bm+xCJdCnYOIl+P2mgXz9MeF7dzgXSSz3m/FPVc
OeBC/wFi68J5be1VeppsuajLxmVyOrY3zur2969lJrDIYuOcSkd6iNXw1NpG3p5Nong27i2uRbDu
pUwcVt89lNzuT51mXgiZITLsi889Icro03LXQdH+HnO35uAv9jc26j0VxumvEJA4rj8Tf9kI5Hfx
vwcfFwXkRUHT1xltuicT0uZQ5sGJwMf8cTXp33jxA8aAykZ/UGFxkLdUgOhm2iJ6XZMS+SEoQi28
a2LX+DymGraTUcLfzScuk2MqNaFyClcJgwB859HxjFNBAVXfCEHOJBIE80ss0sxDp0J3OU94HeSk
nU18gaOx7fqz0sc0VZqhVsW6CYj9rS13fL2cGEerFLBmC1pQ3AuA5eTskWX18N+kxE2UiyejDwYZ
YiFr8hMseEJhZmx91Qh0YxcYWxe3NKwBysx1Syq+NhvQFJ2G47N69EPRUkVNmYYGLaOUXGHyCpjD
6yp14vEYNzxGTKBG5mSGHvzYmCGpC//8bJ07ZizkqFbWytlTsmuVEMnAt5/5ihUGgsa05vUxW3Wk
vE9a9kYjKyutuQCXMFlpfk8OFVjTi9kboYyo8Smblm0DUk9lLCfU5PZO47skg20J9QBk8FJFCrJF
Q1OFi7nGUCrFsyd1lx/dUP3nv9ATytnG3KqNS4qyWEQKbDyaukVyfA2aCdOhmdSzV72zWAuiySWN
w3UOSEQCDx8JvS13xZe9gIUsaGGQwwNhwUA4OLaNpk+6ono4zZro1cZlXk4EACoQAyFGx0G+HtmM
41p/cVF+s0EJwWuKLQCW/YzgSBJ8jmaKwhd4o78nKlT78etygnMfK4+/qz2hhKNv/PeEAnvci2X/
AUhZbC9KgBHJyNETgNQORuMP+7L9s8W0h8HXyZQjAHQiFiIn89YJgT9BChgkvCGseNdVHYop0xHB
QxU2ARfyIp+ACBTks6TpVNtbESNShOaPuaywM7sSftQZrtVZKn5F57axO9p1Nk+3mSc2vClvh06u
Y2nLhRaMarYcxESx6QwEL2FiEE9WrUAkTl3qw7y+0Wd5OkHZuuS1WjQlx49/abTIUlh/euoZLncI
irHRB4MbwW7I+1aQhCrptuHnO0phv2fH/o1tbLxFqfjmV8XQO83BR7Wos0Bs09KqrIhf6ndegMCQ
2DdCmWkG1h7xyILnMpCyE6tTmMbtGGOrbPQtqsyX8c3jNMK4M32ZNenxLKxyHwih5lBHpqwKitL4
1/FE2dXE/kre21VPERCxkHLietxOE8INlR3fwNfnn2fr+gyRSVMoW0tT+ZrEznDkzo4dSWLfCUft
N8Y8VpmrDqfwTWwTnVmI4sG+b5N/lRySAH+F49qEqHHUErh15Hq53bItQa5IhZC8pNsjnNPLcAtZ
onhJqhX7qlIZes6nqOiepKank5JesXkWWIAiEP6xRNCQrJH6arzRm0he3/PvGi8hkbtK6txLgGhu
uIlCcnVxLCFuQy07pLg7wMKsHuhvi3FB7B5T/jFDQa/N1pG/CtiIDUQWkkSvHX3ePYBAtuT4oAYO
O1QCZCbjl4Ia1Yl0nzqPQM5DTzfKTyQGzKozkCDN7cgMeBgQk23e3hi6SunYjVvbjY+w81XMT2Ry
Ysx6B6zRGdOK6gqmrgnentsVmw30hv2sCoyxML7Qdr9tbOTGONLlQB3FyKKd+2dMl2BKfOcrCui2
ORfnPxjA1kOuTg22YZ5OeeMpjlGsClnx3HpWOVgeqoXN5JqFyix+wkg8BrLBtB2A76MBV98R/SGG
w9EJ7Gd8rzVjMLvyLpPdgKHYWCuElEGRXD4ukyVJQhTq4lsG5MoejumKd5wx+Sdzd/qx0VCXC+9G
CWj4A+05XwK9NIJN1ZZht9XR3ZdXfbBwdEyZMw+5So+j31rflTc7n+NO56v7c/RwAHY/1+iWCc7k
rc2y8Z6vgdK876TkXnjDGPyvjKQ866e33S2Hr8Kc+t1PArRpyCgutmDeaYPRcaxwhIu2qlG0nqvw
WizNIKBbLLqoqXv7BbQGM+cK0EAZDGPuPLXL7/sCJOfGF82a5KCuEgUBNmQOhoSFgd85kaOQ8gI0
CSF72bmDtMqWla/rJbiBYYSVPSknvCf3mA5t/XpemzdoGNszIDhPOZ7Z5jTTV4D8QqMKqVnz37QQ
xjdunihbYzV2fSzjd7woZqTQXop6qJgI5MFNZ9JiQr0t1oQNFnOIPqABCj6qr2dZRGWHKnZc3vuF
ENAJcxB6sJijpoalPNEiwLF30cDcG9sHFZvgTlbwWwmCcklC38bfuBM9Hcl7Z2AIE1yhwtIj/riw
HRhCt+jA0lNEzBCz/xymTJMgy6ZGHUl7DuYpLDNOg2jrrAdfXO9WIMIMPNiA1v47fHs7xAWxDPYz
YU03azh30lvo13fW+5aaIGguhWTXzYmbSFCKOJuIXYBqbJ6XhDTtf0uxg3HFllLpOeFTb2aJ8yMW
8iAS/7IPxCbrzuNRCDYyd1tQdF7l0DDEwxExFFOpbXpLzSh+acG0VvLMLHIU5ny+1kdveI4ZwihA
iVvH25gzlnANsEI3swOWwlv9Gkv0jnRBFrl7/HINpWXQk3AJ6kKRKbYT9r2ND7C69guLS0IIVV7l
9JFQZ0wKo6Z7E+L1Wle7KX0U8JWvKArUMGQzSsswa1PuhLdOA2xkISXRPjuu5db53QBfaUE8QP+w
vb1jxiQC69cwgzwJ+Cu0+6J4WS18+q3Qii9+R1mNi/5lU4USq9l65eAGIYLIrOBArSYM6KJogqLA
MW86VvYBqRgyxBMZi+0QLWh3LA/xuarvlRshaUF5c/3okRjDxqbjaWa2bv4b8ZK+9Nd3S/v51QTK
T57s61NkLpKxEj/loJOl6dfU/GZulE99pKjl42eoJRvm9Buv511LrQGT74CPJb68HYoZEfbzgzpm
vPkMB7dnO9CD959+VpoJtXF+0RYU+g0bG8FTeCDGE395iICvghmUKHot+VK0Na+v9uUiRFlbL094
5K8UjvSi1fGnNZf3ZmLWS57+WvLfdUK0Ra6FrUDAS4PEdokG94E9MfqdRbQbaXUkjQvUDqQlUQmq
faxy9UzLijfIflwlbSNuqxpXAEdVB4YRqY62aYIEc5GWv7N8jBlK1aGTeIfacil/wzUEmJ9JDQrY
jm4kZNRniAhNu70ff7WhrofzewSzwILmeA+ldsNUB0ONNgCK17UU3ZleKHNIIyRWXgNqDEI9YJHo
wXIRrDWSLSQL/Q1Mte97VOAaS1IemYvoA0u3vUzgtyB/u30cos+PIW4thpD5BVQRptmp8n21LS3C
hPhZkqxx+qchKc/w4yLztGHwnnmttP8YxIfcmvQJFH091jycjRAWPAYIUgI4kRp8zFIBdHRuBbmF
Jl4tMzgK+ETBjx1fXl8pOyOEAKSLbzfWrDyw8wbSo6UdbgdoKQhe/4n3rMM7sOoQszS2XjX26FVM
MiUt8rst+w1BfpnmClsYWP1QoNyaJqyHQLqt0s3dccf+kDrXmC2ZqBRUKy3TE7K8S3UfOzAoPH9I
xn/3se8+PXnUR0WyBcggOZwcFzwVwiE2ZBgrLZaS7QpmLQ2+7UqUhOLN2KZvLn3pkYq21odYtaTX
WYlB2rWfhyLm1usEKs3HA+MJshKMj3SFjQHzdZvk6uqAb7QypuD2AFoooy8UPJSo+GU6N3gz5o8M
pa9SH0vnh3lFL1quX88REBD6SkRWT7sbWhqn890XOZxTA/0wCUeDk7cPqPxrFR+wpRQ1Pdd7H5ZP
LhqMEIg3+9obC+02MrhmSDRjMhJ7uWWkmaUoQn3CpIZ4HTEstIQZyHUfxXnBxKKgom05/W2fseVr
Mbq4OZdfS6iNRKrteIrcEW77E3eC4GdxUZWe7dgIFz0mCYj7GoMY3L3XTWBqD4SIncgpHuxv12Yt
Ghpwz6+4N6KMwOYvlC2j4IE4HMAPWsV8+Gmq4pc9ASAoxSM5QuN2EHXZKot3jOwWiZzn7eLewteG
FME45ash73iU19jNdT1yXc5Oe8ZoovH6jhbqDrhsvir/UNQr0xqesuP3sFwVINgzYl5yhDVCdtfM
ajHPo+BlPypaUkOYMx31fCBdqocjIIPEBBoVQjKUpLYlUwbJOxYAotxe7OXVkmC6b5sk1p1DP/Jy
Q6N/Qfv/rdjNKTcLHK0qxo7pH9chebPTGnVXMP0RNL+Nv94y4GygXGBLhEnoA4v7GsWgiWuJWBZA
Jvc0u+yeiK9gfWs+dwOX2jlbPJxdIWWGhR0hulbWYI4/+deyM33/dSVsIpdTeEv7+OzUgmD2EBZX
eakF6kDqPOeODBEE8oIYHZ9u1m2DCY4v3vLVBiySvv4GGQf67zjDcbn8mfnTKnFdPoLhbbSlJ36S
kbiGzJhrCxMhbcixQQOQP3jOhr+VuWLn7yy5xT6qypredBj7RktkIhlp47yD0z5FiO4PPFOqNQJy
+x+fLnzr2XBAZQ2N/OXD97kgPEryvgni3EGR0Znx3OBJ/jpBWy1SdFs24t+I2784XJyZDaEjN0zq
6U2sMHLDQBFGfaArCQ2zDaPpbUhDC7NHo6qqhK3eGX8RuwagO85UmJY1UJCSb4VnBJrvFPucEAXq
GbO/xpJpMFtvhlOpvGYqCcWxJHfoHRsNLLtG/dKAPQSnnfXvB4MDs/38xt0k9KfVKcYho6TxdZ7n
WHl+SktRBkRISQ1zeMFzswV0FJQQ7D+7jaQAHBD7Rg55n8aqYCKSHEmTyrlwgEMZfjq5QAETzmzl
plGgaWOWtXtKlOXCB3BSXOGTCHPR3nt1NIx45s6J6MFkAViRicAgqiydcJBtCAzn6IilZf/Adsxk
8GMzzkMHiBv9uoSKLWRQY1918XxPYH5oWc+rPMB7Wy+7hxuIi3Mg6q8xG0hmoJip1BZXr8Q7QP4d
mtOZg6QhnI33NqxzyJMSEg7bPNFzEY6whFZA2QppacMAO9ag/3yRT/0VaYit38D80rBwwrjYTuRv
XoJyOx7J4K+a3AsGvk5Q5hkVoynMF7Q/ULCXGrehSJmtjhbvdzNY83p/97POeQcbHLvoYiQaC0Hi
Q+bVgSK+4rQZQ5CDYtRMXemcJfisUZfeCGH2XLbyWB1dKvwLaWXWK1lD0h92XHTbeQNiIxSre2AG
k9m0h0dPH+4XKPzw9hD2UaDqFdqq3tfNYs/KckGNBRIovqrIoW4lfXVQNNIrKDNN9Te6ueMNWORl
ps5Fw4xrSdfaDiR5askJHFBrBWOCY0DkDOpQDIX28OjeeciTvzo0+IWEqvcd4UyDqLFnb4HtvVQp
XxkNTlThXNL4KcyvhbPAQMui3O3GzBMVceIHfevDIWzFmr7UKz9NpI4eavmocEDALMbYIurufyei
5bGEWgOfrbP3odTuH6BO3LGPUSIiM3sYJdcswoaXF/nvvMuCihPYLzvOXOLBKry4sTlociz55lWj
EGLkdvJNnFHem3AW9gTXC8Y4pH3HvWmG7Vk/fsIPaPfDUq8ocgECFlmNBYJgGTUCVDpl7+KMC047
W9qrWMufcyjZkdkAYEqzzFDKDricph0ZH604U3hkrmBn+Wea3kHPyh7UPJ2pIhicu+PaJSgstfyr
nys2NhEdGub4gtB8aFtnYEjmNcVxlZnNzqynpv6WaZIg6ZNC/I8NIqHHwemJSImU2ytNvBhf9za8
TvduFTWZlO5Lm135/bvWvbBZzC1coqHIH2VkaRgeD4u4n2H1Wyd8ZcGw2HUM5NQfRvwg+cf/2mSY
M1I2//C8dIP/of2FdgXeD+evCgTVPnvRJ7W1k8nv3s0vsGC7l5n1HwCgUh2E/vi1buAwS/sCESl8
Posim3HyxhMwd3IU3XATHouqY4No02nFqZFSwvYyuimpIGnj0xamxsTO/bU8LBpSgz+Lghm/tKbb
R5nyqxWOTirU4mnBirx6or9n9wghuL1iQhWeXTcV85qby8FYUxtePDpZ4G+F17p45ekRVoGMaOhZ
yQUyKR/C8TQBq1Bwg0pa+mViXSHvAVUR7u0YxjuQEJMu3550vYtdjt3YltZ29+RbSNTfhNu5mM70
VaJy/Y9pUv+lC4kzFKsZFlCr+ZT0MQonuZLRYUGkCbDfkGhSKuVEOxEnS/6zm8YMoCfoVIPzc1US
djSUCq9W/fvYs9Q6FhdOSamPRqy6HLTaH46P7KOOCesSnCmJU8+t03/ZLnlUCnAKOBHDoVxEOfxT
nBW7MqxrS31913Di6texf42zhpLaMaazB2e75CQ7OuWFn/pLGO+nOW25SybO23+x3KRps4jLiKtI
t0DRDhlIfxbssA6if87lvAkeNF66bGH9x9Tbzs7vO0rCdFhCtgjgAAFncOZ+ymi58J2LG+N1V1ei
CFrX1ctF0IMCDFa+IXb9aKOuYqaQNKfbKlsZuOvmeUCQjwag2ef7j1xnqE5kYk6BBcAIpiqyrmbG
gO3JuO/vopDVrIx9U1h6oww2T17vUekP6ab/8zj4e3HiXuKCLKvWwaRNz426SvdUkINboEMmpswo
+mmb1xyIAZUWgTpuF228YEKF37F4Ahpbjm2PwF9yDzHa4esFT5f0iwra4HMoah4RZVFiXi57W1aK
IdqbUgG7doojM2hwLN7phN3thbv+MNr08K1/zhDzzMaLwl5bPfa6jYwdboeAOEf0YWsWuGKT05RI
CfEDJTTB7b+AuWydCLC++NykzDkYfLrzR+bBoEIOs2m/6VlwIZHYlb2wYM2kpgSQlNWzrj8IUU6g
bzbV0SyTir6e15fUWHv4ttZe7nftpcNjQWvgGj+wf6o8650uleAOMzDAEsg6c6x31rwM+f0UlDB2
EBWiJB/S2cGSs9VlfN2HWBfIIbJpLBdKw56cYr4u0h62jHMUKeVwY40ShzLWmAiTZ0twgdFsoS+2
56BuM+6X0pdnJTzof/f1by9Iuqj7/tFUvIQiHn/pDhgx45PXEwIBkTzaKW0UnftYU6E3CaLNJp19
PTA9mApbgZJENT5f9VkDUAyyceVZ+y7h5GYWQt3oFNyqo6h11J2kmzVjxqpqXJ00AStGQRu0j+cI
ROg3rNMlXU7tt49ysQV79ahbVNGJSYsukEWf02OOMFB3t16PlqeQRFNILyaEqYxKZcl15bO9wzfI
T5DRw11/smdcmTe1NrhobWoedgP5DmEc7TI7Y0+ySnnl3cGZesfx2RWV3swamenghjLe3Mw4ayxT
MUFDAbNSXxPGjmO4VI/xJ1Y/FLk5kXJKX3Fy3GvXms+pmZy90xsA8lkzuoCcyLUCeFXS5F6lZd7l
SHxcjGBQZioNjILlgAJCSBXzedBpaNxcZYSIDhHW4cFzRZd4hJ++SNJJ3jREQPfKlKk8bDhUD91b
VFMWpN3xswsCtt6nWRg+E0S0OvVmb9dqm0IX1zbvihgswq81oJrxhWjagBKztU9IeKAscF4gv4Tc
qx8qweko4OH0RaGZlB8o0MIWKVFp5Q22f/8d6S/0bWRBriy8H7cBhDbmW59C71ZRBS9Mlqu5WWU8
tmPOuFhAZpp99qPWf8byWMovjZRqC/8sxM6K6skFMe6p9uRRgXb1mlpgCwLWSC6VQ+aq5sFRuYYG
gxq+AnY04n105slbQBRq+uN3jV8AgUfzvwpH7NeDE1V0nBzYDB3tXhD4jbERcXJhjh1VDpL+KmDa
GZ6cx2pDKm7LGEANmyDcarqnEE2cgcgQyyHVTg3JoEa5cBf9EzPFxrNMvJMw9PeWrvU6J7DozrL1
ttU8BlTFqbBbmrd1JpsolomdvViRsxuTInLWnRBu6/WlMRpZ0CSauy96LeQHqDY7iSkxMSM5yXk7
YKRK6XhkooFILjpynjn86iWrG9bn7nE+4iH4z2FGV6gPtDW4KHV0/NRxwAFRpu68nhEhZwj8YfJ+
RQUwDkhzFlAA3OrubrbRPLDTrYEcW12V6NolPDo5sAngKBtmF1ud22g3cEKBRyTAmGlUjAEkegga
xyYKypSX9lbsBHnbJLscONoDIMhDtIbOKUIp5KKN9TaL7ozol2zwY72ODGsjJk9LnpT/gWlu+Eql
vLOtcfoE0QwVg2m1up6ZBn9vWfw61Snd4ehZJWivPFF4aV3q3TzBD6Pqu1l+z7ddlK3meqV6vCIp
Tv0ehHEzBkESPyFxniZcNbilKumI7w8bqOrbi5Cfo8aKjctEJY54GlmCJfSfpiAV5Quys0CKnPA6
SIz+8/62UFYoa1JwR9wmCu6OY7TtjG7xMQ7wZqBdUosjS8JeqPrE9yy7dCarWQUK4XBqnVXw4+VH
MTZKYZ8bOHuwBD5Kdar9MiNwCLuCrYprDCS04lBwunzGV9YaKBJ9f9gHQYGSh2pJhVVB6c9ZuCi9
Sgyn+9lEJ7bD+8XCrhaqWPGXm55R/c3PtS19C4R3bHEUwsT8ml0ygAsxa/v2/+ihQUMan0gpt+QW
jsNFaA8fwCa5Vnysc8dDBTueqiPvf602qoha6DfuhFCsZhnjlL0d7rgQ3PALRZ/46bhSeZ81vzd8
Qy+de7E+bRgo4bjCRbGixC+QXlhuoomWMmooSHs4MNh2JhYz1Fuz3ZDZwzGRyyHDTfr91gJPg/QB
UFSGmmHKm1KtaDGD6+CWxZ5IPmrvzleIhgNNu+dDSB7M0Qn5jlZucEuD+4dbdbIeHHktTIBZ2Ih/
HpTnd0lKd1Yu5ZAdndeIP3NEaXWFWkZq7mnNCFvIt8r+0SIzIrL6vvrcng3cfRyvpM0gHCm0N7HC
sQiRUGhZOrdO7k0NYzY3lB/7oDdPuphi4yojSYLH6m6QM5VA538NF+LiHvfr5O1HOuFPokeyan56
h82vcVLjBhRe3RKcHR52mJMha6l6FhVMZgK6rlbZFf9yIXPYYYBSfT+/PAcQoZsagYAjG30wtJ9M
teZ3yd1jPrEjASlDQPtZGaNdGGMypuBKTLj1TFSjK+/Ki9c9kyEeF+SaVjVxHCZShAf4VvV/gJuM
PCmMCSqtDz10ez8ebLJPZgD9NzzUAMvklaS6dW0ZfZ4yo0hZ3HHQmQNK4GzirTJy8+fUXD/BuCfi
bKPbT1IvW1xMWgrUDLEOMO83/otvhKqB9/LS4O7lnBH12UiI/FhK20LekpaOXfVYLmtaFtOlogJj
ABDJWDLthkxMuhdxKWgLtsTzArfiGAodJ6p/BAkOu1CXsdzZNiT8JgfSUmzyUgH6LSB3gFER9FA2
l0kbfmwRzJdue8FHwSaX+kiADUj+ATCDZjvHUGwc5sllgD25OZQ5fIDrDbPi/V5Y/XVOEhSP/cFp
3HEUiZyw6PJ29wUkpYU7Hmt2tiO0os8A7DQh3iP6FPzbaHi8wjGfva7bjscL1MpMfBprDFx3y5us
W4Js51g+7Y12g+B+RwJLL8rN3bX3zTaG0TVbT+u/FyxA+OUg8TYO2rwpDww9VY+llbtg6LYWkC+y
ndD6OZIgp5J4eZzgEv2UpE64EgxgcEkqolPjsOMotcAsXh30KBX/qjIc6Tu6wVagvkLAWVfyzvoz
vXveJd9wVHKqmOzbMmCLurq2qNdyJRrllEmzMpb6aFyobx2XhAaep+imS1+mbwgcxjxDzx6V4Ggt
WIROyaYsCo/GxZ0t8P9mWDhMLqnYXAHVVqBfqDCa4BN5WOf5ZktbNFmNovL5MSoy+GPSdeL2BZk9
bufoWOgFqjPa3jWLYLdcjyfh04AWu7Andibj4Agcpy3+zyt9xguUpjyZgftV+4xMqXdozjZBqj5s
lw5JlhNbwoFWB6bmIeqfJ7pGqbDpSanjucjmkuvV8LMVaSxhZQSHAyCLyDUE5WmqbLzGZC5XgDyt
bIg9UTo/GExThO55yK/OSer/qrxNmn1wwT+r5HsTeIuHznJ2j1LVwQRk5OP9bp6ibZmXIUBCeaLd
oOe+uU7z19JUhd48CQM8rbr+G1TDRV0TiAlaJtK+0XmZPGNQA8UDl3kdA70Iufo46U1nkOOotonC
rngmDfW/oA2gmZJE7LYxEjdZOA/4JulM/AmJOL9JQUKc2ld9tW3hCtb7cr0GGbg0486vJc+N47kr
vu0RbkjTVfh5ay7TbdNVTU6ClDHxKSBE0AtDUAF3mgNNcDzWjsBRx9aaxlasy29Mr2Og4mXPcTeZ
1D7Rp7yEOntqCLrTpjhsZwQgtzWrkHDqaXDeQ+BMHHLkahumzEyuSz7GHYQaQ6WU0O1tvJ3/8qVF
oO9+YSETaUOTkQRLPpgPee8T9iBF6VnlbHqu5Kl9GSgEEg+1HXVqNE7AD1O4r9LT9wRE+ilaChkg
E5iDHxyUzEmVcNMXah9uVfZBpDCHCLGEqZ5a3/6VDO1N1wDPd7JrL9KjOEaINljwfNPQFvJHVKSN
8z9nnVRMX8jGoElgexVbnAius+r5WJi0kBwSR3uQS+9gXKlKoFdu+LhKOVN8A/26AZnS4dLUGPow
2wVmL1c1VqiAx+1Ud1PK+bCguUB4dLjTZ8uvrQteAdUPOq0ZfSj2ndJfQaTSPJdmjNTas0a9bcsx
7xa9QgtMjmIix7CWTo2OiLUX8pSCvnp2sTSCLLrMd6+s2ISps47zkZocOnAwuN3dvrW6R175+ZAF
EBDwVVpaqQfilOLbFL7ZdS4OfJg0S1v/GQq1d+tVWcDRsZdia/8Q/qSbHzDs+rnh5GO2lO7B6cvZ
PqrQBlAurhuDsVBMmL4jxWyihG7572f5dRKovrlhktsOIdy1psx8ZUtZ5v1YYNJDhetY4qThEZUo
Gai4aaWb+arN1KsdIVLFhf12wHUx0v+XZmJ3XBRVyvOqegUnieJu8F6ZfLQKvX8jAxnt1SMMzEjt
1+675Ju8/ziONudt5wJWfBC/3jERi9z9CZFrIylhcm943v6FJS5zqObb40sMKvBFhMXjF72dN9r+
AfmG7PRYFgecP25+I1wMj6rODoU4bgjb3diPWAaLlW/0Nb/HZvUxkIHMS3skM22ixndQwCEsCKIS
3rPSk54K+borYQA+TRZ6gHneQ53bECANe6rKkIUkUrzuviO4Ruea3qiUYdhkgLoD8Iso3yiYTz9k
K615rSimQq3IKXBxgXCfn7SmpDWwWsKTVTzbPCBC5UlX7XkjfVVrHG3EJmLUuOEmY7W8i2OSg497
0koyWerdlLGL8ifYoca8qInsgPI86JeHD5nsnfTI+6A55CtQE89pOORUxUI6CXEgCCExUAfB1tlO
YRgUfJS5H5uXZ2GFPH9QVYbfq39En/qkiBoyQ1Ti9YL6epSAeAudsCb0BB5lL8ji2qYaI1NfXS9Z
BB2/VWEf5qtktus/XOfjaCgMsjyH9JCbVD8auk6u8eZzSgNe75HlgbghxG8hShte6518qdGId3n8
7Yc+5yUZc+TeZdvkR10Y41P4PpZ06DKFdJWF0joTZOURX3jY+K81Mbxqx/ulvAbbfrrA2iJTuzqU
s/8coc7wN8ZvF2Avh9bkTqtPGHtn3gYK9diL6yOs3yhi0r7UmuNbBl3cJ5JeXxcYMuqIEcN5JRp4
yyi/25mhaR4NV/YkEHAu7xjS8sY8JFvzKudlQrsnEyboVMbldPOUAX/tiOlH1WTuDFYV3NSc7TEN
LebKXVURugSiM+Yv5sGotacTnQ8upxtIzeQQbKAdWx2qoCSIh4rncPKGjGS2woooePYcZgwXPiLo
d4MTcaEhzMMDblEQjbdBvfL3SUWS564uCYlHOmxyXsCWGv3NZH+5aoeKCmaR4O3jRKdCYaQhzllD
qUOute01ZTOQm70SEDVRQLEgiq9ZrmA8bfB8yWClvyT3EnFe1aFcb+DEFr7YiaTSfftrWyMvFVA0
W5Mscr5OBmAbvwCEC2ESY2hUvvKWxAy9JN6m1GUeMuYj2j4R/0SpftmNUX+RCS3ToI7/Amhs8SCq
FZWxjgWKK8jLh5Yqa4pVaok65IWBs6Akv9o3HdtRsT8zuyApXLsteCh1/JrEEHlI1DyZBg4Ux8OL
5C8aozt7r5BSqdtmUut/dwnrISTEcEQLVBy3l9MvPpIIeEV9jtR/y4daIUvIDLnXYsqvBJpCXH6X
MUps4on7zzr0FW+ffucLlCudeRIKJRgSRiB+YFnuUl0myjAvgrUlnn/aMVpxoIV7ystRWRTct6Y0
B//McEbQ/juJIeJis0kaKrCYItbQ6IbMtHiJCUSEeaE9Go9Jo+8wZIUgVPJ/ic/uf+6ZNS0MmxDi
yghIOKlN0f2Mse0yys8phPm6I4GIaN7N27ZrAd867xzisD7574qgAqEsJWdyghBfd0+LvCebkPpN
B/0FcOQjMf2kWcAY8dxNwr+1fVbaIbiKTZ+fCWg83jmwuRrpf1+GXUhULVYGFAghhRsX2qxXQVRO
82FtB/Q8ZDv7vREaO58wpxPr0vQ3VXIkBJpCNCFYsufja807OPNN1VzR08CT6Sfz1/WASD2TAkC4
rqphxEy0nvgE2ON5FHmmeA7U3myRTb4qXKICnQCf+ZBzvjzQ4SD1HPm/xVrM/CCvb1eC8RUbVQtC
DItik4k/MPiof4VYGxyuWXsqPlEEeZO/UmK+Ks/0TneoLIGVOhZ1lS1pbWzYlYlLbGm1R3SQKLWY
GgXLhnTSdooQrhRaUr24yZFLFMcHz8+ger6vSBIyRo2VYHCGT6ELKqbN4xANq8pJWykomMpopdMt
fexQS3XSBDEByR7umeOC3MvAdk7RRqyBN2UyQ8B/n4XtgEwByLXaIrx7MXisK/HwYtTpJaQaIt98
PPWNy1yGX245y969mKy8Z9+ze7fYrkIgT/wqrzHDwOC7whRQIFj6I3ccDEnhhqmCC2nOZdgfObmW
BNK4dQvW5c2NTvncYBqw8u1a6NQQhGtKlbfhuXYubJyBh8IckifyQikJZ9XtHSeItbPwmo5swyhR
laJncN4Tp9iABozL75O5ubpZRixzffCFNB0uBppd/FdVNHQ4+QEZWYYSHLR960kuSn9Unj7me0Mh
3jDpCm4vLNlwVcHzxSRV5q/YKKDzPPfzWMlDFkDwoHrXUSrZnzYgE++TAOZ4qHxhhydGa9iD0+Em
eiQ4OxW1duAVQOKz/IlVwRWGI3epG9rkllxsx5TpAxyPD6HPWPzHXJ8pFE8Op8+Wa+oY5OTRu5Y9
oU0rzOLKgqDMEfJvajz3I9dR3Tv0u+yRhlvD4uT8nsc4hFOuAx8KRchtdA+bkH3RLPVygry/ORng
2WuKe0XHx8qUaLB12SjEvwBifMSB7qpPttBYry3RGQdZqWOYcGAxXLkz2Qm6QRyegc4C6NIC/Ojl
sRK3ISvKPmNQLIIFG+3YhVMEbscbT7rYtz9IokAgIqRj7dxHhwCQfBHKIpTM3sQaMJgUNvAKdZBL
UJvdPYmTxEnTNtb4iGaw9UQaafFdOY6C4z1UndQkcWSMOce7E0QifTaRm7dXqcI9ns1rT31H0ukc
DuObbb1npL/WWho8GF9CBYdiDmjt6qfdhBSpcel/E2aWUljqbINx07mPRSLDG87qgufftqqd7vwF
gWNDygjfbPes/JgNexQ2Q/HKtuRiR6vFOs7G3VKFRwVjsZltnFr1i0U6GJC7F5B1CEV3Lyp1kWAN
z6QPsvUlIq9pkQNt80Tll5WerVOnzVh3zxM37fQ7Rjj6z3e3IXjgG/pZ+967ydUNK1Rf6JVhXuVC
LaOOCFx4NhGkP9gZiisfS/4Dm4xQsUDyDoRdLlovoyfiYb3PhQByKYBJW2tzsfGNtTEk60pg/HJp
SNVQgwJActjr1PK5rh3ujfUs3MMe5Vjf7KqEhBVUmNaOgiXFm9HBOwAj2GQ6+B1pKbu12QcOxilr
hcu8PfogWxPC1IFdUvtd1HqxJoD6B8k63zlTjAHYl2UtsuBftmGpGxmIXVhTqzPrvJvGMeMrChqB
Iz5upAgjXoj1UIcPnmMrzhByN/uJSUJ58yjX6ovXerZFHctDG9ZjWzGbk+LGF62GuT7UqEEstshc
ZFiToPUyHFILI0HcQS/8PRjgzmTFrWzQt27t6wVZcMUvC7auw96Xem6SnMsMIdRhftthjy2Dlcvy
H+pEKstlSFW2dARogD8aIEV2RrQXefXVILyE1zH+LF8yw8Kl38k3f0ZkxyT9r81SGVwxcJLdnCo0
AuLHpqi+yqru2NiAyInNhd+4TustkH9/LPdvgFa8EQRkTGDHRPvXEOeJ6dDI+jUwI5Jfyp54Bv65
4ni+m2EiBbGdMq3gyQpHkKZzwa/WJOlR+Hf8Zhez6nCd+MOVRnXfHkgw6OjJkGmFKM4H8MFO2c+J
mjDKWY8K8qG8I2AszG5wG0KPg58MBFA5tk2OzoCFPN9baDcewuUSOaBIY6nWSGD42HCzXAHlmYIC
tZTlThRYu5wDmjDsXThVYZWVlkiL9N/Wx6m7a9V7wW0Euu4+A4Po/54LgIlaJ6o0Tn4AuKhePDd2
kK5oTbnbdXPTWkO9eDtXNV9dDHftZ9ZNXb1PR9hpeghWbvs0oEYbmQUpMGCpeucbbyEFe+EoAj5F
4pjw3gzMwYaCNQrQtuw9ZEFw5g0CKCFNJYdorsDoSMuGqWk01/u6loGVC7Dha7+douFnlh+hx9jN
4RNLudKx+lgzWyM4j+9+GxzptOF8G/Y4bRr6v62d79sOxUJ3p/rNwkfsEAP5EFmbg4JYS3DY9NT6
JvzDFRu80AyBjQWIDiCmYYQF9bToT2DXNBtHRvbxOKSOHl/7dlgpdSFvvBpFJXCaqYAIAHh6aWFH
Zm0mj+t3TZVv3872co39h2YTUitQcL5GANieMARDyD4qSHWoa+M+BQ/Z9hCoiJR5v4mcsOMYAbin
z2fxpnj2C93Pvjwej+OkEXqN3fsr27WRkkJ3L1N6o4ntEbcKvdVeIdmv+R99HedPi7jm9ZYp1mRX
ScvAhGZL1RzfFwoaueVQCyVbeAn0v/ZIDv8pHHTXnHP7KK89MNBMQoca+CsbS+XvHnPgyroXPcix
jvBYZOg6QFHSPBL1zcwY/C0IEATOb1IqfoD1YVAbpgcFDyZwQGQXq41EUwrPI44Aj68UWSHPRG9T
5czFkxm4cuz8zMVx2W0yzZOtDSR8cSz+EFZZJ7dImZRLF1VZNylF/Y0wnvbPuRhJKhR3LANWRs64
njmzq90cDSNhlvbzMsS9dB4IWouVOT1zjmgpbWfjAbEemhe/E/TwXbbzJzdnaK2EB3tbEjsMlWR/
CC17oO7v/J+tGo4bXMLZ1iUZAMC1z3D7rmwqoadZ6E1XnuTDnHvWmILjr/Sh19HpV9GNF0TEeNOy
F+bjSlOeqCADxFv6bFQEynRfYN/JFWMa3Z6TTAKnFwyoD5Mu87znF243GESXgh0//ZNUyNIVXM0x
q+aGkpk6ghv83CXo8WTJFOetcoqZ3FpQPcebGZETTCPQj9d6vcuAwmy5EyvD/kGFxhsFXG8ECOlV
qcYU7wH24NK2u/EKuQJaTFByTZhGwX5lhPwKpGTIRt21rPsjELMEvuxXdRc8hZlYa/WeOpdx9U7Z
YCRWAr4jM5iTbtscPPPd33Omu07iTaKkoUUTby416Vdg4jodv6x2VgfBYcF6m6mIyrVBIru/UrI9
U8W5CSyA2OBpb/BX5V9wnD07oS1pOogujWaItT3BS14vi1opmd8NNYKr7WEpWj5Bs6oXA25n9SP/
CZdiF8JHC2ThhGCRxJn6HoZ5Mn3sVLIJW3IYcRUHU254nDI4qiF/KjIGIxs+UaCOBu2lCpae977k
9Ijg7pXzvoep0k0h/3GB4mouS5+bH/bZTBETpftoWN8qlC0nE2v7mCoctt6mKrmTmx61F5UWcYZP
KoQEX87DSYtclt8YzOlndrvc2Hqf2LzyyUAv3NkttgyDhlkzN0nErIWamm0PtcBElnDebRBWOhMZ
gMkkiLfALlUG+zxiJf6pygpaYld61BptlCYbh3SkXcrcIleDfcU1Fur0vYg2zTH2QhMPuEBJYcMX
fSOQGTicDg0+bDXAndvqT2DSnU2o42Y4m0yL+8fjTdUCTqtXALAAWWqn4adncGwAEr1PJBmmo3/+
3KKCFbd1yNMWTFQdWNFbaN92Are+JHGu1LOCwtpXGP1wP334JJ8yG9puHSflZV0Epr7muFw5Tp4K
ccStgbuFx2frd5TLSsk8Pc3RZZzyOr90QK6hpvqR1Mb4CXJRMNNcmutOBN2Cgy7arSFtymEgoYsm
/uq/QuyXipQVtCtGmhagLJbxZw/GymwAMd64+3OHlD+l3B7jhepHvIDtTjT7OvHi1wkBRuzYWKlx
npXPvC+wGrQHIrWN421qBRH8z8fG/kEFlFnhmLEeqmFI3Gt3u6rfJEmaprBedpQoN8VcHIJHXgwJ
EPZU3PBP1AKjn2tTkIRglvZL7XErGr4h514gpACg1nRFX75yZiNaK/8zamkSlWS3tbDLD8pNSOfJ
kMOKOkwGeCkMNaQyG0dkpN+RX9oiVsUsl50NEyLNfNhYhlW/M3DyAHiFuoOk4dnHxK+KjDbnY+aT
mueeFHp8m9EZRWrc2EVgIhVV9uat4JxRa6i30b2yMK2cMjLe/ixQ8U/cDMDJGC0AhE+mBEmgyM44
h2KqWSMenTqnNbxzfg2CqUtBlPWog0MSZw74SvTNqaQUdkimp6sf86pHUR1oz7nnJnW+FMkfEqnA
lY+7NWewW2moXqpMbe7Htrk53xSMKgwVdWNJtux2uNDiIuaLUApCxaVlgUmEWhE7eeLIceJId0cY
cHF7T8S94d/Tb167Z2VAGyxyOPgMR+72QrZvbZlhQKZQvQ5ie0O5QoZ0Tp33H/+yd1jG+s4sr14C
P41f3+YzPqYeh2t1/YkN19bRCpJzVm4bmVOjRf9uFti2wrQQX+0qdQ6fkXLVBsxvlIy6ub+yeMrQ
aq8V5Y7UuXW6DvrbblMoM6qsIGTEv0KKD51cNPAvbEyUAjlFd2XXQI0supH78kvFPHXUJxpt/047
yBbc4DjuxrKq09keVOxbSq/9MLYeJsJ5wE5xuJ05yTLLhSNS6juzfObJ1tXxFU4/aK6wYYMawU9a
gViIrsnYW13fffOoZfgFJFfN5yu8KOVYRd/0ilXKmHOFcbm4zyimgPMf0YScfQ1Gra/8Sw7+rlO3
y+7A1hwnh3l/q8el/KCoGZvCHyrHYlndR+veZuJy/0fI3/pHEZEayOlwoHODh+FnPK2bzAtO0ByV
3Tz6cawrKnKd1VsYgVwSmbuh8HyJKMcL6dyujJQT0S1hHhuxU/WMv2R0jzcvbyopcSFAY5DQPQLM
PzTwkwi3ZGXWlz+S7tUijBWf9/Hs+kuddtk+/2ixNNRxG/9aR3qx5qY9mH7vliIUEqUU+mk7odUu
5Ex4LKiAgv++GoxKpNcnVUbsBlFf/9YsMIoW08g6gM390/jzFOf1d9+yz/7ERJ7w2Q2aDTB+bGzj
W6oCzOHk5J+v3Nz98uMWyBqP0h8x54YyP9lchTPBReb+XvTplv1J7QP3mkpervJ0IpgNCTu9S1gd
6b5a+Awr5hKIcfdwl4fpD30ywakd0B8bVbbt+/ComCV/J0ouqsmH2tmucuYK8prqE3doJIrlv6Yw
rEjieyYxDKhnmwTjJ50FpeDU1jcFgq+anosNx/mLenCsBTpEX9sO54lLBjcwEjbK+y8N2vMMe7iF
Zz0XMqST6w/wPuO3sYN360HHidBqg3q+w85yXO7BaAXQCp6Chg/1QNALNQKc+qBqSD4PfK/tfMCY
pB4c2oLPObUf0dnwc8hNE3GDGotq8Uv9B0Uv+DB9yMkXF7f96m3xcFQjiJgbGu5j8dK5ncbYy70c
3Qp3O/cfUtWcWF/1Xh9N3r8fCqgUc8+93FmuWuQw3xGLPjSZwoqtCjJOV9dfmr7h4HfhmT+KnqAg
Uo5cRAXJG/R4C8yGKxdp8sFtDxO8fl21JvwWQZJjNr/XQECX0BwTy2WuacTnafe14PRoOz111Xxy
mBHrlvWL6OyBIXydcI4WrqRbVFcwk8EJTbz5l93OiO0m8EF0ss0uWyahf5A/qJcbICmDhkoylrQ4
8SZFId0M07F6USZGWF7AcFEgjfDmvXt4Az4myhm1SvqR00wqEsOz2E6UrDG/aQ62PCm4MrrNEutB
uw2d7M5Aq3JLlmpJwFyoxQWaes8m6BJdDtA/jc3ktsOQjGT30Fdhimi7APE4HmfVnOw1C5aCGl+k
6/aqHx9aCP3JDx+GTSF7XyXUfHQlTWYTZ0x3VabSrDmVcdKoC1/d9Vl5UwlumPGRUgbmKPzE9/U+
y3ut1edOQ3oc2kZOyxdoo8CI6/QYhHbweuYr5O+vo6udCNe3ClrodLg1zSAZe8+a8kBLMRJiy3Jk
A/2QOLt8bPzQcAqJk3kJbi0DTfdJCmG0YrUElExubKRct9kvX5KzCZeAAdyhzUmG4u8n0WPXIaIf
6hSULl8EdbZoOwBIyW6ubuJgnM7ozlrIs1dqxpsbnj0j8I0ka6WLOse/YN7+T4mC7UAkDGdq9uk8
meelMuZWuUPLniCc7eUzTiiKFjcqBXAKVpMNRgNEKPpTrhKU3opBnu8afzhwl392+Yer2BtaQJtd
c762CB3ucpkDm56dLuoxFlMjluD0TgRS1LVdp0Krpo68cZlT7liMqweapuzIoYmHhUIPYtkBdtlT
hqD11fFZ1evwaDRi26fFmhiJehGqZ2BVOqRQbB5rM0rQlfDgRFOsZYu1KixQScpHh9o/HYih+CLh
MC+JHCc0jQiQ4BupPqI3KlnY0dcq+lErC3dVBgREqA2Y2lsZMLlaQ5HxNIaaJpilFCY46uiZPg4z
aU33oWhImAOLUQ5Q4AZlkdrx5IBCZGitOosMMfPf1lNlMAmNRmvI2qbrTnFjSsvJM+4NuX/fG+c6
OQhR3Ekvwx2lSwyxkpBpYcET7T+w+Cgu0x3+H1L7XZq/3dV+LpQgmgSdULYiLCr+aU8i2UqzyD28
xaDppJ3mvE9MPpD7s7XBw0ZltkvudoTuFWN857yGD3Ry00iZ3ECuVn38H5o8FEeY6YgWcOSBDug4
mLlQ4600YeIi/hCrrgAQXjdun1zuYYw0welzmkSJOW2FQHLIDA+V6lmkTFBsuyql7mx6x1Q1k4nv
YaZcGlpAe8dsvdjDuEcF6rBPO4j28kicWQz3nuSYc3O9Tqoshwz93a3PnOKkY6e1J90s4M9D633K
QlRz4I7TIxOO/7ZXUGbBGXXFGXq2dqICF+JaOhnJaRVwtjQ6j785+1q1A/JGpv5OlGc2qBbRODuJ
pit4dG2p90Ko7mzP2gcafsPIZxKhEViDq0u4dvEMMSAHJmbx6Aw0T0yjQhDGawuae7RGARJsULBz
iMe5NyMzkBf+1GyRKQhdG9JN/uWlBJN9lNaDFDQSIF39jxu+Uqk9xXtpokslm17drGUINW725MvI
HLs27LwsTaZuyLt7QFpX7uu2Uz5ML+8/x7Ort9AipLjJ/MlGPZF11e/rk89urIzoFQlNioq1eurv
ZLwBrYBfaxKV4Pg71xpFJTXWgtZeYPZf/zFr+mGB7NMQBHdp9EIf1SLqoe52Ud3WZoCSSEKnnkkP
og+jC8CKbAkdofJd4ZX/v9eYZ+060r79Qv/RQ0Z4CUawQRzOyrMkKApd5nPdIO1XXPGLFDU41Qmi
E+7lP3H8LcQwPG3b5g+IrdtLpsEG+VlKriE0xrvyHZkWpB98XlEYzAzRngD+dG5hliSpOOaZK+bC
TKQKR7foktm9y2VeDRg3Ov1LZamQ13DEcgA/gK0FF4/3k+JBlv++L/EFsaZ34Z/VkktZoNpmK9is
zTvh2P3U2OI19bg+B8zmqRqwNiRfHSrhqbSscztlSUhAZWRI7rd5ordXpmy1dBxJSSjxLgZ2+u7D
0ZF73bw35oyz6nH3zQwIyiTpZOdl0JsOAXuDtMLoCpVpq8/566W4MEy+ATEu7yYRiPAHrzZLgCo/
XKeBV4qYPyv+2ZkFenhpa11bZq6ZfoxUAKX7EULUHQfXtIxva32GaVvDzRQTE0Ui1qyOIJKm67I3
7wFUikAhjgJR4A2Nqr7DaUrlnOhIe02Z+hQMIuGCDtaXLkvcIwGvUscTIkUBH2tyH0/iUu5M6fEm
NROaIYbY4Y/UMYNp9pA0KjQhwcxL5QsQg8CBYzQ2edXDLkpqhmYJkaI/KOWw6H1mimFFFOko+rnS
WsCZ3GUNH/7y17/TF0VUrPy8klaunSITS9ESsrJpM6usBYHgY4ByuNcVkvWFvcEfHcytucJ+e3oe
yBTW2ojKGAn6jbuupKkyGAyi8rRZ+q6/J5V6WBxrRd/pWyqX+mj9et3u75S40SLVomsfnapHf8TN
mFIjDNALGnhk/IeFwhxREHN9wRJ/n61RRqRlQQMU/IIt87CScMF0xuKPVI3hZ2b1CtWd9GN8MawH
QxYonSaETi6xK7cec91mCqBJVZJQweD7vrbqcabDYx9yBNYsABfxtI9yJCObbBOAVKbzCJHegOvs
7mBYPDjmcyW6w0E+50fWDl8+LmIifRlziArWByRH41yI/CgB5L8/YpEy33rDXQl197jWUW/VUbMe
RQToAxINztg3IjT04WmtqxcFFD9uDvRsXAa9KfKA6qMeiROB0SrPVrsgfQvZ8p5MMAQfa5/LExFG
6Ii6+cCJddOkb8PyxYh0I7iXRwEdTwGiCdI/d7PnMADJJgTBBD+XQ8rDsA3OdUQy12hLrlxv8p7z
SjJU7lVFhxpiH0R0sEWYCLAyzp7LY2tb/C3D7K/p709mtPHeQgOcvyuGjZ6xtFvocU+I2lXsqtfv
wUBbY1i1DyTrRSmvgm87HcBsK/EhYnobvT1HxgNy5OajlIoNrbnQFbs7UB31HRpmIt6p4E5Qn+Dd
nMS4Ajia3Ghy+p2JJTUVudu087pTh7yKOe7jjKUKs4uAg5xXArR5ETypv3aJdXfQxgJyNUh9tpGT
k8yPaa6lM06qyC9+ni2FjwXETXBlYirfp9MEs9ic/CTXI8B1d8fXuNJ52Vj5zf8b0g5MbqtiPqwe
w+7qL4qK/Shq5SSa9Ql+K13uSgE7IIg9c2qFU382ChnkxULdCSaJWp3Uk8HGG2elh3YZqIst3ZvN
CEQ/Yc3KzCWvJRg6EKkPHNELo5IFhGOFjpOBe+ds4TQyiv0tX0kfadEwC1FXy1YHKR8xD0nS5fFW
vZuxBi9KhoJXdNB7znihBn1IcMp+8PF2LFw8EFN9EoWqXGEbVv4BY7yewJkgfrifLyYxsG7CCFoG
ePwOHbcCxMmdfy6dngP98ApdVRZzvzmNRZpF+M6DRPF40eA3AjDUZ3Jfk7QK4aDVrk96voN9jVJw
zYfdFjx/aYrpTTXxnYjt/Rqp7Ap+N8mUjXHLVF6ok0XMukNCVKy0y9ybrVTTLBqSRBHXcqefATfP
+jv6rqfpOFm1oqwu94rm2AOzXnLGqd4SY7vhBJBa+hNPvuF2OSdsi4NXSgyaeX2eWftJYdWOm10i
I67ctb5ITfD+PEBwxbBYlfXraCAHHXLMYK772Pslz2cuYC+4ffEpYWYt1VIv2YXvG5ZD47EpnVr1
IL8x8razaJ12+ARxefoFCnyedBlF8io7Wi/uHcwKYcQQOtI3ZMJyyqfVbNTwESARl6zirsxUdBTd
9Q1qVhKvymlIL+oyE4pJWmQmSHtWN7Tws/DYjS85DYiHLgURyYOMr1M/EngERUpVT6hCzNY4sid+
JEYpYA5/SQipkbF2u+gs09Hu2c/EKISrZzCPHvOmaRUlbSGaU2ug0MOyWZeWO8BC0CVxebXh3S/b
CvmePd3FPOi6N/VOakNLVnSf4COH7N1Ha2lfXUcwGPcEFVb+uvuWiJWkobWhRwYoe1ulsdsdsn38
B3WhWasZUhqfC8PGtIuC42EkE1b6euJuQrMxpA6XvGIGkT6qXseS2J/a42YWJa4Tb+5soONwc8Os
VR/sYYm98WMcIA5KZXGK1KvwTtL+YS1QOGQtm9IvTkI1IuI13Q7kbhUYKktYgXFnxKbHDCDxpRgz
X38mqA5xkUiB+j9W6vs+eM7uXrChx5oblfk+jKQkc7JcXP9bDW4xSTmEh7Jawhz5+rZ/a6Yw9Wnj
eFEEeLpH907osFt0OqIRo3a62U2Lmh1H+wx+Pq1GDb9wVphd8UyPEtkq/H/98TOB4b/MOoLXPueh
CE16YgmC7l8f3genVENfPSSufxhQCkVlJddAxr0yR8Pi0f0f8SKeMd2i9yM/WVpittFUlS9Q6udw
2R+XAby7PFWYxdEaABu9vQBGhn4W3SJ2D6eoQdk2NLvq0xvG2ncilIxrtqP5Wcx5BebjdPkvrk6r
yCLqGM2+1dxYFjkFPBGDn1pzHvN701H2xLQxrTDA3ZLhkmQel9CfS+JPCv3SQEiqV5gB4ajKDhGe
d+gsBI2p/xMU1YNE6FPwhkBy/3bd9fhEkQoerbqUPWg10O05SLuHY344WF4fsLwEQfrPncFoPdpQ
oey2hztnC+50INHDUCCUVfdyzI04mhv29mj31tMM6Q163LO7Bb9VkMUJ3p9BWLbZfXL6S3ohUtGl
qJQJ4PhEwM4XBoTMGR6bX8ZbFdNtKpnGAdwIVeuRr00DWT+L+vOR+PlNA6wAu65r356UwWoXP+OP
4Shy7MHdAICEY6jXbp/9CRYspwIUC2vqzgv40uE3Bg8OLBbIeYJh92ZNeBcYNeZv+MyVfJzzVNGk
hlceiytAyJc4yMLPbfqM6bBSYJnEQIPo2w0Spl467Yk4dyuG5yCVSK9xgDpoY2pj64mjb+uHeQ3O
iXsqHbaT/a7heztE8iNTpDWKS3jM9VvUDIhe8h9G8Yh1XOR8WaTmMN5m8PWtvQBNMX/lmszXk5Jo
16vEPST21mPq0ZB71NDqOcsJfDj9T3YP1raDKpoGInZHttvphv1ovSjnikZ1tOkWJsdBrx9IxbBU
dpCb+6gNiJ4X54FwWmU6k1UU5kB9DQDFB1KuujxJ0Wyn4zzBspWTDQ8hSYI3ye3zbzJeZRm3M3Pq
kMQ7KhhYy9zT1bb90Slg0YIBfJjCv7od4FZwZYaFS/GhQI//ja6D6aQoL6DPgCZXVIYbhLFOHWZ7
T2v09aYQQiOhJc3W49MAmOR+XpP1oxZg3SqOlO6C2SrdOSNU32YpqCjyBr4KERlVwFxRTPJQvbZs
uuYtDzmLY7aKNtKsaGctpNTw9TZnGAe6gyDNUhFDJ0hWaGTZ8cv/A0smfLuYK4A45ctbphwfdl2r
sxyFWrto3JWaEPUXgl7DBkxf8+rG5NqJG69YJP5yRs0AeWUG/xgbDALQ1pOcGu8m4T8rK/iPKUqn
NnGt1J7JPj2rO0GtqsAU/lrDG9gHPt6crTqD45uHyjPAp+h+ngR9xncb43jduWRpr3u4wUqExf39
WXJk8XU1M+r1MyL3yfqjnUhmVH+aRhkAs3hgZJrU1AOWT7P1j5PPnUVexU4l7ZUII7rlMuBL2vnD
I4/8EdJ7ZL/zYc2/vZQXBPdnJDz8xEdETjisxvyPFQ3wh1HxKx616lQ0hDrN5yVTinYQQFeHd6L+
0VIBMhL000Sdu8gy6knKK5fhUERHGvAAad6jhWsndT0VqfHyhwP0Hq37YITy8BDHSqLKo04esMV0
6o5/F1ilin2buMxyImP6vrANp/pyeixm4BmsjGhR5AF6USxSlB5aVplgTNliYftrvknaimMnnp8o
gzUpdF7A+DyTPszlNAs34mNR+D4P5QOJsEPTOEcrCeViWwLY1Ga7rJqB3PKmb+ApylhoLk2+A7Ac
MhlETrVaLo+ncUgkjoS7V3uKnRqzLPtJfm2NV1Z2EWgpFouuLwd+Iw3haq2bosVC4YBIfcWi7tFv
ql2GRb84L8UYxLDVzwhWnRO9IrDR+eZqntCpW6ZQSHZ0j6BFxq/02Mpd4hrbGmCp/vKrDlVSW+Jz
LS7G0AuzIb+LceVvA7aummaDueBgojaWWaPuC6b3As2hF+HN/ACqZpCnVeMQ+UrBKtHc6SOdtGv5
dgxB3qQ6W4bx1T3unx13iG49LyTMp0/9BwRWzJ/KpQDGrZ+dZgwtYRNrxLYn7etPakpXXw/xDTEN
i7mTB4JoZctW0VuRPRDqzYokN8HJGu1NyYORnwcymLgoelg4vs6+VkCrqN+RaiNal+R2dgUQpUC3
PPRgjApTiNRi3V7TsPg98PITxHpziJSTg5gMP0alSx4PRUwxSopFxQW5hhJ3CAHQ6lfMK/1Yqq2b
MR8dxhM2qAgaqwC6o+qerWIfJefxKe6Vj0P0lO1yXiMsqcTpEn563NNEkWDpAPndGb1SSWRcP1IC
xKqawThQ0iD/eFqaYo4qie0L58ysOt2I1/N9YZKz4w8sVUxvUmFnon1Q4acTsm+/F1Y+f1PWYCO5
Q6AqxMw3y5vfohXwdKtFhDArkX8/aWt8HBezPbKUhfVXFHMkU2P6L539qrpC6bDCgSz+rGgJHFKu
YcKB/IMQTajvzLXQDhKEVNHVbqx4G5gYMufouI0vH2hf8wF3Qge/8ROXTat6mBkHSiSb9lhXkJ43
B7HWcxnuoEGtPRYhEX4Ic/vJlE/n/O4h2cLHHMhbVoNXuC2CU9DemyQY5m4svQtezl/YQuyzeyl0
EjsHXkAvJ6wTzxMszRu73rtNCKT8JIcAEpnpRz5+rJRh3kxlhoHyW3jxAgc6SVhp11yAA5mXZV9E
rbOInCTIKnOiLFDtqtYUmZgvKFV2W2eLDRocqwO+rx/QV/8HXgBlr86P8A5ciPhLRLlAQo1pYM57
SuR6EvmvVBcsNaCEA13823Vj78Upr7ZQVzEOADgR/4Tg+ltEfrpJ27MRYPlL2DjcUtIriUz4Kekk
J4zdQJVvYZoRgsJmPIV5Iuu8PuP7sNiXOcpawIDSpFUC4R1iA7etmAKCai5uAzhQ8EYav65Z39Z6
AeHtw3AkzFe8blhCEVPLUV5WK4RX/bapyqxnN8S4nvS6Uv1jJ+9sAGHSY970Z4hnVXP1u5runlpP
Z7ZL2eEx4x5IvDBQIVoYq5Ly8G2TRvSB/fp3iUpD1VNnFxt1oe5Jz71vgiDpMptzn15ClaQsz+c0
EZQ1fVgAmiVyPQRTWN69AInuFc9Au95flC7jkdEPaTGjrR8JLcMX+o93pRGEP+S/27qkrJFftFMy
NbLyRHLVZnliLoJNjm0vBc9kMrmtTuOc2U591E5q3FunDhorclv5UtZfWWv8OfcblqdTCVVl0e79
5lvJ8Ua/DJ0zxWHSVIHjixEnejyguyu9VzFCZJRU/GNYGUHBqc959LYBpNUgT3oJclkY0ZTBdBTx
9T62gAW2wBVQAiZubF3lyLDSFRJ5fWO22tnd5her1ptBzO4kTpkEa4pIFbTsU/S4HxQtAFBi16Vp
xTaABOlBxD7IFLOmhYHGO0mDrwjgMbYb8R7RphCgjei8M/ZM/FSgu7ep69RXsXfT4yqrSRT2zvA8
D3ECSNS1+Cs5jAm5fnU0gVM9Maebvt6KfWdz/2iUDkLHQQLYLyIA3ciFLihGroR1OMnUctWDMZ6N
xEjkSpQJTLetDO9fJxIdHjGekm2uGtmM3OjbAYioCj18AvgLSKEA5Y5tfHdD5dfJ04khAt1IuWLs
szvtt9OMemWYVv+6XeHgAZ7k4mmA4hdmxkkmfQUkN8DMh2zc1Fa0O80gV4TjayCyge052/qVL4US
EmdjopiDa+3Y+a6FVaBu6qQYY4M44KREp15KoJ6uTMeqRARzQhNX2IqA14mpLGfxfFVLDUTaP91L
DsFVtY8l60rJ2KJ1MHlOj0XCIHqciwGdicG4TnOzkFShyGZCMqu9ebbAbD5JmoE5jnYGUiw158Pv
SKYkfQzscsU4h9RXfa2gNsyeD23okFUNQ/ehYMsChEXKNt3VWLRCFbtq9OMRh3u/hQsMqS8mwbPW
1motW6HAKBSn1ny4RPlOskKqWWjLeudpgFb2STIy34l/uNH6Q5n0AwkIETuyQx3Y9b1b514hL8qt
+5Dz90mZtEnCbFHGCg8Jb8WOSRrE720XY1Kyk0QLrgajifQZ2wIBA+MOiBYdsdi8lJJxs7TzDNBZ
tzrWZSkxYngNykDfuDM6ui2zyllwmTKIMG1bVDssDC6aP9LGEdmxHMFkY1l5/6f5fidNrkbI1mE8
Xv/RrFlPVy/o0GekyMC79A+eBbwhW6LzquAyzPG3dCE6zJgaZon+dl5Yju2mnvEdmvr8E59aHyrX
aGG327hlXypNsrBLGXgkD53hIlnmJVO8d0KuzyB8kczVOo5DiCHtF5YwdywaWgc71gvqUoUumeDn
xuUuLm2Xwx73zm2Zt/UpTvl1k0EyRv7GM5eJyog41yPywh0mCejMDU5mqpzH/en93a+5718yPuHK
Cc3oHcOmksJtKg4XI4b6Nd0uzV9gIbocdh1b7cYbiSsCNxp0IQXE8dpIvDziGYXAe604OZ68whAY
IYrB9ZLwYnbHVwBJBKqULgE4Y5/FxRN3020i7N3s7ipyNCyRGNdFTh3092YZHzxS1QR+gqD0yKvR
tHYZFXLSQfeRYboG07sBF+RBtrT3iS7GZjVy6tX/GX9S0XyJ+sjYc1eeR0apL+K0FNAuG3PJJBxN
qVnr/H4QmKbVb5X0GzzqfRA0TBEfBzh0P2fwMTuZ6eQ8M8KMo4u33986ngEBOfDdYZPQ9wE2+0UT
PoRQS06uxF5AxniHdM0nTCAUhHq4oXSuexqDnbHlHE4xEWK2y1NAU2KsRu2GLhxPg8Ou+uNksnuX
7GDwKDgu3zppiSL1YegulVzvnxKZMolSjAptfu650tNyNumaLqlNC9LkBye4K64S8iDlVbdfzDOl
GlPxZTgpzTk4aPeUPxadxH7V1ZyMFnA2DHLHiXxue+laD9JSYE1tjuCenKDKkwKHsqfkCz27o+KV
kMPofLILMV/HxYlKKnq6rbChqx8WbIADSdfdUnzlGhHb0BR1zxTOQYQA5PwA/3nTAmi14C0LZAcG
p058UcLIYml5kv6v/hyb0jKEs+8ZlJK07mmgHbXM6U9+SSROhqA/f13gNlQLMrdf7jbVm5elAYj+
G4oAo+C19cM8p43TOv8BZn7LaB4ono9aWftuH5woWftBdP0zkWSFhCyUythAr9vo1lAzXE57WKdb
LbCeRpusPXYuMMgqfF6XMSBRAXd4qFUSF7ooFkcFixLL9whmB/XcCGE1rtXlVgOhanfDhEDyUbXu
Z9osvx1+L3orDe5Tp5pzrGZm4gzZ54duzyvai2y1pgrrKgjwoHbZ0Nc4/kRwNyjDuuv1irQ6Ug06
NTggyk0V3aDgEW7BS3/rFBNi6wa0//+BfGPjrfUhOfhcGHOxv/aIWiqsT7aJ3f0vB3DP+cK1V0fC
/ejxX2T/CWByYGVIfTnoTN+vaULGsopZaptCcpo4Y9+4z8Sj4ibXtfwuaceJHi2wHIRgtpS7uCbb
66b3PJZoEU8fgkU+OwNEfRH0kB81rHw+EOYqT9uWZ4eNwVDLL3UcrxLZYMYnb6STcvZ+/r1jwqn9
tny4UTC76xGUPlih+0kmOPAX7sAoyO6C6qXVtjgVZXcv+MQS9m7VT26KXe5oTnganiy1kJuTGB28
m2sMQlNF1bXW4BRW22/1I0PAHS3pF4P+WWypZFAClMxj81e8icsRJjNAxk9dcSP/uLbrqGX30NUs
1AuuNputWLeY9hoDCBS0YXSW0jN6ttWl7y3GrsXEm88TEUeLI/VCNVXb4BpsbeOzClEq4ZGXPuLc
TS6/H073bg4jZUB+ysqv0zdU0dRxvrI7xaI7cD0k+kjjEGgrqr0Cg38jReppIDAbzEzyjmEjU6Tq
haczwDNDnm2zMIOHWoVJjp6AENTX0tMFaArS2Mq/jnj2JYATC/huz8/J0VAXQh11euWjKIYoOZe7
8wLysy/yL0f9xmajwD7Rtn9c/S82JU0629rfzmN9IsuZAOZlJK1v1O8fbvjBq414gTSVs9PtLJNK
NhbULVF8PPnUWhaqy+yzPA+Mnz2c+xihRRRchfqgSr/BM6jPLGh8Qmq4GuoN0ZUUWRGugKxKW0Ea
wDN7NvSuGHW1AkC1epk8u3/OfYLLKaozZFprl7YjypGsGUULTsqvXe7E32LNxEldhpZjQi25sm7h
QlA0dTYq6TMa8Aa2bdybu+95na9cTTxzP6d6S2PWHi8o+di/bToU+3iar+ryapZdSy+hESSPA+L+
ng0enDl00VgxTBONQEJfXf0/uxHMjL4Jzg5EC/V2KNRqBb536XUnep+GcGMlNzzyTTluERS6ctlC
5EeH6rgthMdiB3sjjWVuNnT4HEjEF0yokD/AZGi3nGGawzUPvqtWAbGOLkyybE5tGJKDV2joS2k7
Gnc16mHWHjyFvigQr0WvVGbbsq+AgpsEQ9hjO5zEz0JGkOH6uC62ELVXsbNM8fZVNlOhRI87fEy0
kFUf2WgqFrJgYnSamlDuiFARgfh6St2WhMVEFBfkDRhZBj5KsDHt52glo2HtlvrX9b/Blhn05vxv
3XIsKIUAfuW2s9r7frzhw5I/6BTo+hfXjwOdGEc1yh+09zT1/LpXC726ZCku+N1TgjpU3HVWWFeG
F+p8W4+gjqpCwdleAtZRuVx3lCdgTjKqd2WV6qBwnDuB3UtW7KvIDaFI1rXNB9ECN6kLZFMR9YIT
ujgyArdFKxEw4m89QUCn7jjghwE/3fBVVHPI9p/SfJklfzRGCsjb+qhpRQsblNuOKxvsqcX+96gi
duPEQB7V/gfFVryEVuptDDnAbt6od0mixlNdwpajWzp4f/hZwE3vz7SAYTXz8SKWQ1RBT5LyXP95
dp2gMhg7nPcg9aaprvIExilewNWNy81dwlOhlmsojuUMLSHAcYi9ms8bUvHCWsY7hRcm3jjp1de+
FjO2otZCgQCX4rcZ/Bw/sShNHkwcr6rD6fe36cDomuyjxFLK0rYwpD2CHobSnQoCXnz0Fx9tdv0G
R6thNykZFGKsF7oJyWq9LFyo52jVJj0IH+0zfV1IPJDS816LRSkUOaQ3i/N+nPQwrKtDSJ2Br3kV
R+24cYS0O0RhDqhTX/1IebDiH7JLZV3n2kedKqkE/RdV7S/HmeIVnakMeeyFhHDRQHyz6thEu2W2
X8Ls+4KvX+tUttNyS87NXJuIqd8T7mRxsRUBZUVFA5CUQ9a8f9Lk5FEXXxbUWrfajLM7U1p8RAq3
Hsvh0DR+I1D2PzqR/K4Vkb0KG5xC7giJ07vCPNmJKvv4CYfplpb72r+bD1pg7KJ7mJPV6fcLevP9
OsMou5+NgPHJeGsfzRMc/mLPMbWyoOM2GKYJ1jM7uADrRXXxvfM75PUhndQ9FO5pX8OJgBZAKJyB
I+6VGD90H88vbmiLBQc+4TbWXHm8gSvp9VmGTLWU6g2a2et9ec/qCJQ4QMHqZBGfz8mIXig0ptBD
Yp9w12ceZAWvN59VkIHBjIYUNegQ6hR4q0pCwzpBjuBcv3Hc7DqJvcN2AGoOmg==
`protect end_protected
