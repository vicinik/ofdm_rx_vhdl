-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
jP14RRuobmgn+jdDOwhgPT+uHyRKFGmy6KEYd8h/990XhzvTQfm7qyDiO7uIa/K9JpljUF1QRBMy
TWsnZ2D8ArAxKX4HwmviSoO+29CkjtlsvTTaR2De4McQ0FKcGtz5ex/ss+rs/sWfuKBQWut3LNAn
+T/KxWOL2Lgjk3v53vcWMUaDofxHD1yJbdUN42dNrsz+Sj/dkcNqcBwbp3psZsKQ+RMH6G/yE8A2
9Jy2w7gHJf0Y845mnNa5iRdmke6N3hqx0pha4dRD8kKbct9lW3DmSlh2oYclUwkVnfIOMExL6i+S
LKdK2V5iuEgwp2MCL7xmB9x7wYtdRk4WhMGA+g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9728)
`protect data_block
v44wDpEDLwajvYB2/UKtfYQrRzEFJJuXX622VqbV0bg1ZfZSq0Cxh39TfQpWJXc+gtBQ+BwDUght
pCSRgpWJoDI7F0jbC4b/EgyGkcsuMLyd2TGGXH17s/YtdxMYcPkwOkJYaSYCv4ELGQ+wBPdzAIvx
14O//EENxhMIl94fVC9ViDoqDmxBrOkc46JwJ4R9kCnjB158u3E0IIGKtSPE3tQgfuZPnBut3haK
cu6KyyiH7Z8Nv3jB4dLTzJt9N2VZI2XUqrXL6XSIqFJgftokUPsizYhy+ABcZGcqFt8rCdPvlG27
JQxibHNPejTwE8wAXbNTic0ZWhfx+7j2R6UibI7IIWNzf2UbX2fLc8o7KiUXJXyY84MdyGOPqXP4
X+lCpD2Sk0qRVW8pVDbPmGSbWcDpoPjEfJGjdBJ2YPHgagSKJbyQz8VvYzIU+caKEmZShNGfSgg4
dD4nkETRyic8LJFoXT7FuvKdClFA4tPvKk0ugkx7hFFBf4Z+M3ajmy4PEkX6kZ2nf57RAUpdWqOt
Fvuadu/BYeoIImVB1Xki+el13+PXTRYfKdohjVG7axAVaVxTnWNzkVIDBLTdmufQps0FNI+FTRPY
kQva2zchHxQkq6Ke8OAwTzfWsaPScXn0S+7uSYaVK6Wy+0ARMODTh6PA0Z15YtkSs6N6TpcgXOO/
7BJG7UUyYqlsBy5HTC3fwABwn6Trt21XCgn74BKeSAsCuxo9pUOzlygd4km1wAcqwSRTOy54Lkwm
J89qLiO+oFQzgKODX1+7wmmjbIjK3qmSTi40Qubh/YpWTchO76kRQEPGYDZfeaYlXd21BOnJK/3T
EsfFJiGMPiZTmDgNQqvqJZnXQJtunUfAxOTcutnyQOKo/52G0BWDPPKdeKKXUVay4rowKKBqEvVz
ypvff6lbK7FFmvu4VAqqMtKe9CG+CiO/uvBZ7Dy9TQ8gPLEsbdbYZQHaijefz9UmwacvHNpBj7qe
0s515HnETbfGHy5agFyxWHlCXthlcdMS+bG0f3/9aWmhINmGv14FZKh5IkTFxoqE8mWVb+kwMUbN
Pk+a6G622RkRxVofKt3ERYubdbN+rpf9YOgyhJD32nXNJF6E7SYcPJYywOr04f1IzJ3NGrnseZXP
Nh+DHzoeHyrRp5Du71s3tuANxDuChbkXPREGDJaKGPRV8QDIDy/dv/0Lvw5FiZiBOaxRaWHBRvpQ
s6zVhUtusULKCCQjMtlm3gxeYqPzksQs/L7qz/C9ljbcNxGZuzO12vFoB0NxgwfusFY+qowgmSc1
klNKLbZW44xIPdhWZk2d8/V1CntXx9K2DELgl6Rs0lY8auPJUSD3dw/NF+oeKJFnZ4NZfHUvSu6K
B2YcyfFyR+2e7SRFPh8sdNDJ75GqeEk0yMN9EcE1geqxwY4jnBZIVbZJz2DcAw1MMSRtGE/tR9Vx
EF2ST/HBrhV61bpGjLRYidr+kgc9qUH76VS6GLoy9J8/0nAeDDQIMs7yFN62JNrag16BiZgR8e/N
vW5Huy3byUHZIKGSkJ12zT3b7PSCIBI0YD95D3CBg84NUYVTZ7QzPBDnlw3YEEwcZl/fZa2ud+OF
cVdmO8MOkQHwCOmYyE7AMmmCJo3nxr+97jeSL/NCVUza440fO8vzMJZLjLJdW57pw+sa0+ZGQQ74
JA6kOoanVbgm1uJQ0arqwd0ARitPcSqOx711aHWsuL9qB3Pk10/eQapU3YzKRJUJmrHIuFhZtv+Z
N/AedfZdKBy7qgOcO55GpI/k/XYplSehuai9vEXkR1XCjnfzCwCjl6/qriiemQJpMR4r5bTNVqbV
WTXfzDROXkeR7GfOJcOqSiXKJk9h2kgrFjSJKwu87mOQHx+uYUlpvProb+7EGrWqd11WRcZs60vF
GBNWBWMbuiykNQudSqcl7TToF2KEe+gqjrtllRRheOp5WG/bwMmS2xRjWkZ3EYeF8MMfv8XrKMGd
PpNI2q/xJjJ0r9cMcBbyFp9AuLqf2QKAFAXTOItMcPvR/P3t3NT3yanVIoskApnP5ocQKaW8U4cv
mvK299Q1W99lXTaO8m3RZX7p+mR+m7IhhxeOQ1QL3F/zEL3Q8f2GMcqk3M72mv5iy1XC2CXoP6IW
W/mLVLszbkWsLlAk3RN/6PdQzAc5NL6XaW5xqoRK/UzA+h0DMBZCsBrjOgU+oipOYRlzYcpCaSRt
kmX8OUwGlqmX/iecO8bQOCyPuREZDWsVG1jGfqgYNFjklTP2n/jNHCDdmqFU9vwdcFWQR/O791Pm
mH04d0zlWyt0nDeVl4FjH2RyqaRCI0D6DxISTwQJA0jam72yMjrxnBnVShDXvyx9aJRI+qZu/FuQ
2MxpxAPFlejikMg/ePlN0HuwzgH8LFnBn1ZN60lh/L3+F6cF9/dJyYPTuAn8iOjNGl/XTSx0pX7Q
9RluJoPeeiVcZQVMaIF8QFpb7i4ozrRhQmJJfPvZpn0B3LebVpoOhrh6pZMs2Athtolm8cEpC/s2
HSA6gipsR8zqWkgg2tLU1eqme05O6JCD9i/dBkcW9VTDRc24udwfzQBrpUVO2DmjUfTXn1I7bF5Z
CvSvy94u/jw8CL1Dw+VvbV3JFL/R1Dzrvb61lUvM11ftfbkHt9kitg0baNkMc/LjI50z+YFRCmTV
oh05pegBDqg+F2YU6vv1ZTLo/30Jg6g7/erJYsn9pkGUsp+OmpG4ZVoG65/IQCSspRbMuxXDZh/O
DIQ+bmOIbqv2KCLYg9cc0NQ8EqoTdUhyha/rtZOvFYTdeArVVTYPDEarlsqDn/exz5sXnOedwaJn
xodCe9s5eA4eMvRyzCAvlutVVHJ52PyMCkSyRBeIoNx1X17oDa6aZbNgPJmDSkWtDUjJE+GbYw4P
Fh7wi7gvUUMxCnRaBrO7kc1Ld1RembLZa2o5o/pkYF8iDx5/j2KfxFqlztzxXtrh0uOW/LXt5Zaf
AKOspWDjZuZ26XwIW8H/SG9hkQNSTg/lYMXRQZFdjC2uierZkhj1yTP636bjK63zSjs5QP2Mywpz
pzwDONchthA3tNJvaQsO9Xhg2ekukZyk1EebI2KlmvISAHEwG+IQ8sOJtk2QJygEQxfXHFGUBCvl
vzKMmvgkJgNUfzOX81yonra6keDLJdi9KVO2WXKaOIW1QrsqFRgy3tmF+TwCHG8cfnwiLfCKzcAt
xTgB1yHxVPU1QaHrRPl6DaG49ecJTXn2apGdoTIq+h3yKKUdZFNx0+/GeSKj4cCzjGIzmLF+eFJn
50PrXof4xCmDaDQKPsBd+4GpchelZcZAHSdAgPx5RzGAa4K7OUbGiXnnJQ0uPTSrVlzbCetcOF2u
APb0vToFE+BaZqyB2PqtG13atEnf2eapOj631Efj2hVL+xOgSXgzAt41oQtZQmkE7QF4HdS3lR3y
1NYp5sKLCBZu46cVanNw+geCi8YUrxfulKAZ1cDtKKGIe+JeugY1HviJ1UZJ2XiXO6MBXm3q0W2i
yNUiIoS9gBCcz2qR7t3VqFevDOIxeDhABxfkMD9OKVauwwe7x3118UnmyksQ8PdZ4giG9DrVTJ4S
UzKJoYUQoH/NDFwXAmYyYxjTd6qmV86LUJU7uKBYtPJk6TqQ32eh5iNfnWVIfEz+LlKcC8uXLh5c
Bw7tHPP4vVWnQF9dbCU0o9YGyx+gu+yLTq9IY6E9JN1SxrjcJ2+ARwJ71Znw8rLfflhIPH3SXhog
TpavPL0lVfbX/hwimcPFppQlDjy36NfCzTxd19Pnw13X8sWXB4j+btqkBG6q5NSCPBHvCF1xhBhB
gExHQvnGe5AO/i6xueqUDkMUeDPNbYwwoqvGb5+3lmy9eWNOCarRwQyss0R80tfSO+YdZRkn69jM
5XoAaOZGb/PZazyxAv5CiJP7Jw+D1+4gaAEZgS3RN9sLTyhEA9ZmRi++YGomlNCRB3r73uGwMLoQ
c3NaWojJG3PWUS6gYDoYKlWDvZcrhLsq976oNCyTDiXKIVMO9CKhOsCw+0dd0IRwKI70ZQJo2Hxn
YlnFHUw8uBGBjOC9qKvZggfmf7xVtDMffXlGwz97Yg3ChE76lPUR79Ul0HWDh5oJdyGCddCy5WQK
jH6MTj3qnkqlBOw+3d7qdcnqrFMB98kgX7De1qjOVnZieLP+h+PnR8OE+cSntUP4gcjGjVSuFeY5
J+etJqrOjTimm3Y+xppBS5lc2PZwUxyRMB3c8oID7NS2IxMBM0oUK4rAMn7hLZ0rDY/PKFlhVzqf
3l2U7mxrIfDbebh4I4dmfXvMmXqBhbbf4hGRXBOMNUVwAajo3hRlyZOcqnkCKTrio+23jRDV/14H
EU/kcLWC+sQ91ce4np/RFdQdCj71DU5//8DH+fdg7XDLAXQ+ZT4tXVZ4XQx1YSRgMrUt9FDqb07c
yLxuJmNa941p8xzUL6put2T3BUKX7rTwkA6JuY5azx9+PyPQokUF/J52o58qaEeAdEYxYX+UNIQZ
5m8poTCkhceOtoa11SpSj4ah3AcxJWMFHJPLClAIqYQe6bnFwXwzeOlCI06KonTfGf307Eagh54v
si7TawbSAmB2ONg856KyeZcYIirBrOG5qA5OeI90WM/thOVRd9g/c1c6vH8oxz+ILS/TSMguQNbo
3HAtKimZrHvMFX4oesdszElfuWdNo1RBYRxouX46XEIn0Z+9v5JnwS2Qd5+EoTnQA5oDdjmTj3EX
0x7K2dALyDaUOiv1jNru6S3arBR49ppVAspkFbya6DxHZOUDD7MOCc6NOurxvKSTJI5AOaVrQ1zU
DZMXHgQagfXlA0qpQdkHUiFwZZkqZ9CpQ+iGwbFKKuKxKN50wSiQxcD31vGAQn79npxWAWWvBeoc
g096X72iyAQpcONuLfvtJgnV4TMrjmVPzyvXL2VK0MKv5Hbian+J1Fxs46u4bhN8MCJxBpz6eMF+
PvjqdAucABd56xCyeP9BDjI24YH0xfLSQKZ2CFdVcoz3Rx4uWAAJo53Xk6YYRSflGE9+ZQIiMFOC
1BBq5hugZEfvOOsMP2zRCn/yNPbc3sKXk0J1uXVgC8WCW48F9CTDTPu/J9q3wMGVSFET+1Xzipw8
3Un1Lr8hP9X+taQR5kc6LNbdu3k/MfGGhYSVAPWIyObEWtfh2vPodRnzi3+mhzFj1Hv2TmY2burN
ArY9OKsxLXct1VGIBXlno99a251gxXDEqB0F4G+pW3htMM8HnUIcktE3dSB4gkQev7kiSUfh+KgF
Gcd/66JGzn0oY9vX9BNXFzOCljGqH4GPFIyNect7KAc8uA6+gynZRqiXVPO6hQdCiSo8ukBPD+1z
fWoAN7i/CxAcsmk18sfNbsM/z6+0qIova+sl1/l5ATQwhrNZau4/Nc0HWa0nSpSAzD1TVDzJjpQl
c9JlBb6/NeuYyLmE+6/AqlO9gRMbkAoETRu7I+w23NxBNAS5VY6UTpP5FaZGPtcwsY+SxQPYmMBL
ZGMsQqQoQpRuSSgfcQsVJ6cY16vhZuMeyEJRNgrNZnVfC8ISB3dd7C/+fqewhjt3PnDMcuzGN/D0
RdQz5dMnhXFoc+zd+m/jH3rhS22TPthfktiEuHGuSU6olHIEZbm7TT5pHmE9uj9wt6qOFZzh/KEZ
+5koiK03W0rTylMWDdIUlpIxl2f6eIVBKaj2eafI3ekMWDIs0oOmrzKwJQuZvHzkxDn8zqlQAQGV
p1yKJCKdK3pCZn6zWgj4/KfqUFRy6cC8Cbe9fbW1Wok0tnRzXOCLqq1h0ysN/sUzwbmCopRisEnI
fNgvhZskuRg+TUKHFz6StIGxNnaIgddA6LGzMFoSeENi2Gazd5jvJ1zdv3r8o3jYgDQ8eixPBe2K
JBvzzWh35eTNUAy9aJ5VvhoOTvUVvuiwVmFbjhP6K/NA/uOp9TYGvgTxJHqYCeLN3e5UkXqI4wD1
y6Dg9pRy/U6RCOv+jvBzYLBmV0qHLGA7TVlEoMFPILM41ld/KVqQJ3L77mhaNGNDokQ/lA/dtafc
O8mGjHLVkQwMXA0U+cAISDZs+1e5zlukqg9Dt2M4GvZfI40dSVQdXh62ImtDHgH/tIYG4Bnyv2tw
J/VQG66r93+2a5hGMTQHS/uwQjJ7QXYiJ0pq8uWovZQ3et5vqSxbpyIP+xfI9CBTFfewuv42Y7XB
bcAoKlx8MSFbwhLsAFrrXSPWHNw6jIzeOEkcj0Jml5VNkwEsl5ciC04TiY219lVDQc0kwTOcMXb1
gjQD/Ee6O+BK1LZ4F+mas6zVN5QTIzmH+pYfj4hEP5IESZoOUsbNVvwFZbY05KBypka6kemoelB+
Wkdg8yCUEhYXSlCaUGn5rkVbwib9oXnaRJ75iRVOOILJARZilQcnSMutcgLOelvfvjIGd2Po5xMK
Y9S7XpLDbVid687rhescZyngH1h0qFyJrsLvCd6u9hrjDpmkv6Gob8xMjpP7tT1cFhAUmNi4/l/I
r8dQ/T1nR9RuIcPp1lvcLGwOR3h9CwFR6qblbkr09fo90LMcRbl1W67VMn5JLtnPCmkMaHsmP42S
W7crmA/E71QX6pgVqVI74xmElbRfgiazoBra5uPzH7denRiefDuTMk1gWPLCcyv8FDdRrUNwvoe9
r1Klu0DtkBzjUDbq0C+5Ew+lJl+8z04nPpbwtHYvNgaGNTlf8ph3/JKKBMWO52Bi38ESkry2PybM
in3u1Gjx5PNByEWe3FuPdwtJHY7W7C7PmmrYSPaytNce5Mrz4KaFD22nFrMyVym27Bpx1FYJaaA3
Yo8QVb6BBRtAhL5z4YrpiXnxNBX6z5tjjTMK10bvjz/haPawIiJ7QpfD229O/14XXK2XRMZZACPs
iH8bg5gNJHIahHjGIdfEEjqy3xgJp+yvS9YqZmCOCY2yPMve7W49xhrziJghtml96pdKabIRsQOF
hKTXngil8/ZYRRWlInI30Aeq3AXLv2nULKFEiy8XcE9RYOBlkJWLdGKoHnIT3OvIr7V5LlHkrhN+
ZbQHE8EIGS4FQd8BU3Dhq5MGl400cMxj7tTPr2bMf91AO1/j/I2Y3TpzoXrKQ30eKkTIdewq37gv
JKpSZyg9zLrv4Ucl2fSzNJC6d6FvKtZguMT2mR4Vh8846fNc05pxsgfgG7DcEnugiFLOUcuwZti+
HSMSr2RVr4b9r8H9voc1kCLyHTMtOX1gnN3NbUIIlLfkflBR/1mjq67q5+lVS0T8FgSYL/wZ4Z/2
ur42EMi/wd9EPfzNnPKdIH5hI4YNh/kGwfqAbWOfxcMyGsAgaj7lVFv6OE0vNeT7LDRVmWAa9k4m
JufDjBY2cVThzV7ITvwofmYdXJN5HLVOneSCKXFLkZeC5zaYzBL85/zkD1/NhQV2Bk3phK/vfPOv
vMFNRYVPSNS466s6lMxBonjZbvgpZDmpRYvg02edRBNLG1RqbestoA3Q1i9xVbo7Ru/nw0q80JvS
h4w9WnPSbgorojgHEWS6lrqGp/vrQgIKGwNv0wsem0/7evS3SG+cx7BgT5oi/DhO4k2be8ndRvWm
ONJFZYYN7FGi+yxhhpwEblRfehZRKlQc74rVB6PJwdAf0DKmBlM3US/qUjD482TkKIwrOXFyWflT
bDhhRA4AOo8EUe7efLDpvC85S3DzBaPGNaK/inagUlx6gQkXUy3RxElyjVZoVKnUqJWZyP8xUFpD
2Le/+geDthoma5eUUJeUQx/DvlrVThNqVwdUzei0UbGtbVssAxZtWVIst01WnRAlScB0jaeCH6P7
iHDnP8MnNYMegDXbJSCrNqvzqH1T/8rtmPTBHGb7L1BHjZpeLCKZZha73a1aGdD1lxnghVMsKPf5
cGLXiYpEufij18VBS7MT3tY/Z5R9z3Lrn/Cbc9ffPQBizAi0pC09JKOmjy2XfWTzOk5Hbcwby1xi
HeQ2+3EA+2s430i34PXpXmJ/RlNIkchUhv7K0bCXy6vZWQpoqs6qCGI6FdnXjceleX+G0kw1qRvQ
Sonw/gyIvTV7a2L3/STaxKM7WgMhjN6MQDeEYTByw+YXfksha/iuxr59NsGR+tykSc2LvyOo7qgE
NxLdESgMaEPlzRvMu2XSzYrWV71dPaqwGmIVHF6wwF0CrOec2avAyYF0Zev3ch/Cy/j0+NRiF87W
1lyMTIkuaixdpic/FTh2BYaXZIzzVrNMtjpNOW8MbwHc92On56uenTYP3+k12dQGlfbxxf90lfMB
pzK4RsAu0WdC9Lw2aMi1unFOyRz24uU83daL3o3ub3tVN8NItNzaxzkhAaBTUuRq5YmvUtYMMlXO
aUMHKHVkdO7QuYzxDjFskeWfTHHkF35XMSwng5E5FEKgyPiHB7sksOcKH8837eirf/1zuMuYgMz+
2ESE5SnmIrqXZR/Hdojf87YCUIoURlYH+8qdhaNICY81v7+P8EGkQA1a52LQ2RT7kMOKDNiE9f7Z
PXd4lLTQflBKEJkIqi9T3VoZSXDxIiukTz6Q1paR8EZJW6kHoqGa3BfIXGEO4RXdPWRNLbt0gYkG
b5P7abuVd8fUAoEi8EcKboftxU/0pPpFrR8UM0pPRhHzut535gy3saLsLblgDkmU3i4/JUbQpup5
5o7lN6r4sdmAELLLqGw/Si7aQKUFN/T4eWrlHwPEbZNwMj3F+OPPXyL+HTUajMw3ReMeS9AftJuB
NUsqqQIbjLMji/QKHpVTOAn6O2ikFh5iUpQ1YEQQM0FsNxhJV312Bo/pnOOvDUyNWaibu2hvhDZc
G9hq8mZgMLEp4lFzbVQ9Scon/4jbS6usNzreKmY0WY5d+et5eHQebIys80V4g5TM6C9P+zdtyBFP
3gIxdS9FLBHgXODj3SEX8tph8Wlt6BLH1aPTtbRiBukJcGZjIXw/9k3E5bCSp3wQMO9PCgPe3mnJ
VRAsUGzk76P4Lt90mdzob175LlYEIcOUClFcJRgKuKIMPfP1NS1de6VXkbL5n4JZGRcwqz9HtVjz
4uT0eN4h6IsweiFhOs934qfxFHrURR11rdiDCNLRjqrrmcpYQo2KPGEkePqOufF48htllfM24yZK
QS53PySXr6qiG+TnhYbmj1YGrhRpnjb2tLe8jAJg2EKP3Y/+YI1BRSNYjQSByaMIKUAGGaEqsXtT
dZRe/8Q6kruRMPMp7v/vlIk87jMNNbpQaH4O7P2mj0w7GDo99N+KDv14JeafR9aPSdMJZUDgIl8S
h++x0EVLCrfKjYIU3kCzsTmKVEyeScsyKvtIdfLrdNN9WWyDa8F/wsjcH1PDxh/s4zXMkJiWH1m+
os2JIIyicXnR4Ckk22Gk6TPNCFM2HGr2jIG5Wbg/cz0ZFp45fywlJT0Syu22obSxROaU0QJLie6l
osMXpgjeYuWud5r0wAdlXnU4i5GIocj0JkAXuE6ZfyimcD9Y6m3JtJrKSN9CzWsTyisIWENmvE40
DxNtrnMJWCYDCvTdte2psaWzWL3inIV0QWhteGE4ME1mlVcCRdiEZCi3MjboyAWum8iqFALeL8yo
SLo1whqb1qpsRNSELzOZwP9j9rEeXX9vc9jdMQ9nHbDZJXdDgeGsBviSQ5OTMGarkEmD160vUh87
fxbLbVFMWD6fzRAI9k6aLshJC4m8GN9zIGaKnGspcLrTLIhQAa/hLPtavb+tcRqpKtbX8q5mwNa9
CC0jZmYYT9uxXTJejlOMuB68rlK/lwg0wCZMOM9ECA/S/H6JuIg88HdbiFClRD1fl9d1Pcnpn3Bb
3TtQd/ptvzJv6q87b77RPFEmEJ6G+S7aux0sQxTtIrJwbHwZmhvSDRj5UXvDBkDqZQJfQu1F9974
4ncUetdsHpVXCBMe9tysBlF1m6TzOAvg6cAkIGZnA6hpKUsORJY5xYSCVjXF/xMNnh6E3VwGnCBT
pvZDJ6WxzlJv5pGZgKd5IPVzmAxUh8XdWovVtoS7NIt2/tsDyzwmnfJR1EBBeVE11Ja5FDcDPyc5
nXq+LefishEoPb29DZgqgMd0YMVrTd1jmQlv8PsPDd2U+vEbAI6HLijccM+Iho+V6IzbRX/SjYHR
2uoeztX7B8CeErLXwZKexAH++FpQhY9VOLAw3yUVPzYei439iG8+2WfkuFLc+/+n6UqEn+F2hOuU
JNUMtOJ045PkKU2SBgRPP62iMAp2yEI3iPdrj+zaUhgCj6G+zjL9uEYTCXE2d+4XqI3peu1IK/Cb
1VqLN5pv3aJ6fXuXxLQ0ugrj1ZtdoMSyl3dTcdBtD157nXgYS8JvTTNhKiTzKA4NKmf4SQf0XghL
Rby8SNxm/ZfzwHxenrmiKQDjCexDSSkluMpuEG/eJoS94CHE7Mln8GYFAf1FXBiXYq/SI9fxEeEc
QnzWdriq2hZiKdiNMAteNJuWZiQoYDjhKkIAG04Utu5RZsL4X+Ae5gCBi1/JDRrzu5k2GZJxGFCm
PDSYOW3fxvtPIM8npQfPKhKpNgUwL3Lr/6gJ/SXG9ajeup9fcojt7Ua5b1HtlaJYlHO8e6QoB+2y
Vh0TVmPiIxcLCwLNAlNuwkf6es2su1+AwJ9YsMhPVUSgAj/JpPEbUaG6EqOtlYi0zF8TTL9KDCJz
GTMB3fTDcArneUuobr8HdPDtTajZkV0z4wPmd6d+d9mmJlCai0WKkDnmnfi4wtvpa70+pUoVHHDJ
SDBI9D/rqROkZZuzP1ksHQLolbb7YCwe4kOMCJ8PeQ1d7AF3VkEQPLWTYo33777+n/uo/+G6UIo5
ymbNb9ec2r3b8++CI03rM+IkDDl2D3H3bcs2BWWd2ZJ2EAKPSGJsQ/EMMCZpua0jIBn2WuB2N4Yw
Da4ASDTai1mU2CwEUdvKc1GSoFEt+P8zF+p0l2v28n8Fv9Wti3XAK6vjXR2hbpAv4CvSTEn7xjJp
7d8m9MGI2YccfWftbqyW96+n0AK5tR82zWowDUYedbucGxOMFbKkIE0DxGnYjVwDezHYR+iAl7Dh
0U+jb6rTE/VeNX4jH9bQs/X/Mtrun4in5TICIFLVayjxsn+cuN5CBsjM3DhU+MCknGVGFY6fyQNt
JFg6N4vkcMj0p/RzDxH9vjhVkR9LdtAlodPooAjoXYqJwmgApEh7D0MsWb5R3K8eqoHG1bVUum7x
/6au5ojYiXLzCY4/5/gT7ZNzi90cWjhI/zDF7GtdvSPffKYyBtCD5/ys8AZPwpuMs3r7poqSleIC
GTb6/JCuJSeFIAZ3MgYNc7vVWhuu0GWaStvX5zo25tEfV708SediSpKysFIIolERUFtYs3prwx1P
EBKb2i0U5xULlXh0VYKwMTnX5x+HIfscytJVdVDuHn47Lg8la5AsgQKmexLpTMaNsCuewWmbMRxh
Q92W7g2W5wV3kZi+J9mywpHG0PTxftS4NUHFocPKmsnXYUhomTws6OX3f6jk8Md0N0bUmhYQT4Qm
CS8dDGemWv7vJUNjQA/hJjBfmEgsm5T4xXwKV11ULGGpjHgJi0OuWkYmB1r7cr78mir5bMdFao/s
qdLGOz5VPOuR+PAhr1V/ytqqEYP1w4sI4XGnw3AZrHj5AuzdzdJum6vtAJSko6P5rVX+6KOshCOW
U+4VZp8COcD/krMtbfbqdQsHUIVIJ2kGgiU53ImPmiMQcho5fOQ25smw17kweFv9uL47m9COQAuF
5J8S0FAM102PT4gmoHnFhQle+1ErBEk3zHNUyNwGPS88U0T0uaY6Jnhms33AnP3Hh2rVPPEiputx
1HwFOUhtJB20Wza0wt6NgW/OJ3vQc1XidlPyQUgsLZea93KiflyzsetZQxQx44cBZsSzim2MFTPo
IGbme/Pgv76pAX7EJZQnTgQAm8civVua+CknlLujnqtGV1lUCfj9eNR2nRqessjwn6XanY3xzyoO
8MJ2NFBBARNCD3R52W6cISM71D1DMy95ndp3hEhicLXCHagLte90bL8whKQt2zp6jEuy7vZsTd/h
9BO9kyLi+U55PonfLh9QQ4trRQmy6VSNeY/GoT3oYlnBu96Wf1Oz+JQM89WaE3tQBfBjhIt6RWus
Ds6wwIBaMw07+vDNMg9TNOzjle8bCvNgahANX9K4raQ3gsyn/WPVUqkdmkQXpEaMn4lBIaHEvlcQ
jpdRPrKgCkEHSjnEkyQ5JgoGaEYc/lu9xd9FcyURcCLFVsjwMBkDt2oiI7p4brvwH3YKvRgi9HCO
7tRB2AM9LTqfceq/a7RJtlBecuEGZFvtu233sOvZuoYO8+e4+jThi5A3/jrei4B3wo3nCywfk91w
aopm9ZimJ26xH9UrTBOvsQa08sOJPcAWUnmKGStiR5ANOQBtC4frrj41l+7eaafGlQfZo4Lrvist
0Oe3kYZYKqYmABSGN5s/Y8X/8di+a8LsjAu+oGpLWJdLJIS+/C059cnTflCFDxs5ttCYR7AfU/Pz
rvxw0m4NN3O9VfftMZnEylBHaFmn+pNNkTBTUnk7W1IVCO1h89LooAWlZXHZ+qceJicsu1xxrQh8
u3A33yYVxG5gINFmEiJDpRX9+d1lu+ryHzZB4kziJdvnoIF1te+rKy4VO6WVSxvfo3+8xsY7Vd16
G/YovP9YGTnQ+AHwHqHoCwtNf9PZetIBT7NVe0tqKK3cNrzyiVAvv7ecOiVL1nDtBBBqokvtBo3T
YItHEOtq1/uA0mNxH7L57TJ6voSzLEepDRf6FXbMZHTjgW0QaDS3T5SxX2lM3N9QcWYY+qJt7p/O
FoRGZWQoEHI/rCKK8iZ7a1Gim1tB1ZmyoDb1aOaeJzlO4jJrbOBr+YDn6OzFC+YnbjJMKpRggkmp
t8TXojsHeAkegl7cK3Esi7JLd4LoLizI0kj26IMNydYffmCXX97PvbASEuYSXNQUf5HOCTnoEiR/
zdGSgWfIKzo6W8SsTNml/VWEcAjRlIxeLxHctew51Sdau6lMUwuHh+OtZEv0NXSpcaLetLCZcrEb
/5J/eoZnSOPfRMPYy1WwtudgPq2oeV+YQ+KsETnnkDXQFpl73MM=
`protect end_protected
