��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��8&�����c���a��8���@٩9�����,n*��Ӌѽu� G��cJb��Xu�����n�8�m�.��.<�t�A$N��J!���D.I���sF�BY�(�����fq-l���P�ٔmB=H���3B��	��o;5,�w��A';�z���^�xv�����7j�;"y���Q�8~��p@N7�˓4���9c�m�E�K��B�̨IN�z/W*�=�:K�U�[�.1�3w�>�z//�� R%����0:�� e�������0�]ĩeKB�mI�у�<!y˜.?�����h��e��zI�`�7]7`ʉ�P�l&IžA
a�t(�j��WΊ���?��T�%C2��@|�e	��,���)��^�!؄��-��PK�g��jl���<cF�_#���8)�4������ ו�Α���aLɔ	Q�SY���$_,��/'���dѥ ����A�ႃݝ���O�?��Ǿx`Q5��G���&�Y�\�S���-,��n�Y���G¹�ҰNuCO�?�.q��x֊}*��F5�q�Kf[�tO�e��y����KX����z"�6�C|k�>sT�H]=g�!5}rY�i��/v��X�$���;7��)��nP���r_��p�fэ.�������m�h1mrx�P��ȩ��3#?���ҭ�� 3S�7hM\��������\�������o��"[�_�eSO�l��T*'ʚ	ԄCI��	��S.?pcF�p>�]@��i`�C˟*ѨkR�z��������� ���e�ݽh�O�KBi�����;�!�����sc��u�K,�`�!{o�׮�ĮGB���H��HÑ��I��k}��H��UU��n��Ķ���ɸ��F����9�AdC�(�����A����e&��&c�ҳ��HG��vK�W1�h%�g��&��5��x�Uw8���$U����Wn����]����}�QN�qv?����u�/]R�R��j��%G���۝��H�W�SX_j����R{����t��%�{{2!����4�ؽΫ�x���|��j�Dp̟�˱��8����[�ϲzA�?�����\�����V����z��m�XC���g�
oU�)��T)�N�j�j�G��#�@����<h^��-
�$��χ�CZ�+WO��	���Y�pI.��	����ғ�%�����b İ ���US�� �dV�DD���]�;4�\�8	-i���w6�'��ن�b�@-�և�r�����,����csG�
y(���q�:-���.���Kz%j���r3>p�J٨��\�Y7� ����!d��
�����@w[J�M�:Q� �^�x/*��}���|O�ᾜ|���%O&�U����p�0���5;�$�/&�{�#����H�������8l& 2>�Tl�3&"���{#�S` '���$����4���~_(�e�l^� 2�&]{I��U�nqQ�5ȷ�E{�Q��zP�Y.ї�/�����1�h�'��������t�O�1p��٩�	x$���/)*m~��=:�3(!�I�O@�E� �6"��c+ɂ)�tf��T/�����5ʧzɐ424��������QNU5�l�a�U-�5�R�� )��2D��;��	O�z���-���&9�����u��!�-���d0㼜 �T{H�P@��揉kC��,5/�}����#%M񰢢��+2��
j
�N��H3AP�hp4�*�T�嚝��zk3��	&��ה�q̸L��d��`Z�o��(1��GÓ��qA'u>,���dP Kc�Dm����9 +����D���`�8:��{)BC��	^�2܋T�+�{���7���?u;��K�6��\��̻l׌%]꟰a��HY3�*v�:�?�.*���[�-D�sD+9�Y��oP�T�=+�Ws�˅Bs���"�/�8�z��$����p/BCr��ٜ�4�BC��S����#[׺���x����^6����薃�y$�;	ؚt�ob�z��{v80<��"�\�,��]�K(�>Қ���|��'���q{����5��\E	^�t@!P)	^/�<1��ݖ�&\�-�v�7u���;�1�j�_�0��	�� 10�ͽ L)ﴩ��kٟ�(h?��@����vR��Fh��r�&�Î�އ�E��Ŕ&:�9�=$����.�`]L����8���A�$�6W��i�Fè�x�@��=�T;�����D��=�Q�s�I�l�
�!���b'�F5�Qٌ�Hh���C\��64Oq��ڈB��̎[�&:��U6��#�-t��m������=F��ySד(l�C�@D2�W�9l��l�}fǾ4�L^���>p�����
3H�Ug�a}#��{F`�+�
jEFc�b�����g�Q8vj�"P���L�_'Ƙ�՘(Z����t���]����/��M-��V��F��vb��	h+#Ɉ��|.}\��.��̀��y)��͊Y���aK���^��nG62/�W|�����;�SJ)�+�����T���uVS���6_���F#
[�}�S�e�Z��T�E���w�_�U؍�����38�q�b�X<�a�]Y�kY�F� ���Չ����Y�ء������A�<����W8��3��g����#�+����׭��22���#�d�E�t/�KF;��ӧK���+�}��#/ך�T�';��'"�d������Lh���P4-&��vW�������;�@ u~�� o��oA��M8/�4_(,�"g�b ��3�."��E�=���it�d�8�P`Z�n�R@����'�>,h�~#}B.����1��L��©���p�����4k���RRq��V.|�����)���ʫi�@��fX����S�E��'H^�q��X:-�97�O"�c�	x/r�z�ԩ>��l��LHƝ���.Ȯ=�܌�:^x��P%���'���=��x���-T����m���#���5�I*s�5���]h���4o��tػ^�C�8�F�-�̱Y$�ު�W꺬�l�����xJk��t��+%��'�8%���8������r�ٽeK���P��3;d��I���<�P&^�1)��Xe�}$��10����MEY8t�&e
'�V�o����>��w㹇ȅU�h�b��>>Ѡ��Sg��ϒzȼX;��y����NI�5��Ep��| �!�%��'Q1�2*w1�I�� wߴ��c�P�\�)2��/ �;G��s9�m�LJĉ=�k�?��)�� f�|�	̓�D:�no@X�)�zPl5j�nv�w��*���#��f�����ؑƥL��ckTJ�ՙx�CRۏĴ�8����gX�E�=(HU��� ����*�V�����V��9qq�]Vo���P|��O"
���@�� /�!݈߷`����޾k��!jX�|�����8��p�mw~�@����B�!{����z;�{>%�#b��%+K+�7'Q�&;f�a���!$B��Պ�;�sry�	�́��D79�󢮽������֋�T�T�h=�r7�ʂ�񞤪{on�v<��v�0f��^~�p�P�cP���./�[S,!��XH�B���c}p�t��E�����h�Z�^a#�+�G{%�����B���I�r5�s�� 0�J ���	�3�&���*��p{��=�j�oؼ������c<�<��_|�	���6�X�m�F�`ɷ�{���"�s\�/^�Y�$���ە&�8{��r6���^l6�T���ȯ��6���Ȃڕ�{��:B�:�.��ZI����R�E�*)�{�!Q��h���"Dq�քf,!0h��L����6�Oه$�m�����p*�u��ў��\�j�k+�$�9D�
���'u���R��Oɫ\�����<��p��R����ze��a+��?I�K��f��PxUq���������e�� �1���nVg]!��|:]�!�0�u�gX�Q �^͎4�,�̓!�� ���}�l���ɼ�J���nU��P��ec`q���yGa����[�����?j	���!3���4�X)���f1��k������jd�z&*�SmKY�X�f�/��N9�oP��y��F�,8�#��고7]��F��Fe���#c����w~�Ԝ9�}�{QL��zln�+�I����WI�+9{��
k���-�d������$��(,(͐.��#���B\�ע�V,-?�#xe��<��!+�p��}G��ǒ�n�.�Jj+gk@�V���"��	�Y�%)�K,�~���M���ִo�SfT����N�4>`�#�ԐǄ�u�ĈI��&��KP����օ�9��O��؎���ξS���}3���B��j%W���I����i4��!�K����@s��7�E��:��}y'�i��xa�B�����(?E���X���8+�uW�N��=��j�l#.ij��"��a��I=���w�S1m~�X9B4�	dW�G3��ce5v-�A
;x |
�Oұ�a��ݿL�S���QN�wG ٺ��<�[=1l�h�����~#(���V4Z8/2J���^��f� ���	����Ǜ��>���Z_�Q�=	����YX�n�:��������
lJ�RVdr]a�B$Z�x�m� �%皉�7)�Y�2se�	'/ψIbP��c��_���i;�iZ�o���)\m{,J��OǦ����/ ����| � K�Й���?`��'p�r�+Ք�a"��y'�as�2-qҫ{��/��E��.�lP�ⶳ�YH�#Οp�!G$9�_���m��A�g'��>=�\:�hYR2��	#-�����G~�k����4Rޟ����w_mס���1`�Oκ������3�σT�UA8d�I(k_2�h��0C�as��s�򹜁����2:s�� $�ܾ��z5����:a�*���;�yca
{�޴Կ�2�qF���>����!���A�����un��iV�Ѳ�Ϙ�-ܺ��3��R�S1?�jyv1�T=]='��yW���EE�f]w�j�[��/,���G��lu��`��0٠���*����)�W�@�3�^�In�Ը���sF2s�!ҋQ �h��M�o!|� ��{7�]wc�1�'����0�#��S+0՗Q��R��j\>���̯�G6(V�g�����`13q8U���m���"��c�s�����?��хux�#�aM�p�7��p�{����CG��ɿ�NY��&0wk���[sO�� m��v+aʦ�B��k��dd��Y,> �|� ���Y ������	��CАi�{�s�g�J��<bB7;~\�6�����KEg,
ˏV�*��A�^`H�It��Gҷ ��u����߀W�T�x/��qS�ִ�~���Ѵ��Ӏ�!C������k�����'F�v��˽An�e���9���X���QH�m�ٹ1}gk�!4�ș���]ڋg%{��l�������<��*>�e'4�~q
���V)	'0Ͼ0O/#����sm�x����N�<@I��>�ɭx��t�J}ZM����Ŋ��W 4{d��.V
��m�~ԁk��\ʼ���K��_�5������g.�ψѠv����dҦ-O��g� ��|ᨊ|�1��,Hd�]W;�+��-���ԭC�~�.6Xt'�ѧ��j�#��64�Ѯ��.+2]��K��j��'����1^�J~�婋bth����(��?��$5��o��l����&{�/�<L�6r����ڧΙI��/�o矩\n� [�c?���{��5���ԇ=N����ޑx�J��{n�	������)aO�^	�d�JCiZ�2|��
n��ǄZ�ŷ�����e���i{����/�k��@u�h��'x_�ǭ��D@����aڜ������5��cM�0�cβ�~)�*����M��ON?�����of�ђ�81��1|I7�=b�]|˴���U��N��([ц��j ��z<�tn��P=r-~�<m�̐ST��u��$�JƂ
 �G��Qyj����>.�<��ۡ镄��z=m$��0���4'�94�\��ri&%�Q�?-�̥ڠ�Z�C�^�dg}������ �_�G�	���eD0K'�lU�z�G1�y[�[�6l'���k�V�1�JH������� ��\W�����i�Q�lwCi���)[��}�4Z���۹��H��Zb^�=&���\�j�ቼ 쁦KQ������sj��bJ�\T�����1��V/�m��5"ڽ$8�Z�o��GmMBk����Q٭�s2�\�5v �r?��V�@�D�⍇�C�]bR�41f�K�T��u#
鿙-� �R!QW�M8��ԙwƣ7���Aޣ�j�Y�ZIɻ�.q���U��9q.Q��hʥa,N7j�3Z����[��� ݪV$N���i1�����=� �+|��J�n���H'���	yE��)P��,_ ��Cv�]�)����(�����Cc�H,8oj���fvgfD��+R����h����G�X�o�i�x<[M�����,KvX�X9��~)���ח��f=�-��"A{����=�z�������H;���ƸYO]�9�O�F�X?���Zh�<yW���~(�?r��\���h�!s:�����*\"�,��mQ?�����%LO�ǖ8�-q����tnnwr�$����W����E=�K�b��z�85�:�졇8'@�s �κ ����L�ȧ^�����m��g�V$0v��&��݃XZD�Ɋr���/��tV{�4g �w�	A��D��!	�Bb�d#^f�J���zl &��Rv���c��\��/��w��+$m�RT抈�y8]I�u���(�������l�8Z
���N/\}��`��e��B˛7�/�7�c�O+���m?++d�ނ���cD4L��K����Q��������p�(�O��.LO���LxY��zn��e�U�l�#��0E�e��q7>h��4�bΑ??݂Ʀ�Uhp��C��ݗ��
#�����kq���앴ف�T
2k��*"-XWDl�����Ý��fz��LCڤ���`�BL���+�������C�S-R����/�xZ�%���y7�k�Ѹ
Nb%�NW��]�oITZ��N�X�;��I:�x}'D�Ѹ�N�	#���6�5�Bh����^?m�z��>Ǒs��%�p�����}?����l9�qJ�f�6���0Tt�ɏ�x͜Ԥz`�>w����a��$��/�������N���DP��H�������;V�E�����SD��)�S7�w�'9>"&�2�@���7��o$ g����CI��o�By��Et���� I�R$�~d!��A4�ܺ�>&��ۖQ/���ie�4�k�ц��x�2͘&>�A�95�9�[��dA!��F�K'bC2$yhb��}��C�'k�M��3~O4�;U+k�7DlQu�[f�C����'��T象
am��|gw�-s[0�أ����ho8W��9�౽b�i����9bS-���?+� �~_$����h 9et3� 흌xHY�����Ⱥ���+)���댫s(��,m�QBf}��#�LΈG*��N�T�oj�-�e���&�;�<�ga���?�-��]��'�]�����hX�w��,f����`��G%�>�cB,�nwo��9k�����+�K�\���ь�r��)�.%^4@N���^��6��6O8{�����1o�a��J|ƼyR�'���>Y�/>͠�p�a��f��gݳ�E�d��%{�V��i��+b0��F?��3Udr}�G�H&�&Xn2֜��N���ڨ��}Vx�#���������z-Ξ�R�p���`�Y��q%�~N��ϳ�'%�!���NO�t:@��<�����
E�&����D\U�F~�/��r'�-��K+	���&��������Ԭԋ$N�{Q��Wi�vpA>$��r*o��3?�hX'/�
��Uɻ��[<!��99Qy��������L����<���<��X`f��:o��
N4C1�"bq��Ā�˃?;0rG�	�xi�7�x��ۂO4곞�C�v�ុ��S��Q!�����?KX>]�齩ó<n\lϓd����\��u�!%f0!���� d���=��*͓?Zt�(�;T���(<����b.şĈ��㪻����~�~�C)�|�|7�{��d4�9�����λ�ī҉��,�1ނ� �!)�$K���혧B�$�c�S�+�xuL���X2�Eb��
��pגe�j?�!�]�6��aP���4�p���	�����s7�$�k�fp��_$�ߏVU��A���F9�g��>��؃�6�}�!��J�7Z�7�>t6ߗ~)h@�pB�r�!�||��h������������*�F���[S2p��|��_Pa�� �j��ɜo]}��<��i�_R˜C��,�c�V����3L͚̱l6{�f>p�,-)?���Q��P���i���
e?��%�tVr��n0����(�q�̖���qMzs��홌��%�oe3�?�2w*�$2`��,�r�5�`ծ<�l�44����[m��v��W{t�6��PJ����z��ͤ�D��*jWE�mF���3��<�������)%�F#x=$������?�	��� آO����m���`5�)�&M-�� ni7̞�t��.dy����?'aQ��/�V�'����e�������i�PZ(u�T]&�p�3��9���O|����b�p�X��}[,�0�ڲ:�����[_�����D�>����bi|8�״~�^`�x�)���6k6x�RR�4�?�4�����tv��������@j)ʰ11L����{�h��g��{���q�WH�{��Z�7��I3}�;'�쉨WgWP�P�_v/�`Ϗ�]yE�t��JrO�p�RS��{y�O���ig�*��G`|���i�U��Ѹ��d3,1pJmQ`�͈����2�%==~�a!	F?��}I��rc���(���H��Z]�&�1'U<*�y�eGW�PI?P�m�a}C��]#�?Ƥ�}�vc&G6�S2�#��
:�ƪZg#���Ŵ����bC�0�t>�J��1�r�L���/��9f�|�B{d��[��u�^3�����)���ܾ�q�N'�Kƚ��� ��F@obi���ҷ��:�諾c���`NW��YOHk���X.�o�<�|�
3�8I���y0�Lh��s�+:��m�5W)"������][���]H$R�1��FDa�v� ��7<)Sb�[6����rEs,�{qI�Yb�t�9��08�D��BW�!���Ъ]�f���ԗ��h�r
�G���RGZIr
"�Q&ߌ?u��N��Qڊ����W�q��w}��uѴx˞���LJf�u��6����������o��+�4��I��>��DၘȲ�|���Ч�r gpYڥ�m���r'j���L	;c!O�1�H0�i���>I�C������SA�!�b�s��׽)� �dÒ�����
&�+N�<��6t7x��;$��G��Nl7tR���n9%��O��1���UBD4� �����e�&�1��3���0kϴ��#�-���-LE˝gXJ��b���D���{
���<8;n
�h��+~4��_*e��b���t����wk���������������^7�|�d����)�M����G����ˍ��$/�HB�D�4��޹��m?!����A:��j�QV��.�]�&ש�8��b�Y>��ul��#xs�"	�O�a���c�ڳ@�@���
�^I�w�b)w��==���|�������	�)#)��Y��ќ��ܨ-(����y�&lKz�U�D��j��ׂ����$�0N�z)R5�JVN�gR�z��i=����jPc��Z+"�?��P��WI���e�/���-�{�/���"�Ց�<��wI����Ѕ�nu��t9"
��i&��{�5���-'���Bp�Gʡ`��;Q7-�h(ós��*����t����O�p�K�'�ql��ԦW@-0�f(�R��� �槰u3u��4�cl�b�#L%1�SL�Gi�D;�m�H�,����,^I����#��F��M��zga�	�)S�~�1E��[�M$_J�(K��k�~zt�9H�������������ɍΡG��͐���b�/���r�m���Oi�@K�����ب��q��� �����,����2��q�d��>M�2Wq>k�@DkX��v���0ܼCW�Wc��+8r��e\�I�;�ܝ��Ms$�yK�7�rmд���,8�V'ې\��Y��;&��D"���g1;�M�o�k��{:��Q����2&�+��Hb�P�h ��:�$m�w��_r�ﴇ)����oɫ�[M�S�<����Gw�h(ə,*�D����?�/��bu�	�[]�P�}B�W�H��$���6Bh��< c��+l�Ljz���`��
�=�`G���Z��!9ͦ�x�lSC3,5�[��*$F�C�) 7���<0�^|U� V��ynR�O�?��Bz%���Zj��F�_[�b�o�^UZ	�Ż[���f�1{�׋��7<���=dJ��ݴ���P[8,Ty�튝Z<ͼ��y̔w����~��or��x�Sn��;�Ow�g�����h�� P:�����"C#��(�(� A�L��co)*�PK�ߒ�N%�z�I������m"W�e�1���1���MH��iegw��!�Sw)w_Ͱ#aOS�d�^�T��w���=�����&Y
�H+�Ǐ��O�d��bc!��L�3m߭yy_�\v݉�Z^��5�{|�{����lHe��e�T�\G��9���@���9��.���C���M�/�Ȳz�]���b�`��n$�T�3@Tf=t�R�xY1Jg��z-d���?�V*$����N�@%�_v���r��S�����xw��<�h#�UfP� �����㺶�xv���:`p:���5��V�I�a�t#��������< ��ਚ~Q<y�����	�*�0��Z�/�J[��O����?�(�Qv���7����^i�|1o�%uJjb�S��y�̲zE��5��C�(���Ӳ�a;(�>���)�M�@��gf<M]�MY�ҌQ�Ҿe���߷h%8�ZY��ǿ0�d�������OR�$4��7[Ɖ[��m��\'y�����`'�T "X -C�}?Y	G����<wuH���D҂�<�I���b'π�F��2�s�7o�z��a8�`�;9�ʻ���/~{�H?���JcZD<��O2^/P�V�����=ʽb���W�D]���2�I|�ZKoR[��n×��ٮ���y���,hhR�:ɉ��e�.�t<���$�~�)��m��P7'gP~k�;Q�Z5�
/6�n1ٶ��3�t�v�mR�O�+u��u-O�e��K�Z8<4/�qw#1S��h�k=���t|ِn���A.Nd�q3�u��%���w�{�u�>����!���^<z��}_�|�*#T�QzX�J���������֡�=w@�9P��/f^������N�EQ���`���@������ }��I:bR��э$9�/3�=8pĥl����4z�VZ4KKA}D���p�&��Ȣ��ny�MC̜`?U�f���7����#\�e�GmMR��@�X0wI���{�� }���JOb
�t�]�g���*�J���*�{��W�U�r<ŵ�U���
�&ia��jO~�Vu΋���2��R�/���o_&�lDɂ]�a�x�y�_� ��(�࢛��C��_GU]�r�^U8=��h\��zN�\�LPpm���Aw"d�ɰ���/�V�Z���%lo���?A�}�0H0�"�-�}w���(s��.��J��H���2W\h��eO�pע���ˢ�+u�B*�j����I�1�^!V�%1��iEM�J����3Gp�Qd;�ސxd�9:�5Ǥe�ɢ�,ͺ��r*�d"�C����H$�k��i�G�TnH��+,�lh��M�3F�/"��&/�]�u��'��)�\̎=�)YxS�����:���1I��:J�������w2K�CN� ��n�]����a#�AFM��*!c������1t*����t4�)9-�vQYJbz�+���=2w�v&ŧ>����N�����^�Eo��1�^P�wpG����%�1VS߄h�I���v���{+��mG2'{���7U�𲨫@����Ϗu��6���8�Ðu�%q8�4����Ùi){e�@>��y�u���P�ޱQ�	-���o$op��ABk����������f��,'`W
vմ�|ګ����q{�q�ii֛#�'�m���`i�V����n	��ʥ
o�Y���R3>��4�R�P6�ep˪���"��|^�h���֋?e��D����Jƴ<�H��)�k�ǚ�8l��O�椖.���Q���a���K�M�`���$�n�U�(��,�qA$ܺj�������n� �i�QL;��\��Ù�;<�r�0a"��yx}a�JS�]>5�	H�:X��j}���8�+�������W�,����d^�Q�Zg�dqX�z�g`�0d�G� '�����!y�mn~�k�[����AC���C��.3��m��`���~���kh�>�	�4ǧ!���ig�_(�@��8���jч���Ke�,��3Q8m���k�|�u$��6��A�6���� Wd|�:��ei��������f3W씔��
گLD�R)e���L˳��(k"@rr�[_���,|F�2c�P���uv�*6��Y+�b��$b�L�����՝q�U�_b�٧���Ѣ�Ȇ^�xx� �#�:mP��	��<��4�eC����*2��&����ΰZ|�i2�ж�z�*L��� /g�w��O�Ȝ�����N�~ڰ>ב���$�M�3j�vPl;]�Ƒ�<w&?Oأ�_���S�x�+ �ƱiL챐�\@案�K���z#�h�Odd?��1�)r�U_n�+83̞�
�.��N�bT ���C�Rm�]6&���$mR6�..d�B��:^�����1@�W��_�ZX�Ap��ޚ�c��_e�� �i]�i�mOj=���.vL���)���qh�Z�ִ�*���F삜A����i*'��CE���Zh�xĉQU�+`�_�)�
��0���-'�ڵg'\��)Q+�H�#��ڗ����f�G�ߚ�(n����Z��zi�JrDҳK4ϖm�ņ��JU����!O���/`.�o��5��1f��1���Y�_"a���=����Ap<�&7R�=q�:K'���v���01:LM8�a��L� ��ϩ/4���9z���_����S�M�����n3r��o8.�n����v�I&�Ơc���,�n�ȏBE#�bx��_Yʍ��]���� y���Dt��q��Mԣ��XuZ�-{��i�[�[����֠����7�)��#e7g^�����=ܰ���vz(�ޅI\6�������Cذ�뽱O���ΖU��r�qk��x{ڍToW:�+X���i�@��@���c�_M��9P�����o���,�GW)���/��̘�Fz�|�<�ΥK��sɅ��lv�2ꇗ����n��Q���Â�1 �, ��ҹ�f�B��mI���;�>���?�T��=PP-���S�c�H� �m�%�"���x`��z�� ��}�Q���ʟ�
����h����^� =�\�]r[�4-��7���/藨���^�ŏl���h<[;�n�
�ӑe��M���r
9�0Z���&���%�������|�9<�{��o�gBq��6�hu�&�E jTN��G��z<���;��#	�j%mN���]��i읽�W�W�@�k<^�6���za��`�k�>KG�7Н�H�:�o�$�R��� ���QY��:�*o�s)�k�e�pjjut!c#{-�;ݓ��}V��ezl��x�&��@I�����9˂�A�=t�R*�p!�
����b�C�����R᥹��%�|I�'�^Go��:\~��*������4]��R�Aj�V��h���������d�.�I9���R��f�����������|;����2Cf	z�c,X��O�ў'���_�̋Y�`�A8s{��x_%�}��U�.BA~�JGԣ�g�"���	-1�M���enkw�f^%�~)�� �;��v]0&�Z���E�ZĶ2)�g"�bgZ�b����Z���ܕQ��;�Q@��)@����:N��S���Bz���_�*�b�������R�c��Ñl6�6#;�d��r��H���3����j�|�NdIu2,`�[�3ч�:�ɬ�.T���c�r��R�l4S� z��A!-�
�;� t z�1�Ԑ7d�a�	����h�v�yi���i��haK�!�HLN(���t֪�౤�fQOM�~OsL��;��MKr��rA������s���$�>{
���\c�3�_�=�;ۓ�C�����eP��?[��k���$ڢZ�􉣝jj����׬P�wj��:�B�O%(W���C_z�wP��U��+���g�� 5��*M�z���ص����z㢵V"w35��A L�n��;�<CzY��F�z��8Ź��i�������q���|��� �u��ܯcr�<���, ��N��>��IE���#���`��/�f���sq�҈uvi��D{���f5��#e�`$\���SI���r�ib����	q�%!��>2�H��������d��!!�Ҟ�!N�/�!Vx�m?����t��.�4 ����'vM%�m�Z͂�V�d�������nצw�.���4�qg���Y�j��j�R�K
v��Z�1��y��/%揓7�h���3s41c�� �9��S.TO��ynf�B����X�3I�-/��l�v�Cd�B�Oý����`/�M�~���#���۱h"���XI��9�1��5C���O牧��VN�,�A<��AZ7� �Ρ	oP�V׫@��/oi>�R��i�sv��N�n�����!M�t�O�;����!y��!�b�ʹ3�U{O%�r~z`�XTV_E^E��
1�`�S�l0I�F�?^�ֹ�k;Q.���$H��{3c�e����L�wg��{T������#�;��LT8���kz�VXKV��=S��7����enq��V��O�W��Z;����:A�� ��f#�d��@�C��w%�{!��Ae\TI]Â��uq��Lm�{���^�>��.�����w�>D�DM/}�q���N���Z�<g4�U��C/D ���cN����J��b
�&�wZ3��+�8�8�#h�pX�$w�@Ư�Ꮋ���</��$0�N�7D��ɸ3|g9Y���e��[#(��[tb�=_��^���p��$B��7(I���з|܃�[�-��(����N���)b|�~C�B'�p}���!�a�2!�ɦi�e7_�F�z<���2��E3d҈|��2��.�y�oK>[�J�63)��G<_K�K�R�Ad��1;贁8N���+�p�[�L�A@(�:�����,�ȵq{�6`��)Kf���#�ք���(��I���q(��2��6�Z~�s��y��d5���v ����o=9��6�:��Y��%�XH+���r��BˡA��0
J4Xׅ���C�1����l_	B�0�rB<R�v���q҇xj1Ì�$���(�3�,�:�����+�ڕ8�q�03�S����JUrލ���׈���bd3�W�KdV�����g�d@_� ���,R��H�V�ggߝMx��<�CKm���d�V��ȂDY��pp�J�<	�Z*N�����84���I������I���WBγ�3S�<_���5�1��3m���︷a�#�	���>����ku14Q�8*�m���8�YM���L���1�ꐤ���φ� ��5��	�Յ�aM�R�w����DCO�`�ɋ���b��P�҅�j�
�9n�2�hU8\���ї����h����Y��ɸ���N�$3w,�`��>�K�\O 
 "6������i�?�H[��e��L�q�p�,|�4���`FY���r�y�ג��v�ְ4+k5·k�z�~� 1�?�ݎ^��2�.X=�١��+_A����kLIy�,{p�3~���Ƙo�v}�����UN��Ғ	X�{�N�`{Y���C�,�v ���o�S����������avi����r���d/�?��M��%���n!�w��΍{�l���#ҁ9����������h��|^[�(#�4JO���}p����N7/�Bber{dq�]O�cԦ���nHHو��Ќt�\��9@�93������1�㤝_�d��[�7(�/��?�A������0W�����Ks�x��]�C���aq�"�ga�W|�������6�\i��t��7��5L����d&�E.[;s���x��1��XyT�3��V"��;q!`>��p'o	�y�v��+e��(4�`zh��*��Or���i��p���1ب���㛦b�H�-g�i
H�md�rX=��)�p|�� aKb�,�ZJ�t1��̥�&k��B�[���A����=���GD��ꁭ��Gv���eu��|LZ�'��|����8�G֩��+��#�]�@*Ut�2� ���qXH����2=	�E�'$�?���Q��b*�8M�����|=*���d��|V�%�|�`��m����>��R,����售���.B�c/������W^lpS�����֥V$^|��뿳��<����o����/&��}�e�a���B��|�� �k	��I���=Hs��U�&���e@Fс?i|XtHJIb�B�ԎCm�v:y�
A[X��5<F#GC��(bѼek��3�!z&�4����m�x�7u��r����r���46l��7��W�&v�+0�5HB����Z��xm2r_�g����x��X�y��<	��Ќ�5�Y;��xW�e���.��B����&�_�%�X��|��C�I��)9l�A�Ԙ��x�Kq$F���`��������s�uCߑh�g���\|�w%�b�(Ik���ʴ���O2�E�۸GZ	SHQh��y�������rc��T���]M�����ӏ�؎�-G�w9g���ݠE���j����!n6����D84��t!��lˌ1�t9�u/#m�<-���q��M�� *F
r ��t1�o"���U��R":��b7A������QQ�t�����������νy�U��b%��	(����٢'��f���V1Q��qE޴�m5 ^���.2������KE�fe����˩h]��܌�=��h�Q�Nlf����6{���T�*Da�"a��f>X��4@�Y	TR�&�ϧ����m���w��y��JJ�zz~{hW��Y�)@�dNGb�,�$1�]oL�q
���B�-�(p먑��ɗ�L`FF��SN�b+z��̀7IV�	�OU���a�B�8���o�D96%M��H3E�Gf�=Ԅ5������Y,��U��?�Nll�	��K�WJP^�yJ�,�e��@��r�$9��l��;�D#Y����;wR�ʿb��,������e�����i���Rth��s H�X�l��dt>�U��2���uv�e$�BMs�"��'QWS�z�2�P�e�bk7�A1m>_��0V����䢋[�R�ϷU��o�\9Ѹ	!
���u�'X"բw�tF��ܨvY�	�ݴ�҉n@�7�cF��	|�L�Myw(����G`�ɭ����j��1��ԍ�*v�;�2b�0��c�	X�8��p�;&P]��@G��}�F�ÂA�<��W�4�Ԓ)��ӽwG��MVնq0�<����