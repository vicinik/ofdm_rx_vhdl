��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�5�T\��s���6,]����Fd�Þd�* ��uCL���+rj�1�Q'�A�Q&�j�3�P>>�O�Xr��(�D䌧��@�Xy ���&���S�ۜ0�$��Hxy�hU�M�8�0L�5�6��Ζ>��LE����)M��i�)���D�����U@L3���������Ŏ[^�l�>�شz|��Xm�dIB����'��E�����f1M8J�1��Na�O3��H�u
uY�¹&���.��;'X~No/#����O;4v�S%� )�"��v��*�#&(��9�Ig�ˠ�PQp߅��u���m���e���P�ei���<G�,|�D�}�%,� ���p�>�#��"S��y���3��w_Q�?4_]83C`{�
�.K|#�;��ȓ�xMZ���=��
���Ǣ�>KKSC�.S����|4
`I�}�G,*V�zh�6�#G*l�i��3S�i3����bq#Y�T��] ��7a��UV����6�Z2<���ՎE���+x,MKx���+�VY׌�KC�_��@�!_u��b�]FHR�47����'uQ��e7�z�N`�&6��&y`�Y�>��Z'�5u2�Κj�r�:6ݨ���נ`<�w�Lr�;�R����a������S�nn#�+]��D>�K�+�l/��D�G�VE(66�1���%�� y���q���w���w�GQ�g^{E��;o̡h�[��ᱨ��fQ~��|��98���$��*È��)R�f�^Ф��N1X��j�k2碃x���es��t-<���\Ҿ)x�x*FF n��8�u�3��)[He�̍/����H;�\��Ϫkr~�� ��YpC�v���d�Ԛ��xJ�]��/Qީ��JZ��}A=Ff�ϛ�b;z	�`4�1,��0R��,x���8�g��Ѹ��8��LqlE9^a�	Ϫ�J�:A�9��j]P��B��/��`�D���ՐC_{]����FU�����YB�y�W/����p�i�7Nx7T����r.JL�3� �i��Fb�dꇟ� ,�Esʟ6���?�W�N�P��'<�r�7��,�r��p̹p���C��eN�
Q���)h'f�
�z#�����Ky�Pj�C)��,QI��{]V�	�v+z�Q�$�����p�Ǖ�r���+�^a�\���m��0Q�"h�w��v�-�i�^&�`����;��[��y|҇�����t�ξ3��6���*�x,!W��b'�.�����}��&t�嘊ъ��A$n�ê)�9T7��~��N�%!�)��9�Z=�������+�#Ȧ>�k����T�ڇxE2��b�"��w��!�J��W��%�OAzB|��Hw�<�W�1)�PJ�m����*ǧCk����ՙ�����}ƾؔ��~��מ��J&��iVKɇ��إa0���H@�%�j��	���r��6t� "���0q����G�R"0ӱs�Y�@l�.om����A%��q]F�)�mzU]�>�Qހ2CNpf�{�ȳB�ѓv��ND\`5�Aڙ��l�1�;]鿟h��5|�G�v^Z�=R/��X�m�����0�.�Zd	��O�z>8�*��W�:J�-#�8Ƨ0.F͚9�]b����l��>f��ߧ'�B.G�¤>mh{D�xu�a^z\�,1e�����=⪋W�I�Mو��m����l�贒A:_�w�x�纉.�ޒB��cDx$��e���}'G ��BRi�k��ER��~�QֶX���n839�Z��UN�B�������h&����O�s��HFd�GaAk��I$T��`�Z6������)�!ܽ��E�z��*��� ���9Z\`��*������w���c�� )M��a�dd.�gNc���Ĉ�O�q�����������U� ��5q��L���!�����f�[_�Է���cm��V����A�He���*D	�-�F�lҲ���/�Emʪ�����Y,jvn9��&���gӼ��o�f��?G#�r�@A.�Dhʸug-\�ц�+��I�@�t�"V�#ۘ���qZƓ�K*��/�����(o���o]+�0�<����?���u�5��Ό�nv5�����M��̪��5ɘ�Q%�q){A7G�J
s����)�DL��1���X%��Dlxx�NA�@��'�Tq�Ndb�р�Mʜ�!gW�F�����$���Tnzb����=L}�t��|��u�p[it��59�?�W�Z>K������1(��Yҷm��2��J	Ԫ����+"��:�N&�4�K�Gt�A#�A������%x�]��\+��<���l:o��S���L��ZK|Ck��cča�N����� w�<�I˵&h뜥?V��ϱ�V���r���W��6����=G�:�~FO>%l����³~�?:89o�uB6�7�qNۃBkB�U���සP�r���	F�t�zv"�r��8R�%�AC �m���17YUծs#�3X�	����[���\&J����G��n�Y��%9z��X�SwA`��.L��1�^��{L�Yr�s�$0��URg&�ם���m�;�\W҅�՞�Hk_�T�;y>F�� �� ����I:�n��'�J��	x�7ZR��N~��i��1�Ԕ��ܯg07�����@��������i��§km�g
U�����k䃓!l�F���c��3av���Ń8œIb��L�'�i��3j���W�o�z��+ko��.-�@e���v �����O[O7Td�ȴ���w�I���7}c+Qt|�T�Me��I�X��3�W.��w����*\�,�K�2�����c_3#߇c�垒K���q`�YR�bO"_�H����v�3߭���#"�I#o�Ʈ���,:�"b#]����US��]Br3����\�(��~���o�rqmQ�U�Ǣ���(�E2L�<�!d��R ���{n��zÛ|�d�ՙT�c)���7d��d�~��Ԋ���|��D�Q�u,��"�,m2vHD�K�'Q�&"?ߜ�����$G/e�a	أ+������ID�CnOg����\�5TM�!�zU�f�-�ì'7j���@�O���t|~1�b;�Vl3�9-v�!2' �4֨D�`	Hb���Vn�p�j�=a6���ڜsB���r�*��'�v��|i��� fFJ�ژ��#����˃���w�_�؞�MN-�|�AY@WH� /ҩ��׷.�`�zܞ��G�(7ei�<r*�R�G=m:ؔ8�_���(��~5'TaYFy��z�lEq�?��?&�]�8&�P�7Mq�ܓ���2����[��"ښ��X]U��:1�P�����M2�"E��=�w>J��M��7B/�y:�D�L�}4�6;, 
��?�����j(P�p�6�Q]zz0�ĜQ�F���OQ.�3ʇ��e/���el��/5� .g���$M��t�ަhlRjI:sT�M���$�+ů��\���!��9��0ڮmbD4a�y_��w��ġB��g�g�(^G>�J#�hȡ��4�ן�l|�-5�|W1#G�j�%����P����D����/]�RI�K=�_d|.^���6�+��?�1�
MlB���t.ա��@}�P��*���es?�o��X0�m#Vm�d���V��7q�f��&�V�W�c�T� ��vlﺫO��8WǠÁ��S����#����b̗�����A��\l������[_ Fy%-oT#ǇQ�$$�k�HtOw�ഴv�m���@H�����,ш�>����	*a=-�;�ŸW��|wC����w�cq�v6�F�\���X��>U%. �\u5{Y�U:1.z��(�>���w���	Ā{2z�`E��A����<��2�bû��i�1����7���׹D�U`(5W��&�'�4`�v�O_T
�e\�6��;6lG��n/*	�Գu�B�(Ɲ�T�Q��������"�͠����3�|М�u^���LI��V�;Ne��$)|�S��i~�oE��M�{q{�a���{(�	8�vm�lLr�R�L�#��9�v���a��;lgM7���:�d��0��\�@�_�L�sձ��+���>��w<��.���W�b�s�ҳ���4�ֽ�ӛ_DΚ�0wK�O���gN`six_�-�i���f�Xz��'3�NO5������"�$��Xi�BA�S�k�����?����Jc�6xYǔ&�������p���J��'���o�1�*��(�=
n�&��=�>�p��Y?���V!��
Na\��.�Xi}����T�K]b���N����K��`�c�o�]�a�Ј��̈́�l@�K�l2�oOJH�C�S�.a��!L?�'+m?���>���esuw�����ٵ�Ô���k�,���w-4�U>!/ÂO�2l���i�f	b��S.�Z�Q�������Ŭd���|:~e��1FX� �>,J�>�F׀�$>�
ԿQ����^s�L��,��u��!>�m(�Hu�ЄP'���z��� �R-̊Y�$IT����3B�� �:!���v�f�k+)�m�@.U��W���I\x>�A4���1�Q�۳�*G�I�䝧7�l�O��|���+9]���{��Eq�<b/GZ���u�s3�"����cI��}��@�������8y[�~�|���s�uސ6�J%%s��x烵`���	-B��T����lN:��<A�cvx�q���Gf% ��y3�q��@d1�$rQ�o��#�[R��q@�<"�o%-��P�I�x��)έ�H2t9 ����Dy��	�,��|����Mk6�詊i��@�,�nU8�!Y��${kݛ(y'vz�f�{ϟD
�c�1]� 0pE@��p� gc�=�I@��<>Ĵ�Ȳ���6\�^�	C$�0��:ĝ�w�!F:�.!��eQ��:'̊�8eL�rm�����nk�*�q*/����*�!x�
g����ec�.�տ�ƭ\�M:���dQ�a#|��H/�M�G�6 �'��r�w��KhzEQ��s�(����X�%Bi�������d�[d\�y�%9��=0�Swb����^��ߡ�`�u����D2EI���OK�do�C�Mqz�aA T�̐]@[�:�����fw��*=��s��f5��'} ��=��/P�4�/�}k�����x�	�2,;�z�cW>g��~�W�D�گ��ꭒgj�X��,`�P��3ٌ���4@�In�Ś����8����w����ck
8I�+���B�hjEk��M|)T�mT#(����s�oz��CH����k�8�i5i7ؾv��*�%H�@3����S(���FМ͠n�C��|���#�7eg6ߵ)��2�p�c�̀(���m��Kh+y�5ջ��ʏgY�ɕ֑�̀��a��yq�ZO������O,bI_.u�I�4�/���_�`�� �A����MNQ��א��
_��!`[��WkX=$ ���\�e'HT�Z'�O-,6x{���s�c̮���<M�H��P5��J�f�⤒D��d؏�� ��8�5_F�8&��߽�r}���f�R�b&b��7�l�M�_ )��E>#�۵E�x���,�1�p
9���v�r8C�� �ҥ��ｳ�?�"��P�V���>��;sE�> �籢��м�[��s�4?�"�'m`����d
˦�-�<�5ѧ���B6�3�u��������>F1�>�}���`�Z`���r�+�M�R�㑿ѵa���]�,���y�x����zb\�}���t�H�.?{�-�qK-��ui�}sW�
b��W�%���g�{��bT�Oo�ά��L����ik��!_)���20aF1����ܛ����bF������e��Z��� �<@Sŧl�)&�UpM;�@ʂ�q⋛�ѽ�;&~�1rWt{�!�M2�{>tC��H֜�y�2��c�_fwХ��병��_d]^�*c��h >X���9��v��I��j���]�J��w]�OJ�h'�x�C> [��Mp�.�:�|�vUbi*�4ٹ��T�+��;�'z����.��<�l-�$hr� ��>rdw0[E�/�]��{[A�����G�m�Ȋ��Õ3�wU�����i��X+R��j�a�ftf !���[ii��U�k�wz2�����Wu��J�7�~��T�^��S<�&�Z��)끂�80'9�*ɇJ)��n�n@_P��F�DD�R*m�{S�竅Y V]���p�|�r{�Њ�Hó:�<��l��'>Ug���/_���įZ�����>53������J;o�Q�1{A��W��;�#Uo�
~�$om��Ji��A�P����J�M,9�jT���-n����ˀ�̕D��9!����Z	��%Y���ySOb�_z{1�Ĵ���'lpg�8�+�Z,��5�?�}�B(-���,�k`|�o(��B�<�>Z!/Π��T����T?&�i��Nt��M�z�w�
�����@Αv�S�L�y�b�����:�Ǣ��$SC��5���R���娿�ȗ)������C=�1#��" B������3*�{جHD���lpJx�����HJ���X)F��x����k�ic��F>����ü0yf.�=u��-e	/ ��!�а.W=bd:g`���..�K��aē�;I�^7&;����g(���Q��1���ޞ���̮���6�@C��?��#�n� ����;�#� B���.N�6S`Cb{�KF�I���2�^�u�N�>`�y+J0pL�ٜ:�����۹5�F��5�������T-7x�-���k��u10��GZkb4-M_��T�d�κ�f07a�o����w���z&�^����ф"���6 �N6�gb�SuC""�,�W�G���x��nD�����w�N���j���7iJ��-zu� U���8���v�z�M�\��b=�fR����x7�R�^��.�k�zG��[��@�/6�3��p�_g�M�:_rIKjly��Z|H^�1G�_�j߈�@g��U5P���H].�����������^�9�Z��냩�l�6D��(�`,���27���kJ3"W�nK�u�Rb8�?��9sp����ُ�$��TDsʧ.�m!QO	]�A���:c#zg��	m��r���g٨P�,>�g�w2�b�j����ΐCѡ�G�FQ�$bp���|�=���|�>H�Qӥ��������e���:������쾲�(޽卝^�9h��,pA�4�VM1w^�B��=�a��������>�U_ �"!��ɖ!��R)=���mG�M��H/e�Q#��CE!���������8eRs�s>�"1s�PdÀ@����O��UZ;}~��'r��o����#�X��O���p�7�~G߬h�d��Kۃm(�W5��J�c��')m�c!хO��Ѓ��ݯU�X )����V�J�nC�oi�!�������C~��t�Ύ;Rl�m�cG�c�%��nҬ��k��(���`��/⼷��y�1߼�@��7���1/J7'ʗ+�WU"S�2�,�_�W��+���o;�k���v6�?���Źl'Z�M�X�C讐*������,��]X�AZ��H�{#EK��Ͳ���El�!U!7�Ci�?��8���AK�a�y�YԯW��$X��y/���y���� 8�j��7ViO v�F.2��_�~�a�W��s�XK��ۨ`A��*%/CF�����Դ�YQVE^ú��ɽ{Y�7x&ڼE����Y@E	WH���u B�LO���~y������$�⦨�qge@��u��+W�X��D�.a湅y�a_/f�y�����Y�Ni���tV�g�t:��/Z�\��d�[5m�,;��e�����N���j�ѫ�j[p>�[�_
Š�3bb-NT�5�F�T`��;[�R|MuF��0j8��r-|��X.C]��8�c�AQ'�/Z�;�bV�����!�U��s�(v�g���O�|�f�Y��ъ:d�����%��Z�CzT�}�y?7��5R�T� /�R�=>t����ۋZ&��3�1դu�G�S*�����Z�������O�a�����hf	յ6���5u�O�<��V�M	��p��\��*=(�BYy�����L*�$ z#D]j�,���h->�R�`!���`���ю�t�����R���f'}wŃ
��|��c�D�'gy�!������/VAL�6�� �>���k�����Ңy���Vr�@���G�ŧ��>R�)S��n��w��򼢰�j9W��&�샣D݄�����9%˚���r�%�c��w,	����k���D��m�列������zn�����c|D�i�w�`!�O����>�U<|7�ܥ���ӊ5����oQ�O��-�&�+dR�:� D�'��OM�����j�{��B�Yu@��FR��q���o�����ҹ�늏sl[�~��J��-��v$�%Р̽c���dN�0^�M�M�I���n�],����`z�&MҺ���Q=E�dl�M��殐=�Қt`�"m~ P�s{_�ѧ�!yD!�n3��%��B��X"|l�Qb�D�.rdm�+
!��`�K(�\��iS�V�6��[�j�����[�8��H���� ���;��J)(_�E~m�Dk��Ó�'c���� ���bR�SW���p}�R?���1#r#��"J���q/B05XTNDk�gց��H��耖T�oU#����JƳ��k�+��	D���J}��QH���3k��Fѽ���R6�i�WJ���<�z��z�Ǵæ�<��:�F��@��L�.z�����h��a/+Zz����)h�{:�Ry>΢|����+���H6�	��	�s��k�h�H���De�AE4vOr7�V7@�#�AF�'	Üv+�&��a�Q��aY@j: