��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒�GD_��Iy����[Yq�W�zr�uj�ai�Q�2�Pm����Q�ox1I�90���>~��R��m�T
�L�o�(���C��o14�%0�m�<ԝ�xz��8]�d����ᮉ#&*�x�L\S4��I�R"���b)ܠ�����_ԓ�b�V���j7���?F��2H�ۏ��<:W,sҙ8��.}��(���=����Mx����*���u�JhR��Y'�|�)������c���k�&���w��۳�W&����m��y�dO�8A�� ���}�U��#ʔ�w._g\���Ǻ|Qջe�����nE�U4���3NE<xC`"�$�P�|�1R8�����H
�&4;�Ϡ��w����o��]��BM6�X�Ŋ\���������������9x�A�KFN ��>�Q���a�'5�<�݆�!�PP�7�8�I�#�|��;i�\�	�b��}��E�U�����ȗTi�,�.�P���s��q"�H��_�\[}Q ���1�˙�l|;0i*ŧ���:�U�$0��n԰����O"I��S!���'�_5,vS�.��ST�����A��� ��C#�[��A��ˢg������*^��Xc���&o�n|�2]�DJ~����ߍ����#{:"d��[�d�UЗ9�=�W�Op�tϻx)ou��Bj���S��-���+N= _>�sT�W�������׃T�l���|HٲPv(�ZO�r�e���|��x�f����o0Q,`Ί$��Ã�IM�dC���)]:�5���Z����U|�q1[�b�%«��w�� 5$>:��6� y	Uo�/K�S~Z�c�^#�Y�y9u�B0ӏJ� ��l��=A%h����6x@����N���9_�nޙ|��3qZ�]���C7�	,@��Z���~:��zS�J=�K��r��6��.���7F]{�o:C�({/��vΆ�[1~����ӱu��
�ʜ�"��X]z,�M?���vn7V�Fwj��Y'm�1Q�9`*�ͯ.l�k�/Z(Il鬰[
�r�~���\��ܰ��|e�ti���2͋���Q����^����!��m
J���w��@7��̭lkȺDH�[�u;����גc�����2�qb���c��肠�,fj�=Y����7W���>�;3���,2�gQ{��'/)ڏ=�!3��&[�u�xG�lq��%\�k����W�����"�x�T��ߥ�}M!��T����K�������I�m�5� �Ο5�oJ�`�SH�X)-�R���}o�b�ʔ
q�`���@�0q�Y��d�/y0�n�!���oS�뱦�nP�\b�M�q@q�$�I���kD�#I;�����f��Y�u�e����߄ 1k�\��n&�g�,�.;�*�����J��JS��{ǎ�k4��sM�p��䪑4xN�� #�sF���b�.��E���pA�|��!�S�^�TV���!|ǉr-9RШ=���,S�DYͅyz&�\JR3�MY���Nc`��T<�I���m�tɁ,��}���9��踍~Iػ��B�L.#���F�փ�N��c���Fk����st�.�ؓj��n�]?��C����?Y��pyLt�F{�֝���W�P'xw��ia.��6��c�Cا�?m�4#/�m���Zf㪤���67��:��oh��"�'���n�0�>k�t������!Ы�l�F�S7T��	�}�(�Ó�y�R )G�=_4�`��Q}H���Θ_��[a:%ɏ� �#>5w���
��az���!��P$8�d�2����:�� ���A����H������L�myw
�`btcPw*s�2et�>r5�y� q�F�����0���,9�9�k/��\i� (�vV�)��7����L�1X��R�_�]�h�)���S���a�~�L�VaEdA@�*��P��`v���)k�VR�0��4�ǺPs�����/i��9���o��Rm�z8�k7A6��#U.�Q��� &_Y�]8"{�/������g�;-��<܂{�q����:]���N0�ŋ��C�,�"=��/?G�{:*T8h/�)��Z�DU�i�}����f_��k�"�j�.Ӻ�6�c�x�>D��L�����s�X�|�(~_��z�#m�� �<��o�M`io�|�׻A�R
BKh2�69�Z�1*���s��
ρ�9�^p�i�.�O��� ܇f���[v_�3��C=��oP� �jڟ#��h�y׉�ڃLߛ�5$4���l$�LaŪ��`	$�n�>跈D��.�����?:wBh�mʡ���G��s|(4q�����	�aY{Ľ�2�Q�a3?�u[>�9����l���-�vf|qk�vN��&Ӽ$����l��۲���P���k6��,rH�l�/\�O����R)�77�eF�Td�}��g�o_�l蟞,7��74�u�'o��	N���+����)�BL�0$Ê���-m0\J۳`vL��`�*\é�������P*�D<m���^ �M$^�z�"Rl�-F�fu�o��O�|	�Ξ�9����n8�GU�Ha c7��>+uQ>����L��fT�y�P(����тeh��[u#�ި�p �S�E��۴ �K��JJӱ7���V%<왭b]�r�J����T���J&	�u�����dњ>� �K���g,�A�Ͱ��Q�8@ƅ	A؊���c&��秝�68����[$מ x�δ�{���9��1.�%�[�t�1��9~<��a@?���="���=�� ծk�(x)���н�D��Lb�nCׯ���2�.�gz�l���0�_Y���s�����ׅ�8��^[���QH��O{��KR�h�OŲ~��iS��c���x������T,�����G�H�f�b�_R��ruc�X�L#S���+ 𬰈͢5�Jpל�k���@Ȇ�3�E�#��No~Jc���h����N
�M�^h ���أz�6��j���D~M&�m��AG�8o�"�kE�=P�	r���ܴ�ǿ�MJ�W�z�<qԉ�
w,��z��ݱ��8v@nNH���T�����FC�HS���*V��]D��h��e����>����L
����57���k�m{��SHnL���Қ�y�~���˰#:��p�R;�YCi/����1�4��b�#w$���g>���愉X��}��8������:	��$�\��/�/Rr��#�bb:��`Iy��͟[J�t>:C�2��v��_#"�������q�����w#`�.�r2��T�+�d��F������l�侒��b(�dm���8�)s4��t�6��A���K�R�hE����Au��Hs"�+ބrFmtW��Yֻ,��4g��_�氝��ssܲK���W���@�/J���A)ų�[�mr�v`�{R �)�|��(@.G�g��F�P����%{{��W�����.s��y���iW��m�e_0̍p_CFx-<����F�k.�r�p�P����n�R$ ��S?1���iKJ�=�T$K�%�p�XRx{\���0�Y����x�]��S(��􄘲����А>�*��rf�Bb�'[t��� M�%-i�._s�T���ԾǩW[ެ3�G���R�
=ˮvQ���9������a���n�������F׏�;^�v1��"S��{��Gm�������Cu�P?)���M	Yc�|�D���rWz��N�z,�����2Z*+��C����F`��"�\3
�܇}�d"�����ϓ�t�{eqw�� ��,�?�OM����}��a2��Z>�ZG��4����9�eg+�k��Ē�揻����>��
B���N����?X�mѱ����LiG]Vg�; ͇�;輨(%$m�j���obc|�W����9�DC ���#%J���i��w�Q��>�o���ʺ�*x��q�ۋ�	�q�L(��������X�t{�2k}������[�:�W����ɓ/��!}G�UR�8��+��dR]��G�/ �N����.e�3f�ch�HtڙO��G�P��Ѻ���"ň��ԗ%���>�-r˹SQ����)�V���!��Xiظ���H��N��e�|��H�Ë�n$.��H{�(d�w&�n�(�����&�F�N��]����ReS�	h5��'n���lrX�a�-ʜosc��+&}�j���B�֩P�_$����q	�ת�xR�(��F�X��u���_�:�˫������X���k��}����2ޭ����rPL:�7 �|��>�5G�w�$
�ip��+`�����ׁ&�������]�z���_��r��Xi���k��,J��l8�7C�i-���^�KC&���/t��4�/�s��w�3�	g�C�A�b��K����Ԩ��-�n�R:����So�ہU߯.�lh�
�p�=3|}֑��*qM���l	��w�Ǯ�rPDZ�_�j�@&֣\&ӧ�Y�����J	�e�Sц�^�X��kcօm�l)�8����H	Yu�Y�_�-��7<��6�~�[{�t�1*/$#)�˷W jх�p�/W���o�I�5!;l��=gF8���K���Zmu�9;�z2����^��-�8כ5^����ƪ������9�w��ADG>�s"]�y q�"i"�{�i�����a��m�b`�xx:Z���yY ���Ժ�����;�|!<�>b�ۿ�#ب�M"�k��a'�NZ�C�5hK ���v���k��la�S1d�#�C�N��J��h3A�^����+Y1��t�N�t\�[�?�P����(��\g~u2-ݪlz��>��Gy��sjS(��,���_��nk��MC�͌NL���?�pp%O�xs��>�0Œ��-�O�2����ZA������˵\M�qK\���o�C��2�6+�CՓ
 L���`ᓻ�"{���b����[Y�B��(�>�Flx��h�\	���� 5p�,/���mgY�����zme�8s:�3��e�?t��۳�qBE�Aۥ+��{?̤|-eLr�VLF9�pi�.O���hc�{�qh,����S'��茊!������Kq��g�OA!�<נ6�V/zЉ���f�AZ��x�.)-�Q���<���Y��Л0<A��o�P��2!0$9�۞9���]l��.�����:)���~�~��|J]蠜X��R{'���p�v�nQ�!��i�@��X�����K�;��<(�`����%;;��Cz�&�3��Դʉ<� �L��"u^�8�m�����rm�ZH8,���~�P����Kn�w)Y=����0�WWV�j�{����|�Mw�6-�WH���S����/ϙ��/]W1���W�De����wk_�i)�6�E�(6�F7�NR�|�$���V�Nc�њ��{�׾C(ݶ���p�;󞫕�s�%6#����xI�TJ��#�l�T�ۺT�Arbeܱ�:�fZ!�H�:��GN���)����-Nkmji�8�&_J�X�d��a93K�."��S8V�'"��V i��Ι���>��e�NFb�<ޔ�Q&�R� d}���.�A�j���T�.��EH|z�//V���W�Ŀ�;�Xd�����d�⎛ڶ���Uԝ����O|��� ߈nǭy��Ϗ�5�g�A$#<W��R,��g�g����2���fid,"�����Aq�n��M{}��՚}���paK�tX���h}Y}��`iPxˀ )��͸��%��ӝiGPn#
�L�2����d�-��o�7�W�0��
���
䦀 6{mcl�t�l+,�f�L�-����q��}s{����cQ�9k��cD���4_ؐ�M���X����;�Q��R�Xh��>��Y�µ�^��IC3U�`LU���<��q���/�fJ]ƀGw�YcE+�$Ús���!�$YM�F^�[8ç\ ]�ﰮ@Æ���	f����=�p&R�ԛ��Wb͉�T
��VW�|������`|]
�����g��&��_d��eKaCę��j���*���&;R��y�T�M�}�R ��3���g������T<m�<Ȑ4���IZ�-��B�����Z���{P��>j}���(�u���7�n�}�U��F�6`���t�n$7��-��g��)��xD�P�6��6>�s�H�C�y����ߚ0 �WJ�U\�E9qy��%��Q��O�������}f?��P0z8��-=pɋt�,j�@�'�7����7�RHzD�E�=�Cr���.��Rn�%���Lm�f�
-�[̴_��~�$��P���<��^��r?4��u��Ze�D���M\�2�|O�M�k��`P�N){$kڃ�V�x�W�	g�Iߚ�;�f7(�,�J�9��>�^�3^?k%�5�ͫ� c� �FG����؛	�:O�)k)*\Ś�CN�xA�0����^d�{9����2TM�@i!��!7��]�5�N���5�����2��بl��P\�j�d�,�"j�}rK_��M��ծ���KU��q[���-�0�����e����b�R�����M�i��� tM��cx_[�ADu���۠qJڼ�w����a0�h� ,.R�~��d�s�L��O���s�Z�+�N�����w�OY1���pC�V�k��Ű��3�JJ�Z�|[�$4Z��-�LO�����y^Tn�~�⣜����8@
ң���D�ʙ�E����q{���zC	�Doۚ#�<a��0�HT�g�q��"�z��f��]1b{c�����P�����񄤭�jV*���;��4o0�3ˑ�~A���;�;�&O���wx�g.o�D���{��S�r��y����Ǿj��*���%����JIp���xv�i2����D�݂?\�B�?�G+X����5����M�����$��:q����'V����ϧD��
�����~��`|�1����1�3_`v�ͺ��m�7�
���y�i��%����T� %F�8��z�X�7�K�.F"Z}��T�2�X]A�w1s5-�wɕ�/^�GN�`��>.md.���>yZ[A_�㢨���L��_��q�2�V�}�!߸5��,N�U�06kϻ��j�x'͜�DR�Hv*���v�;������P���M�)ۋ㝳��;�0%���(� ��nS��ز�Q�`E�]�ؔz�Y��$b#]4�� d�,k�{j�>FG��S�5��xx���?m�M�(pi&}�g���E-[��%.���ٍF���f ���"�}�O�)��-�G�g��س��( �􍚆؂)�p�ܫ����T	��Ӊ�W���Å\cF�L��3���V��)YB�l�H�oAK���*�.m�+�����^k�c9R���EH(�U]�h|�б��%^ρ��r�il�^F�s��pZ��l�4)7;�z��M�4��>7�N���)]�/T�V�!|n�a�>�x������Y���#te��|edJ�!�k����!xՊ꓂eɍ9�	�(s���f]����\�$�>=zRm�z�Pí�8-YԮ�(�b{U���靓z���EE�`�L��'_�Ky�6$~ߏhyi��\��;:��R�������&���⥲({hw�.�HնP_��'X��Uk����� ���#kd� ���_Z�/������xk���W��� ����Wp҈g�jOg8�~C�jNE��G��f��ѭ�g�����Xxi_�&�#��9 �x[Vn��f��$-��]Z"fG�A��$]���Z�E�	BIH�+�Js��F0�}��s��"[>��`����j��Z�']�;*0����'����ʵ��$3�����r��
�+���J��W��R��K���"+4�r�y����U�׫��Г<�d��f/�Hhy/�_UT*��$��6ϖ\�� �{:�.�Ȧ�^�.�Ձ@T�[tzG퐊:&u�-�&�Š��=�1��uo�/>�6�@��31��{�W\<j��:rK��H��HeU� -�چ�-(w���@?��V�#'��&T�O�𮮢P�0�-J�$=��)2������������v����jX ���e�T\����'�efc��5��q3��Z͹��]T�&�m�����`0����}���r䧜�E��I���~������?ܥ|��[�lB9�W!ڨ�Uֹ�@���,�V��^�e� � �k$9�v�Y��f���c���?�X��� 0�M����d V'>�`V������,�����$#���Iz���۞����t�@'��(�|�>p�í�rf}_��oM��F/CᖉX��p!����y�%���l9p�~� ��{=�	�q�d��N�7����]��r ��*H;�m�(��Ȩ���s2)�VQ�JLP����W6ݷ�VeA"L�Uu���l4�
~uAB%�cb0Zd��-���T\�@�B`�[$� �8eX�!�K4��������*~�'tۼ��z���!�pNO�+���K��#;�-���;YYiH�u V�s6�f�V�߼?E�_���?E�D0�� >�=�3�@L��Z�\�콜y����Rj�H�^{�B�]+�f��E$�M�v�E���|=���Kdb����C����/ޅjV�,���ɚN�_j���kTZ59���F�*���8��{|Z%]�j?7]���A��3��c`�<'<���@�)��ƥ/v�<���e.H{��x�g7q���V�5��[�U
o�4��Τ$_�W��R�����&���^�01Y$g�/��=&_��5@�	0�暮��(c�c��Y��I
��~�F"8(Mj��K�ۊUI0���3(֜�H�7HT/IQ,�l��ٳv��Qk�i�Fo�pF!QX���,�}1��,�9~��\%�X5S�ܸR�ACQv��U�5��֟����6�Z��#>��v����y��EF�����E}*S}Z���O���V��B�eq4�R�ح�N;Ҙ��܌���G?��ٺX�k�n���)��iUQJ�V�����i�mt�144j��$�t� -�IpZ)��v�{�zl��&;���y#��T;��1�����O_�MKu<	��%��;�Kg�gT�-]�XY"��n,�6j�k�2�,�Tt&7�S	�fHT|%>*uJN�V�֛�7/������Tq{>f�k��78�%P'?�$��ㆥ�V�~ꊒ�8�"��hBp�t�����A��xj��9��@�`����m��t��0��lW=��.4�v^��0oQ�.��3=A�}�Z����kz�l�b��
-57���!T���l��E�b�N�I�q�4��t��G�G�����`!�5�:�";��e��bT� A���𚅮��!	"�ۛ����6�M耋
�uߑ�bi�^U���2�Kp��� �B<Z(���C B���e�A!�X�7R\��aN��`�5�$��9+��b�K�h�B 0V!�ZlgS�^�݋��cQl*]m��M�:o�j fN���0�C���PCtG�����gB�X?�^�_C�|{�Z�Ky�E]����2G'����H�*^�x�Y�-���]T�8V>�Ȳ��)5Ed�D��C���q�y�D'�o5�n��$�pu��4{�?�;ﯞ<�r���HoRB$&���v^�|���ك::��P��<�Ps_���ۚ5��>�A�����D�9�x���w�W"D �}��ʨ���RߋȲL�U���ԏ�@����M�̖3�0�V6L�j�u"��w���|��r�P��͕L���:pP�vJB\ðC�q�zƴZ�)�@z3w���q��7x/�b{�S�{���k7�@���f������aL"���%e�z�	+�9�	�t���
�!vO�Ns�8�/�����L�����k����1,3�??<W�We��!0��.���`��0����B8.��쏩��E�۪ ��N�Y#�Va���נF$�� k���ҟ��=/�SOMQqy����n[Q�.��:�5L�n����'8��P
����g� DC�k�.��H���ЄHM�;M�Ăq稊���C��8�0X�;�(D��@		��XU�U�`��.c����b
(�N�h�1�æ|Ř�ѿJ���M��E������k�DʣK����)�~�1_[���f�J4r&D�Pd�%-���n1��mgC���)���I�X�%O��d�
��4��$D��7��d���V�m.�����#H�0E��~�By<�v���ڎ�f���D����|���֙�-�d���P(4�wz���~�_�]����⍠�ㅣ�w�i?oM����{�s:����0RH������WIS�3���3�k)��g	����Fڦ���sk%�e��K,�R���&2v�-
�p0ƽOТ^c]�D�Oɱl�~"хB~���[ӘJ����Y�'�%�5����2�#����ޞ�A�uYG詴�����qm�ėPͭ}��!"A/���]K:uhT�mmK�?㭓}T�~=� ��j2����W�S
���V��y�'�ӹ��Ǥ�,[�<�+S�;~�ꀧ�i~��H�W�:�z22o�_L.�a��<3Sj�����"�tB��Yr��j@��K=�.����s+�Rbq�� �:5僭r�4}��D�#p�<II>�Ν�繥+������0������G_ʦk^5��(��<7��~:=1����-��f�4�,0ixs����-7�?f���#w&XuGo���,�!RV�Fa�El�g܇0۳���Ɋ����财Nλ�[����>�;��S�	�O���N�H��3�z�
!���T!k]�%���Akv�8=��3Oӗs̅=���<�1!��,� �^w���aQ,���+rHr�)a6ҌC���x*<�c�x��5�$H>����1�X��9�z:g��`��U�.�WH=���C�w�  �z���=:'����9E��P��W�����V����؄\%l��������%؂�{<na�йl�u�, ��n�T�9�[���ݾ�eg]:����� ���vP?I@�^3$��r��Z�k��L��:��1��6�n7YYdt�R�h
[��`��o�c��@���ɗ�T4/�{T�#�/9£��+TfǶ���#6��GA]>��`��N_�Z�L����RV��<�#}���Ud*���@�(����^Y��VI��^e=�ޞ?��VW,Ab�����G�G�E�M��g}��}�O�U��ٔcKgk]; kC0t���]�q��hn�	ҳ@�H���.��I�H��HYZ*1 /�"P�ΔT�l�P-��L32?��we
{�s�,p2���#[F!N	���x�~�������>T*�np�СdQ�`;ӐT
��+���\�j\�U�+:��zm��1��Tq�����N�r���L{��t��>O䗎"_sN��C��e��E_���喝�X��{����%������+$0A��ý�;�'Ft�ʤ���[��RZٖ�4/H;��Fm����^��(�4�&7]��j����KmN�=C�h�C�!�I4���F�*�L[�a�ɺ/m��Я�^�����~ �����d��һ�����\�j|��t�[TLY�y�X1��x��>>"�.{��QY�0��1Ǭ�o�E"dj}��+|'��U����?RU^�x���XT�nc�D��K�Fy� @��/��^s�h�_���K����_���ې�a��l�n3Ue��B7;R�l�~H�h���j��{ra?���n~�m��_
&� vj湞�����{8[ �,�QDE��JU�2��i�%��G]�*,�n�?���Z <�I�^�)�dp}��rg���y "�4�!Q�6�ַ|:,�IM�9��`��G�+�������N�O& �0�tx�6����*�f�� (#�0h&���������q^{z�1��qu-�&�¼��k�����w�^p�~��.�>������T�4�N
~�5��Nr><�k�o�"C�\sQ�ʇDg�� ^9�xGm���ޝՇnU�50s���2:���ám<���vŋߗ�EP_�u>Azh�a}�i��'��>
J�em�J���0��Lb�"~�I�%=  3zC�Hu"7��X|�E:��R��e. �dQH��u���W��Z��������0ڻ,����6�UC*�i{r��(9ٱ�K<J�~��^�q�����xZ�De�'��(�A���J7,��r��|����B�O�����L>�)���x�kh����-G�t:p/Y����o��z�
����[��nm�&\_��v!��=,v�]�=���������1���Sy��ܿ;��
�8O\��NYW�a˪L��}�^�?l��,�[���t�����!6��{!��۳>���O���V�F��#q�b�z��g��0�[�������L��M�������O�]�l*x�������ycS]^r͉�`��o
�3� ��G6뛃��&��j��g��Q�T��}a�g�񭽵��N"�OX�@�]�<�9�sQ�;AGZ���!�:X��1�W��=��mO�K�?���*��4;&f��j�j�p���}����E�9��a�����0�����q	7�{Ӽ�.�"g�Lm��m���$�"|-��]g��9�Vl�C�HL�tGoE�#��*�0|�h�U����i��"?K����#��2o�Fv�y7u�)�a���T�7�C�H�C�X3w��9ƥ�dI,B�tu&���"HٵLPqL�03ݡs�ɬ���qgE$8T�j�0,�ta2��k 3��W�T�K��M#4��w���oN�[왟�B��?l?��y�I<����{����j	(bW�p9/8�~1J�02�/7q�X��!��[w��0�l�%`�D��Fo���HI�pi������Q�ڹ��k]�q�s"Z� ��X�bl�l�2Y�]�k<�]���*�`:@�F~!:t�t�}�^��׳]�^��Mx�'V��� Db!���h���+��7�@b��)�B��'Y �R@|M��k��0r�H]JQUv_��޾-��`�Y�y�VByS.���׺ �	������x$�>Ȅ֩3�n>Xr<g��N/�����5�}�f";�#�ʓXY�s1��E�'������cwՎ[���9�NQ[Skە�`���qA�F=��'�>��:�����H����>Zy����0��*�/y �KNNDH��$(�������
{��K��܅�M���1�c���F��~�ؐ��N�IPA���	����<���"������PkHf�ƎJ� _��{*��T]��:������Mx�p_%��4��2��]�A����_���V@��dK������0�g����K�į9�vj��,�Q����1��]��=�I^����Ԣ~�Н���ܷ�nо5B?}���pB����ꉊ��� ߽��� �Q<�Q߀t�uR��C�����C�B�
as����ϑ-zL2Rz�Q;�ɣN��C�W�ڏw��M�����M����)�9�a��)ﺉ���w���Vksq8�3Z��[̛` ����T`ڶ���̦b
/t���I���<рĔ����c@	6Gs�d����RG�n��~�g�5�|p� m�ν{� �7���M"}W .���6��H$�O��*1��+��ŷ�6��w����{�ig)��$9�xçcD��̗x�ɦOM���W��\S��h��מgƁv���FU��"���ra6 p��r��zڶK����߀Xnc-�r�}��T��L��	�����,�]�P�/ɡ/��~�
�]�,K�����,��NO�5E�%��,)���)RJ+�%̀jE)���"L`�9�dou	i��6\;���t0j���	 �+I��F�CN�q�>�[c���9"e��ɣ��ts�7~^��}���!�'f�BCx�Bg�����iR�8k��+�
��ŷp��)2�fH��_��!'�H�.��ئ4듫s#�:�Y�˝�?�E����G1V'9��C��n{�o����.�
d�xB�K����K7�a�'�2�oO��v/�f:��lnM���OTr��&����,u&��oKoF�q��Ɛ9-��
�9���EIR�@�@qWi����H�1tN-�xs
��f�4n�PƆ��w�yl�������I>Mc�O$|�5��:&�_��Z��_e�ziX��C=4~��,�� ���rz5�L=��DJ��up���H��T���pF�J�����C�$�d���i�4)�/��q�s|��j�(5���k�,P����4�y������bs\�"#Ynd;�z3�X��WH���W�~xf�Jம��|A��{:����:�zSj j,���^���`(�������3��mx��i��~������]��AS�h�="cq}Z��f�K|�)t��H¿�Tc<��F��m=3�C0�W��a�T$Rg߷ʧՔV>.��dZ�u�O�'\�"7p3�-m}��0��,�����fҭR@�.-t+��A�������c����=��E����@[�ݪ2�$�[S���S{��o�����X����e�]��1��ľ�W��/�]6cB��'��l�ҿ�d4�Xʮ�d�(:s��ߢT��_�ܐ���p|��"��m��/� �!���T��G��J���%�Dť���e��	�s_9�ʦ��ƛ��-<G����_uXx>�^�����r9��q��u����3�!2CØ̄��f��L���4�`2�9ejd�
��Fm6��Jw�X��W��k�	�c9V�_	�&����K������?�4�|Õ���ޮI�f�0ܜH�f� "_�V��d�{S�w��l�k�QW�.z��~�A����G�e�hi~��u�O���gGaV�m�~�O�h�c�D�_ӶҚJ�ضy���^��ajJ��A��K~��An{�=޼��os4��5P�/�����h�
Z��jM�����0����nRX'�l�Gۭ��S�Ĕ�$��(�f�4�������5�'ǃ��Gu��G��x@��~��l�{f������c�|�?���l��sK�.��>�,���O-S �m��i}\����B���8���7=��i���w�'4em͑���@���GfkV8��	O�~ڬ�H�;���(����R� 6�	���Lᄙ���G.��W,����3�ZFhK	�,Av�z{���\qCr��˅���PH�ZL�t��F��.�d��0�"k09�\h9|<����눈ݡ*��1w=h=���<�l�gg)��%�?+�����H*���è��Y�jvO:R�_�Tˣ�o����臭��!Idfۜ�ʝ|�1F�Sj抽vpn{D	��`�ypE���R�Ie%��C�L�L`���0=ױR.��g󄔼�vp�Xf.9�4�rP��,��u�-�����Mk]��{�+�3Q%�7k^Ff��c6����pч)y?�������7y`:��!o6���A���"�׭d�޷s�³�I\��ǑP���CY�7�z��%Ņ7�jI����o�̣����:o`�,����nct��ك��&M�f�'�ݽ\mȟr�%Z��+��6W"lVE�!��(4�b��:�{Y��s#�ϟ���_�]�'PMxl%c�@��s�W&�V~?�D1-�K�E��Z��+9��9�����EJ2;;����\��=���5.yo)��}!R��O|�86�6Q丛	�E����s���Bay����� �t��N�W��4�@:�h�m�����5^�QBت��f} /(�/��U��9f���.���.Tc��%4ߜ��|�OJ��r*:i:�������YQ�Rf��<ѩ��W��*k�j�,T�Ϥ�`�Zw��d�.�p=6��׀F��V3G�B�_E���k�e�j�A�QEi�k^ʋ�Հ�Ǿ���a�~P���(pʺk�l1h����˕6�;��A�W�z�5cZ�2�?Ր�n�{w@��ND��.d饨&�n�����y3�o��F�����*p#�{�<����j��N���]i޷�t�s�`x�3���-�ܸFH�e�g����yL�Y��!������3�B4���Z)��bg�C�ր�j�����c+�Aj�)���zʠ����n>,��������#	Nm��;���y�=C�Kv�� ^[;U�i����G�8C����oUx�ec�I!�c(0Y �2Nn;h��7�������
�EG濺�1�`7u����E��v;$؎RS���υ���a�5\�1�@�"^�J�Y��Y�}�>>2�\�JU[��K�?Jy{�3'��GX�{2��*TTgaG�RJ�xB��u`�I�ce?Y��W>����^\���*�~z/�*�EV�y7�*��~ё���%�<#�����g���PX�����2)u�CɋI�N��'tf�j��]Q��0S�\��///���ت�8�F��Q6u<}�PVu�g��<)�d�.�$��ο5vJ�]���<T�\3W�]��ʦ�|���ngX�0�m^��8�z1�,�b�g͘ԭ�6襀q�[gTX<:x�1���]"3�a[١�������أDߡ��ߴ�w)Kq����� ��ټ0v�Ή�g@a�n�Y>s{�8v�Fb͒�$:��V/7-(����J_5c�Y釴����P^]�� �`�Wl��d�lp��k�@J+%�u�H\�]f�#P�z>h�rx�}+�$!g.�hu�(�����HwhZ����x�(6y��M��o�+�~��M�|6�_�k-��${v"Ơ�	�4bs�^b�K$ydW<�̨�G�Q�����u��þ°�y`�=�HҰ��[Ȗx�8Ź�A��C�OP$�U�?)ʱ?x�`�K�r��:�\nxJ6H�0ޢЬ�=�[Z����Kƻ۫�0�D�-O!Z��
���}?-�$���[u'��	��ng���C�x�!-��(�����t@�e ��H^KDi�'f߷8;�I�v/���
�ȍ��,�T�:NZ����҃#Ӏ[pC��[��$���4^,�`�w8�^�d��p��ee��L���� �'�A%�~h
gU<H��?��m :%c���;Z;x=z|{�@��~��l�N6�H�'������N �,�b?M�`s���=ۃ��=xPz�V�d��Z rΛ���ڰu���� ޿p������8˜����4�ANV�e�I3�k�$f�#��T !�/>jt<* -����+!+���"N�W���i�e�7M�C�(��"�/
�g���lU�@	|9'1�YCW#�|�D:FZ�����A����1pV�낫7�7~�*iW�ȣ:x�q��I�́�=�CSO����>�_�<�_�Q���)�qJ��%��as��fj%bj��n7q���%)��`"6�g�)��C����֨pok�3���87�z���Y/�`f&���3`ߜ��d�)��l�6W�E��)�`��H�e��QW-��𪑤����b'Cĉ�M�5���5�;��4t����'ѯ�=]~$�";ڇKq�'#,�gA�9���o���^Fz�*�cN�����v���֍��\�~�ܑg��Vt�Q:��-�W�5?h!+����� �j|P�o��8��g�PZ��#��<_�8|��O�>��a�х4���@i�2 {8���3���G�M̽� U�v�v.��U��@3;+)��L��������Q��v��8��wZ��Vgv�A0&������Z�l=`�7h��T";#T˨�3/�2`&Q^7��a�]�W$�8e��u��u<x&�j`�p�R��=���ŗ���S�=�pOБ�!;8�ڮQW��c�F��/�dMA���sg��^��c�7r���NQB���4н���iԝ��
�S8k%�諷���aa���E��֋W�`�5>$;@E)��>}?�� _����H>3���o�1�p���@�R5)�L�t�7�l����yہ41�))�0~	7�XZK�I=�k��*�sE(L���%AE�*��7�Kk?l
��X���
��|�V� �Rd�c<s�	�5$F�P�o4��B:z�I��I���n�ٓJ�����g��#@�p��WWЧ� �u���ؾ-��S�eM�)U_5���t4(P�E�z�\W��N�Ѣb)�hg=����`���樏F�(��d: �#�}���%��M'���ÿFa�I��Ί�	iu�RI�0+����Q�<4�])s�DZ 1}[5j�]��a�oً��.V�[J����"��#j��4��7^���Ι�ӡ�{�ǔڢ�������ǹ�W��%妪�5/��!\��X]'t�4~�ߩQb��ݤ0��u���,u�\ݟ��3�Y1N�}B! �p�^�
�zW�~+���{Yk9��,s�zG~�}t��ڝ��'	�eM$n��)�řH���|�o[���$�=��v�=lI����g�
P���y���W�N�=6��<�g�3�{ޜ�*�\�O���݄�z����χ���(?k��;�z]��H�&�ߡ��X�T
������i.o ^�iA7��+�{��g�?>����r��� MEAfT�iɜ��Z8c� M3��������t.�f�p�s����Z����w޳+�2�nA�,�*���:e�'�H�@�i̳��=n�M�½��"Î�����46��������]
�3����5x�3?����_W�(2V�Ѡ�~?���a7r����*�6`lX�J�-�v����aY��e-ܓ$�hE�r��Q�.�e� ��Eͅ^د0\�W5˺<h'w���䃚l�KccUl�L�'UFŢ�`s�z�ɶ�5lL�|��^LO��g,��+PL�1fJ�^c��k��!qN�!�`B�8���}x`t#����T�@���~��à�?Q����+�F�h#�B[��$�O0x��oS[ag5է8�͏���C< "^�Y���g
\d�������gw�C�	��O�'��o���r���������3-zѺ�������>e��w���+f˝|aW���װ��=�k��|����HRY+��#���<S�$S�Wp�[@ ~8������7mpR+aOV�u)v�n��&���aq��"�k�إcǤ��D�x5f���<�Un���/v��\�yjE�(Pɋ(��/�}kj�ӫ>!�t�/���1�)`Ҁ���0ŏ ������_ݼh\B����[��mXAc�b1����0%��&�1~ O|q��$�a��jw���@�X��7��{����[~�T�J4�iuXߵ���T�vVlPɓ��aa��_�<FۼL�z���l50�X�XZrn�`|�z�c��[�"x��9�'�¿��)9�&�ڤ�_��U���~t��z�j�u�	x���g�����M��ܗl����ہ@ɾM������d*�eD��f�^�P� Y;��c��2l�F��BIs�V�{���������m��y���y�mt����-���O����^`;I�c��C7��[ij��u��
���v���vmy8�NS_+�Ry�G�!���YQx�����V��\^a�8���V�s.o�ܓiw��Sk���o������9��yL��C�$;'We�w�"�y��	��� YA�sg���1����^�!�5�.�(�2�m�53��z��	��%����J3���a%�In*;��ǁ�����3y����ּ	�ay ���9 ��+l�޺�x$R�q\�fP79���H����E��\s���M}xMy����������B�e{����0$���L�B�����H�i\��.�����n�������_�r�r�j�w2�M^���V�^ø{4�m�r���#�
��	r�
������e?�L��g4Ƨ���X�Yw�kB7`ϸ��.
�%o�p��/a����7�o�5��3����w%8��	���	����ۻ�Y�=Qef!%x�bÔ��5�
�m��ss���a%���g&O�J��iS��O�����-+��2��I�̂]vl	=�- �<@�>z\�\Ni��Qfv,Mb�2ᑁ�����@��^;��v�)oT�
��q��`%���-Al�����N\���*�Q�Z�˭V1C�3�CPZ�7Hަ G<^#��x�0-]��!/d�
�tIu�A00ݨ�t�����W}��$r��Ԇ�a�����ЪY���d0m]�2�������F�E)b^۟��Yx�*�����>�/rm:A�u��QQjw �j�6n�F({E�F��o�p���!�;�9�<%�,�)ϯHj-��%a�1�Rx��0��>�K���/�h�R�-�B`c:�ȵ�8	���QN�����%M���s4�^��R���|��7�ZĊ�-O7-�f�.�l���ux��֠��j����'�wm���4��}d4�m�SJ¸ݬa	\�׿~N"��GHX���;�=�8�ӿ�e��m�V�;Hb��I����iҺ(Ń���wBܸ�z�L��wФ��eU�÷6�.��5����I�Qd�,��.cny����wK�O�H�[��&}R\?�_� | _'ڊ��/shs�u/gW���jn�t!�D�����)i8&
�똁+F�j2W��L4i8.�k眆�gf�7/�So�k}tԸvq��N�N�>�	k�,y�Ýxb���]��b�ǡz��qE�(]v���,ސ+�.# ��;d���9˺�
v���޶����W�����y�5\3h�tCŶn��^0d\ʱ�Z�2zH�O�z@rͦR�S�0�47��԰�xs	����썴��V�� ��n����g�&�C�kNxֵ s�=)�'^H��1Jmi��+���ڍ��18�����71�(iMw��'=��h?��ǚ�+CG����n�xl��_��؏XB��
=%�V�P�֧�?�~5���G䍷��c0�S�s�r��|2I�h�O/f�懞�jrЅ�6P��s��P�E���٬����EE�?�	��e�!A&����!��9��%/8�D���X�cө��w�qD�cF݈#_!kE��!'�s�+\�7E4]R��$�K����g�`�8!Չ�e�9b��+���ϟ�S�+��\�9�4�
x��G����nG��s�K,��A����E��� ^v�مR[��C���*6t?ow�ƚ��eƝ~���`�1	�rh�#!aĐ������$�P�Ŕ��(sT-1]-��2������[��<d�u0譲��'�����"�$��B��#���W����j���M\jMs|'r�e�M�5R��W3�4�{��Ɠ��.�ЫX���,v�jv�br�ڐ9�K�ʯ���/���a߫f�\��42nTt?�)��{��̦�;/�ξ��=v8l�1�D���A�U�~!\���*U/L���	�U��W"�b��H ����eYV����W����{W@m�U�_	p�o�\�;,y�O�%}\�FN cR:�Ծ��?�9V�ʓ�WST�:�o9�BwQ J4s���C�[��ϥ� �R���y���  ��w�n�=��\<L���Rq�r�v�i�zǉ%��)�!��,Hߒc'�{�<J/!F�2�����6�2
�Z�����_]pK���RX��bI�տ��"%���6��)b-�^8L"Fi��ʙ/o|�M�
~p�UQ�N�Z�l�V9�>�c6�Bj�)�|;�΢>*Oe|�z��I���.A_�v�j.%�"d$	�<�~`�OU�&L�'�>��郋ld[r��	��2�/��_ǲ���F�^S+?�5��d�5�=�:
�t��|�"+_�-0�,sO����=h���.\�9)|.�q4[����L���[���k=��mٙ��hqǗ6�4Ē�M���jA�����4�3�)97�����_O�d��-Mcc/���6�ro�/�r��xNU�j�>���2��Z4}̵�;< 
�[�=,a�!6G��L$e�e�n1U2o �(Җ8�J|c�J6��<����K��W5NsJer�<�h�����?��v[����$��F�a�
��R�R ��� [B��`�,F����8R�ZH����k�x���oҘ8��Ը9:�F񿃎�17ұS�?Ir��,r�'�ѷI8a��.uY�@q�r���o��QJA���������U��ҳ��Qy�m���3�m���FS@�	<P�jj�4 �u�.�%5�t�}�>��ɬ@�D{;>1��q�D��BC(
1F��u��"&sb�y|X���⍕�,4���vq ���rNG���7���<�|'i��3�Z���gco����ZV�N*t�^�Kq������9��?R�f�@.�ڿ~���MH!?�R��v}�&���5+�cCq���͟��ցe��:9/����	nX8��l�;�ukh�7�F�2�Jb�:�f�=�Vx��w�,069;�r'0R����������(�����O���`�x�LRY(1M!�I�]�U�вo�{N����7
_	�8���о;�qM��cԢ55�ʠ������{�(�����U��?�$��2�f���֗���8k����_�i����z��>=i�&I7�Q=��s�����L�w�)Gy*B0��ɒ���=yrz�B�_a
M��A�X�&Al�N��A���'�&��
�f��"z{[j*�f�J"�rU�#���Ɠ�����uwD�5�����:�؏R,N�i�5�Է��3�2%�E�͡�� "!��4�c�t��W�0��Dw�Z����.r���2U�6����]��e̫7�ߣ|�悁��y��YT�.�]�[�x�&ˠp�O,;O��Ix���"vJ0f�qu�8I��V��6�*gX:��y����X��z�p'�v���U����%C���u��h�dX�#}���^���t��E?�h]
&�s	�Tm�Q�[�F)��З�R�����d�E�	���^�gfNS���nݓ���5���oi���I�O\pm'�1R\���bD�E}�H'0��"~1�x}�6^z�-�-�`K|��~�*؅�>��Z�� q��j["�X�	�G_�e�O4�9-��o�p��!�ej����i�ܯE!~em�H��'|��Ԟ�������
�S��ۇ���yn�@L_'�YO@%[���X���o��x���>��qe��!e v �P�	�1�.m�D�m]��b��P� ���L(�HzZDo��� {a��rlfĂ�7���5o���-�t2��,Qkz�S�yJ�?p������`�de���.�z�����CNV�����I[S�e]4������EC
�rK�P�C3� {ċs6-u�s��PE����o+�q��D u�)A�R�<_B���W��j�d��2p	�a{�hy���;�
�����Qzžf��@T>ɺ
��Z>�B��N	�T잍�1��0�"�S�q#�#Q��3�Y����� 8Nk�')�%�'I2P�i���y��pq���g\б�5�[��T�#W�+լK3H%�z₡A��'ː�G!z>�u^���[L{�X�y�w�1`��?�(�����}������������Ny�<��Vk�ū��Ĥ�Q'�	ə������"3�ܳq�di����ِ��tp�&�m�ѝ�U &���0,�3�݌���أ��@�$�6��F�^[R��B4t�6����R�$���+�G���W]R���d�����U����N;Tܞá-�E��^�jG5���ݼ��o���[�
�[��� T�s�[[}��`�p���6�������s�~��Wv�$}��i�Fz.�)O�Z~�P�f��J4�d��'SB��=J��"9����w+�Jb�b{������z�p M���(�Ex;I��w�G�u���o���6=�g��Ƒ\�:��y*,A{o��E���aO�s�"�JV��{�s���,�����"��dw���OL�]��C5Ha���c@t	�W�E);�(��W�f�M�ݬ�#�O�ǆ٩Ah	�VK�S�#��9���9�`���h�S�}>�ʷ��?v_s�{W�F�9;<ksA]W����p�?�=�$K��%�F��:��p�{\t3��ڂ]$\�C�������$��;w�6����C�+Vp�E�T���;Z46EϯI>l�!�Cb��t^�`�]��At��5� ��A 1 y�VlU�ݍ"���͆�ER|܏"Aq^Tz����D$����iڧ!��<�(����m���>��
��]��Q�Ze�����d��I��Fc-V_7�y�V���ʕ�c�$)����z���.%b��E��!���_õ��N�m�w�[���Ӣ���:�;��|/����jF���mkWٓU8��Ŧq���m�K�?���-�N����=�1z��7�L�(@�WPb�[2��^���.c0�
�4TЋS.�m���N�_�T+�'�O��T�7��<3;�X��p�?;�t�Ƴt5�-��d�qw5|��|�g���+�ipL3L�����lG�oBSV%6E�	4��۟7���t�����u��ozf�4�
CV�t{RI��V2$��:��~n�p�x�����9�[끐r��WM�re33�f�7AOD���^�㙘�����3�YGphO�[��"%�q�Al��f!	h����
/3j_��&��et�!���+$�r3�D��7��v��c��cZ>�S (���PU�����$.�W[c�r\�<
�nm���>�׉ 's�&��:X`��௘��l���sf�[v��S�fޱ�̬Z
�&�"��VV�`�M��o�}D~ڥ�f�����$��_�ܗ�[�ΟE��v�=f+v�>��[��c���7|�x�m���G�|@e���"v��.�#f���w���U�F!S�0;7����#�۩�<��"j��[�@VV��K2^����_��0�R͆O���E����e�O!�8��+���eO�o3V �{�n�Q<�}	�������#��9c
?����k��+Lp�tq���V��N<_qGlɦ�#|�%S��<Iaiu0~&�/��ʆR������ϘMY���������SbR!�#�����w�8�o<F�K��hH�����*��ޟ�|O��1�� �M�1����������-�Dx��UNx�`�S�:�8æ��`m�KR:@ș����+;�5(W/Wq���Μ�b.�+�����=����[�����~��Ch,ق�,\�2�[��JC���<Gz�N�y�dd��hr(C�����B��]��~㈜jS�u�_nU��a� �og�Z{���Hqj���w|y�,p�Bd�`�=*T���5�7�!�~���r61��5;�L�q���R;�S$�h�a@m�y�-��*l�67��F.�/m��w��c����s�ڴ��nй>���_��]pr�Ԓ���00���D��C7�H�)n����YiS�]}
�B��6Mb����as��i�}������St	�����(�ٻ�ŝ{����ͣ��e��[�-"�YS��1�.戩��T�l�>�j<�PHZB�Pu����<�|��Gܿ��c&	 �J�#��"
X�dl���owL��-%�eGɗ�$G��S*�I�r���f�J���a�9L8,��2uAԥ�����&�]o��j��9
PJAn/,��~�']�3VH���hE����y0Pٯ?�_��#��G1E��0?r:�B�P������EM�
��T�M^m(w��(��pç��
��W�a)F����ێ.Y �=�n����/�?읨�.�6��2k�۬�x�@���a�X\��Vܪ�Ɏ�_.��(�\�g����<���>7���\��M5�,Ai�����҃��0�P�ۭ�Gīo�b7�v�:�a����0��b����o�1�l���穼����q���x�J���
p��%��I��dA_ã�T����Z_�0-��k���۰<҂
ƻ+������2��ha�B*�(��&�-�(y�P/���C�*��èZ��E�Ϛ<b�V�%���dE���5 Bo�N��S�kPE=Y���▭��Q�'�4��ڋ�Cb6*�Gx�x�@H��i�\it��3��I���W�_�� 0UMו�g��n��-&�3ˏ�ڍ

��@����;����{�o�6�H�B�XNZ�0�ځ2��gW�~"���g�{�]ִc��.�Rc
B&�<�{o:$4{%�]VpY� �W�Ƀ4P��À��?�O[Al��L�*��hj��"�����5M;�>�^��l����6���%�Z+���$~�'N+*�qҥZ�O�}#�����c��3M�_[#8	>V�>k�i��j
�>YA&����d ?�3x�*������*Y;�
=�0Σ��ILAQ��U�L��*"��|�����q�GF�B5�'���`���o>Q�p'�l��J���-���z+?�Y��#co�5KN�(7v������I��><;�(��Y���M�j��l�� FC���̌�_"��+�`��P�'9��]��Į�^K�!�2n��郚5�دp�s?z\�'/AЫ&�_s�)�o��m��S���	B���}��g��;���I���e9��-kx0{G����X{m4����	)��j�I㻸N�|��K�2rF���29���w2%�����Y��Y\�Gc���=�f�x�c�X�X|�ҏ�����M�>��O����p> ;�h�Xj�]޲�%!-��L)g?�㷆Zi��0<�:m=�FZt��U�;HK�$~`���vdLu��C��yɓ��C/�Dh�<��el���Qn~.����G�S��}`hE;�"��}�X�Zt8>y9�:j�
��bb������b�4K"��^8��$��7~ΞJRUe�li�l
i�r�/>L���:?�(�#���*�t��ܠ�2�l�0>u�vf)k���qhp������t9��b��|^���`�^+���ؕ���`�q=mF��\���(c��Ճz��{S.i�m�=*MS'��ݨ�:�����l��Y�����Tg��f�?`�~��L����l��r���59D��L�����h<�0�L�'�ٍ�=
��3�w {P�gt�H�[�:����9X�SA��_֭��Y�E�ǡ��Z(Č{��j��+1�=�A�g��cE���orb�G��ΰ)!�g ȯ3���<�ؗh���c��- q�M��jϑ�5)��Y%;f0�l&�=g��	�	���?S�����p�!�]�FM�Z���f��S�U[a6���.腟I�Q�uA�"�/'��'�Kc$$Bƚ�v�yc�Za:1����^�+�����_�k��:�4*:�p��� лS�#����o��(��2���d���4>�M� ���G���]�Is�����%���ҩ��*�5���Đ�T9S�r(K�&*���SI���y�#��Fu21"�e	TGe��gNS��.�#'ǫ�zI��?+�E�`8��_ �������6Y (�7� �s���.�-��Iz�L��6W�B���%�����} c.P�7z�5H�\��	��	�^`7=�N�ư,B2i��r_/gf+�������+@�x��!�.�s���#6W(7�bq��n��lz�DOk/	�6�ܿN\`��?J��[�s:��D�g�'�X)[��?ދd�iF�������H��ٗ��a3���j."c�+�M���ߌ�WB����*�~Y�v��T>;A�R�և��"d�)
M��*N+]ݏ�b�s����t�H#�A�
�����ｺ����6Z���I��A�;�ܦB��/y_
���h=��f�»�<x;1A�d?�h�X���e�&��r��x#GO״�g����M5�������.ʉΥ������<ᴒ��P�2zl�ЏN�T�2�+�!�&�1�A`}D�t�HF�;2��hL�&�.�ﱪ��h��|g/��ݮ_�9ނ���mѡ�������P�R�p�<~�?g5�0,�:& 
w��`�Zu�"��T���X&?�K��ߍ�f���;�ӋC�uH�.Ԧv�Ń�Ƃ~1ޭ=�bO�e��v�+k�]��X����C�~>�Z�/B�)��~��H���=�A����efz��	e�~j��8���:�,g�߲	�1(ZEՇ��ӹ�̖������OL�@rkS��5�F�6��BE��I�H�kBA=JoV_�yx�O�+�I!y�}��M�i�]p��;��؏�ͬ
��K�tful�2��V��X�$yX�Mhu�i���%)Y=�^]�oDµ�
y��wB�C�����,�s^d&vu5�
r��p��Νʂ#�b�ZR���6C�m����w�z��ME%<�6�θi�(Y�E2�z���1�f8T=��ȷ<W�B�G���H���n�֚��Ba���O�k��EZR��%�P�s�x�6����Y���bݻg
��t���1���-N4�OK>��}�ޭ�Ùz�/�m�oH���d����=�t
*����u�C\ �B���?����s+�����T?�H�<%��d���eya�j�.�����à��Oz������}��"�]��;�i	�AAM�πk�Oin[7�['�Z�6k}|�j5�F3��h��U���34=q��MpD�����[���b��NM9a�-�i(��{��0Us���� 9U&+Ox?����_r��vj�VLb�����Vg-	�u�Ӷ�s��c�ƿ0m❞3���8ֹ}�~t��e���c��Dqֿ��T�h��z99~,�'����ͬ��}=����Px�*̊��m?A�C�Yv'���%ܭ�9{SǼ�� �����nT�7^�%���d�0��L�Vz�b�18��^�7��?L�&�������(�8T�`��ICTo��g�_��F��g?�lwy�o�Z4COV����!�o��$��)�`����W��������i�$�ަ������˥g�3�������[z�\�p
���J[��Cp�7fQ�ݐ��;@����[%(p��Y��M:�;����y��h��~_� ���Q��6�o���]/%��W ��zV�2��t�ڹ�ɑQ�s4�3!Q�l}4{�"��7_#J0E�:��UG9��O5qk�$1.j�`����#�N9�G$���WıӖk���J�4�k�<O�w,�9$P�=���i,x�Ii76����p��������d)�H=��X�Q����\f�D�ٕ��X�Xpa�pi�y�3���_!�:������������r�$��Y[;�g�܍%�`=&�FD4P]����S9�>p_���C��*�-XzF����ŭ�;����h��w�֋.����j�'��{ �l��q�v� �<9d�A\�����Z�$�}#�,36��4�C+R+f^պ�(�xK�T��� S{�ڝ𦠜{6|���T��h����=D��D�D�.�#��Q^��g��ݴ��Z���<sf�)㧆7$S���!�V�'^���gm��Ǣ�_�L��5�Z7Oy���f���Ն/��6!tk(��F��A��q#�R{G�9~�<Rl[%�B�x����$�K���'�n�Q�\w��lOC�A�F��<;n�I�{���K�4���ju�Y�<?J���y�-��>�H�&9���&�l3bwx�x0�YpY�B8�jfD�\*����_�"~Z)Y��F[�?�b�|�}i��k��л��j �0���M�~�>q�^F�(��䨤�wj�
>HsH�K�s��:���MI�����6����R�0'Đٗ|��xb�.�K悷Q��Ր�Z�[���[�MT�H�s��s8,n����b}�:pb�~}���s��l!�X���k���O��G�Z�b��C'�-�)��x}z���k����_�g����T��~	��m��75+0��ǳټEM��a�{[��T�u�!�i�]��T�u㐐D���f띛>!�T-[���G();ce���1�$��$C7ۤ��}�0��y���dLz��_����G�F����<)���V�(� �����0(��"�� G��)v�H�K⯉���76�yS"�5�(������7�V��b+QZ��� }��/��hV�k�[NN��X(6vl3��q�
ْo���hCKZN�`���_]"]��'s6
��z4���o+�s�$�45]�!�v�$|eȩ�ԉ[��b>���q[|��eNW���^ /�Ş��"�/�c�GQ@zUBCr!�0z0%�*6�@��>��`�;�'���J-�1�"�4)��G���0᳛�f�
��{�dq�r!����#J�mG���P�R{A�PZa�=�;O�c-�0dB�[J޹ Q ��d\4�B�������i�y��LLĬ�99�L i�	���ռoQ�P���ԧ�GCQ���I�7�U������O�i"����;C�m+6���UcY���u��n�I����L\���k@ɐ�2;��M��]mXԱ��΍iU�9ɴ5J|6��!�����L��4<]C�ٴ�`�^��kU�,P��5#��1�7��L7�A�.�E>�԰aYq
jQ��o�	Y$+�q��q���o��u�s���cH�IÐ*�p��Ş�M�da`5U��vR�����"�T�&~���-�m�SJ��&�����cw?���1�p��B���o���$R�|�Pe��.^>,oR�p�����u��!߹��Y2�3p1F�BKb.��W��ø�}�Oɹ���T���@�Mf��iG9���h�?�ѽX���5p�A��u�6�o�a1�ߡE�0=�>C}�������%5��߿��آ�s���(<�1��^"I��K��FU?Њ_�f~��8ʟ4u��Mӄ;��݃�5�?[��0��_�B�ç��qC�v�zKh�r�7��$Q���4��mC~��$�j�[���Ľ�?5h����)�F�Q*�/ʐb*���=h
�E3�����Q�B�˯?s6f�SP
AY���f�C�(sW���N��K�VtN3�̚4�F��IA���&@��!�xBk�!���	��l֐I(�R����7Q���z����`�K�m��0�w��a�U.�)����{���oJ���C��$%����g��+4H��Z�⦏Fčsz�Cq����E����{38:�]�����gW��\����]"�����ĉάL�L�.��:�н��q�iWB����
yy�$'\5���q�ܿ<P�� &�*��g֮��7���̪sڶ�{<��h|��L�}
,�uލB@�p�@�!����b8^�Y��2��8M�g�J� ���k�a�4D*3���_^N�:�0�!;�&=���[����V��:�,�>��q'l�m��B$�r?(�SL�����:,E��T|�&�Kb���f�4��4�����I���-Ȼ�OAnrB��`/ƫ����}�æY��ذ"��N
TH�p
Uc���8��n'< �-It�g�}�BC�G��J�aT�e�)����`��%�
��[ʮ�K��Ч��\+|���w�����<�X(��P���;�CB�?t���&��-�M8�o�?�YڀB�-V�f���������gņ�9�p�Z;�;��KڞF�w}�ce�)�ӓ�߽3��w��f��4V���������U܍u�j$ffc'r��ޫo����<;��'�_��b�-7:ɘ�)$�B��
��mx'�![�x|�/>׭~������T{ς���Y���
'��9�^^�x�q�6��n1�����ٚKv^u�	b�0]��`@)�}:���w�f#$֑4"8m�N���<)��(�_�0X�����Jz��g
��O�s
7�gS��&��]_E��ك�l�`#�#lk/{��[g�S�б{B�����e�1�%Oq"?p���Ô���@�Z)6��q~X%��`z��������ځ�o8MՀ�c������Nr�d��ʅ�Do�&���%��T�k��+�u�dF�[_zqs��O������zP����n��a���"��C�G�I���֐^�G��;D��?L��!�m_Gؼ�R$�4�1�s]�|�ь<B@����&8���7���.�Q���AP'^��8�'�7���R:�0��׳�B.�v�	ㅐ6�TX�6\�j�^�Q��B�1l�ܠ�AT{��H}{�l:����i�D�k���V��ic#�ߛE�� �#ܞ@�H��k�;�/�q��˅?��?<�V�pv۱&Kl�JP���f~��_a���h