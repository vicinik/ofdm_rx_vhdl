��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒����U�Y��7g�(*���K�߹4�"�T�P
ʺ�:�W�7�΄gm�e��x�Z�>灓�0y+�j���T�-RP$0��"�d�j�X1:X+խ�%<U�K琒��81�uK�����(��6�����vM�:�
a��"�  �@X�a�ӃYb�84D�`O�l��2��9��Z҉�$nd���5���%|ħ�ybM�>R�;�lN�%�~�w��d-�C�$r��	"��fK�k��qv��T���O˨�����`N�W�:�1?�6mڕ��=�ƣ�m0��-�p�STA����|-�I��c�2/T���:Ktw�$*�b1�8���k�?��+�D��<�)���b�<�4�"\����e�E)�h*��	��V`�%��ɰً����:��9!|��w�\�D������{:�=��K�%��r�WIR��x�<p���lTZ��6wWGb.2b�|8�LU�f��J�#�7S�I��C�(*�4f����t~̰x�c �r�W;hw��*iI�̉�E�8 ��1���6�d�.����@^8�L��b�`�y����[/�ļ
2�`+l�l4ʠ]j�qVC`�O���ѯ�{��7��ŔEsP�"�Z���?�M�Y�o75<#���Ub�����P���[C5��o���9�<
C��s^���ȶ�В��SM�6#�u`?�p���l����h�g}�;�������ӥ�k�']��y���8-�g�n�� Y�o�{�. į��+��}=�Ն������>�o����x-�m8Ņπ�ɫ�}O�M���$�N��;��:Y����Qkܕ(�T�/�Y�N�,�J�o��i�\��$`�IH�S'��'�ѼG���5	�R���z=��$��$͒3�b`}�;��$�\�}a����h�3LiMA���'1�F�M��W�u�eo�]�s�l�� P�8w��g������O�ڏ�s�Gm���g�l�F�hu-**��o,��Ħ6m�����_&���Hf[�1U���I�!��Rm+K�` J!5�����;���*�-�ԉ��н5�3����p�]��%��r�Ea���I�������I��F�Ž�̞Q�\/a��7�.�A����?�s�ʖ�h��ΐ۳;x���2A�i����aS�U@gb��o1�/�B����	c���{>g�-7�=��Sϣ^�E���x�p�)șA��	�x� �,&�EGx���/ֆ�-?��)���?���;��q��]i(+�����h�R�BYu_]�()q
����	�pCi��������V���
����V4T���ֿZ�&�jq 3�O�Y��5�xF.u36-�okv�< D��@�ϑs���L���ᅗ��b����MW��<��-��4���4�+����W7e����w 倰�#=qU'{֝{;����*[J�q̹��9�)�&w�{�1��3v�E�7_j�X�;	Y>zR�zyY��~^|gx+�|3���x-��	�;W���䇆�D!�b�o��]�7�͉��k���n�(���G*:��������ۿ>��-+�3�k(1SN��wU}����%���ދղ��������
���IAu*�;)ܢ�,C�(�����9�����ռ]1.D��QR8A��|ʾ!i����6���4:c�k$@����`r��u��i1�󞩾��+d|~w�q�6�^�0Q��]2S©J���s���/H_R�9£W�������*a*]j{1���]!���{�	�>���%�P���&{ua8N~VO�f�=9�D'�k��ω�6��N�d��Z�k��-H&�f �� ;�ƹd�e���Ġ�z��G�>6/ɽ� 	mඕ�9 bq VB�fE���3�,�W�~��@��;�0Q�	��KG2��&��-���w�����q�1�b�{{+�n�w�ʩX��WtG�h�)3�%�B���T���� wRy^�J�6)�o���ךw�x/4�HB�i����9�B����z�R��e��u�܂h��*��}e��9���#��*b�	#$���#jK��B�;62i���d�;��� �`��|S|WN@y�5�ʥ�k��^w�~�{�j4b%�@pD1�8jVP$��Ś���M@{�:����ܡb�A�^; ����vݲ��d���G"��a[����;C����Z�xKQ����uˎ�dpi���z8����@�K��s������릫��&��3Qꞽ�Z=�TK���Ӗ\��Og�L|�0E`&0`B��쩼�,�;���?k������k�
t�B1�.�ъ�%D�EAwU�������3M�aEx麟��XC�Jt�]"[��:`���e��,̒3�=��`� ��ئ���C'Ǔ��D�w
V�q���/��?Lh|EW���B@��n=T2+�]1��UB��2�-�-Lh���J�$��_k(I��2p�0YB�pV5�3I��9�V�����c������th��R�#[��G�;\���_���~�������7 �����"^6L�g%A�:��֘���A��R2ӳ_��Է@������"�lFy���q��uv8���[v�	��+�u7�2^HrCr�UG���۳��1F?�~��dfC�h�3S��ȟW)@����֒t-̗���29V7�N�!U�t��{T&�O�d����.��Ul^z�
��m�ek��� �b��n���ʙ汾|kq��l�7N���q1�V��;禹�%�ϩL/����bqv�C�Y��+���:eM�D.��5�O�@|d�2ʺ*-��a��SU;���P��8U�J���h��-�+v��,�:&E�nص 7'�_���6�@�$�É;�o��G�Ql������gG���Q;/LrO��������̸��9����qG�ݢ/2pP����(�^�^֬m�?��x������M�Xe�o��TF����	3q	�2q,H8�`^�|#q���g��ٳhh���ш3�81�̪_"�����E�TqY���J��z�p�(lqO43�d���Z2�|Il�^�b_�$;n�'�L���[a&��L�)!�R%)Ud��yv�������F���&�P�POU�[�D1[J&&Tp����,�O��S��^'���6��43��s��uHV�/�΋�ˋ��gj_
�B�
I፲���K[ݾn��%ҳlؼ�0��1��aj}�l�K��e��u� w���"��M��yŎ�v����CȚMA� ��a�"�����崤8�>�" ��:"��Z�h���dxC����� n����CN��N$q�b��v��	
�84ώ��1se Ւ�7��X����H���꧗�}cտW@Y
g*'w, g�4=sgl�F�Q��̨ !�"�y�����K	�����NM�@3���1iy#d��Xع���g$�A��ѡǫ�tL1\�[�Q����Zk Z�=/���!b���Q����%�ɠ���跂:f�RjP�oO��TPgY��}�y�S�5>��џ�ܴq}�"kd�Q�O��&����ew���}�A�2إR-�}v�ԧ�a?̔?�/�>����I���:z���:T�	8h�D�߀2(Z)���盢�Ẁ��5��M�Ny�X\bލ}�&����!�|d����J4^��ط��S���wL`^�J��x%*r�f��R�\��a���Q����դ*6~�فo�Fq�ڛr��yֿ�9��TX���X!���q0'�5�7 !�1�sX�@�2���bz��(B����j�W�0נa����C�	������g ��k����a�D
�v��F\5��8@tb{A((��
�,x��G�.<�~8������BF�p5Ɠ�c)n�6�[ň�m{�!��/��GL�Q������|v�D���cL��/8+�W7U�9���Q�͂�c��v׋1�FO=k��I�7���H�7�?B��
�ϱ�IV���S�.����d  �����9D�~U3����bA�eM��y�V�d��?w�����&�G��G�xJEy��[PN����J�wӶqFV�c˵�0��Q\:ϫZ2�ލ<x�@�и/�ō.�`u�)���8j]��Wp<��(����)�60\0W�6 �"�D�z!V���M�a8���&��X ����������?ݫI��3Jn)gP�F�ߵ�^ѺᣋC��E���lU�C�}eM��Y�r�1�G�ID��d^�y����u������/�)��#U�L��_+�C�'!_�l�UNW����ҳ���p���A�-uπp8�#X@���Q��d �k�`���+HW�":�2e��Ny�Yⷪ��\�p�SӘ5B[�
"�I�{5���AI���(c�h���p�(�Ka���jWvg�i���m-o(�۵��m�2�(���9%����}���F"��s��K�B�5Rx�?�R��ߪyD���#�uQ'�������Yy��!� ��,�ێԧ2 *˂/���d?(��`�3�w�k��ܛZ����24�����)u��$w�e�+h+9�gi���uP�'�-�)��rS ��'K|:Ţ�u�޼������'�6�@�5I0ym>�_>GǪ��,���<��%�"�`���v5K��i�d��m���$�B�<S��Ie�ޏ_~5j��P�	��]NN��8��h}ɵ��1�,�v	���1��&�|�a|�ҌW"w����@��lۍe�����e6�S4X"ٺ�Ƿ��5��\#��w!X-����B��M�MK����VO٘�����[�^�C�C	�ɭ����=Դ�s�_��íq��r��[|�� ��Wx��1�Z�OK���S�~k�<[��n<�ۻޝ*�@=U�@����	MgD1@E��*���./�p�� nY�p���f靱�����՚�t�N�ZP�2SF �������2��L�E�aG��0~���x+��p@�]<mR9_��K�3�,&y���rU�މ��"
6��W�.Nפf���O��3�9�.���P�X�c��Np��aK��w��VK>[{#��XK����qh���a}��j�u64Ԩ'ϴ��������9f�H�b���Y�^՝:>$��dnH���dq��S�sʶ]��B�kC��js�Ъ~��&�Ն&7zJ%_��� 2�~��vh�[�Q�XG�����Yd��r�����#�ݞ�lV������6
=gN,��m��#��o� ~٩�5J�<p�����[ȫ���:(�y\,��j0F:1��K�]��L�ni�ҝ
r����2�Z�b�h溛٠auS���=��4ow�p�a��m�'�P��q�T{�}��,0��R��?	"W��J��dk3?������^y�H[�	@/jsU��$͔��.�x}#[v�)%q�4����^stB�A����#�P�p��j���Y�+��z³C�ₐ+���B
}�(8�y��܅г���i��{2�D����t:�� #�7�G�7o�F���S�L��ӛk���}�R\�i緀��0�v�Uڌ\�eၤoj�)�Հ�,���4(	t���|�<?l�ڗ���ŷ8h�\�S0:���{�ўl��wl����rr��J���l���4R�ף���o�n�\X�U Y0� C�^?ͦg����y�V�+�V���<m��+���WV�J�8fCQ}��^s�1(�*�@`U�����]"�����uµ��cð�N���-ðrZ�h�R��C}"F��g���~v�f���	.hâ6�B�`B/��Dͯ���/������:���>�,F�I1�����;]�*�p�l�ߏ��y��Ѕ��� &'7]��9A�^�Ң��5���h5Yl��_�2� ��D������7�%=��C�L T�AE]��������%�Xn�������_�|A�tl6�w��.������4�8�IA�vg��uU~�x��4*���x'����"�i���ۦ�q^oZ����(�
3�̅�}���X���Ң��
=Z�̰�@~��{83^[x�%�2ިV��ƣ,�(�_I �ߣ��Qeu��[�B������j�����?e��������9*i2�*�4�?'_[(��d�j)�D&D2H?(�u[�N�R쯃(��9{�>�X4h=L����Ю\ǲ�����f�����sH�K�n�X�:�d^�a/s�p��w����+ ͦ�u���&��B+*�a�h��V0 %T��7���ŋ� Ϩ�-���B�2����?bb�vE^��+����Ö(zK�x˜5x$�hM�𮙳�<��h�]8�YËd��[��t�~�o�@�n�BDG;7Y�g�&�,s���k�%��LO�'z��D���H؝�w0[��n��4� ���/����_@�%Ϫ����(�KV���ZՈ�Gb�,�S\yy�NDK��Q%c��,r��e�ִ����`���f͝}�1�
I���hmX�]<a��9��K<�nh��w�kՊ����?ڮ�ۑ�sP��)��P�_18톃���k��,��jG�8�}T�IԙUJ�Z!�`�a)_KOF�ʒ�- Nޮ~�T���i�Fw�����U�)Jhe�NǛP��HQ�O^n�"��'-�GH؈�w���"�JT�[��Һ�6���t�f$�he��<�7@ D����d�W��=��QE���SqߤS�&H
��,�ĮA�	k#M�g8��!�(�^p�)H�5q�����,�fAfݰ���S��ɑݱ����O�]�������M}7;�RH��;_������и&+�����J�®cO�T��q2��gl��Q�������e���F�r;�1��3�]y:�� # � �/�88��%�H(I�Km��^:�,\3�@ ܀�îHwzR)�Ck��m`WH�3maxw��"��E���h*V�k|a��+�&T����ߑ�oN��?Wz���j��qV�Fv��,�laa��1JkԤ�L��3�����-�5?��q��X]��>�"oG�C\Mk_��w�k'|�Yqu��W�̎<(+�mf�����|����h?�Eǿȯ� �A�0f�h�cN����3�?�)�r������~���T,�ؾU��\7�#�Z5�P��m��4���K��X��17��ZV��\�u����p�� �����X���I�?>�L��TP�od�3�5�E�f���o�.:�0Ԋ�7��x��JY=�*����0oD|��A|j��ql��h���hK�ז�_d�?�CV9B�"��|+�f�_�TP�s����R�x��ɔ�6F2�f+���G�#�n%5e��X#�/��=�#a�����H�8�P� �o�22Y�?��QM�Iyڈ!أ��=��,�7���:J�L����Ҥ����nZ�6�T{��uH;��69]O�,0�9��阰#��1��U�ߜ%B��Z�
��5�����Y�ر�O�d� \ߛ�!�����E6�7��Rok<04 ��H�;}��W�$��A-���A�߹��'��E�v�4,�H� ��?]��ƇDx�����K3�"Յ
���Y,�v�Qe� �oW��&�Q|�,��ٳ�趵U��º �L��'���aj��"Yvxe�\���2mnBS�c�b��v��_��v�~�)�܆�!jQ�$3�T���̬td� Y<�/��m�4Α$���'Ǧ���!�4 �_�4rؗ!v20Q�g�����[����3͹��H�+IW�*����U���Jq���z��"~Ə�L��T��o�gOyh]O�.�?P��̚����M}�mO����-��$�����Es-,ݣ�c�/�9X=5��᧫=��c/p�&R��l)|�V����~�\�N����B>�]b�\+�{������ky%��J��^��+L���A���V�`��PL��Z�>Zҫ�5�ӸҰ�9<5�e<(oS7u{{�W�n���W}��)\m$�Wl"%r���K�M_n�@3��u-ŝC�鼽/�MB�g�A���,os-ڼ�yu�ƫ���q��Uf���^K���4�݈�J����tu6��S#y�'���u�ʟ���"`&��������,��]��d�[9#�R�ؐ���H��&�>R�B�应:�^�y��fB�l-H��/�VsFQh���(��¦�BL���q���=A��]6mN6���P���H%�� �Nc�T=�����-�ϊ����`n@�����3X3��;�I|�S.t$�k\�0�	4O�_��s$%��ň �t������V�9`�d
��x�"TN3L}2q��qHMQbC���Z�p�C�����!v�r�#�bi�tf�̰��UPK����9�O'l,�!D�\�[ө��7Rf�}u���g0qj@+7�q�m����zF^J �ܽ=�IB��5Ϫ�阹v�Hՠv�C�w��ĥ�Z��p�c��>�U��;Я��3:ܰy��(��)O�=.-f̔V�=R~"����۰#Ǻ�r|m �8�%e!��7�hݚ7T1������+.92Q���Ȕ�����._s� ���~��Bt��۳��ы�Z�jN�d�����$T�%��Y��*��@�?��`�B�^���}�Av�"݈��W�9�B+-�o-�4�S:Ft
��lY�dvW����ŷu�~���{y�z�ht_�20�c�h�[΅��!�,�F����P�R�6��-B���K�4�U���ȯ����������̖�,
}�"�+��vnR�C�a�>�_J���cV�R:��o�h;����d�o'��`����Y�=����[�v�<M���|��'�[�;�r^ΫC��I���&h	�_^��I��x��535�P����On�}Kx�C'�@Ǹ�,k�_i�t�X%�f���!���	G:�;�jh�O�k�UN��Eȓ3F�#����-�!�k�<"A��>�\���hI3�O�K��Pu ���=�ʜ�
-ן*�dҔKK���)	�Fx��S-m�(0A��R�g����,����y���Q�z)W9�
m�@�E���e���a�]�.28D�fU+�ri��C'�bDx]ٜ3A���J�NlNx\�j���R_�����x�e�����4�dD����r��s����[E�>��k������l	7���=�~���8Y�%#���ĳ��W�-��24����*������&�X���zwV�r�|�yv����v��� ��ֵ��b㱌�s-�ߦ�(i:�Kt_-Qy$�sf�
h쮔�ؼ0)%��i��u���ڏ϶G�ex����%�%��7����t���	z<�a���bN�I��vh�,�ȅa�W���V�.�zv�b�&?#��T��\��������(�YX*�f%=2��h��?���!�
�0#����"�و��͍�(���۠PgʡMn[��U�ēv[&98c ���"�$<M���Kh��MS4�'�1�ѡ���z�@�v{�a���!�n˳�Q2?~��}�h��"R[�ZV���q�����F��##�z-�VT�U:���q+�B���.�_���p7�05r˙_^��[.V��B�_�~�����Ϲ7�[��]��^��P~�G��-�xo ��;b�F�2�S�A��`DO��dk3��-�#ȤJ	[r3?�+Kn�T�Hۀ�3c/�I�x��K�
�|@�/�Қ���+�]���B�h��b�Eɘ:>�r�U����&
AzYS����kPw	�9)���m�����}W��l��gr�7�x} 7N<�Lޥ�٭�=�a75������C4�Ȝ��n�Y;M�X�N�%��]�����C�h�܂�h��q-'bZ�c�g����	���ʶXna6;�8�����KL���!*���x�7��yĜ:ҿ��@L��m�۬���'[y�3���.�J�G�X�C:.�t�I�G�&|�7�8���h·2��8�Y]ܒ4����r6�^���&6�%����"�i��d�����Y<�ԁɷ�th��P��V�2P�60٫�!�e�_nl橹��^����d�Go)b�p��"���dZ��O�<���nq�8�59�S|��f����4Q�#Z��F#[���vnTUd�)z���5�w�N���@|10
�(drۂǮ�:���ɪgH�i�;8��7�z�QhS\Tr�ZV�x��FK.گ��D�����W�����Կ>�:���o��q�o�θm=+�����@d�<���[9���x,�I�>�/y*Á��+i��l�2'��Rxm�P�!�Q��ά�n��������¯b-[�c~ţL�U�;%cO�I��h	��R��.�.�o!z�����ހ;���`,���	�!�i �*�7�8*�.&�°����h
�^��Je�x��_"�!4�\Ny�H�{[	���n*�i(bz�\4Ӝ�L������/�����Ud5Y@������7�u��<��;��[���k���4f�\�w6���i��t��^������^60����~��
�%��1��ґ=k>K7(�(������6�(sa�C���(��A�N7�mh�(
�gi^�/���TV��r�v\�)���!���L�^���0Z$p9�� ������|�_�0�I�N/��nW,]�J:�c�68��l�Q�;$i-�ǌ:�{�����_��v��q^k8H/�د�ˋ�W�+yZV�6�5��\��D�OՀ]�ծ@�Ic��O�A��`d�x�U�i\�]��4&M���rf0D�}u4v�!!�6]����RWĺ�)�V��:�3ԋ��e՞�����a[Y�SӇnʼ�T�aQj�:f| ����]��w�@9��iF����p�ݢ˨�C	S'1���+x�(&�X=)���͗}���vޕ��EIpN�������N}Z��u\�醁"U0�*�Z���9�a(5�:�uE�	B���r|�� ��c�B0��ד���⽚m���fZ�W��&��%���F����|��6g�.�_kQ�j�2��9�'�=b_���:n��ϝ�*\�P?2�������x,*".n����6�Мů���gc�ӏ��\(W�� qe^t,�T�u
��v��6z\Ky�>��P�4��泴�f��8�1uiĒF���zX�*B����$��M�z$x�_M�.�>����{%f�Ģ�"�l8TA��5�|;�H"ha&j��z���T�d�a��Vb]��~��bp�?���;k��p�Y �]�<T�R ��-�����"��:ukm�z������.����9����������~����h�<�tg(�m;�t>j��g�ĤJ�V��Fh��%3�7A��?�	����6Q������h�j�
_W��-��k����N��ɺw#���gS�$=im�^���nս�tM�$�0Șp��LK��)Y��/��f�ؾ�#$�	�p��/shNXn�zu}�k����g�S�ϓ5:9���wbx��*J�v��RW:��:��+�=I^�i���(��}��3S���غ��M*@�Ff��zZ��!���r=�'�)�ڈ#��G۔�2��C�cB�	Umh����m1��X�6�ɫQ�,��7b�����p;�o1zkc�{�[2#�b֜ob�'� UO��q�v}~y�7p��Y�G�	 ��Dt�a��L(��v�+�_�R�Sb������"�nY�I|wx+Y}il�00v;Z*`e�� L���\Q��i��
Q��+�O!��yu�n�,��fXj��Y�D-�X�AA�����pr)�3��7���N���6ߨ��O0��>����%��.�����.+
�ٌ�e�����e�C��R��f{f�@���k?M<з�*��
v�W<B��{�="�@2jӓ	�z����zh~|Ga�� ����QsU�K%�����
�l+R¹G#�;��L��K�Q��c��5�s�Ħ"yZ�^Y�4p,�ES>��i����*Δ�=�Y�@��4�C���>�,R�صu*5�z!U����n~���}}�`��uI�Sc5������o���
�oV�i�<�m�X}��/ϩ���P��Y����l��qR�`a5�d�A�3\����?ŷ��	�(HG�&��E ��jT�:���r��T|o�9PVO�����2�]쁢M�J'�y��=��,܁�&5s˩�y��n}~�eNn�=�o��}j5%�uA�D��H-D�Ǩ���9���9��$�p�������/�K�~3��Z�R>맫{O$���AE����B�C����u����_@�Iݠ]�l��,�O��&�7LҰ[N!�K=A�j�u4�}�q	��@��	�MUl^�0C�,����NC�����-�7�J�e������5��1Ndl��-�h��h���[��47�E'�f���xɪ������⎡%3���`���qO83�x]�Z��U��~v��:���6�,�_���]�l�>� ��\��E��>�K���B��Էp1��2&;PC<�*G�<I&Jp�C@�%�-+�g�i�?�xwL�'��0mw����/F	0�W����e�+��L���#!^��m6�v����-Ep<�jYz�>���|���邂�Y�Pq����: w>��C�,yUow/M�b�i��F���WZ��V���C�r�U2v�xm�<��]`��:Hz�^J*�tEǾ���a�3T��CH^z�ۗY-���5��\-,|�DBI�v��n$��I+W�vS\K�	�eS�luM �by�#طni�:���㥌O��ŢMT�*q�*���h�(�Mv��4�0w�N��:�W�`��팔��g3�
D4pri�s�'P�� ��rz����^��Oۼ|�T,�q�0��dʝ���6��s(��l��P_��&������
{�3ﶃx�����w"�5�:X >W��*=n�ui�K�%R�I�k�W ��T&픜D�$���������6I����j>d�E�x���3.Փ[�E�6?5xj�G��_<;f:���(�K¦/��B�k��r��}�&o9%�[�<��O�@�@�<l�Ow��׭^ɬd'ғ?�.]	���u$�?לr�=��U��a�ٴ:�*^��T�^� �b�@/ΰ��_�����Q��⣚,3�[P(�mY軥��ҹuЀ.�̅��SN�ׂ�Y<d�>��y�޲�`�[9_���{��\�"�zk�|j�:�R�A�p��U��F�h��� [�um�ʭp����Mؓ��<��|��=8Nʔ��иH/ܣ�@�!��P�A��m(+���g��`^�N܄a��sў[��L&��r$Ȕe�bo���ȰQ�-��eA5j�J{S�KAG�}]`T����Sq��?`k��S¿%�}��j��n�
������(O�2���ۀ���΋<]�P�A'a��@��	���Y�U��+��ǖǂ�:�ȓ�ϛr�RQ��&:��H������e�l����h��Y���(� *x�e֩������  U �:�Kr�^��b��0���M�<�O��6����oe_�c�����B`�8c:��y�'�t�F��ԟ$���O�m2���i=����b���tB#W"�%�1����FI v�p��c� ���9N�^^"�ٰ�m��_s�XMv�F��T+����D<���鞄�_���}ON��iۤ�_�s�~;\�R?�;2�d@�dq&��On�q6KN����"�wuXm {��:y��r�����������!%�y�%7�{���n�m��V�p�>��E��7��];󸸳0�vNn�g��/!!	Z&��Q��La2^�x�Ɨf���Ϧ-�l���CCN$�}qC��@�3���r?X�R0����rM��?��=ZY��Dq��h�%����1X���}���I
S�Z2���D��a��4��Kʐ�hR�^�Зg0Pw�{��뒺5`[d�9�;o�,��`c �q���tV&�6��Z�Ds�M��B�ΩO�?����M�$Ґ^ݰp��s�}���2�����J��`~3����K�㬈���Y(I���(����x�G�!��61�}��-`H=��J��0���z�fC�U[��W5��NO��y�K7�h�!�1�?ٟS	��G(4zA��o����D���&o���|�B�ig�� 8�(��@# ���*[������2����_�>�=��YY0�)�Md�G:�ܣ��5TK�"����˥ױc/%Xfw�:��4��1i��k���3�RQT��Z�I�����ޏx�����Zd�g��ā?>��:i�l� ]��٩� ��eZ�����.i���_�xlH�oKG�����oB��&J	���T�ѥ�9h�e�i�|ȫrnei� ���8���K�\��V��_jA-�p��ʥl�W3�L��<ч-Y�$�a�Wknk��rp�����B�vm���]�f�P}���&�ȇ��՚�F$4��[Q�}��\���O��f(}:�{�F�[�ࣷ�����ڣs���i�5��+g��S���ܦgߙ49XT��*��!�qsE�\B�LUek`h�[z_-�5�Z S	pY�QOZ�%D�*B�n ��tj]H�+��¿�A;`��p47�R!c���yd6���H����m�X�������b̓I��l�A'zf� �i�G
��ӁP���8�x���!�4�뮙(��l�?;�`����5���RW�B��Q3:A�j�-ʆ:m��.��';!֞��ֽ���X��%
"���}J^�톥�<��.Dn���Gt$=_�Z�)�dè�@�E��M� ��s7�A��lY�\t�**ɻo��\���N�W ƚ?ʴ.UE����Dx���C7�M�:1'�,ᷳ�1���@�/>�;K�n��̦�čUF���w�#���y|���/�R�(/��/��A�ya���/��66V�~.�Ofr���3x�b>�n�8}���@:��F~�TLҕ��N�&�@�I���[�!އ5���z��-b}< �q�=#HI��vt�S��(��8�
U���������d}dJq��"�s��6��v�8u���e�q�wh#���L�z\<�|I$ 0�1��Sb�b?@�Z�'ښ�8���O�7�>���5�
�i�څ�\�<��,0M�7%2����CS��Rf*ͳQ:N\����}>|>,������֟ϧ��JN�g���
o��&���}��\)��d!,?$ퟨ,���6�G+�,g�b�Z�!���)����_�j=Ȫ�Q�'���3�؞��8Sg�a.ؐ��	(+(��~˃C��� E�b`���K橤O��J ����?�8��gȿ�;o������KL�al<Ҟw�*��O�Ċm���
�i�ka��=H�
u��:�h����Y����LP�l(�7��g�$�����K��	�,�_�HU��r��il����f�E���j��K�DD�F2l��;��|��j=�}Pܪi�ds;�f��q�'��	��~�n���^(7rs�_$6kM���R�,�`#s����h&3�!b�0�0GF�t�z.f����T�B]Ӳ�p(g�l�kd`��d�)1P�Ӎ�r��
�FQ���!z�D��D�~f��"*0���
�#�Vbȗ�`��'�mó��db�bh!�T�E>z����},�u)�c���{�4�g~՗M�PjPX�5�G���J�o]�!@q�3�C�� �r�BZ=Q�´��Z�Fe����U;�E.�H����[�>��=q[�Zq��V��/��Q�j���v& j^)A�29A3ufu�2�S:>�\�N��/q�d�g������#���iX���V�
צ�^��ظ'a�lV�|���j{I�=�u�<�	*�/�����T6��i��mI��KDo��s�á�R '�k:��&��6�B��<����+�e'��`��ԡ�,���헹``����_��X%��x�M���I�s>dq��2��4r�D^��m��@0��]aG�I�'5`S��1˰�.xL.Ox��0�X	�5%aA��2a��8 Rz��������ծ�'c`�D���x@|��������3 �k�$�sT��"ZE�ޑ�n��͂<��pT��U���'b3)U����9ٍA��c�z�'�o���0�M_�7]�����'��Z|��]�<W���l���U0$/@:q��k_���k{P����u=+I(=}�./�$���[� ���:��}��"�E
�6��}n(��e�YX�����%�D�Ũ{�
j�兛� <֎�n��f'�{���Z����=�1�I��>���Y���cIl�D5A��-E�썬�[��{��$��>�n<�M[�k6�L�C�	�<������$p�y�9�Xd�	���
I�x9��_��jL�\��1y����FÁ7q�d��F=�Vr���`��$H/ƺb�Z~�*�	
��OD!a���Ƿ*���z��F����ey+����v ����4�	~5vx=��v7�2�~��(�ߧmͥ�H��Ȓ��ok��)X�W5�B�>�����N*�N��y�:��Mf$�|IK�\S6�C�%T/텈2�J���@~�+�Y�ga{�`�B��{�reB2�m0�\h��M�l��^��5v`)������G_4I���R	��p}S><8�D_
�X�P��:�����sҪmI�E崅�R�[�ڈ��'�*��  ������e��հT4���J�`�Ƨ�.]TZQ�+��3D2�jv�Bb�r�
�\�����*aRTQXBŭ��Uم��ч�!$)�l`	���u�V`��ո7o�^f��I}�T���cA.�E~���pR��SK��@���uc�l�.�8�(�r��o��	�,NqJ�[�$��r���ʹ�
�$re8��;�H����䮎� 'i��C�����Wߖ;M��T�=2���6_�^#(�;��F��a��§A��8V��'(r8	�E��eDx<�$�xΟ�hZb�6���y6�>����E�_���&�eL2N�A} �f�H�����KFq��}�U�93��k�,9�(!��o`c���������<�A� ��k(��uQ]$��͚4C�<j��6v@��4>%�Ϭi{Vp�O|�����n2��M�|��d�V�L�
}�J��5rw��ew������4�\�v��_���y���e�Y���}�){	��Q��8-�3�
�>uW��ܢ wQ���ȋ���E*6o���EOf�a	��}?����G	����v����R�o:�ر��Q&1��x 
��~����~�	I[xXg9����w��7=�!8be'�� �D2uI�k�m�D�����l��Rܰ��r�����}��|cK^�1��+��@D�-1� �>ļ���S~�v#.���T܆�0V����)�'a	����3(�}@��Жԁ�����U�¯�Q���8�Y�`�w�5��V+sU1P����:Z����Oę�A��\��N�I�U��d%����&0\�����H�.�c�%�*r:E��9l���A�b�T��"�#@7qEqG��G�l���:;���/��s����D8 ���S��y�mr漸��t�o]�n���_[�ς�6g��U� >mI:�t&Gc!)����e(��I��i���M2��JeG:oZ�2�j���'��mO�iW���'���}�6�� �ߔ�CG�s|�F"�f�!��(����Q+�[y�-u/v-bw��j߬o��?���!��a��[��z-*��3�!���:����J>Ѝ��$20������[<�a?;���L�^mb\��!��1e���� .I����B%1�Kƒ�f7�bj�p�Wx�~��7:4��o!΂�n��}:u:�|#}��I�C�m��{KBZ��M8�Z��f� {Y'���Zd#����h�v��s*�N�q�=t����s�b�LG���ʼrǁ҉���#��/���~���25K�E��Q����&�����,���C�г:T����,咆'�I��{��|"^��Q~LR:#vV%\�Wt!�.f:}�d�A�D�n4�"��7+�* �]U
K]�Pչ��d�듰���/�O,��w^i���C�I6RtW[��@a��q���c� ���r�0H�e9���� �	�Zr���u�sX4ϰ��/�t�u�ۍc�{|�4�Q��T���?�G9b�'�*�+��~��\�B{���ԌX!xY�0o*���<[�=�ŀ����V3��]�е�������(�^��r�l�R8�7��O[���.�5P���C����Į/���Ԅ�@�U���&x}����3Cpx��ʯ1�t�fU�̸8ma��ٽ�s�-���q�o�H��VT9J*1���z$�߮<�����g��q$�jB�l�M�d;yy�mێOpw���G���p���v	��8_�=l+�um��9�IΓԹ��Т�&D�������1�ȸ��(LӶN��^"@���^
�	�[���>���ξ�~�#���y��z�Q�c����8�p�oԴ�ߨ��z�~r]�����<d{M3�uo\�/P���K��_�&�������b?�'xp��!���f�5~�5,9�BH:.���
k��������*?W�'mZNɦ�u�ށ����'r��T��-q�pwc@S��Px��H���:�)1i��bI�~�����p�Ϝ���.$���]�e�L�1	��7+���m"��W����x��k3UN�[Y�aՉ���A��!I�R��MiP8�:	v⳻#,�7���[�����(>��3��Ǜ6�2	d0�,kך�����#������۔_9�NȜ��u��j�->[K�,��̨T�զy著��F���wN����A&�ˆ'��9ɫ¼�w'������x	����"�xH2}����)#��r�B���t:]V�xO
�����K<�,�
�`�Ӟ%�~�:��[��U�t�(,�xΙ��nD�0K�'��G3��5�=^# o��)��y�r)H �e�z')N \�WS�^�և?N����Z^�Gl>m֓�L ���5<^ʉ�e�i�(���jz�SR?�;�m��8�[Ń��l�1�?�l��j�e����I__%!����f����VwB�pɦ"���ʺl��ct�;��ߜ�Z!�:J]Rv8jr�YT��!/�� �j��u��6��l�u�q��Nǥ�e�U��H:��l��͔�u78��}�3��Rﻇ '��Ъ����އW:�-g7;�_����?����DRQ?��ܮ����T�FΚ�ð�)�sL�I"���mں�����ߖ^��V�[W��������3Byo�9:��+���N��}�a���0�]�j�IM��zJ�O5e6\*�{$���>C[E�?�_v�~gw�፻N@�$1���{��)�i?���`U
i\o����֪4��\�*h���,��>1��NGVU��)����LxQ����% _Z�{|1�,���F>9)��7�%ϽE2�M���^;Q�F�j�8��DC[G��<.�s@cE��g�X��(��9(�n@-i_�u���^�7�	��g��[*H	x�9���W��p�U�jp������۔��f|=fT�LG��u�~Nq�ndx �Ht�lFU%o�P�󱙭.���>���g�=��H�a���z�&(�0�S��G0>�F���s�ƞ�%��	'��7�����9-�\d�ᢜq��~�G޵_u�/��:7�e6����^�2G4�L=7&�\�%���I#�Ѡ� ��2/�U�n��+Ԣu~���q1̝���t�!1�'W�R�F��5�b��g>[��&EF�5������b�x��K���{��k ���h҂*���Z��R��9���ʿL����Hk;v��>Ap�N@qc&I��{n\1wn�����g�	�=|���{�͉�Ԫ$v����&�J�>����UN1&��[|�OJV;�(y�����7�Z��S����/�C�Q"���$�D�{��`�]�_X_%�+'�z-��&|��˓q���^���d�G�����v9-JƜw��v�d ��ϰ<(X:�����#�<��EX�c�s9R�|�� V�yۢ��_J��Q-%o�����N���e�G�CS|}{�U�t���Z��QB:A��p�c:�����W���6�~8P��ᖃ���c� ��3��Uz��sD�]���".�.��&į��6Vq����jcy���~�]i�È������o�{	h�t��m��֭X#�u�񘶙�ϔ�u@��0��
�DDHU��b�J	iǲ���?�����-��Ws�6���k!F��/F��Ԟ�M�dU�'�f'�h���Hk��\e]�ϞMs�CXu|8r��DTE�G�ٹ@Q���3�6�၇"[-���|'������y8��i���>q*Ƃ���S�ɴr�Rm�S��+DQL���jCz����yR�Pl�殫����,��B�[��]v�hDn��-�r�C�?���_�tg�*�/�I#��������0�vVF?rR/2�}|�r�Q�x�������)�!j���﫰�����qj�9�+���M5�	U2�AZ��ꧪ.�c��u��jK	F��l������ ?�MO�'s��~����}�s�~4<̽��_X	j��DPқ��Аū�Q ���7Ez3N��ݻG�49�H�㩟��!jH�3p�:w���e�v��{UyB�@Z^�Z�4��2�+-e��g�~�+Y!�����ol4��c7��a�v�*��r�~�}a}9�+�f+K��k	��8�͌4zP3�,�Ӕ�{�˻M󀩴`�+^�����.�TΓ��`c�0��Q��	��+�/��¼g���b�l�)���|g�{��eG&����r�s�d$4:��]1,,"����K����pB*�Hǝ�'L�S�M?��VМ�����RB��1��ͬ??��ws���L ��sݕ��*���VP���!�^$8WL��V����
�=Te�I/��(���4س�� V�=gՠ��(�*y(:��4Nd��0 ~�	�7hJHh(���x,z�1�nh-1���ȆNM<���rc��cj�5/W2�+��%�uD9������G�&`�����)=AӜ���i�TU�����V�^ cEC��q@�t[F\�dW��a	� Gu�|�3@K$��ر
PK��e�@���Z����S�o4]�bn��k[�ƌ�*:��>.^s1�m㉒E8骃�g2�b������P�*)y�J��VNP��6�T��:{�=�'΂�8�L�0݌ȅQN��[�ȟ�2
��F���$���>�S��|�+*�,�����md5�ɚ/�lf�~̠`&`R��A�Y�KшK(9�%���_k�$b,�R��w|���Cq
���z��b�v�n<�}��CS�^�ˠ�Yp.�����e:�B9������%h�p�Tٲ�o���,i��fb|��&��+
_(/��R��VɁ��E?V\ȼ�� ��>�q���&�����K�W`�	�� `�7N���LP�o�0�-�$�ԎfT.ꝧ�6k^-�N4S���m/3�D���^�����te%�<Q�X��W�O����)�ݚpGt�U?����x���{�]�������\�"�|`�bT�l26QA\O*>�ν_G�!�4��,�@�B���*��C~����~'N��~z: ����o+���Z�j 4=���o����'p���0��Uee�e�ue4DqӬ<21���w�V�gpr�El�6�&��@5/�b�5���K����<�T�U�_o�w�TaZ����n�FS�6r`�w\���H��R;���H�-$27�[���md�e���D��#��GNNp<>��:�����ȥ�?��0�7h�w�r^[l���]f��% ��[Fs���ɣAZ�NyN݇�s�Ka�N����A\F��`%|�i�3��K�tV�d���ǛQ���O'�~���-^��>_A����K��m�ݿ�)ם�sM4�8{�����y�ʸ��Q?�h�G�N�Z��DH(�6�Ųi��Ip�#���m*��Y���
��y���Y���+��;���c;iM8�LC��&�S"F�������6:[�R��/G;kzk�\{�n\nWa��#,��t:-Ac��]�l��̔���|�xz���D��SkO�#�D.
Ҕe��@i�a5 ���d�6��.����5�X[$��N�2}�;����j�����������'�q��>�t��O�6���êlONww�O}A���}�Z��I��6�U�.B��KY�O#V.�H�U�v>�����-�W�B��X�l}��R��o�y�2�l2��$M�-@T�\E.^����J�Ew;ɻIr|o�vӣ����N��{�x�H�a�'�ЁJ~���6�&AT����ͪ;������P.�5`,�x�yuX87H�������se����[[�G�%�7B�4p����2��wfzk���9��ض'O�6չ�uNjs���v�7w�?F�������>:A�&����@7rh-v>�e�O:%�Ie�Ċ��#�V�_b��MM��2 ��G��LJ�ZCf��`�w��vߊV�<����w��l�[��=\ڑ���cB0����aLc�i ����ӯ���k��p'j��,�C+���Yћ尕�ю@���|y�\=�a�yS��F�@()�E_>���6q�%����X�V,bXJ`#	�|���hIZ��!�iL� �zZ�i��5�'�	|�!�Q� z�s���� ��ݶS�gk!:��	h�L�O�#�,�>�G���|��,���,@���>�U�D�	���U:h@w@J��g[�����֖����GL����_ߚ�H�j4�B��;���hWSF\4 ��yo�F�e�Bd=���ӴcIW�� X��\��s�=�]35�����E���� ��#t�Ӯd�2:�M��ң�F�#�&��D?�z�7���!X�uweק�/����	�m���~�fܩ�����T�GA�1�A#v�8�ߴ�a
ʉ����>G忎Fy�~����>�1�v����?��$|w���7b�@nb����.����L��.螊����f��gϵ���:ѩ���S�3v�߬�������������_M���޶Fx��u|Ȇ`�ע[΅�������z���:�Hh�4�8��ǌ;��єdmc���å�$=��/	$��龦��"�؟f�s�@�T�<���S���j��=���%yG�߰�{I4�"�C��nA���j
��_ˬ����wZ�=2��[ov�A4��K��ָ|�5�L�9qB�̲�͈,��QƧҰD��T�����u)_7��s�T�>y�>-�8��<
+�-ޑ�#X�C��ޒ��/g��Ϫ��<����:Q-�Q�ri��%�L�9�=ڌ�����{�Z��F�� ��V2V��Q3��	����$��6R�<�%T��=�417�+0��D�7m� ��>dn_��+�Ŕ��w8A=��+L�+�5@Q�6k��p���Sm���4t]���ʵRä��� N�Ox��"4嵷`�߼C��(����#�i�eԇi�[)��������k}R�k3ϥd�p`Z<�J��P$�[���w��}O1���W?��#�KV#���Ie�&/�Y��s�l��V����%�D=�����*����l{q|�eM�� �E�:;�����%=���y8��t�f��s-�0]k*���F��s uy �9�X��"�t��6�Gi�� Λ��Ɗ�{/؉4v��Ht�(6���|_�i����X����e�I�0���qN���lt%�{���>�ʬ���	�r^Gm	�#��lü���5,���݄p��Ce*0&8��Jy�.tD�0B�\�kF�ӱ	j�҅
K��������"F�O
��W��	�(;����b'��O|<%�̑ ܵŜݝ�q�M/�l�z5M�s����ȹ�%�����a�㥭 ��(n�#"���sUs��l=(�-�P��j(y7[{�~G�+`H����nP2w8Y�ʄÖ��n�l6��F�(k�ۤ<�s�w���U����ດ�y3Jͫ��YGF�R�V2������.T�޿x�����+~��qH�#�������p��@ܡ^c5���u����������A��uF�tb��+/�L\�	y@Qh��>���]L�R��F�(���5w��j���32�,mK=z\*ZWI֩��HEg}-h��@�R����`��Ⱦya������Ł�Z�LҖ��k P�z.6���j> [P�c�-�"����Hh�(��Lf��,ӓP{6�^[<'�>�Q�c�7�����+��&�H
�3ͪ�`�%�⃉S����j����e�.N\ ��Z���^~���b�9��qA��
����ピ���r��h�3 �ܔiRzفd��E�':���Ƶ��":�eR��Rh�I�݌�r"�|~��ƙ�]p�@V|c�v���s�;
\���s����.$6���
}���la1��)S����\���}��Vi�`9����bcރyn�
䝋<bJα�/��H*cLA�܂vz����I*�-�1n���'Y�i��ێ]�ׄ:z.v��-*���DD���_ �J�^*��Ni���-� �Q�,�S����'�
���)M��ţ{���'���ߐ�X��]sk�P���Qd!9��/B��u�������:Q�w�e&����-I�Ń�Ea������y�!�0�"��S��R鶤Q$ �1�CP��
�U09j�o��o�e<��3�Y6�w�[䂜+�Hm��l��[_X����y�@��tA]�W��`Pڗ��ǻ�l��{�!�Z��<�&7��Bu�G��a�(_��Xc��'������Ҟ�M7�EYm�m�@�����g^��~������ýp����{�����.�O��`�
�C�v�\w��s]���}�1��X
�3�'�c`r�K�**��Zv�`��F�6�D����h@�ʆ��C�d����^�"ˊ��s0���i ���R��@�ͧ�!��i�2y�	ikA�������7�U5͙�J���'��Oޢ�s���]9��~{,_��,oM6�iڶ���dDT{���V��2u�Е�,�>��T�ac9���w�bSJ��#���.]6+p�Ii$��\��|0�������@�\^ʈv��q��Rջ�����-5��9�
)�l�L�0�g�/F�Q:�1&ũjG;^t�������I�֝ML�,{}Y�����.5�A���%�~-���/46jA� Y��m�BeJ�6e�E0��=(yE}����#���Ix�u�:לzF.���f�FV
�݆�@IL� 2��|����GA�1�"�W��ڡ�O�:�Қ2��w}-6M���k��B����8�3�Ǭ��Ԍ\�������-9���-�A���Ԯ@�h���H��٩��{��ZTↂ5h��+c���5+a��u�������:����,.[�m�9�Z���?��T0	r��}��g�n�غ0���A+��uo��\�T��L���[&Y���a.��Jt�vM�3N����"sdup:����^sOb*X6�S�x�q�j��$����5��>t)��$if~��|w|#����.2�,-����P��9��g�5��+�����ԣ�5�\/M�Q�(���b�帙]2�/=@�����B�6|�i���K�_e��K�גu����w�dw_I��|mP��Li�	/ЮH�F`>�A�N�L�ɜ7�J-��+�O�Hl��%�c[UB����+�d�T�I=�-��92p�����K��8I�`��xU8�����5	�l�8*����ܧ,��!���䐸S��n���Ș�,C$�㏂�j�>�E�5 ���g4��>hȮ(� )�FoO`�Ы;pFM��H44�T�)h@�Ef'��Y>�\�/�4"�n�l�=��<��K��a�P����&M�W�3|�k�i@�IZ��G�a�>���W�tN�ơ%���K7��*Jݓ�B�"��Ѐ_Ϸ���D\b���_�KW cfȴ<��Q���Q	���T_��s�N��d��LpSpm���K3�
/p�#���쑇!�-m.R�.{F�����\��]u��S
�M�M�0����x� >�"S��M��B�����P}lƓyIek]����U:�+4Ʊ7�ሿU01߅�����/�^���DO������i���`�B\P���bT�U����g��&<l{�9�^��i3�
Kb�t���'`TyZ	�_y6���K�!��R�ʆ	��Z�Dm�:x3*,�ݓ�qV�+P�'*P�W�m�fl��"[�)��O��.Ж;��¸y�T�*���k�-K�v��U�8�/c/ x��>����^���S��u�0�2Ƽ�����xǂ0Yb#=~4���~�R��z Z��z?��LΙ�1;7�3���(Q4rUB� s�^u˓��#��H��ת��k�
����F3��%i�а{��������S��o���j�̈́�W����l1X����PDd��Ǳ�J�����ȷ��.M��
�[��_�P;���.�	�b�rN	$Nz�9��V!M��ŧ����]R�©���}!=*4��cos��Ҝ��D��^KX��'�Y�)}��U(j;^]H�h�ED�t�"���nR�D[�[ 0۾�)��ϸL��-����I���o�n�,Q�Tkk��8�A�6�3L�DY�����߰���e�X�h��� �^�9L�Q|�О-�ev��H�/"���0ϫ��Ud��G��1p#�9`��b$�>�U�\��uP��:��WJ���)���������i�|y�O�=�.��K���w&� q9�8�r�|�ven��{!����)C�q�Ȟ��!i;H0�Ñȱɚ�%ut�?��5~��q� n唙�U��,gH���xYw�U׺$ �_W>��U�x����p6�^�T��E����呵�q=�̧��T�����w���6�<_��vv#Q)�͕vj$Eg`�I�E&u	ƥ�G�>�C˒�k��l���L�$-M�D���Ԉ�k��b�7B7�y��d��U{ve/":I��MtB&��a�b�~����w�hK츸�
X�T���DF��prS�J��9=Ҋ{j��ר̭���t���u��418�����65`?���WH�&�ˢ���H;b �*[/��3�t(_��r��up� $�M�r} /+�S*_���=��-�����.���F'�d�h!�'͒yjTD�2w�_�_�����r � ���~�)GnC߉���5���ösH^c�2ԡ�� �V#+Ҏ~%��}�BE����:�����j�]�׸����_���AЩ��k��I���X�x{�{(�oCde9~�VR�/��Ӧ�2LE o�B����8��O!���[�?�Ox�~�����{�cpfɺ�!��L{�諸��}t9fX��H!�%�����ZIP]��K���'f(��\����Pz��h�6GkfI�xfм�G��L��M^����9��\["�&�&)d�C�5���"��x�����R����G^����#W=q-6k��%�3����b�:�D�������,{�����}�����
������^'�mH[��X��\�d�),�y�c��Q�xh��S�J苓��LU�
PS^�&ќ���B�i���-��3�����B8��,M<\W�C�r�L���� ��a��ǝ$0��Q�ߣѹ�/ړ۵ݺ�4��~�-�ݺt�&�����wP����ųR���jii�y(�y���W�@r��*q��i��<ClFw@]�����d������e"売����@�G��QZ���i�E�,��FT����J1��9�����;�N�oJ�k�'���+��6+�0�c�^zB�������d�?@��x���2֘0��!g΁��yR
�r��������0c毚� �BqO�:r{���g'1�K|Yu�{�ݢlv/��;lO�\���abmq��f��э�0Sz���.Y>�	Gy͎�����e���>;w"ڂ�rJ���|�v;������Cm����-2A�8��5��c(OY��"rb�Hރ3\�[�%��l��:�^�jc1W<�&����ҐQ�)�TPC�����ak�r��H~i���S�V=ϯ�=Hi���K��S�\y��Xm��껆'�r��k�a!���b���z�s)֛(�y�@Y���r3�֮�z��O�����iq(�0�wY���Tݎa�*69C=:��(�f��S�t�{K��Q�~��15~�MByJ`�'_�SE?8є*���a$�$���Ĕ9��K*�՚ ye:N�`e&@�!�N���ۙ͝OlS�u|�`�OɃ���9~Rh|Bw�����p��^(���Ai�Rċrn՚shnX�|q1��w[<�z7l}f�;p������lC�uuR�b���-�Xk7���/�4��O��׶� \��ë��+��BX��'�p���i��l�d.b��iŲĮ��Y'���R���_shMyȀ�_C)���32!]�i�X�J6Z�J�'���a��N�Q*�%���j}G�3�s�ywW!|ζ��~���kC��%4����ڜ��`7�	��z��8|Ć�b2��k_�2�pf�c�0�Y��P�4|�l0�Я�`p<Xy�� 3�0�_cɋ��Ϛ�N�3Ge�Fw fM��o���Uab]�`o�+�UCb������T������=��lJ���0��"⯅3yZ�܃ʇJ�(?w����g[���rUҀ0�2ak��K���!3���� ���ב���琀M2�����&���&����\~V�������ٝ_V}������B,[BT=��I	�i�q���������w�����̸FX�R���j�'&����{lNĔR�05�F��'�D������;��|�m�V�ۊ���>o�@������˙V	C��8-�**v��O6��zjF�hH�;�}��U�9:$�@��}soCw/��x�u-J_���(�C;d}ܚ�(G��?�S�J�]0���i����qKN��؆�:�b^�̟=ꊼ4���ؚ���?'䝀�B#t�?
��i��c�ٌ;�A�ʐ��%dȷ}�(nU��p��3*HWp�QWu��j��X�7e:4��8SH*��\ؚ�j�����]J�[�X�*j��neN���$g�P�Eiu�4k���:���.��0�*N���/�2�DM{��XdH�c����q�H<�rW�K��3�P�詀��o�P�����6��g
�{��ƒ��߯�d�*��}�z�tˉ��}��H�^څj��$����ܹ�=��7����[��U����3��U�?��k���}���ؽ��ؠĊ�^����D�x�"��0��}8G��y���%!i����9�:�?���Z��W������f�ʅR�xk��h����jY/Y��������]u�c�AʳI?{�\��qH�<{��FK0��o(�-�NȲ�H}�؅�>R��͎zpzj�M\��F�ͯJ<\�Ո]�u�o��߅��|��
���̿�n���JR�mdU+,�*� L"|tC��ǝ�`T��E���S�'	�5R6�7�ӛ�G��XXe�w2  h�nkU���&�n����4��,��0 �O���[������P�ړo-2��������{����LN�9���������_nQ��s:�wܮ�nZ�ٮd�6N�g{8z�����P�בu�?�@�H�5
Z���FLmmؔ"XހQ��3�o��}ޏ[���^�뗬|�5�i��/�l�[��Ne0�iL��s��Db��h͏r-��f^U�>`�h�}]y�L��v� �@2u���Q	����҆�X4��R%��_m_9����L���v��0�}��t�*f���M��n���oU�6!�&��$؄h�Q���ȵN�-�Ɍb\��ӂ�&Vq- �#
�x!��^c��KMfy5�t��� �����Y��Z��ȅO0
x4�{�b���l����Y�+ @� �7Ϡ�ǻ65�{��!�!�(��އ�1���~�`��t�"+v}~��i���n�:"�%�Β��0crj?�PW�Uk.�����e���
~<� >�����?���^Z�<��>o)��7	$��=���;i��"9+w�,����%1�Н�� Y�>�m�\pn]�e���f�kK�X�k_|$�	��L�N���]=s�������6Ӑ]�x�絍��[�7K]�y�C5WH�#��ǇƵ����9?��{��pj�;p�0@��!�et��TZ�U���~�ԉ��f�; �+t��9��:an��r���&���I ,� V614�g��N0��>���PZB���O8��uf��r����b�&	(�Ž�p{(b�q�gZ6Q}
Cׯ?%I`�nY�+�<�Ɇg�{ނ��͗��/�����\l�m0Xc�uT�	�N�?��363˄�3`�V�=;>ՔTZ�cN�����R�C����!���/���-�PwS�jb7P
��}-~h7���=Q���bxVG�l���8@DQ/�na��U ��Ԫ�*���6�c�=�NK
'��0$��`i�S0*���ai�����%a6
��#�c��8�9��\�"���̀��Zwz�wМR���!�VoUŌ3�����y�5�@`��/���t~;��(̡�\�
��AH]#��^�$�,m�/J����e�g�ʁ�/�W�:�v�����rS����T�MR�-���^�Y?,v�2���`J���[+� 羵��?����}>9Rb��C,o ��8���}ԋ�i�%N������������<w2a�	��&�E��3��u�^�3�'�// Ϸ�J��$�<fygd��F���*���*85�#l�l#n��D�t�Ig6��$[mgv��h����cҷ�$f�t���F���+e=�_[;���)
�h�$�1k�q�4�ũHv��;ZA��ʙ	N�$O�jj����TW�Gl1��I��^�#������]��u�ڽ�,\x�?�aE'"�]N�Lf���� �z�ߢ��0�E=��1:F�һ`I]z���O/v������ؒ���W�푢�qt���,q���uTi�����e��[�˘-���YP@��l8��w���І DD���]�a5���]�x�~%+�0�M��mqf��z6���QX�W�Sz���9�s���m8+|�18��$d�\#�"9{�����g���6���c_f�czZ�\�n�'���'�	�h���5aD����U�'��nǜ����5s�fPS��(�S�Tg����=����]%k��H0%���'���{�Zķ�N������d^���S%c�~|~�Z�:һ�Ҝ�1�P�(
y1{fӲg��+�B�E�%��՟�bͅ3B������Ό���!�5,���(QHn���[���h��pF?��pG�߇�p�*X��r�P�r�����E�ټtIɞ��f,@��xYL<��_@�G��y�^�����Qj�5 ����<"�,��3'�g���у��Ƀl��[���@y������c,�~�O��#c��egTl�������hM�<���[4!`����Z��Q׷���۠�*f����U���D��JH%@����[����;�εV�^Z�w�wܙ��4��3����j�ؕ'7tRB������n@����Rӄm�ƈT��N���gB>^�1��q���2�Ɣ�H�x��mT~�57�����&B��9�/1[�z��w؞Ab>��,V��Zq5��Kg�F�_�r�g���t��,�����x,�s�G���q�a�)�@}������=+y���*�:��8���>��ͨ�4l��<*�Zpd@׼�L�T��m���WUwvͪ�%G��+�[C���ْ}��DM�;�k �@P����1�r��W�N�Jz6��]5��y"XW��R�rR8�U�R�D��V�}��NZ�Q�4�wjQP�����6���3X�BWu�(&��a�v띕S�.���.~�խ粵�Ë����B�������٢��|$�?������eN��&�m5�8�9vUR�(�m:���Kn��a4 Yx+8W���M�qA�R���:�]�iJ�3$ �W���P'�N��Pa*�E&�pk�~�7�����i��s��e�%����c>�j;`������f:�u��xP��|!�|�g���#wp�K�c��ҵ��#�9<��ގ%A��y������YY���c�j�Mp���\u�=$��m��`�ձ�A D�&��V��{5�3������I�d.�eU�j�o�w� ��t����ϐj�W-)˟h�LTƭQ����~R�|�6�R��'԰d�<^%(�,��5�C�S[=i�>�����"1:�I��FeB��rf`q�(���v���F��+���Y�RB�k�q�L��[j�d�K���U�:� ��xݘ[����$#�vM��/2s;^(��v���8�q��4�N?<+�BnH�x��)t�.!M���{N���EE�x�?�&��D�_��ʚ
&��j�,�`���P�w�WT|�ނ�h������͹(F dt��ȢS�J@�S٥��9�-�B0��T��I�˪��vzZ	�`�\��R5�f�-��k�I��>U y���Zt�aOr����3����e�C^���$j����s �м0�v\���!M]}��8X�Z�n`J�gcg�L�VЪj;�I|O�	� ��
h[�P�:Κrf��Φ������P�p���:�@���?:әY��YEc��m� n9H����F2��ڬVδɍ�xt��NV>���[*Z-��W�J�;r[�S=.	��v1YN���m��ҹ�� }��Sȱ[Qn���U/d�Z��}ldH���K	�IS��w�t&�����_uJOh�	{��%єÒ2�ufӉ�@Z:ukz����a����Ga����_V���8��=�Lw�UwD��
=�a��J�jNvl>�����: � eR򃛘��5yJ�f�E����G�H��E"��V2��2��!]��.��+
��ٰT�g��O~a�D5�Τ��t=��qמ��K�O����8H+����6�C{�S���Q����u*�,�6�:R�Y\�(�%.A����t���f�2rr�_5yk� B��A��1+���ጁ�N��u�6ۢ@�nf�ߞ�~�۽v���@i���RH�@2�9�3��Z���
}T�E��_歫5�ʥ,�TaK���40��((V��-��`��d�A�Q半t����k��0Kh��d��\q�D��V�Z7NI��-Җ��ሌ�0ܱ�*vUz́��_Щ�fh���g&����n��uN?���Ě����@�Ǌ��qfm:%[�[�^�Oz���dq�m�@P6�wA���z#;m�s��-�|F�&��0��`՟S��ϗ�������a3?���kɸ��3�:C��S#����U��^0��\i%�t����@.��z���:N���18�汵֔?����@ɷH�*�s@\�%���ziW����G�J�PE�K�=��5�f�&ntr]����E�l��A�������B�(�.�����d�$��Y�)CI�] t����J&=3c�,�`	�`r^Y<�Mp_&�#�;��Z�Ϩ��%��/���� 0S6��V<vن��X�#�P��fJ~;�/+I�I�@ax�`L����z$��q�D`��Rی $���N������ڻ@�y�`��oe2�`��5��o��Ypt���=�W ����T�+�"���?k��.�eԓc���dY2�.]h��vMN��d�aQ�M-	�q��-��LFL�9[���֭�0�	�`	�5)�W�t���:�9�����~CD�P*�2"|��;;��x',��4�/��S�[U���&����QC���H��R�{�h쯀0k�k����U�p�kbW�>;������ʊ?�ػ8ly�+Z����-_2xB,�w�EQy\�Ʊ�������<D:@�o��L���2���&�x�<8�������?F>��V�8�V��� c�����8l�0��Ɛ'?Z^S��>ZR�0i�F6ފ��֜J[O�fwz�v�lk("f4��A/����.��WQ��n';�����C�ƹ\�
k�NM�[#�J_�f���q��{����0�id����kS�]����;���`��N�qz�Qs7�>��`�JylZ%ǝ�(	B��d�Q(�).ͪ'+W��Axb�>�s��*w@�*EN�xi���9Hj��F�_ҟ�h��#Y��{�,*rW�z&z���~�Z��@v0N��A  �7X��k�KpQz�#��%#���LBD������iP��pT����W��-w=���b�L�f���~6���V�s��9�����q��=X�mY�
z���&�M���MuVI��8a������j<,�:�Ԃ��������t%g��8��eR��̪@ec-Y
����{�Ƙ��/��y�޸<��q�y�S.�x-��)D:���2�nW�O���q�f���xa�1U)/(h#�/��E��|����r�ݰ��&;1ϲ0@�=(�6�踍*2kv�He����
OB��(��ٮ7]�"F�p���ܐi�dl��Q71�"�-�OW�g�0dAI�G(]�̠h���;|�+�٢c�i����HuRs�c�r����C|K���(bט1nM�0������\ᮈ�/
�8#�K��A:-���Kk ����~s�s�J!�$AIԜr�q��Gu�
��h��"c Ў�"�b���e#�MբEy!���s�.��ϕ��S`�:[�	��5~���2mp	������uM�&00�D�^�:Ćl�l]�
T���m���.|
eW���!A6��-}�z-�8�|��Ȳ	G�N�R->�c&J��)���Ŝ��7@����h)M�����6+������K좮��ʰJ%������T!�|O-�@��H�t��=ܜ��i�?�L�9�F �푊0^w0��1���'W��}�V�� ���')���3^�Ə�|��L�� �	-8c�����F�����_ʄ��P��2�K/R˟R��4�>fv�����gg�!�B�WG�;��7źhc��t�`@�'��������c���,���Y�%\q�m>x��/̬��#��V��]r
�Ȭ����@�2�]G��J+@Vm���m#cE�ި�E1�(��:����Ҿ�bh'�z���M׽�e%�Q�{a9�}��ކy�0ɭ��ULq���l�6G`8�CF�0;�n$��c.�:b�g����PJ==�,%4�ٓJ��`i!̦f��C�& _�j�ڎ��H+	b��؋��Zf+B� ��7zPBe"�O�A��2�IN����wg�)���.6'^��]_*Ru_�-�=��p�oV��P�w_�p��Rn�&��Q�q$SG�2�$Y$��^j�N/���M�W:荙I*
ЬQ-q\�z�y����%/�9���	����2�	��,N(z�P*W�U�$䬃�_�a��M����\�z�u�\[H��7�@���Į�;��6{����P�aܚ:�Hu�:Qu*m�7kχ�)2v&<`��t�Bʟv�CB�K
6N��X�V��~�}��/��]�G��Ղt���ٚ	�,�&k���.��Ә���u���|��1���feX�M�7�R�����P��V�y��]R��jUư,|{�H����ݓB���C]Ƥ�@��^Z��d΋�FP��m�~U��ޣW�J��7y"�3�����ַT�s|w�$��={�� ňK̏�݅a;8?��H[��%K�j���"4�JJ��RE5��}#U[��P,��'I��@ɀ���J��r0cW|��Ǝ��@��r���Pm�\�"Y��l����`k_k*^�����uQ#�`�A)x�\�G*�T �>o���Y���A�#�VN�1�p6PJ����u�{�B!=��	1öB؇�똽����%��9�	rX��	�Q
Br�b�=O�0�u�w����}L*��Ŗ���8H�s1�QǑr�� �Ve���m J7ª\a�j���?A�$���}p^�PU�P���ǎ�f�q>H�ʑaIX�!c�!=gƊN���j�Bb�cx�=�DÏ8��+��T�bԽO�1�V���5�eU�N��$���
A���5D�a�?$z��,���?��/Z�7q%�X)�q\�M:��|2�g+�eU�W֍���7�{,5��j#_��������lU�_�`���*<X��*���j$ �����V�O��#���]F����\���BJ+��Q��Z�<���U�-p���jo��K���=I1{:�Ԕ	�0M_re={���K�sW�]X�DZ�Q  2����p��2Ss6��P����A���d�����GӜ�]�F
��]��R����1hp��ս+E#mdDaN���"��{���}��q�tC�j�\���$f�b<�Y�Z�h8�\-Dm���l�(4�4�Ayb$����b��Lw7w��u�L/���!.BB_��|ð�:�l'�ޠo��	Fx�oH�a,�ޤkn�*����r������I%�[�tP�Z
� �B��>C���������4�XI"߈���l�o�+�ѡ�����T;2qo=_2I:�>ʖ���h�$�h����T�X�k߰y�\P���ЫʆzQ�7�Gb���ɤ��Z�v#��S=��U���ά1r�ZVv��0��UM�R�Ƿq�ަn>�Yb����d��%HO�30���bl����{C�t�,<.��u=Tl��DȪ��?E��;�۵y�f�n�{�N���ײ�FM�LX��gS�A��2���o�+�g�����:-��K��>>)û/P\O`��ɲ��gT��r���5��(Ɓ��Rx�L�c��T�*�"��y�����L+�	y|�Q�R��~���ii0�=��q��|:+��NA�7!x���ԍO��&�:F��jb$Nt]��2�!<k}�ws6���%-�&�l�_�0=�qά��X�7;�1z�G�Ax���g�XX㕷ĸ6^@e�	jX��;��]��ʂЦw��W3)��7�����
�>��v�#@	�?�P�9��b 
��]�"���S�!\��7+�u{t2x����jU�&�-�:4nf;���E��#��X�?M����'9�R�ӄY�	IjC9tk��UN�����b������Z�2x�&���5�jwz}��{�����f�(��E/-���]�rFn�U'���(�ϐ�:F�9����5R�y�`zC`�����d��c��Ԩd�?o�?��#:s0����~��(��Rv�2�upIiӰ��l���#@Dh��PVp�U�x��G�HG<�3٫a���>��a���]�cA�C"��Z���=�#����{ ��n���V>'jSq�jUmiK��� ���,�Ʊ�?|P����U�T^�؉�+C�ۑ%�}����S�NW&_�
�6�.����h��G+�]����G1�*����sEXC�0Iی�=h	<�"�ݒ8�l���i�2��ɹ���c#c5?��6��*���Xe���Fiq�Rd�s�%�ӂ����Zk�7�w}���=Q?"��@NY��� ��԰��� ����Y'�q��ꅇ��U����'�w.��m������'�i���?���n	Z�O
�����FV�nX�A]T�&V����P��t粱8��.�8�����խ'��Fh�:��A(���"�C\���ʼn
$��~�j�ƒ���� �Y��Bs%N�=Ǖy���9�נ� �W`�lE���QW����Z-r_�k��+�r�=\����wn���D+�,J�����r�g�0Ҿ"�����	n�x9r^�����XD[{,�:��8���`�C�%��Xq��(Yټ���,�])���g��0p�OެdT����Pہ�{��/l���ik
u���X�8��������Zx\�J�(%q�P��
D�v�8�Z�4q
p_{��s�]�X+b��Gp�8���H��ᜂ��:��U��zx�y���`�����9�;@�&NnSl!���@�W�,��8Li���������ߔ�AO����tN��]%lр��_��r�.���~�/����R���J�G������WS�H�4|'����5�_'AB�.��܆����'���?5�=yT�Ҋ�v-iۋ5}n���k�����d���{u�$łC�S�nT�)f$����Lŋ���T��'
[�t0�ȭJJz�����i����d��0�,l֙��0���U���5���|s�-@���k/�i�D��f���oO�/l ٍz����&J6���Mܢ�-0�z$���q\)\�Z��=���^�`�	5�a�P8��|AZW���֥����w���#H��Y?%�j�2�H���m:I�h��'�&���'�[�W_П��W�b	v���1[��Sط���H�_` �\����U��P	2&h�|����q$�����b;�Z(*tw��~�N���th15ԕ��c����g��õF��P,��:붚<8e�@��%�����`}�F_g�8x���4[jG󶉈�8c	���"���Q0|����O��"i��Qcvy�b¡3�,s�:2�\�#M��92����.�������l����1�q�\4O��%Tݹ�z OKY�Y�ӛ�w]jV&�H@ߪ����إ~X�Yحr^�,�q������	Z���&�7�5k^"�AI���K3�v���D�9�{8�u�˼aFruL� .��(��M1jq̚�);�j|�/˃���:�wZ�k5#1��t��+ޛ�X˸w����p�z����	��r�)�)N������m���n�"����	��u��[��`rÝZ��k�@�IJ:z [It���m!;u�m�SM���m�,
�KJ1WIBռʃ�9���w��K�dely���I�^�����0�8o<��j@t�۔/g�������{>#�����1��)����������]�+)2�"�����pI];��C���սBb�e�^��
I��Œ�jE�x�(2|b3RGFgt��b@i����Y���;�/����0M9s�ҥ�p6"Kڵ�?�J�0b8.��S4@0��V���M~"�8��W�ik��D��Wt PE�8>��K} ��P0��x��C���A6�e�	D�#w�tN��_���}�3�*¦
1	/Z�6�����M��lW8�{�͒���D⠃a
+��'s)�6~�OAB/~�2p`��p,U�M����I�s��:S��-�������w������B�4o\�#g=��h�mg	�C�^ ��4�*#^��2Xw�lz��'��F���F��H���8J *-�6B����(��8W�ʬa�$�4t�}�#i�B����{P��t"6V4�E:���^v�͒�A��K!㬇���.\��(�yRh��:n]?�����W�4~Y��}�M�����XT�OBU�:&�ӒͭZO/}2u�؍/B^&,��)���%}���^��k2�,7�Ռ��<t�-�t4����0]9��S䗞v��5��@�߉ �\PW`V��Y�Cd�A�:!�/|pM�'}m��V���6���/�f��^�':��hg�E=1�촊7��� v� ��V/��$�+�{9/ڐ^z�	+|Z;N�r�}������+�,�S������7S� ���!XD�����l�P��	%�XKuS�"ښ|_p�O�az�F�%�t9'�Ū{�<X
��>W�;
mF�h7�����޺D�(�~�|�!�ɶ��O�F��?��ǼW_�(�N��	�w#��]qU�^�?)ܴ;ogo��s�8Cy49Cd�n�4���ϸ�f�����^�ݰ��m�ܱ���_%SE�~VE�s~�mk�b6�"f|��kc���ͥ�O�H�_c�����V�"�v�!�cnd�E�~"_&)A2L� �W,U*�M����?b6M����V�U�o�@�Ue�2��P�Я~~>�|�[��Z��<�l{n]p�:�g��r5��T���)i�/�w?�l-��W����� �Jc�,VْLk��!i�F�,��[����9�-��h���![]*v��a�����D��6�|�Vtf��'�|���� &���Eu+����γ�,�kY&DfGf�R�z?h_?�$L�%��ƌ�cYe������/�PKQC���n��'Car#���C��kP��	��{���a�2���}d��U}}��T���[��bN�p� J�e�р9��$�xO6�C~�=Ps0]�U+p��������������X*��D��̡���X�>J#zRi۳X�������Bsj.��M���P����9�Ӌ�&�brc�^7ױ�EϦ��� Y[2�ꋶD3Ӄ{uۘ+�H�����wgWj�&�&�Ǟ�����G��c*���c�W�<���-�Q��X��h�s�I<�O��M��z���{�7��bF��^]�	�����!��<ڦ�c�Y���b�;�W=c��!6A��s�g9\%��y8��Z�}6f���$���>dI,n+�) ��3�<8�����T֪�����" ���k-�o���Y�9���^¨틊E�M1��o���Z�w���PTN���D����Zܬ��Sy^����xV�̋+��n��6���+lF�����Ŝ������&�V�L�9�p�vj��%z��#��`>�,��X	�.n�o�Es0�Ho�[�%��}�f����ޣ��9�6o�v"jA��Jc[c��BQ��"R"����>����D�(e��e�	.�+5�_S�8nPH���'y����xIBv��$]��v�8�["�'?�U����?N ne�9��4>Ÿn��_�b�����>H��m֜�f�O�2:���.�±��Y�Aع��1Ǔ�r+�2{rv��r�1�*�r'?g⡼��k���@��L$i���$�.6%8b(!���^�:��KV�i䏦��ACG;b�,-��$LPr��W� �'����Vznl�撯'�U�v��X����G�?�?3sR�6�"R兮>�̄�Hͱĸ�l楈�TH��6�4���������o y�dS3`ٚ'���|���mW����}�8���em۾/�1DE$yLֻ:2��捲GO�P��b��.<���\b��41��$�$��y��v�P�A�I���WW��&zm1.�� t�Y�ɨfA�%�TW�<3U��!sR������L9L�����dѴ��;�>[XkźP�q�e%�-#z������G��'�V>���٨4��F�{`�ӁCE�����s����l�/b�w�� �@vz[P����Q�}�����U
�z�6���5-�N��ܿw��'V3K� s�z-m���Cm�7yf�=*��I)0L �'�*��q第D�g2<A��e�VX%q�,^ ���K2���p��U���K�̽S�h ��Ut�����؄u�����Q{�7�~oV�}�rBy�U�g�= ��I�^'��Y��Y��c-٥��L�OU
v�}�+z�R.+��D4&����Ϊ�=ș0ȇ�?��'�qF�̭W�d���g�AG�g�,Ι�!M�p��;���'&�@�,+6�� ���������}S[؎t����/t�k
�_�}x�$in?����[�3�eP�e�D��u�tD��?5
��)��9��%��~i����T3�PB�� �8��r���K�Le��^�r��x�?���E����r�}p'�]Ӹ�s���~ã�5���9Am�����L�$��<�dl��r����e�Ę��*��0�ٷU��XH���o�U�װ5[�T֧�ºj��\6�0$�S�͘���r��g�m3����5OS
�"1Mf��Y��y62�����@�ٲ�b�9������V�2m��D�y��)�N단A>rn(d���v4zJ5�����3jW?7���hG]���҂��`(0�ӮtǨˑYw��X	�ܰ0�)�2)Ύ�$�>ab�1�R�8D:e{�[�,YJ��
"��P�+���aM_��x)EyN-7t�O�G�>b�M� #���ؘ�!��_SӅz��^�cP�6�f68b��u]��_ ���\g��m��i�4;q��K�"���7��?&k9���&����9��F�?�U�h�ڤBt�ϖ�ͮ���۱z��4�_~��l��2Ak꟤[�[�,�����x�����[$	��Ɍ�g�椃mG�v���t	�b疪�c1���齦{n#�ٿ}�b���S�#��'�����L�O��#t��۳A�|�y ��jN�aͬ��Z�#hf��1 ԡ֢|Č\c�I9M؎�4�#�`cɁ��7-��r .�A�h���4�^�xjB���������3�!�[(!q�ׅ��Ҡ�U0*]m쐱O3�ƿ�S5�2����[` �d
�^⹔�j����0�����n���}��95Q?��A��Gk(����##���fM�>Q&�Rh�N�#Wqh3�D�w�:��Ʀ���;���;��g�P���o�Sߟcr����Su��fA`;���-�v���ʥIN�P(����2�2����O�M��h)�w��9W�st�0n,�Q�^��B���A<䋯��4uQRh�Ѯ��9��k���+���CPe#	���Ms��Mޭ��A��7L�Ò�7Tɵ���I��/�({�ӫe��q���>�/��I�^�J�`%/H��i�t�ʔ�+�dI���tX��]r��'aXi�CϺ����&����l�/��U� K� ������W��o��M�2
5�� Ӧ�x�S��vWr��q���E<��*�!�r�T�pUvJyk�Pk.���E�E&ls��kG1]j$]0j����w�Z��`���i��WӋ��	��H��q���k����HP��_�q0��N�q�4�/4u�]�\�#�^|���JT������iZ�Z�܆��"�Q-W����A�"�/|>�_-,�WgD��1U�g�O5��O�ŦB�8
�"�������WH�����]�����|龫K6��?]̲}9�
T	>9@9E�����b�~�M �LRQ���ڽ�t��.}�¼�U����,IW�PU��6��f�R��Ƚ����̪�H��$�E���_��3v����y�D�ܗ�d�����g�Η�;��L���1!D�(�Y1L�ڊ9�XS��UG0��0S�2�/ np2���#���'���3@��4�e!�G�`i��b���6��O_Y�@37�S�E`�o8��}����q�D	�PM�\�+F�����O.�t�������	�I9C`���)�B��<+y��0�Z'S���iH!��1�1��IV�h��Lppv�p34�R��2E�-�����OS����-BK1�
�rRT+� ������"���1X���H�_sϰ��v$�w�{`g%�/�����k�G1f�)�9^�էR��ʇ�1��)S.qƪ<�$]�!�wSɻU�:^�VJ�������'$ܶ5o�%R��r;�܈��~8�[�4�����ߴ h]������b@�yԐx����m��,ٺp3ֱin�@blqc��Ӿ/�����q�J,oT����ͬ�f*u��R�k��������HW6Qjb��,Ew�zA&����i�']ƅ�$�����
b��@�|o J��DU��R�p(�ѡOz����<j�{p7�&rp|�R6�"pP��2�>�j�Ž
�����ęN�9�n�ێ���o����,܀�0��RlQ�Z�j�t/�|�:v-�s!�T�&dd�>���2��Vk�ޖma��?����ۀC��	�ku���x�2�6�D?Hc7�����s���A��P���J Njُ�CTBOLV�E������dw�a�F����o��~����4��>MTc�v�hY^���A�0�k�ˣ%���[�Q�xgQwX���O���_JȐ��K�z��n'�^fd,�Js`M���=Lb�F�%^]Gb�v�y���^$!?�����P�A��%^5?�*�Ť�_n5�(���s<�m�9*��35`�7�Z0�WY��Gf��}"��?�}���U�8È7�=�`5��`Y߿;��ł8}��C��
����J\H�.�'���L^�����l"������%�E�U/'��%
���Z��9Ɖh!��X8N!�
j��h:J�ԭ\�G����+��&G�	�����Χ��X1W(�IE���r������%k�j�k>��\��/���ﳡ���4�dIR�R{q��2H�x�I�O4}ˢ`����+�PT�$�l=�TU������uޝ�,e��}?�`�@{Y��+���ub��RF�/d�+��{L�p����*S�S�ކ&n���@�n���L*�'��>���򮙂l3�돱���f�0k�#����b
���%<Y[��\O�����[��I��2�eX�l�F~��(��9+������u.tH8�.U�Jg�&
4M$L,0���Uض�Պ�'��w��.p�.~��� ςiL��H�q��$٪��`���B9P�l?Q�z�<����ۨ��p�(�r��V�����8($?��לk��a?�]�w�����x��8�e�^=&�.0W9wG�����Z��<�jV?^U��}.~1L�_8���N;Q�yQ��������ǸfgR����a��K��e�Zs��тi}�T*�e����wF[�\�=%с��plU�EM���/(wm+��V\e��8�����q���
˞�ؑ��/�l""����]�)yc�I�)��Cf��d)�56:��r�G첀�fbI
��u|\���;��{�6�s`P�O��u�is��Or�K�9�N(e`+d[����Bӑ�+yv�l�r����,<�ߎ$�x�$���A�B��re�=<���0C�W�9D���'������߶�@����L����ѧ�N�wVa��
�۴��~��*O�STT�^���<��8�Jg�~&�ER� Æ�ue��fdܟ�3qT�q���m�O��<Ty ��Y���a^~�*����^�]lE������~sNK���g-'�B�f��-}l��?�<Z\��oˊ�?o�����^>D���Tz`�7�C�QT5H�k�|����έ�i�v�ab]�U�I��Nn���m�uMQw������ �:"���Q�]ɝ��X��42f?����*�J�p,��d�\��;O��|A��"��?�������>�G��F��C�]�7?V�AӖu�1���I��m���?���/ϟ��wU�{������W<+Z4~Hg�z��SƏ�Hĕ�%m���:�D��f]�6��Ǉ�w^I/9Q�6�Њr̖~�n@��:��A��s���т���kG0j}>��ӺM�y��췲�����;�/ѭ�T�M�an���x�T�2�^��^�y�vnˤl��R"��W���?h��+5X$V�D�F�3m^8�֧=�H�h��7,9�~�'un�2���L'b��� I��[oz��䵘���%�(��"���s�B6�=-5`�85;�����?�%�A[��X��?T��(A�+��~o<��T+��G����Τf�W"J�/���D��JIzg��]��K>O��GQ�\/��M�<�L�z&�>�;��B�٘������7����˰�6��3�I�Qm��c�[)����� �4ܻd��WꜪro����뷐��2ʮ��0��1���h>r��0"���6���>�������s�α�/�C�hi?u7O�BF�a�"N3p`gq
��HS�En�tdr�����T�iH�mr�)���V"&tWDVe��Je[]\p���T�oƈ���f۳��l]�+�c�`7x��L_��vh�+�u����$f:G�O�I��YE�n@T���;9��;�ϺI��������s{���VƤS9�m�TH���p(��{�[�3���zشޝ_ �Q���-rd��e\�W)��{�����TL���x7,8;>�|%y��I��fK�h��)�r�
��  &:��p
��j� X�?��q�m���/��x/�`ck�kC@�J�V����ul��G!��+��y��v�]S昕$��v��SZ�Eè��3��!�e`��6�[�/e�+�V�"�}I�J�}�W1$Xxj��w�H��s�u�9����+	9�i]\p�.o��hW�����D�>w|`�3�~�لH��i��K�o��	T�����a������C;�;Z7����){(���P�Ugf:�\�S�]�I���e�-*i��iE���8ףw7���F)�E�#b�)z"%�=��I��8��B�'�� Ƹ�5��<�
Q��s8��AjhpS����-��4o9��b;Ǳ�m�evy_n���K樕���%$<�vf����o��g:�:߭c����U�w�'��s	cz<��&QN����?�7�
���3EyՄG�躞�2���@��|���l
�������j��5�Ca��u����g���s�IJv�6"�K�{̏��0z"�K�&�͕�~�p,	4}(o���!�� ���.�҂돩���[��DD���7�d�`>�et��1�h�0�I�VB �·E)��,�\�6��V`�S � ��LO cD̃$�tC�� ���v�$m�,�p���j�Л��qy���C?�/P/s��Dlt�=Z�}�(;�=큀/xgѐ5n�/��;���	�cܺ��b�E��4K!���D�m��_?M��<aCd��ww�HI���R̡lI��H�a���ܴ��x�����/=F�+d��#�����W��d!c
d��|�D�8$��ں��.<���,��:FW�nh����#�pYA�����Ԕ��Μ=�=!7�#�Do yv��j�r�zp�4��MİT�7�=�#סZ�^]cZ�g�v��XFt���d)fV��
��R,͓��ۻ��j�S"w����5f�}e�����v�诇�ex}H�dl�������桤�j���zM�@�5qں���E4�A�*��ƬJ|Nj�W��G����"��??��˚`���M8<i_L|�Nش���`CW��@���䋚�f�k�0�zie�cߕ��3����A������*�����u�~�^:qF�FA�e*�yn��N�-R�2U��<�)�"��Rӽ�v|m)�����+W!<߂4�*t���<B�BV���7���)���U2��v�Za9>��Vg��F�"d�Q�w�Mܤ�����x�f���Z������e�51��ò
w���y��2�8x�Q��0��x[�;�v�訓��:�`@����[��
H-��Ю���lܖ��.F����u����k}��2�hФ��p���+F��u���K ?�7��.��ma-�t�`V�Q��F��7�<t@��k{�i�����߷Ĵ��t������	��o��<�G� ���Ћ4 :0aț�]���3l$"�C����^ý}τd��S��~<�Q�m��%�Z�
�4�:��᝴����v���ԨG�J��#�y4�Z�-)���,�Z�._�bI�7�œ� $�yI�1���H�����B{
.ivH;;�J��9��@��,?S�������h}EP{�[�.1�m3&�~�
�z�h��wJ���ޏ'[�9�l�xH����0�g'����D�Y��!E���>̜�b�[9�"�x���>��1��-2~и��_dCH�$�h�|�	H�qP��G&�u���D�'�Y��])=���zg���^�W+0I��B�w����)�6i鍵���[����t�w���k����ƀ}2.@�;
M���d�/�<����}	��:��`����U���tq������8��!Z���y|S��~��[����١��f2:8[g�f���W_~�����Ŵo6�X4���qpQ`�Y�������q��?cO��$���!X��A]j��{����Dh+n=��I���;ݛ)�7�,�~Y��T�>���̞�ꉬԺ��6=�3��}]Wb�L�4�дC�.MI�a�iK�j��(�*���j�:Y�A�6�)o��.}�G���,�?n!ѭ%q��^�E[��QyX�M��z�Y]&x��JAv�h�Qq�Z�Ӹo<����z �F�C��	���D��܁,�;����5��3
�AR�Գ����+������)�O�;p�9K�����Z�����z�֦���>ϋ�vt����{�����d�M�ԕo��#��㉻L��dC�x��/�)��I*t
KX'�eU�@��<M�STvc�L,փ��K<�����`�|��2�x�s>�h3��(�	>,*�R�!KwY�9��ނ�����<Z��'L9�W6��P�tK��������4?�ZE����`x����^�'{���pu�jx�zPL��3�J�t�����9���+* �^?fb����?b�Ɋ��Qr&'��0w�;�M��!��j�f�/��m�����eY¸1�ԥ��|k�Wt�`uag��1�}�S/ъ�dM^�����(X�!��c��^�i9�%>���s��{
;����A�<p�7R�H���_��R+�j)o�:k��&FQ}={6x��_ �c���Y�͸��m�S��I�t�AY(~c/8dڠ�G�a�}�w^��C���&��8�u2 ��ܻ���oʞ@���4v�o2�c�S��up�l%AC�]���Z�9��ot�w�Z���08�E�BOq�N(7@����ⅼ��LK�q�����乼��φ�"zk�r�ߔ#���4�U詈��M�M�]���^�D�="�#hz���H���Pʟ2o�2ZmCd�*��G�P~}u)�zy�}�UE.��nl�~c\ʪ4�A ���x�T�!S�*󃪣]��;X�e�GE?�R�母(ɡ�e��U�4�׺����&j௴P{��-�As|���^�M�`��!{$
di�푞r�8��D�Z^������?��`!d�+v���|]��
w�J��0)6����R��P�|~¦WC�v
��7~�z�>�����9�
=�(E�����$�&�:�7-��9H�sfwβ�F.��؂�J���lx�=�:���
���J��2zص���i\z����z����;q�Gڤ��Pӓ�V,��o�׆46[ϼkQ{찇kmp�Dm���ą"+t�x�_�;���`c��A=�q6=���&�۝���ǣ�!>,j�~Ȝ�!F"W���V��,gB��y�Ҝ޲>��r�J|��hI#T:=.n�`���b��vMN��M�k�bh���E=^y
�:F�=Pp�P�؟��y�h�N.l;����p���d.�ڞ�N��.���U�=`n����wX��1�[8�CX1�ײX�v?� ���"e���f����X@�9ujr��BM@�)�뵲����[��M�;�逴��.r�֝��<����na�� 5H�{��O-��;���s��b���Iü��Ѿ� ���E�_�����.�`t�� �L��K�)~Cdx�`�,	J2 y��#G
�Y	P�|�G���ч)������ZjvDK-�m���O���0��G�Eٺ�$m�����ud�Ϋʐ��q6�q�p�U�O�|=#8ѐ"� �CNj�p��!��sG�ȶ.������x&JR t1
V]`���5a'+�̰�7S0~�����#'2�zM� ��{v���A���*mW%:�Ն�l��k�d�;�6e���~��ӆPGP��k�d�d�2p>w��e#d~VT�k��!��^���Z�S";+����y��n�Pא�o���ۿ����� �إaa%�`�V!s���� �#o9c�@e��k�S�㥺{m��~).rEh�ئ��A��`�{��-s�ͅ�f����b��\w�پ�M���(����[���#�s�*��_�m�%9G=��.	M��G�n�R(,� �:�'(JD`N�ci����{^�����ݔ-.J���
^���k&��_Yy�p,�Z� m�wh�R�$�_F+��&��)�ø!�r��k��|/�ٞ�6x�,Pnc��7˨�_7rD��^�}��P[@�b�L7���u"a[���D$���-~��Wd�2.tJ�|�<O��w]4R�7�$���K��Mv���_e:�%��)�t��KdRH�j�{j�R�n|�w�������P���f��� o��nG�h�R��pX"I��t�+�=�ԟo].sӞ���пO2��='��J1��)�Y�tkm��a��2�	���Ϙ�H�u~"�'Û�<�`�S�Ш���@.�!ErB��y��Y���Qw�Qa=�A��S�	�?�)e4��꾡z�	�}#8r����p~r��:�m��b���z��ѩa,����sA�/��`���%�z ��u��W�`3��Wg�;^���m��u܆I�^��12�:^���Ի��Q��n�,?��i���¶XtM�'��qN���):��i"ہ8F]x����*��"�&#ΥXZ�t���$�F|�~���������X<Г��-[<���q�k>��=�iL��S�h���;��pl�D��]�4�s;�(2b��C���]k�A
��$�䵈��leBs|�<���KVT��IIpl��B�����|8�Ѹ�v���0J^�-�՚*��c�B�}���V��<d"_�p!�a��<�lH����m���F�إ�'?�H����:6P�Z�":�jFڭ7�A���%A��#�\�p��2�#.��Ľ�!�3�H �0�AB�Y\����O($�j7l���3�&x��ɱ�A�ݹHN��E4������,֒Z4X�^D?�,��hD~HyK�3�5�(����޴Í�̽�m۵W`�>��q8��
z�tI�8���G���Aa��3�������H�F�)G��(Zt���|���l��
ҩ��\����.N�76�޻^�@�3е��(W$����a���9����J ���mY��&��h�����+���3�̵ք���o/�r~f����kפ({���e0�'��IM���cZ[�g�, ��ZT��������Σ1��3�L<�'��X����G<�S'\��\}�"%�o�C�'��	V 5_�����T_��	s�-bA@�aO�U�K��Mm/4(���Nv3�~UFma�1�S����?��HtPq=ԥ�<�ax�2jtrj����-9��"	wj�W��Ope0gל)XB��V �&;8��B����� �F�'�[��&j���5�8���y��̹q�]2|xy�$9���9���8M&�(U��;0�x�������0�nz:�Z�\�r(�V�K�F�k�Z�U����`�_D>mz;����=D��b�$.<�zeE��M����z�h����x���~[��$�;{��I.9g<K<҄��O��qo��:f��?'��|�-ѥ�+$� �� ��It0QLZ���!���ZY��uwv.+��%������@m*��g2�Y�\'jHC�*�H�[�϶j;~\�>D�o��������8h)>��ؑ�m/l��KVY�O���Z�F8q�j�
�Ѯ5"M��DD(*�jN�8-�~�p��UVQ��[�#3	$'/S,�&�'��L�NؓCJ��<�2��ϬÙ*lt Q�(|x��U�\-��}�n��ƌ���(,�"_o�[� ���>�	�3�&y�����H8$�ET�vb�a����Rʣ�h"�&��Hv�1?�uLЍ�<�}óӋ��Է�R�)sPƐd&�&y˫���T'�?N#� �����������?��>|�V�܈�tcu�SX(��NZ�x@ɥ6V՗B���bt_��1��!��,���Emߕ���eA��l��S*|�c+N�F��K{n(�5���.i�_�.��kc��=�P�ٍy�����F �n����VΥ%7�>3�����������"��c��H5��
�R���0ؓ^�f�o��� .j��~��,Cf�l{"cAWb� �ʇ��J_j1_��8��,ȉ��(S�)S��qp4�s-X0����Z�������e��v kC 2Y1��@�;Ƕ&�qґp�R��/y}VV
i�h%|��NB[�2�����/نaޖZ{Z.��)�9�l�rb�JlN�WI�����	��R�����J�/�+zf�^5��"�jqwAh�c��^�6W��N���|i�5Ĉ�V1��9|���۵�p9�,�T��:%�3xȹ�9S�.!`�����|��N��R��}V���x�u�bxn�"h��̻��)1R��P�II����01��8���z&�>�>�s}�8Y�Z �����>�_��-�� |�^g��YZV}��+��h�����lw�0a66B�vVo����'Wb�&�t�iW��f��H�Y�����
ͬ�E~F<J�0Z�͌p¸�'��	@$����a߃����BB�¬q��,�Uԛ�f�u�?T�昙����-U2�[�
��o:�֮�W�mt%���pL~�H�{)Ek7�۳�˙4-gkΉ����!*��
k���z��V+]��y(���/��o���i^�I@�
g�🌐�~': !^a���x�Ua�:�X^f�e��C��73�����A��_�O[��x/Ѭ�{,D8ۃ�����h�ApۄO�K�5�GǑt!�~"x�j��ohF�ş�M��>'LLe��e��:�r�T"j��1V������;m��/�U�:����y2�]<yi�b��<�[��S�����2��N���<��/�i�������*ϗz`QtwB��gމ���=5�e��Pd����&1�P��c��b����
��aM�ʥ��3wQ��Q��"�^�um-.OytZ� <��b�����u��F�}S�R�������-�q����b�aZ2��=�f�aqD�����>����X,�O��[������'
4�N�|xKD^�X������k���C��O�MP�[�o���Ě�:����2�-�%�ƈYq-�ͳldO(��Y��V�@}��e����T��-�A��*I����9��V����[���{�G��\}��`�K^���7jS��m%1Z��������a:�j4C�	h�΀����`���C!�p��1Ը% ������|�A�3<��!�]�_�m�-�"6������:���Z�+�e,�9��Hb��+�����G�b���YۣH'Q��(��9z��@Y����Kf�7=Ї�W���!i�g0d��?����Я��B��ߐ�Az<n�/ʉF�J���&4��<d�� b�Ӻ=�ۙ�(��TIb!�0�_�����nA��.ڐ7�P!*@*��p`�yi���C������M�W_��F7��
�3E�(
v������Rv���&]҃�ak��&Q��#�|�ܾ�xR�B�.U�d�e�:a�<�L3��/4'�Am�����O���
�!3C�W��K�Y��e\�
��Kw���'a�Ꟍ4F]d��ޫ�=Y��t�
�tY���sH�-�����O��x����U|�m���8��n���v�FvƖ1D����V:SN8�ed��QW��ϰ&����x��Ix�]mDg%pB�]��3:|L�Ei3JNΦY�$n������=�P[6.D��7"s���zu5$�b'��-�/���x�Rc0FGZ����s�Вx�B��2�O���r|xe2�,�ڎ֑���~\��ހQ�ރ�1"@��A},$kpc8I2�����(�A|tq��K
3�'=�ÆF�8$��v[!DTԩ�x��y�G���h�I]�Do5b#�B���"��o"�k�q0����?�lFdUV����s��(V�0�����e����.���*A�V�I5�j�݄�~.g$3�p���F�>/�}�Z��W�G�u ��F~�C1p �̯��F�� ԅ[k����Fb3%~4�:��@��i���z\ΓX�4E�K��M	t2��P(X �1�2���	xc?ㄐ��7�-�H��d#"Ԗ�3�<^U�̡\}�g}Vv�WWн��װ"���Iq���
% RL7�0�����#{���_n����]��Tv���*gc]��")�vx�D����3j��S�bH�%'O�)�Mq|��yL�I��z6���'�A�8!���S�Amy�1�����<j�
�A�H�I�^�ӣ}��_�b7�s��a��c`�k�?ǖ~���w�f�R���B�gw�0���Y��B~�U5٢';h�>TsO�լ�7��'��_,����p8:�Q�eee�';@A�)FU���~~�#l�&��D���y�v��6���tȢ$[dU@9�(.�,K����J�%���5�I��۱�7+\�����4PcY$�W��]6�����0aRHǈ���P�a`Ps�O�y�[sp�#�U_���t������4�����Y��ʝ�����q�5�����6gB$-��u+���k�`�0|=W�qċ&t=H>o�_ A-sߤl�/�;����u�Gz���Geg`6�Yb$Oq�=͸P*l�Z4��O�+y�����#_��8����l�?�m�����ҷ Q�?����<���E��F����hv����Z��j�b�*z�U�5�r���6-�۪�����{e���YP�\����L��D�Q����=������	��AD�Z������p y� ��X�7�ŝ	��"�%��������a1,$]��rYu<������Җ�U(t������mB7lb�+T9 �x�:[3�B, >�mǴ+#�&��B:9�4ey[s�g���� f�\>��lFȲ�FA<�Ď���6�)�0�+�1^�*�`�2A##�hTQ�[Lx ��e`%Á�G1��՛�*��@�-xN�N#�ɖ�(�.VC� Q7$6���D�G̀?	0 !�x_�0:Z�Kh�o���C���ې��o��cU@�����Wj�5_T�|G���N��+i�lY���1o��m3���!�aƝ�)�)�:�]_�%�G���v�}��c�y�������	ɚX?B�b!̝C�7\e~������ϧ�|3s���#~������ ���ɤ��N�V��{�`�>�!��ʡ�`������ď+���U@�$ �c��J��t�n�n|��>y�<��߁��G�+ԋ'��O��!`���T�W��T�]�-[�zOE���ş
ϛ���Ɨ��#b�[͠�f�??RTv�����T�/�Z'�C��dVYt�8(*I�.��"�/UƊZ��8jy9!�����nFw�.)8 �©�9�yri>�H�-GŉwD���eUƲ��g�z^@*�V����,�,&;O`|ș���'�И�� gE(�K?ȯr��A�&ӨWo�G�3S�\E5o��[������l��'�o�g�"���>+����J�z�=�E��U�P���!Ф0�&�B���=y�8�+�e��$!�	�_��弰�PĶ���97~Ū����7ˎ6,��A�ޛ�XV\��hI|�;#f� n��i���8�@e,p��@<U�?�5ZA�Г���z�2�$��2�4lY�%�'��A���L_"�������@a#�-�F��2rs��N��'i��QP��h�����*�p�ʓ�|뵮mL������l�o|���1}���DB�o��"L�sҔ5��c�+��O�W�/�'�2�e3�g�2w;ԝ��E�Z$b�U� AP���ะ~��n��Ҳ�id���
M-��ȕ�]V1r��UT����{��KL��!P�#5�3�*��������x殍�3��J��|�&Y@|;�2x�X�w7�V�堒���/z�F���7�*�i�&���Qdr¸\�'�	�T#q�a��02��%��}BT4�_ "�v��W���e�*�ZQ�i覈���D�p���n;t\7g7�~�j�d����}Q�"����S��J��o��6�,��.�k���ܕ,���ż)�"�TAff�갻̔��Y=Q�)#^��Z �d��L�ǽ%��f�D������sY7���ٙ��&���x?ێ<�7�q��͊���38��Q������ɠ�` �r��L~�n7��Z�N���n��9xS�ƖD���c\^��iE`b�ȫ��&�@v&�˚gG<&2�<�����ҭY�|~�Vx(>(���\�:(lq;���䇂o�
�oڽ_8dmgF6��&�Ӧ�#�܈�-�:�.C�������a"���󽊓e�Ad���^�Xܛ[��R'5Fgt������Č[��-�9��-���ej@��� ��&ʅ%���|tA&Z�1�5�6	�~r���B�Q���#Ԙ5l������Q�h;�ԃ(oQhUis� �����K|w�']�j�/H�uH���!�w�́�uF��X���I���Z���E���O�4�=1}PQT��񆻟���u�-%��l�YEm���j\ⵁ�Si?X���|6MX��]��ղ"JrK"ǘ.Dq��uWbTf�2|S �r^��P��2�}$�C�����ҜC�F	ҙ.���]͡l!⊢��ڷL� ��Q5nH禎��{#F�L��K���8���}?D_��J�j����J
r�A��)}L�� ���r��rbn|�nf�U1+��m����f-G`�^oM�3��K �d,&�\���̥�&�ҟ�t��&m�"��9�}���C���]�ub0��uYƉVm�}��S�q����'Slov�u�ǟ_��-o󭭮��c��r��b`k{1��Ӧ!q=E]Qø��ϦE����0�/H�t�2x��Aڕw6�\g��ǎ�5l-���#�3&a�3�X���� �����b��� f�'����/�IE�qp)r�՝�1Z[*!�a2A�yi�������(n�"�� _�Ђ���&mu(�����C�N3Ҽ5�J��+�(>�d����F�j'�r�����u�IZ6.%�g�E�)*��C��J�������f�cX�艣iN�n�Y�Y���{��y��߃6V�0�H'[�(S ����f����[Л������J�h{;<�c F$�t�⼋���i�6�h1+�ڼyhT�q�x��-|����B��ev�y�R" j{"ő�c����*_'������p�ʶ�+˖��}�J��v���l����S]�bV-�^ǧ?�e��%��l��\���i���F�^��sCo��9B���*���x���VC���s���g��a�j��%5|�m����\ ���6�i �g�0�{�=��PgT�y��Y�a�5��zq8<׋�l?���E���]�8�je|�E~��|�A�3��ގ�'�����-��d��v������� غ�PU�u�slzY'�H��������S�F{��غbE�T�@��ȃx��n�N�vP��>�Y~�LI� &29�5A�Գ���d�p�.Ⱦ�C��rX,�_Q��ޯb��JϚ���/�#�rJ>!�&SS�6_S )I;�O�o�7)��6:&W#���Y�� ܶ~�a�pK��,�a(���HXa1�X?�`f#���	��j��>
?Ջ��}pA�k�M�10PN���r���iCaZ`1�zb� $�HK�E⃈3ڷ%���Wl�`j��X��K�
ǖ��+܈����q#?��>/�����s�=b�j�L_�WQ����|JK��F8��x�;bD�L\�yW�Qvg{�]�mC�M W��w�:��L�3j��ô���QI.�1�<�Lh����Ï}��֏���K�G,��Z��n�tXՂ�8���S}���W�V�U �'�P̕/"b�3���Z6�2��e�Xl;�Uvz<Q6�b����,�g�����]�(��<�0l�sR�*-�?#��_~�.4�C P���WR�f�d���@@A�u�;��'9`x���gY�pD�7�r�����:����w�����=�hUs�*JG^+��1�!�Ⱥ˴�ˍ�GC�)��j:��꧗����f/�?k��o'�����_�_n뙜�/7�3��G$���{���ˠ�bA%�+9bQ
����*���sj��!�����sp����c��!9]W �rX��)���*�?��v�����%p��ac^�~���� �f���L��gq�q�^�2R�-k��OՆh'�E3���ק�hߔ�0�	��l.'�^��$��,��	d�8���cY�%�w-E���W��m�e'�J��a'Y��)�AV�C�Y�s��:NS�8�P�HM��/7�{��ű���h6q��"=�i�9{Zzg����H�)(�}NBv0)/��W3��#�9�ya���8�;���R���{+b�����{��/���^Ύ��׹����+�O�m���E��|x��$��g��i}�ݔb��^>V�`]:T����#����7K�3����H�5 ��_o���vX �}l_���ڡ�1w��ۺ���.��	�|Y\@��܈�j$�S���m��!���?̡ \C�.M�G�r��FԒ� �'��~� �>��م`��5�a��V�~�O�	�~�Gٯs6v붠=2m��4�=�q��CW�1}[��];P��4�[�����Sk�j��b����D����D՛9NU}ª�d����v�gk�x�:�ʡO𺿞 ��m��������)+�`�Υ:�Ae0��;�>x~s��d5���5E�ɨj�k�no���j}l�C�5Ob�i+�<H�\���&��^3V!�"e���%�a��ۜ�+Ofl]�2XsںO�9��˶��4�J3�aiL�O�;����ǦLR�y��$֥�_�D��Q��~�^&�	˧�'q�S\�����������G4P�'���U��#�1���w���f����ĵa���H�n/}~��Q�uo�Ɏݲ2���wV&�5w�>�7�+c��/���j$N�\i�j��U�k	��ئ��������myL���`���a�K�x-|�w`�O%m���,�+$�� Ǵ��Fo��#�U��:����5��?��0c�VC1^��_#	�j_8����t��-�uf�3"��\��,�=�T��'Cg�.?6�DBu��@�)��;�2}V��%F�4�6����wqp�|M������0~��6��	!�A���n���$y��K���7Y�u�9R� ��@?�g��tr>n�]v%�#��7�+��A� ��54ƚ���v����p���~�CpA_?	,�fB�C���~2������:9�fF�"�Lo;�>�9L�$Dw��k����x<�,H��1A4쮬�C��x����̻���ES[4�{� ���nX / �ZC��h��g��P�t�[Ԩ!NAf�_�Bڗٕ��%�Exh�	�y�r�WI�s�_Y�vƞ.[CAh�cW�mq�-gs�DB�dzD�LĆ�Ea�	��7%�%x���	�:N��E��v6����~�"�)�r�Xă�O����+d�i��cN�_^Ю�݅�_T��q��f�����+�Ctm)di��&�?\�%�:��19Y��TĖ@��oș��Zε~K��q&a'"Zjd^n�h;$�_!{Y�����Y�yF�~�K�!�Ɂ�xk�c�1ļtvlE�4aX�'�?��1�[��Ӣ�[P��Q\c��]�~�2|CQ����yA'�	�8���@q�S�PR��mX�F�:�[��}\MG-ID���] �2����W��QS+c��8x�U?�?����ξ%�g��CƄ�V��7w�B�3��m���`��y���B��2q{�z)����� �9\$s�]s�+	��v�)�S�g���P�]�<�ZqWA��Ά�ȳ�8wE�Ȍ�0�1.�����;ʢ����_�w�� w��$ѣ^� U�_����m��o1�wB�|�l��AaQa��d��:�s?f������{ZS[H#w|�/?G������r�yt(F�C��:yF��KY<�? g�|�5��@3@[�ů0���:���PQ|D� ˟��:c@��~��#V@G�����*_�gz� �{��T
���p�
T�((0z v��պ6����S[$r��r�+��m`/���V��O<k���H�q'鸦�9g�/��>fh���hqi#��^����g�C�Vto]��P�9�?TQ�[��۠D����j�g�'�,��"�.������dy`�N��$��l��#=]������<�H�mj�XK��&ԣ��U��;^�����Lw�jmS��яb�1F&��,'�z����;�O��|Yubp�w0�%kp��}��M<!^Tk���5E2��������rFt�3�
���B��?��DN� ��'�|�!}yj��f��,��[jL��i�{�7��,��#Դ �[xŢ5V��[C�A�#b��L�Bwhj<YڂE��������ANT��;��-�'�vLA_!�&�� �~x	��ԋB�����S�6�E+��l�GO�L��
;�[��-:>�}e��/�wOf�ܯM�x��q.0��e�-^KxLD����y"��6��\r�e�U���*������{qn/`�p���q
V�0�d
h�X3B�uo�釨X6��<]f6 A�Ã�/��5��t�%d���C�����æȍ����?�i1,���#�kM���Ү��Y���������NK?GB�X_s��s��-��]��+~��J�D31��g����P0�^(To�7�����ׯ�4Jȴ��u�-bs.¢YH>���^ߥN��I����tt��T=�7\�/V,�b��Pv��Ϩ
���ôX�Di�D�a��K5	�p�ñi����!M#HQC�6<"�,Y悰�ΐ������`�z�`d q�y����z?sX��kr:!E~RF�JR%P��D#"�@�iT*�b�d���0<���|Ϫ���\�fB7K�!�3ܠ���F�r���p��x���k�E�����4p9B���L}����8��ת���A9,��\έV�9j�5W%,TGN6��ӉS��R��e��m�]4��q��+���V�!�X��+S1��R��,o�w��j���>[&��x4��}�;L��.�,��7u������f������{|]{��\�E�S>��M|����*�[�FpN��F�'�	'�/�eըzi�S7���>xD�d��8L�54���Z0� 2��޸��6-21l囬^�]��	�@.��)N�}'$����Ș�#���ԧ��>薉�u��Ġt�36��@ �A@W��U$�����wM��P>�l��z�Z�1̲�\��Y��E�+;��~���4I��ފݡ�tF�:Ƹ���!t��^=��� �ׯ��@�럌I��q�O���#�Ø�gt�0G�\�mS�������F�*7�%kd�>D�Z���6Y�,F9 *�#�9r�(B�ڂ5	���t]�7UEI<�xj<ݑ[���^�1k}7��(�؀�ӽ��h}O92���Nv����{�zi221�g�L�ˬ@��*����K���LUNqj.4d-������_�ɶ\coF��m
)ڝoEl:Y��I���a�$����W�����]w}5�rsZ�ʫg^G�\����HN���F��=}CY�Is�6�{+cbS')�3��^z)(��U������9䫧��8�	���?��Y���UXs E�<�#�@�g�j��
T��Ek��`4(cH��y��_���0z�48:v	'�ք?�7 M�������I��S�d�E����_?� ���w��A^@���&��Q�I[�E����cH=�2�X��"�k���4[b<"������Pp��ᨂK���C�®�o�wP��Xh���G&�٭[����Ȳ|b$�Bͫ�{q����ϙ�3/����/�����`*&�ȆF�7}@x�!�I�w�<��4����e������6�F+�m�4F�	kj� �b40>H�(�~��p�����K�IH�(n~��5�b��0��hk����1��0�8\��}��=sF��R|��	pM�r�53����"�Lة� �e���Jb �_����@��4�>��A�����������Ү
���c�18M��,��r����\��F��ͭeϪ���G�\E�6�6��؏�~.�+����d&f�fm�o�f¨T�{�����_Ѧ2�W�	"H�gܭL�8)�CY�]e�!� (��M�%���慓�WLG2V�p�T,��u�w}������gi�ާR�}P ב�J	�'ׄ��L	S��6i�Q\a�`k������P��!��z�Zx0�~�2���M<���uEv��\돱À���O*@���E�/Js�@����+�Y��"�D�[}��쁣�p�u�ɬSF��pKUz��z��:�R/�%]�;a�	���0�^��瀝C������,R�y��()�V�'�g�öJ�ߠب������R�k��G�bE�bw�z��ò��6�3�LH7�����5Q�^g1��)�T|+���X�)G�ڨS���������UMi�VJ��9���f����MZ�^X��о1�ͭ����ڟ�_��ן���DPN[�[x�i�0�a�	��ǦG�A�x^��Hah^�S��ań�C��Lr(�
қ��]���tX7p\��!�����Q�AF'(5�j\��y��Ñ.ōA�:�)���x�H�̋��6���)�at�|j
�|�A,��gL�1|��+�p�n
~b��ۭ�x��9�c�tLY��e:X%*g���,�$�j�q�t>?۴�tB��K��d
�9uhvƨ�[��5�P�3������pg����E&7�����EwL7�|QM��f� �O�h
����WJ����w�����p ����8;Z�ȟ8�g2��ԋ�'�Lr�R_��h�T�����\	5R��bs*n�jM��^�圍e�V�8�͗�˾]�ֱg���k�����WN���	��f7C�X���_"MD���{;�+��g���W0����K-��UDQ�dklI�Im�1I�=�:з:����Y��g�wlHX�Јc,��L1 �p��X[>�|)4�!ꆹ4�Aw ��ן�m־A���7��4FJ���LH�#ѥ�@\��蜶q�hKǚZ\>�(��ysm���7d#�Mv�g��a�sg'��<Ԝ�&����w]����w�B��#�i��<������XS��wIz��-�-�8�U�3k��BR��u�{b@z�u
h�Q,����m�r�{;�;���̀�5�'��Ի�BuD���`[ؖI:�3��,h<�p"�ǛPMp�E�N��Oٶ}Cp�*�i����ȯ2�6��l�)M�ݓq�7�]DaLf�}�����I����$�.��!����``��!����Z͢���k�qF�LW�P"��ǧ���.�>�E�h(����YԶ����ۺ�w#~B�:�����G<�1G:{�bl$d�z�[�㨦��2����a�J��o=� ��撢��^��>|��:�u��s�Khc���ѷDN)���st��Hw�HJ�r����J���Rݲ�1���=,/���ba���Ȫ�� %9?������(�ẑƙd�M;����1�ٮ��rų�B��Ge����}`�;Y�>�x��]EZ�e��ɇ����k�Ф�@�`~w{LJ�� 4/�#�x[u��c�`!�nB��@�E��w(����w4=��`[� i��Fa��|Ţ���Vɦ�G��ƷJk7�\K� ���v����H��W�]]�H�r���ۊ׷\;N�����9P�\�`��3ݛ1�����0*#3\�Ǌ�G�/y��£��5)#��=g������H�\�Z��"k�����G�워j�%�<��u�Ż���:F���]Z.7�&Ԋ��`���GS�=Ǽ-�lQv��y2�>����}ﰶ�JO>�g�'O��~dNȆ2�n�K�:e�_�hfdrDE�˥`�.�Z;B�G����k�6Z�f��,uꋿ�P$�it&ԓcN�6���;�A�������U0�}"�t;@B�T��5ؕ1�;���M>�7���n�r8�V��%��R�����9����l@ݤ2As���Ԇ���xC��P��w�T
�gՆ)����׵�T(~�(Kz
��4�,��tal=��]�p�>R�"�����^L5�|r���B��J?��Һl��+�
���²�Pr��㫄�����_���8g�t������������d���؞�?e��_�]v3���|�c���Aܤ���I��p`SX}��\x���lK����|����� �ȣ��e�G?�/�l�D:c�_��*�4w N,x�Sp�
s�{n�詘���/V4�!O��~zA��ma���(�u*f��|�Ʊf}�sdUR�������E�9X�	��\�H�n���Ez�	d���7��j�2��}�Ԋy��h��]�5�����h'��?��_�0I���U�D���k��`�om��S���&u���z�n*S��~6b!�e>����IΓ�Ghۡ�KvF58��(pD�IO�8����f#�}�j9����-vz� �8j�*�C�=9�¾,���kn9�� 偉"��hW��/&2�@&��I�ϊK"�2�l������9�Q��rQo���4�|��4@Ң�0��c&���ͅ�v�����Lz�?����َA�%}��oCM~&�l=f�#�=7 �ҚQK�֚���Os��g��I��ԃ66� #���K�m�3y�&��Γh'G�����LD]�"� {���j��[�d�C@�����#�A�C�<
�M���Y��f������1(�Dir�T�[������8�h�ŗHj���"��(C��v������DM��~�KS�|�2�2M� w"�M�;b��+:��Z˒]G텔�����IY|U�n�T>H�V����t}�f#FcI��܏'
�J��H�5.%�U�hyI�0 �"�5��<&���0��^�D�F	�;��Ms��d�Z�s2���?����A�+��$M���l�=.��(*������o�dHw6H��� ����7{�p�T�|��;3[I��}ፈ��CNL?U"��K�q����+�S��)3:~��u0[�����&{E��m�B�*q&�$�	|�{;�M�Be�&��M!�T�)�|�����g��ɂֶ�L���\��E�07P���[0=?
�)�N�;�W�D��.�>��I@�d�fl9�4E�V�*N�<Ga�R��uE�i��k�ȫ�fbʴ�vXp������6j�g����/�nd%���[R�Y|�]q%<��Ђ�n���������LK������B��xa	��|B)7L		��
���JO	�߽���Ml�F`�r}��8%`i��>3�ȏs�/��*$���賜��	�%j�ޕ��S�Ԑ��������ԬyU�FE�^�O�~m�G��x�R�$�4�
� i�t׆�����η�iJFb@k��>�p�:�D���=�]�e*d�۴f�A�mo]'�ץ:��Xe�J��q�M�(
�5,E5��+_��^j_�T������#�4��\a0^M�Ğa»z.�!A
b�f���V�}�>j����N���Od��n@�<0��qP�� �$�eݢd�M���:y��O@�S�o���ͩ��I84�H`��E�q����櫧���6��֧<��;�(;]2���0箤���m���3M,Hd���$�{3�D�~Uñ&<?dB�d���z�B�-M�*�`����̥8�[��vo�a��%�&�z�\�3�P�&q�Ӆ��g�[Ч�e�ex�}ǻ�Xv��A��U�v���`
���JC�?ދL;�'9g@֝��Uf8� ?$T��dCJn$�nd"W'���B���H;����)�5jɓ�9"�\��]�OI�p�}7�M�N�ꞡ�Qع��\>�3�>�ܚ�7� MS�؝�����r-��hȬ�Hrc���l��]ij���&���{8�=�WK���ϫ[�t�B��SL0��OU��M�{��d*�(�s�x�%�z� 
��{yh�~��D�u���>��W/�Ig,�*mGKS�8��3�����W�`�V�p^����c���֭��-z��@�>��XR�1��߁Î�,P�g�4����qB�H�.��E ���k�o�i����h��M�w��\3Tjk�&#r�M?~�,:�������<��sZ��
0��/G�2�pz��5���,���� D�T���
�����ʪJ��*O���j�׌=�U�'f �5Y�3eKWǬ���
2��_��cj)�G�F�J��9�h;����7̅h���jDeŵL��2�I��m��`�����gk���C3M�֧al�ʘף�Ok�"#4:B��x�(b�fF��(t���%��mF%�{7�����-x�1�v�w�����rȜ��h�E��~�X���Bi���T��]�X���Nm����{��U�ԧG�dif#��:��c�[��$�8"M#�|[_�~��av�RU��j�����ɀv�O3DW�A�-��w���i��E����bb��Z1|�(�{��P'߶��]W ͬS4��2��BD �j_�8��Iz!>���E����e����P���:�}sx@��>���'�� �Z����+����t��>Z���\�8xxj�Ck�0��_��47ҵ_b�.f}�	�)�b��J9T��إpG��h��QX�4�ؐ�䑫y�'8�B".j7>R�Sr�~�:�Z��\ύQ�$���X��f輐�O�|4��*�26��(�ҧm][)<�^4�U����|d��84�Xv�k��$�0����\*H����y��5=�E��(<d����}�];���Oaϐ�$��^��i?���Fs�ܢ�8�ʟد�C*m�C�}��q�C~
L-q	<�̹f�3������>�_��]ε�����?�36e�f���Ǐ�=�R�4����p5�4Ί)O��j�b���%�䒟�m�E�@�Ҙ��W�-n�|����1eTծ�G]M�@e��u�ұ�� h�<�J ��E%����4,�!E�zp*�(u[�i�'t�8�(X��݁%����]�����O�/x��Ӳ�н1��6���ɕ	E�R�zЩ`���8?ܑ��+����}��+�ќa��ť��>�Gd��5�a��(�j��m=f�4�=��?b����C첼[�`$~G0�{<��U�A�@2(^�V*č	������r��A��t�k����$j@�p� ٻhL��Oh�}`�L�ok��dp�/,�������C�!t�tĲ�y���{Yi��)ʎj$i�]r9��Qe�;��?\�,uV,�WƖN�J�3�!��ʬgh���=�s3��j}{N����f\
�r7����,��yx���H#S��O�H���94.�E��>�t��fO#�IL���_>��i]�	׵�Yx[1jZe�,�����"�_�[�^S	�%��f��Cً5�+ߡ���ڠ�ϣ��+�V-9K;@/=�/�"^]T�P�]G��.׺}��g�]0^�e�`C�_��k�fO����Y�8g��Y� �
�=�yB���O6�dx�G��w;��q���4�w+���MMl㏎��F(9v>&���Bh󛽸X���}7�:$ 9�#����abqvV-9m���6r�`3�4NSV���~�K�rZ�v�2�>W�?��X�/Q$c� �ns:p.����XL2�fC;����u"^�M�e
\_ޟ�p�����8�~���F�$�*A����=f�d���MJ���	�ƴ�q`���I�q]L\鯍���I��_�)i�T� bs���hE�Cw���8b�n0A���3[�z�/�'^���g�H����U�Ö�csV��.���6�}�_K��f�hzz�JTc��ߎr��AI%���5�)'��i��F^�٘�O��<��q�<a����#>��|u�0�����K�Q@��O��Nb���ۉ��蒛�(.�.g+&=�W����U���1�&�`z.R	��+�!]�p�8�;_�Hk1��޺ُa�;� o�e^A���T����G.���v�~�wǶu<�wF���^n�γ�Gy��5���� of�v�o���a�!��{wv������2�������� �4�5�:,Fo)���ٗ,f*+���%Iņ��>%3����0�8^��`:QG�}y��(Y3�NĊց8"vo ���ux����[��9Z;��$|ނ�;���ɝd\<
�Wi���⥞�t$�We���ݠy%�*����x7w�*i1����f�q0i
�UO��F��`�N`�.�� 0&y�����:Z�Sb��5��*�.��٘DM����G0�FS5�w���18�:�ę��X����fe��JhW4���! p�M�	;�&���5R��������#T��[����8���DW��yw��1Ɵ�D�E|��ce���=��g��_����C amtd�V6�V|��������~��T�=�� t�s6v���d�(u$"�,�|cgl��h���a>��nͷ��6��Z7��G<�V�$���)�R�Ia�:O2���0mO�!�s�ۚ��Hv�K$����^=.��N.ṍOb�\1���Aw����B��+{��^()����
}�9�u:�/��P���� N̈́@Q�br{��\'T�����/�M1��B���y�Q��^T\`��<��E��(��H�ϐ��.V@+Tzf�#�w��Ξ?՜r�+i��i�KI@��Z��7��vqq��i7&&g�X�C�Ö�y�f������.sx��y����Fׅ5a�7d�Ҳ��7�:�B$ݎ%�����x'}1E�+�!@��ቲ���~P�)]����i��K�h)]�L�쯄����@32t)�TB���0��R�¨nwO�d�ч��@K#��Z@;ˬ�n��3�����VvQ��\P5��� jIӀ-�S�`"����uR���۰�ZoA�~T����T�	��>o?}ۛ �t:�\�V�h�}��ͣ\����s%�ui��R։�+1 ӕ٣i�m�]	Ў�Tf�z���(��M��\���O��'��L(��{� �&EVKc���]|�]���A��K��ð�]r�_�6�ʮ)H�[���/��e^���= n��w��f�i�1���ϡ�����I�?6y-�iup��$�82�x��#�Q��؋��Q��X����iD���ߤW[+�NMd��/V�`��hCr
��8~c?-u��� ��pl�+KT� ���Q_\�x��A�b�@�.����訃���=`"�����fj/J�P0]����U��II��{�F�ߛ�!��y��ʯ�!���.be�:�`B1�!�5V�\�I�o�<9I�G�U,�!/O6�(p[���nH_a�!���i�|��K�d�>~n�.��k	la|��/3{�iqv=Y㙮,C���G���V�	j\��JtU�G��� 9�6(A�Ә��� �8` Ǔ�=xe��%�Ǉn����xZ�7��L�.�U�P�Pȶ��hQ�-��F�Rx����^h�, �=��.��"_#��+8��.^�m���*��l��)��E�^� �����G�D�#�8�	����G����إ�������.�;�t�h]�z�q��y��:y���U	5�ƜZ�Ɏ��=��H,�Vu�|YfA=�"쨗3O",�x�J)%����+:hMP�K� ��Ũ�jIգ�O���5�+�Q�^ÿΕK�����D8�b�Br�D�;i�#��&��NxD؊��DT��p��2�e	E�323js�Ș�`i/���/�*��mAS(D��Ζ�p����p��s�`��ػ�<�g��y%�P��ǃ[;{JH)�;&s�\0���i�� \*\�D�$��P>�-����÷�Wg�{[u���<���<K7���/ȭ�Ldp��d��Z6�v=��q��Z���L��(���ox'�
��o����]������nPɉJ}@�c*�d�?`ҭ�g̹i*D)�_'P�wH����D�}��f4W�sԠ�Bm�&P�1����t�������S��Q�������u����jg�����;
˝|#m�c'��B~X�;���߆��V�i1DyT�HsZE�ǩ�����*���iO�����J\���%|:�昳z�9t��r`�a'�)S\ "r�ݤhz����Vٻ���4���c��q��ft,vs-չW�?��%k�1��o�W���&���a�joA*�JOm��<�C=�GӐ�X�i�o/)(ܚ�����k�G��q�H�| �D�R�\���#�j��9���z����3J�nM�o���=�ҧa�al>�{��9@8����9,($i)k������^䢧k��^ҵ��1��O9|�շZ����2�X���}�s��O�SS���>�o�[�0l�ѳ�����^�v��r��Q#Rr�Vʐ	�3:ߤ{UeUH��Sm3K���@��j�y.��'��E���v�(腸�O�2�o�;:B2�Ly�����ӅL�l5���A0�5I��%��ܨ��5�3��C؎�h�``եv�v~]K�b %���6IO/c�5�V���T�'�9��G��8�l3� g�i���s�c��K�ڥFQ�P&ފ�2h��!���C�KP��$Ѐ��N��=�u�\�ˋݿ�M���$��=;�m|��ϭ�D"|�v+�u��^M�`��:�ʧ�.Y�#5������x9 S���hxWf6F�n�ll$�4��ӛZeh%��:n�U�FS
�Aޑ�b��(1�j��Ѣ	ˉ�B��86p��a	� �Q�|�$����5�Ʌ��%��gHN)ql�민�Sߩ8�����Q��R�GU�������1Vn�ۿ���\��JI�6j�:�^��f�ad�Rխe��{��"6 yi_���\|EX�s@�eQ'�>�je��h���y���J�o��d�u��T��ڽ��n|\f;�Bof�V_=�r�����VCHG�V��볰q��9m�$28��K�k�����p璛�d����Ք÷��3���o�r�ߪ���z�0'�����E1$;l�\�Wګun�ߖ�|n�x��|�"�]��""/}}??��̑7�������s���J�4����8э��҈.e�(��\)}v�qK��0r�8X���`{K<�+�R�m��DSL
֭hW	C������wI蜬]s�?P�E�
��u ��q���4�0�& ��G�;4��.�gv�k^%v���}s�N��X!E�)�+��ޡcj�W(�x���L���*3X֔K�y��)��  ���NS����*�\�
��J����(�W��gˁ,�ƕ���'����fl�d�>R`Y���k{�)�|��0%�[x�.D��'[B�Zj��״�Dw��>�q �ꦉ�znn�H���Ю6m�M�RT�F!Ty��WX�'���k�����}��p�_X�;|�|�{}���3{g����'&�*�}e��|���Fh�sF�,^"  `c�:;~F��Rؚ�g�V�&m+k�Z�ҪM����3��B���LJl#��W��U����c�W-)L�P��d9�����?쵪	ӈO9C`/�:���Uy)8��n���7獩ƿ�N7H�I'���z?�"��Si�x&�T�2B�tyAd~\���RZ���
�39��j���w��5^�[�%��N�/q�2z��ޛ41O*�f���!q�X�˲E��ܻ7���3�b�������-�_���ı�\�7�����c�$ɟE�13���x征�l"L�H�w4`�?�pAE �[����L+�M0+�~)�;�˚u��^K%J!E;���g=�Ӽ.ӧ_sS�(y\�=��D���f[ia��������Ԉ�_�3�!SO��-�9E�OǚތZ$d����h������v�޽�#��͸7j ����k��d��Bdο�Z�5F�� Z�Ο�p�S]�6\�08�	�a��o�n����׍�K��Q>$}�ӂ���ENX}z"3��q��VgJ"�?�V��d�b���6/,EO�<+�3��hQ	�Sˌy(]�y�O<�Qcj~���m���u�	��������.X�0%��}[?�V6�Z�q�/�\���XH�����lk�^���<��o7$.[k�i{�o���5Z��Ti�%�L
�i���-�is��p���m��X�;�)
�+H�P&C�՞s��D����h����`����� a�%��X��M��[;
�I��#��HS�_�� ��n7��ץZ��u9B�X!��̃j�60S����P�j
�L^��/l[��R��:q_��D��S�6J���a�~+���Ή�Kp���wa�mӱ�3tB��
��Avܝ���͕͑x����ەo�w٭ ��;�r�ЬaǱ�ƚ��V���L�@b�y�ܫb���O���C̮� ��{�$;es�/_�/�<#��{��jl�Ο/���R��5�ԓ��O{�]�o:E?cE����"w�՗QU�* 	&�TdL�I��N	ѢV��l�~�*Q�Y�U���:�Q�2�\$�\�FQZz�wf�ߔg��a��ssGR���ÒO+�������A�k�/W�d�|!�U����mY��o�����\�_�+7��<s�^�u����(��l�@ k�	�"1��kA���3�R�2S�����uLE
��J��o	F8����pT�%o7(�JxqM���:8n߿#m��!.�3[Y=Af	 ��?��BÖI��C8͐k���K�YI2Y���8�(#�<:P�_Њ^����_A��,�3߃������"�hy�Q��.W�84j �Fe��)����Rǵ���$���� ub���hbF��J_:~Y�"d�ֹ�,�E��V�d�G㵤zVd.[�; �m�#�`oa𸭕=��]y�P�4�����ؽw�Mb��Tk��|;<�-��n��K���(��5d��K|�8�Or��͹�!���g�����N���O������\x=��]g���
�y��@&��o#W���K�@5
� r֝'��@V���(�O�<[�eEN5�Dc�>�z���V*��Nz��6����%�[�����^�]��~��ڣg��$�-�X�p���^!�}؇.)��%`���.��S���x�d����@�TT�Yds.F�0K��X�$���*��?��5�w�a�{i�ܡyI��s��˜��u��7��wխVUwL������״x�@��~��A�$�sJ8��g�����	^�{��'�MA��{�rhs���/�E�W�Y�J�gv)�1�+x\�<i~Rb�a�����8�ˣ�/c� ��Y�Q�Ձ'�ޛ:�	�O�yh��~���0����VB����g��E��ٌ^DD�8��JK�r�%b��]�S��?G7����|����D�2���+/ _��D�9�gJ�vAY7h ��j��)�>R�鬆_-�B}z0��B�/�m~�|�{�X��H~&\?��]�N�(f������1����I6�ڝ1�)9X��9j< �-U*�Kֳ��[��5C{�/.�}ӂ���C�����Ͼ�~ �����*6���g��|;τ]�$�B�j=��t6���0}-`��XB{q�"	[�}ԥ�I�  ���;�H11V:����o���v�����(%������e�d����-�`1�6�!�޿�����g�h4Z��!P��bbl4�2x#�hk��m������b�W�t��o�k�N��֫�\��F,0/(��@Q&�8����lGz�s��a��cn�1
0WO��I���,@6�NB�+]�y�4�U�5�쟡�S|�I���
�p��n�妾�L�󞷰"�\�u���՗��j$�=f��w����-��e�ӳ���M�q�b�@�7#<L�Q�o�p*+�svSd`��n��5�53�ױ���I+�X���;z7F���V�^O7>~I�d���v��қ�̰@���6�:F(̹O'VC�P��}<w���Xi)�Bj�
Ù�����.�]�����e?����H��Ι=k?�<|�}
�������~�)�`�5���$e��j�Ef��X_=4��ˌo�˶��4=���5�Y.!����d�wVC&!��	�6����~�.DaO=��	]~��cz.��{�J��sI�\A��
;����mKr?n`j�6v��=�l�q�Z��F��5(o�5g,8���^�q ��ڂ��7��XCi�yʐ��R�^���t �R��iS�b# r�j�H:ɰ�|W��������&�:�.O�ׇf�5�$&os�ںȏ���5�1��w9���sCz?�p ��h�=cmTI�"�+�->p��L.�/�K���q�#���^PA+�o@�,`:6T�`Y>��qy��l4w�'@粊��H�,�&6N�� �_Kx�� )�L�]��r��l�6��S~
�	���7���+H�:Z�D�����wph����fv'� ���2���q�����.���;T��K�nVт�u(��X8f\�P�=���<k�MR�5||�����$��ձ}�؞�,�?�D�yc�Z�2 L����u]0'9�2&��wP�>P?�{�GI/�D����-��fs@�)B��I�{Ff����;�tɽ��>���^��d��b�Ѷ�R%�k�^���4�������7tNB�pI>�]0p?)���Nf�&u�ʕFƄdV��슝�||7���Tl+�pz�6d�����V><��гp���J^�ɴ���qF��֕WmlLC�[��T8k5��+'2�8����RsO�/A�1&���*-�\�ǑC��5�B��d;lgS�����-R����Ϥ{�jC��W�1^}�i�待.�`�K5��rz���@r���)c��:ad]�p7F8p��C�'�-�C�_+�]Z�m���:US�.�̣$������"��m=�~d�\�W�uUs0�� J�9�N��T�Jv7�"�����IHe���ꏤ0���S��B�Z����sis�1y�/S�%s� �;~z(V�}�

;_�9g�5�������U�5yC:�h.���xhb����?�}iᠫ�g����oh(�pu�!�cao�B�3Q��b���L	$��L�6��Ŝ�O� �~��-�[Қ�M��z�مN��[�9y��6�W��O�Ʃ+%m�ބ�r�1q���\��ihK�}bY���N��X���Q.��Q�s<9h���ja��n[yN;Y����.��B�I���]�r�Q5Dj� V5Q	.a��ō1M�q+EŊ�K4��.J�'J5��C*�sY��m�{�c��0��9���.M5�3>�V:�D�ji/��7���Q�O�g�n���+����L����?�h�׽����~&Q$ܺ�CmxV�C�g���K��s�陱��H�[h�����4� �����w>K�<V�.D��ERZ�݉��i�O�V@���U�Ҍ�u�][a�L�$�FH�7�v����.`	�.���$���Qb���[�⌦�G�*j$�vU��]{l�$ Q�c]��۞�lcc+�s|�<�<������g��>}��5���о�6j+_���x��Ĥ���B����=�?�J7=B��j�n��~`��@��%�MC�ס#^�hC4+F5�&�k=�A���H\��
���?�ި�Z�����\���1��X�����m�<�)/�	G�aؕy���>0?�^Ҟ�G�����y؅��:p�1h)�f�OT!��Ng\����D7��V�A%xdU�.��̈h|��-�W�s��6�N�����Le�'��������g�b�	�|���> 䍫b�"�U'��p�'d<38�1��|�@�[���?�n#h�I�F���V���Rm̟��aʔ���vI9	�g�$��CT�
���bX�u�r�W|�Q�,����+׆��L����H}����#�jpz��Nѧ�N+��#��`�7W��"7[NO1�
��E��L{@��C��/���g��Uf�3"pp;��{`�l��k�rY�k���:��b��^߃�����T�5kT1Z�"g�߼)��v=�f6)\�A�9J^�$Q�c����Kl���	LR��i�sqo�d�p}W�w�;T�,�iY�}x27�����;����ǖ��c�\!U;��C�k�،�>i����{�/�S�('ѡ����8��|�TUn�6{r��
ތ4 j���{^Ty��+#cƚ~�@�E��͞[�W�p��;sx0��J��&����#�2��w�WL#Q&���E
�4|g�v?3�^��*��
���Zn��(��L�RS��A�9'�
��%��f.po��#jC��Հ��� ѕ�ӵ�o�V��;N������y�V�y=�^r||dG'3������b���t+��R��aBEM^� ���<NT�����v�����/�U���i!����-!UЌf����nq�k99쟄X��s�(�&^t. �]�� ��;E0��~?�(唞��;���d����m/�1\ �kKnE�;��ު�:]Mp�ӝS��	uרf�����W�h��������Qv,�5�$#�4-]��۝�d�G�,�XQ-3ily���6M"2��s�3�WCIK�*���d~��� �9벓;#��Y�~�F�l��j`�C8�)�6�׵�o��_B���O�,.�>���k8W�*lP>�WR�����#Oj,2'<B��@ EN��5��:@��`i�npK��raK>���!'�u.��-�,dr�K1�`��;P�.9��7����O�h�ĩ���7��I
n
g�$L���Z�vK��Z�\��|i��zs]ɞS*lq��i�+U����|	��&�[~P-jM"(A�,��9ȫY82ׯH�N�����.�,�仦�4�`��똏إ$EZl}��\P���=��^��1o���ړ��pё��_z��[.?��n�H���![�B2Y���Z�9��T��-�R��J(e�I�����:�']���7\����}J���$��X$�VU;�5����R��TA��/x8X�	�j�Ll�t<��)��N�s8�5�C��R1��=KI�x���~�ưqT{��	��Z��?'b�tq��8����YyN�3$�&��'�DPwg��U �� n��Wp�UZų2�6چO�8�!:���^S`i�v�Ca#�`�7P9q	��n�iS܏鉑���Fb3��٬_`� e��r��"���K\5B`��ks�����Hޑ��|��=��w3B�	'u敢t�X��qYu`D�5�ڿn���L����҂�^Z�k��b�䄵�u��cK��O��|�R �+�.aL��-�V
٧�в��$�$��|����.=c��8��4YQ��ĩXU�Z�K��y��Ġ�ۼ�+G!�1Vh�y�UV��4 ��5�D�<'�4b���*j�VeS��8�m�=�ca[)F��Rh�z���(�"B.fGÌ����aF	��%�Jq�v����i�)b�$��?�CQ�Z���H��/��I:`�x��WV�2�O��'�m�fT{ N�:E_!�u�RꝨ��x��� R��=r�n2{�y`�w���T����T�OByL��D�3��q*++$���
�[NseN=nA�@V��/Z�0��e�8�?WJ��z}X�|�"�}��'mIe��T΁e�/���o����zC�s�ŵ�`#ɨ�:�����g�Ԫl�$ے]���#rcA���E����Jh�7�+Dŗ�w�!�k�����ʇs�#��� f�1��'J0�bmR�@�'E
�:���MD
�\�
����qm7�1���z�͒�\ڜyC�r�����e]	���ڝw�n�|�`&"�?1��$r�	f>�W�s5��pG*+��+�u�5�,�+DP��KnJ�b9{s�Ў��)�?���9��<�G,���z��CY�� �S
��x6�"�!���.�v�xl�ds��W�$��l9���`�0�|�~��8#� Kf�R��s�Ѥ�[�X��q�5>9D�xp)b�ξL�bq�T|�qTߠ��Yxɓ�%�������R�no{c��T�rΖ���kj��f-ߗG�Z#@�Y�\#1�ŕL�ЫS�y�ZU�����>WP��ʳ���R�g�źrt:�s�ӗ��Ž�V%��n�a���~�(\}X=3VH�G��
̢q�B�ױE���֥?�MȲ�G ����ke �{�~���[?moT ws; �V�z4U��3�<�G�����b�<0��*amd����w
�������A��َ5;X`��%��ygy�ށ�R��պ�07`Y>EJ����5h�%�q_ց@��������|;��4�����ƀ����q�+�Y�p6�����m�NGM���he�\M�o9�;�D���x��7,����^��<J��8�W�I1��d��>��(�Duޯ���Ѷ��+�:׈�1b�˭z�u�ُ��Wirݱd�fH&}r���pu��n�R(�i��� 6�P��Z�*#���@
"Na�׳�1#�#�yc����Ӹ��)�f]Y5�[$��(��W�f1i�q�:)��,&H	�+�&����dR\Ꙥ��q��:��$V���k��s��Jw�S �G)ǧ��#����_΃L'��s*�v����}�|��)�c��ji��4:^}�WO$�]�$y������߬�/��,6��n�O��^w>l���v�s��{�u����T+&Y��o�c�l2=P�g�ҩ �x��,�_��k٪�*��K(�,����k�����N�j5�}�VOM)��s�����Ҭa_w�w5��[��zoJ��R���	�b����Z�tB�J�P"�Mַ��/�B�>V����B�r�CH��a��v�Ԇ�i�V�	�M��y�A	7~yt�����v��.�rp\�ZV�/ʯ�+{��
�IC%'2O��_��J�Q;my@4���b������*�f*^����T�?�b��	{�`}����8�D6�<�Ȇ���ײg������hm�H��5���B�ZXwa��P]@���ab��w8���CV�Z��'�%����'S�B�(���3�-/���}�x��%����{���4����aFIo�[��.wv����S��+G0��g��ԟA�o�g��}.?��oi�-9^aRF X�#f����%	e�=Qf�k(x��*[u6 �!��+��k`�����{�K-�RJ���ǋ0�N{Rm���^��������RěG�X/���b��냶t�
���t3/ V-��z��=��aZ�eN�,&����{[��a���e[�߰o:�`Z�Z/�=d������S�\��U��������.���9����Pn_߾��^��:��YS�ֿ���#�����y���a�d<���#���`�y����;2�������?S@���r��a~������<qǄ��T5.���v����</�Ѱb蜪3��Gu]J)o�QJ�*�q��@*�9��|w9Un�B���pgI�.X	4"`�M���N�3+CMt �ъ� T�s�q��a�v|;���D����G7����8���4s-�e
-)͌�.X���K2vd"d�8��e�T́Z�S����aiŒAN��!Zz�~�̯}�z�7�����7/��1!w�N�[�4��Uwh���ًQ�������1>R��Y���F<�M�]g/-F����F�G"��e׳B�{���*��;/�{T�_�
���(h��0O, �И�g;+�g����"���;���ZΧ��ZڰT�u�)���!�8��;���D�Fn����V弪�j4�f/���M�G�bbce�FL�O����bE6�~	���������48���ŎȌ$�}߭��1���o����.�N�A�)M2����Cu�yM±�*(��֠h�r^��h�1T�X�_ �kmf�(��	7�[U�!(Ie�g�F�x-]���!�t�L�]�I�@)�}�Ѩ����_��(���wtQ�#��]���le[�˚;]��j���y���Y�I멒ܓk�4~V*�d��6�	ď�"���:�E���m����b�!H�׷�nm�T~	��8�� 3�/�e�XL�k����h��#��R �ʊ���&Y	���n��^�#�a8g��D�Wp��Tz��d��g�D�c�?꠫�M)���Q��,e�v��F����<�O��><������7�V��:	ѡ{���rē�2$>+��uֆ�C�����e�������ި�q��M^����_�����P�E�Nn\U�����p�b{w;������pE��������� ��jMκ�����p���"1�>�k�B��ri9ס%Q�զ:��E�@������<�ʿC.r�m%��D�P?��`	�y��K���{���9lʆ��w4c�J��X�jz�g%�1"3O�K!ݲ���զ�U���U��)K_�ם^�+:��	|3���� ���):X7������'P0x���XUkW��G����ê�\��g27���"��~wj���~��s�SC�S���QZN��0a?��E�#���:�i;�6��õ|���ݏ�{�zJf�kYP���˒�b�~�B!�>5�k$&K����9�S$S<!�d��b��TYE:���~��nl$���X��s�$����Y�D� �3�O�������kg�{�ְ��>�������,<�Pn4)uN~~40Zڨe݅]��Bk���A�qw� �&�Χ��΀ݡ���ro��ZῬ8D�����X�}�K����n9�=5�� ����	R���1՞�,��]�h+g�{8)��b��2ǎ��vl�81H������Z��))�ެ��w�sLO��N$�.j����e�;VѾޟ�?�u|m��XV��F���T�9.�5���I��o��>.i�����~*��r���B�.J�(�+2��6�SU�M�4���L���^��j1y��m��w���&�yIy��ު/,:�`�D�$sږ��[�x�c���1�u����Z�݈� �
�WoK;k�*Y&�i���J�>�_O�<B�o{�DN�����J�Ck}^���!��Q��2�U��R.�k����!�<�M>���ǵ��,�j�|k¦�ZE�t�ZL��Y�Q|̯���A�I4ݬa4>��<�3��E��toT�9��;��ޟ�|��,Z�K[
�q�Goԣ=��(�e��oV�WH�K!��#�.�M����5�(�,Ȑ����kl̅�,�'���@����~6�7�r�����Zg�����Y}�o�/�+�G	�:R0��L�_����Ճ{���M\v-�3xcH�SX��җ/ �C����[Ǌ�ŭ�`��]�eHW\�%i)&�x{�B��:�*��`���f!�FJ�vN:�1�'�����zCdxȈ r-��LfJ�l��֖;�T!�a�dԧ�{�P�Ȫ΍߳Y[i,J:U�Q��o-y�d˻aJ�*T�Ϟ��\��Y0j�x�{<�2t���6V�� `u�྆z�W������2}>0?�}"T�����x�	�Z肋DVW�J���G�=i�����g,?cDM��Y��v WJ�3�u�B��x?^�F��:s��wS�,�I�]��A�V%�L9�)��qn����Zh�ƚ�f^/Q2�`�|A�ы�!n���G]Ϗ%뼴�&^8k������"{�p��Z~-�4H-�P
��Yn��bͶ�m�����)D� ���h��sڸ���	����l�^�KO��Y��3/��=��n�t��������1�R�ب�*L��*޽$5Y?"�[�wQ8�r�Ӫ#��$���X�"��`��{�r񕄵�AS���٠�����o�\���G�YmӐ��"�w!�G���3�n+<	���O���%�(/�z�O��G��D^�Zz��!���37Bh#�t��dJ��I��2������p dHL��0���X�b�.�cV�|����-b�d�`���)c����lB����8��q|Z��b:�v��p[{�xrD����<B^�Iy^�W����ڜMEM�(�_�s�PO��/A�S�m�qݶm��;�`^�������'�y})+�$=��(_ ��B����IVT<��ɿp{���Mv~��ͬ�X�l˂�3��-��E�,֩�(�����Ȳp�Hz_h�n��Vx�c(�x� �P�Șk5&���;����ὥ�@|�-� X�kȌ@*���)�@1���h8u�����׸�OUW(T�p�#�� �棯Koڢ��	U��	��?د4�/\���%�ɀ��EDI*H�����%>(SN�r�j5��@O��R��2����:�}D�i��T��޲2����Q�d�rp��#�8�8��s���Ӧ��JF��D��ԺqQSmE�K��[����Y�
2bK^z�K���ͨ�q8Z��|��]�EM�j]�~a	�yZ,R��U}k��+ʇ�֫(sڎt�=ȧ�91������+N�(��@o���uIj��q���g������V����\�Ѝ������v��vE�<(=��i:y��(���I��&��q&���ًy��|������,(K���L=a�h��t�
/^J����R�FS�"bܙ/�*�gjO�b,��y�ËC�h�P�g�f��.m��G�����Ѩ�Ü]"[u�h�cy�bK�cO7t#�3���rZ��R���t�4w�O��>l��>� av^_!�<ik��W�,µ����i1$q���Ǐ�� ��l*bhD3��RRC'�۴��V`J�����-Z���*%5�T��L�k��1��ϜC(�G軂���Ө�Ro{�,�쥳�׭���?9I�j���j�{V�J��{��v��&���d�o˥� a��9dZ;:����V��y<�b��4�Fx�����X7H�U��8"�����ɝ-�nm?�kJT2	;٫���a��>��:P��ZJ��g>T.|���h�/�]�����C�O�R( ��k��?���bb�*-�ē�P	�`�5���F��6A</�	��GQ��b#��xݼ�ҥhl]����`!w���#1�7>�E���o@y�B�Z��Ż��a'�S��g�ϐ{�����\lv�u@�+��ye�m��M�)���D�
dȸe�FmA����Qt�x������'iw�J0�>��ϥ��=��lց��&]����'��A?rfw����Ur��p'�߁�Y�����ҋl��i�կº����,ɭj�Җp�&ᯟ.w��X6��Ow�pP40.ef�F�^!28b@aW��6'~�\��uv�4O;�~���)�ޙ��]�}�-��g2r�����D�@eR�F�ܡL�# :f(�/��r���G ��e�������!��D��.p-i��T<>���a`쬧[�o�@Tu������ Q�;��Pf5��}�*�9I�n�y�i`D�X.R	�L�P�C ���m�J�~��LN?��!e)�[��8�+��g�9T��c
7�����+�𛆽"��8�@�dA�q�(8�͏�)�f���H�#�@@[�����A����U����F������_��2�kv���"��]�~�Ѵ,��eR{�I�Ę\�D#��}蒶 �*b�F�"�gܠ�q<�tK�#��_ˣǫ�۠���� 7d�Ҟ��-|��ѯ`%��C�J���0�Ӿ�ɔR���azN�d��h*,�;Q����S�A?+�S������y�8��\��qf[]^��4a��9f�H�?��I�i��ޑ��MT�<b�h���N�R������̣~���S�d�h��6X�R�_+ؔ��p�������ʈQ�fz���^����~�&v���F*����g�t*!ɝ~�ꅁ����(,t9!:���7��@��D��z��g�S��I��H)��#kT�0�N�M�*�6�Q��ͭ�L?օe���`��v͸�^�5@�ک��T�u��Xn;=�ug�+�m5����/H���ݦ7�cBd2��\DTz�����_'� ��_"�[�hi�P_ڰ4>�f�VN{(,AUb�P�{L�l��H_#��8��
k�iC'�@ԑ��آ�J*E%����婝|���\��AJs�-�ٓ�"|��8}�����W͂}L�d�$g�O����)杞oدr�6���y�w9$UADB+��	�/�)!���j���ǥ m����Uy�C*p7dY����-��p
�8�#����r��X3J�A%��cM��r.���z�4��UY�J���}���&F��L��@0�]��U6bI ��Q���Α��2D�J&�8G6��y�f�x�xi���u�뼖�� ��	��8�)R΂��jR�)�]�/%��m���ҫ��btރ��A�/���Y�6`����Mpz[H�Z},k��_�\�-�7�O��H�9^�O��8�#�1`6��OgS2�(D�/��u���ܚ��b#�uBv�R�<b5�Xْחi5��;�)�����E�6�M��U�A���#&��C�W�Hj�hxZE���~h����?[l���>p=���\b�g�q��w���/�lxv�%!�1r�Qt��+&n�[)����4?�?��\�1j�f+�PN�dP���,�T�-|2Gނ��ӆ;Y˭�A�� ��p�r/Qx���fՐ�����N/ uW@Rƚ�6��t\��ea�.�wѼ��t�饔�N����pyB$��f��Gj�d�!Ox��y��)�� N�@񈶟'D5�<�ǱX�
/�,Ow9=��؜��^\L����K�ؤ7re�쭊h}��;��0�	K%=(LuG5+���[]M�"��D=����.El:H�NC���(��Hu�<Wj���6�?�SR�fŵ=�+�I�u� �I�NtBd���b]	�p����<M���K~��0����&z�<��[�SffQ��R[>L�`#/yl�$��x���X[������.r؍y��w#����c֯��ӛT�[p��1�@�w5�JU ���1��M��ƽ��c&'���kb�a�o/�����%ov�[��Q��&T�v6cGosL@���[�B~D���(�Х�@�㋒��a�_�_97+Af���hp��}�h�!�DB0UdH1V�V�X�lR���C�TzfQ)�A���Հ�{�Q��y��:��;��|��;���s�L��<^��O %�GU��J��X�ж�!-��/��5 ��{/�ߓ2ɍ��L� ��G�`?��7�e��7V�lG)� �x�v�*�\$v��=D���������At���49T�F��^��Ҍ�o6�Ȃ5a$�d@j�n��q�脤#�#f�Q��άԽW.������@��+@)�I�'1�ihĖ2|�K��ҕ��:g1��H�~� =Q��ܻ1?\�uJ3��x�m[��4܍��Set�c����ߧ(���!��ĒɃ�,��`��vE�6ړ��̐U�7�J�B��)[t�Ӎ���"{�B���巂�Le���g�Qѻ�|����=�DfΙ��πВ�TH�	x�S�u=�$���I@��ִ���G�%?b�qR�����^�L�^��{��Ã�rt��K:2�{t���g��ߍ��*8��#gN��h����fK���t�TO�	�vv8�r�����*����}�q1����:ϵ���Fω2C�#%�|�*i��*ZU@�+oIZ��n����R�w��l@�.�o�����d���jv��������\^�/L��Z2VzO�TM>��rO:K��%�|��Kǻ�ǗըEn�%�iن�dk+�� ����!�m�����U	Lm�1����j%޻nG��%��z}�YaR3[���?T���_�$���d�C����!��6̆�90S�v:^�(�r~����K�Bs��)��a�a~��~�ޕ1�>�$�L�B�V�5ѣ�l%̿A*;r]�����q��rr\�H��8鱇*{"X/��M��Ӵ��*j���\ϥ1�����?E(Ń�^��Pf�4$�t���/�<��*]u���d5o���uU�e<�A!k�z6��\�TX�F�ְ�^!�6�hMo��D�΄p�"�!��ȸ�2�e�U�@#�?���C�S��q�꩹5H�P'm98�j���Հ�9�$Tg�~"i/�x���:��^��7jW@�j��-�{}v�̖�~˓r��y��l�l	j�MBEt<)��fY�t�]k��+r�y��V�����U�_�l����Q+�I�9K��o7��1r5g�/3)&[�$怢-��L���r�ؾp��l�Ź�d/r�C,J$��ç�={YmY�M��*p�6{&1]��'"Gz~U�����	*�9G%�J�m��=k�o9qI���:Q�~�����e��z��$����A��)B_͆<�u�Ռ�5sH���|���Dzq�f�����!m�jk���?��Y��B*�X�E���f>�L��[���-{��9��Q�}Z[��GD�����o���q�{��|���IC޺��Wr����o?7Ӊ��ߕ�z�Y�^�������-.H�V',��i�ήI�{������l9ϮL��X�n�����o�t���|�����0m�RP���D
���������d�_��V���ŢL�(aK�&+�������d�28�/�D��׎��6�
n�#���6��P�zJe�����aW�����S�+�͗d��?h�1�V	M!�pA秮~n�RqcWpă���˪T1?�ܼQ^������yT��/�Nq����:,S�9s@J��.�뾌�8&�n��8���Wy?(��a���)�ne��:�W����-�.�p�wST��j�Ս��fm�	�vچi�����'ef����	��H�n��@@����f���Gx����X��m�ݴ��q+�HW.	ѓS����|��#>�r�:Y� y5�����Z,aޏ�{fĿ�ł�K����
=�+p���8��e�*!��y!* �m��UbNs������fĲŁ�F~��8m�f�A!$~�� f5f�Z�o�]���|�mEu��y��s��7c���=��B�������ΔJ;Lx{
Z�)v�'a�ij�:(mx�3o���o���`�Eɫ,�
�Ԗ��VDR����5�HV��������Kә'-p�%��3!�rK�7_����8��2A���-��
a�ؔlF��G�)WnfD�~����_ˣ������4�ʱ��"��yB����Q��=� ���=�K���ji��M� �,���~�`/Ŕ�ȏ>eC��Ε�n�U�`f]U������/ 7S$(}��1R�̞Ϻ�_ej|D�TA"�ƴ��r2�e�6�jp�Nhgi����O|�>K��>�MC=�c��/K�<�ef��ϠC�r�1�Ũ7���D��or[;�1uw����VIN�Ԉf(���c��:H���G��L�#��NP��@04�Ve��v��ԍ���a��Թi�3���4���az���ӏ| ��G ��|P1�tZ:��I����V���g� .�P����
�I*9�pC�̭�&�CQ]����
Wݔ��v�C�p��G^�[ԑrQI���iK�")��ȉ�O���8�����w���k��v��fC�_���a��m��\���>ӟ	[�i7�����[��D��v�V �Z�������m���_��#��6���.�Qx�Y��ab�u-8#��ՌZ���N�d?��#͊jP�lͱe�������8q�0a�rA-���]�J���7஬�gm�2o�]�_tP�N��4�5��s��9W4.���(��C��x­�-r{��#2޾�Zټ���^�%�r��sВ5����]	Z��+�E���iV�hlK�)�A>	��J�^�m\���f�)6/F��+}���f(=�6�<�,o/O�r�ܭ���6j�ˑ�{x�5˓jmn��~*��ԏ%��d��Y�smF������v�v��ׯv�gK�t�B��;6b� q2�5/QJи��'������*Vz��W1_C��dq���4�o�>�SU�p�.wq��}�PIx�8�q��L�-*��b$|�V=_���Z�8H�~)����c+v����A���4u=_L�v�?k��$���
�B|��W��
gjk2�#����;�z{��sN��^xi�r�ؗ!�>��j���Aȫ*��Q���A�g	 �/�HH��=�D�J.����{"S=Xj���'@�K_?	H-��N��1��h2ћ�P���,P��h��r1�\�k2�w��|�M�.^�� } q�J��0��
lN�P�2aH��Rr��FB=����Mn�;@:�qb P��6[�����t۟����q�����$��A���BB���K�碌Ȍ��5E3~����C�Ze�y�2����H�;d�Լ�ކ(��⮿��KB��!^�ޯ�թ�p�$"(�������z:�U�w-���9v���c�KR� �2�o�k���9���s��UZٱ�	OS��Z�I�%�]����뎗DfȾ ���F˖�T��;�J�.{��Gcu3*�[z)�4�mu�{����{��Č� �i��GR�@�����q��P���U�ԍ5�!�
'A�Q(�8���f���t��t��1�x�t�Zb�%����]��h=7�!�,�92q��N降��}�롛J��:���9z���A�ޙ	�R�9_� 0��Y¦���^�g�|���ޘ�� �6���*����(�r>.)^4I�۠����,�o�
� ����CTb؋��Q� 0��P��5��e"�c�	C=�fb �BqGmT�(��w��Eٱ�-��UX���Q.��]d��G�r��k�I�9�P�ve%�ܼ�����+'D���!�qBul�����~�00�h��;-�y�+.��D[�N5��6I?4�l	��G�ֻ˕P�Xo�{<�d���~J��|�zɩo�r��w�b�-� ����,��^F�N~�#�l�<�H���p�����G�;��r|���"G�0[�agM{�o�tw�k�A��;�zG�)N<UYO&c�y�H�X�r�DY)�MIɐ�_k�u?�o׌c����[��c����
��fT�Y���@���JvF7�%B�P�U�30	��Am�U5}	1�ޖ�Q��٠b��ME�gH�C�981,7���@�T癯5�%���ݿ�w��\�%8�}+.���>�J&���k=P�Z_������{^\q��b��	yvj|{6Ky~���<�f��Z�9�O^��h��r�y�����T��Zw��}�w/�FkP(<=p���a��f�"��J��g��x9'�a�R>��F./�Zc�2T�Ox��̌�JN��m-	�.���5����"��:\p�9.�̑��3�}g��dL��I�&oeӄ=�FL�=^nҚ6����}yt����ա�8��;Q�����2�\h�ܓ:Cs�����0��p�ѭ~\�B��1��������?Sr>�<6t�s�8�>h=,�,n�v���Ig�Ǿe� �����0RxJ� �2~Rx�������t]�ݮ4�'��-c���.� �A�LJcu���5�T�|N��8�RA�p�v�t�Zp&>N�۫�g����;ΎVj��O�Ý/�3�"{��|�I�5䜆���G.���������Zs[`��b��{S�)�"��)&f"EIz��|K�d�ϑ샱���`򢓮�4^�=��s�0m��o��o|���Ǧ��g�z�@�6�sh�w��c�o���55��O_a,i �{�]�Bڙ��5C�1nI�x�I\}HpSX-�����%���x�#oY�$��h#� �S��$�8�e�+�*-C�[W��WzZ���^qSV�z��*bII'1GO�HZ�>����d9�
��a��"�o�����l�T�V��@	���p�?V[1tN���8��MS��E�3[�x��;9�N��R��VHy*�E��|Ե�������PcB��jv�Sҁb����&���K��%���D�j�͌U����~��,w�JGnu��]=�o7�3�YÇo�|���ō=�$G���w����E������D�� cD\�@&[5`��jS&�r���+q�܋J^��H��lF���@�t���SW}��JX���!�nY��m�Y���i�����u/�UQ�#A����x#�l4�,Fu�������@x�r�~z��!CA"h�0� 0��9r���FT����E�� �Q-��� PC�@
����A�@��&ܠsK��i!KOx����׻9.:�ٜ����0;2 �>/o�)D�b$�T"�{\e�7���t�V��WO,�ȃ�N\]���RH>�,F��n��/4=	�S�$�'�������m��HDG�_(�$%q�&�׿�'�zZ�����O���d�Cyt����%Ӎi,��/��-����i(�"Ψ)�L!7���*RA:(�k9��9��zO�x|ȁ��4;/ �=�3j�Z^	�EG�zü��e�1�^�	�\0ca�=�ow�﭅y����#p^ܞ��S������6�5�!x:������ ��Xk.��!�l%Pi�;$���r�R�E
-i��s#9���2�R��A�]0���I��U93g�/j��ʠ�2�bcj%�-�n8,�Cwϐ�2�@��;��6ItP����n��/g(���jp��ЍYM��L�h�B9��Z��]�W�{�h��8���I�R�Ǉ�C�տL�k��W���WՙAR��U����ئ�v���@���s �r�mc��w�VIi[�Y��[@B��i�}�ݾ��,m|"���,��u���ň��	��Z���&$y��e�@���0@�6<�qF@�U0_t*1�q�u�k=��ȑktˎ}Q�8�c#
�jL�FXeL�i��
�����z��s
Χ1���2IF����j�~���-�l�w��*|�83 �Y�ͻ$��Sî렓�C�ٟ���@9U������REk��U�2� �6��%�ՌlSS<~@v�L-��y�p�/G�����4�	���B]ܵ�%D*�Qu�j8r6~�N�r�T*.	fM�L2��L �x����/����c��)���xz^�&> �ʒܻ>Z�-@���d��b���s0�]-����(+���w�]��������=.�v��Q3�[Ǩ���U,�����mQ����*g'}n�͈��3��3��H#��:����S'�p�5�y�F���WӴ���i��Ԙ�OC��q�E�������v���1��9,|}�`M=^�����{��=��R���`�fȥ��,,׀�ղ�O�,��*�e��������]�4��i��N�)|xۈ���NZ�w~	�#)ي}�����M�*�3>�A�m�?�sp�&	�067�^��q6�w3D�E��S��T²��_��x�B�O�%Ғ`&�P�4]@r�n��� ���<?�R�Ƀf���� Z�������j8Y$;91�ӱ�^	����d�����
�	ӑAg�3�d�v��_�N�X�����00=�:��k'�4EW�%��	��n=n;�����r^gq.`��K���E���o�e�m���
1�FYˑx�:� ���$��p�~lR�D�-`�����m{D��B(E�,v��Qʓ[�'���������K�9�����u
�L>�>�V�i�͠��ώ���*�D~I�
��X&�������v��I�~����sѬ���y�����f�������:����Lپ.�֊K/�����%rxG���+Q���3�^+�%�{N�`��\(��`���k�>�AY�4��cP�%���i�ߖ��U�0N�H�2��t�(Qj׃E��Z/d�06M��%:��oM�F�%�d���V\��[�ʉ3�	����1�U<�E���Qj�����a�33�ҏ� r�)��������A&�7�]��
����\P���f�hP�������2P�jgt�1V��v�/HB�~�HI�k.O<�Y�C3eAD7溓B�M��KLs/��|��d����el��]�co"t�̹�;��UV܆7��Z�ғ p�6�# {9�4�TJI�x��-���/`PK+P��s.���"]U�㢱[m�Z$�>�Hz"���J�@����[%��Y=9�dE�	 X�b�n}{�e��`���$�� �&儁P��[=���Mޮ��E&�(�튾�hi�u&xB��|B��O��e'n���v� ]���^x�5gq��� ��{V��.-���Du���3���w�Q�_ݾ�;��S�Fm�mt5��0�)�$��qq�.�lV�d��*�SO  ����φ�V�Sq�X� �b��+�*����ϡ/莎Hp�#и׌��i�|���M���v��=��s���^�8�D�m>�(~��N�Z:�+�4�}J�{��(�]h�ى$}l���y2�j�j���l�r�pG�T���7I�܀<e�L�z����\×k��%�A!�r�tM�G!G�74�.ڸԒ���u�'�'���i����+מ���ͯ$U	�}�Ė��T�Pn�@�@UrB�P���Yr&(;��Ւ@�CQX���m��9�m��F�	0�)e�{�fq�19�ʣ�ε��mΚ�.]�2i~|��p��L;�%�	%�s}%��7��[��=��Ѯ��~��ߨJ��-��	���~?��Q�2���S�����ǝ� K�:wں�zm�>^��@�^���5�ʟ���܇��Bgc!��|���)q��ը��Ǻ�v*T��/m;��
���ڭK�����?s������9�8r���E�ݤH	ʦ�x�� �.��LhH ���me��ޛ�]|��Dy��rke��g��~��=[B?��\���SM �a���	�$D�R�����ؚ���T� �7��Y�h@����ݢGY��J��t�v�`�'�Jd���_�FY�	��mČ`c����rH��<�2Y�J> �)����n��k�^�zC,�h1��<dX��vd<G�"�
�w���e�U+b��٥��ٹK0q�)k�r =�����L멒�o�5�E���^Zht,�nҌ|�0p��Qs��_&�� ň�2��dm�wHE-�t�Sەr�M�!
����Լzo�2�m��@�KT!k�)^x9�>����w�o���ԥ=�ߓ�H4����qc��#-�B���h���L���8�$���}��7��86�l�����$��ׇ1K2Rc�����(�/�*��2���r�k��h�gB��C����0ɂ�vK��gf�����р�zE�=P��&�]Cʠ��8<#K���,_��k���%�kL�GD�Tiy:��d�~��rWI�~n9�K��n�X�<��-؎'˓ĹB�^�Ř�B����Tl^�k�������k���_=��6�3u(��[��w/(l:��鉻?2�H��R%�l�II�jӫ��i��}���.:��^�P����4l���7���D��h�Ht(aϋ�]�'`[�2���PP�~M�3�.k+m��7�+aʭvi���ԡh���x��(#U�w��T�~���N���5K�3���w���f
��x�P�����o�x��K���0l��ŏ�����vP����W�t���.3��9N'�ˢ�d@�߰��� Yh3ͣ*8Җܣ�Ѹv�k,��� ��g��A�_�}��5O<f]��Q�>�f�}����a�<߂���Xb+H�v"R�j-���S�]����"���Z$�K�k�e/XII���65<��Y⻽[5b����t%�9��Ϋ�7OB���+x=�ܗQ�����<	���0�V�o���aM�ݨ�c���S��w�Q��X�y�$iYx�aG3�WX��JK�,Xq}_9	K�3ƮSA@o�D��BK$��k-4����3���]�܏�q��dk��S��X�M1�M	����c񠣸���O��庸�Vm���m�&���U��m��n	j�9&�Gs��z�H��Qg�{�ӿ��Ξg��9����Ec���t��lv�_�?�*��@ιr��SO�����O��(,PL+H&��iRJj�j�ll��7?y�b��,KV���/�yR�wv`p��M7��"�RǀT���~��Ϊ���)侏V>�Ȭ�H]� ۸:��S�,6٫�`&T�L���J>jn
!��W��w�fHn�ys��V�9��L@��p�un܀�a?��MĤ����		.�0di�T@����Fv�!`�R�G6��[�sa$�%��>sN e�J&��x���>��6��#ϣ�m��n9>a�������ۈ�ߗ�뒛��qׅ"��������>����<��5oFD�_��KRC Z8k+�mA�M��!\��]��xS�I���_��u)ZR���z�dZyF*6K�.��LV�@�J���+�t��<�O�a�O�"�O��z���1Y��59TsA��k����N"����E�EѶ�=�Ѷ� �K��<$M����)�3T1��xʲ�Q�a�@�6�#cX�j���{oG��vt��BnwB�[6���v��X),�EU:Ql�/'�x֏_ʳ3a���<P�+�e�8.����/���Ю��������#L�z�q<�B���*:�əS���ԟ�Qx)�@�Wߏ�'�(�|L�%?|�������w����9���)Qt����Ӎp>g�v¶�qÞ�����{��S����s�s�'�T�',�[qf��bo���. ���:?��������9<SI9bWӄ��\������5Z��-��/�t�	w�9�F���L����Ҿ��P�0L{0����1Wo��ը�<�oӄЕ��߂��<r�}=�������5V�d�z	L���!#?E����XF��v��K/<U)p^�u,����˘�D�-���scx3X���(�f����V*�r�/=��4Ҡe��LJ6V)�`��Hݡ���`+�e�
� ����Z�DH��sd��ܢ��#�8�#r��xT֌�y��H��4g���/�\fr���Q�2p-l8l�����f��-�i�ܮK:u����;�ksR�
�E���@�&���4�w�_kM�O��c�1|Ic�Xf�>ˑ��1� Ɲ�$�t�/ns�7z���S]��b�9r> �|�d%H_�k��ͽV��~��<�JA��%}��.����E>;,i�c�����%��+v�Zx̳�j����*�k�S�8�0D�ӍL�"H�M	���9��:��'	�4�Q��!�9�����@Ђ��S���+�Qw�#Y�\��Ȱ5~7�A�h����2���4�U͖'Ua��£�F����E����g��S.Z��f�N���0Bz�1�����&/���J�<���0���N��� m�H>حp��-��N�-��^��fRr6'�8����TҧIY��]�ل=ΜM�����(��#���­����@M{2jƃj$�^A�TO����pp|���x�Џ}!S��(�S��=�*�PQ�"ȉNL�3���/��̯JJp�VC�L��	��!'!����d�!�_������h�>x�7q��h;�����qF�8b�Q<O֕M�������Ɠt�)#�Ʋ/��;�"|&}�'���[k���.t�j���m%v�"Rm﯒XR%6{����䊷O)�P�����"���x"�Uf����=��"�Ny�)5]�g��� ��et��@r�6Cs� 7�]Ȟ�I-�OT��9�@�f4R�n�5)i{���dS:�Z�m�2�P�S��9d;ɴ��[�s�1�S��R7��M���:Դ�{�� Ohݦ`h��S[�ɽ�
�w����'¦�a_�<�7BQ{Mx�Yn�r���3^��%]��/6(���	�(��8��A���.������n�س���|�����K�JL*�����:=,�IY͢�'PE�oQ�2�;!�zJO�O<�Dm~��8�V���p�Ă�`�ĝ���=v��i�)W|��Vw=6�	5���X���U��xhS�bq�P��ӭ���WH�L�'Kdٽ.�O��\�����s���;�޷~�R��:X|�u\���篿6���k��(�
�O���X�ć�
���o�E~~���6�{x��-7&�=��
0`ʶн����d�����$�!���Y��+l�F�!�����d�@���d�s3/�N��M�;꺰�}�B@>�G�u۴N��cB߽JA���/Kx9{ư��q�]�nhU���g��I�ʨu^t���	��ª��?�  �6N�ј9�_�-l
�Ј���P�.\+BSs����D�Zi�ڗt&oX}��%�)/��ǮGVd%<1i!��qcfR�"�ڿ�l��2BC�J-�p�e1�Z��E����{vW�ʫ��|�½�;�ÏJ��VpI}��_�h� I�)����کMǬ4 =��u3��P�������5QG��>�X�1�P���a5~F�H�L�����3�Z���{�w�-��{毵Ž��a��fD�Tg��3��bz�h�OL�rJ�N�+5��
}����k|!�m�b�u#6LV7�Q��<�����&�)�Kʖ,=O�LGΝ�\%��:�
4���AJ1�\5,����r�َr`��{���£�	˙�q��o��ҏ��T���+�o�µ���
�t)�UU.�q�v�DĿ�~7�0f_�.����!zt���r�U�X��<Yd��e������q+���Y��FRFTf���" �D�"lɕ���}Q@'���H*{O���&	��o��y���V:H>�n���Mg$im�e���s'�_�X��Mys�dGQ`��W�UF�h�>�6��4�:Z�e�d�+�`y��zM��Xխ��+C�b�u���YC�wT����Rɛ�x��B����٘��2����`xBE�R�;S��<�����{
�#� S�<q�GB���~Ѻ��
y���k����H3!;����*���aEw1�Tu��NՐW��_�q;�0�I�X�g=��Ky�&gw�-�a�V�Lv:�BY!uVn�e���?t�ʭǅBI���7�о}N#�2���[�E��&v�a��!�?&�(ڕc�r�<z��r�}~}2\������|O�[�T��� �ee��s0}i��Kq�x�}�[���R"��e�� `P��B�:P�/H���quv\�g[�p����p�"%ɩ�hLUI��"�3��Թ��~�ר���Ǆ�{zD��8��jb���1�����h����%�?���H�����/�D���9�d��fY�C��Uw\罣�vf�������6s,zL�m ����NEq:,���u��t��V�;Ax�y�]:q����5����ձE|�WƢo�ߠ�(������?���DZu/Z!a��!9�^�<��.��O]��,�%~)���	���^�T��I�%/�N��Dq��
u؁s����S*A��/������IlN	��e��Q-�#{nE�I�Yp9W{�U�eI����Hc�/ػ��,ͭ1f�X�ӑ�n%P�cY����������F����2�Z�	F���NH��UÇG`�nz7�_��p.<d9�xA�9�Ҝ/pK(c�^3�<���7	_��A7QS�M玩ˬa��A��eT���,����1��v�_A�גj��p[�KbE{(Xl�Ͷ�0�VP���� �B�6�K�u����d,����Ӑu����r����)P�7X�Z���q`ƾVT�{�a��f��yk�
g�k#��EDL�a�{Vf���F��۵j�����{�ܦ��N�PfɅJI�m}N)�
8���};8�~�`.E)�K��f����&gqn/�>RV�p�Z\��¬puz��o����z
PN��\���a���a��	L'�t?������3��;���2����܊��dp0'\�&�r�]�N��Z��#�z%��KO��E�v�o;�2I�)��F��tM�F��e6
��?	3���$9^�bfj~�}>jX��.0�����Z~�*�s��F�M!�K?��"��1ERnp2Q$��<Q�zH��,yה&��A����|�@���������Ⲳ�J9/l�Ρ�6`��8s|�29Y/^�2��p��@�|z��Vا� ��y�w.��O@0��b�)ћ�)t�%i\]�!�-����zh��/<wRS�����Q����a� �ot>h��L�N�09Q"�?��?&$����]�@�L�o�ڼ�q�@��n��ED�?F�`�k���o��EV���/���L�5�^�b��[��*�\x��d~k8Їj�0���:�|�Z0����962�e���wϟ�8! `$��t3�V
�5�I�q�:��n��ձ��6.�:{-b�6")���զ�����Ln��D
e�VC��9��e���67��Ǻ=�)Xɻ�ŷO_�3r$5t��s����n@&e��E3�J�'��pI��]�
�`2��+V� 1������G�h-��/V����#�CE�3@�Ǒ���ph�g���[|�c�?����c.#��3����� ڲO.�>���?����L�c2x�}�Z���8��q^/���^�z���M����HGk&�_Ip>|j�~���#`_}r��詃�����q�HeQfp|���sz�3?�[��v�ֵB+7�-�i?ʿ�8�u�N�w~c���n݃����G��x�\���}B�-�����1T�$f� �ʢ�il�޶�ף)[Q�n遧Y9�R'Mng��ك*� x4�8���Ɣ9V����)d�DݯG�<��� |�Bv0q�i��L	�U�>�~lpwR���������Q��Ε����A��۱�/�����FD��J�i[��X��C�A3e�''�3���ÚVx��d��[gE� ���ePA�.v����k[�tU2��;x�Z��V��*.
��Z�<�%�n���L�x�qW�m7i;�{
2�@y��c}���B�6�Ӂ��|Y�l�k���2�|�E���j�������m�C���@�c;����	N�O����#�ɞ�<n�n��t]ڋ>7m8��SX�Vq@5*	�y��C��^��yTŹ5uC��Ҝ�Q�]�]0�_��y���%���O����)��o�J�,:P���
}�zl0����nҶ���n�!�����P\��@d�� ^�s�Q� �j��Ҹ�T=4j<L *<� <HJ��ړ��W[-�����^���<�S���u81@&	2�ɚ)i	�6�2���눮|(Bx�	Z�}ōs������)�z\������Sl��$���X���7���T���o4˪�[캴��*=��-�Z�O��1\���.�)��)���6��\]9
��u#�ժ������̙�bX�m�3���j���wAsN�<�r��f���tjK!i�4��y����U���5ظ�
'����q�˓E0
�s����s�a�!/����=��i{C�j�Jpyg��)��L�>
nh�Ҁ�u�Q�	ׁ�j(�Z��z5��{��UiPv ē�p,3��H�0�b�ݭ���j{��H��O���b���!�R��>��f�^��̴���˥]��Ј^���g�W�����
�Z���S����=Z�1�KV��>�L�����r�
��3tؚJ��6��!�����~l����w� �
�'�6?�q�6l-n-�����:R�c�j95����*`���6@�3(@�N��j���D-i�~"��׽�Ӥ�8�p���.�{pm� M&�7���-��l��wff��تB}���E�k�.�/upv��1��v������T��������.�Y��������#b����������֭%fava����z-m��L�+%Ѹ5�w����ESN�0rR�*�x�H�Lm=��>��:jg�KV��xG�Z�Ԅ*?v~��(��<�tPb�	;+��j�mS]Y&�!$?'�ZD��tDq��똁C�9��M��Q|?o!�2�4�?��X�\�ExkhsQ��&�E�&��c�*;�RcMfv��;��>y6���@�Fd ��������T���K[YΉ"n�[�T�ޕ��p������� E^�Ʊ5��i�o�d��������?��$�7�>8\bמ]y���,W�>�0�mV�bP�yM�9q��	��a)�2Rۊ[�ٗ>!�* �n�/W�;#�?����3>0�Nf.�%�m��6��c���ޚ���,��:�<����9ЕY~"��%c}(Q'�|����򌇪�bv�'j\���&h�.��D�p�2��t��أM#�Ѹ�J�����I��&�oU���ci�]g��PD��i�v$�:1�N0��}b1=\�x���	�9�k"E�̡>Em��V��ޯ�0i����=�u����`����H8�]/��!�[�t���XհS�y֦�+1�8��z�J�,�V ��XJ�'��	\ѷ���2����{?���dC�wڠ������@�^�6R���>�hC�U�x3�X_�d�}@>QD���0��a�HF������ W�5eѝ��׾���ޓ<vǚ���]W9T�?�p��j"�c��_��2���j��K�d��lVv�pP��R�>���!U�{��Q;�f-]5.o]"�.���H�"6��.��VƇ�ݹ_�8J=��T.�w�s,�~u�q�ֻ8��F���W���5�(xvCr�Ǒ9�ʈ���/��t��Z7��`_�l��)���M�ZIrʟ�yg~��������6­X{�4-q�uү���=���ق�;@q-ľ^��L��2��lrr��x����K�q
��u�ɦ�t���f։��$vX(��D]�sfU�RX4m�V�R�v+%m���,�\��c�s�8�;���?5��Ti�޵'`��	%{�r��M5����x��Ӓ�H�o\�����ca���qM�b�/NRlw)yx�QNV���&v1��  'A��+­�+��<��>;��R3��]x?}�ن�I��ؾ��s�Ӛ��\Ȫ,Q>��;���Et8,SЙ��x�7����'Q^=����C
��cE�av�3��X��y��B5�w�x�	�J��z��rɂ�h��稰	��Fl+��g��	��"L�49A�ƭ�(��}5��8�j�۔{$ˍ-q�syP�c�F:ј�5L�)��L5K�s�.z'CΙ]Gnx��;cB۸�Vf� �L�Y�q�e�뤲�vgt�"%H ����';"�ǟ���߫���sO����u�{�u
h�d���p/( <�g��B��Kp���������_ Z��fs L{�Z|L�LV���y�q�`p�dL��s���z��vRݠ"�&�rptX�Ξ_��8s�Y"�5N=�v<���v/
�ʨ[�I �)��	�Z��J��`a���u�ΰ�|C��+����qO(q�8,=�l���\�:�|�}*-��w�0�A*����j,��uȲ���U��wGO	<�Fԯ�J���>X��*!�k +�?F�\�^b�ä`0�X��:�%�	
��h�����9�}�ҿ�L�p�q��lZae"^�W��n�6������F�$=h�O���:R�)�L���7V����C�� � ���ܗD����sa��%Pd�m�	���y�J���/^�:�j�ZWZ��v�b-�N4ޢ�M�x
-����$�>�F*��)��}���H�Ժ�3�y���g����>�9Ǆ����!�C'M�?�V4
G��uF��iȤzj�Vn�{�&�`N�SKbru��)8��
+>N�4�rq�U����7�i���2���Z�Ϛӯ^{K��ä��.#=��찱�����y[��:���h*�J�::��٢� D���Ң|	êk����Bj��/t)��Pe�ud���˞�����8�c!�����0"�ˊ�T���=����
H�(����6���� ;V�������;��K�����=K8��/�*5}�_�u�X� ط�ɒ�~YM�Qv�S�F�ZZ�W}P��G�2�Z��k�ǋryoG�����p����+<�:�ŵɭ����3���q
�u��^nPtC�۠�=3��3�A�$�Y�-}��0��z�s�tX�����
#g��=)����_��׾%η!"C�}	�Ɍ�ꠏ�"�܎�G*A�o��¢��Gpsa��*Os�b�����U5��q�S�g�������Anҙ��`^���O�lQ\"��!E~!�8�en ��}ݓA0����	�v���%4���8m��e�'Rvڿ�f;�NO��(����Lem4Ս�0��K�+�&ai��TE�]BU4�� �H� �<���
VЭ`J{��U  u?cA�t���d$M~b���ޕm�V�bw����ji��|r��2�=)�������W\s�M�K�����!]"XOsf�F�u�Y�: ��m�'ޚLVr�7I^������P�\W	qG=���9X���������	l�홺ha��ed�-��#�loGޤ���C.I�0'n��p
��n�@Ly��~+&�(�����S/@�O'1��3�ڭ2qqd�m�\�)ӷ!�|n"2�w�Ft�X*F)${��-Ο�M�f���0H�����a;�;[.��h�>�P�[~F�'��'��؈YlJ�ж�8��x�[Z�C��+����ȇh<�'�0�Mɶ�<vv��I���?�Ȏ2�jD��#���~�I㫅��N����VvG`�r	��̀6M�����2)��[���::�8>l��",Jl�!�h>u�hA`:�`�)�Wg�����ꇙ�$�(�Ře�nڦ��|�T�}����Y��ӸHZ�!�ɨ���G�ދwt�68�.��6uG�����)�h� ��[I�<�עȎ�쾟�9:R����I��=��Dr6�	]����%.�e@�GF�;(��vN�h<Z}lޫ�/��t�� ���)���=�Ɣ��C��_rx��>�!w�N�}�[	?tRAH^Q��J�0��UV\�G�9�-�� �*PE��"�,+W��M"j�ц��s�mD��?����R��)r�ӈ� �@o�o���ӭ��sG�����X։b��5�+�,�Dw����Ge��D�pⶕn���U~t|�x�\�B����ák����+�"��4�+�pixB�6F��σ�w�����(���q�s���}��h8���eƘ�~�ӱe�{h�7X�T�y�Cz��zG��).*�� �"����K	cTU�D��M"�*�/��E�r=,?5pUr{T��I� V�~��L��jP��B�8#���\�t��T �	�F�0��.o��A�"CR��(1x	��Di�pD��!WKW �x�m�*�=+���F3s@�l�oC�`�'�B�Q�^�,��o�77d���bmn����k��x�WNz���m��b|���;2f$fc�8BϬJ�*0��W�R�V�0c�evn������I���$a2�D����+NP�b�>�����u뛍1/���h�T�dF3D���	'�rX�zm3\8`@eK��,8І��d'>���X��lN�p�]@��b?���X^�=h/+'�|?����a`��kk�_
o�'ǻ0,��𻖄��K��x�Rs������  �%ۛ_YI�����]h�	���,�|��z�ڲ��"��~��~Ƹ�)��]��}��À~����1�H��q�#Wn������u�1W��>7�����?Da���h������d����G��U�Oٷ�������P�D�p��~���p�I����_���BkJ��߉�|�r<e@�D��y(�C�靯G��Q1��>���IT ��!�������:���Դ|x;c�Ah�HXs)pB�O&��[��0n�ȗ�Ƣ�!�����3�L����TS^��D�؇���,&�R�%ԯ�+�ٌ���t��CS�hG�˙uW4�w�`�]��l)g�EbTYҜG6��f��㮍#��߁�f������*'��T��l����֊Œ�_���S�����
��\ */;i���NM7Gnޢ��nqqT�b񫻓!�!M"��F lc*E���C����]]{�1M�h9kKu�e��aއ��9,����!��.5��ӞD�A;�\Q!%	'���g<����<�'���-��U���r�//�d �,/�j4�m]CzC�3�d�OAB��X��g�s�*�݁L�on���G ��\.�ϲR-���!<���IW�lL�{��A:4^��Q�I�\@�̯��$�,I�Q��HW3�G=�kMȴ�q%�Dcp�4-EN�9k1��W�8�$��Pt��&ט�_3�ߨ��*$��?�
��Y��ja�F�㖮 �.���h^LU�<��L��M�N��0��px:E����lu6�r�Q�[���f���	��8m��avSF���S�*UYz4�s���׸i�;� ã�}���2��-,��A\�1ܢ4墪+������D��z4���5O��`�����b/=�DJR�҇�vP%Ir��������9 ҚGZt'�Wf8�"���}��
�^i��]л�D8<��D��V�g.����o�tH>����_�T>�z��_���8"\����x�d켗r�0`/R�`��8d����I������h�S�|��p���Ew�N�Vɂ�x$B�q�A61���:>�7l�&�	>��E��Iǘ�HL��z�к������,(V����_�݉D�rDĶ+��	��+<�Z���:vd<Qߓ4z��h�#���<E�P�U�G_����E�g��h�M���A��Uޣ	�'�Ļ?���x<HLy;�i�׌K�).�<��\o$G�Ɇ�Ռ��IG�sHk36ݗ�ǰ�M�_��/;�����%Szg"���d%
�~��2s�ƨߢ��Ż�d��C���h#��}>~ Īďq9�HW(S �������}8Q�S����T>���D�>��&BE���i�07��J2A.��;(�-���	�V0�+i��_�J�{��l����`�F$� xal�����T� .�,�B��	{�F])8;�~9��;�p�����c�2kw�u�����kzڪ-��y��ѩ��5�Jn,*Ɲ4�����x�|�����!�Đ���)�6RJ�ӹp��ėzk7�f��z�>�ꌊ\܃H�f��}b]���<��p�����~(@�R��Y/"�<�\�e�s�y� Ā��n��T�w]_�&=#w�Ğ����]�0K�T���xI�(���7�2��W�i����n���[������G�[>Ø:ؕ�=��6��(3������E#^߽jf�=���j<�6���+R*h�x�R��VnS�}�y�&M���0Х�,���I��8�xi��Q�g�:(HK)����s���+8�
C��?.����\�_)G���H	��Qh�s�^�k<O;;��߿o�*)�����%|�x&���*���ř�Xge*�>S���+J�
�9��`;�l��_d#�ȝO��v���u�F(��8��V	i'�s��`4*ڻ����'�Μ3�a"s�9�X8�����Ϊ2���4���"�m ���$��8}�2�X��8p`ǫ��sH�ǴH�䘭Ε�`�rI4�?�?����R2)�`�﹛�7Y��x�J��C$��_.y���ڸ�1�T�~����ecQlo�^���o�_{�rvf����S��D�qNTZCQ,`�0��psm��h����@B�c������t�|QK z�1���=�0O�3�o�����70�r⃮1|�`2c�^V��e�y�q��!�Uū�7ڇ�(�By��wQ�+W��� ��An��B-i��aeq�ю�˞�����d�lgF�+�,������<�a��P��ɧ1�v��xG�[��AN[�����+�<ϧ�R�pe<$ϯ���M�}�<��X��9�KdF���b��1!�A#
1ȨEi�;Lu�P��)#�N5��[6W%���狂�tW��4�o���ډ/�о�R�J�C�y���O�K IT�0�^ҭ�4!$�S��k�3V渹X�D�j��O쏁3���`�#�������&f1��G	����,Q�&��� ��q�A�¶rB��a��`�-�wl�ڸ�1�W�VP��?GC���k�b ������W(K&y���i�3�x]oSIS=K�W/�Q�kV��Z��3���ʩu�3]�QS�9H��kߔ���l��� �ld�Ɔ��D����L4�Zl �6��"���{�E���7�ՠ�
T��Y��/4G����	�3(_�t¼k�)V���<>�a�у���s|$�y-B�U�N�ѐ4o��4?"���_�D����l��\cl�k7��
џ5n�}^̏'O����̏�����\bJ�*2��+NĘ�)�:]d��b���}S�N�3�{��B�J���>YMг�׉�M -�*,@�ɪ����[_d�C��Kc� `�����~bP�Vz��4os�-]&( .GF3�2�P�^�n��n�׸Ο�F������gJ�,}λ�M�����\N��+�7�+�9�∶�;^ZM~ힹ4�l��\j<3@��S�Gi���{{l �z�}�.�.Rޣ���:�w��`s�.m+�F� r٥�:n���9s�
�8�����͂�؇�;\B���D�F��M�lWa���I���io����pQ�l=%Da�yŜ��|�C�9D'u]<}��.�J"��TB5�����ʲ��T�m#WIv�"zE�Lc����)��תr�(�*���07����lm��:B$*%gd?���Ϸ��4���n,ud^

���3/xu�f��{~�q?��#H�	�;�sв/�Dj˺O�c�}��3A��1���D�|�8�n�(��`ԍ��1��NI�Bn��%�n\�YК�]m��$"L�wr@Pb�m
�)G0v�p`T��5+��6�II{�>Q"�B��gɹ�H���4zOvܡ����X7ѵt��Mx�o�[���r� �0���g��1�R�"9�W����Q����}>�Qb����d�iGG1f���D�db�S���7���$+>1@��!��@�*�����<�K;�)��4%C�o�U�}�I�"M��u���E�a��W�z�G�]&v.��GE�����^B�ve�\K����RZ؍����>Uv[��1�A�I��	+@��ലӗ�{̼�U�z�I�8E3��l���~��W�^Wq�m���.�AV�VA�/m���Jj�>��guk_��d|>�
�\+���o�(%B��A��>�L�ަ!�~2'�=�N�5W���[7vVr9h�߈��|F?5�+��1�yk[p�?��)P�`:�=��N�9�����уܮ� ���Aql��joXq�$��,��*�8!�MN�r�A�d��y����[|�	�R�7y���v�3f���0�ݼm��<�N���Q�v��&����2E��~�i.�\ZC�N��(��5�_ U0$d�R
e�BMr��d�(`$���U�ۋ��_Pk���=�m�,�����X6�PR�����^x�і����<�ͤ}z[�#ͱ1�|���u�D�ZB�3I�X2g�JV���I[�\-C0��p��Q�K����I�s���/؊�����	J\U�"���H��Z�o����[��$�%��&�p膘�^{���T��o�&����L���X��9I�:�h�l=�\~�y��v��v]_��P0��Ţ� Q=]闻c!E\�>�n'�J�]�2d-����~U �6,,��mZŇz���eM܊��6��#�W��0<�a���%O
�`Cc��e{��áۋ��tK��U.�ϕ�qSOc�������������SF��vUޒ�w6?�X<A�Z�,�Ts䰶[��gQ�_]�w7�#(V�j���3�G���W�W\"��\;Ȫ�����G+�CpHL��Tg�UB��ld���9q3��U���.L�<-��%����v	~���J�.��1"�-7��T�-��	#��Y]�?�]*y���>/N_ϵֿ�R]\��NpO�t��GR����	=��/���$��y=?1���p�/)�pp���N��yZXa�Z�E��:�i��6lE���Z�����i�eݞ��3��.�Ue����� 9R�jN���7���yn��Ei�]g�%���K���:��ET.ك��s���B�FP-�{uI$+ٱ��[�U汞؀��O�X�z&$0Fj,8i��Z��`c9�
V*曩U-���ex�55X����棜� \}>K�S�|{��>o�QRC)��'$8�Ǎ,�����&�oSs��H	$kz��^���^�ek�أ�k%5���#O�%y�C"ao��d��eq��z!x�J��y.�X�U/�C�����6��yc��U!m�U^�������fݺ���#{�p�	��Y�"[�&�5r�j�M�k2�/-k#��ǘn/�O�yd�6��wb����ӯ��P�S�{�@Y�����T���F�"�U Vuj4���5�d����5H�f� �ko��>��t1�� I����B��-�S>͇��)x��PBRӱ�K<�=�-�V�x����g]4 b�j�z�l��+
����0I(��=���z��8�ls" E���j,?�-��v��Pa���ڿ��Q�H��nr�>s�y�pv.��)�q?�у�5/_"�tX�;�X�G�bX���a�V/@���PKI����.�-��p=��V��(��/����Ye�ڭ� �I!��TI�����\����{�7�L
���M����Dd�<�0W���$rwa�TKE�Uxh����J�ߖS����		A�N��In��|1��Z0���;�$�}����qS`������(�l^f�r�|�xN�K���ִ4���Ӎ�ˤ����1�;�G�i@9�~HJaT2�Ln�H�Yh�R�a��-���ѡ�[�m�Q[�;����e�}�0�����N�m�Q_�v�����,���:��FL!^
�Q|7������;�q��&�s�5��<i<,�B#нB��Ƭu�!Jâ?�`Ɇ������#ya�ުS�CO	�0�����U3m�rz�曆�%8���Kd]Gk�C2K���[2���\0�K���ءe�>�x[��M"�Z���8�n�umi�i/l��V�cߗ�׊�x��i�-{��9".��Cݘ��&"�����l�Ȳ/mq�e!A����W���/�@$����$F�郒��'�W1�T�Z�%�~�r6$C�Lm���R%f�
I�+57��Kz8=��ʺ�HXY��@<�.Fp�Nb���̓�l�d9X�_���:��!U��\�1D������5��o����h������؝�T6s��P]�X�.�΍�繋�@�'�v�[=0���A�wj���
�tۋO��2FOծ�����YUߧXO#��2�O��Us얅8����i�`'�Kk�y41P�@�k�������D�I��t�C��CC;�J��q"^�5���Q�}\iu�z �3iD�.ۨ{��V�+���w�|%mcԊ��i%/���U��#4B�_���N�	�Ӵ��֨�� "tjy���]���?�| ��g�P�B��|R�����!#��9N����5�k�v��+�bM�S�8�w���&jfH�_��������Y�l7�.�� 7�'��3�N�2I[��"���{_����Y�t��x�03�$��r!cp�~|����W0LRGx�?Щ��hD����/Qh_W�!b ����C݈�2\���YG�����db�������Dk�@>R�\nҮvf��p�,�&���� l[,��Ӄ�/��-i�ok�af��W5�a�4�2�?[M,����.�0������j:u���y�yw	�?�_.����#s�2��V7|��E�`b�}���%��M�2� T���}F�H�&5���:�H���f����� 8��g-3�tbD%�M}�\�8%`��ߋIh�����k��t鱚����ޜ(� k���
����WW��֌�Θ!�pл�]���V+C�8��!h eNҷ���ۣsWh4S�];�s)W�@�r֑�� �R3�Ģ0u�r};#(����Ts\�z�Xɛ��>��C���g`@E�m�{V�`_�&�̇��ؐ&��Z�9�Uޖj�c��n����h��0[Q����$�tQ=(1���}�Ooۤ2���S-����0K�6N��񱻆����ά(�ޡ���� ?9
���<A}��}�X/S�>ό��I��3"ӘT���2�c�?�p�#��h��kps��{���1��7V\���4���q����HV�˛__9��S��gV�U���m��Z�v����b4ߣ�q��ݎ�����ߗ��5����l�d�-;�(�f}�z[Ҡ{�[W�M9]�&?�ސ���0����b��6u�ھ�v��}9v	�R�5u�E�o|��X�O�Nv��8I�!b��g��9��u�H��.�m�5���
�b.�R�5�93��e1�%V�q'~��St�r)���*�6�o[���u"װ��,��w��>N��>��ձ �k���6I�
C[@�U�39l��Q\LS1%��F�#^I�'��x&/]��$�Ǔ��@]�g�(+WBs�C&���3գ���ڞ3>:0||p.���țF�'���2�S;!�kq�w�ڿ�d��WZ�A栈غ��(����`���X��q)}�ώ͛5��"�WY�0�#��و�k������?�%��uu����fR�acf����t�Ċ��Q[f�G�|e#>W$�L�,�B�@�.y�ܝ�w�/4�-�n�e�Z�d��LX�$`�A�$0���0Y����٦���Z�Π���[W�b��uh*f���O�l!(��N��w�q����z���aw�a�	TB����;��F/J�bc��3@-���8��f-05[8���]J�?e�I���x��n!nWY�yi����7q�HO�Ӻ8w��!�7Vw��!��_��a�j[��R�ݴN<״���uO	�b/�jp�>������.?cn�xh�3�_���H�_q%Ct e3�T��.�Re]D�� e� �n����"Ұ/
�0����I�B��oV5��B��5$X-�\����~f���7���^*�V���^�N���i�+0�[��U�����3��8d�
�t�\�t��?o�m�<������y��m�q��DL]2��6ؼ��'���bҥ�ؕw�}� ���FbM��O��CFA	��5/Ib�r&��B�g�L���"Yu��̺��9�r\~�������_Ĉ����T��^t$�*!}5sf���}Bj5�7�~:H��S�[��\�B�@q�z���3s�T̔��m� �g����H�Y�Z'S�l�]�'�
5� ��;��mx�� �{�\@m�i�kŬj��#�J�`��b5�t{N����A�v�*��Y�%2����O��sM��N}ED�X�5ZX+�#���#h�%�*��!�������j#Lc��Q��F�DףW�UHu���1�<E���4�:�>�b�9?3j���lQܾ̟����$El�D��I��� ������� ������Y�m�iW�U 	Hf©��U6�r�j�-ͻ�2Xyp>#�-���'�ju�T
겦��TD&� n���K�qVɹ��ؔ�M`��z���J�|^BSǁ/*.©�r:�%gX#�Ͷ�����TŰ��	l�@�?�o\
	���������Ѡ�"��H��Cғ��i���$z'�jseՎ\d��ڂDw�[Aa��m)�2G�5b�N��m*�zV�wvw���