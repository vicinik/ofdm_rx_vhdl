architecture Rtl of CpRemoval is
begin

end architecture;