architecture Rtl of CoarseAlignment is
begin

end architecture;