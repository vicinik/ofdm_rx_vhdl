-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vwMSXp+C14Uqh7kM93gWzcYz1eismr8S8mr1p9KDyLfo4sJHS06WPXAl/j87RHV6RPnxHoRY6wpa
TbxFihrzoiR87hAJuZsdHL0SQOshpnL6A6pCuoF0kfn4OSFZYwZonuryeJkKb5oGR8CTJSsIFH6J
Qv+ZHegX0e8txES1RQUo+/6dovRXdEZnpHsn7IK4cZoIaLqFP8yzeFhR7aFsM54tbUxrb/HKyPiF
y9DZ9RUhPX73EpJUrtjhEyWdc7TauBYv3i8D1vkvfNi0pj7srR+m9u/qEHH25sba9OfhayRfibFp
rfkvBU9ga09Y1l2T8/8VgtPTBVNaP/2v9MDc9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 102384)
`protect data_block
B3uVghPfxmLtMpwmdCiJ0kkjGtkYgKmpgTiLCBkw6+TN3ndW6kR1H1NeW73l64Us5OamvqHJdkKv
u+MlMyOpDYePyCVpoRD4RIHuYsvg5/VqcQfTcXa1jshNhbyZIeKkz7Ne9xMvAcMudeZH12yFz0Xc
Sla6zc00azMoBHNEFW3BOWVyeN0x5WiL1p2eXUrrh0TWkTA1XkMXpFRH4l5CX1lD4WW3URQzjZhh
HUHBkNCTrYUo6hKE1+JHpwcefpj89SyzersxezKlX/as40KuR69qDaM3+i12A9RbYRSDINPiy+F3
x+PjmO1l1XRrmeZawk/Urw6miO2nHGDFwnuocyM2IbtnOUZW+jWvPI8tx9ips2akVYqoA7U2T4VQ
38nYm5PyGeqi9BUrKm71AtXvF56TVaOwLcyt7Y3JeGyoRbivFVeyMltWDqiTXE8mQZ8zAxWoHOHn
vVWRN54QY9WGTf+6dezv9emSOfi7jk8Lrobw2YdWI5fWlQGpxSxGUK43GZY5LdyqmUC38MYz0bal
n7f22WyTiGUpyQh1k0dFx+mDVTzegSyafBizRMlFLXcVeQDnx27i2wkFWoZjmea2shAYQXwkNMB5
l0AyyZM6Z47AsgKs8N7us5KM3291fvFWqjqkgwTdplRciflcL1Rrajs0of9NGyiSyrMR45mZTVnT
q0jHeZqf1xUHT1i4qjpLtZVt+edBRNGfihxTdkpnRS/6elDnkRPHoyDDsJCC9Mos/ZaW586C3wVL
ovh5W/6gEnBDVyQRYl1TeH6GupXOTOyfTyWnKPem9vra4lywwS3mLO6TtJooka3GRXHdWPp0szxz
wKxjQLmANPBjs0IPEM7mnP2Tjcgz9lfI8yk+ON+y+Qw/AyqS8bNd0RTzU/bjUlZ7lqCZ/fES2jhG
djGt9V/T/KrlY8KYLeUvzfD/V3MzeCbTU9zqNmn3x70BPHzqNo5kmUe5+QMjDkDP8Xhe8j0uVoqH
fT0D/eZtlp1IE28De6lAj+L5JWOlcU/BkKhb8FoUPML4Azj7zIU7oPnu6OV7uWkTit9m/WVryN0G
XIWXnfhtMiqXz8oL8T7ll8qs6vq0+n6UmsX3wgei7Cv0qaj/BJ6mHb85ZJ/rGk8P0i42HxfxjLOw
/6IEHi7Xvs/kuHHlGi7UDBlB8GjEKu6YxkzoN321hVJHNWy0DNidpKjsuP3MdVSKzbGstcUcAjoB
IYVWXuZN0OkT9DDE4Av7ZtF9sRztVHtdLA8eFMsOkuQ9NWmvw8WkpqpjalCl/n8QnYJ9iWqgOfmN
FEOXwV2Fd0ZVUIBuHxbF3YMkxof0KPe4FGHJQHkdBhv4gbCpBGsHNx/nXarkuvU5SFTjrxpBQ+q3
uV5QvCZkHpqY3dDBUi9/7dNJFjpk/dgMuIYu1J7DrdHpgaDJDz+IBIuZBmKltFZWjTfaNvLvmMUu
Rds3NA4i713gqLa9O4rAv33fLALNs97YkRBMLolf9/pGLyvvl3crS/ferCV11KC/q+Ci6MUoPRuh
cJUNUH62ViJY07jGc9bGvt7kQJxQtRGn6PAJ4fdYJ6fBK3k5s2Jv4qRQv5maxiElkx8ngVbuo157
T1b+k6RZmYV8hsMhPWFvvkHLg6s7thUhzzR392/AZkGmCsCU4Z2zQOAmyJ3Nh5/wVfzzm4NDFE9Y
fKecszWOGwntwma3PucbQ0a7YnnVC0b4vrXMz3I6KXlkbAcWDmR844tAif9bzjXPhH19g0tGKNQa
PnJb7jtkGK6wVQzN1GntABwQYsuGPsoU1l2Zl0fSuERKWBcluWPaUYRK7eRgwrw6Q2X28mVPVysp
kF9+rGnW7xQtVYXQZHLy8gHhglVx+j7VB+OpWM8oc5nxozYEuqEvrtz3j0pn2xtGwxAEArevoP2/
0hObLAXVcP3xWDLXXLTE78dOeIoRVR47FI9dcMvG4+pCdSQRWixXUObMrScbngq+3OYmxhHCddb2
ZR8NOWBhVysc0oMtAzzK4GmWVCDiyqVbQeDcnz6sshGkc/XOEAtZE0Vyjw2C/2CrT6jnAbCEollJ
v2CvAnSjRwqSfCM5ut+fLD5XbczzxsKZ1jmpeykocOkBDn96AX+qCB/AKn++RcEV63bHycOmxmVL
q6PMVR3vLuD49rOgPdOAKeNt4KS+xnPFhsr5VHeHlddoyZ/vIWZd+PZin3rUgoNYay6XQqjx+5HB
P2+8ort+07uPB4CkYa2fp2uRst7eHJfRq4Olb4ZCQKlVpZ1nAZRGPufWQ6yn8IASQhuTFRflO/J2
yNcRW02p6F+cAF6v+Ll9InUIfbN37D9yfka/IVbwfl1nBlHMmjob+9cvysJ31fsnAWhM5qH6ZT+t
vBKIWitKSckteahtJEAEIlA6WKZCfq+zhFJ296bWP2o43vA0UZcClvRQKxjuMQQ6MoUBFrqngZv9
Xe8kY4NZVjlB4N/BSK2OoPPRdM6KqW1KFcrrWXi99GjH9teF/wwMyj9MJpdbhzYJKHC5snAMJFYK
mZyyqn0j81HsW2fTu7b7vViYxHcBEThUd8BuACSqOY+/aw5xRp3UIsLWwJ0dMuf4m3ghgSlyHZMd
ScYMnPgQdyxVp6cmlVzlp8VdHM1AOgT3250mpKn5Z7N0o60RQHAiQwFOBW+JKYGFCeG/CUFAXJ3m
a6u93aTy+sun3ouP/oiFLjf6Etf/6uE47dmQiK4dOyMBcGq9W6O8P8P/QL17QlvyqRhafFb4sFPB
Doekf9nH4R7PPMLCAL7e/hNQBopvNIVB6NhJyFTYtsJtfXUlNYBtwkejoE057pK3zV719wBvLNfB
CZRcBjEjmm+pKX8RLAJXKUS15Yn63xqdDZiV3tv5BuxCLIPOVRwAxv2MdO+79bB0HtU9oSQBaymB
m7QkKuLdM++EIUI/AG9qiw0DF9GJsVJMlRSU3MBcCC+HWl73huEKDPwQsAtY3Qh+CitRHS3w4lCG
aXKSZIgHc2ZvLPB+vph7inR9avqCJ5AAevGWCcpOQ9gdGqnK0aa72yBsdDkcQvQmnlNbrqRYkzHP
Y+6doweWdpOO1X1txVuf70r/V/vn4hInapk4WI2wYQSpFblBWTpUx/DaRu/wc7ZLms5OhKXD0YwO
dQTfbuCil+n2q2O0EekaT/obyyInOW8AHr2Owc+VzARnkrykqW+qWBpG7JYqPAvAvVQTe0KBAqAr
acsran5eeItbPx4Bhecxh+iBpq9xWWFfxaRdP8mOPDzKqYQH1mDWuAJGJ/HgKnBTAuxLzAXJzc1I
2o39tP6ZhDILGMATecgYdYU8f0/xtm5mIbE7FN7fyHWYxuttj0pP8WtM/8sSJCF5t0PcOO9dzhDZ
SsulrnQKgILyMknRI2V1LF+CpE7J125Z0XONwl6TQF4ROcSUEF1QLsqn8CB41UuLze+q4ZlkGIoT
ZQrGkpHQtRcxzPIe0zg1J3WQyHhcy/ZcQXfD3h+6csGCdLJLLnnszBtlD4deXsQfdyVrF4cs3qHJ
3SGsyn8LTJirhFdl2spE/SOteM0i4K07wh/OFgBQL1LcaJLQvTA20CSVp3Z7F3cOctOPm0bUTVAR
mo+XGgAnbFp8iK9PAFclbtjIIyswLrOg9ilpHXmt8Ua+yL0D6k+4dt6hAh/tPLAbHm+TTYbqH9+g
5v4Jhct36RBV5dD/rDgJHXhChG5IZlBBSuXeUk4vp42lOJGbtWCMMvLtukRVM/l3KR3YGC1wG7sU
0ULd7KVidPVahfV9xx4ij8QRxmO4UtNPj+wtofJGrCP6gEwPj/ACXWI9ahmQ+UYkSkDLQrOFJczq
NK07A16E07Jod4m+/E7/xQjc0JweuU+zFGIigL85VIVTTXOfzCg0spJIz+dfBg1BvCNu1OEk5qfd
iEfM9y2Ep5wXhD+fR5UypPfTIPngcsbXx4xaLflAa8FFGeZQf5x06Zk17RmViFLpSBhx6qPN1S27
+ZtpCR1Fi4elSpYVMcID6qm/GSK5mZ+GZ2LJdZZPeIhH1v6uc+qBLXq0ef6jTkSkrAqK/VZj3H5+
lfM7/1cXGA8viTwTGrsYfTTUIhwqPFw4DSMSvZzhgJ9c15bVJcAczy3ZCrv//+JiSkXs1vCZOOcW
ZLJpz+kpb9OKiTuNwAqjbpCPQCcKPVFzx976PBZdiYl7IDTgo9U33Udju+ICBJtnAgZeEUyEs8rp
XCZQusF244r00PPpCE67UCg1OyzItdTgWUqyMTuJUUphHVmtlddnWx130cIwi34xJFO46HZ4F/64
wekbq6eLxDOdazIdpB8EtU16tQaWriDS5F6gz3bHErAswzdfVf0wpXG9frYb4SAowdhbuo4Xi2de
Lpr3Fs17DrX+EoNqQo0MCUJQguwZBmrKaMX9LrEhKY6teqIGJpww1dG5H6+hFcuNqnIOP4XhRuvb
frmmUg7K7WddeS2BNR4Yyd9mvlcVolcQfkzUnJSwcQD84GhQvYqBVcv8AEukliHSETqc3mrZgSWc
jIH4dHbKwpxMvI0jBX9rGY/TtzDnI3+j/JGxSMfVxMrB9KB5Mju/tBpa3Ly7hk6cMxjyEZRnReJV
qRqtAQLHWghPFDlCbDuDHacxFzpdTnP+Lc6/Jgh4OUiRZmVt3esVfFLqYCDpCKgx+FzBZ605dhEd
CO5Xn/Cy1dks43iu+8L1B0pGogcxxtMIJOBXNFe35hEuDfZvABRCTXd7AqjaUrhgzLqbw6UJbX7K
r42qvnPBi7gehNmuSE7wwbfu6YqrvE5g7anrk3yo31WwnH1PlQg36jpkr6dR3gPeG+0Xg+OQQrAV
HSu1lOwJ4b7rrVhzezVlUPvnMiMnHSN0i5cXZ7OXt/N6pPeSc0PDvankKCmXoAEBEJqHzQXhH393
tHm+/k0QaT2PWb8N1CD/PjY8SFOUQuObu9c5fF4h9tlv6rgafDNo3jOnlRpkklJph5F1IkOa3xpO
5xFw3Pw9bXOHiisn+0eQUozsvjwJncWnTDPSYFhLjvJw5MD4YNJbJp8oerThPCAqgNBcne07hbNv
7ih8bw7iRnPhDCILdQI4Cp0lU/agh697nXQBR9oVLSwFU2SjptyiVjMY/Zc7C//g2XoRhOgnJnVF
DACGqFcma6CXJjvBH6M2Mq7Gn2QLc9vJJCyHvEhNwtNfmVS/hMGMOIjuh+IE/PrAIk93IA4Vccqd
Fhuv7rSgaHqsAOb++LMGozZGGRdgeT0duhoTA+lGJu27Gi+d+tTBZPNhuf/cEbfTd5dWWFiAXnm6
IVBP9QasZBXjgYRFQyL8HP74fH+tvS/fq5tZT21gxFM1OcygGbh3WV/DoY582alsZDCFxS9dS32s
RfbhTlGgongjjZNq9sBVBsbcoNjOkznlsJ7DT60Lzf1H7zEyMZWtQxI5ODMLx6i1vIu07LdaMSoG
HRPSo7Eer9lXyTCntTbn5cenLt1yqPn6OAwD8I0mHzxdfpzXybl5auwXFarNMfEYXy1lYSfr/bej
wYEpQEo3e36fug3FGt+jN831aobtTO1N+iGnNP0IqHnzeTZs+MBumrEQyfUHQWdFrQJKiamyoZf3
FjOPqf5+HWzB+jXiGwhDo3xqqBf8XGphUOB48eizGQr11OMRKRvImI9TPIbVRAFb24/nbAK3gDYO
h5w7nXvt/O5isZYiLMlbaJWRZfqVGlrXjx4JXmMxXg2MDMvrzwBP7JQ2PAOEA6mmPo1usnV8NyUi
lml7+j2P5SFR9suOydJQlm+8qk/luSEghVICdWWvB1TuXqio24k0vIjumfjYc6YcBwCiV4FibOKI
JC2+mBvqFDsAbSU5hgG1VhQSolKJq3sHpohklzDfDOl6SrGIzdXJQYHLx86jyNh+gIFJl7Krr8Ev
yw+SW8I4j/Dot3V24kKLmBH3IZU6wpD9Tx+SkJ+h+Kz/pl3nGuJ7mdUWGglXYeGzVqPp0bY6Dsfc
iH/NZxqV6Q0C1kd7Es25b/Xpf9CuejqPAAmZApXf6pCLqnDioI5JQ4KrUwxhx6dxBLb5ik55HUMl
PiP5avmZVx1XI7kqDtskNOAZjEK4SitvHcgR3aEzFfyCa6pOxywI+UGsI111VT66M2E8sLqHH50d
RLuaF+ObwqyC0HOGiufiGuwUYWUM6X0A9Hlx/JXJZYgjH8padQ5HoqgvmFQmKVorLe2eyry99Uf/
pOMVMvFz3v3D+0gk/NiSy0MWfzV5zge+hBk7W355Z6wOz0eHTVCaCryLZIUsZOMxzjtwNh8ZKVTX
BVkWJ5TS6Fm1JKUY40gXBiOSQ3ECOEhWfnHlGOzJKtQlC/287QydjNr54CGWo4CyinpuFMwP3zAW
1fFt2e80/L6Zrf5C0TxWr7P8T5kEecb7Wf+1qcAUXIu/q7KcIs9c4As8s6GBnZC1gQQ5OzYfhROb
u8AvO38DKCzF//JlD5Na/urwowFGstQodtjvqGAqVt3TzgNTmnIl7/+OVxZt4Vv8oqt4ZKoW6Tq1
FjCxBpPYlU+VCrq/rCHfM1xtWnSBgFp/IQh+OjjZ7CanXAJn20MacB1k6qFqOACc7dOTwXwIGUZA
yQnqokO30wWqiuRedU01mL+uEOsAQxrnOwc2r5FT+dSEoU0UqKyrzVaIDYjv5YrapNuPeLJkMSvj
/55rJNNSrsfGfe7oT7PrcW6Sp/EhsHlv2kct1hac7Oqfsb8GlFxZWD0PqGSwAWw4ZOGgYK63peo5
KNCVbAZ+w+qflB0i2ZLzg1IQoS+CBFnzMVIlXi/GaPMr3pSKFHUOD/Vez0FS44V7O13O0dm+/m4z
a/jDwVU8Kfu8ThcDvrY+b7KuAJKNdQ49aHgIPnR0a2ETB/wg5vACB9u2r9/FzzsDLhbRUNC8nX6M
MDq2xALKaX4MhMv//ufVmDV4ccsw0pDK92OeBh22myJKkGPC/9TCXJAf9WVEn1ll6HSRYaGAJo5B
Rx7m/sFQownGDe30u7PlThLDtv/uwoMYslViSqlOhtMBsosXJEin6Se8JJkiR23qlu8CvWonpXRz
3jkGIs0rkALrnhwiAAmlmIlrX5elTxWOJ/ps0z7YvMdpMFr5DeIU/zhbut94F5Kbtf00cuzsTTYH
4xQY5zOEs4EKIKqYDt964jNKBRYLkPh4l7BNRJkhS0rILEyqdrIRPmt0j1T2zxB6PfMBO2uGEvG/
e/xuLy/f08ry9x39449lJ7BZjV00pK6liiIuhKap2ChWYrF84bWLLZ9j0bfG+5QBc7KccSaFRv2n
vtHaU+S2SugjWuidxRwH+dDQ8MA8ujvGRxjZj1RLn6aOUZCoW2MjYZCGFjNQ178OHi9hvON2Qvyo
KDW4aFnIuRKES7Fcvh6hOJHxmQScArptFjCDliWXMp2dKbPPNQnscnd1/6zNdfRF+bUbZEzJJz2T
Yq+56sUzFbwJuKfZ7rEezUcctBdYouz8AGXkapwEd53Z/EY9Ri68CRroPGeSTuiR8k/YpnEsLM1r
QISCYYnInGkpnbEHvIBeSAlBaPYnD8IxajWR/l9ALB7sy7TwxmQCM0WLen4Az18R9e/lOuETGgU3
8f1m+tp116QDEFtEQ88b3wjBGbgbFCgLLVajm0qbUCg6mKuU9BVQSAn8BfUmsCaBFJLKQ82n6NZ9
V7gqmhtcLJ2+k8XmA0k92X/x2A6Wdb7QNLX7aAPmLQ7FFNbpU5rLn0qaKzSuuYRTDmbQkZt32kwi
LX2Qg7CT044Uy2LFHxoLaNd9KvtbOCYvO0IBAYamv1wbrniE6ztJzrEnkPagFh5B062NkjMJga1t
5k8YKp64WlqmStSBy3JxRZovb+7RDRkyu2slq9rxgd3eFfyQlHbYeuu4TDO1DQG8iAHNZk3gCFga
vHE8ftz35nV8O0dmtcmLGD6PNOql3mXH7nkBXJaC7a7MjbYuHqBxR/WYT+X/qWL+OSfzIl6MBYVr
gEdBVs14DaDXc5yC6K7jYqXtYdzm0Pdr62Vc5qQ8ZD+BuErAUiVsePO6fKNySFakLhLPfq0zNfWS
NYXDAOvkZyLyposfk3btfRnyYJ2sJI6njLRPEjYlALxYnZi7+nHGUXQ/ZJRLki/arRLYttGd6H9b
tFRUnPTypkDz1Rs80Si4fwo0AkYmXeoIOVNMzPRxuMmCEee6z+vUp90ONjcNTINABaDZOomKzLVz
HTWT5ZNyEiJa28VR+NAQrVU+ciPFsm9oKox/fIQD6TLMVpkzRnGDjqVcPvYZFtPCMKK7z7/lMr08
VbAvGLgpEpbOvXO/avNjRbbfX+UsqlWlEWVBqrJBPS7HrLduzcEqoPOwZQMKHe0LztJ62+dgpMTZ
oBRRCFnj1mRk4/RvL2IcCaY9XXCKTfMbvyu8FlTaM5tz+kfsIxSu9C9uMvIYLde2m3xwcfYxVEf5
TIyoEsetfcsycjkD7+IJ5hXjFkg6Xrn2jkTtgFzLcl5AXH8wTlJVWHknHAlFpsx6AFWofqdMBxUv
Ib8yG8zNa1P0Tg+eEo7wvv1GtXGFaXLBdSkpu3ZEXOVui4HrTbNhrbEiWewnEsQmW56bFATeJVVL
QJP3b/bORFtjtqyvH35dpVxkQhGIbWhdp34FpGk09VdTUpnEE7zVO9B7rPTOEOmhQj4anLmKf1Az
e6gymm2ZItWZrCzRNQKyQpWdydudltFptQ/1IwluHD5YnsfLjASdovuadbyHVeF7q7gF3HxnxSEE
DOswP6CgWG/9rhlsAV4QWYuq0j9P4csNf6DV9VpumlxX7cOA5Ile/Fiq0yMWiCmKoFgG2S4BP58R
DcRFBIGyfOyZpST3p3bOEZCFfu5uVopupvDGp6+AmD6iYBcfzelnJieUgCIiFlBeUKCKU5cjHX10
QFqPw4i5eXAtLZCKO6DZ5eZIpWS+uhi0Hj7p12SNfqcg/tIYfW79fFYzLxOqkDuiCSNOJUkcIcFm
sY4UPl9bxQuMf/x/BEfCw3S/pOVJ3T77v5A+yanCi+rlLLf7/pqatGs0wHyZInLykKzKk0PsDwQW
ENfnjfwCQXmC/vEFP2qxKFira9wf6OZ9MydZBc7YS97x0bfUepOmJ+q3Q2fX8xSGqaBMjIs/Z2GX
pkQjRcvWGve6VEpr8+foa7YkXhQJORTnm3f3EaswajYYvCpaLehOuvzDRdP+3Bfb4W0kspKfsveU
+wgHjKD6a060YC9G3b/lMZFFgNW0OsgrhDzt58TiZthG32TktiswgEJarqD2bCCQYUoLaMnT6WCE
RpyeOHWhzXLXesi1P4Nr6Yd5R4xGKhMnd6bCTIyCX/HOUjmkbFAriKl6xYl9RSeGnXT8QA7gEvB7
zFRTik+Fb64uMaBtrf7s5uXYsWuMHeQKqVMmxzhNhI6sfrldNIXabBhmXuBeeiykWSilcJJ1NauD
t+8yZrOy0lc0ATUUy7y01C13enuADs8i1571Z3VvWkZ1yGycGu99fpi5PVIXgInD0ovrCvq85TjM
PHDgZRyIKqvC1K+KtfDqyZUFMwh4SXYbrFiUvxwLfNq/fn/xbDBNFEITimGqR5X7r5whOZTPjhuF
GBFSvEqzkMnF15pxzwSZ5nCVp2fwbrJll62PhwpO5pjWR5MuAoyXot5xpXKfmSEfYYVLNaEs3Yik
hZfaLx7rqeuE3Aca7hW65aHml1DtWMtDPBCtOwxiDkr6qTgCx2kM1Q7IX75myXo06va924WcFqkT
04oFk456XphbAgG4PSvnwCDWj0kedZv/5L2bbgTLwsusapdhiAct8DeoFSF6pe60fUM6AdpeJErP
ORMq+d6u79CF1P5z86BU04Z0Frzvawb9r7Ln264W0mQl4OwPVT3a/ssClLHFnxmzJqs1ottQ5J+O
MGfGL2I6J4BB1KKk1Isn/3aqtq0fZoTRWh4CpQaLXPsdOkcfPMUJcd9+VrxQYBcRrmom3lm5Cecx
Frp8MleuyNY+FH+5yoXxk+wxbtlvqB35kO2IrEUmt52nmosw7dDEfTQGLSQF/LXgHE6yKZIVNfbT
6hdpSYLMHLa8sJ4QtyMqShvL+1sbzawuSrEm+BE7VbEVqso5XQ59hqBzpfB/y+AFrrr5TzgtNv0X
37QMMnmQDZp8mmit4FIp4wW9Kg9XWi2vDgCr42Xl55PYnxZH9Za6x+5ni5nRBtl9tMZHB16raQbn
W9TdU4t/HlDTtx6WEjCGUbATeXBkV8U65HNnX6xQFuHlJEoP44hr8wj338SiBXbrvZA3syMpx8Jq
X5Of0QFXpQMpGeodGrpUcvrwBcJJHZrD+JSBnPRXaGs4g7KgLOtNqnaMLfk9x4oe3ZhLy9RMvUWq
rjR4lVJlG9x/aP9VCT29tBAza6pbtfICsuyZ/XW5rjnH8yMM3BlPX4nRVWKzS0efVjNtcu6Swh3w
E3ynbWRwvaOqZtzmprTOBt8vLaegcaq2jIi04M3pRTQ8TIe2LXMtNaa/5z5tZuJIDmfvW/jryTz0
okrYru4vRgAunYKcnCAhyyvD8mHpIWJGVBsciyHliEA7XAH2gVS9YgPRmoywcFGIHq8O3HXfxtlj
FIMbb7Blzcr9cM4SrSwNrmE+faRtNgNtXa5oagXvDfCFHWizGwYuQ6p7aUR0gdldTM1EL/AstEPz
UMdSm5bq5M6dQdI15t5RfRab14wkM6B0aVBgi+sKyJwZxsLAkMyXxohboVNTzgyCoG4DDKoo4iaS
SNSaILeTikQ2vbc5Ip+MdtEeQZ8Z0dZpxmCLHmSYdh9KOuQ4fRGTHQuE+uyC0nMeriKRZEB8Jsuu
cCV6MAyqUzdHPwM7ASu9g2VOuDAfadXdHcUIEHzqLC5Q8NpH+HKC6QOPrNbTvHCHriyXh5Lco1EA
SELMpg91LEQCk6vl4CEqa1xdWpRadoX4TSCLc9QbojPgF+2cBKIa6TzLrS6A7PvUGgRZAgr34TRY
XFzml4HCI/qC1rTvsY7csSHtbSSfa/49+YKl0xN2AzJH3u4A8sgQ9387GJvZ5OS3gX0HYK69dUF5
eThy9p3M/d/v3R7J3YlX7zRLMUZMhzZyFKi1aFLpzMe3ZYncVwA3cMrt40vglU/9Qa46/SBMpaeu
UbqFePedXtd7ffW8e5DeFWfIBsN/AM55DdgtF1XZ5zW2e2EAE49qc1v8pMP2lwArQdbWC7ac0VwS
eS2On5jAVyGSWknFk53YnUt8dxKLBTAf8euGtW4VE3UcgNzgv36UbrXa8a4QTHWDlRPCgFrSTuTG
t/p5omyIKDxTemOoz/hgIuaSXGxk/ljjlqdFk/C6JGT8F9L90mn/dM8wn4YOD7VmOe7Ffky4dMl8
uUjW4zW3xJ9HVBbkpv4pqcB+Oc8QCzkWs7h11V7vdPG7BQPVl27SMt0ujgtccGABDMweJrfFSADo
iQGFLwzDsPFK9wXhVCI+EhO5J9vGn9d+nQhWr95sD57MT8eQ5bAK+Xn+aBh6A0qhsexiHT/qETlW
iWPAdwHF9oJrrkfSER+S8mc8nY7voRo+py14j4ZzBFi/0Zzq+fgM90/ZnMZWEzgjEMxDJ2F2Eomd
FSymc9f9iQlSGz3YzAvUAjX25MG4bfwirWS8caIEJ6PZ9+dqy9dOxa3m+np89HR3w4atWX1O3jMz
4Oaibk7uzlfkNHKcw8QwlV1dXQo2E9XZsdIIP0bs+qJXiFC2ojXpf3zCTkrqeSbahvysvQ8iQ7v5
tNRFkVKRabnmEsut3FtvOO5FOFgA2AQi1I+K+0bdJGRbzset4id6OcWLk6GFiD2v95hJLUwmDGAO
biS4l/+tJWtbFV1USRHoNpuyY7G9iBycD+x7FKfMikpu9Un116plZ8C+tX3VWZlIx7+qSLHRiIab
LTaCqAFiilNY0EWQyn3FvkavfmZE+XBcpA7cCh2GzES4AqhVN4fg0Cy2vG95FdCjwzW4MJfj4ymN
F6Efp5Sb1X/3gudnTRqiTVAogK8YW+pVCElyXI7KA/Wx70A3Rw78VIsYP1CYen20ldrtm4JH+DJJ
ctraSse4AdECxNHjiGEyKLreX8c25gaDJ/J2+r1ZpZvvLVcr+NQImTsgetjVgp/PPcWdpE5Sja+D
kzY3WHw1yoebZ3X/rTITpMeCRIMtMJiq12+9ks+jUd1SexVr3MsZpbFDfLfzlfHsGo3MseLq9Ude
UReyrbvlRzRaH3DrwV87MBeR5bZY7Y1aTk2QXAd5uyG0/d0l8BcCJ4+B/TYQEGF+w3Cs6iJescin
KFQF6n3d2MLr1LX7rNQMq07GNvaMGggEFFHZlzxpc6bvkK2hgH39+XdisbMXVgCQjtt5YS7vp7Mg
vpBsvlOV3Mz3sxbRx02MCBUJuF9J+ymjZ3xDXqMQR+mf0yZATuXvet5a/c/uOuQKEX3Z3CRh2A/2
V4ncWEKl6LHmnyV33tp244i7Lgxz2/uYjH4fQRxSLO4Z5kaGjyAS5OvwGmVUAk0SobrFigTLmUrY
0oGrRzzHiC/6V/oa0TnPL8vPTdYoZVn7ppO0I83FsumbWbXF/jshbT44CDeKxoqIAoAMTWW2Nb3m
7FXthya5GIwkt85IGdOG6XMerPMaSosdrdYUBPR7DSrXnkXGGDeH3m2VmtKOJJDTdxJ6nhwGYmDk
m48EVYP75luiLcaGF8KDPwuwklRw0u2IcWZsCFXNiA6dEXY5VGQw/2ob8N3JBikLKXXJFMDLhqb8
hBheE5ZQZVSYCi20/cnbf8IqXSqDYnkie6I2kcWpwk+WarJeU3ZcoUSeDnE+cVOtlznK9U/UdmR3
Rj5kMlSTF1QkI7CRN6OEdoYOYvPi6l/ORxeQk/S/WXqmak1WfZcLLCkRBb0ujRbf7gnSmL+AyDQt
1gSpIXd+gzzQuSVVoGVHIbLBrJrSrTjzI4yKZwurXFLTkcr5iYuLvGKwLAxJ9EjS4Cg62FR0yn9z
jJlW4dIhbRAvmbYOuLhE7Y8cKSrROeUTMPqu5GTSv5N/Bbem1uSL/IMybSabgrcInmLF/dpw1IYI
Aqc11n9x9uwIc7ifE3kSXy0ZC77dL4hxl7GuKABogsOyo6AKyVZzOd/L05DIcUFNukJvTEqXfnAd
lPIWvJKj2E6OUBUyQAWsD9L5Q4kzLmSlP1a9N1op6Zu0xJzw1WclXjl7pgcKsPZdfpGHkdYfZGMI
bfOP/cZ4hjVr0sPvqF9etojAO7Okks3aRkd9bL7hoPzBhDaTpGoOsZx/sm55jsJGIWYQLUvrSukA
u5cCzX8s7Jvyg+xyQMDCvsS6f7aI5l08ft8+wt7ui5t7Y/YaoG/OWYOGOK0mG7Lc/ZqMAhu1/+Zd
D0qISFKIxz45+2ISKmqwSaloeSvDT8eFClZbijrXbEIL2mnMAxxlNBFOO4loIqlZm/0JzjE4SvT8
VRkIDciq8JmhMlssqN+TLx8YolJAPn7GlxgZd0TTyWOF/fMLQdPG4tqIG+5tM+EwP8+rf2st2Jdv
wjctmMghBCzokLEkz8H+HyVBbc6MHIhrLK+1s4YSjXGiTUOVDUm8bOGhvmp1OxFNNFz7PGRRPE+x
qz2wuo+QYLzMAadRUHW+ans0Bli+kwdrzVIQMHfj+UjjuePS8FZXfhNHduvsrSW9flq20stjoNwd
1DImjzn5kRcJdbc82H0Ms0qt6/VdyZjY31UBrxfFxFlRQWCP4u14qCIaEi/yh5tGhw6BCgt9p6Xu
vWPqqpOQL7XCTu76eqscxIW94SgT8ZiR/HEfobBJsywSf7QyvL0phnQUhB8iaEh2/cYXWG3Oo/Jv
gP7RPGSncqUtYNbzbnB4kv8lwKOGJpFnJ0DQ9PsRlTlaQgJgETxdnPze7brJ4pysefx29Gb0xypT
H8Mw76bCfjYfgogHiJ1noBXicv5+1fw6yUZ/1B48ENHInEDQKz9NqDTfCI8teF72XeSOQ19yE8xj
6RJlZJdBZAqKX6EHjre2T3DOKctSWZ7QoptEOa09+FQ00B8ZqA4nG8iZMvDbUbXOvmplOVAtgV7R
1WmDjqKc1tZcUemcQJrPy16uKSbxaZgK0brBwYpzmHLsCuEjAI9UvBah1xZl1owkaijb5sMYdrBz
G6oSbOk9lOdaxzErxX6w5nsqGT1DNtitMWtP3NE1XOJm7Ryu7HcgNBdO2xs1PQi/9+33bPMCtM6+
9/7a5AWUSPQHcEOt7HRd7+MNPkWs+rbHPK+6Vs0OKNj7cVsn27v7+zhE43RW71XMKDCq89cbaL4t
/bZn7NF3IBW2TxNaJZyar5ycrlOVJDLPY88lfnCnh65HMt3/N/uKz4h8QbhdTLVodN4UUKVigYdI
uVu7D0GiIOyiczP9FrUcX9gMyidT3hs/ZCKE0X+rudnvLUQ3iLG630tvXfJDOXUWSuMJoMYgo7jV
ws/2gxL5t6grU21IKMRzYVWb7q+EM0/zFXlbLyFirlRHey6mMDukWu72/+nyqj6kFZOg4Aunilwb
IcLgTu15JC6fnpkKHuJk+N5Zt7wzE3WLZh3YxSgqcu2KrK71xfj4KqVAjoPB/90x6jYJS4SZob1Q
ZjP8ExJ0cG3XepEqspIb8EArUA0gbJEU3U8aKvVhFujNVWuoiH1mlFRqoByjyvNOFFDEPNmp8qTW
btbem6bdgsozgRwYx/KAJ0LmM9/BXUEsMmR8/zuqTSJztlfIRKI6HT/6p64SHQrjAf6q2sdwId5d
HdzjdIwa9oor9IwboQbd5fCQ5aI8+8OmdfgMqRo/wMuQcZ2Jut0wNaYDm2k8uWk71S547/dPJNR9
uJIIu0YTT5P8aGZYNAY60quOWL9eOGjGtjgj3tth4nu1JeEs+WNKwT+6pB8xDzowvUdPaq8TqjWC
UdL3BlSAhGJy5zP+F51nEyx36uaOT1Wd/FEsEHOB7hn/12jDM3svfd2j/ZzcaCfE9F8odrIbvONi
wU4XVco2ZXktZVQBVwIvRDW88Sp8n8MoprBzNx1HwO4Oy5e94tPXxAAvBKTDjQeC3qf6ftBw+uT1
GyQBtNsj0YVadRsDU31BCHmM3yxbvLXeSajkOsHxuZNlW7vTfmnW21A5Cuqmmsbqr1gA1ALiC61S
YROtzKKrW5sVcz3jZOueReuzTri9nW4INQhkXHJEJ8Mgzwzff71gi+aJOw9i75ZXgCAm5ktqE1RF
ADw+5/7U4EOQt+mNlYOH6UGyNTa4dl7L+iRClVisY/dLpjbP8LrarbfAqLBzsXuFKyJ7WdrxwDoU
HH04beHib+ZJg6ud+mar61UsFM4pA+b+G6CsGAnTwXgEcMVB4WzqPshCoerd6qVncOfrj4m9nsV2
/t7wbw+Q54LV3xpNUMHTO4xszgMXAXLKpf9kAwpF34aKeyKjoNuP544vwXqIkMY+txNKA0IYlhOr
4gc98+BLOFES08kL/cetjyv7eSLwwhiYz7p9qb8FKpa3kzctPWiDyHydoIJgCw87GTLk6RwRH1nd
7IXSFzS1hAJrwH4fqJotzOGXryok0612or2PKDzapgkLIi4gEjY8d7ysaJvhn/vriJC+c12c/GQM
Dy+73IHAAPXeKVHPOPpha+fg0sZogr3fpWjvWrWatTtWqLRAEtLEwsO+AU3ptHy0RlSKseQqYClW
USTQBwYAZk9089HlOq9ZgAdbODiK74Q/Yon6KGgJcychVqzwzd6Oxqj1A743XRPFhogXutX+lQth
yTlORkD+b54e+EfURKVPpI4l1II9kXez0iBhyYgYlZ+0ROZe7z39dypb4LW/pQfSJLvwiFJMy4s7
BLazJ3mEy4+g62zW6j9uiX1PCmOkiaWLioTqfBUzh65cmqT7e19Vil8Ur20+pn2FKuOf7KXb51/n
SkNRonbV3xGPH+IPCeS2TUG6Y7/dQ8gUWNAUOKJHxqD5HdNLUggcOvoeGBOsVkpKNuBWcXnzDhKC
OYhYwGWfCeFFqhdC4MoWqFmeZlVnhIs9auInJ5cepDTdjlZ3u9Fpu9OgkD7rm5nF4XC60baDnwQw
nIUy3ifPszJ/vZYQ5eqGyGdnxIdvH+XmDwqJ9AHi4M2rhPDXXfD0kyJJYd/3U5iArEcl7BQFMBTf
eh4bdnZVII+okypOvyLBheqNX06AIfgL1LnGA0RGYw4knfeiChOqpSOoYfAx40D0th8H1Lt2odzc
tYI1DSUPqF21v0it5MP1NXp9Vf1VBmxpDcja9RSvOUe/rQ4pzqXWaOU/iAGdNlr3nYX140KQnZFm
3ttNd/yF8GAVAFcFv2c/vDVVaNLlVGZa1Dkia57wiy+zGCKua45LtiPNeW1UxcXZ4sc8bJypSN30
NJODP9CxsDRTOR8MGh2T1yTcsVS8dl0baJU1fYw/qYOpoxTFb4rDK6MvfHQowMP3Zu5aO4oJr7LW
h0eQiRup+BnsL3Wc16OGhpouX6/2ySLdwGcPMdm7AfgTlpXmmk3gqkh1NcVpW3XaKeTYe2STYvV7
198qtgQdI9qRBftoAyTLSmAjyToYU8NDJQldJK2lCzaaAepGCzfxAcbe8XAH/DM2ocs5Lh9yLwVT
LgxyvNy6fy4N/SQuwPqZOK/K+QNSz+ZvUuRwk5MBs9iupYvFR3R/FxYgfHsJNd2U+JVFMPuqf9aL
4uYxwcR0f9mti1opJ+/NXkaYUovBOHfJMXEknUU8cjagzcfoTSD6ybuxprvsBLXe9DGTmFwYCraY
BRMmziYLfV50bHJOLCmTeJUsBHSh9W44SId1f9ddhmd3grcq4HZbKqpZwa7DR9VEoYQqIYROwfak
nbaXJNEiZLud+6uws/gkdNZYf+ZCwp9YtugsTzw/DoXIVozFLLgY+nIaeqpPSsSnj2G1pcPwa/0X
CVEHhoKHFqUMjyF48tnE0uQipCStQiGJN53BdNcW/A7jUFZnbaXLLLn/XB0TTbJpEsTVF8E/rtKd
hfvPxI7y8IMW5z6HZR7CEPPu7UH0RHUlaDcQus21lVIKfRSyMkZLGdbyeCrDoU/K2Rt28MdRAiJD
IgOBAaxaQXRQcrBSlStZyWcSyK+i/oxoZqfaLbBh905eB18fZ3fAQDgySkNWd5jP9y7pwsudwt0p
Kt9kKOs/NeSEShk1zlTETPHrKDcXYK7g11TXahiEpSt2ebOxPIsAPV2cphBJa1PZmKbcnP9DLjPG
daNE9TO052xupDcgbq62pG74jx1tksmvvTaxqRRm5Dls9a4qQ5omnB6X3albCpHbn/KGJGCHKu04
kfSLksfFKfis66GI3lMrptNZrhXqd9L83hUALczaPCh4z4gr4ZLsKFOlWaz2URxs4eC27znPqq/b
dZziMaPPbMORp1eoz0ZYICNxM54dwZI8y8ialoNZg+6Wb2d5FCwT4iIADQ8d52ZtNL6swSvIjTSq
ly/jHidt4uWnU/KpGxsV1ecCWdvrBz9N1EQF6Eiom+a77ERJePhmxMeSjpHTA0LSiUUTIfw3TtSc
oYSkHHkvs/u8hcC2EnegU5w6zF1ntnaiMn6NTmIrcFJAyb7z7iWZNVX4odeia3SIrdYprubmhNHd
xLpMs9w10aMFubmYtnzxsC7lBki9GcO08oYb8S74vq+8UtlL/5YBs6uEoXog5xXaXFokXHq9cPIl
dx+EDddY4RFrGTWrYoolh5hPFUVjY2B2WHrk919sfmjWvP/1yx+WA1BoTT7oVVenNvJEBb30niUl
te/o8YPZkYrKYWH/7iaaMZtoFcAeVZ2xkV+MPEeY5QyoKiLenzKRe/SQJTk/eRbiV0ia9JJIcf0L
t/8J0fkhj939TY1fRYoRNPWdro6nna8R2Q7d2T/O5FMxHl1M7y4d1z+G0pfAjxsxHLvH82U3Skuo
GR2VHxPOnfV0OK5/zlk6fuSchiYNCMCNKYp4uWCNYvsTxkrs0GLdlMhomI2r2engkjUxleWHQuCX
mKMjbfXyoe7aN9b662GTqZKXKS0adS+HHCq/HPJvHuyvYdPD08qxxFyOm7ufV7F0x1zqtFJLl0se
vfXqBAyhXM8sofbLhRTOBFtH9ZSnrbD6spDYdo6sPMotieWC0LI893axE1FVif6AV/cYAxEsBo8P
NwGAebBxl4nb8/dYt2hSdzpGZ8S+MG+XaqgZkk896oiRhV8ocVz0RoUovxEOhfWuNeRvb90UawcF
g9hbwGB9fs/OkOyN3ahoEIjrZ/0KQycUPTPZEXtiI3JlM/0BOF394W+rr831idFNL3k/ZaEExu6G
v4lGL4NO1TpEposlRyDA5d7dNjX6ZJPPzP1xyll1Fo99FqlBTEOpML7ggUuy3xEAAOAviLwAEOxd
c6HoVUOOz9erEdsA/OWYGbHwem2bSOfqS3uYiwviqzYW81dojFEM+OLjRHOTSfcN1D1jhUNBrswn
RIPwZDsPkOYm8u9931sYql3v+qZ0TLexlYkkpJr6JciS4MqYFzSSCcSwhPd/VTBdoBwOs+7VHMYb
jWodg8dGIKA9zB1ImzqLlBR9+wVPgpnwDj+UEffqMXZCi3bP2NSfpZ1LpTOagbj57pZebLtF+FJM
xbfsGY1sw3rtf2pKkjE0GrLNayy8BbeD6xctHdJsfekNLSeCDRKQM9JP5To+ngVuGa+Wbh8DcVwX
miqI5qdXbv//ifBD0DcCZnMueJXUKEaM4B5qHR1wzp2kjVqNzc675rRqSBoiw8R2BF+8eUdkDCUM
PXaxahzoZ9uQ5V5Qf5NeP6kpZUs+T6pwTv8A941phT/ouDLet/V2RUdz/RsCYnG4k6FzyPvpHlb0
8mIePj3UCS8FgVU4UEApsMKXQjiIRke9pfvo3n4iN3KyhOFK5HyxxFY1hAeKX6mhBfCLO16CzjQN
PiHNfaaKZtF8BbA4UxXzPs8KyZT1K4bv1M4ixh2i6nLTCDY0L1jX1Q6U4ox6tPY5YixmcwcFt020
b4Bim9YLN+9UWJRHo+50LOZCK7DAUGnMRaE/sqUDLQmU3+VWuXP6Kyo0i6Cpx/VX50rhUHYiwPty
UN8Lj2eUlFEV4wAFNU6YDCTeX0Msk7N0qIYY93arB3EF8lKMqcg/4rIHqhU3fA3sBis2smWaNEpn
CwgMslj6qnsCddt4cIBY86AdlWtSD5QBX9SKzQnxRESKxlCI1J0xopR3pvxK7ffa75Ishr29thik
XN+v5lKQe7o51UJEsjLQiE5ufRlsQsWkZZr9nWIToXKMY4MMgrcI0m2MZq0m+XhQAPmYLmR5WvHp
AxQyyjj/gqVbNeSejST/4DjZSQpgCkijwkatnODAmgbYtNZeoOXjsqxGw2m4rsDAbkLXKnIdplTg
CpznzUOZ4IddOv/unaWml2sXTHspBoAsqltUKR0oHxadx3R6BrnTBmo2ocUTWRS1WrqWjrk/53Xa
XXp5NPwCxErMj/yZRmzUVvSmlm75OSJ7z3F6NkMiG9HHuzc0x8jFadpWYjh4PhFm278qGZ1T9/iV
FWnQqMv5Mbcr7NKkxcy8x9gIUFuvBJ1KhXOh5cUzpr6mIO5S/EOWupHAgX3I6N9iyb3WBCoaMrBk
iWDvqXcdV1jV3pty56IKO5wMU4czh+TGomSU/qC7OmyLaAZEn2pJ5Ff67BWQdvvpSL6lfivBwWh3
8ata9Uw/gqt+ydc2PAmL+aGTSjXrrIkmWwTLYd8DvKkTCoQlxG7IZFhighaRdosuV4pU6N+NfI11
EeziWgdTudlF8l1MhSiKYUgi6agfz3QCCwfk+Dr6Lb/rcLC371tKHgfPFMhOq3J/d3/almw+BHlC
SodrjQ7oo0YPEEfGLb1sNt6HtKLve/ejo4uKiETCUW67J6ztme2DGVnX4PhURT7K07cnCUhZq2nf
rZFX2sCKeXPhY9niEFLb2McXHb98o9y4+iWkyNank7afX4/QIVXRKjeIyOGnfUZ6dNhB5ymd827o
FpqOL0rL2BEfQe0V+tJJYEg+08nZxAVU8Ls5oLALqR91A5iPpRdxZ7Zp48ZO0U4krLMVQ0v6X+U9
XqIzjKxAebie7UO0n7S3UllaNa3t/tNwXf1pgzXGe9Yv22DU9QxFAkxl/DZRJN5EvOE32Df4aPb5
ptgObPc+Fc3OwaXozgyZhsj0//NE0w/RFQnnKWl2AeIkBslDwkDybSdFbJhpgAhfkhLPL1nCpvxy
DHdiGgn1PeG6wyxiIzbXDoWvTVVccyHpBt7O/wEMxUP2JsO30xGyNmPTNGwfNpEdBkO/FmCfkHMo
8X9iWV+Vaqdi/20EU04tQwaNUO3bQ0a1Yf93AT+xDEUr3Ls1/3OiEpQ/CqWZz2F+DVFWYfbOI6cE
63iEwByeeseRyhF86IMyQg9ip3W2oS6Ub3BJDqZbIxdoX9yC6J8Uj7LDpkiXTc2hfFFu2hJC9+JC
a3GHLtzyMekCQp3o22zQKaPOEJifha3G2MzOPRQqgCnmf9idwYa/reZgbRFOkifv5S9n8SrxLSKl
w1kdosA0UdCid4JLTtoY4zqTAdczY4cn8h1LRd2t1+7jp0md0VjZZdfrZwnAKFPAT2YvdkcZNaUG
rPD2IDp9/YxNiId5cnJE+pd99sl9iTuhYkbEKrEH6JiCVxBvK8Qd1PxXbvcSdE7R8uzriZRGIbzP
wQJkWqVXQdaNham5z43LD2UdqoeonRKwbWfG22Ua1JAe4FFbCKXfb/ymLDh+ZVbwBXNFJ+BPYiGw
boTUSJu2LElRtq15husi+8g77vXAbB4odJW5IJKQLYzYU7Kb3eOFMWwYLBA0VWDqJsopfz1iW101
0mzUhtb57GV7apgN5ox3790a9/1K+tsQVJov83Wpi3ws6tH/WLp4RLfPNv5eOfAyZeL/PXfLlfmK
VCBildmPMn8ZJjW6/8CLNCoUwBnTjW/PKu+zAKNY8gUlJ0PazmeL4rQG7QP2hpWOohpmooXYgTrs
D9GuKi0tEonda2EI06MiynU7w1BiOkgjImjfk2jJYVMguHXoxJDAdQ0K5fagpPPg117wggtvgsMV
+ZkqiDhlDmPT1CeI3e+U04MfE20Pbdv40s8ioWSw6b2pheBLajdgocyhDIWweS8HA82UpzM6aC67
nQgl0gigs15+UvgskQWm14Q00DZyEzju7bP5NCnWH+I5ZdHFlZk83MGAnD/3uTVjRctB8kIjT3LK
Ylc3YcLdo1sWcgPCDHPpN8rLBY1lPO5623bfhNkk1hsOCSlUfEeiTTxm+N5Xnn8Vc1OV8EHNPhvI
WTV0naIBAzLcogo1Aj7gQma/Bup3+rMOsRK6m1+/GMh4iVcZiwecq72FQ/mKhrXp60Wz4ZDAagyc
2o7/KwIyJj7uGq9KBN4pO+axSG66tEn9QZO70x+Nc8GE0etQjGXpbYKm74TKTgQ8ZnzMYSGoo8li
Fnk8KbBhgYdW5g4IhcOh0dmkyYW5Se7xkmghb7dOvWZJzG3CrfhdhrJSue7FYygKymmdksNL9WXg
KOyTb+CtN4xF6xsRW7j5gj0luTBVh86VimjD/muokR/9f57J/2K7ynxoRxvS7thU8Ax6EN3Laq37
UlAwh4u13aOZD73dxAwWH+dIfkfXuL+HDSvBl+dKpD54PkJ0r1uDWevkoXjgZazWH3Fxk6vIbcbK
PsuGrdlxbmJsApeNrtf+Su98WY0PkE8vPCC/ecHcHIaU73tVWHlVOiLBSXwdbEHn0BBzJkFpU0+g
ugXBIixNC0suIS0F70VKnLryo1litT77y1Dgvnd02b0WfoixeyV5fFj7jzfMDWfLhuMaFvgTg+PN
zJDQiZm7300zfPd7bXIr7o19WRX8XhOGq2AuaKndzzz+QoLVNQJc0VO7E48b+Spj7jgdamcyDyGE
P49w5YystKTVy4/okzVHsScflApLK9bTWi1ewkY/9A8uUQEAJ+6I5CTSQoLGgCwEo+XLt+Et3LF4
iarTZNC/igRd6XB1Q1X5s6AdDaeIpbyJB18JKmC7tI1vVh+iAT96/H332dkJfNAE9MJOYVXPMfju
b0sSxsRAY4Jvjqmw+4ZwajyLzRoCji8/Gpd3S/dQ7vFt4agP5sV507CMl0mxKJ0qRUEHYAIqU7u4
UsF2PXgAQGFlreCud5MIX4A4/TGeIzYarPtBIIMtUsNtidoFeEmiTuetRtcH1gPZRjlQ1px5D50h
31uF3s27+45Vs7d2Rhz8UAm9nnzzzqRwK4xfSTtgstDLsFwwG3AWfuibABexXuzGYsGDbZVzr09x
+UnUJC2YGkrZWmEFtMGFJpzRvXISvb6sluGvxa/n3HPoQyQqclGL7ShVEHxO/amHp6ZK/UOrsacm
ZaUReAE7+HBBjDzAAyPqFV+YGhbDwHHk8Y6yy38+Tk0djYpbs0AszGZR0MGKSnHE5HIENy1lkL9X
LYAOIFlxYkozYnYqWKQ7OfuiU3jy5efMMVF1Opk6E98p7BC2/yRuUMawi4LzzDuqfsTAxzIwRLjv
Ja1ix5OtDbXpzlTKOuqrLhdeOFPqHi3j2VmMCQf9Kd5/nUFLMzSRTQcsJ63r9jpq3pNKyPFg1oAZ
PVz3sSDLj+g3bchT1SfX2dmzPotKeraUlA7Ej5BE2OwPPfCeOqkM4fIvN955rKAV5T17s3bN4514
zd2XuS4Y5Iirbql1GaB08I7+/2FZTHtP1uOiS4OG8cFCEkWeiqOWBaqDUdwAOAUB3lHQuDGkd1Ht
OXv54aL9dcH4LXQQcACrLkQRLxKd4EKsRTminCcs1rH9Yxo0LJjQL1uvlG0caV+/UJcAJWBJ59t+
ps06P/jMWb4sttQLMHz+lvINIa11EI6bfTvoslMJZGiP8QRtHTtdMWp5ovgmXoF6bugTokS+mhcE
AeRcqFUVJO29TS6YMtSB89mdqfjc2w0CUfvtivxgTgJER4sKq/+vtdzx+EidX7j/1FmH6NBiQ/7d
0HcfNDJMb9UoCnsnY+yYO3ddlbLT4/8wD+el22bwPKalY2LhVFOO1GQ5jfgrS0FZjM2wBJgm4btg
Vu6hiOYG812A+Sgk9+NPtlmTHLKMFY9LVKuUcp8eDKwHbk3ZLbFycv7/NhsgGLvRvfsUmcuPVTrp
pqXfNsQvzaROeOzS6yUfeqQzw6BX7Zx68KFYlpgwZXxj+mYpN5clg4OUMCPsYCtLcF4Zy6jk7qYI
ta8BnzABRhNnopjAYDLgaXh6qg9VJeZGVEvTibZQFb2730b8S1GnnJ0BE7GiuU3mdxaQP3BwE043
vNx/e7pTMTVdzbriM3QhuXS/0nK3VgC8R6C8Q0f8HDEYkBrIiz94V12ZeSZJGSCER/xjqYNkSIXx
xLV3JOwMNg4rQx9mc8cjGKq8zMblLTpNb/ny9eU8WJD/x89K2Mq7AV62dQgkQKCTk2BhhA0JX88P
BgCzD9WBcnXBqqVcTlY+mm4j7dAxuSY16tjYE3p5VQdLtemt6IWXIYUCUIQWGVbxh8ipGSGR7myv
H/DQLvBCejPiyr7lWK6wjm2BRRJItEd4iJ9kM9/31PghctTESGWhI5MUfDZfrRkEISIeteBHJsmk
NcE5u3zvbztkgqrQRzNLnTLJ0yfXVgcpETICdigCxOcIULtIGTd+rccqZzpIpIEL+ByLuYahNiF/
MBYhtxQsxWzpa9cWsXh1ck9Y+cK/B/G8YoUdlFqAqRD+7zzKHS9D8EWmzknKHl0neJLaXFn2x30f
7eWF6GCf9JErn+PV9bUF7zEE8vRLzyVKXaQ9hpb7hd6WdYaBc/JF4t0JN1U6oPq8I0xd0sOvQzYb
kEoaZ0GGDbKNkPftgNaZr/F3nXSKKW2xc299CuJkIULXjlAGJ9ygfTOlSvzw9iPT9KhW/SILthaC
mujU1OcgHEfhHal22T440llmKthL9v7DDQU8O/NoaytM7sW2V4/SXvOW5aEOyRHP5PqW+ddS5afT
tY00fVPnDv6u9S3nn+KcU+ipTGzUZhiCosyJkizkohILysTyiuptw8Lc/cTafyRmWY1KX8xO+dvX
SLffoF5347ca6gLe7GgpfO21sgKMoU4Eb6bO7iT270lRiSZPPcdlR46u8TwAYRy8UVpte/ElHdrj
j8DKsYBUcgHSplkP7OvkURPyiZDjy4JBDOnS/799mAyPSiA9Rqbwiatkw+65VqHNP1sAlQFe4vLE
IIFqL+j3IU3teT6V8PQOdn+IcFOsXvaEB4k8ng1rDC+9kWegbTY8xcB01GaqPMjESbb7BsZFTBs/
7GAbya8qoz3ubyp9T4IzUZ6AAkM8brVvsp55SYH2G7Pik8gxxUlsuF50PuUeUaIqILx1tyeFPb8U
XJzBL/fw7pU+ZyNSEz6TFEuRQQjKKljQ9XU0Om95/c+Z08loVp9TBjQkzy3THLWaJHDhY9D6D9Hf
FXDzTDvkCePzJgjH/X49WLqLsgemDybcZSWy8CZwRL0Z5CY4KRFUMmaawAQ8qi07ziwjFiAyaWSl
t3+rerfKplgds3/0VVVg1JxHhUdhRpvGETexNgz3lfn1uWqmFXGFAgq+IPWnj58UiOiiwWrcCmli
XKqisbwQDAjxBrcjwOA9sBTtRcDp4ZvMHjR7TUTF4kt+B83hGU57Y0QFabKrMMnqgklHfADU9kpr
a7IihJYicA1jw5w6GDNPjDIOypCOQK9Q49bGsjtf9MSvYINg1ilb2OeV/Ui851ifpY0X95ypjnVv
rTesW6XNhm7ZsWcw6x7j5po2EQ1BFblQ3xNUJfXcX9Xybm2mv1Z2XKYTWWVziYG3R1hc7ztoZVCV
Lw6kVFZioQ49yeb2d/RazIzZrLPD8o1v2RUSMVcc14WRFvJ5J2R6Fth7H5LQKIU8Kgo0zLC7WfcS
07laig5siXgAHCMZfwHq9lFPdDUgxCnJbkgjMP1Vb7CYIRL5TstvgDrcKyu91b6f+Lb4D2Xsb24Q
XFioVdXDvSUtYX/W4eg/7xN6DzDMBiS0Rj1JwpesY9EHMxIyXxI9p1tMjagEEVUlBx8jqoONCq1i
A12pWB3ViPhlNIU+4kfAp+aee64FCYVuTtZVVJChRkGhQSswqSnrSbFdiKmSpfyBHKLuK3Kj4p+y
feJ/lmDD0CLKpf2KgGEMUAsx/lVjc0RM9QRSWi5zrmwBxOurtUwkDMoyUVTUpq48RBty+LoLJ0V7
5wK4Sngg6uPV28nkxBy535xpTp2sCk2kthBxfChfYI3NbttjCJ5eLdbLoHX1wGg90dfzDbJMwIl1
8ukGMZzj+paZLnklnDD/ynrjW7chM0GJ0YLboDXeh8+Q9oF7wUhvCYW43svkwvy6i8bXRios58sq
TBI5ncb+rbVIuOSsl4U/zEsv0hbaLm4FngnozkygB3gU/yQFuh8I6KCyLAtHbIvyQtzffvIB6LSB
eREAvwwO0R7k5Bdl9+D1BpMpfOMydbcS0uNGTmr3GLPMKG563QnWIAuYAq8Y+HfWl4OzjvyJFHpU
EtLec7U7aWLRVrTOxowxDPdCqbxlo+wniYV7hQTCJRsiRPZ+5BnsxAAbhieuazGclONwKIoLWztl
ztF+3mIGkVPNq4yc382fjNmPxxae/9+ptiKci8/hRVu9q/eLylEjh9U+UN3SpeCBRRLxnmu4vy5J
aQsu1+rydZ701dQCW34a2gb1EiBiMfBNRho10q938CVRYrhHckmMB7wgsxZL+ZUnKCuIdCzzUpNv
/a1KIS5BmCkV66wY8TwSqHRaLiMmq5xYjXIbqiDa66g78zb85C4jXiHRAGz9IsoSgEkUCStLb7n/
F/H84BXTbWBCJK3AyojAIHGBCfNVrkFLL4M+divz+zJ159jHekiYs9XwIOEhYVhsPAsWsYdpWyHh
IuAYnXYWP5e3sYWDiVo7iPUeMCOzcZXxMjYoDtO8lb+FdCPKmmCZV2a1m4TGYRCggVx4E8ogrBzU
co9n8XXrK0W6CjB9OHWwUmqylmsbXMcGl4yd9xjDNiARKMr3G6vCSSpe+Py6/zAzfGgpbqKZYTsx
zIWEic7gREcSf28fHXYAlQPYxsUOa89r2kyhna+diF9egKY6iEl4ltkRnZDUvnnTS3vQy22nMlpZ
DzrEFCy8SvY+1fg0+otKfQXlYgcas5qDOXxMHwVWEZCQ8V8wDuAGAhc8yAngUoWjIXpg5AH20QNb
IIkoSczIBEh02u+XR+jVScZGvvC1ldhgNAsMrYUD6Pu9Du1ACye5mJTGCnxmvovog8YJDIjODX0h
hKEU4sZPRCVjtSTdCmGefLzhjG6Xs1IorLwPMO/iGj8Wc/dTYfXey/sgEdqOrovWKB7O/u3+MWvK
dkDJd5pY6yXJCdjLFe1RCIqg/jSqD4G03MM7Qfdxd1cQfgNa/MeRNFZSg20Z0+Z5M7YUbKwu+KgL
8Wq/363bCshNTuX9tHYGlMr8ckZdJbtIZQt5ahR1jjMqBPhTPtb9aB2tKkTXdLgy1XmQG3Y2FO5e
klIniZupDsYXUL0EMT1DKOdspvx/qr/hNQEvSnI0XLJCn5zik9sBgzn0/CA7z7B1b5J7wO0IWmaF
BeFfoyAYw653NArA137dyCkX/VRV8h0K413r6UdV6G89xNJow+ml1JyljE2168mRFg4tAb5dUqYl
IRpDkO18y4jdQlyxWzf24IwM1l8IrR/vA5JergIFL/xx2eevTI+H6kjMjr5WC8DmCJ20IMBHwVPQ
9r/Vr9EcqcbCaT4nztPVWtXZ4T7gaB4DywCNdT+z7NjPefea+t0DsPIEnyayiCB4UjQ0qhfaweV4
ax4TBPd1sH+nfNdIkBbPZJda3FgPjfIQRMfaVwpGvaj8lzY44bdgUQHxfsilGPNa/gDZ2vThdJbC
t5zYvSeip83TLlMvThzBVIo+pqKsi7J+O+fBvgwdj4mQFg82nsnmbczqKKU9OEKOLO64Nv9quPta
2kAfmVnsY14T7qH3XAj9cvY4xPFvaAsTTi7laha3Ipn7Jjb1e/DpiTb+NrvjrOZTWS8jiPmfIUWt
yrrjMXXza/f4O6Rq5GVp61la9A3oLoTn2LiXSg0JcYrTI0pHEEeWV5ZJJD1nvIWdZAclKEryyBZG
jW97rqHsnhqiP/0jgUj0MC5ss77E600vANMcprl+cAb3E8oaLYpciwON+hpf3PIduYwMIHF3RGJI
o0pyL0RIgJGFjMDL7AHGM/7keg4MbBrgBeHrZn9Cgi0UtY75mXs7cbJhrUtw+EgiKKSSSQqZ4PPx
9hUkgW0iU8hyPXnUA/xbe+7mVvzyifhxHa68KmZwg1BZfefjXKhFJrq0y1gIyB/hBhg0ljwpEtgC
4NIna8IIHCKBVG26NVr2G2jscRxClpT6/8YJNQU41T/ie1Q/cUML7tT70nlv6xb16rmefU3m/TuS
vnw4NHGad4WSHlxJ9d5KL7NYnG4pZqpvVbmwf5gVeeiumA1L++h78O7uUT7X3DxZfJuDgBOo54qN
Ep1J7UWu0eCIacgsR1dlrsSNVpKrT9an/MU3c3jRpuOiBGs7nbWQH6wn5+zLW7DJREYown+6L3ZB
JssG4Y98i+e7q1N4oD4b/IeXnp6smCxP4AD5P7Hd5XRBmbk0R4kLvvepjJcIbP7GWTZzh26+Etbu
L59dsblsBmKxAWY+aSHBVlmqnSsoGABObCGze8Ax6D6XewX7t4x0jcIkmt+/1AgcPdkUoUItqLh2
5o0kwUaGKOgDvlev8fC50Lusi5ceplYOc8XQlzYynaI22JBEtsbW7sBt8hXTcP8aXtbacfA+zux5
pMugJnj7JOMn7OMzZG4Ji8yHH0YkMA2p54cAfV7oVdbMWYh6vMSjgck0V/+8HPZqsQNEkAYmmDA5
AMuWXx9if+D+rJz97YF3SO59F6YNY7QlSQ+fNoSEqwxP02matiqhefZLif5i18DZZHl0tpaKCAlI
JVUvux0ugiiTibVuqM1VKso2OjcnAYNlfneonSfE1Ym7r8LZpTNAASvtPrAepW4MeOo5Hd9yhZBc
3e5xlWrg0e74187IfLgohU1OWvIsApOeA5JIKQaDCeN7lY3/3JwO/Kly/KVbzQ/MMoyO2HgbanUB
5KXwCUOWDIuPoaerqj8/CmVpaFm/CXG7wE3x8KeVmhzQBd46fPst1WVwnj9E93Wlr9X6fwFJ/8Fh
mxGYPOpiF/hpIHQjpum8bZzJ4aXarX+Qqs+ozbF/7DlKb31V4n+9mPDiAV2sNs1Gtdt4OJSh+knN
k4hvwtJg2s+IY+KMFv30mPf1XxtskqB9EXFTrxYEQQbUeNEhFuTrjZBQWIyD9b+sExWyjHSpD9y1
TUA6WN5kPajd3eWgBQViFa4LJ1YcMm5gZGeqrvu1yAwE4cQkkM5lm4iMsmUQ5lAl4bRx/lO3UK//
+oVtPpvVRrlhEUHCOg48NWiSLuURfn2oVmewW26Oopl60dhwIVpOQno1d12yG2TBHpYUDWJaxJPS
qJyinn8QsZs7wRaMzS7cxF8/RN1XB/slwh1zQWQUponyRHNILTpSvr0a6vL9m09I51t2kLnRGQjk
jYb/HYwrXaV8YhQRaMVSQqjCorD3VmO6DdD2t8Xz5D6mdykzOmXtPgq43Qb7GjqCROZ6Txd/9eHM
NpJ9enQFYo1Hfiy/bctTyo9AIvjx4VrmCfg+0EeAoL14j3VLib0TvP46F/lDI4O8CPNMlq8EcQ+V
2KPyQnRYU51DNeFa+oAQ68TZODgu0oDUAofxfjuTV+UfIc1w9g5XFIdmPH5vGqN8R+0a5/jtyuPo
0MAbgeHSAr12GljR5QPxxNLKudqd1f5iV/d1OXQdIb1Xc8k3K5mMjCJALYexqCuDUbWM+sVdRBc2
BhZto4FxVjhp05NYh3fggEte5USlR47Wjm8Z3fZBGX2TXLQ9cQFtLifYcd01NKlHDIqJspwEFZXZ
xmIYtrBkXjEtRrPV7wqGs5v57G6znrwzT0lvO+NTyUW4sDiZuHO/lamVttKANuBV03Q2CBkkTaBY
/4xizI0e73pWRfObLV0DH5mkUvWc4xrvAvLqhXe4lC0GZSd/0mbYI10G/uNIyS1kjIOkS4ywUDaM
hgAiSnHkQPqxw5+BWlT8ZxObzKAeoTeVz145bWSaOtU1LzQ59ynAIBQj/znFGWw8K01FeeGy/xsO
IQUPT7H2tJdppTWbb7TxR1uPJfiaeMLe9VwvYius6SuiqEwpIVm4JnVGA8R1DUkyrCoNy+bBVj/8
jOT4KCoNsdexy741ZvK8nle1y/bW2xybaxHoScXL+dsXG+L+yrbPykOutELdmaymS4axtuETxtiU
KznXPCSQOcsy8QNdOhqXAxNPpB2zTpcLjjiAPbFK0vb3l3iQbl9WZ1BzLpPZmer3TH4HJT+KSuTK
b0Hp5tmQ0hFbx71eNEfaXC23uF3MF6bW2vOijZjHn4u1KmNz9Tlwa9MyW82ADbnBOynwoIK9EkwP
cfmptc+nbJYwveyVheltCLEcx7A8Ow6eqbdjykuHBBIH+REZLMFMx244cVc/+dlBCZl0QZRLVVwZ
w2R4mLSVxSAIe1wgEGNgsN9Iv/2S5wCa7NuhxJ2IrZHX9wJs9sZdXawixAoLxW8w6/XD7kqaT9bm
PJptvliNyMSgHXIdinCVJtZsB1Zurxp7OBmYpyBowqFYp4sBn00niIuPDCeHbhBfhLgXeNv5ezJ6
IjZMlf5qHwjjC3EAlR0hVtMJkWBqfuqQv2St6K1cJiKzUMZs9HMo/oQUWZODbLg9lXwOXt5XSJMP
IWRgK83xZS7WgxaAhpqr2iQbtb+t04nH3v5Vfi5z3yaiAHdjK43AR6cD9iXR8rN06w44Wzk5LxOs
q4w49p3yLmRqG4RyIWFLc71iTwN1ALYwMhMKs0Sh+OMJuCr+Bb3DjHRkzIjQRBXP0r42go2df1eD
XSAQlYyXy9qyHI2ZR3TafYIvhFLs+zUmMIqkHjL229pA0tfsxvA+E//vRFQQn/o9EtE8KBLufglc
5gcXO1KY6v8SqFWSw7XjpKioYJ7dlAIKjkkiA2nZil/xwfxj7TfJOT4Y1AeLf7E++8bxPnfmH29Z
bcDwSSS+INEMqfFkHfk+Vnp1M2gzLCIYhazk1C5WaRCn6TGjURYNBFHoLuYBWTUh0ixFyZ5i01cN
/xOVEfvH8247CBDORL8XBO/lDSKCzlcnbYISaP0rj3UW9yEEVBmUpin+dBRYPfLsjbA1Cxf95OCV
Ph62E5SjfQ+dcRLU4qqFLhM8S8mt6SoeqBx+4WZa927rj9jmeIik2DmlOsQryAoP9V0gAfKEBcFs
hVLQr+z/KvmtQagWPMcsrO/hJ55S6Vnw6qDfDfq5WeyE1zBnkq38DCsLIEo2sMZHqtk8I0C+cMOK
FmKc1VexakLAKE5a1/NakwEbi3vcWCYKLzfIBNuJYWMsbwEUTRzsrD68Zg2Onm/l078n7qZ7QaeV
MlTHP2YUXkZJvheMfkgDlrgpLEWy5gIH1sdaIFnjQlp38pTCfgqqFuU0zRvxWBQEFDOV1PQ7xapJ
oBZRnuMgLf+qOiZGcGnGDR/lIXLoxst5XnwacUC56Z2Ghl7azHkASbBgAVmffLGQcsc4tF5NAQz9
YF5668A3sSYFvBWd+bcrYM4qKbTkwBSOJLm7pKo/zWLDimXBipp/y1J0xZrieMf4ELSp8fa63l0z
oE03lxGY3Ym0Rume4d85IL2j5KPAQjzHdnq2rDcYLLaXudRBXjHTdl/P8bJ+Fz4SV9VoQfsLbEju
daGfYKflNQBjQJt6qjRztSEHoMbSpwGBA+nt4fVQMBagwZFT79UNJbo2MnybDpipqxwduAyEGpgj
bKYJW9LUBAbeFSB/WQigJz+Yro9+DYGt4ODqFEfgPo+oMezTI+gdurRzhkf3iAWW6p5HFLlgACNV
8bXCeCbZKVAxtXnfyrYDNVA9Lrz+Lm3+zdH7OfpSOWmeNr0tcC6RE604ya4qV7Wp9P2SZ6gQ2pqc
CNAFYv2puw/pXiT+R+DzczAGwQqASPixBSDmIk8TUtst8C6cDX2Jw4TeCjRQ5k/WH+nRxPni4h+M
zDRpKRGjq+PP6q0pgQjS1GAP9L/sCxN5xBFo4gi0FU7OQSK3YyDcWitFLO6WmgxrAwElWe/H1iAW
/qzrG5Jx7royAv4J2hvZGbkaiJLMDTVPqIcdy2l+MzL47woEICqEC46Hal7UoS/cjQcLY+Lk1MvC
bTImssPc7aZNVBjPQRJkGPt1rvnbdBieL1x4+mN0d6JakIjwlzWMNVyqtcDsAjC/BVbLjLOC795N
8gMHQ61OmbYBaE+9TNm861rfCzsk+2ZoWIq3j+px9kxouQPD4E1vlh416WQVN+5deA34B5UrQQOm
+cyD8A2oBzj7tBpwOGLjJFBxLBLFmsiQvFLHnz/oIMRJH6Lf1+xfUnwrCf1ir+Na3Mw6Vah8g4+/
+eomQCqGDLC9c9qct0s2edgCPS7V2B3EDXk1Sr6Dv5lz2tetqHW/TJm6N5SNejxQm40NEy+tILep
nYtwIDkOch0BYIl23HeGpm9L/2Z1Bke4I3RY6SI+ENYOJvTlPA8o0oda1bbaEO9VsiGyiafHNPWV
4rwXnE6RV+NpqbBNT4snVqaHRUvXSgXJnJ3bjIRm4vw8Tuhxkq0lJrsDR3ntEdtyU9zzT/ojfW8H
Qh3maZi4g78+9DlaCG77tkSYG9XHmFU9CEhHqQmmBNgxHES97PpueMH4kJj6gf2M9taw0WhfzV4H
n2+v4wRgWEJJ8KOPFTANBvdQXOO7Xv7k44jP+2oLlp7iTKPhlzHDFGKy73ek950IxVhwJQEd567Z
sbR9tUsxa1kf4PSUQT4rBZqqTb3HpaKQX2vtOnYGAGyuxSC7DdAiHbzXFlRVyl2wY13fMRmS12f0
eiRwAqgHTr8wQhz3E4GdYU2jK7VKuzLn5voMr6W9Yaz469UyjseeQcIT/nUaYH9ziI+zh8B1M++n
QBAQGTVz7NIBAn611Ew5AMuiMBam5xAMDjDPZH6uKeooNHPpApc2yHV4jfLtQ1hJoRJL/urb3TZf
AFH5p88xQyK7W+/UJdl61uK2xzhiKt1wYc9y+VDv1R1JfBj5RQjs4SpjfLa+0Jy+/d72MNJqT4c7
aXxHCUT0gWw2wigihwEDnKGlbi5pGBVQmwavv9Bozc7bbaoL7K1SK3OcdMWXnXD6bDR19wiKvt+k
CQ2AEJYTOwUNdBQdy+VpnRCc2JMOM4xVW1M1N5nSeVVuGp7svy7gMjTTg4GK/r2Y5+J4KxSk+Mdi
uFQm5YbNOa4x5Tcl3l4Kjt1AMF8A+DppDF9Ltc0osmr7+R9Ef216lb1S1ljMo6htn7tyvZAl/Vd3
0L6A172St1JUKkhWc/fC3y4loJq/GzsZRZHZQwGGrUaF/cR3LvUR3sJLIDaLoeREAwreQy/LS1nq
E8me9mt6Hpk9I+tR8xX3SN/0Vt4mKCn53Qs/9HvkZ5seLZm4VbTMXrQvVljS29PkLTW2jBEGkz8O
CAT5//PwoS6aS864RQ57nB2L0hOTYH4qAfiEkOMH5HjPC0Thl5eDq+YIZriSeXP5su6oU2pjFEKC
EwPHyH6Be63fihX1q7LZRJpOGhr5z35kho7jA6SM1701odnr6eFV61ZOG0QaAT0qrmO5Ro/Z2wnO
X5rhVQ/FeSD/QFCr86+b159ufyLs9p8W6nIrS8ytiiVAVmloKqejSwM2MMaB2VqUgjr2H+UoZ7jr
Ggh3FrOqZHHo6sWKIkYj8ohEv4cikYUMb/bpjHGzJdJvGu9USVTiR3gzz9Yt7Bv2lfWg3ftuuESu
9KwzFO56YrvjqfLI9eWD4gF6RVIKhyrN0pWGCMuZq/q+PoRSJrAHGtu0FkzS4kuiqIb2KqO3nxzX
ZJOfuZw6nFDWH+UXCidvCA9y7nxZkFaW0TJvGtPBzKcZeXtaUpXJ9ImnJ+jkqWeVcolfUfV+7up/
7awssgKQ0MGxUgO1Cz/Di8pUu1aXvG8HcC/KPmIDeO/NHzemPdTV7DeczYlV/EPVnsW15YjAxELl
6e+QeOdHelyM3Kwh9I1OhBuzZT+7/mhji1kMNIeATxLFWXxJGOsjf4Y0koAfav0GrMcdXgEnG4ge
zUtFodu0WCsl+D3DvTSprIixfFZwtlEbjPBg4VFZzSbivPieA2DIaMkUbhUttTIG71UiycXbKUyB
MIgABUOoKMTqoIQo8G2Gh5OgZRtMXGGaI6H3XHlz8+sQH3ybT0apRaTXaQwzytybcz8GRDaxLDVc
Hu4u6spyE2sn6hJq5NaPpQJfCSRku/rXQiKYfI/Vs3QuUfCBb4kr+wBhLFF105DT/02YRPLoy1p/
ewXLsfE/1au3CUMv3oixf0wf7Kb9DhgARRQ87vYVLzzKiA96owbaIKvdzLiwpXXAzo1WC+Vbj+sz
Kuith1hbj3jRXsj/6uaBewEw4KFYOYziWwgowjnLhUsvqKNcneB5+M/n7NV2Gsyak3zJaiMCNYrw
b7BDELYhIAxTARDd30QcNZQBr/tI9ys9HSIZJUqt8V/l8eYymyXtpNWcK2/6W5AKUXm8ltVFq8Se
6iheNMO9J5LzDR5E1cnOqxFIYqqs/rXphUYWdp8uaGoZVWO1hOQ5lDPISTITrllfdUvNawWE/Lj/
cCp4m6gnEYHHLoLOcI4FfSyVRjMAHt14+wy9uIlRVFjbeZrKtvMFXNfqGBOTrj5NmqGPcHvnjixZ
7GVj9QYk1NXnQoCAOm/mM50Trhnqa16jBAKUdWilyAMjt3v0CbfpQf6oWlTavtUihIi2ATbpZvYY
BU8n0EN0lrN54yPoiE1kwN6CtXGg3WxlQXfspjpMJWLeozDlk/D2J1q9igcMRMWAmnM59t3dEn2G
lRayCuVsHV/M+kpezjothbGwNOsnqHvQULtoKsQ1zE0aJOqZVeKeLZil050mLchUzWK2pnZ8H9vR
W5KlQjS2fkUOsjcxX3CAf0StJ4G0N//gEBs9pj1Cz34cxD1f8N7SXsS+ZBLzhOuE9pm8dKjtuASC
g8mJfakiEij54VWI2qBWzGXxuNq9hKNxVf2U1Yg88ezpYsSnEAswoGQr/SpBhltQFoAiv74Eb3ia
FNHWMpie4hCtVG4gPO+0XcWDDB9sWWdS+PXv4VbsscWRlIR2cTIF/HaXIrLWjUr7QSHynZ30GAr4
f8/UvdwiiUcMO3AmFqDLnOCRvczXj+klCVcVI7VgMsTcQHkzaIN3ixF84p/SB4dBVnhezguY6Er1
z9cDaIaebzv3MsXlgijucSR35ryXtntAUrWFdx1UFufbWP32I8tw4MA4zspngqDZzzz6Y4XeQwRw
PImT5WHflubDFxKQzbU72jYJH9s19FE0mvLC6WGbkaK+LCjiJ4GDACI+ppWx3yoWAqxh+ARcbUeG
U4FMtjdsmg9/uw3mVGQdQFtzfFMhmCd+ez5+jkR6eJp3rmRG4495jq9x5rFE1EOf2voSYP9i2Ey7
PwALX+fsRftsmrHAwZhul91fdUkFg2J3lIFWTxXtn6ZgJLnr3fSCKuNhDsWcjrJqy15LfH6zuX2o
FSM3MW8lT9iDom8LXM0GUiN7obZ9MtYYKgf6dSWhQHa8reg4t6WQNwgRxDjnHVjNB3RtRHY3scVh
rygP5ZbMAT0JM/P5F4vntCXVJT4jQ9hOmuOUOvoONmwMIX4ibChhBi6GQeUaJxDYxmIFhqIVIViE
YqKAEki65eSBA1TNMShqai78vijNMJ4YHdOZWavkK92lF6dHxjmiGQQchpEGfSQvA1PbgnaGIXa+
EIzLnxH/qQQG2liokKunggoM3alq/eZs7eI+q59Z1Fg7f/qvbcFoohJaBOtNa3cjcNCAzf4/SdgS
An6E7bp135U79kJsbR5GalSv3DaVVuVJXtTp0TIIMgNIfJR7isDXnZFRvzn0Gim5B2iHiZ56sYl3
PHKDfO5ahvHTW391QQfqivJNSQiqsTEVJUvrqv1IMjH003kJ3mHf8VlcHvuY8KMRAnzIJV9RdYc/
D7q/EA0DhGrczmq1FHTLcYrR+5MObDGy2Z70MgynAynYR0LACn+ogDtjgohXd2DBxK7hZ5BxfVXt
wblbAh6C1Orq59FSUQaD1a7pzDedJ33AVv+sgahgfdZzkpQVJF5B6nDmfm086gOh6EubXE+EwOnR
Zs/zQmnb/K60nCz/9S3Gf5odLv1Et6trgQD0mSQOAG6qeSYhwuALZRgzuxwHyts1Gd1Skwu8OuJB
OG21EUzL/wCqf9hxC5WPfIEZ5B1Heroov0kLkSDY9N7iS29cI9yNIObEJb+cL+blN2hW1jNiJIpU
UKO/v51j+DDHDOYVZ9KI70TlkQEiGRTpEkC5v6L15wjJFJacotxBfGEwdiN8CwdbhbShSPGoo0Gn
astmUxW8Rjm1qy/LUapikApN2Fl6jYgIl0DFe/U8buHzgbfiPH0Yijlzsw1HF/XRr6F4dFIIg/ff
gs9pPpWTRz2kOdApxRIGVWmLW8GATEbQ3JERj+Bk+vgK9PMA+Mo0AvexziDtndMt9N/m7iqC/MbA
HCbnj2YYeArBFtmUUi47Rq6anq4MYDLC0ct4JdsOOK/sAL9q2HPSYzLlUsN2nkyFdvemHICh+FWl
fySpZZwHTYk6Nt5lAnKFpsQQmslNo3+iatiqcQkWj/vCLS7MBet9nfl74mMuN09B0he6bmxuaZ54
vDD5poj60ypa9eQeGcMjxj13l6OlA/6tQ4mIdPNehkNvb344YStmZ57ESQZZnbVFm2QCitsSyHxF
YpECCagaq+ELmcOxTjKm4wtS+5jBvZdcFu7JEK4+2h6IF63rdCvNK7TOkoiX3X27SCuG1sVtuOai
GSpn8FqWzF+pV6fQzKvc0CU9IC6v3q3eIo2UQNTYfqP12KUryQ6lY08+gvPkoO/prtYtW9tCGdN6
x7OUeFcR+FC4AKOaDGZxLBo5G4wEXbf26HUWlZQIZ0LRcaJSgwfSCkwiHhFoyodyIgC0t6E3IZWa
h2YkKX4V9mL0T7F6fwtW951XTgKxaQUF/RScPP4IPMW4gmKowbpmLdZgPsnTRidvPa+8GDfD9dec
UPhZSMkZzirqn4sf+bDsd6tohxcTn0EAudK1hH2Te/CnT9+j5YAp6uf4JLysqaW3m25xYhcg/hTd
JzUteWA9UOMficG5PRw6IXYTvc4UrhiKYMHKkZiur9gaK52YOD3bYWZ0IGTAjy+6eXZtFYA3hZzp
rhPz06nj4dYzFW+lYpMO7gPCSoWEDCpT8ulbVVo1SLBBpK1W1KnJGUH6VJeAbJAlWSqpCqlAuW1J
sdVSPNREbn0oYoLt/mbVEjZcCIIQfMOxWm8kPGYy4klnmaOxLw4kxgbszPjp4efH5RmWFkNeYK9j
v81jLOLNT9FeLkvGsLT6M6RJuww9eqV9KYGEYuTxlhXxr9O4XoGU1TjwaScdCei92NbfQ4yok0HE
L0NTv1/c71vmKVBFulwYxP+41bw9XZnFwAnzgNrCz32BObyVQr5jOrnfPRYyV0BVytVMH7XS/yGk
x6fvLpaJPMUgWLEXgUFkGsPqbuP7f5jyTWSYIlC80Zd8yu/2DFMezt4pz9ykiFC89hSkEo5CWLgv
Od25Xz9BiDdlPv+LpPKYqd9m85F4zGdeKKj8plXSlKg4CrIfYJ+S1d//Vk+TCteWEa/Z8JVuWlPc
kVs7fUo9CGYVUkzi5UkvAdtuQ/ntIbrZwCarr/NsOkJnxE5ptDqRS7mLzsCIalMAYUgxFMCrOEh3
O0aZyAHY474gFC5h8yh21rFNv2xWhwOCui/JcVdOUxL5Z8A5WJ7o2CYGVjLjHNCfYAuFecM5KdB/
VJr4YFKL6aONw1SSTjsvKk+5m/ltiLXn8nhY27ScevPEc1iKVBqI4P+DO9r3gxmgiydln4qWQT38
yyl8l9lI1KvUXKBe/Tvsr8ZoLxIZ2AA9rU6soki17KSGMriWISSe/J90vUinAdCvzSY0NCQwsRhV
+le3c+T44zA6ifYfCqvOpZMi5NyKclvyqKs2zhDWAQkUEECtAj8QJfnRkq9+gqJ5N1Ik0SGljPWc
WfQa2OJROFwdchcPridMJ93Dcpp/qGshz5GgYW/eYHdT3+4oo0RvJXDa8DuVaytCLbVERBzQBODg
FThhJm0GTcwm83QuT400PNmQX3kRgCtJGCCN785DBKTtj7CW9ekF1KmDh+t5cObZiHBRgp8m47t1
KjOVcXizr3QlQ8VfifQ3fd2UqrsehX8xdTiNXdQ4i7i/F5sLZeqiYmtuIPj+rJOwoxpmDYW4tmni
xXssr4YlI8ST5cqquHNfruN5xj95oidWrv4jK0evhIIsQt3FvGGgUGj91A1g/in6lopCB4IVpgjO
lNQgUiLiUXVDz5lKZNawbKu4xFdmuarGrZO1nIciF8Vv4LhBVKIDDD8/k6+GInF3dlUBIb9Zef6L
5J9uUBY2vllfPBEurQrD03vQCq3XlNYF0JOHTOpreYyp44wKZpCe7fXBEgjICjk7PPqXblOEWAn9
EGLoIcp3rYaNu0+ktiReAWKCQUMXZ8auQSmLslfWXJFTM+PsUcla94riyaOeaA2zp3ws7zvyKwyD
b1QabjFUs9PgFXXuXm+R+/YEwv50JinyDjd9gkM3R89cWZPk9rulNnO5DFtR2/FSpI4NGtr/rKF9
Kot0s4RjC2jujM51P4qz9YmCjCEaJ4A1eKs6Dwj1THadwhO3wxPI9cXFS4KgitNez3ZAeiakrXal
NgmRGk/C2dFxNBEuY8OVXZS3o89OZU4e0/6oE5EFFzkpkeOs4RhLIxuppcjWjO3YiPJ+QQfsfPqP
3eNrnNOL7zyB+luv1BGxfKmVj9k2pJl/D0WIKhVrIZgLDt9zQcmLqJq6c4UC8TyVxINtKawqJuXV
HEI118FFkVqe4IKvl8+ArczM7fnJjiOAq7RLpt68bTLtPANE0IN3I+rUFLASzM0z9TZOv7f0owrt
CpdQaV6OTeOBm0BHeceuO0u30afRC38Q2bsPtmVSvUwcfkSvwKnVGnmWQaShFaJNBKYq/5uSY6xF
xzk7HdlzSO6bU1H+IKQ0ojE1xnsQ36FMCnK83SHp0qSWkwQ9ie8nKPuaKaBnGgow5jFxYLWBnDRp
I+Hl3PkPbkIcz3fqbrtZhdEHXGKJDE3Nj/Wgl8JWUYfs/c/gfHCfjC2Nheiib9rg4fP/1EsHHMbF
p9jElB/rhwfgDZk7fbKlWUJJIe949dryiPyTY3LcGHiP7luwcVDt3OoO4DvP+1DmxXCpbYsGJxLM
rqAIRYAPemKgBeO8wb2hx/E43YIR5d2YPpGjODu9g/JVBYjxam1841JKFUPdZ9WworbOODLqf8Wu
d5X0FEKx0F+P2MULBNmlG09oIiwEu2gD0Mp+Yr5LLNbCjWV/QSQ/Bdx1IDDKc5+6DBms8ovuAgI2
4UQrHidVMFfVKAIe8ro/OpfdAYtaAZseIrjs3AdJzrneQ+NEMdQvebJ9KjXmubeMZQCqALaM9xQS
dJ+2rSw1HCT47lXT2r6WmKpvaEkmbajpSRomK4B67eHY0cnZKdA5CEb5f9u8+9zziui/ooKE/JCq
KSoiYatArNIvvyhjNTlYmUzNtlSv1v/yBD+SN+E1odw3FIqsrEvM1cxWxCmFk1aA0CPjdvZZN5At
N++aCLwGgje/FGxU27DttaFezX3BsIq+VpLBJ0CcQZdw5WgSXgOjMm5xPbg4CAk4SmfiXQ+0vR16
QiYwr3hwPKc/I5Osar1mphqWh7asDgK4RdEIjgxoZmJzNHfg7eFYdE7pMyfI+MM/l0Mk79I3300J
7jeK8Usc4RqwKvRPoex2VOJkIlUol2aKwfaWxMUwgIgeFCtaRllESDwTdfLRfUuS/ZM9T0KCmwyT
IZuLNhEBOq/Yrt/GefAk5IinKFrd9SiblqoY+Igal5yAhBkovRiSrijQi5e8wOs0zL08zuyo8Qap
fVXmUf/PojgcHBuplXnEf8AOlfZMkm/H/yVU97CCUQ3FbyBZogviPlU9VCWxtD4uTjEqJ529h2Po
wigbb48nHBs5fKMZHVa6w1q+DURSAF0hmJg47ANlTVteIqICIY+y099ulbDAkcOMNjNTCdpO7pG/
emaL4VHAmUqTEBGA8Q2udrTkX0WXJsXov51sbqwqBmPv12SieX08pUiCFTuvfmyefMBPwZBKWAXW
nnkS+oHZWoMyFO0yxW656fUj2a6O1CF/B10h4QmIy7/hZJtBacJ0AwwDwzy9HSSTNNJQUnjkk06l
iX8rjoI7BQqMghpsM2fqzSSR/J5pp1xloKvdqtJTZwr6Ulumvi2xvb+87z209PiNEFfpPGPA0nkP
xE8bxzQF5PJ678OOyC8AVAS+5EwWntNM6feZ2pl0w5zfpEl9hG/Jp2DGmsFBUmC5xq7Ogw6OTVcI
KYmzJLC9lbPtwqz38zKWTpqleGBZWfWhuJujHV7DxLnDlhFdcihMr3lRp3XtCwu86lx5XOjzAHu1
O8xBIfYkPXNSsnVTftiprer0V2YrXCURcUU4034HiUrSHCy+v/bAWztZjm1YSjTfNwwMZNPr58Dy
DkX/1QlNnBJYTpi4mN6dcS7f5llVHTbCaSAXyBtUsIPJqJOrH/uMDjWuMm3hKIWrUcbvmRkRG/Eb
O9CCvXAMV/SX2rmkY160TyBctCiXcPWEgFnSUpyXyfIVp2fSU7rbG+Gruhel366Vy9n/JbxRTRnD
X+1DbsIpiqQXE1CdR1awqCXnoi39YeUu7SI1a3kBzEuSrtpi17ifK9OKAt/kslusLL6hyDf5Tfok
XYmAbU0SViCgVrahG3dr/SGqPMqJmVs1eD7xL7P7TqpTIeazDzeBeXB9QuiDb0oX8PNPLBzqe6oy
ax2gt4Fc85+LUqAEJPIJLlqj015+5WbXH0PN24NJF99W9PaIIeGFQPfJU0yASnP3K3asAhb/8Odn
+GJ0tb052BiD2XBgu6nB47G9NcxTCrnliKV0zRNe3avPXxY7hjJRZKfPNw5zFegkkrDZxAAwyJI6
/00n4Cf7vOPQos5/Aky9xwRE/qSDBVQsogijUMboZaQqOKe81TbrTVAbdqr8UK8DLR566LG1Skpw
cwC2XJewT7zG19D34H4Lpo0oL3B7gJ2TSxaMbBzjYlwaTpEYjRB9FiTeyeVf7KoEpU6ToK2P416u
0e6jxbJHQtrerWA6yWy0Rig4T+h3A8PZRXjIvZKOZRNlvH6fajqxyKSu2Gt0milFmI+5OVb+Xrbp
FXLBjj5WbZixuldfXslfjzqYIMTOCfe3IIkbgp2kOWBvEvdnzEqoXl0RLV59adL8q4WGzL/cVtP/
p8C9b7QeDl+SUVJHPDtSX2ndRYIuAYFKJMqJKrRoHIiUPdBdHBbNGhE6LwkOTa9lmUtHIGA/OhWs
7uPQrxNRwJzO7c6MQslKpaP5mNg/pbcV8oSnNysN/YBvYM9X3C/DuJUiLhlsEsDNBn962ntifCF4
OHIk32oaR+gQYMBc6bfxkTquqSNHKprNGq6wGAx4PQtLrRvpbrR2E7/66b5SCK81lr2PhEi3+9ao
J+2sJ34mbf4xvnkOAok96bg4fXPrWXQJa6Y1LQM7Eg6ApWibbxbafZTesR3WWlQNtN45E96Kef/x
SPhhKhMDps/PsopLsN1NUfAShgZ+kAFJAeFx2YueAgQF21lrLYzXfxuZXf5QmWnD5oUNcpo4hmf0
+3gPC8X5Rr5vF2nkEMVCrznXBFMdtuU28PH6A6yJOY/4wQ5IATwVVjAM9CSuwIBGLNr0jwUjvST4
4Ox+KFIM7xCGMBre8sITgcUlm12Gj6HteRMJO4raCW6jy6IfJBjot+aGO3OPGPb7geoRgpFmg78U
M1FMcvRPTdh2tNIb0uRx4rlr1qPEJmHppbAEnjo/AhrMPrpIXxsT1GS1uo5EECF9g0yZlRsFhV2A
xE1uKfxM9uzKoZAdTrK3b9Gl0VvYQqD++cnLqRdFJMZXFVIs2jb/8DF4qN8jQYLHDT+V5nU7nc8I
ULGApk1xsG6Q6Z4uxLggCHPU2UCV07eGLASxjMk/Ye4c3GgTIPn9TzROdqfNDRoFOjaOrQmPjJrV
U+HHlhOtiNBDm0KH+kjVGsbLOAF20NvZSYJE0iYQ1l6ivbyfWXulp/Z8lMBNBHzYcLtsdfmJguYD
9CT6WikNDpesY4Aw7Ox1dR16EEa8erw5oRAvhLariEhJUJZT7fJRTAXC1uZj1VCb1mQktSoMSQav
CCTq7Kuf8VhUB1Fky/PH/9jTXqD1iaRba6jWly+ru7O7eAWx40VKCMUgFFjBMoDf8JF7JFh7hnVP
DIQyNf8qvX5x7G3AELiSNTWc3rdpI+DXBpJ12B7xWf6D2J4Qn5VrA3bQc7jZ3i0Enzi4LzzuntCW
4xTeJ6zmJ3zsWEi5YTyxrUZ10eFKeMK20vae2Y/jXpAhhvmMGqPwT8DehPp+jZ4QuHkl3FSVRX1R
1qTIW1lmJpU/J51N6SVua/QKOb5FauuqiCha4/o6x/rVgdq2S2IkHYPW8iiU18Mh3SHZt6+I+Mrf
ZtsYotkpxkp+Ts31XNxWbESqr6m6Noc94ZuMRtd+FVpJWIlA5047BClfKBmL+q/NKczDhVbFdOP9
uWcQ4pYR6JsJ25PNWKyEyOjI9s5CdNaic4kJ8VWaX/oZOLmvIxsQLZRit12fIrfxJ7RFaJTNDLe/
GFb18S/X4jLyjHwVM/+9M6sqlaY19FPY7NYNfNc0wyMx7EfoZ+FhsI/23gThyHWejdX5sLeCxrPd
hh5u5Llo+v1igVVf0uOozRpkkDjGOJAPnlMx5f4FfsUFdChGiFT/ia5tJ2R7dbrqZliu9wvxy4yq
dYkCHxZRKPgUyY6+a2z1L7z4AYkGFkhZFwprxDvb0qwt6YEjOePDT2Tr/cA5KPHGi0CXCF6a04rl
pHXZ1ACqFprBBi/GFS3BoCYpAncpRgYSwkAVSgTjOwg1t0YgJAaMn/v88uttiCmMyxBAP6q0WRDc
VTiftev7cWlJlphZSuHlkGlqx+C9ZKv1bk5LOv2a//WrbkiO9bi3POWExuy5agIuIAX6DtFvVAR/
YuNs/Qf6B5UcPBNPiGHNhLWJF54W+HyF5yJ0CMnJs7VQcgSqky9BCOo0zkujr/BtRMPuFQZhz/+Y
yDb64O3dxOu/g9iMk2pe7hrrwdEIYBLkFakmw78uzzwbZ2rwWOqKdL0rBxX0dpfij9waA7XT42Qv
XJZfWiILTgrLnUwa55VG/ZwC3cYuHUNCcVMiqP8eTxUM7mLmNaZDZRJyxpbrXe6rzCra8pEDuoHD
GUuqNYnsLScfPtoRYa33jvi0RatqaDkc3tw7LmncIhwa/nqb0E36gES0PqC2DY8E5ygeWbVpCJtx
wCaysqCkzYLdEUyZA0jQB5qUQ+Ytm2IjzB3oA2THHXlsXdEl0duVT4TGIXVQjTrGbSPNTL0f2Q78
UeRHgbiXysk0oHdYZdLVEBLdkRpYtxSF8ZOKit/vo0ZiFAsEwOZ+yltyPGhJ6FNyfaAyFiK0CxEw
1WFEg/alg8RCkMFL5HXFr/Py5W4hoO8CzLz5gPOpYc31AfAV7Xn/AhBA/QvWk15h1/kwFaPxU47x
yiEwZ2HiX6zkE7lTXexUG6Hfs1xb1xbkYhdIw3lKEhKnkaES5BLet4QBzN7VcbupH06OpU1fVjqj
D/Be1X6+hrwnL12BrXXBpGdZY54zgvs//klimj7Z6Mi8XTjKlIIUliWQGAXvyDx83NYrQvslWMp4
6RuBjVY+JONu/Xse0NYsvlsa1J5W8LCNJz428lSwEgK0wkgh8Y0FeFLvG5ITiS4DSQzw0aNX1GWF
KR/+uV1Jlh7CRzi2pQQHjW+NnntypVCWGSeeSMVz5qnqlnKjeAj90vmfVD2bD2jv+tU7ZSbZriE2
W0XQRvAe2JYSTGFMMQ1P2rfw6Ogi8lfniPktDN2g9pagU9v5w6+sU3DF9EqhognVSpkSthY8DlmH
btIXPd7X4aJkSnOGkogXY5iQcAMvhuC6RfK9KoreKQkVcNv2Z2vCwn0mrrbXP3a37YgsgoJHbvcL
LHQTGINEiaSFiApbh0ueh/+/YvdHLN1CZXWq1cI47xfBIIERpZV+5MDigCsJhKfJLOuwpGdl+JIO
3SBR7PhGtVVuaIHlswfu9Pzxbo44NfMKqBZzMYYhlyCr/XutQwSyfuVICjNZlPuIinOtjbBdWliu
rg+cBrKCl1E8IybGKzcOMPD2i7D6WSzQmfszshYw9SSLb1y0fGiwTtqcTlKvlzx7D2la3rSFZn99
w0ULJ/yr+fg7de5+EIVUs5ZvydWsc8rn0epy8lAusJDA5KPXFqEcZ9QFB5K02kjQtBgg0L99uazU
fUpJQ6eVVgMEpKiQK/cOCpMYXW1FXGDLgDlaP3U5PQP3slffj0lHpP9AbW/tMsUASXnBIU7pJpbD
xY2MTuDTNz7rTZwYsMg66j3twAVQAvGiO34hjOIwkfdVk/+UQ9vGVf6ESsBI509MUukapalihkYX
A5Snb/PdcSDOGlKxCLawVzbIg49r3rfv+YBAtiF+JI8O5OW8cq1LRLnVD4Jvhbule5oA5lTv9xg0
5Cqa+zyHX57lmQi1LAE9lX0U2alwQB6GiXakHzm25O2fe+lPRHdZcxRwagmhYiX/WHKqoLIsJfEf
OBJpByByuleg4brlvRGttWRy+Txh0OFNGduqowceP2JCmoEPiHmOLTLex5zT3JV1tgVXtPBHLLCJ
PQb7u9Gd2cqD2OpNmAKmg9p1GI5WGPBTLm5kor+4GtkVZDCqU2B+z7RBX0HEgzUmIJ58J1Rfal4M
+jIv2TZUQylKca2vW56oAtV3jCwUEjrSxcQfDiSxeVrZlqkEzGtVctUWjXAvqxNExAuWGzwatQrQ
Utyjans3pyR8kQGeS4ngT90BYFzFQjgZ0/ih081t5ml2p/kqp8wEEtaBfMTTcW0l60XJdREPVKt3
D0ljXBAKrkkXOlGIzBzhJv2RrkMJPyX1Vo+ANkQkto/HNbsquzVa5kjqTcMtcSoElIGDGqmPcK2R
fa7SHX8bKGmC8zA1AHLKJnD7ynjJUNxfI/yS6PQWv0xJsTAinO4tBDZr3teCcX2Vg28R/v53DtTC
8CrgygwyaFIAzNT9sHs6XqjVOedxsMg/kzNfgu14kadG5sY+KWxzXB+XBdUNcgT8044spgIfl8Os
1i8WuDoDpnOdGRwQZwBgcH0sqCv+mhdCy9RCVXgEZykFgwA/lcTW0OsjNMSFCrqdesntnrEGuhPm
gUKB0jEcPc6HfUS/zMllNCf/VULkrv9dQoED63AcVrTZI9k/uiIy4uYhBtxT/kB/6vLT3yJLKVa7
f+Q2ZvRd8rNc3i2OAd+OYTZyKSf3h/biFyxLXd+e4/SVkSl6/GX7mLOVeqJeWDMKa2Q7vdoypK/t
LAHZuEFvDq0IKqSk0ggWPl9apvf+N2XzH5lPBwn5bLlCAHWWReXjiMdwHFLXA+o6I/ouPFjWXJYt
1C1XQwCRqp+720wVRag+7zSA7SmVWD9XHypOWNYLjaQ47arWU41ON5pnQGI0hI4gy0JI0NSqv65h
YMCi9kq10hh3pG6aPHnNDzrhKVRJK3tkRkTSsxFWAG6q68Cug+ehT1WNsqH69JuOhQvQNFJe2a71
L+hSWeWqEJWDbjNUUumoU2Fd9LX6YsTR4R243N3pC4IPTLZFg2tevGTrjQAl/fQX3l98Q1zPqP/x
kLQylQPq2vb+yT2aLjrhULi7ZCyySJEk2KMfUGip4qeklhE0V7wMSt3mIUqsGfnnVE8E4zlad7Y9
LMkW1+iDo8ijSJHUBlRMj67f9gyW5NS/W1Plp5k6GBGCFhKV6/Gj277GuYFJMNKhqrY3XgwzcEhr
7HkEg12ZrxVKMYadnfUuvskrLkeDDDyGBey5yJdsYiDMcfGzYwK6YL6zwm5aWN0K3HUKnQGXwcjp
mha+3/ljaWLYBRzrEsBBdJS55qkzSTbUkJHOj3eKMHyzfCO33WSh4Th52WSbd5hzuQwjSUVQeUG2
h+BfIdYWQGqkQZWHRVretSgNjSrs4/H/QxgJUtYgsJZdUmZn2r6JJmEdisZN2hh/zTExZ5E99yra
pyhEDwxM/dpyXKgTpJf3qrjEju1zZ0boZmLZO61j01XkXkeJel9Snkor8HHlqbzPZBdNKczTDJxV
BFbiX0Epw1HnNZxzg5q/ui0lWFKzV8CdqyyOziqLzZMnCdFWSBiK7wRBuCiywwD9lzEW2TYXhV5r
eOeIbMl+C2EMIopa1rRuSbUv6l9VmhFZMm5DjPZZz4cf9K/xRbqKC7APUvW3bVIAB7Z/iotaShDk
ogVjJpT+ry0/Z2ojAPrX7sBzHs6r15YSZcBKvtBlucFrZjTTw0Yii1XhAmt7dgBsgH6tcDRe/roN
r4kJux6obLlu4CgE0Wa0NGBtDbG/jskMH1OtNHFokLuphzIP/P5pvKZv2s/aF575IPbschmvq/Dr
tVJ56N0uSvYvIi5sRbsOHb5+mv6nuKVpYjU97T1nlW4pmTgReWXYMQQtzXIWoF2aVc+dn8i4H/SN
wfjwHYF7ucH6zn3nurjkow9EMeha3w4Gaq78+7qjCVi+KCx97H5b327AetbS0mvzXmZWm6Uf6Vm6
ZWE8F9fqLG8earqbnd1fvrZV2NEuI8ZD6N1NUvW2dYOif1ZSqbcuXD+36Dxp8s/Dp8QXkw75UYgL
wN1jTYnDZ1vkCp2BvnVqjMDPEyRFPs364wjK3CVWcI1msQYxGE9k/UveYlj22nf4iQfft4Y8+qio
SD37sXrc9XM5vYQ3YXpk7ICFHlTSadhF0Savm7Dg/Qyi1fwxjXaaD7zWL4GirFCZyMDBazdNEziB
0vFx1S9ssfUC/K3tTlTU6lNSafooYdB42zgNVBoFIR4g69eiKpVu9jdb5zs8zThtt0qd2rMPv98U
AYpiIMmMhFFXTwFk3HAgRTfjGWOulozlZNEp4yeJWM4EUktSMUrNgYqLqHkV6xLASdI+3/fXGG2b
qElXnnfdz6W0OLiiHHHOIZOGmJS1t76XQlrm5Ljh9ZbnDS9ueixYDKjG/evdm4EMxWODn2imDqDi
Ryqi8NRjAY/s7ZRJGn+owM1kBQVVn3gnAP4lu/CrWLyJX/4eXZq2pmz9ecii4eupkDshlkzagG6S
6ttGIc9x2KZUzrIhnlTRsqfGhoYS5bcQN57qDu7MSVXUW1gXWM+yjevZvIWKLtMda/FeQfzL/tEW
BDPZ1dnTIsaiiwUd2HzNssM4/if2iROAM/dpegWq8af3qaOYfr04MC0VIYGcYvFlg3LNbLBH08Vv
BvbDOKjXMSd5i6xXBup1s9YFds3hNsn55oow9I5pdHZXYQ7fx5LtmsGuMIfy53Ch+8z7idYqoeSE
oGZnbpvBkTxCfqTwiCCPfgmUXYJmzu8vUHAWmRMKUBWI1YvqtNWwr2BqIBpP3lsgHge92XuJ7J1o
0o2i0zdNyxIEubjOe6h2AkeG9u8m/8waP3zXf1rLWPFJyI6Ru9Vg4WGhh1vthivgtBYfhKzoev54
5KBYA6ZhPnS1fgpz2KiAY/Ay/ZTe5mEpld6QyfKvNGu0LuVh8WPceYntgB1+kfdLtS7VB/E8sJ++
QTqomGeS3OHk29UvbfWnCwMpFLxER57WeCXLk1J/wTYw0+liLKcRSkuRznskTAkD+1qLwX8t8qZz
mHCJ7giOOp9SjOhzQWpN0Mb3Km5oR5+FTF5KuHECMdWOu6BwqTz0WCY8Y+o74IbZDBEKvzP3f7lE
i/Z9quipvat79n7WE3UiqknnGCWfiLWwMVlUAcTUrRmnob8DEkZp2rP74OqrtEslaEtKMSbmGWzj
rTXKcZnxc5E8OBj3v7bCOyG+zxbpgclc/dAXj2qibjn15a10uXC2vofK6u/ohjnezz3UFCvr/Nrf
dOnf8uidfqFv8xPJ8Q8jRlI6KxQSeoV7MgHWXEs7eJ5aQE/ZYHM847//0epsYoZVoO0Jttcwna1E
nvTA+hj8jBt0GL2n8Hsg5pnn5MOToRklkfQ0dTcqnRiIb9XAWR6EjDCuT4AeOF3X3+MqQ+o1cnHg
Dg1CCgpqdvn+HGiLTUn+WZ3rmT0ZI4X7KRhc1pdQTJmHAfFTNTapJdqlZM7vnTrYBocbLt8cdzj5
LQgG6T/6njwQQZS5IGxmocDiOiwna6nXnkQ9pXl3TboFQ04kYgSYC7yTb5I9Jsl2TAa9zPGHOrh0
xeSS5O6BQsmxXwxRy1i4d9duaQcM2wghxY8hHNqFJvbiIgbMUbygdiweYV2HVQyl5EmJ+FzhFi9A
Kw39QS/yF9AMZdfphIPyYTD37QS0p4IawJoArs47iAGHjYKxhlib2RqIVf4OKTkYYmXoKPXULS9D
Qi/fEg24Vx09/SJrxyQGDmsId/cwsIhY8HTjDPKy7SbKqPDDGx0qMFDlTK9dpmpU7XXXv5FSCWI2
0UWWHIYKitWI9h5L4n1pmWjaUgAraxMiDP3f8IX7PiLr8rzX250Bwhv4gcljRhZY4vOVyt/vZrXi
ZdUYHeI1T3DvSrULi+bWEYqOXvezeAN8XEKfLK43VSP6LAqqFYABufig+PpGPVfgraVOT1vQcN3I
1wnQrjBrIWeM0CQ1eeEXSJPsr7eFK/6vT3eI2frRS3Rtt05p6goWAh1rg3KvwerDsVlXKk62iGW3
sz30ehrJVWjfJnFRrV3I6seBaP8bJ9w7kCG0DG92XIqZpbOfNQkDzd7QYH4Bs0+IqaqBapt1mX6l
fl0FZ6/vZV9vbU3Tr/Xp4mknks2gyZhWeJNvbIclaO4zJfnc0AEgNeBC4x1vs+Zf34UzSLdVHFAS
U3NT9pK6koUE2HAkk29Qm/LdQgQ4GHCnYGf/aNEFK1haFxlmpMkar5H0do7WkObyeswjBB56JHme
vXKxT1s8+Om99waRKj78g6xVLksOKi04lrcj7N0BMmodVuM1r3HQ+TzDn4d8FT4W3pC+w1b7JGBa
qusjwkTV1w0YF/xh3zAP1I1t0fswO6rjapeXuXejPQOHnvg8k0scbDb/xRvcSVH/YEq+hbXrtLOD
sh8q7B95AjTaDXRdGli2m8jG3pIH+tcuet5XSG4BUSD240KjZVzWBS/lZ4/tiU8bLbAZ7UNSdXM8
SNOvQ6gpttyfRnnPRqN/vRzSiumaIDljKtzdKH8HHwBAYVONS9FPi7HSbH5r+73JV0oH6/cK4z1g
ym1XU1jU+WQckgU+yLgYiuHcD7eSCTh22a8O70/5LUIpv0iDfmIvOMHx6JXZRCwMeReyO50+5N1u
Mee//xE7Te5TR+ijJVYUjc7HWHT/WAQaChInZ7CM7QJAiehf0baMNw/uPMSDFnBP5qT3TDEWZIe6
4KlOB2VKdTQTRkBTms7MmAfVS8CYydGCXuSzfXc/0w8Ph/9ViCduAvm0de1fpHY1vfBjXApaZr7i
dwc/yYReM+/noTg7ww3UBANDsdpvTrM9l3UWHF9n40ICJmHoaNKVWVut6nj08XwANEjYQpiBTZ4t
C76MR3W/tefq+Sy6v5NGt0TlVd5l7cmf+ZDl82Gb0+4w8QWxQW9aYpZ2O9I07lr7DKIKDpy3hMbq
xozkbwT0YPGC1EwQGBVt7GJE3611xnfUAsMWCQ1D6QAUNzt+RzxvPXb7uHnmbI7ddo9Z1T3YCU7/
J0goKxWVB5NpT68XGg8pggqqr2pyXyWdCDEnUwYAUnAs+pAcl5CmIO2B5uGPukZb62TzM7pBN+rS
L1UZERFVwfgTJlKyF9ewhSbCa8XKWiiyjTkuKgCksOdBa6XwC4C3sH1wHQssUBDFd1FleZxcws4L
IV1d371EXgpOcJgnDB4Ej+F20mMCCLOX9wqkQdptZQ1kK1bM7zB5x8XdIVRHTDiCI4WUhR8wdPJ1
qH1tbCtD+sxyVDPgLodZsOz4HAmLu3xIjV7ZDre0j80y4OJOQTBJ1a2SCdHbxpYQnNV/psqoyJSC
ewCjzZuy7Ug67AWJBq3iRA/bMcdavTehJiOCs1I9qb8QnmFV36XNBVQpeHj0Yyy5u1S0f9wI8S6U
q09nLavKZRZNWJEl3ES3ZfNHc82xXXTB2FJOv0/EUxwElZFoSY7cVXH9QIj/dOJGAXiphHQqvHa8
vz+4qPY3QMm21cMiC8D+0zTRkU2cnSazwY7E+VkOBVnjih2NDeEt1gmasFcVA68PEffIbMpvjO45
YjYkB7dqz/KvCaWvXw4jlHEjwcRmI38qSmG04qzznwCo2YYMa+4pM+indjj0Sr98+OYDEFW7PP9p
oXq/xHHeBsjh14DING+DMTsK1dz0aJvGc0eq/LCZ03LjlDycUaQqr6GIjaOIN0t+lLpsr7Jd8RSo
+GvQPiHfWfv8dUfCagHglIZd1WGgsSjzoyJJmj5SCXcfivRT4mpcW8uJe6cXxIGf6CjfjvRl0DYZ
spDMiqsn2APXK8XT6shRQ8Cnb951VA6TwRqusB0lgGUTB4inn1ZZwQspym/S2F+EqjDi2UQ01LQC
OuvqKk4+U/0YCzg4N2GsT5E1fJBvi4ouhDqJVhWc/y/LnSnekbcIpDxloWrj8UNovPb+xibKI5nJ
udG0BGXnUeMW9eWu+oC/NKDuR5g2TGN/xY99+r+Yi0UGFM+AVPds7326bu8xb62JsC0LSwf2jNnJ
uzRGDy0ykk/o2ygSTdSmVHZDg9AoOBdZHTdmrB9fgbJlUHowqFVsAUdnTcJNZvfd4ie9gpyv6d9P
KTOnxwn4BLxIqFgvuIBCAN0hczGt51RoajlxA17Oetqihbg9sOj9gRJJpnUTK3cYvFNP8dNTsHAX
sMHHnvu98JSJguHWc1UpsvVdlzDJ1uZ9LJ/jU/hCAgxmLVp2MwrnNtdaCtdsQ5NEQ9fuK5OKjoZY
7KPVNrt1ZAsY94AiTs95jT6Y0ihSFaWKyNtGoaFCI0y0kR6Z3mDVtpPLxWkkE02mOjArTGZ8IcOl
ACKJQycSp9nil0zNX3xITW6ZzIFLmbvAG7gVYoZ4TCuHshkuTHwCf1ALZBMv2KjE6r1oYOJMw72d
Tb/wsLen5zJ19WjE4NU8P5sNXZVAd0Ly4JPnP1NyOTcD4VK7hmTrSyJ1Ayt+GVKmAnJyjo2L0oUB
Iz+tqB2121zp9CGESthSY3Ya6DvA6GpnCN0z7RxF41zHrkUO3fHEcL+Ch2WlC/op3kMHn00RVY0u
ZEiYlwG/C5wKVmttp5WFYN2SI5/IabOi/O7MQOZ7zrDiBJVp5eZGWXe2gT/yQRcXvYt+6F4aNQLt
/stud6u/W/0rjADY6Z8ne6PnaaXL7eWt39t60y8U41Dy+qCcssKnv/7Uda0QhdJmlOZW5T5FJ1M+
DquZ5oBnDEPZzfXxaq6X10ZzHAGiwGUJtly94xLZgZ+v0s8acIgb+DCtFlgnpmqI/nfxPk7NOmpd
NqDznSlWSHaqwE6JE2uZRSWl0/zGgFbPXrKA/X73E05qABWmPwfg51yfmUvPA+RxD37xhjpdRz+m
BLrd3rbxx2DgJncgYiAZsXPRZL73r0huRKoeZwTpp6Em7EUYTcJBZhzUUKpX9fckSwlvr7lr3kLO
9YV2sBP8uyFXNVVod3DLy7F+IexL4hjI9kLYH1/qXUQcg0hCsESbyz1uDV5vDEbQPhObaycm8Q11
1EFpN1j80YpfX1lvgBaP0uLYRqVV6g08Vin534y0xgRlcKEcb16DVcGTDC3thqLBmHAqNynCV0kX
sBCriTeN3HorLWfYyVRcOgsLI/zlAr4XqHfiGJBYeB8jDVdYsJAtWHnJcHaSW3xDL9zRunQuQJVo
EGdbq/0lsg21T3yCc6n6nRky+o5NtNONhqymoWf7wkWs6dNOjOM+z8nwLc8+/kq6V6S6y7QmO875
i0WHTHl+YcH1rH0RiM8O8U6PoUrfTdgj6gU6LOM3nPLC6AysJ3LBGsAnonemAAyQygWfkjByttxd
zHvK2eCllmyKro24IH26FMIw0IRnNiZ5zv/f7loH5g6c+CBYwbPMgkHqVNBEnzHN3O2dSFnHmZow
KNi2AvdIotfsQQWlwGyDYl2xvAHFCW0WkjfQW4fscEtveI7BROGwgaDSpkI6uWgU6YSIYGlNLCh9
7sJtgqjDJHcUC4WHPuokTQAZF5/VUhf3TVXBUtFuQuebmREi+ZQf1As9JypVsDa3uxkqhxN0PoQ/
oGCfMh83xyTex4PTR3RHykEumeiMT33D+rQvGyBz49rmzKapUeEGFpZy1kfJiUhpojtKDFtKCnuO
OaBeB11rHer1BygpH66Qt7T33Z+KeKB9nTwPu7VWCtjqKk3yQv+WzlJkWw+fqT2QUB+FwLnNhgqY
H4vP7x5ZXyfMrSbrQPo9XcbFUizm2qi3LZps24Z8cMGnirPnpySMG707nrOTdZcD/L9YPI/n0TZa
vzs2xsY1LLHEL2dK6AgSqLm/s9l5i3Bk0O80vHogw7N5Vm89fv1TYr8Hde5MUjHqujUdfN5Nfr0u
BBsmNMfvwV5oDX+SeqqWumVuvUWTg9J2kvjy+W1SmjynSHyQos/Cm5q4+91OcFcyT4xia3zmqUwh
9NrKhB/7hbRjUPUaVFHlkwNMtQ4NOZZts3R71HUTb5YiSor2eRA1+7gbaZ+PGmZ9lVUeUl2NdqqU
7cKnbQ+YOUMrihV+R1yz+0mi91k20XpuI23FFJyCZ8A9N4mYJ7DzAmCT3VEWO+KmEEHJWAJp+hX7
SHHwAsoms9IR3ZoQVGVPOTcYz6c7E09DCO50TCDWb2xby8gEJaakUL9EWPwjBqhAjOxTOIAmrtAa
zzx7OVWKwDW9a9K+kTxV7/E36yfUMyL+mVp1ZX1U7zc6u1jS+M1zvGjfvm1lWFmNkdkDmG+godY5
n502+Vn7c29LkAWsfxppqbV+d7+jJZNBwbK6izSVWaKvpmuEQvET6rWVSGxrh/0GGb5w2HaBSKaf
3osAEbUM1GN9/1kis5OQnniCQp8S5J3Rutg2xj8VoAcVjrMgwIp+IGyx1fdmjeNmAKmqs4TLGXhy
3iwgyx3LPUzpznzf+yarH7L9l/GgPIh/mWOOGRdLXCVfvYykcak/qMtOb1Bm43efDURX3RY2bre7
40vJ2Gn4jpFVD84Eh/JKA8nBtUnfSrvgx8pkqvh52ze8rOKXO31R6M8Jkj8LXTBq41LWbjRoYIj9
IURYrCx1PQjLlhm+3+7/tc9DjN8E8F4KOHpep0sE3dqyUVZxfy5PV21EBJC0vCJqxcmgqdxTBPnx
tCNjW2yfRYf0cYGrHzt9AaID34G+M8OJt4VN2yioMUkEmURHKCFg73aE2EVk0nqghGpXZyotomfr
O8jGX/3sv42UXvPk4L51o66OsZ/z7wQaRyALqDA/UPJ7iMA8xwK8lTECWiVD2qEoTjPuIXqzjcYW
UQZxFMHCicODDexU46/7G0RiltJdZOcpWVjjMGlQtk3Z0vAT8uvVBvvEhaQxi7LD9o+nrWQIBFX4
6sBXvv8FVFkZGRLW9PUqPjUXLE8cCWBnED327M9RbeLslkQk0XJGf1o8e3KhVWstz3edr98fMFyw
bFHFoF8o/V3fEHBqk/hAbdSG0tEtF61V4lBcMJ3nNhGkifSRexNOuEaf/4SvZb960CZSls7rU4Vf
z2f1//5AvqF1a9AAc0y5UNUu3aCyrEUvEOLwlMu+74GJ7np2QQLHqDFD3PwqUUr2HofLWwUw1qpl
hWWfRwkEOA9NfDLSJcT+rxlJ01nzpVr4Gv5wzcTZEeTiV5yk/a/ZeWGjNj0P6XasoYtgd1sH9PdC
umjPD+/DtONJMOMnMlVCQeWi43oz/jIAHCSZaQRgxC86g3FqA6a4H3mW+K5wYIR4qZsQeRN5cNk2
GmkZxavv+9b7OyRJLTSV7u98RPnKEoZ1G7XdVmw/6Ixt3WhzCCDbQzNhgdxTb8MCRACfNO+kO+xX
akb8vXg/8+9/vOeAN1Krc/OMMD+JoxBUIf7qYu4utqpgF9moqPiSEwnxvTBI7kvAmEZ81Luy9Ue/
PPdnU7RV3m+cvuJNY3DErXz/k84cSKePuFu4cvFMmVNyiSRFvEClCqZjzmBwcVKIQHweTjtcSNN8
7tm0tZYEA/Tdk+cseXeQQInb54SApPziSuDkSlBlLUWQBCKHQw0dYUc+hTxWtji3IqQTHlvlJnIN
0L69pgCNRyyldcu6Nc+vdSLkF3YWbSSzsMI4IEkQHuKAP0jtUgjL+i1ylC/FiA4x2c2OrZdvjGtp
M8wqjwnCzDLvT/QV1Nqedzeli1lTw3so/926ey47YZJ2PYjKhKx/NDTuGk6DIf+KuM/P8A4qGSwm
bNyLaYhvxYPeffvVhHrEkwodeI9tP5isbMmISl2LeCHD5rxb5F7etmxVdY0P+wIKHEPjY9hp+73H
rbg2rxba1969KL1GAS9bVNo4WwEJ3cUPBAhCZI/V7lSzdcodW/wJ+U3MPeDT/ZhzWO7ZQJHDN+uu
VpQlUryTBf5wHkzUSCPYxa6at1UQeAd75/ijD23CW1aZtK6RZZY3zDLlK7M1dyq9mDWK1u6cFGJl
3iHyqyhYJkjoirSmBfh2oqZzumPKvsbvqJTQ/+85RgewRNGzjM1UrMKLE5n5BGsmhMFUj8plOX9V
kS/Xk+A4+KGu4ypAoVoPdoW3fHrmwm2FTOdl72BOse45h04NGGh5bn0ZfnMUHYte7nggIRBcAj1J
49cPTinYnHzXMLqPEX2wOo6PDiA2M1KdyI54QA3nL/nHjUJT5iRboD2p46vmgicBuzecqEqjY1db
MYKRitJpgMuSKp94pQw8LtSDfxXR5GCJBz2weFbWuf5RLz9L/XGq5BsZq5f+I88OHdQuDatLgI65
Y4Zyj/+LuYUsgQzKjx4lby0s/tWG5L0XLyBGrps1UZ9kmn0Vv0v9RnDg0f+p4p0TP+lfRAnEConu
1cq6P5E0lNLjHQ5NhbrqGoM+uY6DRKpapjE1jYmnezDhAq/VuPoPFy2ZQywuSSjoeySBZYtsKYat
BL9tzhj6YAUm/LgvzeMlK5KcRpDytX1468MPCXuEbfblXgEML2+3gQ5zFBYxsUD98Q3ervNFyIYk
7obk/ovoGJWIiXVLytdClk/zd6q8cC2M5iskfxZWuY6Bqe3SO9dv6mv7jygs+c0gMSe3IxGBG84D
aoQ/RE5RYKAAwPAEshFWWqlukh6tGphwPSzzT4sQGtQjRWzL5FQkgimIstr6Ny+okS7NARIIr/H7
81C6VmcCIzk0hlQYMJKBP2K1il3xCBZLv8DoloQ5nxEQtdeGjUkeutnAr4fHq6pLOoK4AK4lq732
J/9pAR3lLAvJ9xjavlJb/08AFNJ0Yyhg+RoVFMxLFbk4lA9jLnkt10i6dCFXHwG2xDSAtW/XG0SQ
rWSrDRm0geSw2+kH2jDWNRHWF8j/IUJ/9ugzVMKOeMD4pjcNhX7wJ3ouOhgzUdgOZxsAWObvVSPA
KbX9h060VVphC+rgz7tve8JAffvc+c0g9AEC6Szi1x1wDw8XJx369d7v/ILWIWpBFRhKVwgoZzdW
x7WJSkfhwtdhNdEJV/EZ/ZDpej26bknwxZKVIlvE2a0+NAzrIC1TKHTrmGJ87yvTlN7mgVc2/jS5
yrIUAvAHLwW6mcd2EwKrYjqEyVeYRZqYuR6LD9YGBtMFHpxkWBKJLfE0TX09lBh5cZTgTsfSGeDo
otgSgxFQAoeQgmQ402Tk5j41LXcLfJy2mCNxzvj49fPdreHRmZ5nSK/M4dO5Zeo7XrsyYML0jdM7
V9fd81EZ4WzcPY5O10Q3CvGS8FarWYwl30D353Dx/PkpXgDqFYMCO3haQ0KInz12WKP5ObWS82wT
bJjn1yINofBOdVMCHfLaNmxkWPKMCuvSk9j4yoWCx0GgAm0pxy/Fse0V+rYLr/EdmVjV3Hc5Lf5w
4XukaeR9FVp2u1U5QW4vxvXDm+mmkBCfzSbwtU3IHiKdXfDrkapYxyjcLWrYYSARN6P5xaZs1s6c
aCjbuUsogBrXFUrSSoUhBd/CaV3RLNGAHJtn04nxtusgLamreXTuoZr1C/pGHbtFmwFbHUOl5wel
f7Uo+fo9Lj0OIzq3t/1L7tjaZtxKhEqsBatvr23r+bY3INeHSZHk1oPdKmw5l2tw5L+vpJnHVEln
tSiB/rII/TcpzOE7Ib7by33l3QFgnYQDnipJPrit4UaGr/8kOiP8Z0thB5AnJ0FqT6tXrhnUraFz
Acxnz78efEUeg1D1aDLReVhGAvLen4XKzo9sp/IInd3GF/RZ56qijUEtMJEHnavNWzXUj6ybsYp0
S4gwQvJXmkgrwgRPWAIPsBiYywrQq3IaDH0L4qcUFkFnz8h2v7jk+n/US+Og0FSMbTULa56GK82a
CFbX2g64dVMaOj2Qd70kD6TCBSvC69Q5t+4yu0VRx+jIUXagb3iqet3UtTAUozas2NFoM8EULxO8
9m0KeGxDl4WuBTCQ0APSbt6kwjCSX/X3RtE57ovWILt7O277/kM36t6jzVw+h5xlt8HOE8KnJlcG
CuADrPUMkq5D1KhtSZHakz/cvW+mIy9YKbzhwmeaMIUXA1Xdvzp2V+WynEGdiUQUxN3VCd8hgFML
TyO6RJUiz4fjbp/A/1tyxPKmdOcmhAiaXPDJ9X1K00UTiyNPGDR8u5KtjhmY/bUy+VgEiKwW0zdq
GwU7rkqEJMks1RHJUd0VeOO8GeXgbGKQxFzqf+TydbdTQA4YhLd0nXb4F3BdfZbEW4XfOucCoynY
ZkyCrELKgf+iwcDjEo+nTbByT6lhY+6OxZS0l7adWHppEmcKHxVCN1ZNrVikwxLmMV4JMCjDc/8H
PNQdvobXmTwNJdSsYN8/HeaxtYylnlujjt2TEwWnb4MXxUtRmqOPUhdn6lLh0LABndQpqyue7NRH
MVnMyxK43fBDjqRqAszSwKnS2TOTqxFXIbo99rrY0z+EDdLJmN9l2IT2jM0zYcJ21TWVNwb5dAeh
EQHQ+AJWyZcIDoD4n2nCx6IFy4LjqvLuYoMh6RmYBO2TfZ13ICA4lo2udWY71/+h837rleXIHAU5
l6Ykkq6vDlxr/66ylhlQZlM4n/NIypR33XakBnRXrjr+Bgwt8luodATmXA8SL5TnWHOOBpLyGyt3
RmI0nW56zGY8gRNCjfAiQbyV1Dkm1svGUOdUv/000gEc85/jo7RnRBCSJbwIbIJg7/B8LuctPJlf
Ad6Q73shtXjUxLX7JPcwrwNLHHAImxeW6GHkYc25ijcBRhX5g4ynKS6VLcq1wub4CrnftFLO8n6y
hQql/aKFqNYvRkWrtLnEZIFydkLez3iuTtzAomTVC7MPsUeAvEI6uMZEqm7zFkTAyeJGxVreF/KK
Kj7v9XYKtPTN1Q1POsKggR3YiFB9+87Zdd6TGp80LrKk8vu3D9wC2nk/ILXEMSnfAeIE+qsIFekA
HtDi7uajk6LI1jwMqkEhO9UsCtkRAJYhQwukyFVKzb8uOFete8V1TfJU0TcDM7/gVwlPpQ1kM9rT
pvrYWrmTsHFNLJ4otJ3DCjdEBgoHDDKL4LKD/DtKQP4WOT5iHHmCFn+jq1KWBq+fazobwKftpfCE
/BVATxOt7XoZ/qaQlro+XWgDtCtrxQdSQxr5d+yd+xmWaYUOcPbm+pIIA3co6/c3k+YyLIxC7QVV
C+GOY0ba9X1UMXnErBjtKI3CuuY22U9eBnHL2EiuSXzsqbTrNTS2w2jRKvt5yJvIalJAhChY9Skh
Cm2PEh1y7JD5dcb6S6xb2Hz11oQxpjzwsOqxAvp1o+IpF1mfe1GR7QlLJkIzIbU3qd3YmSYPPYsI
hXNgnegdhqBl2VrrY9AXhp/+k6qAr4x7Oc/ABNrlV+2T+aUgWvX5vfNULsbf+6efiN9GYOXScjkf
qqNNBb8k3yozUHGCW9wXc07erntKNCqv3zl+ktb6OKQEZvCZFCZ9GTW29dJlOgDGV2L2Y6AW3HsG
sls2287A8FIf8nAXnxv2WyMOTH54tItjgRKi0R4xbhoPorClpcqHr00gpEpEdXNq7OnzplxdUPpk
DT+P/BCuVy21yZk03BUO0Zn+Qjf1XqHbjZYO5Yez4F8xavGXD0BbrRYRNuI3GHWyHLrUzg8Qokrp
NVKDlxeeLuAD5xWbImmqEMDLeZa18ASFIga0DjclDrnbSQA0ZfSc+m7zYmDR6ge4UHtLMupppW5/
jr16CAoKugXXx0Q8l1Opn5Lb7+WmqHGTOHVK3UnCFWbC2J4vxy3eDNlOVIt37f9hEVII/XXzyfEV
l1CRlDGzXOzLr063LjmyeVtcKTnO1BxhI0crxggVcEQXdNsbuTWdo5vfznJsgnMD9AGCKopqsFil
FJ4V2O+PIBCL88jq47vSn7AC4GlNtoSpece/vHM6KKikzql+U1q2ZGQ1CUjBVNnDzzklgsqVXc5Q
6pDw98nGnGDUf+PpZttfTmWQ8S25SuOfw+acDI6Pr5MbSAPy00v8gfIHHwztdWCSAS8IP/tRQH3w
rkBE+vq1wm2OD5tZKUAkxkqZTZZ42uZVCb0GqqwgwhczRy9NOahPL+vKx+5i7gvnH+vrAJGe9AnO
cmwWz4SCVtU1v4TMJ1G1eScku/PsBvTxFGrc1jkJGNjgb30BwWrU7t6G0fqEZJZQgZuYZGOU0OmD
gPkSFeB5Pg44G8wE8eSTxobf4q8dFjOIu4/AaKMCSKpZv2cCuDehnxR491SJMaRRYeG9Whfesaw8
/NTzHLO5YnC+dPB14fCTaNXG9AL0bdchujW1ab8I6PHT4qad5Ufh7VrEcQON5BOf62X23E1HoCiO
HaYQKzjknHKZKaIyOIewmUDGUZNlvPiRW/69wnP56haz3etBDYPZnU1NLDGDag/L0sIzgqgRFE8G
p32F9sZhySd/4xDn2ZIhSKb0g0wS8uiGh74chlbpuUBPfuhDpNqSQXReeSSti4/cXpdXeCM0MD7W
HgiSAK1cs6eg59o4S7fsISIh+rQAWTQ2sAqGEQ0th4NNy0p75JaCVNQrVXqu6q+kdlRsbYcNVXej
ZXcq5PDli5IgV2E4AF94fViSQL/7rkAt7CNicDRFe7MX+pO77tyOSMVHPUPbIKP8HvSqkKbs5yl4
TYB/EMXblesD4iKsqRE2ZG/go+EooXumML1I2xEDPG8Q6WeFUvw68WdcMaSTu+fbCoc3bb6luOjz
vA+jXCiTVbHgFN66ZzOUfJ5L7V0cfPBm0WWdGcFZ5e+L7siJ/Kd+2nMlZYHmO1AoV/Dv6qs8u6EA
NclYZyRHMf5DABim9xDBTXdt4TLNQSKM/RdSiThNhGkrSOLNU2/hp2JlLTlukSMRufwN1oE5FcWR
P/zd3rrICAGMV8266iOErLmkjpYACY8/6KYMueZ1fX0ODlKoKumuch3lnGZbuwroo0ZMAORIP2uF
eeceK1SwL3hOLI+Gr+t1eBJb+CAx/SeDFNdvCW4diAprxr4vo3tU3XB+6IToZ++K7lwQ/QTDIIqW
Y6h6GDsVNUcjuLqY/1QbpUuyJ+IEcCQvaKu4pHLEjZxdIzCiBAMk0B7un8oivHwhZT5GZaodA65j
K/WSn525i8wHqrL4aIpIjN/tI4rlu93wjKZddo88B1+QlA+WTJ8WEE1mmPLYKopBnwb89xGSLhXp
rTvvyh/Z8Ms1bLqqQqKGAk5ba5Q3DvB+2i4j1490/o2DSbnF2DcTBT04PjbUvMhRYw4c2m0s5V+p
lnw7RyAVjT3VqwCvpst+fn1k3paLtOHbt2AVr6KgbilqagPOJb7vbhUUcVpWF8t8wMG4qoGJywsH
WGeb8RnftFXev36BcrEJ7Dgfk4kOFHnPEOo0M/CTlRRo7j9QamO446VQcFtLmaHyzA3w8gyh80Sv
ankAy7lSPa9QQZ2eP1nJd5JVbYTvNE7XQgEKSPER/X+t81QCePpsFhGqzuUJ26gffIvoRfNfxLiG
QYus7oUolp8kU2Njj0GxmnJ8wg7fMO9pvXhJi8lB+StOfqkWHPyb6mVY2iy3/b//PmmrSXaZBGCR
mFDdfe1hExVEVKEYgFgGoBX6uV5ifVDsluh9eQykcqp05rJpKDN8cmlhFWbBPDHYlTofxs7/8XB8
1209oGLStYoSSieuRnZeewPMISvyn5UOmhEx8ZqlTEISaPAzYWWv3TBKF3TSTJ9IXtrm43hUq8Gl
5xdcYKymGvAt6ymPgIzs4nh39t0vIerlRzYpEejwyQEaHS7GBR4I2Ul1PDEgEtTPgMfFP1L+GZW7
wEMzoottUCTAHnOf26Z52aciqxjbBXcfuGiV5Ejq1X22heOtgU0d3D5fvFVvR78b3Ha4DauOMC2V
b3wpYvaRDOeb4Cx37e2ToHUs7gijfbSTDCZg0NnVAtRYU0ge0ldcPaXVs2dYN2jApdg5fLXx9Dfv
a+tyns0HyfrziBBBxpSwFRS7/GbjALiwUOmm/LJnfH4W4VCaujberowN57m3SxF+2gpYyI+iW1jI
zZZQOZ12ddbGVfM0ZZFtst2OZEJKSvjOjBaMKHE8TER4S7RCQRBInkDUVl3bCCaqMfrCor3iSRRe
4+mP4cH7H+vITaK71kfOWKMew6bbhw41fpmAghJLRVm6gVM+TqorNArviqdCUUElgwj+nByHiw/5
uY+JJGb7D8ZtWcTnKcyll0SrRaoroNbR6IPotNTgqmcWOW8G3WrFLFdmel/iEj4E2EFsVogK2rc8
ILPf4xaXKdIU+Nf9V4mMmqcYj+uJMbnUYP7xmHZj79nGR8O2CCUTZgRUR30FH99U6uQ4wPmlRJbs
b1FbcxzKaajmy5OfUq9ow7ZCNyMOFAHlCqvJ6C14d8bf1tQJhK/eYZYw8sl5MoxWPmwkQtwPtTT9
tR5n9Rr4CYPqPGgT95QVC76rsrgUZOj0ARZVPrtThgvyK174zi9W99fvD2gounzXK6EQnE9oBDha
KiWNsYLGTugRtAO0FHRWqeG9tFVLbhKwAze/PEJjhjmDMmoklqX2Y47Xm8IxXYX/Od2ukCu+K5bd
PyCp5VxGiouOnXHVdO4jnojQb12giUJBzfSF2Fo2/AKhVj3haBe91iKhMVzl8HXEWeZG3MUx06Px
dphWzG5/kSbo945tbbjhroL31/V9K9XXsOQoP2APBsiosmyYxQncVcmjRaC6SCmY0z4D+idJl5To
tUEeAqs60KmMxmoqWRGRqsO2JJg+QyPRrZbsNm2iNOVhPwcvXJzYeH/FK7FH9F+n3WJnKF4rvgew
AJWiYEvEopjnmz5Usgp8fjJwNasx/4K2JJeSyIT/I0PZsETJllyZPBqy3TMkIlhxEz8o+Tlj/Ngf
LWkX3wwR+QIeEfC94C+834oWRsRAtc/8PfEQUgOi2046rBqiemkZlTgfa/dfVqY6+dXa4bQLZ0Oj
YBa+nJLgMS+82HYeLTE28JIy9qSB5BjEjwp0tun3bn2XICcAWp/1Cp78+E0N4ZQcXp4pgZVVAaNG
LRa+kQl/94balDPXzn8b/3mYxKgSlI/VWmCslKRhi/3P1eI5o3C+MlxO3anQSbSC1EdTpepPdpFh
MHI8cpt4nvB8nJ2HKRwE4siINdTRmWpGQupI+w2FIrNW3rSY06ZZOACUVRlT1W+WsLXGFSlkYTtt
Cqp5Qv5uW2xIn++vZAg2As7cx6F5Npvy4/8vdc0jNatPl071PS//XUQNZRTh/83cl/geOHMGwlD0
Ng3/OJuh3kkBvTLC3kCyn921ZLPgJ/xYo9h/kDNUMoHUiHo7vcYhUJU5MHZsXo2NUzF6rAL48hf5
UP6JWq/fOO20ysOKHPDnpgHmTf4WijgLhT0lh01yJb+X/lQwCJfqkbOV9JjoVb5OZox7fm/hTNAx
enkKdoe3eYDUF3IdtHYsuh6HrRMj56udno43N00zWJ/iWi3JjV2G9UhWCAW/Bzcsac6oKJ6alOUZ
JB68ugvBY4HdJ8iMVbiEAfItbepxPhE41H4Jx6wPRPArbgXjmFzt4x8yRnINot+JbtALYLZq2LoK
bC2JBc0jsfJGIbuFA2pjK/ex2NIm9i0uKVvGZGuwKR1mwWxf22gFGCrDFyntHhvC2p7dHFR5wzfi
93W6o3WlvNYck2Nboo+p4RkluOwEhQLx63DjtRvw7uF6JKGNna26tDA5bN6o0yjKv81qZ+v565Hb
PPTMs17atm2U0gSRNLpyZWm4a1WljVKorbhQAKfsHT2PqycII66pKAfcAA34276BQ/uZLPqpdpCm
q/d1lFawUB2FxmXKyaaxLzSx29bV92xN5YoOPPlGhcDQRtK/mjIgVAbBFBzv2ALSBDJv0DywvLGv
LD7A91VRr9YhgdF0bpZ4niGN/oT4n9k3I2efhSWcfLMvYgTnBxBo/vJGGWLeQz/LNmB5H0s1UEAJ
RHTBaC/C1rt6h0qht1onfWvX9DvbwyRltJx2eUKxRrbUJdcyGWdni3sRrIUtw7MqM1u6QEpqIHSK
KPOuWSlSUcuDtHnxPoLKeCVLpIyoWSI3NSp9C16Cs/cQMxMlmJfNAuakO/BAYbyGgmFmTknVmUqh
5Lp6x2dkhtD2lcVG0GXgqn7ABDpmNbjEcyHkWdgHAEXWBRBJctQWuJp1N9qUCu3tfOdgTo7QtWBF
vDWqQrhnlwWvu77uHSlnXm6U0jOqbO/WfuQhW5rKrBHWk3IuykcK4wNHXknIZvEILMOrI9omjWfR
QI9DneJ6hOUinWmT3NW5CLlJEoDdVzzaNAcK3VWoulwJ2P9+Iw09PaK5XGwglaNUkgPclhwaqBmk
YLfmy2KX5BIZh8v8Fe4fa/LUmwyjrNVppk2Bd96HanDepNXGZWMn02z/vnqoTLe29FZhh1+ajOEG
1+OB6F39C5Et2LOa3xRxMExMMAvvGF0jwip9fp5ud5QjcyY5P/+PgFVWGZ/okgnnjCMNZAKSw3xh
8mIhc/PRZsyNfjzpM66iXwm6omcG76Qx0u62RrIiOT56byWDo0QQ0mfsXBTCibF1TA2TJldg0n5e
PkmvSABw0T9X8H8I4UhdYwLSsJo+PWkrN6hY+avDs1tBkgm3RZNeDqqYkD76QqP87FAhEr2xdc7T
6376KmrQqEhJZY4YZJ2GYUpqAI4KEmKlG59upeegMg11I2lsmjz7ggZB72PEGuh+SFaRIiEic6AX
GrQ0EyujUp1BZ4Tk6zaPw+DJXQyD+qBkeYRwFz2tZ3bEmSJgtKzaAFy71XHJO3RtvetkuCCf4vWv
XtiO250GIlh6gsywSzlPSZG3mlsrv02v2SEvUYZHOezrQh0PsdIVMUb2iyIv0U7awwvLVF3GRwHf
0x36TmN7DUD2w3APBkJnXLAkEkyILUG3+9jFlhwRH50VMNPEl8aqa9xBjVFSjVmeSlf8c6ySitwt
a8senq3MPZMH2B7pa0I8/uJSaIQId2ERASHMsHS8heOSk1dOMaFL1/tAHhDzVKWMFahaZfcjQMiZ
ho3vIAlf9nah6T9QXwdPrvEj8yxnxKbKKqj6ieGTcurWYEC7QaeO+zw2xS3eURhE1w3a1UVmCtK9
UaJhbg0I8RE1yflpW+lLNVzzxP1SXGNXNmOUpd9jHJEI0FVHtwBNP6lT8DdUP4xLTd1SOmZDSabr
nVmwBloyHl01diItgOYN35yWkTF55JkOSYT48k+oXDp1T8YTvyI0Q2RgBTcQjfm2F+OTYXHxdSJ3
hfe2exL5QFfP4myR2VruJ/LNYAw7YqW67SGh6ISFanIBGfagz05NQhGZznFdWxWPAP35lJqNcwu3
ePTcukpLXLAqTRa8sR+uFMK1+AKrdz1bw5ri+vP5DoSNdEyV0PjsW2N8d2CyUl8+tzRRy2wnra0N
ogRNLiGr94c73FcQ6GHCtmbdzOcwFF5r/haW/KY+moAGBoieNBcCzWihKB8LQnN7u1cXr7N2cIrP
oZiQeCPN/Ue2gYsN0j01OfoXli+d1Dh29I+IutX/tnV03OseT+HNv1JDF8jwXbbMXFOI8BVfO9uB
twWVk5Kt4eB3KKHoPN/KPN06tdB1BnRZcf0hBSwJqlRP352LpaGd0Oda0yeAyiUyWcc2sMhwebzq
LJN1qmUmsj3LjjDLv+oCLVB/vbzgCERXZn3fudwjqj2BpS3y49cSSwH+Uou1T8YEzdBusKN7xUbT
fULZgwSuQZmeqsAoMx0pXdlxq9K3p+9kNJj5bAvUFgDLoirYYzUULgWSBu88RN4sqzGR4VU8Ke4G
7aE8kNVg0gU6qsovNXNSngBdOGOucHW9MJg0UBOFZNJaQNJA9vTLVMEBhZikuO9M4FgizkyANSZJ
93eiMkMNUhVDzdM3sVCZWB58+ABupSi+MyysCppJth2IEfkct3f1QcZUvET+PQSMsBuHOTewwr9H
aEWi9LRDcRkxAGY6/c3EtfptSKxO0b/Eu3x86TGL/f+9dSu1ILTPnBddgUbhs+QE+FSQSVwkuDqI
6vMoEwJLjRCkexjyjBlqAoiYNlD7sOkwcc+xuy2JbmRuutoMozJY6ozcHmSInSaWOV3qM4C/+NEx
Y2VywzXHiBw0hT+WL+vW2RVwY8N73A0m5+RXT+E7mc0WTROPvqdW9VQ8dBH0MpI81IQLvzbdDy0i
ZOIDAJF6Gw2PvHqsMjBk8EIazwLug1ppRe327o5+D7F3lAWk//8Xc+cvOoSzZ+mKrENV5t2YKanV
nPQWASLVQpVCS070HWNzWMBpror4N5HTsgKHwaj3nBbQ56C8SV4fCwsuimUklD5UTQiF5E715hDf
ExQwsylPhE2jhGQMDkxkdo5VZxd9WOEOFBv4+ch/fjif9O/z4ASIkOj9SMBq+BnwUV0pLP79LZiI
cfOIWM4EXsJmZjZnJ8ywvzy6+WNW3i/VzcADgHbcdRfvGOPw758y0QwBLQiI2BRbUHSg2Fy/WW+B
wiUorFGTJgYpZgZmcqO7/kFCqfoy/3hkdwiqcBSZvSbxWGvevRrz/epB0cgx/sxM1LllFcCRWv0d
okj8GQ27qkNSAoO3EZlJevpffBl8whPZ6Bd1fto2ODQ7MlOeWkZimEKCaLtCcRvPFd9nsltyCFvM
PRjnd7zy/BqopN/i6ynMuRrVeVQNhyf39aiTyY+cCDNzsDT2An4dZ9UMH0FKCCtq/kGveXhUHwmv
9TSSyBJ23g4Oe3KCrRnQGlIAOy+9FDLvIPFx15wzwUA2Snc8SAbZyGPy8cxv3fn3xTLZ/a4Vgpdw
0hxpPhXlk0fPNfFVDyMcxs/ynVfNTK4wHTAIO1ReBaz46cCcFrfy5TTqZdBapwYX95yV3tdB6I+X
5GgzZfhb7UHeqZSg3LD6togXxA+tYCi75zB1b4t4QRbu7pFDoVdFYTfcXg3FNA6fndNz7xpGA/vI
qMyshM83C+o6QoxKw+7/ceh8j/BEN/1zar8NhWpe9WjazazRGpnqxYRWSxQTZw/8UPaQUroqyxw0
Cfh3nDtTc7h094FN939+gC/rQOxmUGDZj0+BMTSJ4XWqWwHWNXs3v0F9Yns/tPLXMHPUg5vN0Lfe
4TGa1JFYUhGYHUsmQ+/Cof8pcAKbVstsom7UpMHShec594axnLICT6qPDCg67GazZRYsoJcN3oz2
YBYbjrZpNY+vbLXODRmJfPoK6UnkKWrfXvLUbJc/yzMsdZegyXkLCWNMVvMyahGIlGjP2kiqROT2
YpfceiOFWsHFTwcnKW4SvWLUQmz2W3CvH8bntTB9r9ofRCp+XhydDWr9a6CKPjrI7yf7aOPb8EjG
KJzg2awvh/pcLUibkg7easHUeng62Kbe1QnlCX0X/i8w3vGI+y+okLhezEKIy88b4JrNT/0d00DW
mDS+bq9UcnjYT5CiYju+w740i5XUGmOVuj7vfEYdpciO1P8CJXuBpTq1IzfkuYZkRZnmf6LhfCFb
uk4nCjbnxythEq1kjCdY6+e7/r4LwcocVN7O04wyaBZLELGZ0EL1/Wmz8Xbva05eIIyMzJqJa3yc
smuVRcvY9nRDWc9ADikFWZ/aPRqo9fJW9pmoBDxI1Rk3Y/kUbcCrCuagvyFN5EZQkdL9a4nI0zar
wk0IMsZp5sl0ebvI4BKCeV1bZ22ILw0hqVU7HIrkXElKQ83li2tYTG/0MnrJaECrUVhbcPmGTWbl
YGTFLJjL2sPbdh6sRvFdm2SDLUcLcylO/zhVi9xplmsSrklgyLXDDygRqMMJN5CDPbn2p6oLKBJ9
+IYirkbh1+2sHKrmkq2b9yWuI/ea+0XacjEJiMysWdMZDzPdwrjBqMMpRe9dYLVMl3fcm+HeRtwg
S473Ys1hJruTE6FA1q4pYipBfYL2mp4S9VwNeJ3GXuxaapYLcay5KGCwr4nOLxmRpA8WFoFRZTP2
9NlfKEW4qz206/DgkeOVNCEMirXOBU4bRFpMklKFnIczx5cedl2AZoj+tZpqD77oreFlLh2hH3e6
l+R7PX4HcSF32tvWR5bRzMFIjlzhQwEiMM5ndhrKbvycRP1kDhcDUSUYeFRCovB/Z00QoCPRGxXB
x0T/cl3fzKSdKKSJ2V1Op8mWJ1RgDoucc3LL9Mzbhv0UPSJzG69oipzdlH/ibUm/5RAFDPWt0aeh
g0+/CDqiW7HSj4R86R9nTUWnoXNo0JrMbp/py6gnP2twCPwLn/DKjo7lDYb1lCScOxssS3FBOTRF
GkdC8UIs6s9irzd+hTqtqbP2TjCDVfujR8xQMIUpjyzta7prfzDYvql8CPC9YyunJKDN7kgVRKli
BNbgyPREuNXNGOeLhPdSXlrRXkQ//63S96fhJSEotAh+pJCfnOe/c2pgxvqtSF07wrp0FqMz8ZDb
OiKQSuAQFYFHrq9LjPRZYV2pT5VU4krbfrtrtkYWpQpF0hqIFFmq61e5wRWk3zUddvhiKT2WFAYv
YFxUJmFIQ4xVoplykO3sxSIzqVWsrem6QFwE6/D1v00t5IuvYeRx8KHB5P/k7bW1HdpPV90kBBFq
gmvgAwRx0dvr10b/WtLsQnRi+fhGhOe9/KGheqDKc/R+bJ7cvJwWQqnGWXN+XBr8zYZXnBpVIedY
rtO3ZKLaRzLC6ZtdfGNt0t58LAWqq0sGe0T1QsbjiDahLa6/56rsNyAMDaWxnv6VPPOMCWFqPn6Y
r8gdoGYAzcXquSbM/pwgIwbO2GTea/mjd7XowTwOG+34+Y4zhNb0l7OgV9zKDoHLOqRZc2K4qHXH
9kuwIUxfcb/fBIpCZpldbuvmtZ8wClxz+UwLpbn1qfg+QUr9FcUovq+xMawSBjDZU9XO2ZXghIOA
tLP0QPGdSVjS1ckkCcNaRf6ovf9b004mCDUjcDqa+CSr7LH/YKVniQSiOVPmj4JaG0trcjK1d0FT
9XUkjiGAr6cfuCH7qk/AkcmjkiCjAIGYP9RC8mmtwTgamNjyTEYOtG4EdAqR59WfF8eOkoI/3ScB
feQHjqIBqBa7Vk+2SDf6dlLXJPAbeN5HFIpR2IIHvLy5Qe9h70d16Y/gU/rnuOut6ZJzziZdcw/r
s7MfDBniPo6w4DAGVddMrTvPb58p1GuGe9zfm48120OHnw8WajTZUhlutZoXzPt29LrNJxuDcHXe
H2aAgaNhB5KhZTTQnCx93HIiH3qFpfZYEkZ8sF2OPpVIyomzBZm/sup31uEWukYI8IPbqRuK+wxw
XmaOiM+YVE+VeyqXBEoyQP4ZFRJkl6ONa8PCal4YOlN4EZ9GZiUy5DfgLVSkHpe81YdDwoQjskHK
dbn3iH+CUgOFa/BH3FCMv/yHKWcMZPvCDQT7nFtr68rMJkEEpjA/HunWniu8z5/8BIEFBxM+8Z+B
5ZPV4e2eNcSUTHzbcGTNADJ6rTlPJQVsg5MeZ4gmg0tg6SdisS1FS/c7so/6zdBkRDi0U9gACUzw
dWCnQQXrtIuK2yT9DcMGchXv3fTs9snKUal5fC/FDZyP9ttUCD/U5FQtdIXNkanuO2QLVF1g++K0
J+3vyCEYDipzJ1aaqaUzxbWeM/YtAB84OX0vQTggPCtV5l5qMcQYB/MlN1OsAcXN7XGdweLLYeJ/
UXoYv1aWM0ZR9jGyxPBNv2MLhqu1r3EkJSQX17Rk73ltOZjtVXLaL5Ws1cEGoj6al9igp4ZR8gbL
Y6IzyITBC3HEAezoKECS9IzmW1UDCriYJL3Ad1BFBatwB40NATfNnQueHrXDwIUJtZwnqhwmaV4h
paI4F75WZP0flIy+QRsSZVa8owwIfxwh/zfHVkOjC2nhwdNHH5hrgIfKG64gwG3oM9S1KmUxrk3q
5ND0RDgnSfomB4PZiJLb1vxI4IiCXEHZk2Dy6x2PWlivLCpUlILZVd1/mTNB13ebApNP9blXnaRa
w2F4yy4SSiyxtSpGL9mSvWRNh4BIuS75TXU0CdH2LLWXXYn1rj12aSUVSpExKsBpnqPkxGmcgKmF
bqX6GE0b2gdWNf+LfhiabElmkzCPvRSg5xe7Tym1ZJpeY47CQWD3cD1JNSja/MB5fd7yB/059gwL
HuleMb8SE+hVlN+zZhbnbQXd79hcaSyjsTPYdYfH/Hv69RZCxVgYyxkSibCbsbLFO5RFx2WUXcbk
sdannFnTcc69jKEh3wdAWbxKou2toHvlKCAOcArtg/cWJdOt5Khd47Kwb0iaGvSefXijtI7z7vEI
vyHwbF+e9BolAAHaK5/N0LAEPLvnbY2Lh0bInt+HU17Z/Ril1rih6C+W9HkGupKfXs+nz6ctrmuU
e0UUXOzpRD63BXuU+Z9Kx1uOLNKbsmG0+wO3OrtimhneETgAKfWynM21nsuRD/bgP68n72ItXPum
Fn3yZWIjz/F6MoyQ7LPCs1ED1Md3OKKfuhofQctkU78H1NfonymQdInNsDc8gXf33N1hWt8BH4YL
Lkboi/LPF8O8VXtsdxcJ/j1jmcd5wuf6I8t3piV6E7mt8rAI8hA/X9FWPnhoP6FgZfPzq1F6k8jH
GemKwAVT5oNiSuYRlsx56gd9EMrPq3hjA/F0fV3EQDb2gkCjD0DiZGIx82/htWp5+wyFNnds3fj2
o81KCqN+Cw4do/f/Qcj/At4Yy9e/DNf0aHBOiWhTjIyndUCIkZZAnowtngPbJNf2z40q4HiHZUD/
JKCoMo1hZtKlXayb+kqUV0opj+Uxn+nlFkVFueNhK/xf1n4wTiIfSGVG3q+9ThuSLKMoCAzguuam
H/xP0/4ZrKwfSKwdrYjSaNipk2k8MFJ40GNtkLQx/sSVZNl+oj744n4zjowjVd7cB+wKZ0sm+I2C
1ViZDxZWYiVIb0uTFKiKwzgmQWNe7/ECcetIkhgaFizKcegqDkq/nox4VxDhc/XqAPlAwAwlQB2p
gEtQAsqR8uzlcRak4vCfPXj4WRsD70rLfK/XgHVzlYP3DznUdllx2qVHj/V0StxQwLR4D2Vjn1Fo
dVzve3ZfCm1D+9N16Y2PZs6YJCfsW/hVZOM1qtooMNEI0kSqpJgGxnXrKEnkC/yvIZ+pofljEXQS
H1hXCAHdFbD3leJMr5t5nziQ5ZpX6KcL527KM83tvyCiDf/8mWrwrdAcOVjxueKieR/2Kl54Ccqt
yedxbG9XDEyMpC+sywImMkHatiWT9hVZtcTghBC78DSJv9yWVSXbOEqbpd/KFfSjbinIhvJmAIx1
ibQHf/EbEKw21teJ+PpBEiYE4EYmxeB9sFhRt191xSBWNHvD/x3fBxuWvJZbuX8pF18gKqoU9IO8
BvlpPaDFPhaC3+pivZ9mjNhZbZTK1azFnvzNh1obAkFYCn7qJedx6+/0lO/9CpFUSs+2nsShMaY0
JFDfJxZQewlGvhR1+//kTglUNJ1RIGEW6hRDL4F+6PaV+WqVGwYsNZQvhirlAk4JLrnyYC++h+eT
y6gGdrjnCk6NfgApItogPUV1xLiK4dwzNU2gfjYMZXsH+Ki6P9TwtvrPBm0WscPg37weSHA6VZYv
qeonqdtx6WltzJOkUY9DEOsQBrqZ/zZOvvF0R+tS3cQvnRNW2XWsWa1VPaoCHcxqmUWJQHTUgdDc
pVce9bFJb49t1qpDh7uf7MdVY0V/MwPOzt9ul5a9IZI68mVS1qMhvO5Cps6K/KCkd8l9AAtSTf5k
dT2iK/m5//KivDYDy7wMkQ2FvoAlBQskq2OekuXpIJlP+aGznMOJXZ8GEP/hitqnOjlAzK8q87iz
HQE4iIqJjlFAgMyf89zKgxzky9EFCGT7MkW5ZDq37JLpE42Z9Abi/pgJoDhMYoTFafsPq0V24/TQ
yEPXQLlXCDSP5a1H+gcdBQNW4pCl2qCqI2pLQDPpOpfQbuHOqAQqGLcywbhgFD0zL06tbniKHbgP
I9CmAPbm1TWJPpbwARCko2/PNbeQvl+wFOW3AroVOGWBfHlmWRHV+WIhN57oABs3CqVyd8yqYkjk
kLXoh/go+/+yY1OEdNZd2mj88693N3xtF8gGFM6HfIYBmo2reHslyvYUt6k9xxKgAluUe6fRo06x
VjEx7SxvOsxpoJDHnxVfYTNWmaScGOz1/2Ir7j3PS+AZqvmwhdcYsXBqhs21Zt7Q80heCNv/a4cM
JNbFMUH0bn3Hjx6EXBdTCe/QmuGRmJ9eq/Dkfejq3nay2eFx5EHzL6uCkjPWRUsyh/NCS8cS64in
H8IQtEL4VxTf4uimuUhbk8UYeFrEXuikxx5hwi1UQ2yBH0UORp5M/YkvtjADJUwsirgQssVr8zp+
VkhSIw1mCF/glNzCxX47EvDa9+bZLjaVL8vd3u1Ah9+LnTzI9R8BJ4NrTSARzlvqWcq3ef//PENC
eXv20bTE0wzI5kHRjS3XfxHbrsjvPiGe1ccjIHOTJ5aAaEsNVAOXVkjwdQnq8xSLiK39Yew82NjP
XfG8QiUcoAMZwnor89Aqkqk6qlgWdghRnJ84lt8BV56s83/0W8Dx6k6vlxkuZNssiENOUIYY6WR6
llbVuYplF0sL+dBHncrUOixwbtmyPalWaE7qNvOiWM1iNIzb7XWxlVVVu3S1HIkZHt2Jk3pFzgR6
N+V/KcJ6xHNd2IG4Fyv2vliwOnO/2UL4BA/3I+UXNtNUqtqk3rTRW+wXstc3KzIAVqQlzyJrx9JX
cSMlDRUb/k6UYgLrkP4soHl8QP0CsbuIr4pAGCwjDdtqJUUhSr8Z7wHqmR3SXMeR5/OUHwfJgvaj
OoSUqeRRPC4JPq+SVfWJUqEXly+kttIbDCod9Th5XJBBLMk1iSnyUwrNHooWO84KZ/G6JBhjqg1Z
W2M+Ov32vUopChuoAvzyBEjFUuM29C91t2SMib4Ja9HZJ4rVJZh0Xh8suFooPFj3pvifX1LMCz1n
5Jb2gsxzAs0xBk8bhx33PSy0FxmFzK1atRTVTPLUzPv9eQbmLRRjkR04WhDmZA1NS0qFpWKcJteC
i89cfZyFbBhg4D18vBPoiGDLSnny15K6TCjNM4uCEbSgEDN97rrc0Oh9QkggjrqU+eT4OikaF2GL
lexdbNJjeU7EEWVaVwi/5dMnt9nKz0IWQqp13I1Llh1u01gIRN/ObktzRFxQq3alzNzrw7MaPsV+
fpgGMI0XfriHCvEUMEdSGLBRJWijd5/Nq+DmoRTuLJ7wS3aztPeoZGxD1Gulpe7acwixNwgK4Pw1
bz2lkGglioQ9zOHuD96IRW5vya/jUuyTimxNkXJfDIQXPdOOehbxDTZM82hn6gedfBsdPX8X14Cg
6LSxauf4X2AT63aCb8XrLqJ1v5SJ/rvmVuIs8JpJPJbgpr94o04JuZVIg6f+nkBM7gVdJL0uXVC5
nZ6EQl21Lde3sTOZf6PNLQ2QhbRCMjJ5Y2kk8tbQuBSS4g9Ffw6OZPJWzraGXO/YoL9zMvaaDF2d
V9dzRVhfvJChrYuCldWOyluvdVYXT0XWhzzkHJsFi4JGMXIjLm8ltNnreomJi5fxUOI6xU8fYcFE
k7QkNs4lDwqeclX4aNRoLsaMRKUTmuHN2Xy5BLybutNlwko0aEUMMFMI0S/tlXB2za0V04Y3UKb1
JssgOI7EzaolUGPFbvwR/Z14bm4GNX+su9twdP/gb8QhA87UlmRGt+yzjT/IfvsUu2emdzRSBahe
jKNmp5O6Gd1p+MZru+2p7KHSL1VwEsGtjt7irF0b/OUzfmvKJEMQ9p+ZEbMVjFWQGCXTzGOAePZn
VoLl1rocQPBdBf/D7c9K4Sfo89Oovx8YgbHKBjJ1DBWbIX6ErSF37KYtdBkMbVj9pS8q+4/P7cq0
xkAPsNR6QTv9rxgQ+OLMxifcEfauoKzGcXGEu8AoMhoGunykBJ9SLfz9e59dQIWbt8G4Z1sVmeUm
WCcWQHM811udGsnFZeeaDNM/3X9D58J3Y8ccsxGcIO73c+RN4/6ktOPWQnndWh3Kt1xQhsUk3LId
xgOTGx4FU/qyXWa+7FV/8Y0jo1nXyLdJEQSwd7Ff0KY5Qm+WBptjurhXBa/ss23iUflo5zfyMeS5
bo7lIyFp2drUPtnMv0ZhxeGA2ZAkF1KJPQjhCmhJTPgQz+Bo4kke2JzORxuXatVzNR7k7rYjmSwg
e9CPrqvhJSjWSRK5A550KISTj0zQpPgH7GgnmqEjyvMI1U6vn+82djRUDHgyCXzsL35NgOM2h+nP
xsbFuVSfGtijput+cp37jzLNw003l1a+sSZ5ByO4GcUnJELAK0/FgxTpp7jAWkiOc0adznZWx3Fc
3VyKKAWoPKgA95P6k30ARJ0BdEkDzWM44Jkphwp/uonY/YPfECbFOerjR34S8QWynx1RcY7L3GTw
ojbbu8BXNhwkrzvcnFMNioYEPrbI5Wh47EVTwv77Uwk/KjxPujBRiAJ7tx/e52e+BmAKcIBDbz9C
O5RnwjjprWGVtJ7aztlT4d7yhfmHhvjbqwLdhh/w9RpCFjXm6Ewf3TcxCbqSFIgYArY665MTrzf4
QZIeXQnph/TalvMOWHPogiGKRwHlktlWtoypae+Ftbqp2H8iuQvEKlHPfzoFUNNxNiWYw733Z4Rs
62+Zr8TN3eWhGbdXu93iW/OBHvGpsj2/CKddN5MH3cKlJwxBvSZkQa0h+GdcZ1Pv9VE/4hJ9HkrS
gR5k7Z1BRpItKGu1CnMXwhfMgNOrNNyfn2l1toLPQL7xDxzs8a37sfRLscOwgzsudz7P8GiTdNLX
KKL6CJg8bK1likCdVM1k6WF5bpk7V8cmMGrjGLZ3advPIIk4RYQMOmLj/0lPKhDfxGGEuCe895sw
Wer31xaRyOfVLE6pNAjs4u2uVo2WZTu4KYsaCXBQY9raQT8LM8tZcesOxg8dBzQ/8wBlgWYDW0y1
btYphqh7tYb0o6WB7a1YdWPFnKGO06f//kLF7RGTOR6dNVvryqkmtf6pkTRyi2RKJnjz+fIXxols
QjmhoLiwKkpZUPcIBtFSg/vKNjTMMoLeBRCwEIjG9m2eeyyj5uJlN0tioa9fBXJFj/i/JTaeiCPn
UvqL5h7T7Z4aYBC9hsRagSATj3Td8fIbmmjEC20k+jvmOp31tAv1maaYornt9AI6H2jG7quqTNKj
Vf4pN+v+U8XXWe2vfkfMDfYPIZHQGr05fAHEaTmQ+h+pC3WyvgRqpOupJVXv5Vy5nRTzT5GbUQpH
cO6EbPhNzcTKt3KHNh6C7OxpDaIZU48RDQAmgfZWQFd4orWoKse4uMQesesL0h9bBdRb/vJN+Mgp
/kTm/GDmW6OcDAPA8PajtyHqs4rgcIPIBx3OgDbHEqtyzVqfa9dJBHf4H1S04x+sZrIuZQXIvEvy
pRXgcuO77bAA6XhnFC5Pp5eMcULL0bbR9svmGoava/iJr10Ygb9f3RYiVVT/kmV/1rfbQLzQ95ds
+gnpHukuqveFyxm69pPlN+XU4nn6+ULuGFwR27rYqf4cJ7t7RhBf+adKNdwUt6YlMrKLxKAsp68z
PPc6Y+z7InLKQWpOQYjNm7Z4qCD5/SXyCOWS/0/PxcMXioe/9oQrPGdOrqJo1PgHrcqKNyIX2wM5
+8uEiMOgV3+bWP/c7tJrxCl8DIiPGARtk24MaUAhys1XyVixK9D0QOqIqAbPFJ9JnUeIynQwrVTz
WqYSNdHQ5nAvlNHmOpxD9LUo1a3bbDW/mWgC+vLwSLRjnyQVMWiKvyHxzjF5PGaqaCrWk3X+mpIw
qIW5iT2uSMj3J8EFAfijsylGXyY46Ly06AXU3mHo60BFtPaFZmzdAVdcP5/+SWHviiaqm0nUiyQ9
nvcnJTQP8zHLRTcfERVjoKEtv8yahFcd9u4PhbdqXbZQOM1Tz5UuAO4ECqiboxY4xYdcquRH76iP
Q/+eHH64UI/29xZW0CHSdbPON9hygeYEVx/C7qDOz8Jj6EKorW5ISLRlBZe3DhNMUTRoy0cJv5DZ
8jhPRmiPEJYJvJlMoDfpkJOEGKWmZvVRcCRUbfrWwy6rISmMsgR+BMrSO08mynRxkIY6P/3cbeaf
kemQF/p0LstshGE72SvsLVYB0USsJbSSL98aXvW5D87DEYT99dkrTVOR5RteW5HJbLwsWkD/FYXl
4jBaLzZwSY4ZnJugclIj8ebgKtZ3bpfQQGjQPy4WVQD2ALOFCdyXqvbo/rTkrJFhCGuwZY7LXUrJ
XcpHS5HQ0N+1eLVT0NhQYkI6Y2tZKh6+QTPBKs3UnjDXU1dJ6UfaFd1ugfftGu8K5wRAEv0qdiNC
XrWt1PUoaMSMQ34td/dNNlwFIsShWkmQXlIk7oaEs+G43SF0jfHISktDB12xBsB801f//urjbMvm
1Usreur0HrLtOWwtM0egn+Uu3ZTezA1zHzJbCiMPunIdzQ2PN4vM9sUxO+Wy/etPIfmaLExM5IZD
ooT4n56MB/15UQcI5+m11EtAsBWhtGP192OEC1Wjj8PtM13cl947hBA/bEXOf2eCAlPTXQuJXiL7
1l34XcTn4MZno/SKsau/+3EjjsHHxJH3pu4uFpGX79fiLR34oGJ+SO9ZQBfv2LTJ3P4LcY0x3mg8
IbOlKRt+vR91V+la3+p0yffJZ7MxcPCRR0obFN50SB/TmSJwsr+Z2AMBUMhKGcIy1CwHC9RL0kkD
ZgYEspWAUJ9PVQ4rq8/c7dtoq1Mz0LyCnwq0Ubdf1n3pBFbYkcJz9jBlR7OxdrH5M+tlhIEXYq/v
ptVmpu2pi2oH/C/D2hiWakF5EXTL37WZdmA1QwkOKEl03SldGygN4zcnlQCAUmHJh5K6R8sVHEy+
TkNCodiHlq50+qVbD3ynXAT8qLomFiZ4pz2hE8fYeFCz4ey5NSfZlvae88vOechnnK15+Gb1RkOM
e/2GcQACBI6jyo1wZYRfOKKiOBVQFffDz6ApRgrCz2boi2C8sEkVkhJsAuD82nmabwryz4HYDEpK
5/3bAohC0ymRiKVvDzMUfwg4zYGO3F1M1hqeoGXG/pszL51a9djv8r/ZvZOlBxriXoFol8vazRJt
MT97XnwgYsyTeESVC7CCH3U8K3STvhdqbQ8EL6671H2kvm2mHq3xSSrACDCu0otvuinZsP34v8ct
BLYeEvc73nXWjjHf9J9+cW8fyOzaNdsOkgMu3QSjKMiZXcYEPJFyvGcfXw7JD6c3CWd7dXhxsBlm
4GpaHrtd7LsUivyukpGmuUrjkBsLTe11yGHvoHB2mevKXzd0eeJg4FBxMsiSpNSdZKTREhQ3g7oQ
onO1XE0au4B5RUypkyGS/PSWi3Ik/7W4kx8bcwx01o5Ezht/g+YYw7dBLWqSmlKZcOJ4sysm+kdk
6hijMQX6q96pxdqpma7MHbVmqjXbflnHLjeKEauWZpZoktZLIF+27a0+E7hI8ZqsHiruGv2BfK3I
HiWT5oz4YI+kqWnvy/dtVFLOgEcYGm4crBIKRFZt4jAsdXBNl2kXtPntRTQCYd58Qdl+436b0I0e
QJZkiZtzXKqnJdAJdhATCtcwJo78iZwP9ORgJoonZxeocXbsXtG0BqzRNeO+RzAGSwNm4Rri2nVb
YiLWmeFl96/MQpP8PgllqqErRB8iuu80Ceao6EjCDpVNBE+SB6XzhzndIPMzH4pP58R5LOJKEzmn
7Yv7gkOvg9gg9yw2b06nspYF8VBgllGi2un9kq1fxhxmeDwLj31UH6HR+Un1L/+VOX/9BLG2yRyZ
/BuG4+nfXkKu7yhQiGHPFSzcTOoBmgbbXJlOaKsYKhgN7cGwSFZswEd0WX56ia6mkH4ookl0UscV
MQgczrio52qoTLAHFXqpQmghHB7NPv3ci7OrDNDhq0zjW7uO2xvqckaNBLd2rXbTAyyleoihA2Nr
GN00N7mFY7b/xCK5/l1vfMBdhYXbaWXnl5kre0kJb15brNx5vuBxwGEVHi74aIOBgI4ZtxmBTpiu
Hgp/RPjZVxgsSAqOYSPQAkMbsP9HYyQUlSbURnLAoo56bPVyrB3/vGb7l7ecxAqw9uqFPxfbJBWT
7G9bzw323X9M1oRcOR2t7hX+m8t9pg23Kx/30yE86nbocvgqqY4p6T33rfAHvnUwR9qSbtlj9bWR
H0GppOeipyUDCyZCWT7ixU+BYtO/9PaZisFAFx9jAcBUV4e3qG2/DptWq/BuW0sFBUY9X+B15+7v
eFEnuSu/Lo0bno1qs6tXPI++r7Jpm0SGm/tKl+OSlSB3scy6W19vJVyaMuNn4phDOzmo7ix5YGoU
loaPDlpEHMorMnu96JBxPoq/KsZr5v7ijLE+stw8lHureRDv2PsQyzNiCFd9Rhu4RSXhrDGhq+v3
fBAXgkZJFvyf/TvX6BBDjJqDaa9CUI3R4c0fqeS3EFzkl4XL6/191/O+VQeDLRd6CjJbDJj/BZer
UN8nhaUsQeavwGbS30+DHeWWVdIEYU7Zog4Y2rRVYY/QxKTWD7m9A6RePJmb3UqurcYB4QKIt3xs
bjidQ4jClc0KG7Cxbjbekash3M8wvrAKn61R4oloZgMXt+7vrg8mgp50WylQFNGuTAJpQBhHWXlO
pXok3d9B1CMc0rMYm3wSl4qUfkoy1J0WkzDBXk7Ql2714UG5ZWXbvT5Jy/7tCrJas9Sa3mhDNx3R
/YlGgZyfvwC1Enh84Rey+ou9QIiGMXJ+IFzg1hZmWUiE5iTM7tAkso7V8Rj3DIKr5M8YCmi73Jtd
3hZGWrCLw+jYwsn0FtGDldYPFkWdX9cn5wfRhn6pyd8zmH+H+kI4YN8Gru9sVK8R/xv4YQU3bD/1
Q1Yf/j+BLpFcODgtSmfmWvzb2QZPe8csPdbR9cm5Q/3mfXvMQ9JLo92EPL5LaqH+seeV1Wg48kez
h6cqtmGiNAzyq6ddRw6X/4mHbkxjhEX8ohQ28Tgzia57fRgcyuJUKyZcmo0Vb/SCyYPjpEGWJkDr
ZExzl3+S1lVDheSA2csC7CRc8+7iUkjgMmAlrWuXCSpsAxsGVtBE2wWye4WEorunADnyhzm09D7T
ULjsMY9XaXCB5Cyhmgk86nI+v0IEkuzHEBaa2hEyA7M0ZIieki7hFYlAxaux4Y3IH5YHoBhGTb2R
6EG1s7lRP3FX16lfe92rySFxligvzFLHv+X/qFa04uT/Kunj+qgnYaAui+f5IQ0XAaMMmAoEV/5z
vuX5hS0L3HYyCwfBrBZSB9vygLVihF47yvHU3pgISkz5o5qEiz+74tDHTRf3U42DvLojkf4pOY6g
QpUsWsLGiebT1LBW12r1/sxWvJiJXhXvGA7Je9XSZkFZSt+YpuiCxEim+3zp+vm7GPtWhGJq+Jh7
K52sNuEtXZ+ZeNEgUCqt/KfNa4YbEe14KG3vOL6TT5LwCXQKywN0oxXdseP+iF7x4Jv+S/H0VHFZ
8NmNTMyj3h9KV/6k63CP2l3OEIl5N7LPAAmH45H4cf0WsExm6Bmnw35laI7Wpp5NzHDvlmnwHw6B
Czn34ZybXhoL9/Pa6D8zwWa3i7HnGMJZP6THjmhYrqPEA5JhniOVmd6GO38vb1R0VyP/COUSwBJI
okpeza5cW98cZFbDIEIW3t+T3fRszqDalilPHQipC7/w2KN+MjJUXbZM45msadJaEx9GOeiPHYGK
FiCUUxAg/mDWCQ6c6fwGAUc32DlZiZ1QV9rKd24m/YXpqYjhrEu5J80vdrEjq24b+JdkG4qkQ/UZ
kYwFLcxvDIsMgE8dCURf740D0QWQCkFjDiEWMfhsi8hidr19hwsOEQP/9m9gdwN7Jw2jX7ckdHvh
DPOoTQBALKgTI70E05DaQo+PIzSGAejJ8FQhrvKAOocykQRmpYAZrB6ELVbMSjVKiVZs41kjSpLX
731ctjUJRp/nYUMld9gA11q/B8FvKR42JoeEgwQYIPizTYjVghGuGNV+xmZYdkid2d/2jOkAEQG1
JdQrUjj5CmQYPxOSuXGJeLz3vMPLXpq0//DtkjxIUkoqpd5oFLLZEC52VTdXCeQvrOhfAlBYrfHJ
S2tvWyZ9Zxwnbw2UiusWGoGXu48tDprdC+JhcQWNxQjhcIRAPLRw02Fv2sFUljEImxDoRNgOG4Bm
S+YIKaSz+ukDzesegp4oPmnB5OBubh+9bEkzfR7UhMHUJlMRfyc2UNSJeXwEah9QyhlXGfbxXFk3
5UkO+pwj62K4zI7P7H0gYXVVJcDtOpLZJx/ykRjh83fAyMi40yeuGUrGidkqB00FN7h8FahggfQv
KI+vBpiU37vWHyXarZPi7lm8nqUSXa8//3f7UdLkgETowwqUkcpUdIaxEk6N+Dbr5igM41AWkwmp
3JltCI8Yl2wZr/1Mda44+JQCoAqymWE6uXN1GMlsjcC2keUePY+qtCBUoKC9YHdN7n1RjjmRZK2W
eVNsxjxHiPhpCQelgDoBy4NOphpoVzAosGIXNXd8F6qDOOKNGJcSqj1rkelzciqXBWQgt7kXX6Kv
LMoe5j+ORj6g/0ZyzS78BXsC0u6mzdHNGpg0IBoFBHYnCzNCx4WAh3dPAYqLRLhBYAOEc7aXRXBB
cJ36qhuS6Ty0ER/1JYzJQcciZYVwoZ03FHCkjKnr+rPKbemjWZ58X4ue9G11/FHn9iaJ9HhXnuLx
igrwriZi3AecA6NEg4Y0eqn94GElq/5E7/pn/VYQZfVXIZeuLwdWfd/zJ298iLghbw87Nnj6rM7t
CZltkG8FyAIkNLaszHYn2msorM7fUKZOixk5tpjhzgt09u8Yt1w8ITuh0R4K8N/o0dBhFYImJ6FQ
+FXAXjSJw68+NhKUE4yuvabLvqc/QPw0YBbilnRMO9liUAwGyliFOqYq1OLbu3oUj2LdS+XIj3is
AeKqNCLSlln8Vy77+JtIClJQyiFl/y0sJ069Sdy3Jbh9kTAamTE4T8y7EuG6w+D+o/Uf3q5tUFM1
CZOp3URlmTqiypeQAVPz2ZAJj55z6PgKv23Or2v07lH54dB9Url52H/c7Ydq76ZtHUxHTN9sQVZH
uazpUefy24YlQlgLV0ap0L/SiIlPvtbl/VHnBuiH5sMhSrw4QSN3qXZyXDu0IniEigOhs71vINSL
hW9BjQXusfslKCyqm+pcMAWc6jpSk8B9MMqMa1x4kP4o+gKuQfK6VV288daG1+YJkbfKYaFBW/m7
f8hBRs4XmhSDhrAjJWIhPq0nFtzKXacs/s5MYq8v48Jp7FHUMDYitU+dfKPiRj0/nmhqJ8X+r3Ax
MvIBviT16LVcwxr94iqEaNRkefQ/uehdeeuQXbpApXI4Eosoa94BDkZexWIEWi1E5nvtKDb8q8z+
VviWdndPrwY0151n27hhN3AZubf8c0SDZyfUlzNIguN/4E+wZjQw+WYRvILqMLDnDEjAVEITaZA4
MCowZWcte0CxV+r0ejx7z9sE+Fvu+2iZSbLAbLKtntd6BatzH9hD/PB7Lz1nt2jERaiSlsx8XzIs
0g9IlcJgmnr4XrXOFIlHmXc9IGLVJsXHc7P8Du0f5JtS89sBqLMkbJnlJaQ9PkxXhXJCnzDIzhBc
AV/VWG7A3zF4Y2v0Jaac5yfd7kmUAGKDRTAxsWW/sUZKIZEG/k1cSpT5oxk82BCYQZRznxloT2+c
AtoMnKix/CeW5MYzvhuts5Tf4ZIwWB2sRvPhzdv0kYYxwdBSZrA7aIg3t9+dZJ8DrZryPN6rXmCa
xeSqC2fIqG6UhUfusnzcbXavWI2y42t+GNMi9ubVpBRu/Fo6DkIlnKmR6iYvVKTWJ7yNCaF8gTcg
nGSFGOdtT1jIlHHClJtfFxQyFoG+Lc76iHqonAAOJ29af2EocxOrXy1otxBopR7UeMw7TtewFXHs
qGctcfdSaFAvjwkzRzgzMKCRyCoPsnYcMgI60hRqSIgWaVvt8rC5kDxe2AzccffBTfA92/LO6KOF
pevLnRtrB7H/sWJAvcIiJQipRNK1/mEJ1lSjNFxpgfvvKvn/ZL1gXNvhWvZKD36DMv6VCT3XzV8v
7Tj6L7bwcxIVyHs5PbjX5I6Gb4D9NzV7pQ2uqW0nvzTEmrmlPOfbgiJ5zE4T3UiyOYJzizAXxJPM
VFa25h6twxlzAy4MkJu8uisx2in5vfaDvc1eRjX4F0wWpphpV0NO00sVqJMjcmgz3gD81BYvtoJq
6+CJYejOZzk1WXSMderafBRQOt082yQBCp4t6f7aAirNTwS/bNoCAxbTgFxbeS3CYqqwI1L3E6wA
u6ay0znunjt5x66mNSAc9nVyxrxg//6vFhuIV36zHFljKWwanThkU8+WToQeA4VwuAcp38GRfiJG
ns9bCvoeHHnvrvgvxraPIn0OJzndleikoIi8EXSQOe4e/dhOsUhNkmkQMmQL33xlnpwCQpD3vosy
HVvJaQmJ8A3ubs+YuvcNiaDuhpLQ09aGBN8ll6oDz2US4ScL+n6hDY3V1bZi/ZyBJWT97rV5bAWq
qdh8k+gOjkq8LI4y+O3ugyfuqqFLjmB/sCoEcgHmf9SHDqbchRgNOYey615eOWknoLzHosVSd1rU
CFj7SQC+yU4i2UIBfZzPgYIkquPwkbImX5YE9NGGp1JPwCNTbBlJj/AyjrkZzs/duzBzMxPfQSHW
05FXaEtPwcx4BQwg0hI2wIROXVtvxMYeRXwpie94rfMQlgSwB7xYndLjAtKKx3SKnFM8ehc+NHIq
1WaPr8Aq3gQJyYY/bwXY09q+bWu9SVZqDga408dgp6ozEz0KpCvH8kRShlzsBBfRZXqTC8fSsk/6
yYADFuws0CIV9iGrloc2RfELyCd1atutTlxTB1AZwT1gp0i8Krsda47QnmcklLDPvxsar1tJN8gT
4JusOHRAtE6PtVb7UtcjioC9nMjFikiPAHWrCXdyMp4B83/SsJ/OsTcza1uH4yD3G/geOVXeiAsR
468FDi+fAFg27NlKpY4ysXtFv3h3vWJt9fOmtTfCNrw4MMGDS3nCKJAyvnp7xs9w0GM0X1BZxFaI
A9VDIjqrX8h3hKxhgI9Wt4Sl5DI3wxOsH9I87SE0rzOwRCVBaU+HV6R1CTtgSpZL3vly2RypRU+m
eYBBpWUgeHWlUYhbNIx9Qh/rI3JzL2bZ/t6yScx3Q2LKfLmjCHLfXk7DpRZ7eOeYHImKpIg1qqSA
RT32UcYWKSU8htkeDlo7CF7kxfuJ0/SnUgPErKe6aLyObBQvCMbTBX0jCczd7EiZ0EWmU591unIC
6ekERqf0H94zzhzfFvhg3wNVVx0EjlF/zVcFQoBd9ev2O71RJDAxSFFCtFCkWdOFdqXz5EK+Wh/w
kk//XdKLWuy9vZmUmMTSkky7TGb/j+N+hnodpJRw+NCCaJpbQ2xkqiG/Xn7XCvDOmP9SyJN0NL2q
TBcwu5j+PDgUkVCRASFbMtQx+vuCvy8KUOa8MYS5etN7uMdH5kT3QpneHmVi4bD682uEGHmcIwAd
NWmsIdq5K2TGBGsBNtS1DxKB7dLzY3DlDGYli5rlq1xHd4a1Jes+GlVpTvEM4/og2/AGhW9iSsqr
n7h+AqQMqGi2O2UXvqCJLRdd15S15Yjv7KexwGQqJ7R20hamSUcCPSU1pcTP/wbn6SfMx0AzHV+b
ga3lwaT767Ptb0qE1uKWffVxQXm2Dawzn5PGEpi3wUTCBS50QBcgvYR2b9Ibxjwt5lnWd6ATSbv+
oKIbe+7j5fEoZVea0la9IzQNvpRhdJpCNg46xIgwqbzSmvhywUgE4GRiXOVCz/lTh673FJ+cNmNc
BYZ9ysKOIz9+kjEnZVOEONinn840A1wnTbu59To8xeW9J6wPMZhqXEM+BTzmJESyN1DY8WfsDquH
Eo9hhofvUWQ5WIOjgus8ReWkm/nyMzZLwcc5AjF8usDIP6SbRBo2GWjkoIrBUTX8qDhmvlAY6vul
H3pyBADcuRq8V4N96+SGa0Xg8YOOh8CTqeqbx3EsXXc0WUyg1wXrcxBUf71XHc3I4k0FQ/76sT1r
0kxqy3ktqSdtpAwRKMSW+VpeHZDKKXqXhz0o4EmOhRWPO3TFWXAz8WzL4vP6hSGDyTP5fvN1sF3C
vSNo6mPLJxbBDleSh6qj5RJrHFzSfk2V+TfD35ms7WLTVF4p6qangB6aC9NBh5SzvLqkqIjkumQO
rIRDYvTQ/9iKXf2tLYrPqOIDagCR9ctyxNazCltQc33ADGcKhfDCRXfbKgFK1TZzV2r1PeZ7za9u
h7zHSA+2ev5guYfmH/7rySD3waXN7FZWm9nUp7zpwDW3Qr5KVNK3cumRY+IHeJHUy8DIc06pXDuS
R6tndRppUXxhk0bSeErsNlUSVcI1WVNFpg2Fd5kG3QfBFTp2yX4X7gcFjPUneORcg0C7AdYMgzNl
ezlzLLjBn4M9A7fVdx2ZTRSNI/VnNhq4RbE7r0SXUflGkyH/gSKFPo5A2YxcIqKFif5pg3ULhUQk
P1rGAMnCebjEGzK+ph9CmtL7+LB+XBJPTAlyGVOldvrsm7/gbZtBRSjGiyZT/Ks99t9w/0opHWAE
7cPLrJBHa9z7K29Qcs9vr5PW4R1d4CFmibalLqdp99YxcTeVeZ1qdrwq89dM+pdLKYnSztm0O/nh
S6B5cUWEnKA3uasb4ygV0KtDYAdXsg3NkYpC3zdtvLfrdVw+mQ5YtPnYicxaDdSGHJ8m748V13bX
VCPHrc2oFRMBOO9M9MVdPPbKmrfSuJky0s8e5zdPjagyVFPuHpTq9x1SHAxPBz+87OWdAYYpxCKR
RNmihiTKW1Ox5jOmkusXaLqEIg0ngJFYj8Sse6uo7yDX8rbvJSZX95yUB77TkQHorSSo1OraAEqk
pE5kjuQ+zBLayc3KrFo5xQnGO0+s7Bm7Q7k+kz3eEPnuiwm4dUXhPCZXRVomPKRR2NYDyxJKrWns
/X29NkMuwGrHHKvL3UR7p4TaUFfCnk2MJwPX5yw5u9PovwbYDmJnPVXe2OEuynmH12bdrwxFjPqw
PDG1xnWArJKHPO+olgnf3R0KTRZymx0CR29QtjCa0s99QAb9rg3fVmJDBSzTDIyiJE0kz0t6NMDq
j/zl1SitdgdwghHMaOUELb8E+ZOtcmzd1iAkbsabaqZkigdKgD3uHlfaonwVRc5E5BLVK4qD4aik
/x9Qlh5DKR266O38GtU+eYMiTX9Y7LPWOBUfpw0GwgbD5PhHP6pwznYh2eP6vmvSU4HzvBKymtV5
zQvYILKJEuoeMM33O0hp8DhHriskDedl1/Jmcr6KbFUxzLvM++6WbzvV2flwFa0WIr7LNaA7xCN7
fl1c6ItghxFH6qKRbUXeCLjxYgXJBUz4+fs3r44vqD87kyQq01o/AnTXKgS9zo8QzgmfZUP36v17
cZ8jgZH8MD1zKGjllUNGaXYxfP99nUxwAetu+uMzX4cRQnsG9iZK8wKMn+YV2ryMN6YU3kUnQfq5
+DWomFcR+ZIJ+YaBseYtyV2b+iLrFMfe1BUVzwnkb0KD4F5jROhxwPipqmP+mct7c+uWPJ+6WOCi
Fw5ZbA9PUIfoJGywNai7iEBDYPDw5EcEsJLGs15CHshArc3P95Er2O6FHfL1Io2hwq9N7iHDweqk
cERGUb9HEu1PHF8AYNOnONPkkHaQPD2J6ICZaJQSmdM+CD/ZS/VhNPgE7vHz3wZkmOofMC3557lo
uI92QrA74/ZJG3CjjPp4QdHFsWZsRbO1ViBx/H9W+rz3MH1UvMU6mgLLyTpSPU7pOOoQMoo2Zecg
WECJ8ZdcMwomXGtuiiP3pW0ANc3DEBBocMDDyJstBnebrei9mDU9Rk3vAN9OjYWda3/3potbZiiu
p/um9Tj6T1uP6r6jrjqW2LVKdmxUze+924NHMB9y1dhVOLWjsjZFMzAHPrUJcGLlKFI3lMWxxL7Y
q+al5a1VSXHE+ihuj2A3boe0PbLCMbez01K8EbnHllVd0a/YCD9otRJiF7dlmGrrIknxaHXcuETz
hu0ImJeGnSEg4ApMI8uzE6iv7vovvYRPBhfbgLtK8sQ59aX6EtlM6zuma2gwTKfldqqbL2EPokmx
NCs+HYp3DSxtgSp3CQPqStqLeI797bywvy3PnMmJbqgHwNfyae3/cHzBMlYIjuxM4t+SXr9Q/1X5
QPk9SQLjwMiIqqieBKHdyMQ5QBvhrvMgLi6Tdsqj0NeqHJmFBgpnItUC3+InBjQYm2kxm4wi5gKV
/u1plu+bXsXANDDI0XZusm1kWa8G5HlhApccHiUUEw6Dqdde2APcHi1ZNLHsmOksBCOZ3nwn+z/J
MIpdIWCLQidWfjt6X0s3hFi/zjqPoIY9kFYN1HH50874yN4Rb7TDYFk6eAl6PRQ4Rg7YmmoWOT9u
tyu3eVzdBw1m2tIZxH2Ee2SCQ8ERQcBDa/4cw7U6hEi88uIDrPY12g4DbHJ+CWvmC/AYqn7tP4jH
OomUwXsFMdtzyO10Y/CrqnqnjutkgAEgD5uicaRmttLhMhzJImR5qIlsrHzpuwfQOu7uSMl7Lriw
ABPkBIzpKsGYyimRdfvdrS/bu3h/88Q1o46sABxFqgE43PSA4pVP+chSYs4Z6orPQcKw7DAGLDbV
kZLyIlh2LfrnjGRGM6Cta8Tfa7hriGF/CxNzGetpUofXiBglOGAJbwak6oKnSdjxX+OdRFH3NDbL
3TlGq//ZaK04kY09AxUtUUqXHt5yunIIRM8fdCk5FPTzJpLb88sFpP5ZsF+Tyd1g+FQTEOBhBbHl
zMmdpRhGme0Lcw+Df18Hul/ilRucqvnJeSmlTWqhyEtopTqk2uqEHWOexc92ESJTLIJ22ze8G3YJ
RvcYNlC07TflmlT6TvxAkBDYgagb9X8luxAOp0xHxPd6yAwyxOEc+eAtH9UWoLhHP/J0Wbq0c8U3
SVykP4foFbnW1NRP460McbIOYK/fqRmApe7Vbrjs6g17AhdPjZz5FC/DptQ5FyUxw7q/YARQ0D24
M4Q+TF6RTfSelq3TQvLabLtA6Ka7hNIXI6nZsPnq5QhcGK1hS+7ad5+pjUqhx+xQYurQmstxVMhn
4zveculHgsdeLlyxuh78Om+QtaLHRzE0BVthv5BGjKVrvk94mSZ1WD+G4kIMtHXAwaCTmNH/ICDS
yCYxX+ySY87WrpJwxzUizjrhOmHpR8SYJ6DrhGxPPP0vVx6fOcFzKBzCb1vjPFsmI8G518fHQTQk
4zdWonljBNHoc1VWfVNs82qQ84qPSZgocdgBEku+r8yTBrE/bAQx4gybyYVf0UtqupZrerl5z4EA
StQ9oVBRwvH348Wh02pCGyaPq+ydVRiI+VOauAtnC4X6UlIBcGlKl/6HCHQEdGSA1+Ehrmymnm+c
e0fek6ZhjvOEwPlhK5cn8ohzlBb/IkVW2zrSkX9TQOSaDWw7OC59Afk0JM25NJbtS9Kxc/JYwPZP
RRwJuRrM5mJch/C7CViljtzQkMVhfj355eTyWa/LyFtIQQJ3FD8DeYYDgGkY0/vz854CaPziGjCG
vbLpM8HX21LNtgNx7/JcZucy2zRSbPf5sV+gD9+pAFS15ZQFRqlDknfhmrrzUd0bOSL+CYvT1dZR
/W50GuhYSibEHtA5gqK+R3dytaMNxUgk/5NHQXbUJkyktwdQ4dTrNK7qxHvzUgbXGaNwfZ8/12iS
1b4MehW1QCI2jHBjjzOaTPsIniMk7m8K+wN0E6btWalYzq2SToxupHjN/T39x2Pcm5wC+zNMbfKq
QPily7P2yDuzswpCBtG974BI8hNzZuyn/drd9oUKHcj2DkdBT1jf0BmarP2E1WGz6qnkJ7Ehk0ne
HwNSoX2FRwfpTZy6rIFxwSNtZg9o6CBU2esOsfEe4bxAHGBa/zupdJB8L9ejW409dD6j/Lo7vnUJ
dNSOuwZpn7vaKju+5sbX82FHOKHNyD1GBhc85KTYw5tLDT4zgeRHWAE4EuYT4Qk5p3lowo3cr87j
9DmS+rr3jj3M9NGRK0ae677+4p1JemGit9TLBOM3iPRYBahqqOGmyi94Wn2vHHgw+16q/SsR6hF9
JoKgdwafj//PPVebY8cEIu9UZAALzMJr6KiBuRw5CcZMO9bGSjWWY8720yhsDddDl0loJqojTb9v
s+7+cY+jdeDKON1s/TSjyv01e2X4EePn/TqkV2koSrh61KbpLZpQYFnpRT4snXmcxt6lI4eW0d0Y
0YOVv0KOibYxQqUIQden0gyz2bS9OlfZwMt00OADe/pU4h74kZF1ax+HCtY98kbNHKy1j/Qss69R
hFpPUZ6yMFPLlowxGOV2Ccszj2JGg7Ckqkj5JB0F5n/zpdAekp4RIixsygxBYezhA3ZT1JdQ6n9E
0N3CKocEnYjak5EahIzUODh+QLuxMmuGyQLoMU1MXMBJweE504HvT8OPk2M48BdgbTfAwn6A1nmL
nfYEUgaKzkD2K+FYJH3kat+Y0t1aUCSALDI11j8cany/cGFbZDmzjIvX0JEq8dVtLUqn9kyOVCQy
U8UHtxm4ucPkFMzu2VK2cCvTZ0LRZTvYye1Ho/G5etzUZu9xGWDi7+g3leYuhRxR1SLb2tWvVzxC
51BU/+mSx7sM5mVpszzpElUa/QiPdJsZD9ElQ00A5k62YHAU7bQvJFXe7IDNof3JIaauuTXvFwV0
HUo/aAktlqTqcC/quw+J8OkzijZVUCOrx53+cAu1bLD9d+XMVhy8gz8yTvFoqY81oiAFgriARQvZ
9KR0ajlQV5jGYDc+xxCLU8Cv+0Iz9DR4IKoxwFZ9uaTklx0VnpwGiGu5333HJ/Y1wR3pn54Wzab5
yYGAQ5qocWz971p/VXCtj8l0WCH3z+xEu95LrpVP4zk4iwppV/j5zk+zfmBvIQbc5zLnisjbGvvY
DmyJ5GtTVZ+5vpI1kd/1q4Uv4V5pYTfC5HGfcBYJTKz2lDyVcHACOBbGxGlo0Opgr7aQJdiQVmtz
ycd66/MNmPkro/F/+rGMYhJadXgVL3S4OpssG3as0SmoqmIkfYc77YYrGAxKQkfa6B0Tic+gkR06
OahpePqbhfQKhWzNo0Yzkps823NrXHIWMRC7FwgiBYo5gsWY/lTfMtBIEYV9gH6O/GzbGtu3sz3E
+pDPWRqf4OnupF544byGejqxSzyeeCGGEqfyvVHn//uOhZII2n+F20Tf1ZulJFEAKUBcZqMuIz7Q
hNLo+fN3vpQRVFTDI/AU7oMQwGgtpOH2C1mfezdJMvAltlIQwJgmiLXdNE/NYDvCGHwg0iJDzARE
+2AcIMKpW9LNf+yNJNC6X5sZkLIWcVx167V0+R6qWCFCQrIPIvds6ZbSPfh6fIhQfHSyNfW22Kiz
cubvyM5REQwD/Ho6ru5USsHQyXUoZ2g5YkGouXdkTc3pB4BDiv/2ccnQtgvOm16qnRltZNTSswXe
WCbmPmVABuK2dTwuBc1pYXg17+ZA5WeuELvkXXfwszHuXpcRp9sel1xWpN4joftiIc/5BUcYEv0W
3cUrXHPuQzg3OC2xPaHNTq2WWTAOXMOxuq6ndLjYZsruB+sVBXG25oPouU9j1hbA6GUEKKqIA5JG
PE0brjxL1A4GbZvENTosL9I9Lx+jIzWUZ7L9hwBnIXicOSSbdHtyRpQmvGJPat6roepv2+3Xoryl
tTDATqNImk/gJTfgGrVdBD8msCsHQwhgo/hLKhITw2dTMl16lPVFfJGJWLeQBmw3gTdyPyBJ9J3G
NJPIYhXqpcCzKhvrgu41VCrGIfpb7IPChoDQNORc1KZAD4dRtYBssx5GDEUGnDzRFx6lJm5XrsXq
j3j27SxUuQ0qTpPhqArFXWoTCogMOlLKm4mBT+ww0ip24kE29xAyigU8UQQtV5a9j20M53MsiqTe
RUzeK/1cbwUvlw4yXCTGrFnxlzDvO/kyVLeGZl67w29d38+iIgwjsUJNa4xXJtGsxydGybWo1zhD
jZNFOz0XeRhONy61ne+pbI/qOJfd96+6/8UAJS4Q5eUC257bc1a5wIjUJwEobhUDdImPdEXzqM6p
pRJX60FhSoEHkhnOOPsmyawfVLh4ntGk/MAR426U0abHBGXJCD9i7z82a4xAN7g087rmKqAaE0Pl
G4hl9+wZzIik6hkPJsG9mOe+mDymJvbn+JBBxlT7R4yvhx3kTVouhyckX2OytvFKfzV1GvjoX8eU
0lCNzdf6xiAPsV+gRq4poEmnu4SU8dbr+IwJoUxkzig00OgAdzEuiq0Sw2CO+vEHqQk7bniAh9+J
N2s3572FAnGgY09v+DVAz7NCZ6w6aSsCj+gtdBzwUpNYhs9Pa9Zgit6L8LM6ZV29akHsC6AWcYbJ
6QtvBywxXwj66HrCx4caDlqVVr9EIlSXUXik5Nwf6EaK0djRcVlsiLsE340gscAqaBWgcslOpF0Y
Cjy1TRA9zQiN9jccufsoDNE5yGq3HyVSvWO8hEjh4nhSzsNpW9v2S6Yimph//Tg+nETeZjkhrvn3
rozk8ESl2+Cswk4+KwjSzDGdJoz/yMdrehe3cxJbw6A4L6yDwDkkf+pGyTUb1MtbiFNIFfxxhV/M
33gmQA7+18uWkTrOLoDd7hgAPU69/9IzP3xddYDKyQFJrU+lCQ3ZtbjTOh9MCnT6MZCD7ICOH2Vq
mJG2MAXIxps5UBAzGtC8RdwD+VIxwYWuEwBh0nPPi12qfidZHts21V6PYtIkodWwHh59xxp5MyCC
pZ7WsJbpqtn6z+YYSbutcNpEZuEZBeqVyME1CgXN7qgJlA12XgoGGaOxNTiwo127MDtz8JKybq7P
DX6kkZE7uTUpnCxK6InHxfbphIeFSo3YTNl08Yj42eOYB0GoFr9nc7EWFZM8gGM486mebKMD7k0d
hwkNbcFa0utj8VcAquK6earxmVf+aaSYGeIhLtbVfCTXHFDNDIBAHWGQc2UBRfz61+boX/G2Svpt
vO/WOzkdlz6wHkEqaInIjz5Af6NMloV5RsVh4DBEtyMmck1ZCapuVVZexcZU871hTgHVypU6Mt1v
J6q27lEmiBUTZde8vGtINJVj2z7hrWqXwUEjzPyNu++csXW343V4hHtXdseA7se8uVOmEb+Ka74M
S0fK0yopeLH7mTf0LmjvMUTFIKXnYBaT3dXrLeLH95nV3fUec4unLgOyclkevSpJ8uz5vvMfitu+
OHatKGL8B1gjlHPVNpcuSrNgNLK4zO2rmHOtjPCiFx/7JMvt3EMbC7KjtV0Md7tVhivY5+TOF2db
kZ2yciQ85W6bCcuaivDMnh59zg+D+bIFmuHn+kvbkKct5l5OQQZPBNyQx5p55+WD8osf02ak+RVN
bJ6MzDhFo3C1YM4FsMxGBc4pqLtovoZfUukJuQdPKWoicjPVMRTxSHoWW5i9JAdZ6DTbOzOS8f8S
7M9JF7YsrNKMwoddfa9QGoLmk/qWgQU59OG8jctF7EQdDNcO5KfKR0OZltt13guzcYfePdTLVUn7
U/J7N4NDMCGS8kCeCmZbPlpvioyrlZo3vbFyDfB8UCeoYwvGDLM6EfcdoOnDNS1lduI7stmQ7Y60
G3VPCREggibNvj3AKC0mXzJwcxuoVp7T0mNfDeK2bWwQsfzW77gvfaV1UXbQ+847BugdDb0HslGo
/QCRiYFFPv3bNrm60mkQSyQMDu+eQR8MhH4J6kVLqurB395GXBK6fNJksSfNLNIUPodamdbm89OO
TDK5U+Edf6c2mh+drvq9tZxnnGUNbhsIwC1VX4TRytyIvRor88TPGCXevl1lmuzlQr6rZ+GlizcR
Vnx9dAMAmZ06/2Fqma4UWhUu5GqKoUzXMZ//U4Y8yxiyG1exoRQqURKTni3jQGgIuHpr/tpUZchM
KbzhW1hN0Ii3fTxhgMrKzoHQkyBhS+wFLiHVvkt+sw9Gt2YEU79JHMTp9J7OwYbOrfF9YvA9QO3m
xVN2I0pNPT3rvmo23TfvFOuPzIAmlP5LqQ3iE4BQrulURPYd/6MTt9pUxqbuMbjkblBSQqpLWzjQ
4moxBVF5H6jSbLa3Gympv+S2TEx88r9DAFO4r2rUACyBl5v1ZbDZNc5K9ukQCMkdYir6rh3Mcj4q
OiRno5ZiJj0/QdJhikXzu4UQkuA25cl0GgDN49wg8Xorb1rQ6CB5oLL0r4WBlzHw33kMSPqkZVq7
ItQnSeYcyhPE8quPwY6hg0twEVyiu0NV9wkjzByN+7qR00R6cj4oKgLJYJV5iWrxOjETv9V7EOKu
0xn22p35Y1N9MI+jwKxVro+wjbl/skWI8jCWBJcvyz/JZRJDpUyEydTMGgGiXgX7YnNyNrlYXXhg
FxilbkTEehug/gLyclGq6hvkMMhF953fiQmAJoLEkkm14P2AUC5Do36T0ilWYUvAIcqIdcaT8b+N
YaonMxTAx9wPnVbXz49g08728n1lspCtBptY4W7heR1ZI8KXz+Bsqrr5xBC8al3t+vWMRFNjoJRM
qDAArUSgk8tnh9Mu1+HDGomnKKRtfoocEhOmvuEGkgdhghNnhjMaZZM3h4D/V5eGW2hjM4OB/Uc1
cX98LW4TKln4DB/0X9JtAo0BE+7LacH+SOTHORyoqb57WDupad0O99BFkXoO/jfEVdp7J9zSy1lk
qBBefQaRSHaG50V4pKyZ5y8IHTXII0R5NSr5nWcvqF2afmYK3hFIaAu2hRpPnQXOx4TcfNFLPhrF
uLEQZGpmg4XDXY/11n4ebTiW/rU5scF4GXbcN2mbN5UJKm81VXwcAVHuDoTRneReStVlavYFh1C2
zghk3N2q390A1c6jHv/ZL/YKXAPmRd2Pz0ZoH9gUCM5K28ZOAUgwVA/oBG/oCXdEbCTjMjkWmllw
4enfw/2QGvqgIaMp+KkZBsKpYYLtn7qBPuoKG9UYTZ9bMCe+r8i/4W8TJOqjrQgUg4xP6ybQZmYk
4hhy1kvJW3Eh17bDi9EhvGVYoB90BoPnSwFLtlDp9LmZgEzemdPz1tyGHg1scvbhenFnTbW+4DfH
0o0oh70+KVqHy/ckzKE2IU3l594KZNgleGW3akkz4r44RoEyh9toChXuq+DeMtaOPDBjY7gopQzy
/VEoFri2W/LJ0hOnVZFGg4wSXB5G3iDQ73ycq6AFttzuzOCBQ2oBx7vlu6oR4DqVvdoe/0HiQJuQ
jm5fuBQGfr7QRYMMx8KaYTp0YKUreS4mcipRuun6fLhIvfHELOTOvMpzX8VOjhQ7lE35Z1IUygmt
b1QI/VaVs08Km4DSVfvUS3zpkLXjhoC9siEEPtYnOnkoBVCqQLSo9jcds+ZPLv2Lh2KgxpnbfhX5
2V8Z5vG6VKeMw/Pijqkp3ZH3L2jXo884vVCY6WV5xAbKlRR+6B1TErVd7RmxFZzRoVPaVLLRQ2HL
DrnpFY3XwbCFePbl+KNPR7IaYH9ZjCNednkHXa9uIqm0jUCeGmsL+MMk3tPebYu+XXgczyKsY6Lm
zywrMc+TH6QHXUhzBwdfFt6okUf9QjVksyx80kq5SihI0PFApdAhdtzq/v6RTDPOW+fi3y+q7tBh
1uchasl/Vq7oHmKPrscToVc7QPKtVuDzToDr5XcMG/wsvGKZOI556mgkXc50WpX7+ADpyqWyuAXX
gsbAaxcazBhkoX6SVG3gn1lQmOSUkWX2+lFPP+TA8psDYeF64gs4FRE7HjdhD0KjlFg6kbtc86Gd
Ng6LhuOKY64j7Gw5767Xcqjn/ByZdHAK/pE61nDrAaD2OvPNHrnDwyyUi5dyJivfOVBXwIli7UrN
UkR27/EcXDAZ6RstPE74tIAIK+NCuf3wBF+M+1+IUggr6geRBekb0sIUEht5N8YSKc+X9xF6ksfQ
+StUpwiq+0LB4X7HvwZSViLsgIzYbG5V/yjxgsnDbOP0GGnp/fUYNkxPxNun3CkNHKT9V8GENC3P
jVn9qAZK85shOE9/EuEoXZ/RquBgLA0n4zIkX1VqtQ3Vn7brRUBQ3VeDi7sDsxKLOxjraW/y/g1r
yPw6ZSK2yy+u5A0zgVfCUe1WyS/PlxmissS522gGhTI/z8GtlpCJ9uAgiwD8iv4NNYeJ0Ot9IRiY
XU5SESig5554/55mt/PJBEKW5wcWJPCZYOikOqHfzqFC6pBRUbCl1yAk9zakomq4PKrddQ3lTSN7
+1R8r5xTtFPq9NdiXdmz5qjtQhqH1W5NxDDpeM2ydz7xAMTiSQ/6iljjCkdDaxpm2S4mOS14Derx
RcApbkzWluLaRLLvBWaDH7D6VD7P86Ast4CcnzhEOG2KStfDWSuUf45Y1dwzWdLN/eaytphfZO1e
r5RrPFq11wvs+eZYzPSIJjzQFajenbzFa5ZbN69/ObhupOORYGtQEI/2nG4LYaKQcrCHh9n+11P+
Mi92DaftKQMoMS7zDVnidnzGEOBv4W2FqrGZcjGdAupF80MeERt6vY7rhb/mjm+53lFT0GCFLDbv
DLRCi9OHsEJj0ua7D945B/lW4hjGFWXaxOluHKYgBt4zyrJhqRSRAc0carZ1U/A/JgUDuZQckSmr
5XyDk2F0Vrpwr9H9ttxwzvMdNKCVolYlVtlBs2uGIPuLNNaG5KGceM3KHYgjqZ09+8HXG4PwjBz1
1MZ2Peo++4gHKCrJx4ATMlCtluLMM8ROtCmq2qe7PhF1DsfjImFu4EIpxbNSXTI83H7n+fHbbmGM
5G4XkqZ+O7Oi7OUK05RZIx3+MORNdCGAV16NgnFRmghbN7GuY68vf5zWoNER617134qwzkBpRu6D
/IWWmpdWk+jJeeU1pVSjFw6usCcqIVGSvSGRxzeMwLO9LStlxJz/yf1PCwPqMlPlGrUNk/hY8hfF
jLo8QPlA/4IOwJ1FGgsrKpVj/KqrEW+LnFnADRhzeWu3U4Ws4g3FHxW6FQIrh/NvX+ULk8CzpUHo
bPDcRvvt1d2isMiawjsSfAj4HDmEO7T06CVqXUeIWR+9RBeQDY9xFDJ6G5BjihIPg26i5OXUmy7R
TabuT7mWAmURmU2M6HWv/jrhbHV9J0MAiT+9gTxf8VKogOhWvZOOcFpT4X+7kTM71OERIVnQX5n/
gIAT0NBe+E748di90OzO5OvwpayJaD9pjpf5E+PYw0pZmR5rn4TYnP1PvasoTPq2F5huitu1LLj6
OLX3z71EQThtSsX0KPwhD2ujQV9aG2vzHKrWC4E5FL/BQ03LeErpKa5cqkViwPPn6TrJQLJdX+fJ
qHrSiYoN03yQCkQ/L0uz/Zj0NgkN5sjUTCHvFuxAFmlfs6YkSw6P8ArmGHe6kTe2Ce1yzHu4JwEX
w3VBnkXSB8QIkMOohyHmO0uiB9JQcDkmY4X3OAEYCycAe8W/erC3mJswN1EL6Vh+RpQXzylGV/Bt
mCGbWGVUNPaMjO+nLhq3MLHAhQY0FeyfNmzDkdv5/2rGB9Q6QFPvq55jqknTy0puGrxP/1VCYsv7
rQ4nBOFHfJjgzBn1Mt96wEMAVFnjoiT+n+DDF+M3GNLuMsdbTVZzINbAMo9sLU3v1XG34zXasbHP
WmCPPiQi/NcRvyzU9m2RLfD5MY1rhbBUeOV8/KWcVcXtC5p5XTbgP5iWoVk8KsWPicMGbTyR2uIp
6IRQaQs5bIN5kkW9qycbYf7AjyrVRcocevuNKJUmfdr5dMuhnbzw4Gza/F2aCsr5JP1pXTXC2C6J
mAs/EgHNjgWAVS6+xYOFgiYdk/GUsNSwMEnHo9NSkShgVkmJ5yeXoG/duK5gxetaBA3OwOlPjKPm
DndWwsILNLTR+AYplGx1C8pJrtjwCmSjSARxOOK1mr+iCBJ8YAmgzwEWtouvVYk2eX4DlFBpl3+f
j/vYVU/bKhOoKq5/TPacMVSL4gIva67SsDo4HAL1bgymHODvq30wp3vqK6DWptuT87GfnQKsLLGb
ixiVANEI87tIFELKSRKEnSx0nx3W2anmz8DGNZzdSJ/81wuCPjDapaYLGVzvQ5i11fmRE2F2p+PG
oiBIcZymafFzydyzIprQGwppg0kmKtehGkHz9L+tJnULJeiJ6Ypr7+8xRKpuLzHTVFw2ZWtPRVfI
2fboSYu7eOUz4CSJ/tcm+I3hj64VBvZyfN1cFubG7j398qziyiEzWXW3lYjxZfif73e3dLIL4SM+
+MygkvMKAgMSgQNGAHpA82yvuwG5+fX/VuN6JxO4eabhM0oaDH8MTYjVSQwIl7cjM9VjJ8x3NTDq
jM+0R2NubGUyXg4k8LH4hc9neZVcnEcB9OnA5BaO+H3XofOHL4GR/w4e29sV4E2rtfWbkYe3bIdb
RV+X0fveFCeeoMvBnva9T72RqQ4oDeCPXp5IM5AqLIgCRukLlXAM8i5GXBXCtu84ZcSkH0+OIRFB
n3cXytZim5wAmgJr9pyrW/SHrtOpTm+S8RpnxjuEbUSxvYSl+XjttAskpXEXu6IhePKw4MhWNsWZ
mOXKOaksdeofO9fsjIz3Dcprviw5cS91t4Cqyr2CeaNdkSk3WCdT/ZjkoKbe+CjYiOCMI2srUs/P
Nj5WoduWPkFzD/RDvlGTjglIIOT1aV+HU0vApbDBVTcY/obr2muPWigcbxcMBttf24n44H56fXk6
Is88od3A9qLoFhGe5rNHnFlRWPQ7wlOsVjjw5fhaVxVXQkS9bXPVpHEUE+NcnMIKZOmO+1a2wmhy
WjcM/kDKXuphH4dB+/F3LZzqazNebHftrtrHhxk/ZbiVwj59/pFnXPsO7p+kk6yWOLsQgFJtjGui
2SzYkAtlN9Xp5Ei175Aql3mO6pbkjeOkLw6BGfJwwdW2yEB+e13Po9IJi4do1nC+KIHX53COTR6j
SYa//qpn6BAJ5uFjEvhDZwAxJNTIWJZ6rslEiKOiUb+7JL7NlG7263Br0hjM1SFZ2wmM/NJLDGeJ
1I0n3317vNpYLTEaFt+2nAKe6AyNQ3xw87en+6D7qJtD/T68M51VdXco10AwjLTKo9xKWYWoHUvx
HsQdT9J+QcNe/1UAeTVj3pT1Q8R4jZtKlTC9XXr6O2YVE+O9JDSDj2qx+W8JYK+BQo+9V8ifqaLI
SlaUp27vT4LpWNdIfixq/oybboHAx2zkRyvHoKKmDORQvB71qSN+ODCdvNXIs406DwR+W4WyyVL7
XuLNYzg4UK/FSCVi7cX+oAoSIuYTn2mfz3MK6cmJ418mNtiNATd0wvM9l0qEZiE3/7PXAGaNPnyI
qimaU5DHiOQzgTI3Ab0/UaaPjbpF57tSojUxy86IJjIsUY0hFCJ9DX0r2q6xPjLz4EQ3SFZL2gWt
3nDA6iDnfrGNoJFC/FSA7mXPF2KgTKwS5KordKyC3s2Z8PRsQLXhcBt2Hg9R/F+AVpKQPPSoP0ZL
NnAanQ4Yb3zLUA/BI9wWvoD8oZmJMJPHmvfSuroHR0oTDxEmQ8C0TwHE2b0QHPPQEMvEG7SAfKNG
iU7KsgqGSKCVSoWaDO2T8ewtN+WSe/lK8EojcbGMnt3WR/KAiV8X45jRr8uFGQ+VsOH+mobzX0lg
fkFRwS/xg4FnivOLOsmqTAR9vLlhZMLjvM9ym57+nohLU3qu2xEI0Q82+wBJm4npAlTSrOClY6iY
EXJcMBLnGTJaVXvk1wfKJF6nc1tfjlXGTU8F/4CU2eT/P/jtY4BOY4j8i7aEe5+cI9sTrivHQCMU
wT+139NbrTOTwKZcJOipE9pTPTnDsgYlgexP9JkQiY7yGn75Go8NXjzNJvHS8LOg9Mt8Gb3TG1TX
xEDQ86sMTgdIquSexERnUIV9eCAaOYvyzUv9s4gpIgMbJpIn5XlaCzcj67D+2ZWP6KLVp4Rt2YoF
5A2W6Nfgae6UqpTUPyv+SEGqAR7tcnrXNTIcLWX8rwuj3bhLCl6PXr0cL48309K32ml4w56MN8DD
JrVgXFWrdosdJtZID9pPBLwwCOpwausKNjIe79q4T4OkOypwKzdLVWxd9bLI05SgllFzflSN1aaF
PouXFsdd0dDD/VQjfIWJ7p7kA1DussvYlVxL7WYOLiibkIAG8u2++SKAH0xXYOBQP0kOlX0CDyRO
RA6QNvQHAvFJefAtmNkKmzcWkkhpK6f4q0aOt2/DnPsAJfhbLXcMwzUsLOz8cmau6ySK+u4EhqtY
d5uYQgnfHM68Oph0a+K2LM06ijn4GuZH4IbKqYe7H6aJjy3VFxmtfxH9Je4Bikq2Vx45WXjhG3A6
ZpYsEetjQThYWtqgoCv5sXJs7xnk8CNyivfwdlRaCy3CpsRF+8t9BJgHnbPslbA4R7eEZPFAVdrf
FA3iKUBJW9bRv12/WcLBvzVrMHrB7GyuWrYzBW3pMprvtqZ0D5EB1Q6rwGBEFeWS5HLyyYCHg7vS
fbvKBO3eqtvlxqLLg+VoQG5ChhiF+wdWtVQNfT4Bh5XvLTlr9oza/Uchhg7rS3LTD7rBXHJtTyvo
0cQWIWtrrRzNcq8NBmO0tR3r8Oqx0mjLWiOG6u+eyA1WFoXWy9TlUHl/NxGEbWz5xNWTAr42IW6f
H/bl5ONGD3TGyaBsWjJZhxtG4SM8isVmNvBhjXlzlLGbwu6ZKTIykVCqBzJeur683VrO5XfdO7WB
Dyxz55l+UCanqANZuig5gU5ZEadEdnDu/EqhdvlEn1US2/5WF96rVCFq19Y1CGsr6do9VKZ4UeBM
YOFCep3/KDPR+gInPqLxYYIfC7irTzBOB9L0Dr816XEhcaF5REoN04oHkhPbLufKiNzEhfPxxXM9
G6lNEOWn/EyfarN4TLODYiuJb/oK/9zLFJo5a+Am8hTb1wAsH3ej0qI2YYIRyE0Eb0xiALXNyQHq
vn6X8di6l5OBPkaPVMYvtWm7s8Eo1XvZ49axOb+hf2tjCfBBqLVMHQmK+th6HtctM/I5Y7aR2qnt
k2aDcKx7ItrXTREU2w1dUrjQZcjAiJxl3gB+E3GpVVulOaMD0cCPT3yumTM85pj0Iyj0/JFNI7RX
o817DlK3yTi1bltw3sh1ouBhIo1F5vWm45NWLYcZd4Ll5ur/VjcnL+yuW5AHdag7/XnXecdO1zGP
v7DTNPxEC1NsfNfxG+5Rrj/Z+9JFpOGlg0ufGHunRvwqE6ifjQIhhgxjOXTWdq0KOs8GpAf2ZXRd
hrttumQIUiNJm5BOlh6VMzaM1/OsKALxNiFn/xCCYSEHSYrO/z1j1abJ2w1vIeYGkkEfJCTNmIdp
DvlfOU4L408FAuWZZBFBB9AUbd1Z++UDU2UerI5ihZjx/Dn4LKL76jBcHmdTaM6hyjzY9zSqEyOt
FBa2efVikouWuKR4YvPDdlfqTa32p09dPrfTJ2hDP23e7yMOPyIQkjUDkNGv9UWZh/Y6N7Sl/u2q
6IzcZXXWQ+RXh8/iXGU0sesDW1OP/j9qvxF0hEFUUhLNCRRb21SRQJPGGgYGfIljDJQBwaNzcz9x
uk0fVOCRBDdxfKIaCkCoI/F2EKYc/GLHstoLu+7bQqr8UrlcgQc7kcJTwYUaDBuBG+WjteMOg3Gk
prt9/JP+lpn9Qrwfi2gJmgtKjBaEddSJo7kbIjeSGLibOjcsVtRt4NS9GddqTOTHNgF6sKDPXES4
cRYMqeJPRu1sY1VwPYRQnKEKslXALMfepzxxq1qS6rBlenU6i6cWpmsi8Lqo9nO+IOMcla4RqnKd
lH6E/3v87eqLKj98rqZIB6UEhjYITmg3ouI27ycyYGm8WnAHzRPw3PsyF0bHYfKC2dTAKwRcuwsM
FhBF7lnOn6c5SvJ7snTPll2GuxN3tdlQvBw8VA8Reur4uuYbohPmFvrjFJNh4dgF6CpLXm0gSEv5
IgatwXgZpjz64D7wXTR7DpEvxmE97SGqJKV1OAbLk+aXtjAh4ThEhgU1K3952gZ5cujHAnf0em09
8wWC9avCEFIOnE9OOox5u7J8WRt4H8cyRzgsq4jayWvtrKED7jc6I5x0ld4q6L6r2wCwrMWjypvr
pkZhzv4Zo9YPEW/KzrVVFK0ER/9D1gbWm3os/GSwnxXXfR0CCsbXHaEhG9spLWVvCV6ZQtPNRzcR
pC+7/S8xlvsAciwawOrEF1/gMdg8aKQ0bKgPGeUMsz4pvm0tK7HFTLIvdZwwLHxs8BKbvDRG3QLI
Exy9pe3G83CuJ6ghvfYoeui7xTv/o/v2SEnrFvvuHMTdpvXcLvkzG4UNXtUpq2VwteZcZYZ0GI/S
huSKgf1GGbh6zvN300QdJTRr81UMAk21ad3dDcvUhgmpdPhEu5MVu7Hz3Xc9Ax6H5yCnK1BrcF/N
RyTkdcC0xG/OOnXGuGsC3XCfrZx3vtz05Ci+MNLJgDEClbB9dAQs3CvvV53sH5+swXAez5SP/n5y
zxmxIpZSFQcDfuqdomHutByk9VmXN5yuOCqbrU5a1j/JIKKkgwQk5QULI1F2WNF/wu3OF/l6dz0I
TiKm1NYEfSaqPck8eeckYFUO3tU5mzsRo/Plv85pzvBM8AL1uxhHIVTENjEAvOOW0hfHe05Xt2Oe
gMD1wHB2GS466aS/9vF0kCRSTYqgPuXgvp4eCryTiIRzSX51rFMHifwvlKETrO25AiKiqp3OqvZY
SA1EDpdOja/YZ1BDIIx+CUHXM2nqVZDKRaeqLex3i7pqq0WO9oovQO8RSKQdMd86Ckvsd1hclPh1
adE1ptwOMikeXNC/QkEL4M+K4knQ0Ul9c3YF+pj++xrEO1zAAkQWBiomcJqwo5yp7jGocPkaW3bf
iXhQzZMvGPPMDODbvY3RsVdtMhaGCpzyr54Dr1TRQFDdpZBeQ26rbtA6L7NHrNczpf23/rMzE60N
JYDcvcTF02qZvy8J2GOH8FJkhCZIUJ4nSOo5XyrV1uWre2XPJXRx30zGQlXLCyxcqgjaH0ZZSIO3
D2HtSuyRTvremqllm/GKbLahEdzXT9NhdG3MqkvilbR1zy/GhZwO/Kf+zoQCCD4IypKkbHi/3FOL
NNwRRO0znedzvTJzsNKuaFK3ANGuSdHq16xyxVQ8ph8v8CJPyfjX9EkfsRp5hsFYJzI6D8qhXl5j
X0jh8ryfo+EnX0NoGMr3FzcWnP8qmEocS7uCt6/orZLxQYBU/FQoiM8vrW1mwokImzJcrXFPMfEI
JYM3QWSSE+T+opqX35b8gOo9QzwPpz700wxIaY6VU8lt/FcLVcQVXZjYjMwFUTo/LWvNnHHvtKSb
MHkdbPdzxVySNdw9xDp+6Gsj7w/r4lX7PxvgPPGTAPZQIwZhl214KcoaBJW/7uqEi6PRRfijessu
brShDoKdEctpzqqiqGVXq+HSl4bs6cQKQd7cNJbMznCxGmgIy5bBb7AxwydDQuX9mXJKz6gWDzUO
Smgu5HR8FTRPyEDG1Gk8hbPO7egmow491SjsYX2Kummkdnuy3/VnRn5SV7UbXsf6UTRS238ykg4E
6DR2ICgpdDxQ3YoEBn9QlvV/+b+5+8ovVmxt3Ug1LDbuoXrpV4AFB8ncm0mguwW31R/TLxib+b3Z
8o/IVWtyJ5pC4H5lNmV69lk49CQM6vIyQ7j0dO3fmsnQL/j/hlZiRKswPXrsKctcTrS1UbZzl0mi
TZCemGlq8Hv2BAuFikvtJlsZf4xBgjvDFGg9/DmKV6p03+701YcS5HmGUk2AiqffeCfdPWZGYh0K
zto+2bggOf3NWz8ZpyJpEHi81J5Ua+C+NPNqiXyUNgJmVB4xDLhRQcLswBEytlCTfU3uY5X+Tg/f
snHZ9RPnSjlwijqxfGFcs34UGV3vs1Rnl8ERk/ofBJ1vmUqDH7u9Tu22NSdCze52fAOvUGPuSviR
28hbFUB2PPIHG+utIqPG0HEj9ZCHISHBoBAX1RwDk1rVOkhtzJs6BxF6qhQrIoFT7Lao5JwkTPh4
Snb2iGM/R70cCqmxEEuWhswZReaA6p7fvs5QvE0wH5DZf60QRg745zmaWHoXJFX3V4c/mjVgykMr
4klL4xtFx+Ab4aYZWKXKkS42yBI9y4/QYfmau0Gv7cqHd0wICE7ktv3ZDKGfs2C/XHHyYlEFXo1P
wSSKXOBImeZ1wrp8JY8yqTxSqAMc+am71wKlY0QB5mEFabzeVP51L8gWuuLWOA1qQToAmWKws1xl
WBeMZ97gZ9oEkmxRQl9u6lcmRYMDVnDQkC877ivL5A2CIr84tpv4Y9I5JQHmPrpqHF8n51Ii6DJf
tG41wl7dWZ4GhEfvFybhrzp9rVNPHxUuhShqKxrQOCpnLGKYjFoaFT4iGJGPGDddU43jIXiaEHuN
l6G1T8JT2rRF77tLwm3WaCRWNHVDoX+LcJu3UnlufOChvXU991sDT46mv78S0F6gv1RPyFB+nECj
9KAlhb922qi0PTb3y9bh6RQotQnMA1mU1eX+YRoCSQNmYD9jw/YB2EOzUf2sJsL3AXU51Vhg/Y9Z
4B2iHy62rcnskrmKogNmBVIxNGBfbnxivyxNUMevj1LU0NlwG1Hi0Guzq77ayMpQMUUuamO81AkA
nt234lffBLRA8f4S6MBFAU32zme0MiXlBNMAa+GXOIDs5RISDpMbMdF/WQsw3AZeD24CK4LStlgN
zVrQklnnKfos5zR93lFN+PjYJADaZ4uZ7FIta7MrTpx8TAJmrzqpVfB6BLP3Xnzt7W/4HsLaTOQP
nGZGo04fExrmlTk1c0lc9GDvKuXFul/JMQ+l2/YmfbxjNdC+01CzhBkL+xHH5gob8v8ltslKk9mC
66yKPxYT4eQtcWqBOd+utea1vdNn60N0/BFPpluaOT1YV4KdTakG8mOuv9/VJQw/yifB5fUU7avE
5+wNkmw/QLjQRAI5wBOWAi8rPJZ/zNQKYtFgQEdPbJBtii1xaSmnR56mDWSTF4HF4o4gcGGrqpmT
kcqw70LhBixa3npNv/ZZ3dDWCPmecL3u8Gl/bkFpZ19nkk9s3mWBQPyWKOHhWxs9FtyjOcAKUtQR
anwNVzNNR23TXtddUV0an6xJDG3GnLiUSjdZmSsla4YDfVSFomQ+uRwknwccf3lBUdGVohKTyi2X
muDu5bbCrUVf9ecSisPHVgxnVJVCngcWcQ5IMdzIw0hknfFyx5xRQfjECH3mF4wTyXdAcjraHZna
ZkgS+ZlJuIvylcAWXHGF2IcyEJcLVHtrZtzyKrH1t1uxyNA4P44+UAxOeFOtRyW4xhtLOfythy61
1dkQdJBgwSRm32Run3sZiRFM1WVdlLTAJ+ZxMFWMHRwAQmlJTrPQitV8m9PFQ8qET1ttNpmm140x
hioMgR/rBS8gJ6ISWgf6Aa2KVpVIgcBsygmdfYhBvAbPnnEdgnrloWJjrFb1Rhynl+94zm8OZsUO
JcZhZbqpELTHEHl874aL8gX55ypnXk9BMHP+zb7fYTdQ15yjEKtQwvRBc5bsfNTeFFukslpiKiUD
+1BtJ+5Ua12A+Ok7rnmNt8089859TE1hcth7eCuSwAs0ZevYe9wAJG3xm28VOzJyA+J/YCsrww1a
ZEEyRuKNtqZ4xYpJZBVONm1rLvlhSao0KKO9k2/gFWKSNPIOB0t/LUk98txc8kwaUDzIzEyOiSSB
rHYb9jBd12zExm7jqkJHcxpMtmXHHjQPmx63A1AWuS/RpjuxXeRsAfx3MSLog3GmnlyOuj7Ayrvy
ZA0r6ggTiGUq3XITdHrt5h1gNpI7Ct5m0l5A5tSiBRhyIRJxJOCZLiAJLikCg5dk4nbk4Idk85Dn
LehG2nFTvDkvLbO1cfxeozqe909qDXaO7dtrsauKglkkwKtNSyWNFDYXaWDU0TLQOeVZyZ7dU6K9
fRIuiSrFM2TONljAlOXLS0EbkTu5Xwd8Fp6OIKL+SmqHbqCMBt3Lkb8pwgTnKkX7USWV2lo4xOh1
obK4SyZ26aduMtL1ijE1ENnXvznio+oLlwGosh9QU6XLpuwJ6LqMUrAOuIjtxm6hDJbiX3nA5qTW
PWmGL0kBOxMIhGJXn/IifJSMgWS92ZwhF/4LgrRPiLEGlt+83+f9Dbk/pZsGK1tSMdy7JqgXpyhC
dDjrGIn5MFv70XE2IqFY1BYc1hhibrQwXSgb3TkhkmYoyt+5U+ehHYOSMY5hlBN7xMMlRrJtLVEw
Ennij+RZQK+g96FDKLtB2CMTHwjlPLG1u70iKEQh1DcHo8gelLGRn8T5P+bHCOkv6iAF5pGnXT4A
7GogstUrKBQ5PAkw7QmrCSz5dM+FRO2NbLYmuscOmDLihZrfQgxlrz++bG43X26l2T6qymshe1WK
spWd/IobSlFwgCG9H72EGCIJ12l0k5mIza5qvm9fdSdi06kyQywY4bxHxwR2eiDjfNBYR28vDKlr
XnvJ8Hjv2NIz0I+BFSb5Z5C5vtJjOOBwKqWjhVFGQxn6SQbZCl0OOvI0Ij5ENK4ipl0MdcJ64bW/
x1juzyT4b47IyvyxEg2IvFSaDJU790kmYm+96HqXPJqx9DzBd5eUnqn6JfuDtU317YJAGFhrHQAB
/6k+emTqvm3TPxV1WTfvIP6jFrbdWpmteLXiNmzS0ZV9Nqj4N9oAa3GbNYYK3b2qjquloBPxt/Xx
iTc6as4yvfGKmaoyYTd9dPfZBytUI0wTRA03LyXY6AkpxMwmvL2oolCiJDzXv5fneW60TQ6PLSel
2GU3ywg9bSUnqMVZGen0tsAGVnAplgTdsfkesK7gz532AF2SbDprd6JJx+CR1B7ztXha/lzJQnlx
k7tb9CB5R3BKBCCMBB0lIJzNooI9rl3TI0p9+LGYjvGoIAt4K3JuNz0jfNzODdaMci+6IcVybvzM
w5iusRSMN2bogtcL0BcU7ES13BDgaRWCn45fhAhxA5RB7C5vzF1lF9N7cVocNPNs1nu8yn8HCaIz
Uf2H9yKGtCMbG+4uomi1m4giu/imXri3Qc9gnQtM6fu/JDp6EvtMA1/CeFIBGl6c7vMZkJ/06q5y
lK1REx9Af9sYkhkaJyWLqj/bhurC8DxBEbKqUqgHDdofsfXDPXtZIt0lyX2w6FLmqZesHmv4hxpG
rzs701GBXh784ZorBbn7ALv7pEsMDIGfIW5ZBXr2kbM6Nizr0W8JimhQMLja09yrGwVaB2JTNG1o
FC8F6txsKnP2JUhA4FpmayIO50t5NR/ex967pYrNMaL4QPDVBebjLW/O2ElHxOVnlHKaEV0aZWBH
iSzNAHirg3h2UQynC2CeAy/7cG/Qgqa3tksj0hvSXNNMSC4H68krBduoPLhGKvxAB256KI/i4d9n
BBzsSC93Jjh+Fptk6xkzXa4SrcbRSNyVLWUL3BVt84GpAGwoy77blr6ST96dUhSPnJ9dlhdAq2WP
PUZX/nGjalT34GkZJ4dbJTxX74QbBZOoNlcD0cnSzppq5JNqj72JxfjiYBuwy5gXB0iq+vbZJiMi
YzS4WtmvzO/7dnZsXMAQu91RK+KRbeKxicnL8WBZh6AsWid8m6uqpbOuSvcqXuZHCPl1m/DgX2u6
KxySWqMwNneY3C7JEzgqXQpS9NNoIizn0Ehkci2xFR9NE8wGg/sHPDjD/XZUgqLXZX86GCSEUDkK
60ebJYR6O20cfgEll0BGhaT1GXS9SozhHkIgUzF3EhgrQzJsro3JSGgVO3a096iyY7xl1mU2R2Of
HlAN9k7ezqeMGPeiXL4Oh20DDtoh6+cbUejn3e30T488/0s1q7s5q5aRvgOzY7iMeNyzOmJH+tjP
Sx93coZdVX2akbVQXgfpKjRiAgK6feSbSp/iQbr8IjrNuMz1BT5m7cjH99SdKuOjhEcxKl0T1l0h
2aHcR50+9FUDJK6OVRfsq5HNFSAOOS1mUaUhjqztxRa6N/EGOm0llxkt9hYm0QQAlBszqkeEr/Tm
0TIm53UMomWVF+yDEdscslopjHItORSNEyJULX51Wt+pca4P/1It40zFD38vKHZbl8SNyk41rG2/
Krim8WJtiYOH4Tqu38JE0VgPgw2CXntNk3IEPR1ez4XJxCWNRtwV0f7k+GAu34ag7kopn6BQh82c
mvZyajP81DRokJu+fmAbLWfadJezpKf7e+8eowsh0B72seroOw/lrmpS8iFOVK4S4ZE0HkCFkkOZ
JQU7O0cntxNu0Xbw01coJP/gf26flu/tthZ79aLoQ1UAwVC3HZClVevuI47QCBlcoymSG/rkyJzs
Kepwwjpd08STegJJ78KsrbiwEU9NDEk1B3shobx+7C1IS0KXqjs25eFBxYsxtJ7y3qcStG/a1ec6
6846MVWsuiIwaIbcoxzOhnZ0qtFEK1db3l/4inTi+tExHiBdya+rHsr+2S35ILNJKwCDQS5o6jy/
rrQ5FiiYKK3H8NbLW9IZwQIhkSLi6RxkZjxLcuiAipqfjzEUZ8PDzK1DZAIlqMy5boDwXKmqJvue
aXS3z5qAxRk9q9/Ppjk3Y4+viWUjJxLEKsOByW7nPj3Mwc7/NYW2hYyeh+7Ci8n4BgQRJtumr6nB
pQykCpBTEwIrweGsG4d5lBlwDA4UeZMtwIO7BzMWgGioSCxFzc+AevuSIAFfdO85JN1HeLlm97L+
E7tm0zr8ye2wsColetaYME35xAYfkJSFg/khONH0DIOZGtQvG7fWG7UYNo3et6yBU1byCn8D87Rc
+Qk2orEEw/uhhMuaDR5KXO4UMya+eV2BwTvum2GD443fNYUo7JsYSkBT0n1UHRYQLdgm25BLjppF
uNq0G9bwNghoBEL7Y1ks0mo7b52k616Vdimea+B1mpNtpS652kjx683bbUy3cnkRUvhDYSOBHqoZ
RSF4Q7vUBweOA2BoA0lJWvcvE5mFGAF6TKlnBurhZUktVg38hRufpcaiPiRFOhqS7fxtf8+6p73q
U8ewyr2zj0zIDqslHHPzke6KgfQC0WY588xRnlKOQthJUJee7bXPniHijb1L3HNo2Q9HMfwlD9nD
UpDe+xfuidqEG/DctvWsji67nw6k86bh5w2TbGdFFpBGC12wDEhwwW7slOEN/oo/Qfzi7X1d9VN7
+7F9Wlovpk3/ucYjy/r4vCXXmDcSxh/4w4Otfn//wNX/aVHSuAI4SspxrsLDoEasz0OUgSISPeuh
Gzwi96yyEJ78QtGr9cbAmFc/UXocPe36C5EiXILKW/7bnF/0/PTXVJlT+PHa2YA8ckFQAXQwvwSV
gJzD2mIkkZgzPeu7Xe5IM5FSivfFW2WG4A+L6TuBr+3c4uxftaJ5XqyUsbwPA4A0XkYYRYr7ewta
Tu8cPW/ZBh+rpEuWEMwFNOt3O2NeHK+QpPBtti2mlABC/PWNaIi4PMxvqJnVmw7WjaVnbvOdV6FQ
slTtyoZ9dy930kxKPRncMVwvO8GDUcF9mvK7l2M2cAh136ISDCBKBkXINyc57alYurNYjWdlKHGX
fU63RsHuZNFXdXiQSt4wDN6nnPqQUIIj/1GWziYchkeBvf0SHD/fbYRpFcirg1qSoVjXNBZi+06C
ecUpV0OTCucaVjbyoGhOdY+BmYzrN9hJ1XB0O8CSNuwoadDsQ3p1x///xP8TKjTt8EGiCNG8VDKm
JOLNU9U6rt9MwSpuzjsIsshIZMgx5P4we1NcZ9BdXk5H/gqWVQ30C+nsTSdB0JpUWTP5Wj+I6Pz5
UC2nWW/dBdUqanqkbtp3Lo1WcMIqZABo3oPdlGMllZvQ7iiUyyJ1m2hgM0QOoumhwxYhZSI3K/G5
UOAy57b5h9/N9KZrYeBLvPfaJoqvzQFE2CwwzqUDdS+Imnla7fFW8gDNHLhv8WAKXGZS89vEblO9
RsLLh0jN7+otAJP4HqQbfJeIBUHfCHCOjbeH4H2YProWnCBGzAYL+A+OUw26EvJ0E8VVuvB/mwqP
sQSie4T6czISXeQo9xiQq4cVbV2vxHtnMtvCBLOh5JLIFEMQu21qMfaY3Bmm+dpOZ7ZAIwwOKVkT
L1+Nt2uYzhY2K1zQX+5rv9orkLIbCc9Yaqe+Gr31a6oJqhE8tFWVUa30y62XL5v2S4HL57b7cEd7
nevR/TNuAt3oXkQMpctQAG8bHlFh5jPa6LfLUxwqtWad5kT5Q9UIQ6POA+gVb/HUSJmboEZ5jvRb
5nIjOKsoEOGlFdlYsTAmE4gi3fot/Yt5gkYjsgGl55Nr+/Kc1fKOBPeORtJJwYa5Pouidhh4yRPL
9RBQ/rCusRsi1LpuAKoXaqnMA6v7es5C/Sf6PJdQ3vmyy1sRTkOdRQ/ovl6QLGT1WiFXWIfFb/H+
eiMz6caeVu9TgX8ot2+F9CfQksnhEhN5hbo1smPZCpoWvA+BjCn2Qjub8iefBYBHve1XoRyUD1tl
8BEhzZQeFrr3O4zXg6OrscY6cl8+bUFN6+9OhamaSodN1WNcsBU+vdCJ+ryZDmGzPU8f1keZ53pL
Z2XVw3QPIXr++2tu//SxIAhcrSpVJ7yQsbqY7LwYwYzhRFfmEREpH3v5QiQzU696yi3rAMS4hD6i
4LO9/GjA5+lcvJFspLLwiSlysEkoK87arLjK87Ib9L+0cNFQAnQtP7BLu1bgkUm4FYqkexIRSPsy
rUMqhwUWnUb8sIkhWL1xCEc1BYbtaVJxwjKyA8v9Qzf13Rv8Wxs97MbUIHr9PogeHodNEDuWKGzk
l/OQqb7eM2617q2GkKZea/2qjeHWPQhf0azaUuYSJC1BfGLxr4jouyvwvbMXa43uz0x/6ov867fo
aThGXzRplEZgUJtM6TN4p0OalVonIiQyftACrCJYCSgZrOrmkuNGS7m4LQ1OOd2X/eKYyQ5o1buX
HXk9kO4ZfhXKfTNoTLir3YTJdzz8cilYvcpSImF2dS/gDGtrrX0HkCM0orsdBEcHve1A2XQlwHgp
feWW6ATzqFR5Sl/rhY11LMBdes5ZdvmF/2Gj9Mi1mufhpc4SxXwboa0IkF+kjkzADcw6Xxtq/mL4
Xvy8M3xGsKETCH4YQG9Oij7UP7fCvVHed0nxhqbo1NHKmyz5vKQUD6jpvxfQrWmf76F9zHurTaDc
4uRtUnF1qwSLoI4s59x+LbSPtVWadfN1a2S92uPuFvxn0/XnA/RLYVFfew773gMy/VXjN28CuJmN
INi7oyT847NmMVYNiObf6BgPQuUl8cRO2GRs219460Xn3T9lFg+pNyyEgo1tSe7DdznNLnSH/3G+
XbjaWeSBRJ0Q1EUO+pSaWnt2hOqTh+GUINlnRERBULe7nwMZ9lOqkZMvZFDAgu+F5DMgPirendnq
HcNYiwikr3kW41MHTmJFQ+D0YropQfa7Yj4ghnZvuj8jxQXaR/MrknMHrbVuHa6AZ1krSirVcAbl
1lE7UUDChTwQUPoV8YwXMWVp9EtzCU/XK9fggW3HkKn2Sk53+pN7qvxlcRqhm1f4LgO0QluVecWF
O0167W+egKiKbp9EIk2U439F3ahCsvOv63kpD7O1sKt5jcIFcC9lnHZcWevmp51Q4HZc3ieP//wK
YPiMZbpvElzdtluFjOEsl1dQ+IRcd4UAvoArTCP2s912F+N5aGhDFFshuMfaILVbnpLtASd14nnK
t2/fDTO/k/6/DzmZcEdgWAnFDvdDi05T6syv1IEC/LMavpp9uFVq4svKuL/NQahCNgyCXqXHXxby
Kgnh74Nq9x7fqsu7LY3K5RUkswC+oyaANlKPoy8ULmfT+/L9iiuf/qx7oHBKT8VcsvEIUc/d+lBV
FQSG8mblAfBPGJtTxZ8Y6ICGbdqcC57Hsq8nGJNZL9W2ogBFaLs6q0aSI62nZCt9+r/ouXnj1voD
VICA57gxKttL8PITaNM9w40Cp+iXTRj/rn3BOOB8VAuUABwGuKviu8uV2IirPX3eph089s9k7f2l
WZze/9kqI3BxFaXgXg6E3tC4KA959llKt6HTNzXTTsu3Jg1JXUiN8Yt86m1il0XBFaQnl+m0NPlT
rjiAok50ja+gRXy8JR0wpn4r8E/T2U3u8LzeA5YYP/tzjKUIG0Wd+rLXGb3keHfNNcfx25oWiGgk
4vd3ZDVkHgf+Zny1Z6ZznRYz7L3jQyJRBF2YMeFnxlpIoQD8vW2pYd0Sc8wjvqmmoBqsQ9XspN7W
vIqT5HGTV4dI/Rz3DmYXiwAcuVWn5V6VXBrhYY/UHoAyBw68fmTD06tWK6w3MSLMyS/+gonxBVLc
bzKIzIXSubQDY1IcTgzjZKZjXt6PJIdkdIfuzkGjCyW640QRTm6bVTCOSWW4wtlSt7VLYumXhSx4
rY2hEwN+OP3Jk7DL5PNItiGX2+IentX9BgWVNbbys4fe+3yYN+6hfGhpTPAGTc++lywmbtFjppKN
G87SyKXcen5kjYHR939diIml3z2sNDZnuxnmy4mTFoGFFjllMwhCjlJNmpb85xsw+COdxa2sBkkp
bhmTOzlYcZtsqz1Ky21Pr+sq9QZZVFt/sdNQbyvDezEd4tLTyIXiBgVdhPMpswlMzwWiWjI3ZHaY
ukVhuQSbvG9/3LOL7O8EF9D/EQyIRuuOM7+YLrmnLFBFl/qiM/kMJ83cy0H4Eyy8/z5jKeqjZyQc
cVo1vUeq+Lav5ZMpU6kxyPMBZG7Rwmb3ijb9CmqhvnKdI3i3wx5u5V+wO5WJhFQIelFnB7JvnE5W
k0yErlUHn/jmXtjxd/loBTCAyQ/iiJ3BpN4O3LVlrWThsw/LMvpylAx/9TRq8QwG7XvVquf3l75g
Iug99oOWWpChTPG2RdmwaXEsxulupSkpINCpJnqFGNp6kxHXBLvEAtE4pzEhsqYjFxt07umWrasQ
LRG1m6Rouubr3nBS4ypXqGg8Jlpu4ULWHrfnZfxLwJzVht1s/CJ4+p4AuqfjOkkNexV9IqKv6+YR
jHX2FDoFgzMtnmYizGZK1dhLWFI66Rg/2APJaXMS7UZnAKHbGwHERLBvQ+VRQXz+lmKl4NN2Jt9O
Ay5DvwVEjuSXVj1iPlwMQtvmtLzlKOq3N7UOKfLUA+0fAdtp0PRtH+urX9pB9Bbx/mxuYAGcEjRa
kkpgT7ctqN8l4/F7XI8pRKAPY/gNFWEah3Ytey79hUOuJyWJzaYGREe9KkFm11KcujQ9t7hepE0W
k7VGq0Saa2a91pYqdJGhw287GEcZNZxC7MHem4qe4sJnib9LE5+FV+yXdtV/NC+CnrPsNmBWF9cQ
XsBSJZbxlDTa4/P2ULItigti/66o4jcuQgXxnNNIrRLGCgBvqvOMPF1w8uaV6WqO9JKL/s+wn51/
Jgqo+N0bo/e4+zx/J7ZQCCUzQzFZNXnAGxzr6jxEFPAQkpcB84jDUQ6H4m2a+WFpHorVtNlmc3+J
AY8sF5qqWmBeYaargRV8Yl4zO+Jmo2YJi/7nQyTwh0z63Zk5mTgU3e+S+9cqEPrHw4XUbvh9jmog
seXhshLimeIpITEwJWA1CVz21R3WNdVptLrnNDepCCuMlP65pFfJfX2i3ntzq5T6il61HWEtLmAP
Bs54efj/o3fb7vWR5i2jjZi4xNz97VFAFp23qCdVVPSIxvgE/Ftv5c7Eov3WZ3e/cLO4F/CqfAgO
3DTJ85O3p9ChsiZQQ7kdQtqvGjiqv03j72Ya+pZwlhGMdyWlG43G6avry4ryNeoXl5/gSkLIW1Y2
LQ7O4Cf0flXJI8yDU/sS5JjdGUv8ThRy7BrVSk7GaDwhRbEjb1rsThXHz8b8TH70ersfL/8ALlqp
I4QxJnhBUBlew6t1mtHJZy8xMpvY1NL9HCObO1q7jJQiJmmprW7GFItpDVz6T/j4ZZQP1X1Wxlq3
aFsWVZHSFZV++aC+r8pT+xN9FwqgfU38ezqSpQGFZ9JzfisStYXnRMQ84lZqzPeNDP0459vOUcUh
KQzdKUFviPcFkR0WhG1aAl5Twbz7Npq4ZFv6AMnK+jnO4xU+cpyOJuzimr9xtLwCqDKI8cF3VcCD
LPRf1H6KEy714Oz+rr2NFF2egIZS+gqCtGcDXx6gZQ9P5s5kGIqOYC0HHFw8X1xa0iuZ721d7l0z
gK5p9bLa1ivucs+rwXpInUgegulVoWSwsSMpMrE8H9N/ZF6f6cJ55L3x7mp+xoWrnSHJWKWKXDWD
Cth21liNmAACBgmLhc+XbnezEkXRwOrM5HXZLBY2hTUFZ1TpyZMt7LGyZ2xyiTmN5f05EFsvomZZ
ivs+SGBRGwXssvSVplc0d4Fgd6kapumYpnxkROFEMFl0e26LgmZ2OB+eh5lF0oC15rRzJwT5hK8t
/8//prBRwMbkJsMaAhCjurfFOGhs2SGhngfl3PkGYXaXoN5oQCUqH/6wt2ivVnIl+yeWkVr9m+Q/
0JfYCXbcauA6c5a+Ow8sCNPX/nQcmITxgRfoiTWLL6GN2LmIcUNpkdcOBV3ghp2AxOmsI0KhJzPp
PHAQG3zcBEpN3MEWIhe5bWpCFmWnNqT8fPGPqWvXdyUj/Y64LiQA0cVUd/zWUZ5D8ilcuFdDGznd
Ek4wfUE3QTEQQcuCJH8Gms71bm2VkxBCShUqdd//DGswDVTLSbBj4MvDUKr7rEpx2G15D65qc2RB
S/W5grBQQG0iCg7G+hONzv/HHTqE9+rwPX0ws/ToGfWAHpC53MMTaFJywqmt7W8AuwdoIIn4KvMp
STF6onz4lWdabrVuWN2iqqf1u98N1XLTDPtD+zy7APpQbY+NFfDQ2iUE88n/MdEd71ZisU4wNgz6
XyIe+yTVNN+2wdGQj+07MdtkFaWsyVf2I8xTsbbhxU4V3IAa0dIHJeSmeQzVK3CMSEUWwhxuSS8o
6REBWD9oRcnld2ExETfqdn/jZaByWj45gqdyr0cpzYuxM/D3l1OtKVSuQF1D3nosLD78V2CzLuE1
8IWdzPBBAM+f4J4rdeYgq8x8N/Vqqo++s4YRiPygA3v+Zb8pp9pAXfg6+gxw67lWZ2R+GkAUW8sz
uROM/BQ7kq2e0sUi0Cum/Wg6ro+PRhg4/JdDK35ius7NJgu1VN0xIXvcSMW7dk/ZBPoskZrMPRfF
3u+ocMgBxyQLG7QLLvlkfTuKqGgiwAITBZHza6YnYnHlkFalmqo/6x1G1fC0XyDmBw2Uf/LmRYHV
u/sVpZ/H0g8JaKViKehXMdyjgmQtY9XTiqhqJ1MADj59whmoCF8DKG4uSw7y1x2S6dxHV1K1A8tk
BZ2GbOx4a2VsYE6XGLFnmXnRRfmp2VVxxXsYUFOfbtqdxIqTXPQPySEAzrKXBr0RdsI4xmVezrnA
snjUhr/YijKCA2iGWVc41B296V5bXn7p0b7e7lEIkrG4CvbJJCJpZD/f2KCLHGkJUzu9ZoQDGVHe
xY30eQuvw4sTjx2JQugjHNn7adcGwTItsNKchgOQcm75XeSkU6bvC2vh7e067Hg1lnfqKVfR9T3U
WNRoPQngm0mmJvHcTcZcq7gFhpZXeu0IFqdEJeHWX84J2mHxdH744zX+mG9RPmeAEyiW4Bm6F8q9
qg+dHvhTivDFA45ucfNGddkbFkeL50qDpNsVaZpA9bRhiPTfUebtPq3vlTjSn1YSCcpHMm90r8ub
kCcfgcgvQRpM4jag0soG//TaPhH1kNBNMPlIeIS7JkDiVKVAL8p3Cvg6cmvTvjxTr7X69MOdwOVJ
IUoDlAzDQFzaDrEM2zg7gXeK5iK/ElZN35czejI7+hCbdsFhwyrO3MCHvG2fGHrwTErD4RAyMR4W
s7eOzBqEcyHE/4rHwxEjsTCp9XYeugi5QGG4FnhMKq2wWvClGTJafdosCFFKlFkb3AlVcC98caGu
roCkKMUfo5aTQ0Y1QZB1bV9MFl5KlmzZxeVwg+sMU4sPBcIrBbOmUL5rI5Th1z5tvcJSwiD/MM7G
+oSwBWjlM+Ic+mpvy++ZJ7MXgHA4M6dc3/W3IvHClYvY5enxRNvXFEoZoQ9piWdbw4lvPqQslDvJ
56Dw/WhRQkQuv2R1mMmRaDY1T/G5fzxxV1UPW1oNt4nek4RL1sYVw8tbH9mkge5PKF3YZtg1HAYZ
2VZuCw0U/OdvuPJopcRo5G0dNWHOPZY8cbjs2QkL6FxOR7MdTML0V1G2029GGgZ96Cy7edGY7FCt
H7BtgYVX+NtfR0fEGswolKcXiVTln7MGMFhD7COlCk1YhrbYkQ6vtJuVX7WIyk0nh7OCm5I+K6fV
yM8Zf98MFKO5e4ju853u46SyrujwUiAspWUSjvalicdI2BXelF/s7ih4OSM7vL4mGG64RdwdY0Qt
nGsiOfJPWuAelK99OwR5wDlqbtY5KB6JcU8/+UuTYqkwK3BZ06Qn4U3f6fEiJsLG1DPCwYpxaRMQ
WnumXMVmT1PNglF3caDqYzbHzx7qYxhCJNlB2wwzgREgTlVnuU5g4eUsDz2RPsKy2d3WyD/KUVUg
tJCigrCvtajacBsxQOtRSadpX5G90/bfZGO+V8IUue8u0DrbizJl82FSaIho0VFPqTiJdXP4a9Yi
h4PLwd7844ePyn9+c8zrYp7sVN8gJEzliLbAW4X1Dclv8NvpnejwWgmodzgafJ8vSc6tNjqIzpjv
R0d7wy9MGs94Z6k+OqbINEb3LNjO3sXlSLWA+69zKaAcVb2NdN/OJWlEktC4WoMBiCkhxWiylasT
EN0YxHPh73PpItyChWUPQE0XsncM4ZfvC1VHfU2wrtHNkpvm/+bAEGsi8J3noLdIaTkhNUlCDmFW
fLeF5uJToZvbLyJfRP9vN0SPADTPuJuScoirPgwFrzG70B8YA6L4fgE1VlWfGrCn8JZraoY8FyUW
T4V3j/GFqI3qrL3EuMLSAWSJ2UC/2CzyhV+HLjke49fTLDOXzT8JzqK+5jKsrMK2CIyiXMCZyN+Q
900d73M//sljfQtLNw3Nxz2B10DuBmLDnjEzxPrIgeSHfxcHd+2gxe4oBYxuUBeyeNXUXuVg75kD
ksWPP7R1tY2uSBn4ptZkz9t2sp11WOi6yd6QmyVc685++xfCheThrWH9IKbUFxf1sn1d4tM+0iC/
dkq2NahQv+Fp40jT6JHTaClZULq88Bv9gX4seWuW+tt796DsbkByLKfgkC393FCRAsCUTHnMEsJA
ErKzmpMZMsHToqMI/+YtdHaLlcNsgPY4RLAHYVlRMwbMwqT9WD3cmQSoD/O6Gr5FR9nwzvRUeAyP
5JOVwgl540Q88z7lfTs/qknM+RltQuRu3Bzr9Z2DYD+2XcCka16akKM/3VCJj/kF0srBF9+nRex1
T+1GJ0GOm/m8WOoXZZARW7OHlqlCAavxY/UXZoJQx+92PLLf0YvbjlOssDkm+EpHeblRTmQ2HL12
h48nY9cSEyvR5hEDz0imNV6A0GwT452zVw2mJBO3msTawD4kIA+m9B6KsnikfvZbqWxeYnNYKCJi
YVf9FcfnxiaPJGeyrR8Vegwaqx1fr3gCfYRQvJ83aY4K4T4uUro6wANTnHgl4Eoyk26LLhRQDGnD
IZyT1HDzkv+5tf6oYo+9NoUyBjIjUvvUrBYIa5TqxZ6/zlrb7M9ZThhOr90mSd2MdiBGg5P5P52s
nTqLzWFYWnIBN8L470zqcwMm6JBuDgblIGbx+P2SNgL0338QJoAjt5TCAcdj/4u7zjSAIaUQFuQG
HV5O/2b8/qXs/G/bEOf3IaI71itV+B79kcNLnzd2vuapcQtzz5PfZBC5G0tzhfB8PkPFquFh7jit
S4Ec4xajx+i2rGpMnIkQ/63v/gGafE3wiynaFjliiHQZuIYV4a0DdW0CQbxoaDwYL/6n1XTaBCJx
6dQnBHsMRRsODzkt5bnsjaC7vQTYi0J1FIOpZndBsRiGossXK/m7l5YUGoZpwUQ/UHPVYqpINrU8
sZumrFAW3pl/Sds7lX0hYvwqOGOlgp4rODlm48hdfTiYDCDhDggxi4OtcA8/RHMqR4mxRoj8jsZ8
v3A7IsYUCulGwFAG3+yEbOFB4Bk5Yz91aKGjDsmL8876k3coKr/0wfmuP7ZKaqNwRKdiq+90zKsv
YjAPBKlKoilNKZS4y0drc4TtHUfDrhQHWGlq8JVHhq0IAmWAtlv4bgCHzYbDpuFFp5evUV3sH5SE
G17s82BHT0e+nKD+oKCmh7uSo+rZ1tvEbf1eBkPkeERl0A1JuO0zCBSJY2486oguy6dAqCHJP/j3
cDZEtYDbjiOW7UtlLwf6ZOm53CmwTA1vCbPJS9FS4FV1NKn7mcBNC42AcOFg8YuASt5aHqdrX9F8
g+alsEaZS+vFQyDbodrlnc07Pf2KZjD1hn7GyYUbBo9XN+DjCtGabZPmO1TNv+33wNkm6VGL8DPO
C2JV0MaKXwttZhzULNVCev/I/e/0YokC+eLDVjgCGlsGkbDSL5sOcycj3TGihKZ6RlScg5ST8qnQ
3eBV+z5VBeoKF1m/sJoJSGEIi6ePDkrxJTJr8IfJGLab40ol1sSre5mqCJDfoKjYwOvX1PXqoebP
9rPexFblka8+VJmkb1Nt4TNFR88VupZp+zQOqBlkOyQb5ewXgM5a1up8S4Q4pbXfaqmeLKh76sNP
EyWENmy6Q4BPyiA+xWAriVoDltgAKC8bHX7SYbJ/0FacK7CZt3IHagzMcVZm5O3P5/fT6jabQ10V
g1H6u6jczS/uPtkk8/euXmnHtbzt/uq1dqPMqKX2l8UItLfIr46IJj1PPwtjzTjGBLbeLed9TLKF
nowucb0HU3hVSQWMJT0RDvWPtazglR6OK+LCwIXB7zj4QMve6wc6ZvShAV0tDfhPRfm8AF+/snxy
p80Xd49CpG/tjw+qx5VhJnHL6l8tgO+iAPWyrS+HptZ29FioBsTEt1z3ydbJ/K/oYxX1u8PpVw+D
68HIOIoDOG+/1D0TzDo91DYrpkNhoYLTdzT8v8bfldEmXprjOdeT+Px5LsYvR2g5Nv8mlUFxaFnY
fjgBo2JwcMpldnp2JbhwOcnghmsxw0EVa/BQ9whb6NC9uMH6mWN60AbkeIGQeNEz72gA4Md7cdhW
L97CF9fssCseHQxGgjE9RKC0hGL0zRgHZzMGoV2TPsRStfYVxKZlwWRx/baU31GIn1aPJtI93L+a
J8D7ZmB6q0uAtBr7ea+lyxfB9QF9V03sjFYLdRWHCluNHMk7p3hBj5zUxsoHu2UtZ0enxTYiKnSy
z/L5/r62ivq5aWNEMWN6YsCS8yOw2y8Nu+X9WnWAieJjgFEMm1ocdLOYb42mvoZsNbDGARlHE2IP
p/8kt5oOonDlaisFrLdhsikAo1NZmvM5kowRh6Z21hXhSZoUPfdrx5fsJVEIy1dhw6dkTWHxWki3
T2qy5//n2fhcwip8gBNW9axmVl502CEUys0DZ1xSn3oionlrNpNWiMUSEvLSVc1pnWdhHHmbDMwA
bTifc1bMc3py5lEavlcSH/H9iWUlSFkNOYm5UT34KPdBEuiHADAFUMyaJUAUii8fSzV4Fp4qzbF5
JWbgIZXKa3ObSOa1FFovOJRlXicPbzZ0Naq42SgHSGS9jEeEftAM7rFP2JJSmmdFw+t+51ANDU4D
wDJx0qXThVzolTN+u/aaoaAaB9FtHRi5RwQLxcScHZFzLQNKDL9+BkiF2Dn8dkHFRe8vY6XrEC8V
KANUP/6gTNq/GmW8h7lLjRFYcFivXame28fM/9IrFoe82Ch/YHTKZ3og3/CJ2ik/T7eBCI1ClCNw
WmniB2NUvEJt3CV1Gsga4Ibnr9MX2bM6HHJUxCRm5RJMD5EJmJqAl/m9xTD782L65qko3yRwtFsP
HvMqiNr15MKpUwFJSAMGFzJN/Z/xEqYkUw5EgryXGA576k7Vomrqbwj20qRF9HbR52EQnn3W6fFa
G4bNEHYjBWAEHX2nLFPwCmxHwTwn/aqo0WuzpWjRDCiqkvXJ0bv07HO6UC3J95XtXA6q/UUFbh+j
79aOXLQzdLpGWkC0Pr3JrvVVjEh9yNtsJNVbeGA1kPChltNCDFDg5AxjG1FGAegy6KMtbSLlidmt
6q5Blm/D0RXDTeslwVzBTAC4dRGqf/ZlAXA09+1TQz8yxHOzHEN+Dldiyw4JcRo0PWUOckiuLsGp
UdKVxGUST8ZmZK0TkcO8mwbaNJ4oRiI8K2/c7ZGb3/ksw0V+KpJFSFjRlocx4Kvha+72y2tHIrHI
g14kdE2wZfc07jfdbg5uSrxjVa2n/zIPC1QViQu4Vw1Ay1+rgZcEPvkcUygoJT8kB4E+EzG+sqgU
C+InyQiUpVxmCBrj8WNOu2FSualJ7JAZBAIrrXRmgbf8vi+Yocpes+5LUHKmaohDbxLpcbFSsM58
lxU5qOL1HCCJlNxRpqyTPv7OEolg3yphS6tlpcINz95BzW3AN5cQAFP2dr57dw5I6hVqUUo+r3Xi
r5g0ayifm3cAbLzjzzyDit7G0YhTGN/l/AEwjl/KxejU3Rpfqr6rjRpiyiJyV8EPN+K2QUqblsoP
nic81loj8/bOyyNSRyABQQD45vdpRTFSnClfJtDSUBFDfqc37/US+Fos/ZN92rGvC/8j9ZNfkWLx
wRKimH5dcIImHmS/PkmSE+3qqdxCAc3o05NlHGTqsRfluFUOCp93xKBJm8vhnwjpRNrzz/LbUtul
HRuWA9TmBDcdABjflL3PyiuJu7PkJRDugm+i/09D0VdBcyQ2E9JAE1ZlYdiypafhqX5oDycdaJMA
Ysdx16iZeB0wX97PbB/oTWKkmpVrdYZqRFlroUhmoY1ZFLlawTiaKRnjoAFdxMe6QLrDUoq1TbIs
lIKtSnbAezULZphXr+MQkidHrZjFo7gkeAbLdzq5h8NH9gBI6ydWoRD4VpghTLcg89C8PsqBfmjo
lMx0vv13q5e+umFO1/sEztRbKmsC5fdkk+Yy32PwQ9XRejXEXk93pkqq0ah7iMPx6ZoqrIjOz7P+
p+/BfiWhHLpgETMkJFpyfrxwiCpLaDGV+VEHNDmVpk2FQ8Jo+0bLHO9jyxfx25V+V50LzwiUIoc4
R06ZmYoPRSpiSE8q7XfyDv46RRmSnm3eHcofLGck+IfwEatsypl7N18rSSBP45ZS6rJGU4Nmpwfw
yGjSdLYvVo9Pf2zSfkMIFxB32/CZNTkypLCaTMJlRQzCLgeavTPO0HjyokzhG/bnUpV3PyBzq+Ph
xOFc4FIJxZs9YFNG0Tzd3eR/EZBU7ouAYXqbEGpqc2RV+ZzvwQyF42+BmkP1ML+gfVxTQoeVSk2Q
L0ll/ahdpfkcTDkPCJBXb5JwqJk0a+PaWCXMGrhWknChZU2fxHCFPNODUy3rNc/GHOHluTnLHvVf
S+/mgtIygP321UQPuqSPWWiNoajjKd5w7KtQWpdHB6nfoRfCYFFYmR327xFUwWouuCGJ9oEzResu
LHeC12AiR+lyPfzMVBe+oDQwSXI0eeDSuOncypkb/ahExpIwI4msb3D7uO3iJ87idgx343OOS+DJ
GPoSHUuo1yEmKpADnylxXu00P3vxi48vloZCOFnv5RXbybCIszilc7zJ01BvrurD0GDObopk4Z1T
7jD8eFiPbZAbky4xFPQz9HwneHo2wH0m7eDb52KsgwQPL8C/NeIwLgzNYYWBmgLg52/bAhZsiF/g
Dp4Y6YklN3/S8BEG1m7qqVl1wkBgNirw4/g1//GCmPV94FygHZmktOTgdMT7C37/pmqXvEEECzEc
3QUSwhx31zwcTPSyZc0U/spb7mQljgDMqzBIrhpUKMUZsOq5PPEozATZH7e2sZDNpoBQ+kHIXUkl
hNPt0ux2bZT8L379gey3h11+JuCOI1KXJK4xx5DVechw9/rgq1NtETgyDn60UVdSDU222+PJXRRs
N+v/iOuhSUfujGiNPeNjEgW51z8ASYvO4bf0LzD2p7c6UK24vW9xlJ2p0dZSwd8+A1PeHW1lpmno
PKsY5GmDbme7v84TJoZdLafxa6yYiKkTO9bACUNf1CYutu0pRqca4/STuJzYuU3rGTRDC1Q7Fvpw
oFuEl+N0wBRD8iNoGDg4/Vs5/H9y+4tPT/SgWNd4Wqu7DnZ6AXf/VTNcGQvjOzD/KrPGZP+3PuIv
oiuhMxs3MpdcQpMsAvY/hwzWcp8a4F66ATPUybmZ9aJ/KGkaHqdPfFqrgcwePW6l6um2qE3WJFVn
Xv4VVCwt5MTY5tDJUTrVZCZzwhTB/Ul9mYyipGFOxhmzCL5eKRh0zSnSEKFCdZp6Nsql6mQkP+UL
W7uKva3Vy5WlAtfJsGouzcSKrGsE9YeOVX07CJQVSsb1wn9iX/NAOPv3pa+O5BetBgoGBquTuZNl
5qA/MSn6O5ey3o2JHjKriffVKGKxZit3K6IA3151ahXD6zouvOnJpyjqhS9RyR9zqH8So1wnY8N7
gCoVTIc+j1Ftnh4NJqps3bPm0WhRr+Sok0vo+adM9D+ZNxQc8WbdXIHRa87MVidOzOcJuBWxIcTI
Vff37OOVajlCYPNxaZJmVNkpQOvbU3L+JszUkQIJuZpN6kB0GaXzNhkZUdAlR3C1V5p2Y0jlG1kB
ELYQM912gKNMwh++GdQpsArm1NIVvSvAAOJga6+qzCKeIfolSpdoD3FV2SKQAqV6N/cVE8EBkNh9
MnSXXOVRSFlhEQk4zQD32j9XBuzacfHbXCrOPXUeDgOfrepr0ucUKfEiqFloezRs/iickbBHK/O9
RRY9EvZ5uhjFDyale2ixkeEX0QWTZ/cYOUBiE7BsjPQfSZ+CsrTC+hMXF0RIrYe8MY3LzHtDrYsI
KI5Ow1W3oK5sv88gTwN2fxySHm6w0hcGJe7DAdCPY1CNaYjzpviqh9Js0uL8fbTV+V7+dMPmlGFX
a3pRDjh+ri2Td89XJeAbyP81gNd68MPb3zmM5YWbUFJUKlBEHswEb0k1yVi+NuffnJdYbPBAUiHq
BTHlv3MD2WRA0+9Eep2VLY2csuxfi+kurD2pp7C+1MxMR8IQxcbGlOYDtIMqyK0yneX+bNOInfwX
H0cmi7GbjiH9ng7mA/rSnM4QdJ4s2QIJd119WL7TlRHWa049156cQqlyV9qqyovSU/WFqx2kzI7d
WbIRd6PLzpZEEF8/A6pVBb0+25NXpIYsepCbW02+r/9NqLvnnJtCPo5NahLZ6tuo9qHMeyKTRnTn
Q/p4QU4xRlpcq9SBACe3VJ/LNRr0HlQWBOcFFtWWUiVL69vPRH6HFzzVJSIDAQ5Qy7kCXV2XvrnQ
ek4YyIBDobSgUUymp/rwY59QC79q6gcfqb4WC2dz9yZ/iigDr8VjjiPVvH1gkx6bpNpPTggmQDCE
L3Ez7VOBU7jOzp4nQVXcePpH1ZmIIQPOsSNU5XBfPnFkRR1XUW4GRG6QXyrH5hUP9qwlU2AOpjmX
SfOhagExTRr8Dm6dvwp39rzzmEClz6Wv3ho4TR40TB+0Ii+0E+pt0rxQE3xz40ycRfcYyv2OrncW
XJ2Dbl6W070l7PI3JOSV7D/L4O5264YJ48zkw/lu3JO5h0Zo4BhjA7xt9Gg1kCQcapxV67TsmC4a
W+jjLU6vL3VBU7Xa0NDuP7GBtgXQkEU3Mt15rSo8UNWVTGBAJstTkf4AcLAH1NZuFc3mip3yNkYX
0zcr5CafZaOkm4hByAGwhz3baMklQqt0+MKD/zOAiAz/VB9SIjUClEuxH+xAj/+DXzkDiGxN31HS
ZDWUJsqosRTGcOkyuwWVS/SDaIpItdUKVCay+uDreLkZlXDaA4mM+sahrh/aW5XqUvHVj6Ss/NmQ
n8fIfjdrza1YDNzTpuntvZXStDQSonJ0qgbYsPO5bzPV/yESomcq/KzR9ee8Z1Q0/vMCxGadlrc3
7D49URO3VDyWrh8boojW6XjQO3oW652vS6i47dR79kmJ5XU5CuxHsrAlTuxAY7Pv4CnFVpPsjCJX
vqcVTj8Ch4drlzSJS1tb5OyWshDVqCqTJWeKpW6SUH7nthJEF+ovxF8QLqh6dlIB8uoLoyo6dgur
LMkEi0NvEPgvOyr+XYPEI2KNczIGdjrQpEOIyN0G9vPh/BqAgXHQo0q9GIBX3C+ijlAdk6jn6JBX
6rJqsDiONF7zoGZ5ll12z2xp1AqfeoQXUeuBWdZHoTjyNADgmf5mODsxrPZcLzE/67E+2iOG4d3G
S2teW59yV6EtAmKvV5dLDc8yO6zqFSSJKAQNNtxHbFCwFXcq1vZP1pkeAejq3SENO03TMJLChyRm
L+BjYYaN+cXcI7OXjy1WvkB0Nw89osDubHKUA02tbQvcwtHT1PViI1qKlaNqczEvZbC70TRJRheM
BdF8iZ7OZSzgzGiBUZxvfuXuxJEabs9xC8uhPEboXxP1De0XymQu+FFFxXqXWL+axdbCZ4UWbQu6
M7b/7LpCPQmZaUOEPhggtly8WHJ9ZRQyKMK0pAAizrNr+YUbZsexkacUraxQYUYu6z1HS2Jh4OtV
nyi8667ykO4j5+ihxIDCGRY+benTqIW9QjbD0GuS73/smXCwiEiL8B3DEwG/Tmevg1egf71IKoJg
WCCBzRTxvlxiG6CDM3/QTE0RGfXRbe4TUTJJYO7YGT1TwEypFMitClw2KtNRIA7UaptKFcrB0dUT
wcIwRbgm7fEZFd7eMMZ5POxQwp4ramMYwRTtBbnloN7VfwHhlwlyLK6k7CB+5VMLob4JcUe1Q5ot
WfNKhWnXjzqvMPiRE+5Zv2hUzaeBolmj5dqGwHq1+bUv4xRZf6TOBm4k1cHd19Hg/O4fFeb+tlCl
QoD5aLXWNhzq6pCVEdlaV0QjUBgJVGcLWGQe3JjTnnTlA2CqS+O6JkZQhDfXZS1L33JoJbAEtjC/
89tCXqbTDI5xcdJwUopxXzdRdEpiJMfOQuruDKXkjWBH+imbcHYHX0ShLAxRG+W/PLJdxyKPezc9
BAX4G6zlPg61m7bLS4fHgQvTAlyBZntodL2FALNTLSF3B7qeoSCunQWRAeSXjnDMbVBNF6M/SgjF
DqM/jpfa7jtFzScTQhhbJ+RG9NflC9HITbur22SV78EH6YeFwkUT8KZf+4ulPuadFVpiDMExm5SX
h+uQt/urZLHs9vSrFWVf89jZIzSYnDCcuwtszzFrWoB22VoUbk7hdvA/CWWpkmJbMNtR9UiPVf8r
c1+gR7n/jiD/UgiklBwlJsd5IvdXPcFUuViOZIjuCm8I/gZECRc4zq8rG2Q6PUGlJnAXPumPkvaM
5T7Tr4379yTE50Jbqku3uJ/sU/CdOlwlpkfXC69wuRCmmLxtGXW0Axaxf2/SJR9rF/VJ5I4J8D1a
HBfiTV+MLrqGQuVFXsOAUO67st+1mWHQxg7mjS/QxopSFy7M2U4BMTfap4Vrt/3L2+egzi2U0rBg
VOE2+e9v2yrdtU0sKyRaw8HK3im33GUsiAdWC77gXGzH0K52QwzIp2mdF6ggNObt2hprOzXpbVzs
EZq8ekVpK6KL6k26u/x4KjU4dmBv4a+mE6yLNeDX/GiBIKT7c6y5eOmWqG5xVkCv2464JzsKe0gY
qITt3jqtnJzS7FuJxqfC2uUHByzOEOtB8dlFfgAZes1XEBIVfkQyhpItNjQRGUYg2/hvNCmoa1/U
P0qMgA50/DCNsG9scTdCK5Aw4dwFiPH+aXineM7qx4FORQWnG/u/Inf8qtG+uhTH/8yNkXBNMpig
pDKBui98TQadtdMFJFaIQc3qZecDyw3jyPtfMgPBWr+eFgXwc/QsEKTAGzsEaIbVi3eHuS/A+QOY
5X8Gng3LVkPuEW3+9+FbzxUH5cTNWHHcmunUTg/mzOauj4x694+wq+OB4raFHHWrEhovfaThZc/4
4M2URJSs2JCQBd9NQ9gt1GyXSP4BZQHTQrZJKJkmxDdFPbluppdqXFxsMdcLrn3vJsYDGLW2LgDw
/VrLPqkF/JCFQbf49kIGRk7K0YbUYPJe3myie/XuFQFLMKSLuZns2uF4nxox3SzWpA3pxp5qhDb8
QzCgqLURlcPegjz18qzU50TfowQC5eetTexCazOil7m+lvm8pPbftnnOU7CHjwY7UIXQAjAY7ZXx
mwSc5KYqxigqfE28Hc3a1RADHJu6JQHcRD4LrFraTjf2pMCMt0aOSEbxyRD6NwG104Iwj2B3f/ky
8+gAK9oFX+kZ3GJbCg+GzIqM/yyNj/EV4vLp3FC/Fovj9iSLzzARJisMzduKAIr1LGst29PtFJrb
Ka9JN3Ot34raX6WIFIkHH+/AgLDftDMxKJkRsVUVTw9cJUAUeRiwKD+CAwBMmZrSS2nFimDuCELK
iHOMLTOPg7yw6fK754nd5zT/pWbC6+IXbwiV8U+y8aVwK+KHBkf9+Flno5LpSfrVCJvDvFKq+ypY
ygrF/ek/jSBkq+HZgfYV44a9OXuadQd6IBjAXTYtJJ7unmwWzeIwB7zragHUFFnHUXVQpGegJleq
/Y+uKMDoDPpwTOZYZ/fEQtPCkO8mEfgsWLQoUCJTk/hLq6CZymAAElm4BrzfZeEyDR5vRCLvWMhu
1vOy934+nmSMVW7PHLmtuluDBUubt71vc1ERg8LFCFbPd2mDTx4n3cphLgDHWWeUoTpVeCj5lEka
RZkSzfeqcDIAEe5d9rARBUg1ZzV7sQxqOSuQ4YTnH4ay+nOewfzUahs15OZkHDo1nCXeGlWbJc21
P+LTGS7XUEhBapIHOH4RkJfjsXv82qqJnsIthLgF5LAciWX0pIQju48Hs6jWn8pX7XOIovGwauWu
lVWcQEl8TuIMc8QmDMlIixZxUZibm+dVcoaS+DJjUEs3h2rV9HEQhdjWwEE+MJAvMWkU4y5lmlEC
+DiF+PR8GSsXsAuw5FIutwl1IYdO6S0+PdPbnsn4mIP41FfHxNQBJGHE21RmZP7Y+ykRXftOG+VE
jRHi1Nrf+yCfLgEdvOKRvISRAZOK4nGBXPldp/YsV6jl08QJzTHL1RUl95PpcCkxO8fxxS9845bI
Ni/yQPTq49OpmBJb0KKve+SNcm2YopKIPGxmsRe3epkqes2dAdixokpWnlGal0dTK8ufOC/wB9YI
MvlGs/15clGmevma7TYQIfaNaNbWiAyKtRXezJBpBnp8GO1wnbNecvx5Sr7Le54OuGR/g5bN68Wt
axOpkICErcEKaiDRF4PlpZHGPPVaEHqDm0gaj+onipiTXGF/NuVM2QR9qaqImFlJuK8HY1Jhvdeo
NrDJ7qNU0foStP2cC5VVb0aDwtRDQIGlM+qHcnADQM4NTDK8+toZx2YvdqJzdPUgwa1S3VxO8Rrv
x9R3VvTIvattzEPhUKrdVuN17xWK34ghYDnlk/XfYGJjkbMJhbjJS5ohaAIGC7o6LC2WUf73XM6n
5eA/sWut03p78VdmJ0N4Ma1MIPoIsQeMuVtJgAuqjqat+S+jBdGHZpee8P6rX55NPDuXvX/DXrJ1
x1sdGT+egx9KQL3pFtUXfHHNGGrfOd9jPRr1PoZ9tqq2t29sBRHYDJztOQaBVdiL7xxh40Az3itw
U3XuG91eWLes8dw7KqtH0ZB2bk9Gk8iVC3pKeZWJ9JKZKzZ4lF6EbNuXhkOeav9940DdAZl0tdln
YHzWnZ6pCQ7Auiymn0NmLumGzzl/TYfXTvk1erY57B0y7rJI65Ij6BxKdGvvpE4xxdyZREDOxGYT
N7NfvY/CiUOCj0LoN5ip5tV2idqbCRkLBsZ45zk2KNCOnq2M+bX+J+zfX1TZIKIXtMlCWkPZx1d9
oI6xLw02xDmMKohJCaIPuQ4o5pXJ6F76gp7IzdInCPQND+KDTEKa2Y8IsTM22bvsUK6a7bkPz+1s
61aG+FacNblriSZNE2zcAe1dgnK/FzlS4ZiAd0jkXTj1lkr+WIIbBB4/bdi9t11Gw0lXP0xABmNH
HNEEcT62hQud1HKFEhWhrcq3ryA3IcHV7783q+DEzZqTligk4vDRrFGuO195h+GP1w5y1l9Dde9/
hpK6LsEwwrebmQC4JMSUVH2QjY122LtF8cEJJs3sBv2MdbRUU1v4y/wGBTViCffi/ulB3QCi3ADY
9H3hZmMDzYQ12W184smtlfqvM8+JAN5ZF4uGsG12Wol5O7zHcYEKNlZmstUwg/DMVhQ94IlMdLFz
4ru2lyWsdHd9idLT6P1vsUNa2kjMq/f6mA8MLauFzEehVvW/6GxpfyWd8w5Jwor9HYodwEiJ0UQ2
sjRO4yayx+U1a9X6e/wlj38P1C6Cf6Hj6BZXVCLaz9kukL5urcxQJgaipS+oV8bIV5Dk2SFG5c22
rhmZiDZIev2T0NAFx6HiUSZyaYonCIP6Uc5k/TnU34LeWPXHoaZ1AwvyhmazXqDmS8Ddn8c4I19B
sFEANmcqfPmzPIUViNA/2vJFS6I4px+otoD0KnEKWlIagl30inOXovVGZIUBoIiC0T39XcxVb/A8
ppk2AnNHx3Lv4ovkAP6PoKR/jD1/GcIdJU/cu25CFY+1xGFJvl5dPLj1CRxjqoJ5+28818KV492o
esFLQdHZstithbgf6Zm52dD9bDxWaFHXm2occ2oW90G8RAgBVe7ITuZ6wLERDROH/+NTfWH2JNfH
TEZyGni7iwPNBAaaDtUGVym70jGkaP//JBsXjTP0F9Edn42nUhCTy6SRA5dEFQxYV31aGirE0zCm
7XT95IXXxGXUpX521ycp++utqI36Mrlh6/9jegDMtIaiytkqBOzGuVz8DSVzdn2M8vcav2xid8PC
VbfArHpTZC1vhnG+9ADpynewETkM4/0kTv165RcQp+yde5X2JJ/e+bb4koCVOnZxJL4BLRxQvDjm
CaQOzTLAQcSvIxhPWKyGfXpd99ns2jsYN6Ecog71Uaj7ByxvFpsL6vDV6WNmG7znEQu3ZNNUUSK3
OakPu7cfIhltRPJDwBjqudIYQGzZI0FJm0OG9EHIujt1i+8wkjNY5oNCLOimgGURhCUkTxaIbhVo
fLpVDSMxP28cuzR1Kf1+Ff2065gqvzVesmZwmCExJLmGQAyWA8us7hYXwicri844aOLzw7630MoZ
zlVZJuLRpwZP/Xf4qCrLsoRT73Oklt8/0jqyLWGPbGEtN5YsqG3gD9e6zgxeGgf2K2cfDHaM11Ch
ZPPgIBzXXxNMASLd/V4qpwWtcKYeDhbRFQmCo1lnDJqtLbytQQMGltx9MhF9vS6cGV83Wf22Tmvd
Y7Rq2HwH+CkxYDBx8U5PQepoz0z0W81f6W52Ldm3GRKDuIkUKElKCBhBYWWu2h7kwA3eADKHJVWv
M3a32CYSWxET1WaPDbCSlBiZbsm6kwe8O1NSHqU/5/DgkjpJDZhVxUr9xvwPqtZ+vAxDgCP2w2BI
aTzeApi5a20luDCrWMKTK85O8EDEdLzqTjfVf62qRs5Q/KJqqMxGCbgurnVzCsiE+kjP/ypfa0CY
GxpawOA9rCOTcTvAmGrbNx5fj0vqqbunfwBPTLet+ZhpPiMMlbRHliGuuK/W4nxGEfIQlfK7eCav
faSCYXghmP974Kc2V+uE8QvmKqzVibIOAODJaEQfaC/hzzu/iJB7rycaOWMg21Ahtd4imc5siefM
yY6PMznYIPQIlZk1yM7zKWkBOdyV+R79XHJguaRDVlbTvCs3HSbHlR2hFx6ysaRvevMLyW59JlzW
ZYRyVg+htgRv74ELKMl7yRmm56JcgHAYNEIUpC75EaWh6dZ2mBTPbP5SXdmiOZ2C6D4o94riwghC
Z3EUXv9Aompvsw4DThjnttNIyB2GzvC62RDpFcL+91MsMrBVZDqZr2O2m2B3fPqSrqQqLJxqgU3z
knRf9C29hxhFYSubfcMaMIc6BeYysvdn/213MsQ1HgZCg1kQl3i7DVDFkXY8czhg0l63T5cW/e6d
vqHEYOkxfO4S8SrcAwOlWPgC1ftFDrWOVdtw3tMTjCYeiXKv/fiwBeNo+8zBY2wiIErhKZd9fH97
+52qnGRr6t5xtGFa34OgFcHAsM1mHJBSJk3qzfCKYZxu+Iw+Fsw1toMPR9ekauiWlmPPBF0hYA4P
qigRvaCy0QHlb6iCywvZ9tyCIHeyi0KOuqGMVb6jhw29QNz8Ffvcluvqf4C5AmYltkelo2N7TSrP
OdVsoEOKM0lmP+otEgVHjJkf5e+LFBnqHk+tVlG+HvIzIcryMqwxrKcRyvY8uH+ZcwTKLeFeG0iz
ww7QZjD/3sNS3boNZDj+QVR1A7fKpIeyGNZhcavU43YM2m22Yi3YyBnFzfCXJ7VXZWcQF+2pHEv+
Gv+ijuFxQElCQ1lZlkhQYHkfuplvc+hyDSzOZEySzC/AA/cZr98TCxA7YI/MeW5hVIgZsan7VM+U
TVGTo6/I7kO5mRanpuxqJ/72HNU1unj0p2L/GgUAaTKHhxuY+zmHPTRpGUglCfKmEZT5xeuoUCaE
w3PN/mJzScSKY1UvJDSCsTS2avIlmuPhEisSRdFF1septEFDgj64Tnz93zSxcIXvfVLFaodDtyhP
ZBrokDscDBuJpk6bEfhickyTrimMJFcCUOvCGyTcZElpKu6uerX5eOb+tPAH+RKNSG6SiKw54TPm
K3rV8ltq1CFSZJOQQsgq/fSn8nXe6Y9HzD4RzzYPfCOTG+D5TwAmriqj3c4BiVq3BJlZk6vwSSX5
A5QfyZRWgoeigAcdW/cMv4IEL5eXcdXaXOQRttRc/cDW86fsONpIUH40aWMRSfxC5XYFJRZB2KrX
6ZTutmht46mAML+6BBROdHYWAd2dNA2XH8Q79latHGhRLQWn9IppuNVCJ6qd1aFsc5M33wyUI4v8
yEvI04+nHpCwYV2czZKePxBrfHo2ULGPzj5mKQLYd+JNZZHHDbwTZk6nuGislOXLcTIuW700p+Oi
eJdW+HD3rxjrhz/oeiML6Rj7pP261jM3cu9qY8OwF7+2AoksSKSJG1GHXWGrK9im1jfO7owA09PD
dn3JijFlmQK+D0y2Z/wGdajDhqd6ecFcACTFbx4v3XWZurn/y15VrA++nwWv17qMDofMjmPK2svC
GOdl4P5tNDcok9CDHKnTkwSJFCTkRaXwdSX2Xid8y/L8HoKTBiPMznTs5Ro5RGBYjyTGwDDfc858
kF5rRzfzngMp0/4HigEa7NkPxzRd4HnNXHDAPvIZ4PzaL760aDX2IBR989vA3ugIvPDDGfEAde1b
WxDJ5Jgccmkm2LzdsH6HW+AMIFl+6hwTCZNKSwr/8af60YYdTFzNwqxXNtCpGG778lLcfFuTYZXI
CrWJD2rL2Ibj/WLcPeUqiIbql/E3/11EN02z5plB3M2ya78PVzuODsRQhI5usLtzDgJ2Rln/u1Z2
qUrWs2KR/w4jflHC4DNEGDoM9HodVXR4cRyZmsPw+sE0fOJuuTN6MPN4IkrUqnoChzQfGDThq0qI
fS0Vr0i7sdTLE6vZp5v1z09FOg/eLw1cENRffM0CYmScjM+/EETA2GQzLYabeBa7ZeiczdnVzGHj
+5ON25k2XRRtrKkQ4nZnrDonmaL0gtXtBkRPBgGl90C/jvN8YV02u1g+s++v5jnW+Z10qTrIJ1dc
+Y562JGZxwpz4HOVubtYMYMt4rD+rQIT7KUnP59nr28+8F+UYZgeFEn/uESFPXaXMVYzZnUIywAl
q+D/RO0tn6F2xgDa7U3pWIV/33l5kXcve1XeRH+lbbimwVSkhdycTTFhRS0IepzIjUJzhggPH/Sj
LGLJlI9MBjY9X5QWMdUVxy3DaXuQdQnh+Y69dRY7nZLRnW6u5GXB1wmpOExBbD6wT4D8IbrW9dpv
fZhmIRXIzs3uXpyooTptnsbwheMcFQ+KlV6Z4K1oGY7ZBa1SmyQuLZn5y41qJOoSyp2XRRFnYfJF
9bJ+2VkHf+XGoZlPDFutAu8iSP0VfyVcek/OC/w0fWDJH9ogVCJl599tt7B/FpjsZngSfcf8h64Z
Blbk8nzpRu0cMRwzIxeSzeM0btuvpVNg1bLsUW1S6UXo3MZI2oWlnWRTwLrTBnl1Yev+JT2lpQEI
SS6mlDKjmbPAczdPNa6I7t3nfvIDQf3+nEyQ+uyX84kV+SJRq4Kcy8CG2bca2xuLV5TUfzhANMlY
K+8ExDGd4ub47Kj80DjulHb5iTlnAYPPPmycjEZJTfvvlB5uCgllZ52usVYuR95wWk2239H61Amg
s4i1iK9DE0ePmpWz2LCen3w9C9sS5OFEyAescNCyVWzsIHWWwbdctuDIRyKlpzobHclso27pcbAe
7GTf90Iogg8ZfPwICy3NONH4II4bAhuU2krXbHxSC8Umfxb6KpGySEHcTilihKxzYUAwqGjlPwHM
9RmBhZHucK99MN0MkJ679Kl3YwICNFMhofGdyjunndhHu7yw1oWJOtfbwE9Bnr5p7Z9tphnq28LM
rJ1L25sg5aARzvUOT8FM1xzqfiIHDzYlpAKRJ6Kw6JoumTJTshVRgfkrEF9NcwyFSI/cOSN7+Gn0
6u1R2rknSnsaOusHceHmrbUFzAyYseBTS+KS2ByN2WvMsM5+KukrjdHda7/rDIh42EbRPdmu9tlj
8AcjCqSKrKWrWfdkNarnjexWkA/v7Q8HFvyIcmftWFpFyrPuRmTmciw1bT91zhaS9LnfPxCTLdhh
vHYDe/ZsqW/5vA2kDJ99exOWRaWerpr4fNWENBjvJJfwU5UkAO8MsoIASdkdtPyQ6YNqKjJ/1HN+
GCLhJjennj1skL8XVq80w88tjPx6JwcsJEj4qiWyhHoDd+TMLAItFYfvWoT07UOHovsl6V3H/6QD
scI7W6Tp355xxJxlLiBX9JBKN+hae+jtL3oHReZcq7IwIOQPM2d0SVidG34oOcXZ98y5gq/8k/HU
RXwlq7POt0Owb+SryVKh9ikUBATMUfsY32CaOsAL9i9GahlNCi0qgkjzuQvI1u2htxclr1lsoVwS
cu/0dd8mhIXPsjiubaPTp+2K136aLe3qOwIlUJe7/xjIJRVgtmWMmTCO0A86RjEAhKiDskEck+Xn
62gLz2S24hHabn+Z2ldhaXz4/7y+LdOFQTkpy6pwkdilzT+/6ad1IzrB2C4DjbuXOth78/K3S43x
ITxMB7kYsEzasYUlfHznr7vRArUDXuewSQrv/CYKLOYjVfWA2D2r6kQ7nISN3R84n7Bb/NOsRYxu
kgtosq5TLznB1zZVZHiRlzfSzleQ6U/S9jmndWsCyqqig016Yg3sc+vWGbTxhY1DkNd368ctrjD3
vGvQhZdqiPhdZJsgrERMGIMQ2kh0Dg7Viv0rgw6djlSaGFvOEUeUSUibxSy1CDBNCTnqBCgGhlaU
sSt9q18GnTAaO4vdFXKVeIUjjLmszyCSLBia9eqqUOynq7StW6z2MECP6/aVmQl4m645gL9ddm1W
dQcZvNR1A1alrlWXIHDSbmIddaxc7kzgPCr6NNdWyIFhauMURxeSWNosY1wuvvIerx/5OfB7LJy6
YMZdEeCzdFbf5BHoJAOhF00hwvBrgcv94CBbluMTBu0i/zDiqHqY9mpeBToaxUDRYsJ1scQr7x68
L/mPMw+ntH56r98b7r36hjpGJbR4f7PlypDbX5GB1IcKiVt+RbxkTAlpi/5Y4cRl+pfe+cR1q7/u
1ukuKit5X23a5/wlZuEf/yL6IsPpnAdyIXaPClrUDCO1neDL9kqfpSQ56po8zUaThwBqli1U+dVI
JbDfH7CBzIMcO4+ta31yARW17MHvY3PeqAbBjkFUGTl/FL/gmNYPLgT8qOjUn6QnuogQ2VT7sgJU
+dc+S/Tk5XfqQDoae4b6WBHpFbaalqaL7mKjE1/Kgkypf3QKpJ9PmCtB54ezIwcKQzLKTpGP/peF
Npe3fmVQTmPtC35aFJmbsIgR+ryPQfs0YTd3tzQQi5eHSCMLoITjYZClMll7t/nRLS518Nx8+Ku3
MJ0vq3UtWjS44WjDgqz0KARnxdPaA7S1XP5dxCCEmFUpRjjLqhY7TGhAEyyZclWinZeVTo61dxCP
vuRrgQlvATIfHy6fr9hICXR4pcIWWCt3L4dzJe6tYUlJ9vTNp02oyXOGICxa1UPQ8sG1Bys/q+Gi
bRMWNyhYS3cqZaAKKDG9cf+Ek50gPgKQtLD5Koq3VZwUT2mVbk2rP8ny/Eo1adBvv6yK3DIG0YE2
3ciyetv961QuMx/W8dvoaTpvPg+L0U1JXJVaN+0yvHZQFxCIEFnnuSXTU+kxopJC+CoNjAaeYmjf
iKKS1CDEYl5uynUZvd3zXVk/oW0exyHh27SY8IzGyggb7+lq1oh+k6sE67yi61f0LOJA0QWXpsho
2GlS9Isr3Hx2N8I87NHo/sgSSgwC3apc2YJnWCcaJC9do1tCm7nq63XpvgrEjCvmatSn45CrcuCe
u4/+nf6pVlejXhFLYl5AukWywhx8inoadDZ3510uN2ChwrVwapYQ1r6dTBkOwhM843NPSTRLgyhq
daKKEHC2/BHMfn7xKnt7hMylCVz/KXgBM6RsSc8I3098UvnfAFDLbfCtJcmuAzerHSrsfJdM8Q4j
Ha1oQEwJDwem/rbmfsYJvgoN0FLmQNPXG3bjRfHZ3VQ7EVAsvDJtBE8oC7mQ8m5VgRmf7681DGbf
8XJ7+1OdJhwvZPgMqR6bD1GLLCQMq++kd7T/QxgY9U2lxX7WNhaHeItAUyZ290uVN9HfVWq0EufG
vWdgP7a/ZYeUKhf2rK6g7UAyE2NrSltBZOZPBtpBeJNIyZQCxjXOsQ/9URj+w8PLzNkLzPCZzvEu
oO4IB/0rDaK2SKru4x7Uj2vuLyXeR/hxtiVDcRiJX0cR9ndvq/eV0NIeG+8pfVJqAkVqjNECBD/u
Gd4H2Lsd78vs0nNxRvTgga9mfXloSVplITGxZmI31b/4qH/v0nNULjt10PC+Z8KnBKRfFDvWrgPR
XYMu/7Njmb2Y39Zarx83U5ttvWcvjL23iiCTV2SBn+L6BBqj7F4hYBH6NYBAF71p3+IeRpWDaMn9
FcfFWFJ0+PO56KYRR0RH+lh9cmhBW6v4QRAykoGABLpFd9yN9aFdf2zvgbk42TkdRTYYzl09EPER
NMP7wygtaX8r5mtYfWO5st/74k+l06WVBefuXRst9OcayC7cuY2rIs0dVRXcVjziWHF82kyKFBzr
U9wDbPFWOTVkwFDZ0GF21RETUt6aP9INLonlp4BYaqWyUNSaKwkqY5f4zyqtXdpW1z2CmHEjiq4l
sIR5DWXuiXx9aqEun001CVXXczYqnbgcs1NHxB2RyIE/aEFMovSILsoG0cfOCmHZu3VXX/KLYqoK
0Puqrkl8gLKrcwLwcl/Oqp3fOPdbCiD/Fjv3wgmovs8mT8a/sZSToaHr+1/HBgXYamCS+OXfRqPw
6uqwmaWirg2gfeIc6ESJkWCdYnGW2DWqvrE6Ma0q0eaYHkgYsm1I9uaS0F5KAm/GzeszNUvH7cf1
0g1ROl5VbKusAmEL4VuWBdPz5mQIpCGwWe5J8ZXZ//Acb5a/7PjPYn43IwZZXdVQCW/bN3DLaECE
aGGcfG4jo9tyIobqr2nDPv37D25MHnyM75BtkAMZVVCVIhp6J5sl21YyAx+IlyrI4Ikkf4Medilp
yTZu2ghKhWUBXMxKoeev0WAfypNQ1SpN7crzfX0QmFMp9LBW72E91VzL0M68KZre0rhm6P1RKotB
n8osMinlgkO+2m7qygrfkl/7xiMzn1MdwM+F47BjkxijMaPQudygck94nEzV55rTCqrqJNEmvQq/
3jaUi+IzUU2TOMTcH8x7+Q9Rjt048SOUPqZvnbJhye8TCCeQF4m0Jdix1O6KpKeOXhxlfxBPDK4C
sc9DHma67Cr8V5zOVlJJhaDdS6AYzUcfo92Lm0vFjm03am1DH1H3AbIRCajmcZmRxcrYFkxuFAU/
bQ/crn+nqWhOKZQGK2pEUoTkekfp0PL+8eo+YhuhMqwKhxhP7tFmy/bJM/dR9vyet6dXecNqTzLf
axBBuLKuv3sDHXK/HmOOfImFIhZnqXN6AXBiKCMoYQ/bqmzjYrZeq9+iZMONcE37ATD6y8vz11cg
azsEaFr5xIz+sYV21mjEiYlmYEBw4tkEpXta3splYIGSDL+Cqg4IRO9ta/Qr/gpjjXlRdQAO8N75
gQ/fkhecV7VhxPGEfcW+ArEvD5T51n+i8LIbGQ/vWfvLb8vLjSvutFmUFoab1ZELKdZ3NLu3fSWA
URzIzOiIcX74FXZsRa60OJG6yjeqeOXvNkV57uCQaiZAEV5MTCr4IGs2whMoXkv2Ey3dFiavTyuE
KG0KS5e9SH4HKilfjYMRqm219/VfhIyJl4nHG6/la+RxwkdCWrZeObUPvmvDu2bxNS8dxTEDaUbt
P5A6W0OzOPJIKuebVoDWSx8GrXsy+7XOinerGzsVEVzJQIXQVQANrQqh+yYP4rYokfzEowEeL7IR
cvt3iuchHc8ZQLksC9dRXN9YTe0XqNq0JeWi08ov3gvPtMB7aO0QwGTIHugdxJsxIfjA6KchwZux
5gFrZDKNzjqYIl8FDgmqkAuIDTUdiy6ya0SvxXAuFgw3OHIIWwWEmov3xWkuX79+bcHQnx/trLDd
54ovGaIwIwPfuxdBfkMVtCjeghbx033LCXmA8LzBd6sMh9fbysexK2MzspCItj7QJ2j5kzur3IpC
CUO1YB5UehsbOja1oqNKdlEd71mxBdPlBxO0uSKrPr1gwt7LV62+yj9x0UM+GW3khuK6KsMbXjyS
UV3ctQukK0vhsNpM0kNt/WSAxzn2CdnL9ddasUyEAbWVFI6hvplQu4Z+ZsMMIgBond0R2NykKsrV
bbINDpFcK31J4wabJogYFn4kXF3JaGd/rLJS0JDhRDgrBWxZjWvGBELmXFiD75r6ibDcdMAjK67c
YsnBZD2Y2kzokL4szHwrkmvV4pvZpryS0LN937EuyexFogX+mRkdr7nrajoijuURxqBF6DswxclG
Lw6i5GJBKFAGwOtH5gboLqJEMc07bJqwb2vFFZVwCWpPCagC0G8SxUqPyIO3//NjfoGvaEXIEIIP
MbNoWivUPUUQH8hfwnu0fCKILT5VfjKWyEM79PbGTKlXqU5lVbnNNWEoJJ2NLjRoUhyUltUIUz1J
1RLlrz15V+ODmOhH3nTgSWqPwijZQua3kOki4AKGz9Qx/cfITppb/D1fmFPmMBYsbHHQIYhEm7EQ
J11WEjyO2e84gyYk+8Ckn/J2QPx87JGVAtJawsmsTGeCSeBXIu7SZ9qXBPxkUEgBbjRmZPH31W49
aYklwtcYn7Hd2lOurmjxoUU47Ne9ujIsYgCKr6+B82hjltVlGESZvq9FLfGj3phOEp3q5CI0/Y4t
hl7B1keq83W7ozv18sDFMMnMBKVvtcdkHdk8TQWdcghMzBlU42gOyzGN6EKCqbfboeBjtRURYfHV
NaKJ3/s/ZV9r8LwPKE2xJ5uNlwoetsFo96TZBdhRqilNkjITvBeL1Pp2na+8ixkF6GeTVVnKANVF
4sufqBZapFh3ofZCTO2fAAKXlkepM1Y8c+ZwmxwAV/CBnkayvykzwbPeI7q7qIBrH+ccHMsSYcQJ
cOVzDglr+DO4CRGD608OpIhoxM1s1h0UIF6D5lWyXR+80TD7I+1dtIRlshvTGWsMfH1JaC3knxiT
aXXWmdPUDlfCiVe3JgfN6LGDKzgqgF2bP/A7+w2flELIYl1o2KkgvU+xwZLVtT9JJALPZ7m4SCFQ
dvVlbSNcli+VdG601yq2MqugQXRdrg37pYqpwlffiQq0F4Z/MLn6xtg7pyg0Ij/ikrM56TOcjNcX
0X8W8lA7/n5BAwc7rBxQ7UBJcQFZbqqEdrahQGAid/clwkp3enSZ0UvJwaf4IXCSS2uKugs4GOWT
jZc8cj0vWeWEDNOaFyO+EITmBCDHY4kwn2Tz+g3GPYB7OO0ThQNAfUjRlXrb0zSLxnzDDZRmGuXr
p+YcaXtKZ4hm8lotaFERPSoNyy7jcGuWmA5SpC1mwRXfkR641vmu9fTqRBlzm33t6r+YwrLnJH/X
D5T9CKMf9ISYIO585TXdDqSG81bjxX9SSpyQtvQP2z/LjyqHoyU/TqrN1h2S8RygmfBRU6p0exGz
jVppz6PwLMKzKthON9RUyVMLuHQ5waKC5OG48i8IKmvG3prt7cg9c0l8k0qYJkrNyf6KW+R1Zy64
rR2YjHvDulKk0WcFwl2DTpRvDydd3mqlro7BOcpQWVMxIeRE9iDD2E39/uU6IZkKcLQ4s/5NDYf9
9rj4zp7/i2z0cgAm/j8VIajkOrckxGe0MA8oRwrxbrafTP/etloM0yM7sSiyqBFqZXFvu4AJYIww
ugXSspicXzh4xTW0hW57ADG9BU9ZH1SonQoM7ZcZFFV6htc4A06Db2/ui3A99IpMqjSFt9n6ysFS
mrhH3B4QcHVl6i6j8Ql96uczzpdPq1Kvs+kq/mIkl47xpPZoPBoimFNngcTQcBce3vBYfsG8KTJy
KdKx0kcT0ylkWO6sxn3OqL7S1pL9IknmsnudSINLasnE3UAxBxUix7M2yEwHJRvBjRMPgwAi2Na5
fhbiYPlAnAajPI16eGO+/MjbQh/Kcdl93faaS4lg2SaeGM0bLRMhPdlNrOVVQn73+fHLkqR2foVw
B8AP34Gph0kjLjrFxXc7i6qT4UTjaqrX7GME2jWN3apZG5fdz+VuV9PbyHDv1vnojzJoK6UL7kWc
GQsvqQ9L75ztj6JkyS1r/6c/FK3YkFOv8l7G2Gr4E7c/U1QCU/HHpGZJALh+ojB/iz63UDapD24y
KWwtnoC5+YgsqbPPBLkjr5YJhM00FPfdasvh4OtJ7EVmNGtyDCcptKMPIT4HEZ0PHKmWOk2/6huX
38r2sDC97QegYAaOSNXbg3reVyiHVvl1uagzMykATm5uptsBL9V74N0sTWCDxa7qEKQ3CJmnr0Pc
ApKqmk/mQVVKd/dHb2X8OAUPkG5RXjCgTcXxlCyi+zNwqtE3DVFa82p8TxwT/zUcETOPBPUB2HCA
9STcxU4ucvJZUHDmE2L3deOVYzweJSO+jCiwHZ3jsLGA2dxUNUAcOGzgf35JOJaikhjzMD88EPqZ
Veb7FzNuOy6AmgvfPnEUo5otAzwElkRczfgqV1wb0KK8kXR8zYvniRpvqsLijWse94Tqzrn9AqpS
+9m7E+01xf0rDKf0ZUrKeUEPJeXngp10WN7a+z56JPBe2SIFdjG/0jtE2592oy3ZIjcSJvH+uHgF
dUdIfQtmnSoR8y+QRuuU+ufkTFKkTS0oKYqoKtUugx8Ic60wQnIw27Tu7nQbsDkO8JzpWTjvLT3a
VojRgW/HymH9gcL1c4sDu69ZeqN4hajaHlumJKaoybI+hct+MUSfBNswB0xtOf4Pzqqh351HNs41
y0l/HCszta8Kx1C9xs9JGnvBAJ7TGpvBQ87j/71UIlEhvZoRsYGiLGs7otslOhDAMXZOyErhrdRL
4U7xXW10m1W3PMmfERD4wp8NKTb8Q0Re+2Jk4qm8hU/7qa+p4dfwcI5zFYfk3JX/klo2aCqg5P5O
zohe7P3K9xfN/geB2PLKjWcmaLfqseLjLTPI8DaiPSJmn2IKZP29uwmz9Vn08xGqSBmXRoNpjnKd
kOGOFibhS8ts9+kz5xMoIOCqv8CXSaW+sCK4Uk+EeXzW/csaYDR2NPYfnqZV0KIivaCHBh26aC96
bGvgCxbeiarqsJ6eDVBGD0pblJchg1sNXMewBC4d2/VLEVoX2NwoZHOCjRw1ZuUMSQkKf6CJJp1K
cWzQ/OqqXhL4igV7T7tCBwkDrxJw698gjKMwHgzX3mSBrhft1vzIMTrO/hImhmQqhLAE25xQcDyz
fuz8kRlDsJFQvtqNnPsjZb6FySpOqZAH2F/ZSfqt2mcLEFKaH9LDl1jW/5tMfP2gsulKSCTA1/q0
wzgqP7VF8Yj/WjbZ77z6Ll5DI9mm/dQICPoY6ZtYcrKs76oOoVakiXAxiKXo4W0GL0Y7q4MBshGt
XJWbivzLJrTrNZMlgO+mdWjWO3LbBu+BcQOGsguVlD1hBmnDxTcWFbXHdwzLPdPB5FHHcy0Founf
1oYXYXftGPYjz9lehjmoDeZLYsrmn0NVcal0pPlXjswvjFWjq8XupYRajmCcdcGJ7UKeSit+2BFj
0pd4ct3jFQQJsikhdvp1RE6+iPBWiVwinTXdVIk1Nj9+E/4YInCdQGIBIn4g7ZXc8xiNWoFrgNUx
ERW1Wky1eFH6QYmA68Fy49KMGUwkgYTYhJbB19ru400w+wsvSOC837N0jCX3OmyWA36VeCjasNuh
oG86+2maJuTIRC6dL+jQH51iNnAPWlrGB7RwAEBlmE4cCOZQlmETSwhl9RrvaxKEOhrGZb1TWjUz
5zALx6lKfAISxj7TRAI5+hCbjnWUeUojg8SQM27fa2JM5k/WeWGjPaCnf3NGlr5sMBbNShqdXzo6
DFnv03fcpspzFY0D3DoODBaiZX38zhrdBaobTkiaOpxXGI6j7kUlHs+kAvTAZBJyR12+TkWm3egG
8myikbsvPjF2v58SQRBNNJxD0TrziaGALm5deiRJdst4uvNDmkki3nJY45l7qn8BsxhHATFxInSG
rR087L/V5wbPek70mVMs8VqGMvv1VImWMj4fNuqbQXlULJuQXgEUvTnU6fFYUmnSBiKM6A/1nST3
WdSzBU3vhMEGRE97jAW6osWRNGHonIR/Owcqwb3un36f3xIjjsdWx22JCQGKMYyksZ6+NdS8bOxk
FGdJfU0kvLzs7RavDqBcs1UJTBRyvewYdzPkY6ct4Fxfh41H25JqbdC/6pnj29z99kdegAv8TEnK
7VbC959HMEbM5tr+uic+sP8hv9zmlQwGEW1MW15FMSQghpg9qzIqcg7uMTJSx2BSAecpmGrVWVfB
ndBkfKfKRFC+zbWfnEJ4TcBO1px1PMsilavGYoS/XW61pDjvp93IvZ8lnTo02G6f/65xTUJbC6Tw
0QTkeu97OvzuuUEvdX1JkMLl33vPzgzIAcNYQVoj+DVRzgUYeUiksfahdG0XvKuVXG3BDyqCOB65
hsz5AQBDFSV/yaEYT30MZIF9rp/4KHzfDWyyQS33y1xoyVKv7OxojKEyY7N/iaTWB/EGR5nY76uA
bLGk2JY3iH+3RAZ6AD1WJSjzzjYAMSqGQb2ujtG89HLy4UXPFkmh83Zp5a2koYakVFhXVBQDDTcV
Rm4pYvB3TIxEE2i/mnfjq5MvbZCJFMV+e1wZEM/PuA9jxl8Ni+rEU0SDt4MXFFdw6bjqt5r50XWL
CSqjhkcrNIijCddVXE14svNS6Tec83ysGrxQyW9uSw5tVRjHxE/2jCw2sS4iKqaV9U7wuJo8oxr+
NRo6yiXQMXUSiGpGvBXEs5fIOq+m2tCslMX3dgIM/vxMEabtKhcEZMQMNk3/ZyV+75cGWh/F3Tkn
yBImSXR6KOekjkgf47lDJn7rEH75+lkZZygG51iW9HXeSyUN5mhfk28pGqejHZESYT7s/rgnYaqt
5hRHEMnFPRSHNtDM8GrGO8ZCeBREeDrA4ytJ5OD9RcSE2v5oZVcwDASnfHZ25leXUoPVSkBD/AAa
BtLCJbnjwUTaphdl0AsdiJKgJ9+1i1XbwA/yw+dRbrnMU6TyDsAidaSvtRe6CF6DzpJgrCOgj1Ge
89kXAVyi1s+npnY/s4LU9Ebi74ZxZYlp3jTeF7fFPj3+9MinLTee0cp6ZbUgHrqEGgKFiX9HRCUF
eSqAhDazr5ybb5eFGVEqd4HO/+/mL8l0CryIHKlNthg3Rf5U17On+PAgmnPkT2EFouT4L87ecBIp
LSV5qeoMH/Rsb3Ch
`protect end_protected
