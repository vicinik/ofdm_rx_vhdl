-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nogbwKZzL4F6tM6LB1k2HFKDIHcRyM0r6+hWeZS8mq2ZNWLYzka3ex0jAJa5c37+XOc0JlyadazT
SOYKQjZJGzkdnA3DwTl2CoBDzxZ3sTdsICj7bxqpMOC3YroMo2TzwM9CuftOnVlpsEl0e4BvTXcr
Qy86CrgqCbUJba3f6LBbLDFEHoP/nuS00UibDePC/2N+Au3wKAG67P4DDCGV0ucoIF4LePYd6v4+
y2r4LQavXYMgdaD5gEAk2FZO3Fx/d/fMOlcYDVSNBxgGAq6FQnwwis/rpuz/Tylzo+J5i8pjADUq
IBxKikuMejR33gM5NtS4nrq62ZIyNo3rIiCAQg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114400)
`protect data_block
imYOZIWP1jk6AukBS7Le/2eAz/n2HquniTyPYMZ8T0uKGt9qeCrwSvg/6n5KLvnXSHn559twXw2v
vHDFK6udSRZZ4EafPXtbhqKUYk9Q4ohvo/wPQYDOHg9/Z4YtrVQujV6pKTlo418tVDZE66klFGnL
tvz3p27gdi4l0Jjsbm9qmP+Q/Jrkp09EYsEtX0LYBfj6FVWhDTubAIDw8eKBSIqD0oqUTbygIr9Q
WHkIPLPGgNrEO2wBWUrUI6WX6Af1HcFrdH7PK/xS3OW19XY6AQ5E/gyfyqdWim1HehXhmlG95Nt1
/HgwXsx08Bg8QnHMrjjSupNWkZcjuiLfvxZg4I7jUNal9hGDQNutWj+aEDs8/85b3rUibVCxOhLT
lO6zuXi8eR8j78ZDJiaOqjSpiynqWaI5P5wWiDIW3N5XGi7EU3gjF6rvwqzAb/1KulwqhVgr5qjl
Q2Gq1d78UFzYBK0CvzTWhhJ2sw1wpSttncXtRjSDtT8UKl/Z/+URxJurUny9AKx5lQqnsEvjtt0Y
pf+d9cX1BA+dAXuSw1iI26qDz/KozzgoLdpT3fLvmfIAl86AmhYRkvsYWkB9fuT7rgWcr+jvX4+M
qpVZrkpWKvlz4jTZ14iCkQfZPSnu4RWQ3piTZm8LualikdI5cG20G6NeBcztmMnG8YaoRwuT0S8t
GrzgCT7STspg5aji6F5jWU0xNKnaLGH5YhWqpzB6kXmBDb5Kvl0fzLuMvcPOPucJI6LkKkCOqFud
7LWfx5b7vn72huNiQtM6DIx4fHQD7fUvUSVE9ThfaHc9lsufop+bgIYIiSEhRO6TAUshh4DQaYvc
7KHGy7KMm0Y4pSV+65d2EOfaTXiq+7kWkV8kk8nfDrzmrlFRHQRrtPT2D58OcFk6qgILeQ68g9I1
mRy5EqtZnu37ib4BT1eoAQWjciIQOBTk3MJ4WouCOo7CX3mevxEMbDOBudNIwWFkIA2PM/9ilx9e
5Q9zQvHeeHSxRZeKTGTCAjf1J9yudoDy30Tus8qZwDRWN44SP9VJtkxIeE5DUhWCTzLifEu6VTEE
DCiGuYAIKCz5Td+KPzECpC2NPHK8w2GaZc5fTYBqiT+IjtsfV7zJWKSepu4Y0E8YwBrjC1alQ0an
pgmZr340LkSzhY5GLSTz/6TQw5YastcfEAYt1RiW+8uOD+vaSP79D3UQUvWR2d7rLQCauZyLTMig
g2I1hRBAM+/IVh1nB86SHTtzb4igQdXEcItRVv7KzX3eE3DfSiVd1r2kRpwJ3EZc+KRzqULFGdRD
MwNISLMLYg/XJXlrHmLpazpUSoSO3id0tJqnuK1+D0zRzgxElRrStrL4rpFKLpMKsOQFUfuv7TTD
87MljuSF7uiHvm9H32ArB8c167OLZPJnTeVSXJfuafFo/4mcNLZ0eab/O98K1UopCsNIq30oSY7i
q2BFRHf4XL5mDDFIPgYLTGOhLpNdtiAoV2Ya05o4vCSEFv97N0hquSrHJ0z1mkUwHVDYWKMDGOfS
BbvoI45BR3qWegkEi1TEEio+W7kjPuB5eBa8pfTpm4DginsVL6rhdjBSosp7huuenixGB0Y2WPo/
4KHJU/ZapPfBEbnme7xLbvSnnwGhN2lOpw314t4HQK3PZsLA7O0aSqyZYe1UEl8s6p5S9MyP/uc6
ZtWgckmmh+X72Cpdp5xBcVHKIZ48HX9VzoRtetxoySuKaj7uXJ0ljxCO52FAywkOD13w/6Ve+m+1
QQe0e1pn6w6lsJ1a7rEM5mnC6561qcoxxy1m5gN83KWMNI7xXtVclGKc4D2139qRIb6aZt6ZW7fq
vgr+fe/NTAcIj5+joaWv9lQzp9/Qme5zmlzr/lPkVeORzEKUIPHWoatiAzv0HnKQ8jNdoBiotuy6
uQoFO3OlGQHf7Nj7BQ2q1vnj2JY+TxWMm9UnsExXPY40iqPHCnT24fqinoThgDpfWmdTVquQBOjI
RcsyfyYX9yAm5o9rfcSi9QGQ9Q2PbuYd1YJk+QtmZ5zV93y0f6bxA8q80Sxel+rMBe6WYM+zkMge
05iYzpUm37DO1FiFE1+tdx36MSRjsztocVnW22cWoGDqHsh6vVPFPEP+UI/F5cgd4tTtZxlKrspW
l0KHlbzWNDhD2BGiP/bGMwK+dv1gtBSA6F080sm2+uWRRmGCO+fQAE0r12GGg+s+z6knjO7j1vTq
Msf1EHsEESG7dIyS9ygIN/4oNoDnLAwr5E7gzZV7u3COTaTXb41V1X6TL9I0+AykFydI8dEk0x63
PqtdN51v7/zNIKeJXgwASGDLtRToUsJMKqUYkIQLunUHRD4KjkX0Pfo9X+PWENlxXqQRYPrYEhaC
r4pFfUWyGpyxoLyI3T531KZwJX0bBdohQN6acX7lXwm7X9aRbzFAwAKqQKDTtHKi1E5CSHD2RqUy
o8SSH8DuAA6rBmUM0xh06n8sYdGNqGkoz/mldqrDy72MmP59UxchdYqKzHP37ar9INZQOp2X41IY
vRizt1dojewXpZ84HfsA1VsJXR0mU+VCUo0z0+m6/r4M/DVlCzjbsfstbKz+RioIOkxKVIsAKFFt
ERU+uAuH2BtyImPRcTzcmbeZvnDHwKsTHvpcSAM+ztYENToLT7rQof6K3FUt0JzlM5zJl++2H5PT
I1bIxsZTRGdx5NTMg60Otq3m+3Y4K2qg/y5uzpvtGJQIGJDFg6I2RXjHNRJYVa9Tb5nmUF/I6UOF
t/f0al5vOCy9zH5M4rabRL8MgZVLtXWGuwZeaS0qwiNhEZyWc7NFa4IiPFjXRaOtIokbWP4DLtVO
MnfY5NyeBsw8pDcGzRQ4Vmi7RMA5pLlY1HNsbE8d13gGxGN6v2kyOMc+ydr+6HyjT9J91wOUFcJg
uFoPGT+bZv1D5UG0KrvFRxifFZlZA0NCAOThx9MuFwYXFn6Te4VPGKbnc4WxV21jMChF4DwAzN7q
3jhgNlCAxlyV6kNk4zphS/bvRNv0tN/GeMkw/DLI5Zcl9xtwIs0/jPeHJTO33lxueL9fbX7An6aq
2gl4rykODrNgrXgK+3aJxrGqnRKbuJSSiCtWFDyc2UEEMjFlcMGdRwkxR01GDKn/3cuxBVK/DzY2
18q67hqXfZXNKa3xA9pdU8GtMRToxqKJt0gEE/YS9AA5dIbZihcnpBliqn2QBao9w7QShVgDDMZt
jDtCMNn6xdarqJ+tB4iPeKVfGqCXpU0noxGNAxEgzHUgouHrdOoMunPNxCZ5QdQmPYiWD750TAX+
Tjk8SHf7VnhmOKyxIXT8PcDb2GIT43FCfMmUPZVmpqUMcM8YFYMw2ZZrs9XwPV3+gwJeNklCkFD1
VKMDTyCiuyb/9VDAdb+Qlqn7Z8Z9FVMtaHYdcHQmYdHNrKibcRB4CkGfScDJwLsLNDtCmBOfGg/R
RFVkNc/nDLG6wGulH4GbAqZweB2VkxdnpQ1jpUnbLLl0mK7yK3df8KdV6HI2MnjcpmMswF8hH12a
NZhEDhapEKz034PM6/F5EKSOuUrIJnCSw5Cmp6UD44CpxyZHg9uM5zSGmA+5rW3VCHGQmRaXkcan
KPUiAlVfsHsJ6RvRSHZLar8fNXI1YlJD7EgswEdqr8n0S1QLlFdLr7YErLhIz+jm0LDGXhurpU5P
p7NJX2e2PXME3FBsrXftbthxgjMNwX6Q6CEa+fPI4uIQydHaCZyMEzirPQKcFV6EqWseTVhDJvUk
515PUz2RgpE/pLuNk/cFmRw7A/RrBnuFbA1iem3du4B4KVY1viHIPkQjEtGuUOVkwry8iRGefJ7T
nBB4OWwwdgk1C9KT/f1Td6YxZpZ8kxYyEhJ3/ZQgqh9qMK3PR6pjdG1kE7eKAUhDvmg4AF3A8nQg
zS1soURgCoxLqjTvsO0RPwPy/OxxYFlzakArVBvwSIAdbhLbJapibVlMZvjqmejjCBb1mj8yqPiT
NygKoeWJ4rRRWUnDbbfQwXw4d3ZbHkwpG5Rs7+D3JFNEgsRgC2KbThd1KQosCTKLQ42v04jDczd+
tEn8Mv+di9Drtp5P1huv8jldvOKuuGsBNQeY8llhG2kdZNhnSchxhl/5VcTq7ApS0fIbC6oIEC8L
5FIknzD+bTdOagBilFs0nxQd6NATdtnIlbhwTP31Ys/y2+i+j0+yInPriYbYU1YqCBn8PRSWzy37
lk+lKEdkiSs6bvsK0JThzd1K+Gc3YH2/ACTrQqqSQYbWtXDxQTibMIJR+N+Rj/cYvCmhVEhza3rw
QKBkAhfSOdooWLFdeMgyZxAmB0T61kvJLxCBfmO4fYQjwt68M/P6mJNZ+Qo77lv62p0Yvc+ZCN4U
al6thMD7r+QprTH8HAM2i5ustfGefVWgjmgTIdFdyH3fUR7cYpTUXORtAuzfJcL9h5Ppwx+r+7pa
kPJ6ndNZnNL9iOuUMQNpIhbBFTSmko2//qfGkIUAmGtCOap0JYHKgyrTxJ1BYPbcEVVPnqzoHjio
AzCcjoCArRI9QsEdWu6dppzlpmCSoiKuW8oN4ylQUTe/4h122zdd/RDP0QFIIQxW2fegkAXRMUMQ
znkigXC9ez0VqZdhIInfQEx4nXGCnEBoy8nJDbPJkUw3F+fl5RPcKK32/Y0hTBvMlMO9UuN0LtN7
SQ1abYrzIeJrcw9/Fwlpo+edRqmXxcQp6ZGBQLBQDU9PPHyfK7aFDtnBwfAAHCoKSGbmXqzpmef/
dLPx7/EjgXBf3KdFGDNcli9eiJy6W00auvBZOI6uS2bj0UCBn9+Sa6CTSmpOgF6o7Yulz+tKgjbZ
8wsBYVggcVMCcV+8lFW9WZ7zTM32XMLWxP5iu0J2KTAq1cYDay7s+ajJPwX5EoUO1ymRiouHdXAL
aenpoxtz7RcBfcGlscHtAV6ypV9YnIPCIvCDK2g70Eh6cT9o94ud69c9aKgAMqLErE4BHdvUvSZo
gojGlr0MEueKB1uDSU7uW+IkgxAAjlJ2Djsr91JFvq7AUkSdvt2NpLPWXARmqpp3AfKs+rP/3sFB
xEY/QBHOrheABzy+/x/dAIjealekz+KKUgaKUeSApGPtbyPmsYYFz2ow7Cu5DrIXaQIHnMwhC6nr
kfBBucPEXvHZhOVjBf4SyCo0J/gU5OKmZv5BzgtLP4W0vkioF0kOWWgVwwzAJ2DyGmKgwmDZkfkw
msQlQ5XEwnhHbXkKD7dSBg8Aoxl8BVtmFL41f3MUMWt7x5CVPKrWZCqpwQgqHsHEUh5YdOpMIDfq
pxuAF/GlfCD0UyVFEGxH9wcjw4/B3/TLBHOhYmLpTgoJVVlT1g2fZ68Tmo8ZFmU5wE1FYjPAIU1h
FWCdlhZmMpipR+fs45no/HcwWELR4gZNVj/yiflHp6yYF08l6xd8RcVviOLnyYq9PYO7ZjZduRRU
KTog2avWt0P+SaAuQGnJ/NSo2NMDNasRoBVBJii3DgGCr5VGx4FzMIn8c4Ddf4jc2XuMJPO8Zqmk
KWNPWbWSl93XfsGXZx8UsSAQy4Lsa9mDrTirDk8Xj8LnfN9TnVnCyHtgoTLDiqKKn+z9GEjJT4pB
pebxPR9d0m2FOcXKfIuFpO5tl4MxqyUiE0+P3Zhm7ND4+9XEKDE/EGcexM2xPrspIbZUf30JIr7C
+f6ZOGQnOq6R922g9XShpzu2G6udl6GOOBhVSjE/z3BcC+4vQHMywrhB7FPcwLa9BHp8RMt+1wQr
gJNNbHN7UZH5o21UX6CfmKQur6e1uC41goGFN8YwHU4YMxikRQ/v7/+MlXG3WQ68IhxQ5BD/LY7Z
YqdEJPh3rfxzLoM4+x1amqzz3YM11d/QK5CQe0Bse7KAM5RCJ3jw4s7bIksTGQ8h2QZZpwdEwVAx
P5GUcqZMqc8zYzEySi9l8lqlWPgWIsk8jpf4io3lKL6QeVUzaxhcw9nMhnGQ9mgs7mlCnUXkdf2U
JnecTrhy9ATZcciD6Tmo41vAfDWiv5I8zYUWVCZN4F8aqkc8Ww+keGokpxdkJXgGoM0KihwPDaM0
EX9b011P9L4frak9xt/sPQTlO6CLuVwAtwNIfEXGbh1AFRLSEPi/pZ+2c57DJ5NhyHLo2xp6Xy/d
PdQHtgSCRFAy+HbTL0xg2dK/PZfY3k7BTibKwF2N7II3G6SLpDuvqnat/IoBE1bqGtrgG0bfZxNU
IQvjw+ipFUrOhYwDznYqopfB6mYQ8LJ9wbpswDthGUegh30pBZLXKpy9IbtPdy+HapsYKTg6uxPA
CTKiMheyUMek1WIA2WuKWrPCF3iMIUXZ4/lrQrf3h1/045ksviCCH2IihM/SZFwzgDAsZtlx6rj5
E9xJUO8CSmyskucbp91HjCsAzvcfOWII1l1R/ZCa7DDpI9z2PZFmpsFMJdgMw/GL3kkCfSE428me
Jkpw0EwEe01TmvcupfptUT6Hx2rTSbHtczFZi+ax1hStXSwkUIrlGHvu2e8HMqXSulgbpl05TCmJ
hcYo/lvHPBj1iWHO2MD9uaJu+NK2mGY+1uUxnp18a1f7JFzUKmsH8NbARMsZcPc9tR0wM5Iuosqo
nFjIXY2xqQpD4M+0j2JVyYa5Va7mM73ShLbMQYf6wMvWZG4S9DnCkfteB+rV3XOGjQS+W75NuYv8
s8uFXM/4sMMo8u5cg3hk+o4ISu1HtNOYF1VtoYd9w5ugHlFDmCEXhk18cp5JfIZx3mNedqCDny9k
72EA89G3/z4ouwTK3lzdmkBSZUIOotBUrxpalw0aysJ2qTPh2cEdBPOCHzR183c2G6Kn+RVcr5Bj
UG4Y8vlz0L8FBzTaI/+dOqgeMIEYMFIouwCwwGxmcSsQl4XnKGsrS3Nw1skDer2dRKFRgIuCrCdT
vcon4N92qOlWiMV95xvB3DGLwxsgfdRyViv0tz1VicRbyZW4pqLWkda4U7s8/Y2O2O/AH54dlGTN
BfOdJF+Ft9o+Xxo0a2kZu2+23VjPnzS/5+L5oI8SY83SyEilD8GPjZTe1FnxIz0aT9nl9psRAbVd
oXdaJyNxj+TnlVJ3oPtXsbAN3gTgwX0jfrbAEv/LT+Mfk2ElzHJGFZiRisv85ZTdG5OuFwGmPonh
jDq4wPn9tKpemNcLdIXU9F1Gvr0xwOqcMG5FzXlNAa4MxIKNX5SQEUsGMbEeJT54BTzXzsVDikIC
pploxDdUygPbHKM4Vrq4XG3rFI8zUWKS4jEz7WSaw3vVw+k1yXu8IUIMNCzJyepffD0H5h/OmTai
UTUV1754Sk8+g3P8DfGKF6MjGJFRGT7YO5rWc984XU5NK+cg8Ome9SfUtqCy34dNvWQICCIAY5LX
PIHJ5TC15/n/c9cwpICU3MaHFYhjPnelr+aaJyX2trSPqxOkCioLX+jFJ1L8GH91NTCR32qxFZSJ
fQhsmi24UB2N0hLubnNldUVrCsF8g82amEjPIb5Py3YHbaPmovpHgXpMFkTi1hGudUs4D18kzTsn
JKDhysUN4cHHJP3dDC2F79f9cfYY7RfnbTxUgWsnvTXT2lmSBMHfq46dF6RqrRf9qDXCmR4HNBml
zNQARPN7bqM45+GoJwwpJvYgM9AnbdMWsKvJAlHV9us8Y8MXupAR+bDSsAEOtsPrHuo2dzxpEhoC
uitvCgWByawb56LW+M8Vpi4O2JN/FCXHZi7cP1tJU2T6s8b05fO/VqMXepawAcpUB3h36MdV5ztl
INQ7iutCIed0NvRLyxZiH5/a5Z5hKh4IGopz3Y1DZPUNbjgJIVq0FMAVDqfvfweq0SKE595s/Bhc
MkG+AmUSQ1b9eMyVgD5NZl+FhQavzWoewJR/qKV2WM8TwJX2oon0F0WHHh4IjrQ6qN62ekyZsykL
Xe9I1Ahp6wCrQZyLEw4IJLQusanYBpbq3SALvbXxGv6IxYX003xgQRL9ju5ONF7o5540DSj6Erx8
Uu/jsDtmVTvzb81Yhy4J7ZmdmuO3Rw5BEQUJWPoFwkO8CuagfhXeIAK+TzLlAN5uCJz3jhTpaEP+
KkGRBRZ1LNigGTxbVtv1qEWfVH8mcLQ73A7FHROZ0O/EgRU6NgnakWWQIyHo1qxjAsUAcw+53P0q
GmgoBm0QUcqB6FD48nWpXpHBLTwaO4t69kRArd2OaRzU22ah8uE1paLBgRoPvIhb/xIeFlLG7jK6
vAN/O5yQPZyykdCAnCmatVy+AQxu0qW3x89ZAD6XkDItWkowyDvbMrDcIOilCRW97CjZJDyz+/Gw
Ybzmtq3O+oqqXZN5w5hxCjo7R72/TXAGdn1x43MgcB61/b4uiM63hEFM4jS8Z20zVG5XlshH97dw
To/s+12I3RLyS1fF3Pd93tPmv737zOzZWxuzPFtd6J21roOWz00agcWObz+4Nxc4Cv/Z2nfpC6Bq
bFMv57YylKN8tkLVe05M0H70b5qcExqbTRfg9+iLDEIZ+g+n1Jicg3w83WAbxzfNZigAYwst/Xgy
GLFxNCVFN1HCV6F9H/n03KzrzGfSe/WjaonPsdMDB9T0LkY1+9XqJAbgy2PcsuLmlmdZDk6UT9CD
au49ALs8AjcLtNhY4yr4vq2669Ct7NoERyrgHa7sBVC/UzfGjN1RTanlJokAE//Xcg0iFTGR0z72
Tzd91tnrTYITUhqyMRFkpzYtgAE9+KJEwRQq5Tz4mdSbpQY40+GvNMaYESlMo7OsFBk/3wNdqZhl
FQfsj4mWGj0tFhMdflNKUb8dN4ry8bHyZHKQIm4N5P0shDKO4vnvuiK+8x+10AxK8zDR/Lhb8dRF
cCQtZ5jkvF9XcXGrA5MPvnml2DizLNWaXo4/KKcc61po3SOskhaJ2fCV9WvSXxfRR9GbiSdXFlIi
1aWEfcq7IK6Y3rA2HpMEa6jStHGlj//nxPTGlMobbLnIjvZSBiYLcVd+3tjo1axYDVhWAGNOjPAz
/YPtIY7UKeR/jHiixrjRZv4U5AZjNSATDK8Hb3+1BQfF9crYgdq2PnTuecsb5cztQDPzWn+Prpl7
gkJ2eqpRd6lMEW87f9O9dS2tFAqpDjiLtmH8tsaS8ZTx2jEOoSlTGs5RwdeXh7PJsBpbyogAFfRe
rr9gx+z0WHsfzMK1dKJU8xF15HusJdCCJ6yRvj+mMJ0R8TklRxJC5p5U3/n85af6stxZpJUHSrm/
4X3xHoWgcmbVZSVWXMGNdQ5BNaX/yMmDbaIr0qpDRcOq59dvYLFs4LFI8blabMFqojbGXKGu44rH
zlE+KXOvWD+nP4x3mJ99CffJNDJOnZkdMDhepvXJxp2QBgXNgaiQko1+pux33d3ECUI/DD2f3VbY
m7Cnub7m8elYryfUQnD0v4GRYe3pk90uZxnSTOmFbVbSr5/H0nhrO9alGjzCmYpGWIy4Fd0bDWBu
kctArk9N0hr5gPiaYMhly73anroEhckyHtzA5f9bAeRYea4EzV3xUkIdmLTCj5xxKzPIc+EMWYOE
/LmlLEhWXev65tOrYwjiORGcYti63NQ8P6+Hz1UDcsYkOxrgQbiaLX4RuOQzj++CtcAMbQ9YP3J8
pXb7mloI6KsufmrMY3aXHNqi9qh0XAB6lMNE0ScEu9Hnc8Q59cqZm/RxnRVynv8O+KBQT7kdbTsS
g5mHINvM2fNBgdBlrCREFLFZBn1U/CI9t24+iTQooY+rd2WDzi0yvy6zWrs3bVCQqq7Kiuml8g5a
rq+MFclRPSS97C0upI8GGKByb+CRWVge66/iHNjTIdq/3isVKk6B08TCb8yY0N/0UwM/GT3WAeuG
mG03fdqUuowPYdv98GPOA70t2Ty3UxBtnGxhWPHhzhWq2ATKZa5tW6iuuutZNK+G74l3ogFTyXMM
tfxrjjHWKk3I3kWpNHDNsMeg9FxF4OjdiyBMQ+uUVkljYhuqbh0fGctVJPnP+oGHnfp4E03NWfIg
kXODGOP7ArS17Db3rzNTdznhJMWBrvq7DRSf0S3qCsdVwz7FkHs06FAglNXwilJikvhcBKuPyedu
UE/KmeeHAtD8ZZ3ykZ1X/TNd9ggbYTbBk1tY70152TGXOhqsisOK3/iR29NmPiNhV1Q+5zljwh4v
HA2hco6Eh+K8gY9UBJ6hzy9gO2t73v4rgbYxq9F/xDiHfwd95GCrW8TNUVaN6fjPzcz9A2kjP+pH
KkG4gt4GSHAvxL2jJ0s/SBTWK8wpiFMmDxPn7Lh2eeaNYJzw3Ck8UerBsq97PdTMRPVMC6s+6ndv
inr9dXPZoovsF1jmDEY2Gg1VRUcsiVwjT9N2jpeJvqnnLZcKDcqp5QwxsSCFfid3Lgqyyq+Z+Gce
/IUCBzb2wPLnXc9c+2tzLp93GT2x8HYavu6qBr1w0h2aTyegiLH0hMHIoULgYpH5Sg7tYiO0JX+J
MhQJkRlFTF+5glx9e6LJ6PJ/7iD5viAoGPpeR48iHnlXUBh3mWl3nzLl1oiwdCVwyVRRm3CG4Dn9
JQS1zQIReMJnx83pT2Av8/wYj/AvQ5it+0kOQZYo69mak4riX2X1+k8EW50mS54ET0I1TFrxCLr3
B7L6BqJuraoZjQ4TqvecPGjeC4Yp2tQ0YfP1fTi/A1ZtsB/UNiyhdQEXTuNqycIqjmKP41W4bmop
ChXPR6Tga/3h16/D9TicAGqpRbCtTBxrOEVmIuEbo6qbxwG3Q2UCH2Flzpv2OAJ0wYFDOseJU07r
XiL+ZiM1pgGygfz5v1BXCMwwbWkb/M378KpjSZe7K50wORe8LNU5jr8coz0jxWzjzTGOGJBo7VVy
+9euechsEGa8rxT1tDNSJD0kczwYVz5Fb9b1V/ASCg06xlEPVbTl7c50Z/1mxWSgW8MdgPkBGB/1
7nPRK6Yg3c8bHDlHsMEA+mfLQa1NpNpsN7wGIpl90gjVfFS4xnjGIkT9Axfzx4WWseMi5t4UY2si
BhAixelscMkf9nRp90rOyQhs3NrIY75hHcpxb1moqVoVeptvQQFtsRK+oWscShrR/GhsAA0jtoMR
gExlJ4GS2TmCk7Hn1qg7tQ0I0W/qZROtJul9abKT56j1L0go04lEsP0fwqijQQPENKY6eaeBOKd/
s1yoLF249uXQMc5j/AMVdpjMwdvzCmkVW01N9DMXD2tdJ2NbxgAVFPsvFFLYPTLy88i23InE1Clz
e8WUXtBP15o8oj7uKT4pOV5fTpz4gUA2jEIdwFuNiMPMYaoXqWpi0Hop/6ylPesXDSOZMp5LVD+h
s8GyYs/9BBGUnZascq1pZNQ1SJRmSFjICRYMi8KhvRgkBjnQJSGwBU603kSWIK8R0wTJHjK1nrmU
/orvCHE54Gx3m+LLxSCpyExnhKo4u31HyW8y4/5WD3PMGFiUu3tkK0UCK8cZx0ouhWvYP40i8cYX
KU+IWYz//odQTD8HjSL1J4VUWlCIs4rqEpqjY1cvyHckrhFWdBPWZJ0wgaSIJGmkbeTXGH+35FXk
zbZJYm+0IfD6LbDmCFmvhaIlN6JPvii8pKvNSqDtBq5CiKziHPnqTitEgzWCzBNpOALv06C383e9
aufnALr/uxGbyQMBYk1s5fmqjlqms1spO4+IvvY+UkDajj5SwWWU2OtbNZrLHgbRRq3NS7hHtOr6
lP5emw0HFj7zHgqURoj3wcV8bdB4lKYeTtAJFcLsCXXDrCagXomsukNdt/3bJDF8QTK1xN9DhoMW
PTeM4AZOPsE9mIHTRKKpysrGCkrOgE0teaz12mVLWboDQU2kQ3t+apXV7k9m4omJi1v1iFF9QjBQ
XhIKOzdnbGgcRZweUhpHkbgx1z/qL7sDvGC0Py+HOVfuWYholgET96lmcJHymbzDsX2anl9gicCv
QRI9beXXaKPN7ATKJ+cUaZyLIliHnHkrDo42v7HLFCTcX9lg9Mfk+TajBUOpNiDuKMHia1aRIIY6
3sn1neduRRNNv4UqZ/nv7J65w7mmQr+XIq27wtLTaY0XYzC59t0gBOnam9AnJMbb3FwOCxuwXM2e
XyC/u9Nce4hQBDj95+aM4FCpJBRc0bi8bGoOxQL8U/6nvY/8lJF1X/M+N/yk6Q/487KvGF8TL90z
W12XGIdv1E4nyyelxPSvevvuHwU4s3pnRF3ijNWWWVgklOhMY/obQEd5DmIp0CDEtHWxWVGjAXyP
V1iH+K0smVnueMXqKHlP2iCovYSZMvTbseTmOT+DvY2HyOpzZg91cjlZLq0O3rzr3VSIvumCbuMA
YXlhZQJ2CkLpsiqkwKBdFthdJVaskZKcuDZub1+RdoLo/A9ojANKEtj8K9wVzunhPMD147rUO8wF
niJvVfhG49UF8lpUGeyZbPtTzI5vuRSRWnk2wI71XPtlVOrN7PA7TRSqlwMbFOsFwWBmjl7Jiko/
aEyTUU+paEHipr1hZ8yqrcRavTO36w450J5n/35P3NGuw4Rcki0Yi7hIHQqUwQx0I057PHI/xlVd
VzOcZTozEUW7IEr3sET+1cw70Vw0wP3oVP3TVgFX0wX6NUr/BEuPKnCmjypRwdNF3+3Uum42yDLE
mrN1R95PKWdI/YNmT228AAc0t0mGoNdsBYhlv0pwOC6iVp+PZ2AGbhS/aNMfAG3L/DKMAPeWw3Dg
ieuBQe9Qfj1Gf42td1X+RAMxMYrI58QdIndfbU4UFVFl+GTEocPbQ4dTDtftF7Cl399BbC7gKVx5
SmxMB+seck4ssFDSZIUibnq+rj8Y29quIlSGXamZVsMdz0CFMaii5aK+btPBixto/lIhT+TQev9W
sBfZrGUCPWb50RSEg4av7B608SI7bqWG7Jjo5FUAWtJcc03j3jzhCoZxISEme9FICTC6i80MUJlZ
3t6V0UT8bX9AVTxaEjxNUa7KvEqdHLPJzeAEgJDYPGThkGH7QyGJ5yjeowUnf2nmE2XgJaR3rw5Z
MI7Ow/Im04PAtTGGYE9MPEB9kBLjoKW9pgYbfne8BjxnWdUAoHlC5JJaFvN+CiGsi1+0c6h5Re/1
MqmZi8vDaYdyOQ5JoXb6m7GlA94zWV4ILH0ngXnuU3kL7cKWQHxEFG8DNhX/4Z/ecUqi0/gOZUst
ssVq/Un3csSZtvtPF0B4smxc13VW1d6Mjgh1fa1/A5G9ZbKnYF+27DFN3Bhe46T0Csn76W9S8VGU
QBuRI5pz7IGVJnZG0uFRGMsT+Tt9vaTPwGaITeBX3aiRUWByJwjrpiZZ3uoUbSQVms6bwfiZ47Ow
ldVWDUDH/LPK6URArpcd+58ck2eFOnBqJNG3y0/rCqC8ZGEBgMmEOnrLf0mYj6lVBRox5dIwS4ch
SwAgmPrwiyWLLjL3mAVFod98jw/zXaRGuIEjDRJOon4BSCQF55zVQtPEz4i84IQoSDEAAjfT3gn/
S0GP5iDsMfq8kuhR4laKdLT2Xi5908hc9ijMUinyESqX8+qjvApE8VDp22mQQ/kTPv0mIluMaI16
0YAuM9VTsgezbULYY6RusDrw/cGAAN9Z1qYNoe12CYdsgxsxSO5I4nNLRbbH/T8C+X8J3+oLxWwm
mPgBOrG2uxe3f0avC2w7wAOJSgTcRLMHWyKrctUYvv8Mk3eFJ595Wtep23WlRaGRIRP4KawL+Ezn
ryKblWbAfTSHGBSwnjoRdllRqZFz9TLQxMn4MXHg+NTuRi06oPiALcC6UqiSuzH/dsMQcw5mdyr3
4FwVs7aCRq5bSHKub7hjNn0wNNW8VCSG/qzE4La36mpZtcAAuuhg3KKsrKWmJWe9V1VLzqb26XV2
kSRRl5umGePLLo+tav5ctFCjt1NXv/bwcSYodgmJwSqctHB/vzTeUk/UpIaI9penkYKOGsgq6gaK
3jbcDlU/ggvcK9oUZ2WI49DgPlLrMe4w/9WouCwg1/HjYSUe0Zd3YMwRveJL80cKccVGVaiF2S6f
cHXUB41IW4ZhK+E1VTep4Da9y3gKgS2S5CXgadXrZM2UBlaZD3WOyNgoZdgMvw33e6QFCo4l4Drw
ABiYO6yT31R6vJxW1RbzKHjaZknR9xcF5kg0s3CJNrxxNc9rGcdhBKVAb6f2TtiapS1206uPacYX
lendfoM4INO5ancN3cLHP3qXyk1pdOjCdNBPbM+FDTQIvM1jsZyi5X2RtdvCwQ3ix/Q7e+y5Mmkf
55CRV8+iwc8MlQdPyXEuoHFDynMN7BO2cyXkx5gnh3fHbCfRJ4hFU+b4QP0xAGdVKy5MumU/IubN
j0xiIji+/UMRhli7R++uMu0eMs/BHXlMNQqJH46Pe5HVXECCDHxvmzCz6hb12Ab315Ql35wtnw13
2ZvB09hPvsfywk4wRM4oW+QWV6uVGQl0+aIVLiBeZD0vsxHde/B5p/nOBrrZjvij3lHOJkfv3b8V
rO9pit2xSB4GNiHIm92ovsfOwvieBdZO3xpceVrSGtxd7tqkAgZaf9lFaGB3OGGAnk+Tuoe3lNgq
1zRRBhXNe61rbloLvGBz003tDPrj9xoaHRBVNT1FjsnrXsPgNvubvzAczyhzqZAZQr50PqxR1Lq4
30ecd2PXO05N0o+w+e/IVD4QaHh+5Zd4NepppB+T8E30ZGwIHToOBpQcDV6ldGxSzY4PudeTiXkV
SRkpwt4NI2U6s7+VsWrANRlM6ns4sSZG3Q+G3ktffC2dtfYKU3zeTjf/TgJRq+USUslj8XFtrErN
UBbzJCQpubNBjuOGi3bpSeUT+Ezx6Rmyx7+eSCdg0Xeuy6FMrzUU4sRodzv1+8VCLyH30MkZIqGO
SzlBC7M0/Nt6jTxUQxVRsaQkBgl2MNSJznM7PJ7IRY7rx8HMWmlb9PEkF0dXhaOpzjZDj1l3YKKD
G29INddmXWAmc7ExGXU3RbHsJt3JP3kWcemZQtLMNYUVn0WKUSI30Zx/RSe4yVum65Fr+LmjxrKZ
/+GLD0MhJt4OOx9Lbghv0q723bhJFFmlSA930EEdPdpImllCZHvQsPNM6BgqVADRo+FDmoxPPIGL
7wN4NKmAVCNbz99dZ+GpFRQA4lQUQPQiRTAXbT2PNIYQ0oCeJANOZqpXSQ8rrXGdJIa0KVMfh20E
e5xs/AVJxAdn7EZy0Rltkv0XJ+lL+UN1WWXoYYbYAl25SOLJ30R1G8hq8sqd27/Fy/OJKUAq6/IQ
Q3sUgYzs1UVb8GhZ/JuEG2aLlqFy6g0VhivbfiZ49Z1J1UguM9EKMw9ACkPxYpmT+Bd4bQll137z
swthQsMqMeOeXzk35/L5l+FsQmHGePvtzyAYqGK5mhSYcDYqwX/nLSpt5XsqgCoJ2ImGFdcivGzA
UJrN6j0c9tUWHCC907UNQjazjlTVz2DqO8Kjen3MdJpgfQY/XchU7kFtEVVfaqSZsHxjgtTRkxQ7
SbPs6i4OhNnvsHhGfRnEth3fSSRZZdSuF5ZuyhJiKsH9s7id7o8Rt6gaTzIQQySs4RZ1a0omkwWm
Te+zwDsJpM64hNRK+xAvyESL9tbJkTpgGfvi8dSw2zs9Nyz6YiNj0+fg5Z0mp2PL9JWs3zlyUv4m
dPEZUd/KLeQRKucthNYaiKR6a1ZLCuCqJlECnPbpFbUBjBrQWMui+G+3NB5J4zJ2UjdFxXEd390g
kmvws9VXtKEuCMGOcqTurG/QWIo6FyeKrS7HU8vTegdaG2voL1sOLMjvLIlIErXDx8Ldi0F4u1hX
v2IKcEAweirgf/geFj/wjI+QOyfnfu4Ms82PByUmq9zA/bBYdzrW0LprKIuPNFlQ/H9puRZhIxX2
SZUn9IUeyl1S1RWH0tqdCJDXYLrWF3zEC3VohLR91xT6b0GrIs/woAFG1qPgyHkiq6X2sOJXFsHt
qHg+z1q+k1yS4vz5dJtbJaWZB6YmbczXEY8yUjWf6xB/bW0yTEJVU/RC8bBid1F+ulM3fFdk5j0+
LPUkMYY5NBP3G7appw4iKT+9Wqadt/wyxrofis5FQS/8aXfrMxlQs+MRjsIdGjftlJOnJavNzgXx
D666QrYHLQ0qrd/ARfrUCzYPILMf+wvd/obqrvieJZ3JkJU4AjspU7aWaf0wDAaiHlB2YdhuT0Tp
VLEP/AssK49ndbYqFpvxLI0FIiDj578wxMzMLV4X7taQgKDKrbiWJ9dZgMxfdeZAEosxRpvZxGGz
Lw3JkTLBetPHSI7oP3IhoDWqNemMIRtzlNujW+GY9ByKH7zKCqR1KmzsAy5Cl6e2iGGix3/7tis9
EXzQVqTksJe22fu+VxD+h3tjcI0+E4ctMZ7pUfzB+Dfs9VnHq/oc2uIWdqbzGVNl33I6Q3NRvaZu
BxG+R6o9IH6pczpV59fDCj8DZwMnE25M8tBIrg/qtnhbWsYXsY9jxV+36fbOkFlA0P0aQY/k2tSe
z/HwvB0h0L5aitHG+gT/yb7TWgI6+67UDnSj4VU59kPgW7/dxG1NbNHDN0UdQoaFKKaj61j5LdPj
1+pwAhzfA6qyFf9t0FZbcrhkQknO0B5K8WtmMU/wXp5z+/3fRPDKMT+sYvbtEaNZFjSdYeabNT19
BXprz7icjjEBpEneLsAwBn/ELRnG+rnrcn+IjI8KnF6p/EFa/WddWtk7IFdrLMp9S6Qq4yx+oFcI
5vqc/5UUhOo98xaGm2BkVl/Q1RA27A3xtyuWLjxzw0rQXRrYNNgBiFYbLbikREVtV9AEtAWr2TTH
hLtJ3uFDkffOxt/igCUMrOaxF5GORYmiAGzutHfFbjQncnfEIpQ8y5+jOupcYF4wggLcwfBYPejd
/ttIKLsiKTmGZErAbPI8tG+h2I3sXMZgcgYt/QBkfSXrAbaFbAHBxLIePXHQOoBf9m9mv7I9VqpU
en/EgMXyxBrqzf0tavJ1ww0bs/qTX7aeHM7JlRD1VeW9jorfjLH0AGyULR8l2hRUlM9KJi6kXOun
69XNuJOORGUQT0Gp+Rsh8T0D72owuxfyDGM0Y9vWhamC4ONIM6XQ+uDYQ/ODwAnsNdzxpucgd/uD
tDmwhsRsPkhH+Ff15SIBKRSFdxbC/bBBkLmsNYtZ1iLhhs4ukxDUaAee2Y9RXQYIUT0pJCQbbQto
chc8zWQj9/bWn+YMsyx+f1YTkORnUzWRqk1BeMLFNDtxaSM0zJJwYg6D4PsACd+oN2pdhsTmzOOo
oRj9RpKi5fZe+/HfMCwYbrhyAx91LBKxndOLDpDQdLLwyp/jEHF5lFy2P2SeXaVDerzAdOZlZVOA
PUyKgXm+6g6Qf3R2XjhMY+xcWyEl0T2qyOK0KNMLAHvwKyst/EkG2acbPyXyAS3pZ+NRo4X29iKa
2zX7TySxRKidrybfWUv3BC9sbf3ZxC9AAHhfvSncXTnGqUBi42QfsdxZoqLliO3txdT0y0t/6E8f
BPhwjWsJkyHFkTjERCYqetrEnhhuGv3TdGtuqWoMb9XtVYnzGQ4OIblPUQwjsfBDd7sLVylSjrr5
7n66T6LZMuf1AcWu3HybM8r6WGZcNEnOe8CiUT0QHONGi1SSlK75gNU/e0cvz8BxSroPodErzkKe
1+3egcy+eo3fvTNAsqTKoV6YBjTpRHu4ZBpXFymnOTt9VrCxnSDbwlL3uZYeHW0u0y9Q96VmZ1fq
W6vUJdNDySBJRB97ozrJ2ws05qJwGr4yZtP2w67qdBj2ySyJc+gyOIDV4l2xw+WvuQYICTKqEX6P
YEnfnmW/Zs08uyH1IvCZg6hhjVbblzzAw6OXESDanOeDLv/w+T8qN9yeorMkEAltWKYFtEHXSJgi
GgW08EjK5B6AhJh33TqfgEuje0UTKg5ppCBeIM9Hnt0bIGoA/Eq210EoGkkJ47//5FmS5XxEG9ki
yzWzMJbS8ZGkgAL637oA0hMSV6N3bsRZLmDAwYaNK9UTVsgkp/my8j/qA23jgVCQRLQVP1QLvC6o
IZmdoooA4+1sLGDrXSXcWowWf+QnlWV6+Ozv1kfsSR4SK5NDuH54NpwsgT3QgSq4m2QTw29sU9W6
TNjwhn+x8KRu8t8WA3+8/ebfEc+tAWDZFrJ5I/mT8bbMnddpQxiFC7xKv1LzfoQzXyn1z/dv2fBc
BQzz4poB+gtSQWdckLeBlgMWjJnF7f+MLIgRYzGYcud2C+Jmm28Rlab68NiEGWAird88Ay5Z9DCO
UKIBZdmnSBucU+YpCFjjsCxxlw/ZcE7xi19F7J0qYMXGE/UomP9tWehhELYBV8v4mr6pYR77zgme
F//xqiAvTOkMFXtQCIOnhZnZRVK0W4xb3b8+dztk+Omfwy+f/70sBYtUEgCVEQIc/g/obR+T0QjC
miIIRkwITtbY7uSKEyXayU+WJBVtRTvd+9NVRF7r5a6L/kBAFsKUXX6yVn8zFz+LHjcTN7WZyDlT
cYRJ/K7NyrOTsxJmU9FItwcv9Ydp1wwkoHcj0D6ai/In8CZCSujZaGvoJnst+lqCoPcCNhrclQfD
S6W1LJb9IkUzxOYYXYcyvVy/OucYZJn/kSGdG6AbeaF0/EFzcP1d0povUSNOGBbPHphVNBP/3ysq
TmBzYHBZWrBh99KrxHqJUceD9L79Og24JYKLlIJvq4DbXMr39GRW4OYOZoJeh5KfFyKXmeXLiCFY
MuzpK91QqFPsfco1omrGYF0F9Pamxi1gVtBjFNZANxxD2sCUaolhyhD/H4ZkEkHM6NLm0uxdHM/t
CFr4eqCvHjaaYmJbU/DLNvViNa6du5UsjBvZg7wTix/aBN1L5l+pwznE0JC+B6iXyii0Qod6YXgg
7vIp8lY0Uw7gjRwsSMGzmc2pomC11DmJI8KzJp2hsQjCDySAhppUgLZJa5RTESy1e5hFFe//feq9
yfelvKwXPjvYhCGJhy/XDIu62oo+8prVEr2zPcDeL27cyDuHpZAZDKnnOntJ99MmWxAiRbIeF/Pp
Vkky4HFhRB3Bgvqjw52UgsrRv9LkH5wcZQ/k+u37Qem1GRmaJJgFniVifOsg1i6NRAQd9jlIbBoJ
YC3A5F8gXorxfIdUeP0fVeIQ8+XEb3oxupsJY4uuZ7GCmXcQ6GBFmqU9VcAiCpUeERlzlDSNf7Rb
0x9flSRg0yAFVp75bJqpbL90/9S5xB8ugI5xRR8JjvzG5OYlvOkGpHHeaAvUZkwQrOqI1iZv98Nz
wjhtqEZK3XJtPgfe4YYwDE1nSOxPLU5ugSlQaTi/R8FTuElqy3avhMzu+tg1qU4XUUhH7RV/LjKk
N0NnlqHtuHYc9QCqEQb9fgRfQrLz4BPDNyJ1OoKT8icOXOBAY4igmGKJElue+QFX9rIq4c+3a7HX
XC8wJxcCsxHTNng60LMtUg9Cubypy6ynWB81GnhVkAhVNyO7zoDC7uq1setx7WrKWAyZsSKkTTDQ
0mlpH9Lt+G6alZ9WlLi4StPEnLYxsXLWS2veFLsjU/WSkIghk1/fPLTt4ym0l5gQHrWyj+tloIve
PURZG/KF13QRy1hdm3tFOgLM3IKhF6uIQ0At/tQDCHfBO8TYy0k54t6uuIzSvYM+hvnBIuhGBoPa
UT+WeqnE9KKJbXHWbQaygDbFFkpXOAu5nuLMsbksjCnW8I+Y3vIjQ2+lCqTKvP35lave/YLcZCFX
wPAQOPdpVAvdy7gfxw0J+bi3i/ch14GxtLuZqrW4jN0414W7F64JJ0z0h+vwQ9N/i9dmaVqsI/Hm
Yl40+UT5i4nZ+dEDqk7bvfWjLPyoJI3SvZ8Y6y/IvEy3r0fc0GZ47maWkn8XURn4Sy0zQfgWlxxu
b0ObLu7Z9eBuM9uqVW8FdAu6u6EUcgwqdGXCqkq3qwm4kqTLvUxioUM3xmwSEhaIbxS69cVLlJZF
QEL8UOgSkHG4ujP5kfOPIACO6eSBjPwkJRxzO9b3wVrwoJlX33zYF3IdcKs1PiWV1wz6D3Jz/1em
UeHqdzPRjHUmJNhy3R2HqTN9ZP9B9pP0lVAdZ5pd7lKAvpHlPhPLWCXKtEiVFXvN4LM31eJ02vbd
0CHYlVwDMJZYNjGIXMWZ5VhbPNy9PPsADdTxu4McD2fbQk1c4XZPEoO4/B3TMuXRaeIuv0rJOI3N
RHG4fLq/qJIkUwy4w4JbxHMxmVYEBd/YNCZicJSNsIKxSL/Vai45JjIySpAnxGDwBGilB8SLEw1z
BMRRi2qgY/xYoGU1jzWFKMC0ELayQQZPilADEZN1MV3/kHcbPiXSqSswRxBpbO0Uho8uuNptgBKG
nsD+pGVjKllC0SZ+YWIRMDzUEWalKjiGI9xnh+KseeumUtBea9lpDeP8I2W7mKe+QPTQGfVEN49a
tEezLnq4MNADNvEuotYUxA8YUTn79KCf1bW7vdqdhYLSiTHKQzLh9YKsZ1YfVV9KLjZAEz8QjSmi
hUOENQSR30uuFYmXpKTjLkPCPUvB9MKkx25Z5jDTTMLxcSC8GqSqkhPwQiQuzG9S60yF/BlrPU6A
qBu+BxLXRCPVM40nqIbnHqtPhWaFtCZ6p5SgE3UmPrGptTWP4gtEVnIy8U2U+kQaMI0uIrViHICH
99FxRkOo5Wcj1IB94yVJE68lwhtQTe6afHvHWMjOL9BFhmJ+3wiGGbe6DGlpBnHS2d4YzqFIR2JW
b3g29nIiTNe1rwRpDFrg69LYLM+JYBI8bYPZ88Q0kC5dVSxONG/+q4UDBeeXk/u/IDJ+4iUZKX8o
1U/0GJHtugMFJRBaOwftGr7eTXqTuutxEzAm5PROJBEjbzqUXgCh67ntC4+rSGG7FV+4k6+oDKZG
1vk8+fvlC/oW731t0BqtnUI36OnF77GAzTvSfcki6fqQkU+G2j/4bBvT1kDn65YmrVhkZbINLH3o
bWeUE4F7PPM8N9g1zugVyXvkztV/jHHh+UuJau9xDoWkHFmc6YettvuaykY+v4lKtIuN6Ap3cLwF
BqXA454hidfR5bASHkrdKyXz+a76zvyfkKtXH/YbZl25KRxLkuVq3L/lyeI4HOC+rWD6UORvlM/u
DmdAqli8MoIqTYYUqJTnPm8iKYlaY7bhLyphlt/3qCJZqWPrMUR6AGmBZsu3fOZDnxoOdG3+Wg2G
hIOZqz+cXy8v23Z2c96zACq/9EuHxW7M3pflwilQ7Sci6XWLhv1BDkTqicbWtDWFwEkNA5NoXMgK
jvrXFLcXy4u4GIRDZZaZhrh3T5K9Zdg0OTjWYRCYVt1LfIAlBrJs1TtAe7v/nb/Y/1boq2AIRt4y
c1MRbGp0Pl8e6MAH7gNoOgaaZGJMKAmH8JyCb5srDk1He0rT90PHbUGzyL77glUfTyWAkmw1iG0O
tZcPjE+rfZUfgYkn+FeBr2kh4yvgkNH+DMjIW/0qZecNo6vTjBt3Ri5Eh6R7MS7XuDWXpR8g0aju
JRIikIthxPxz1XpCWLNORN1ZpQaB/MTtcTEW/XMpyV6p887Ou59WpXWI8o9DHvfzhBJ7NykX7xtc
InvnZaIDunrecu47BcwegSQb+nqnccz9ZoqXRXIREUDedq7WUq2FvWbEewJkW6WJfb7hcRuhh1ku
001yI7fU+MDgGbBZBveGcRpKCL0FmZbhsQyc2ippHrS5QiGzdxpIhKAw9LjpKp4fjiBoUbjaNEcw
vscuW3I3qT/WE1F+euZAq1bQK2H3myGWWqMPC1hLWYThde+FFuGdQknt9O4Zl8ICBaExrsJqFXfo
Lhh9fzja1sVYvMQTHxEVqbPQkDEGFFKN72GOyB2kfI9KOXeTv+hfqwg3jzvumdZ2BOzhIvpgM48p
c6RO4b76UfWmFd/83ouj8wyIUXGEypssTu1Q8qkPIlEYB6pmQByZkMRiqNC7qjwqwJBhXN/bEc2W
4WksFxU1sofMd2OxOoHZ+Z4MH7dPiKhNL+nYzJdJCvMFyijVsawEh4SK/GmFRszjb1KaYfMmwMN4
ndW7abIJ1FlXGLKGr4gSH9SFjbZpItlYe8AK8zpnOYDvhKZs1Of0g7u3vmiABPHMdFm9IH9rALdW
qfcvHswuiDKcg0Q0FkNCHUVbkCZwwOue/whdEPySmI+hKHcEKixVoA6n7I5s2/tsApGy3q4e1Tt6
9+sYjUiVFo8DJk073f+mi5OAoiyUwEPRmGTJBpnl5AVcqCHjp8TYuU36jJiB5Zql4Ev1fLbhkk+q
vy2a+PM7ozHqwew9BmBYeF2E8oANNtyNgq0I+JfPw1ukmFOUsbWylEOmtJSWueiVGBnbed92FCfU
0yXR8yBxXAnMJ0ypqYOrkABSEiJAXkULig1dJdeorFf4DxiII5GHf9rH9HsUbZG9AaVl7ZPzFpZB
2C17XSbop7z/bUJ/5d1r9T3HCakzp+5gZLcSmLggC/5s1ugHAmZqprjsQ5woLBP09enejzOO5sMF
Vdvuxhkioiht2hBD8efyDXM0dlFJjUp4yYcdAJqslE8+213kFroigCISQVppOUTBMT0xT6qTKg6P
BVCpvXBbC1yUCf4LV+7WUPzzvV/r+xkHPw5Mg5SGUye3qQ76/jq5ya6Ie/22hxRHaAMc+6f/NLvq
ej9ToDdJ99vtdjYiYNCSnbseQqJy+V9EDjNFSsqA02h8YQ3fa2CYnaL1UCClq01VEj09JqoOCkg1
wLlsHKkeLBuxqqJwBUG6w0LRvZRhwYd9anc4jxuBiqLAaE7ce8wL0+BJHF1FA3e3fhdPadT0m09i
P6AHTHeBrsBiQJKp83NhiGW+Cp0JqnHi6M44U6atvA3GIZrx5yv/qUMj+8pbkkjlSCaS60NPt02z
2rG65YVs7/rko3j12JmAPtTm0ErIKjcOqIxIqlWts+NWifFP0ohD4x3/mDSra0Jj5icFuUOXmoDC
vFITCxR1P/UtUcm98eWIaJEqJ6nqtoui9QHGs/3er5QslNwxFdR8biPpsZ/h37mIpxm7RC7ShVrr
N19YScAgNRXJVjHvhr84s2gqCl0JLuX6TwQL1VNBqfXC0l5nUCKz25AMoHaip7w1gHLjI2uFGw0A
07eZ0KQN5/0XlWTv9yFxFZg32AXs9GJShbEYKLGTAZyp2KWIfO3qafVLeYnUb4WK6nB5TDtdrBbu
M98i3PxRU8CsrgIvazJbszu27nYYqFpeJIsdsN6rPIfyxkPJCyl9McJhHUtt58CUPUDBJSjXdgVF
hvsOPuKwqhhr7GK2me8480unARlyHBxXSC1BOsoT8PpBH4sz04wIDh2aVWseixgR35VxOuhnstmk
WZ4GlBf06W6UPc9hD/qqTGM7bLQtLQqM2iLp5iRgSN21nzOwCRHb8mrnMqBtS6WIgInYdhnJgmoi
+AGYwg8FaXtT79Fnv8E4d1k7vRgKOE3P8sxmAqAyRVPVVBmSE82wN40TXLDZvACSgKanq9A2wGIX
HFS/aHHDMSM1nurI/Q8GYom8wbbXrmIlXzxbntK8JaOj5oONODSWONf+WUfubtl9SeneGW1EI7SP
M9BYTXPOtgNWTeKvrXGGplgxrWBy5CVIvw4vTRTTkvEr9HLHLEhHSVOj2fZpgnsVbIFy+c+sVE4q
LAApXd+jZLR6QirfizZqKBwQcTrsVVTa5LXV/SwzdXBJcomwt3Y8BaYkfFlw6v+uUDf+cYBx3hoA
mD0rPQPWL3qmcOKdLQLj0kvS7NneC+KfQUvP4SmZK7zmeqlUFf41bCQ72I38ouorfxv+bVDWnweL
ETTJNqRHxkm3hLKaui7XrOgFNDsNixT0n3Gc7xmq+wTOVxX1Lpi+se399fYzqbPqT7kMet6IpJJo
X7TYr+qDDrIiBVKsNiI494nEen/Cl8+95j6jHUbGNv2DLU7d5iOtkUB/p2Tsj9X8ROyyqCUi9WFZ
qBfhn74pggJ4UGsf3vTDgy0FeP27FdE+Hi6Ycw02rqIhpRlNjYA3kvTMcPz1SYCoVAY2V8mzGJiw
v+y2vjt2FR+Gf4nIVCPib/sJJZGBF+N6C9r6pNgeiTEeYiT4FLuizf8fqGKjq1kstBTzQEsXvgy/
MuKAkHEfrZiioBDLfSaVptdqlp4B70GDmRU2rJ3suCFtPV0OGhmO97cEDu56SmI81AUxnkd3ehP4
BVeP3I7rpYDBgY/MFxfn4EQ+mWkX7wI+PtNmyjKVHe40IHCf2PcwrGPsPDx/pvc0fnH7fjOCWgfL
Jg2yVEfCCwc+5ruectjxogP+ylBxu0gDyYD6gGIroz/ADy/H40OqUWbXf1+29ZbeOI35JSEEOy1F
NZrqNpKXEofpnVYtyjkpVk4IEB6ppflP+wZa/M1jKqE+x1Fbhrn8rfg8ccrVIcf0iQlBT1tBQpmY
Xcs005/CjSPOwDO04bHxuJx3WTrd+3btK63+PxXy35SSFBcPKk/52I3Fm0lkjTm5MGJJ4DOAq+RS
aTIIRfMvh3mNhLvBmQ+HL8gXvWtFr/sBA++/X2DU8MxYQbZMAth0nmAKTxa4a7zG37r5LCPFrsGb
ZE9heMHtophn1MviqpADOvq0ude1M3udOANMkqqRsoyU2sZvl67B+bTjtZT+iktFsM6KigLESvm8
2hWTA2Go7qscSECpFQG0y8BztQkUIWNfOsh6SwmhAvqGKtjmBX8hPp3n8wW5cM0iXpG1V74h7rqs
bBKv3SRZxHHM27L91Gtf8mgZGf5udyYybMWk2pezCkfkuV7m2MDq9PjJyUi/LrKboSumZapjF4Ub
QF9ZaoAwOaJ4Fqh3pA+mFB0GELRAlEqRsEPnjD7uUKoJgl9KPxnTDr6klppspr1B2QXVYOvPsgOQ
sqelHE1pEkj8C72d62oPE/wFFBarGW8wxZLW7yfV0BbW0Em25T0OXDJhvp9eUDuB0O9dmPAmMi+H
DajhEsb/3NQT7inLm4SZRzyqRbXr05OT2X//W6zlNw7L4A4Znttl/sJ/6Yl0BUU/00Lz8tLCE9Jm
zhqzp/v/S46ewtVOtKDh47JqCPj4F/6kFJHk0Wsx/cakgBNCvvI91BCAZckzbnvGhQt2lEXnuiSH
IBZGrDSlRoc8vZOgfSmbLNKXOQZN2UQTvTpw1oro59pWupC6Rc42CQMvMfeJU2u0FxMgCkwEgLHQ
PAbr/S+M/ffaD/UPOq/cPPANmvA/xm+PBvtr9kBUXu6himEZiRWbJVgIPCZNk9+d7jGepPAaY0Pa
wsc9Y1pRO0mRmXlW02fUH16zHu6gThBSaK8d0oHiXj8njn34nnplydNochb4/PilzZlYjHKVpcQL
YiSEcLiyG6Bj0tvvKxN8WA9GGnh30BJYT42LuqGmUNVaZeHBhvdxIvJXe4piuY66hkRODOnoIWEn
tAciW1furpXdaKohHSZm7ZWEfTGMSZ/hF+MdZg7F1gQHEHMrkHpv2QENKQCQi7ckKhihaQ1J8YT2
vXSWEiLTVy7KwMpdfzPjNnbcA3HRrel6Sf8XtQj1SDVymtGLLIw0zBxmpfbrUMshloa+kvnHoGlb
LcSG5CBWLDupvG+27NwtzjatMOH6xx6WUJ2EC7MIM9D823p3xWzztBqddunPS4wrtgc6bxGuHnz9
nv7m5tA7txyaQL12+g2mj2itxj6bRuT3gJIz+b89MZr4W30POqp+o6A5batLrdMhBR3WpC3xc7Fs
+zJ3asksNPlfZQ3YBN+/+fOfYmXF2ESx8vADWbqbMbqZw05hJx1n3WYm+o7MIMtNUoESRBu6vP31
KdXv/B3bn5ZPkxx9Mh6wlI7L/qO3unoramvTZEy3G+rnKVDJ9G6MZm+BfMGRO/gEZWm0dMuSI/lL
3ykrWOIuauioGCwPxKovmsLSc+xiGsYEEmjPjFEEL4Ggl3Edcv+N3SFC5ClE3LXNopYA9PdV9jNr
WubNoEseu56CDVWoKinmWJsJE+0Ep6fG6ZVIW2MXfciWt+k5R4HPAYxB6ctkUtCm9blhRpU9/TBZ
LLAfwyB9zQ7nkNHRKTfBm5yjpD5XN6zU902tmIM3oRo1lSGdkONK5k7hn0BZHdXXbsdDTfxvfANX
w4CPo6ZMXcVUhHXa1JrelShEmEtPoftg3hCoEsi/uFcBOgH6tTplI188jMsYwLw/6HzAwavNBz5q
/iu26tSy0BzjhKZf3njL7ARJML2JRrj/2kArc4TVkCTGvjdTNGorI/dvfBzWjhSFokJtw+QMd2Q8
id46Lkh7tPb5zjRv0lMSui/zsTPReTSIThI4BBhsQ09cJ+5obHyAbifgAp4BN/VLufABT7n0/3wz
d9UBMgShiVA8mmHkX/bgtkj5eXtIN+YyKqqG5CKq5GBQeUSNDlaAgrMEEJ6mI/SwQQXmkkSBiFc4
9xpjV3hlVMn53+8ub+OucyXFaeq1U5vq6Kd0ejpOZaJKkY1oziKxbsStvsNG4Az+zAfKsymCSJgz
mTPVdDkWn32+FpouLGZYXDXMu4YypI+bqNEL2PdCMbCR4O/JJR+pqn1NpneA3lcFmqID9d3zI2Xk
Fh/vDDCop4SSrSNojYhJJ5mgSPXsyfeMTS3VI7PBrFooa8vg3tiKVWolxlp67r5TLoc0B4vpn6y7
3ifd48ydueFK2WzXaokUc5TNPZK0YcdWJ8dKF6G/sP74fcrDTpvqF1ov1F7zvACrUA2yet3ffyjb
a4Kn02aMEP5uoo+GXMsHfaJ7ETr72ErdVV7VUUWUK2w0PYco3DytXzsmd/f7rrnPXgkS7MGo+k1c
whUrRr7ERsfIGLrLGt47nhtAYyTrGPVteF9KPAEbOl4PJBnQK3apNmquR/eMJ9TQA9F+Mf6DOrKn
LZNczHFHtrkyczVzPqZ885T1T5L4vynhKEjoNrz/6yf1pABbs8kntF1TIkEEFQhT5QWMz6T3YR1O
ksZXtDPVR0a/CcXD/BaOJ1gTa3ClTUwQMm79jlU6O+k4uzG1xo0XwEytq6aBq9V+oDTBKFO+oeFQ
XeCpazafIP2Mo8RSX2HtUMKggsMgxUMOgym42znuUO66PsZBqLVmRMh0UCPuZZ6GyDdZRXXpRH72
uPNECFUuwvexjb/rkcQpeEHuxwCD9zvglXCaa44FfpXOPMPOREFxhGYt3p2yfiPBaKLbZ9L//aqK
hVzzms+GNNdpcSU2UdOmDL+G8OhyDfJ1YwnTAVCI5GWQTdbUYASVWlybP+JEvRtoyfutfs47+lCw
eKRd6Xeo9YHQ9heQWhv94xFgfhyD+99fgpWvpcwr0uMxZvPehwHROqvbchiPT2nr69xXAz1v9HVe
6pjM6lqLEMNjxnnL1n4Uwey/eJPDJN6qmag+uZhIkGCdJ9m810M1t8rgODHEBUQ5Lu9QOs8WlkAx
lMfuBp2uLOe0jit4DV+TyKMfmrO8Rf10/grEhsWS1ipdOeErNEoVYcozhA/3ASKh+vxyWUoq7GbN
UE71RGziNVstE00SkaGSFmXwNq6Mxa9iabUc5kEM+JMOj/2f1bzTmIpLzSr/Rj0GPd7mJoPQbi/r
xAW6iBKExUl4sOGpLj4YTJYF3ExjquX0iiR0V4VM7xhf/qVyYXsC1NWkp7GEikyEWxREag3sm1iJ
lTWtx4YywsmdFVQR9LyeqPjJXyVNzQKHFJ341nxklOXxzjfZWV9FeyRZap0N6EzMPQlQnX9ccs6Z
OSdIu2/1Wvtj4pNrxoV2lGirdQlBNxkU7QiAbhVn608+j7D1zXPGDbwv3WcLopHl+qXP6949ppL0
rLLaqAuZi973TCiEYEPTSETBCkCJfpYLH1uaeN3zR59c7ipTNGeK8xd9EhtJL9B2uujHqnIszKNN
jPVSN4lhvF5Scob+LsTT6e3UkPb5PhqLmdHwTNm8gxq+vdIZeHBkMu8Bah8AsYTrG1p38xP62X+8
/aQTT/KV/blnm2bVcpDyIP/UB7r7I0I/V2T3H6WouzfXswCCAxIgjtftPhClTjjv7ZHMBUjRZCV3
+jGxclp+WWNm259WFOEXB77jmItvtUiEf1OmF/Xf0lEtj5HYBiP7VMXR9tmvh7DGLCW6RtfJScxc
CvyNvMCDN/APvwiXsrA31spWGtl0s5DEHiSIJNQD53yKRgXQ7WGKEBfREK2/s5VMORJcM5p4kfKj
93FR0QPpEZ19ruQIIQsr5cNhbMhdhjfUIfjqmkV5KwtSEJcilsKqI6Gthv2MUnVGeb6nnU5R8uy/
Ry46/dni57AFDrSB551N7TbB/WK/LiWSADksbm69v8qT/x05SYDScy85g3BEiPyYbDs/mdlh0185
V+cuL6SxdA1HCvhtFU0PYthneiU9EO0N02udVRrOg3RCWPvt0zgiFYln6xThkwIPUH/yE6hZ9wbi
Dibsi8oRG+VL5HTR3LJAkjnxOi/bj4oXOOAJMt6/z/zQj7mK0aZbSP4A7SyxSrFcILYHQ7GKrfXl
JF6HoVtd66wRyoqp5Old0Iavb9mTjK+yqzfWN7JiePYAeqbbJWJ1nuOsYyj6KkXIOHJdgPhhxl8y
CjObnF5vmS7bu6aN5tpn3La7spW5sKsep0LeWe4k44/MqEDvH5s+Pr+1AfZMP/RgAaJUuJcIiQlH
c+w9XIYx/wRJ31ObrxkGpZ/KW+cMXQdO/TTGim+JFhwWHSuJngiCxewi+PFR/QRyqxTZoeZoe1H7
diuLxAyJA/x0toj2tWx+QTueRvd5xVPju48bDkL0TiNIBczizHvmqgASnQw3dopCprr587p2YoWj
poWauedxVVrJxB2Z5OpjkwzxJSnUTUjRDv0OwMiBZOfoMhrX4cmvjplGgtR1unCzAYv0uVdY7eTD
eQzzNhr9zrRWIMt9B4bHpfjDPB6wV8ABgZNnSvxPaFD0WATyxmjOUHsBAcvqN7N8NMKNhNj8hNJr
yqVdNATrLtGE+djQByM9j/KpgH7gYtVhPePV/TkZ6QD4PiJK80KvFJRTg8P5+kSsRZL1Ym6t0Q98
+iXmOaVRa8IeeTYpoBafV4lhXnrD8wYbNFckU1kFk8uIU4bt3uRM7aQ4QmPyjfoSI5OMdi+VlcpF
bHzEY/24lDCV7kZgX96LXH08CycULuMjgw56K8SjQXPYCrBSUpViPEa2qx6RgxGJboL5Z4/hquaM
p8CtdI9CrFKJyDojG9aDFiNMOVmskl59A1FLXdHLDhE5L3zSARPb+n1wUI5eWIwnP0OQHv5HfO/d
I3nfkY/F1fKrPtuZSnuw4sIzKJpdeE0qEtgLNdFY2608tkt7n7LUeLTFlqHi6qmrFhSqkEsYAmVq
qAZkIcAgpQ4W0HUnibj5pgQDd1RKLfM2N+7B19X8vWtn+jF0T2zcCK3yefUWfURisEq/c3GrJ5Df
FBUQdjS6bYEywQUdrMVogHPERGOytjSIH6eNzgL98lOP9o9SGVfyMbKWpUcIEyGskhBvw2gEDG2D
KyHogLZ1VXzewmk9QIbldhe1lIeXK3jmAATI047Mj3QJVatpLlBskG+G/+0auQ6JFzb7uiDj1hbB
xbo3JdspOm9LdQnFwBC/I21MHxM/yi7dBfATkUKnS5/oobYFeIIRNzdoX+rSZyvMWXQV288tCuL2
yUxCO0u1Lx/E4r5yxOiyzu822tmOx+NUKo3Pi/XV2oHKmWf6ZzZQL8k9ACHUGIDnogiT3lFcqgvr
0CjhJ1bWBFF7HJahOn43UomBxF/rUyN4JNP/tW+AiF8F5Hs727UAypNiopC/WzSRnRO9ZbT0k34F
y5TAEzcNwM6QfXD6DIFQjxrq2UTePDK5y5juIWvs1uNu2FtVEKsMnEDDYwN7sL3PXum3Yl4B3IXn
vxERLqJ1YiXRaNPw5qOSJj8oqCA0K4mED6x8kFQFafBwHohFtxxr+QFs8cWmG0UI4x44PvIVRXkQ
oGYYk6v4Q20N/W2Bqxnv0iMCRmTUmh1qFdhbDa5iFq60AavlaK5rGOsdfuu3L7WcLa6jpXAN+oi2
OmnVjSvf7CCfnbYxWWSUQ1B75RLjf0+aMagFl3vGs/FDqQAn1CLzGY4/4wuxvqX/c8XQPfS0mUuX
YEmUxVSoVDQyyOs4l4OcncfS1Kh9Ciekpy8yGSOW+2RK17y4VViFEbC/TOEonRz+J/A82qnHWqjp
VQNyhSN4SCKeFndxJlOXAlGL3aeB8HVNkK4uLH5sz14d3Hb7q0f38BAQVC3wC5zeuhMfkQKYnenJ
Qd9Vq0oYS1A28+8M2IJ8Oaw97BdNjFnbiRQbbuFY0T5jt56hsECUkA+PWb5w1xe6mP08amwwmuBP
oxucNhi5bdTN6W8RXYbfixLrAx+rfVSX23WoZ/q07T1Txp7jxBj6DgZxnisDTumO2HIeVkGck+EZ
MJgaHcWmpbT41zwQkdZjnAzcyv19U+6hUEbo3wLZb0ptSt+3izJdTIKNSaJPAMJl34sn5ZX+8x2C
Vkh5N9bW5qw3wjSVPNYnTCQwXGqlDWhGOxHmnJ7oYP7pIwc6H/Tcgy6PlMKUV1li48Gwgxnr1ie0
rv2FKY6Puc8Ssfi0WNNTO9kHT9v2udIQnMx1wZ26kqEx3oNvAepzVGu6JpDJCscyePB9uJGWTXJ3
fbOdogQQGbUUH+bp4IiO5uJIKi5fABr3WjoYoyUKeceBaV3zZZTaiXNblhS/L8VTaxUqFVKq1wvs
3HIWm2wkh9kJZSHw/RKTr31AYp0+ic/jisq+rvqC64TOibxBZn56gcBaT4HwN51NXqVobGHadAga
obtvtQpJc51RHl6wi4peMOmNfLmoeqRCgLICqVxRURLBhx0/pnhFhIxZKWQEKMzXcEKf2jDFOurN
ynjlW5O7dCFjVrpJKpnfZLSUFiTFeKO6wG7l1y2+5I14sp7DYJL5iwG4NRh4EB2nCYF+zWreKBd4
d1Z6hyUMMj6QM77R2FdVpIxBwngAPMs4QTBbRPtoFXlvAO2aBbFBe3nkelb8Pl4F/sxesDxObCco
7muq2aC1mf1+zPx10zPuqBcaFj+O/YJPJuZJg0fbxFckNsGeqPy3bSJZvU+ekPQSofYPUokuz+1I
EteRgs6iNcR6dq+bG7TRvps639UgFLfNZDPSfSZDLX38N/8CvCWo2fXpsDSseGwYzuZTbA3nOMl5
M4yNen6DUxU02JcnULg6b+U3+T2jXYlx4kdtlYaarF/pmPdWThGUp60jaWGM+gRAdLs7XNHEMyJw
tu0HR1e3gKbE667eFAOJ2ODCyLqZlTAPLlnK2RkFNxlTK90DGsDFv9XjrHI2JF5XJ0W5qzufP9op
OxRC3J39twd++ndR8KlxSyl+0opfqI4UsR8cb0oZGzrIu4NNpNg3J1/+zjFvr2g4L4LoyscCcE+X
4T5lJlKwbQq3A9M90/b48poiQoYstrHWWDvxIwUTDkaVP8Edf4WcLOVr1hVUX4LwDDVRadUGGXc5
CWJDDQCAcWp4ADaiAp/KJk1M5zmutm0eZIKpfBQNWVljoR59oxY1LmKv0Xf8JWNo/Z95YqgAgSoQ
a9cLLF30vNSYx3AMstXVtPi+3bpCncxliZJ4POROykbxhYy7T+92hnIWgivIrHEkECYcFUam4ryQ
Eh6jp6t5Xk4mH/CFFqMuKgSlMETEqa3eVPTu7xO9wNuh53JHrBQ1iyTXeEMDBml6c09L9rhp/2bo
j8wk8ZVmJpIS/4R0XDdb4C2LPW1GaL+yhQNZimbgEWfkLkATQUxDTRLfuoeboarf/KwqNgxtJ+By
seyeJNy1fSW3k4EwBRUuCv86RFdzFvBnvelkJoTs/2nJHJlbBQKaV//T79UvilyttlEG0BIUhPOR
uVeD5ECp/mkMsBO69ZNGk677+C3M7dbBmMjQ9ii2uIVSAAUEVeAPoktHSBUymaY9XjjR0Q3PRjXQ
bDjCjXjlJotsNRHzanjs6A6VNLfVBMMJxAuK1x7GAzKFh7s5tUT0d/SzdyNlRkh1YQ9kyIAq++Vw
1WeFnZAibeLIwS3KSfjrjGxb8bLTxIbPua0YXipxh+2dZNDATJ1ResefefhxvcXxNG6hqjftcuKl
2l7XEVuttB2a7wC/+UotJTi+HlELPhYcJrSfaR6dM46+8CWqiwZuTbS3xQWNsKo2npxwDNsxP9e1
bgylG1rsBQsMO9H57p5Z2RQiKCmxs3w3Z7a/40X/8P0bkc6h9EYPAXb81GIHYsEH1tuhp8iFcDDL
hkvnW7azRmb87PFNA7MW+IhPSYXzcwbrm0TT35xMjVQqI07YBSlcH5NyDiOXNQuQ7RkA7rxS4RnY
VKHxA3ThquHOlJVa+055EuZ8FRm57wf+h9nok9lNKeN027ao/wcg53JnE9CDSgxxPucIADJ1vFri
Dj+EWw1DH6c8NP/a74TvX6wRKzw4QljSzPfr4qfqKFODW4ZPYgPAZWPLroTQJk12C3HE8q3Pe9bQ
VCRWI2Hl3immvVFOVdfHpOXIetlUBuBl6VDnQPFFBKKfsSKVxSr7yAXaIHavDrVUlmKODIc7pQaW
RAVmPej5ytxGC8ZSHzGBxoJGbqTfafrzJ9VbKlOw3gArxdiMkGOa1Pl6Hdhdt6S2/ZvCkRGf2E5+
3o5ktm1RrpzphRzqh0c8wb3bcqNWVf02B4azSoyA+WqxTi1tiYv1G/9kUOKsbSf0XDEHnbaE5jdf
ltmjNx428ptWcgdj13qnpxF42P5Td+m7lAlXa05mVJ2EGAoNMc44hRuuN4Qc+Hz2z27JGJs9Ezby
I1O15wdq/bOheDZFubqhMzeC+oSQ0HBNp4Wrj+ZvRV0GjXNCI7+6qorGLVp95WGLujsJq2YEXRBX
fJD+Z0gI0eOgdUI0jmw7QilkxSO1pZCFcO0ZCfQlEpIHlTks4/phECVQ4uw6TjaAmZXobijfmDZR
3LePUPRlXVOQpSSi3kSes6EKNz3jLUKTJyRIVSeEQfAq90BfgeP0uwJbBum1KslXeLIIBoCC0sSn
mTaCtFbzyqADmoe0jQZhdXncE00LE93r/COYT4ZP7uxWA81G1+9Hiqm4Eh2eZAjotaeWKaqSHxpY
RgloJGHdyQLRGp9ifhJFd8wL0seviFis3NKg9FxXQ3Yhtvlqwc2fzyQCazcNP+NdtDM4oVcxF0vP
5FSd1oQr7k/mP/tm+r9jRVWjaNsTsRWnSNUPEKtoyf4k9U3b1C4SRcV8amdOwGXCkg4VuX/HUF1M
sGYVs3LUMWR7McItCBQB1HFLekERBEM4WEY4peY/ZO7Nnq0UM9JBhSINDYKTOkcrYSKmVdQxTrph
wE5qkLIlE54gqnOuo31XY/IX7AEObYV1XCXoHccfX763jwgg+b1jEvrfw1t2maSn8HfoUn3oGDcw
RIPRPHSBqLNDEmUt5Utv0a6ugUA79L424nOqWJA87e6WR96k9W4B3nK8FrCT4P2DAdi1huXVQO4N
T1BB7aT1dS9P4Pg3x6NEmaploJ7583VGj15PCIBZUeSfCH2mrhXH1tN0sj3pLoPAcuQLUExyhMx/
g+qoNbd70yznTMfjyebQTbH3ZJEuiOmK4jNc7NfuOM/4U6iW2Nc9P+ZqM49S/jXY1yeoTilFyW/p
OJJK8LLruTn+eGvSMQBX2aPKShFnjV5R7JqiZaPJsE0aLpTR849UfbygNAr5+a0YJy1vYOCGMo07
WWRsh7mj7NdsdOSbPcuI/Bu/G8GiaEt0Ml22MzPkPX8P6ZLH72e9u6iNYZXbTLii/6pmsNzZCg9d
Dyst2wTmD8QTzn9/AUrHljqPML1pktmA37p3qHky1LLrF26DtSdLDCLzWafIlzvIm10C84liS8Pz
j+YB0eOc62p42k/BH7xgk6wVTaxC810qhNk9ViX+C6uEOC9/OxrNR5TiXsGQiRhoYMf5YYaXwLUk
7lY/n2UL+LYtuczdtZqA5IqyzqTwaWjlpt/Ax7df5Z8bj29l3qnF6hlR5iHEd37+VKteywMTAoUM
MC0B1nDi9N+G0WpOPa9tg6UDQytFUEoPq5rQOghv38RKt/U3arEG6bYbbdX8tJ9gVSUMGRqd8tVP
NKmkVl8iofJ1SY5jbz+d6ISeJVW/o0QZNdQKB8SLs0Q8qnUVOCdEtmyJbGNls3jSiwVTwkj148oj
JIoUHWkpzChrmnOkCDxlSQa/jEncCCIwnkFIT550IUO66Rdfiqm5O8u+K9z3/QqRdN3kgR+aunG+
cjN/nQDKvOu9iUcT4wHPnvlBQVUw8KxtGuHs5mvGDfJlUkzQxUlss6PoPtoXFku7dzXM9OMFznaE
Qs646qAKdDVGMhNzwJnbpU05uCfCnHzHMY7lXBi82GfeO9sC1TmchrFSj2D+un6mFtoBMNOvvTcv
OxFewXRA5pCXiyKr1q45MX1rma2ThwyrGyhmF/PmhL/jWcLByyspUp4+g8EdUiIJqXWWljnC53Iq
m89Q/N66OyW7CYgX5lEEIIuUBGP9NO+Tx0S4HdzfTregoF3ue3lngEgETYtH5lqUOoxE67OqA15M
iwB2UdgsJpqY2+jXR/c3MUp59EHnHu1k8vPctSNJ7mw7ONZoQiPqUhM2ilDDnJ0g3tV7mIKLHnNo
Mq5jOvIQUIx1NkCE/ang5Gpso8+2kgePbQbLtu75TKj3hsVIqFO/HvGoG1HyYDXXCURdVx3bSuui
bfMA/Fl6rDb95oozsM5vk32TGxjYoThe2D4qaOy6EO9osCjur8hKXcGoSF3zrIVwXxkUQZfGg55w
0xF03dia2eLx6GF9VHXrbSMnalrug4I22gBhVB4Z55Ue0ldFyHfLoW1aWjdRFoqTvFBe3VOhOsTP
ur+lHY/jFJc4znc8Jy1AuBucnciHGQh23tCJlWTJwvMXiWTqdjh5ADfKO0VIjsCjbA12pUt/k7F3
AK/t4/NMCAtezjFCTF65N2Tce5YjQE8DH2AkqN0LFJT735satDlI0+v2id66cZ9Y0EsI9hG15uZK
9Lx88niSaeYoNjZWsDzWahTRbLukEx104xFUjKsDrTngQlLduFHL+2BnjirBVfugFwwFUFcFRPAN
pKHWRBzjHOsPdeaj0QF3YrAOHcByTaLYRqca0etiz1ADludc2Vw4NRkUcce2EC5Wm7p4cl5g/rlM
PmpCFBcsmlIG7L0dWZQXQUlZhHOP7Niws1fWLCkfTCCVVSWYiXR9bSvXkSfN/LdPEvsDPKCjEy2t
bV11hbkjBG/p4MpH89gizCEGY5SaVkX2OZZkC/5Bpq3TZsr1MuSvSFd6uoTOMS2zS1S8E3C8uzIz
XjT41Z8GtQ4xJAzcRVOnzP4On9wVTsC7tQKXuNLbCwE0wGmjy+NgC4wFC2UvP0SMswxNvWZ58RHk
ZRYVreIOsxc47WuZyJd/x4JINtu+6anO8Mq9RUFlW2LpfG+bXVqVhYucjyWXIAh+IKrDwgT/j8q0
jaS16bKsH8vOOyYvhZOOh4TBIXZ4auOpXQ4f40K70lCsDsX6OGfyYE+pnSar68R1RU+9E1cGcFsl
lh3yZ/s/0snUycOHEY1V1TTao1IX8w1yppj6nLxwMol9aJa3IfjYy+AjR3WxHk17h1i6aqNAgGGv
NAcrNntw0MM4UTVQBUVZ628XMkFfgSjs8K9kpsSE0V9Wal4Wc7WUs0O62WtplgP8PYiP/5T/4UZA
tgrSVz+JqWKY87GHgbX0cGuRWpVIuE4Mz8PISEFwxziioa0QESaXlv5/8HnheYsPKrPvHx95OjMx
OTy211+NUgFU+ix2yiC3i+spxUURmsfAXmbobDkQZ5YVeTxvbPHiagHLB5/Riww9R1X8mk+IDYVE
gFjXpFzdmIc0CdwBFlXyhXZtHMYzTIityZh2iFr4Z9MVnDsxPrl58qWMNKBJmvQS95VCwoRxitPV
A05XpcvKLljo9z24cu0oiGQNPngsyQGTrdJCiUDRaFQcNQ0A5PjunCfb3Ez0cz3GA5PHA8BSbmQb
4xRZWitr30RzZKSfb1D5XmXNAXpn/wIWnbivZ0lA55TuJ0J2OT1CSUE86jWv7/HgZJtn0bmOAEJE
MLOTcSEvvpaYTA2RG+h9/KF26qpu/RQIu0ryAwtoRBmtxS5JtoVyXN24QhQd+mtvYvdAbigP/Y1g
RPZjQVzefzn2BjxMmAM4rvRUmS0mKTNy57B0SSUhKPwo1HITrQTbnXLgQHIXyZE5hVbuQAzK2P/h
xwhpaeZMyxC7jF/qvtnjRvwAc8qgC+iC4J+o2lkrYmICuYYXiv7SdcnXxDks6cETYbFTwrgJJvuf
yM4XkQHj4bY7H07PcpA+JBMfDYaUuP/0N2ouk0ZRcWZuIPwC4WY1i+zgYHs2TdZm8oprvsrUzcya
1i/CcAkWbIrvVZrd4fgnQh9yXIaBfOmQyCzgRWn9e6zA4nGOWPGjx+ED7pSSnMzYJwntD1JjCjJX
SjZsMHgcmIAmjmMrA5f+mbKH9zoG0wD+E49giH6snCObuyzCUAbOVQ2BatNgD27K8oJjaOo6eB6U
zCSQGf74930ixj1+wQB0IaEaGigeUPAArK+oz7wWa7n59WYm8EdRa82snXi486s4j9BSk5x4430A
FF+9RGM2OoyXPle4TaWCD8a/8Iodux/dXq1cRyA3gWE/wjhW97s7CKWc5zR8wzxNU8bsHqf6y6Xz
bErqSgFDSlfUgg3QM2Ej80VTR9BJTNFaeyEd9KhSuj5c9UqiRekmvCbEeWu+yiG3DpPDJDo4KUu0
e9S0flJcqwPpwQsTFSdBt63xMc0wud4Vr5DFHi1juNeezShjmBuFWF4+p9VHawTjtRbbmgdNDR96
lAXTaHa6iTaZ43+Y87TiOpHUvk2+4OJSDVrZ1O7k544QX1qbFcwZqIA8/1/1yR+thWHOGsBkmS0/
FPXWvqLtB8CEZnbnlYo+/O8CYe3y4pcg11tG0QtyBuQAJYZapyhntoZDvE/MTHPr15QjiXLT/OPF
O/2cjGBi6S96e9uRrlfe2OuSVrpw8Vp0GhVXw6i6X0J/IFR7a2nfWeNpJmeJ+gVOa5/R23/1108/
Iaa387/EpmGoRZ3SXQyriqZmgv2PTrYNaagwmz42S39pU1c9Juaf3iFSQ1PGTNmkM0aE2omsfPXT
1/742tV/0WyJnH9P4yj8YLxtEig4ELEfQMoPDzskiqBFVqKhqt5DRtrQlNkThy/vTKIuU/mADYyz
9ckxiGVC3pmciBnvsnzYoykvDSiqhcGu1jTpna0fBS7MICfDujIw9425zear42b/gjEn0EOH3+Gj
3+nUygRhWqHcaO6yV0o4vRVbAgX5KHL28b+s/NVfSni7OlEDreH7Kc7mLMhDxhYexYomnuq0sxTv
UB23DylX+jpnkzxf71qGNisC5OPCWTd0DMXmvgR0FqtMQA6tqU26SpD33hDrcUvOWPz4hfXfUIms
SuE10afm3ijmbG0rvXiP4BlVhBbHj3G+0NC9BDIg6NvBizdJrPjAwrAg4tfnyaog0/JKgrBH08Yg
O75QKAxBZkfvHoM+OEd7cDHy8VScTDUvkNjLoHmdKjdMZy6puSIdpVdRrbHg4LUlE03YBofUPj72
+T+oeyxV5gmeL0BvBuxtA/ZWCHGtUXQOyMbyk9k8pchCCwJIyU1Of8hE6zDYx5QLS+FENANLlnfE
ck0zc3plEElPHIX1UkbS9SrlvLEJ3krEJTRn7Wy0sIsi55jWlkzS0dMM6yV+IkGvsJxCz+bAFn4M
/GYPKzMpt0VN4eROg8a/x3ROoY/74XdG5QqyHCRo5/wDNttYx8rCSbBJd0f5HlOLyE2/a+Hqzs8H
zY8mIvj6fZNQ7b1mAohDDz81KtywBws+f0Mpg4IfTJ8Ap0hEwhSM1nFX8cD/5AwcKK5ZXoiTX3XY
ZXsAyA/g58prn8GXaZbH4q0bm+vDNU7wy7Ajc6gwt8dgyn7oJL94Sy6dJusAS/dvQhM5dXUvuvgc
nLJictxoBOtLR06ec5aKdmS9Xh4HMlOWqU1VxSu6Ehd4v3UY0RO2pKxIRW45wpmHbskuiqeupkmt
dqOcAqG4NEmzIIeTWkyME0RGNDZ/xZkTliBt4lJML+csShai3Q4/ByfoBrKi5hr+FYaxQf0K/taf
g0s56tJD2BD0QeoPsPSLDjn7ghQif/rSlQBNwUZQ0Qh6AqHgEvUZyP2kHRfIOvKAonZLrl3KK/wP
sO57rb13DKCE1Y0uXXmOCQY31kTq4Thp+E4s7l2h+gkaghUuUpKxPJnyjP+q+5Ge6JgyxdREt/xF
NfZNORVdEuBQVmJO2jH6vzg6tHo7yKdJ2jbaAlScb0az7qeZWipEoFO8pDg7wuOAjRr3DDwxEU5g
kPXHNA7/jTktYyK74rSxQmYRKCZv2kvA0AhvUF54fnR0zSh5+6zLYt6mf2gR0ANWn2Mvne9peDSd
HpQ9NhyNU3/dwACaMPnfJbEIKhD8QlRYFGT/cdnwGWBX5VCFG/JZsKwEhIebYoPdugYj5G+GojJl
yC0rZam7XecIbfbYRWiRzM0egoPwVUEIPS83Vtg7dY6LN9ycrhfOn+sHFgXzoU/SGBrBeK9Tc94K
xR5Y9233njYxb8uu0b/I6G7LpyScfZHWSBq7ID6mODOx8lRisMVF4DOh6kBJ1uLxZba79GuLRtNh
f9Uq6VvBw7sE9HDo2jVv0Lcy3RZMNeHG8Td9NODvZ3WHzm0H4sOnP2XTyK9c3FUZRFn7VYEPXkKu
pDeOUcn2v42oJsLjMN52Juh12pJs7gs5Ol3UKW3urZ5eKjQ8k6Jvy1NrfZKxCdqN9S9dCZjUZXwI
sH+kJQk2B5bG/CV4ppYitWKq1lQ6kFiV+hGq9WQHkWn5I2J+9PgGP+Ay/1xH0KhQp9c41Kyll2X4
3bas2gnzTPJ32AJXmwWNToEvZLlbtHXvmsB270iw1CLtF8m9P8dUDI5uHd9Opc8CMr9SCrTCp7XR
Sm6R/wbeIsPSHJX8JXFBzmeWUqBIP9FPdow/Zc6m8i6898ck7l5x6Xt2/EqZoa2SFj5xkhwZ1Que
XsJChx8F7yhDOeZ42y8Eqs3LMLuoWG55pMFN0UlymOf5ehOtPm5XBliSSWH8FPoBp8Gpq6mX5lDM
nEqvqEysufv+WrOD0zp73Oo9V50sSDhc+NqjvcLOXntXs9Q6rH0CNLZ+hamJhcdChKXFrPcxlzXS
N7jtUsUbgHRMWwz/0yqDaOnWT/DQQAlXymyUEeoS9hJWXXeFtrPZeVcnY5EaecvTFwHcbaXTxsWK
fhH7mNqjNvXwIF0kaaHkvTm4umNA5tGBCHcnRaKLcSXKiAPVegNDBBpQXO5AYq413VotvFtmfUPK
WuhlDErSEPve+eZsdwFEYBedKNTIosuvwn+geYFsWcSo6CEW2taKH0/4FrDwCyDjwPmfkXXRwuOQ
R3Pi9eUOv05F23rCHQVtjwsdYOvfNkDv1gciWAVd05jE7p1J+HC1xWOYOLPQMYpYorGGhiu025vX
J2PKe7CN0CENVLjxeHe/qayEpyiWdDAqZAoRuUB3P5mYEPI4DLOSsiFwqEdQTkP2YGW54bMUqtnl
tTXXKB2GOaS1J3HGFKIOmljvhqQsN/fNN2fD2tLsvMzQHpO/qaB9+HcLYL3DfCTFInXEB+XYVlOk
l6k4N6QzWoBZ/dz6gWokbT8U/sg6tsfHpDxQaI7HD+rxV9u/pW1M1vm1oVOWGyeGS4oqTYjNfs7f
0MW2CQzLDdy7Ur69JlBmfmhcVkWk+aIrUj28D2x7erbNju9m2nT9AGiI1hZZ/aRKbX/UIO7G2ugh
5VkZRcQGzpDo45qdoR/3LhbCB/LbwHT/3a5BMTyB3NtkZurFcx6D+XnEbToUNjkKWFLKKyv89EyN
hubRsJQKlW1RCL/+LD8NQ27BCd0NmxxE/144GptyvFCfgPEebHH/hFhd0t3lJL3fml9JszFnma14
gb2L7Rrc/04KTAI+4KA6Iy035g94WOCB6YrQv7njza64iQDaXF0rvVrBeLsVLa6w12LCGGC4dJfm
JeuiZW0PqUF3+wvIuQQULZBy6+M0Bu5cNLLSDWxIGEmViiajKK/s0mEqHFxJBzIjdWnlKicJYDZ5
5xgp6Ko4bRKW/c9V51zickC8Ff4LfHrOFt3A4m0HyUkEyOf8PZ1tk+pr3CuvxX9b0e9Ru1VinxlZ
F8GiAoZijgQ4Px2LHezIYdkI3/51UUJXgDqasKbh2d08WqqiFU8GN6bUiemoMEuENpXUZFV7wWnh
Z7br6uREZ1FLtaE+5a3qd3S48wHFDYxC8rnpM3/wuw9pRw/fBtKtRdoDUEQcicc4E9oEHbv+Bipk
5/WvJ1x1sRUsbaKS7yDtyk5Q00+ygCdfBy60MZLTInQO51a8nvisaSN5D5yfrSJi3GAOOZSJok3W
hTmvY/LQBGxmLH+0z5aPb/lU2XAZ10bD+SwsIB1gTRhWWaMYT/IL6+MTrQp0ZXg3ixvXSbY55pYU
64Cxa/EW7yJ4BFw3tPZs1dEs3qu8HvdTxIUjpW6NkmQMpI2GYnBLoaV7ZoP1+d2RO34isvTU9Yj8
9CSvJFhcw9leaygIJtNA9PFJVjGeIHxUksO/t+PZyt+MWVICARwAKgvnMqAwCSgEMHsE/bIydSlX
Yu4Orh7B+c30L/FL5iteJHo4ckC8tbQnuNpJHrZEzsfqXj1vYuoKuvX3S8HFbo6/AleHb8NDAdub
XWEYJJItXqDiyl9po2T69flCXF5QOPfO9wrvQKBUrAk0G5GQSka5mHjzwCrOtoeTd5ae5Au2+xww
3zfMNz6ELjR2yjNMrZyxTcPlOyfRgUKwIfdJoTLDObyD4Ek0v3xHOb2u2kNfS3orODBzJAlJkYW0
EXwuKF5Vu/3otbiJ0P4bxAfLg90CubnaWxW4dJz6+6Q4A5q4Ckj5Jcp35bvi0ZPPD1udUpqVUhYs
6EG6++2Zj+nCGlqIXKlXuPWwKZvO7SCtPDJuHU8zG6fl7fdO2l9ZtnZrw6tJ+D8v8imdV5DUHMvL
CSfXJkG3om49tL+fTbp1TKvFROJhE5GOQR7pOkl+ALcg9vIRSeRskYK568272DlaSpb/k36ON8HN
GR6MrD0aqxdPCoIelIKtl5PIQGRO3Draxam5OQfiwioNrAIS2WTkwlAnrc6ByP9/ejbjViK7fQ4o
PYQLwYvYTrgaQJtob+eSgBN23btptZTtIICgt8Yw4mDg8X0ZrxOXEivQxS27EbJ1UDVDTo0d2dP3
tosWnQg7eaD6owQYdH6lYSsLSlxm0WkUKz21QAfPl8yWPx57PG4baK2TqIDRmzFIca4Kt4hkJVPI
Eeu/q7I5mpL4mm035ToXnQLeSJtk5wMsm1ZmtKNScxoEqHp38uhaGtbb9C2eXatvrbGxOOWF3Fh0
xxk46xUMBfJou5imlX51yN9yYWDf2jWhrt8oiliDoOJ2FMzrAvg4ZZw0H/oYgna4dEB4+T4kSk7j
aCORkdDW3wb7ZeM8/5m4D/2WD3c55aZZ+dqRQYGp30mWggp9eLqqO5JaeoJafgP4JPHlSYCRqZXR
h+x+QibXFE6EMOkXkOdSrQJCiR9rbOwu36ixdjqvRqy3OpIDd6hvqoH3ntyvKwJo23Bk2wkKm7ba
6OLOKEfF0eNsy5W23diMyrhUUZq+2kj7M13zzpFsI5K77/b07YKehcPnhvOLqbSzbuiWkinoc62E
XU8OzZ2wTS0b465eMnrU4vh0UAL8l/+E70PvPafMDzB4AawwMvVG8jKdwXGCB001DO8EmjldCahf
N6hIixU4169ecqxgiho/eoMTkH5kpcvHAV9zzWCrWCVlwlP7rjfuj1pT0WQcIDcaeM+N5sTLT4e9
jUTy9JozSedSYGh5hnNy597+3gOscnmN0i1g0gvvpcPZxu//Hbw0zPb7Cg13DLtk6bXRlab682sC
9jwWTlmKFW64chlU2urrEIt8TVi3f9ep7lZdVKHABnN7++2m0vjoWcJS4VmwA46nsEt+JHT71JHB
eHO8bycToAeWWx8o1HImqhuZfx7ehOvD7wmmXIrAlBb12nlDnPCxTyIoMDuzN8E5tHggywY9PkPz
zt6QshX1eHZvi646VsDEu/4G0OJZsxRM+BG9NsWnajyIvbGQTOrYstD8kSXsYYHo9noiagqjaPvP
CpI68LP4ckYXpUBbxXWyuPP25JDpjDs/m/4lWwTnX+SWcbqlc1q0vSBuqqoW6/QpYfZey8pzIq0b
hvZFuX38ICSLgxUe7vDazEaht8w6mFp7PEQIFXYwD8HvaDPJMNhZMEZf3lo6JYAKcqYYUGLGy683
r+LvoN0xYriKYBV0KAJxp/2OZ09Wt6VrOpFNCqmoOFY+smzD+UkVJ0/5hSQpWV8e6iADnvpckAto
etIvqynjRGE8Uqy+UIGTmO5BbK0MLW7arPcO5oMEg8E1Dm4pIz584CNRMb/XpvskUB1eIfuyofSk
HYyeHEqcxjRShglnzcaFze6XZJZARHvxetFp5uC+lE7pgiPoFi0DFkh8BqdUsT2gtRRXcDww3Xbs
jSDmd3jZuGLmxDmt3o7kyzQwMM21UBinGyy87mZv6wwfPst9nrxZ9WAxWMxOIrrgwW1CVnq8kZlh
P0KA0vsZiqOy/OKDc0H62efzev2w4dtWFXPQYAygh9u55gDCDjr+EStHHKS6Yz+xrrfOiVUQmrG1
ZnOZEJkOeNJaZE5JqC8Yeyk/dC8GdFbuQLyynQO6o5Gtx9ABmWYMT6hdpAv4xCjSSREdHvO72zIW
Oekp0tdDQ3naftQsHMTTEH09D7j0X0m14lIcxB+KxH2f8+Tg+7xA6wT1j94sDSUcCRJDZ6tkMfyY
q8THEwjHzOyJQZqg1jYLGsgf1+BWH6p2WF1N7wVWEi0ura+t3GCYMiv4VZ2RuUcvSP/626fExQ5I
bIPO2uH9szoWr9ySjfYpjxQX78HdYpKv9v4WRWtQ/jGiBOOCJHUkhT7OhgO+jVBMQpwg5iAfR4IN
SI22sWZZXadh3gu0dBkQblSaO5Vwn3KeniA+2Iijp39QIgvULRbGoRMaHZkpUrmCpJQItkODyiGN
U2sQlt0Nog7P3z3FPoanPBYFGHLxBvZQYKJn8lLO085P3Zb0eHo8XGuviB7RoO40H1SL4oX4fNcS
/KdEyZw7rqlfOl7xzbN7MLavYnyaOfLIq5ZgncfVu0Hfd9HolouVxoS6q79s4bcYkzt5ctruzfhs
ftlM26xh7YESx/4sDNQjAWqKE0ScZyUgzj99pV7iKE0aSx7gojRL9xoXwt57ycy5YAreM0KZgZ3e
JBeKT/OLTTJpN/DjyS7AIa/vP55LLxCJP8Sh6ChEXTBFjeW3iVnUfhyv98aZZlWJQTPosLJ3cPbN
F9GL4VFsJtEg+5DCLGW8QqOHXbXrlGBuJtujt48Ez9gdjV/N7PZ1SVE/8xHz3j/forQ+S6eZ6G8S
JEhG7ZnqZpfNg6S9i05NyZ5AVeeSg3FGTB1koQmS0PAKfCHjgD/c1asKjD5iWoZKmT4t+Rr1ZZYD
oQijt0fAgqXIxzxcbptT5iZMEzSOmAJYmTDKyTsakBFRbMHy19qhwLdZ5Lrgqpc9igXuiPFoghTD
2T+xGrhzAVtJk8K+AsoRrEOYclpOsevWte+iPwkr5SIHGwjXJdVd92v+9Azu6nIOD84GIDhgeP9W
mlwj1g0hnwj4oxJ9BC4RYjpJFwmUgyqNaV6vjS9pe0reT6Dipmecmb7mcnR67YWCAFsbOL000+cR
h4kdAtJF/YmTZgJaRmDXsGTIc5pyafy1DKMWthuTtWBas1tU7M0wg7ySIeqirRFNUMsomA2/YRzs
NC/zGq73gSlng6BH/fX8xwtc/+pLoy5+17SRpSpFfhDDZvNY92gtUaCP3/9HVjhKr1N/BzzkNjCK
kj98ZOB22IMkhMq2Fo/sWNVZAqNw9ysuw9yMTXcniSyIpBs1XYT9Oy1NSM2e1qIwir/LoF4GInPB
De+ZnEVpq5K506JgowJ/+0UDqSLOx1wPVZpI35t7N1yLcsHzSX+FdpdwgAT5UWkZ0SyBzp/6Hjmp
ZA7FRC5qv+ij/n0JEIWdp+aqX98tT47KMX8sWlRVhbJ2+3uqSFcbHcN88w2abRSfD8yVAN3Rl43M
OUoBSL8VwkJwONJYLKZTWLTbUyMttWd82KHrkuxKNw0Uorv0h8K8JgSgfw6xmfslqUdsnD9npFCk
Z0206TpatEb/dRgfH9JH9+g8Y11HqhCEvsYtQVqMAeK3GOQVWVvF8DMTAMjBxesy75cH1e+MskOS
1W8dhzbD43yuG/5W6qOeTiIKjUNTCPUSfpyZr3S5kbmUid+hhS+ZqQizZcz9mt4nANP65Wo+a8/Q
bnIDSqK7ucBFyM/M7vlN8oeZxkea1uYtkfVgEtdD6nxp2c9wMq+0vL6IJJRlb1AtE4ZXUVf6gbPJ
b30NpMR+5ib3zr9WTo8hn7LRxCqhyFeyVDVoabdpZptapSdPJfX7Wz+dIOH1puA5Z+1PBlD0FOV3
poHXOkp6Rmiv5/2xquf/MsGvrfwHUN2Va4mLG5wgwgGF2nfY/g3Kc/676m2eSBZA2BqGV6BAvI3s
trVN3VwWA/n6W2AsKXSfc4+hqPIPb+KSmrqFBXxg+UsUWaHvQLk555rC8Ys20AAuV0t6lkJeeYoM
mWO29BPlqZbyWLIk9XP67ywVygp3QPTZmXlrVrziBfDolelAmz7JWi/fMMyAVupRaICVaJsm4nCC
kVq4z93+oB7al9XU9K8iT0VarNbLROTx039GrZDoW33OBwr67vLF5JfGUoOnhzSa/UDc/giH0d9o
9wQqhddFYU4HFTgsGP6r8dCeIgDA9fwbCK0CEqLgX0PLvkl6Z2ca1SMItfUqczW8z6d9onOnH+VO
cBxBisNmdJgOdfwVaXpVyImwZxFGB+WJZ3q6W91oM4B1da79i57PFxMvLLrma4qUBtPjcl4duFdF
peCXMgjlzzIq3dggp+SbUHjwEsqp0oUssOX70LpYtnv2vR/hVef6h8GwYSXCu0ZE8pCoC9JT6NCf
LOhd32PoqlA/BO4t7tRxToIG//gYflfB6ukoa5ei5fLtIh3lFCAH4uu3IwOyD8ACcbzBpI1wJ/FK
ie5mPcpkuU+Ck7Eif1oJGwKMP3Mw5K92tDMedMAgvZabPmBV5viCO5wiTDHXBvdIe6RYzXa438Y0
xSoPVzzP50EXs9ocYKkFhLbsWYwWJ6TAzF9WlyGQ+N8aWf1mrvfl0M/qLFXDQ0wGblQW9XyUJZSw
cgasYEvlc+9N/FmOr6aM3xehKt5XESb6tMlVPyys7+sRShteX1g0lxheKkUAD8Sse2hExTWxqO2f
NhxjsNAdEzWPf/yzZNUKOgCOtbJx4ZGpl9u4rEM017s8hcC/gElkcmsfGaJ5XYyIzjArizNMmEVy
DkCBYRfAJmWyQ3KI0aAHUcShjq4+UKIMpw1OxOVpmOHoZxewdRdAPyrnQbBUEMyF6P1wOqWbSCnD
TWLQQ4AWWtkSPF0/OVdhr2/UVmCSwNFLXDM3cmAl5JJnpzPvwvMm9pxzroLkvkKyZqyKi0TjIRC5
DfeBSVLpo3xHJdxL4PmaqvvkU7gzpWBCV5OOjudWsyTC7mr9Yp7xlDPBVDBZN+jn8d55PgCa3+/m
mro4MZCWLFbTA88T5503z6sJ3SaYQHkPVDDY22t0oLt9pa28fZuPTB8qSiLurGAgOrBo19XraZxb
2u2/p5I3vOc5gFpK4SxmbuLWLP8AItoLd7liqOna04GMN8kWx6d/PJx0AoxFVkpuy3s2pKTSem0e
XYiLHSv5LiWNoHoAbxE5kgzZND7WC5jYRLLE4Xr1endACecH29xmaTmkbSERnNhAUgoCHU6Ukidu
lyvSIGrbnKzxSVrp89gpgi5kS2/cBvVa7dNgMBv0/ufbtpVDVAgG3SNlsNR/HN2+Lt2ybLlDwvGz
7msEAN48zdk6M6z3FKJAHWtZxkT+UrXludaaLS8UBg6gKK9/pxAHB4BXpkyhwaIak0Da0YJphuPV
Dor+Zogl6A8v0Wug70c4LQqbW+QT+P/VD5qWk4nWRsvpTdujNppNLz4VxM5G0fH2L7cPwhMuAGXZ
lrJKzSX+xsrv/oBhKyHc+VTMZ9+2qoAhco2p06Bb3tAr41/ZSH2xHqrvWCgR6qqfuBMNJGSwsxFl
CCZKI7WHveCJPIbPWOWGMVfND/UBN9Do6D5PuAN5wg9T4x5QZOQpm6BtlyHJSulqBMq0H527BQui
K4IAnxLL3C2XFU8Mseo/IW2itw9Y9tr7HmFRcoBxPm+blDBYK/OvwM9MXHGkSAiPF+TJsXtjI1E6
rKtTlzFiFaHm7RsK9XtmYjnCEbqi3Hvz90UtOCJnaSAlgu9avFQ+xGJSfVuq2LC6OHAXkdDn2DR2
lv+j5umct3vWJ1J6M+AoBrfuNzod6doUz4Zd5qLimgV76eQ4L+CIVzEg2s+Gx3Ctl9dMODS04HQ7
+u0MIVs/EGBLJPs9Sw/+7vWN0DJ0JXuxn5ac7yb1RxfZCbzYtt4pG6cGTIQHTGA1xjkzPxyqrTqr
V5pbZLNETrpBBgf+FkRCrAMh2aGVPhaTOw9rvMoJ4+z16qRI6DtlQVdLqp43zrt1excKDtAMG51r
hrFYSz3tp3PZvziEv0t5II44UYhph8R1SpDys5INTfz7vJZuOd+2hJYEGryKuRaKSY5pOmG154gc
frI50BdprkLoX8+HNbEie2L40058ttNivRsAa1eDkZEmMnUjIp9mlOKTR9dV+LxmaZrY8G8/3UCn
xvKWsjdVn+tRdpvnBnYLXbhytEBaHAb3tgPJbq1UVZy6D/vupXIwRomtgt95v10w19dJIBB4q83f
XFrB5AlqZj7CdmYm2S68uyMRzO8fHUrYeKNEFZwfj4kQ8v3d6HsKPIfpzXFuclg40BpN9NMLTGlo
e8jtOEPbapE0snB2IfEp4QZd0FxtQW4WXw/c2JYAoEYo8dd2IJNZdSeSAMktA8iLTdHaYck3zo5J
BQs622YaE0I+rAE+bzyXyzxBL/5L/PZAkMm1QdUX5uFt2/X5QSE0P34W+3qj8i1t+kPgtQE/AvRZ
K3exgp7XbnU8d41aFY3PWdODb8vXnRpCvg2yvGe9jWEEdRsglw0he5Gr6LRiyPaxML1LZ5Ws1nvG
0wu4ZAs/ADPRw7pTGjmXskTo+U26Ff0lAV73pqwPYEwWZRRDWVN9uu1cKSndOuzfqVi8zKiiYPuR
UrR7hpsGMl5pyDAUPi1iLuZVMdFkuZ78jpv9PgWVIkqxSFerqFWzC0Jgs4RaADAKiEzS50dW+JGz
tSxFak9c3GstFlivkRyRvvqY6Z10Hg8nHp6IqVy8QUXYqMJrby23X7Da0eptl9/u9f835lfIuz8y
Rwhp+5P8JSBDvOeKo1jvbE2SflnSipoJQWKvosM2FVH5PpRuaJkXmHUAlp3juzsXbD7S8Kwm8YZb
LFtWeFEwyRLh6siaBLMW3aNrowYpGduKV2eLHM6ogXp4OxVQOpaOr8FIcjc8fAI4N9MkUJpL3PED
vLiKZlOvgJnAD5GZanjqfV9/UwmbUxNBWuHNh/I3O4GTzeZsEfwjDy+l9fsMlIed6r3TR7WBBS1T
Bm+OzFArW57EHdBLSdhCkGDgRa373rTK7u1EYCl5F9ytbBhlRd2W9I1d1Rst5ZZ4LvF8FSCg3/1C
FQJ0EHtrL1QSQxIuKG1DRcslHURXlry+dbs6dEUvgdgMyMbfKhZrpwNS8ABKkAi20hf/YQZ6GUVv
tI3ym6T0OekRXkTa2c9BsLHKKsYgosPM6Fyjyl+Q11LLMx+bT8jLxmFxv7lD3z8zgYivjngKGGT7
UbV4KURZNZoOsd6MyijWHcrAQ4GjVKqqnUUD8xUTNSR2H7AY7x/VcAn1UG/uIu/idabkKygc49pm
+mxmpB99lsS/qqwNkh9llf1lV8FwqGfprciI3wWme5nPoe9qhU1GdcE06LU5D6azEW+p3deWfyty
T/U98MEDsOdTrcwDSVmK0Jo5KnTaiUTxnEcNxi1cxGUDCoHZSWeLgZa0KlhZ7/STRtaIPBkeo/sO
9YkO+epN4EFgOJ9uEAVGGI1INyGLyLzIC7LlUCkQJIpqbJuxBctmUJ+7TBtzjJr4aQ2z3ZSBLyoI
YMNR7uav2Bs0Sp8k/btT4bTOb7Nx+KxzKbcag7jD+UPnG1HAri74NoDvIrW29nvCkK0AOiP+pWbI
YA+fMRustrGdjBRbJo60OaWf5kGWBXEp2inyS4xjuylmm/q094AOCnJfCeea6uViajhrfuSLNYFd
TB/lz2fHvrk4fm7xSwV7ZHQskrKMKLB+bpfCp7AMAi/qcwV+akZADds4SYmHA5WROVzj75BdpwSO
szyoF6biQA4vRVlaIjFrykbo5XNLgrz9HJd/f/HejFtl+RoU/jvscj/3yE4wHJv7iylbjy7L/A8S
uWQyPVcsBs/o8CsQdp7NYIfAV7c1d/xNpU4y/TGds33mBFhICgPF8ga6ef/j2uKhHeoghoLB1RET
qWCuv+XHRj1zUBIIlrj4vHTWpMMgcOZ0OkvWbZJbu/4ByGDo5XbT31hYKV4C4NbEZz+3Av5YTFm8
QgYNrx7jWCdPAIaf1dDvBqAorDj1dFZqEsOmP3TJsj/HW7DSkkhdXGf/EnfhY7/nU2b2i8iK8fjk
g6Jsk22LglwuN2Jk7C0LnzDe14xWQEk42xWjwMq+bl26bOqN2KWdI0wn+9EeGPHOgH9Qb01Vk0Fq
uVJgzP+zGMXxmqa8TDlBNDhnOKRKaYiWPOG9EiLthJuMD/7SMNB47GecQAIM8O6WxI3Mujn9g2dJ
zzny/73V42VaCxVIUnjZJvlxEu83bYD8UmRUNHshtmE8gOsQU3rKn+d7nO3C1y0kZELGCrS+TOlI
0TAvv8ZLzuYza5he8xMAODdRuyFjM3bGk1X3znnAXDg/sKYgFBbuqwVc6aOLshBr6WldYfyxA4JI
d+2y0PN2qvcXyAe1beBxQy9qkncZ3zCA71nporXHR4uJYSXjIWQuURTgSJ1v0IfjYFoL8L1WKWPQ
Ar3r7wR+Fa7Gr1Z5iEYZXAIg/me2eg6LWgF6lKGy5UUUnP1mbXug6Zhjt7kabsnsaQcNnIzG4HxK
ICNeWY4+0CpLdhJkjO9JTMhyjl0zNoqIoKbZRoflHeVsH65WXNQuXXvkXcLIEPeSzTs3iceX32S2
tUt//8ATaG4N50P6dQxc0IPFCOFNBOhmS1NND16t5mo8COEN3/dbtavhT9dgA+17bWzpQtBHA1bj
OP45gikqionlQN5nkbp4m+F3/pUzLO3GHSP4Dro/FGcr3hyW5Hsr4OyZJXB/Of+wQ/zKotmIiTTS
ABE3qn976sic+znvfyiNaXjCnLXh2AYjRNqVNF+c/kTpJTVTbNYY/3zd7P3uTL+JPlOxq+ZiDsgi
PwiE1YCjlQf5HobeuYaTjZEYofwP1F3lz+2SZotoaJeMWE0ueVhHJvBQF31VTkjEpbFWrdusH+RF
dGeHq2sEzGrQ8VHWETHfVzeeu2JrmavtQ0rt7yUAQB5KL6RpTUaxgZowBe0tVmOsTPHm4FiLItV5
7FsXg+7Yyg9ErVFgR1LT9hZl7iF2IMQq9YW4GBhPoyZjNLVZx8m0wM6BsXxS6014X4oDFX7j5DEs
p/fB/kQ//h38qDaP2ikKh/E/DY5Ky17aLFRgr2jZYrwJb7w9oYtgDJ5oXLkJG20SW5s9p0eSObpk
faF1zlsg50akigZ5zC8bAkaeq/BzuqBn0wF7OmJjCzYaZT12pc+fcuChfaIt38VfGU9dEsuqiFdC
rurvfCcxfuVuQipQ/sI56TpE6V8v6+7eJcdU1OBIlL+EblLdpkIdMg1BsTz6v5Ykgm/XfocuSl88
nGzIZJUhjqIuUizhwKKU1fWeFC0boniTO1oikrnTDq+1DZkBpbCWGg1ksl6fzLjkdpOwYoJeHCCM
cT//ZRVjPNSu0lMQwY05RbGH7Kg1aYRE0m21t5cfv45PzRI6Yhb1HjrXd2nD1FqSvRYHFrnLjr+m
MuL5KxRhmIZMWgtWlGENgWvvYjfOREedWlhIpV4g11nflAXswZ6Tlo0GMR20gYXr48h23ZLLtOTp
26rdiqEZZ17mYBSVwzlnhwt/XMrU1PLlIrHJ5li2gkuTB8A0Qtt2mWzhTgcIxf6EgM0MKIkYIpv/
inH/9rADg2LdLKuHC/9aU/EsyzC7gHVPEEcV+oaErr3S+1SM8lKVanfcfl4wU4nT1ZrNqpehPJXT
Mpeb8QL+o/g07IOvqZAjw8mSBBZ6tRUp4iOCBNiC8tkiL0j10bnKxCDdIsyVvLmki07DCxotrhnR
/OPIfhCcN4wRIAG64Q2JtXKnY2nnaSVgGVoWIsemX+1vmPaR5lld7uIJXwPe5U/qAjrvp78aBM54
ifcflswTGirSfP5BiEMr0DGr7bcFulrFhTRBtEJa6PHqAwNbTOudxi7ugJV/0GtoYwIAEy8fg/tJ
KfSNPhIOpgaOBr3YyeAXGiLCq0NhS6vUqeE4+AxGkqI2swBZebnVK/K/Rppfn3hItA3l2xqP13Av
Wq47e0W2TfpZ6LYK3By19AgS0VnPqQpogRvljiAfVj7LwdOGY3zntXXPYFZeVq8vAONS2mIJ2K0V
tqLHn4fEa0Hxp55qv1+7d8aaKnzUuPenkU4fgL+O29IH8RKiIY4zWcJMkASDV60AJrCrNX6bcDrc
4WDLHH4yFpgHWKGJpj4s3TbihCl6mZC0vCIAKqWR5oYXgDrnSbard0hB2oAyE8afXGnMRBVA6WcM
/3sQfPcWhuw1kN0zW/E5HRCGScdr/4QYuT+/O1mYx9/nOlrOyEvqXHEhnn/v/InttEQ3TgEwo9yQ
zRqrl9G4xiZLlgD0W45A9RaMFRDHuPQhlyGRqwE06G4f2x45jBJQm0Xaxt4ZJXv2MSyihkiODf/A
Rx19oF3dJO566O1igIfJ/CSEkV4Ora/mlPbb3M5du3dNYwzcQ3MLi5jOv+/leZM3CnbeacVZkeoG
2MwBysj/8/dLsUBKhrDjquXzV1htVqnHPrEHV2raKLxpBhAAvtzM08nPfAvSHuiI8SD9WfNHkGwx
jlu9hPyAg1oWYPu3sgX0f0+MKQpY2VzmOdgAKFW+Y5ek4wZSK51NhzBmbHFxaP6iuhGc596g7nv5
qGf2wZjQj6xiyU5ciqyfWkvPlynUf+SUXDzz6z3TbNQropQC0LZj/9UdFesLzDbyeLH8MsF4GXnE
0pOSH4uSIoSTXd+h/ZJ56dZySw2gl5yfYG+EadFUObfQ8WSq6Ox0U9FALppBqR1c+HDrAcQBu91g
ihjdoM2uUX3rQruADc0HsR20ZWTDyGxM9zQVaLwh6GCsm0unFdChiOq0LtVyOWOQgSwXpqkfw1/H
dpcNCTCsM1lXDPt4dVboEm3XSpRTfemOF8G/w2feXNSGVV/82GskwWX5GBBeDmHyQlycsjrNwZ4A
FI8XMaspmW/Qp8M/lhMuCALJ4u633osgCMxbZLcbXv02PhVdkGBipjbT+ZArsnfBBwO1BedsnxMS
fhRtL+A7BKCM0wyO1EWBFHLaJA5qWzTqKf9DAF6TEMJXJQaV8qblgHDreXaeSW1GCnksg90ZAiLQ
az4wg4aKNVV2QyUhpGPVbnASUnw0Q8HsFgH+5LoN/FsogMV5/cLa5fl+RheYDC4gghmtuu+UZYqL
OQkOnH5t9HMUEsUu7Ue+V2MWyX5jp3zjL2YcwnYo7Wat0FdCkG0ZC5FJ+PCy6QNsY/SIfOWMFL2m
x29OVjeoreKHNt7zbY9CruILyykXew23Jaj/bdELg8EWyZ1PrEwaaJgYvwza5KJvxI8T/DsGdgth
PU3Kw9D42HnUVJHnloM2nzZnHqUxU7xL3tu3TYZ5kBTzn4J75tNTi7gbaHjocyWU4QAS2pZY4av8
LTIfxaw/lmVe8V98Sfnb55ziu4RlhB7IyWE/4Vk0iTIW/x0NrlBsojLYfyiD0IRDMVJzB1WrAS2q
Zg8expQzIDnkU1KwXRnPzD9ggmNxCMOmsV/iaGbYebDHpXI21+V37ZpyDoJFN1sLPWMV8ZtDAXqb
Ik3V4q7ori0q6ljHfAPQz0qIyA/P/mfDHZjUM2o4QJw6kEDmTMQkXbldNk47cntpYQhs6XSDAw1N
ilW4J79ofOlZ2vATLHaIQ5F8Ot4q5xcNJznhF3Xc14I8NSl0y2Yj4R0byRaioendruEARxEZHB0D
5Sy+SVHOcOI8M9hmyLX7aVLH/7mnNa22j8Qc0efWe5S+HeaguM7DI6+iELbOH+Rageg6uFuXNnSh
bPihEGh2+FjEhVaCt3wbtRnso8hgjwQzlI0cX5ofxGUVN3p9XZ+5uANG7FJC+aAeY23unxOxIUic
61y55lugwCkRG/DyU1I3TZg2LsZj0KGOzwThwnd36P+WTYJ5iT89XwfX9YwjZ7dboqTwL74uQAn7
BiHVKODFX3A8wXIKGTsdz3SlEhj4MZNYlyPVaJU+ybudjuetjrajIsmdKyxLSrmWvWRfLYZOfLqo
ntQoF8Cc4TMzzIfRrnI9kh7tNot5XmqDN0kUgKElDhN5vLhy6gAiHzcRylYAJMuyNGQjV0NT309b
1a91utugRQ0kTGWg9Eg2lpsUCUE+ybmDDandmzNqURTqKB7nFWCVbjItxhXLNKhdpXElBcQjWZGd
KdfDnQL9jlS9m8R14TnsCMXaVNLCId2rtVYYN3xj148PnqQsbsql0PLm59PWPUpOAumVSMEdR5d6
zvThc9IoMQXYPm60oxXRLp/n7p2YWrdmxKAwKDUQMo2gJWI+nbTjK7+Iyw3OW9snxij8GnpVtd3v
b4fUeyrpI+O9QKN+5tXK7Bns61ZrYzF6+5rzWJ8FsV6UeozOPt6uIeV2Kz6wYZa0CVBqSPwNF3/6
a6U9nrM4NoTJTw8jc77NJFHH0wgmhNgBCP1u73kX1V6eNSSAbzahx7jVx/9gK6vVMfapDDHXDQm9
J4JZ5iPWqDCLSF4bf8+j27F3LyXn3CcV8lCJ4HZY6ezgwexr57Rx7l+Pihbm6caU5dTYvb1teXA5
YrbXiULuZJ0j1iwfqyonVx9ssa61L7CZhiSmHcIx8A0eNqrc1K1MHancA0kP5rJU1fw6H890lBEe
gDVQA4JzKlMb8ZIXMoVwTOaL1V5Dr1CUcrNt1IOlu/uLX7oLVVJB3CtshBlbV5bO4hOBntHtZiq/
aZdp7vQ5QJJSmnGLIj9IWW8j7U9crceySHS0dbUFW4aQvBOEFmMA8idzSojZaEilD2EaLdNIHe5Z
hBuXEmuiwucSkSMCBMIAsuG15rnPccxIwtlLc0VKYug3wEBLCkH1yAUVfJeVZyfEW7nXtesvcifz
cr06WKX1EB/CpMHlExZ5NiwDn2pLeiToVN48nmJu9JdNdQ7bxPhF9KKsKtH2e12KCQRPxkXuGzJ9
4C+MxP+IIm5HuBt+2TLWTdBfdLDAVcO7XNhATPSMlwZJvNA8T4nSzrPxwrXals7C1JtZtKBW2dUB
VRgN+we+MwMIHCRC+/xAv1zQKgVjwbMDTtyoLR4vugZFcAbfm86mHZ/87QAenMGRlOHQhKMn89e9
w00Jo6ylVTCERC39d7eKHvsqEqifVaEzZC4VwiusEfAUtb3TpL35mp7RVTC16Z62TVAvmqmPunCi
nNAwCq2GZTd1RASCUrwKBd8gwmZFSvhFUIRMnfzA5pvII627QA0TNzbU3eeM77T9EYp0VYblfFK9
Yv81Ou2Q2AGgC5uGIK31aAWkifp4tClxdyCOdtngf+zjth09Lzg1IXHXuP4DJtMFgfnjSdpKnrYZ
rcyvzWR29bt4TSU8DqS0zBwW0N7jKDoQhG18NcdzONyeq21xLOagO7FuvSZNGCyviSOpqirUhlx7
YbCpoSfTd2cXP+XMseH5JVB7CWcHEgOao8okhrHcwTnhe9sw5OECerVqDoo0ICA9Hwef/XxTj7IN
JGBiFJNCiMHT72gdVIMpdGtFVfAqZoZAhefTucVB3UZ6/1DHQQuv+nlregSOEqw9K0lExdu5hlJs
UnT8XfnAVZjOhUfkvLu8YMQMKq+zBCXN5cCnw11ei1qUhyo/Z2r/zYZ8VCeU4yEsu0zKUC8FptZh
+RT1+KxgOBNKFrCaTLXlaymvy16ypuZSkwxCwcg8z/U2BHR6vT3IjOGqeW4Iwx3JHx3XmJHd8uL2
pxiXEE9EsaYvceYSDdE5UNySp2sFEzjZxNq9dc3QDxp31t4EHAYztc1fyaSesWVf6kdw9GPoUTI0
Hy2CxlZaq3iF6qpGqM7wr3Ly8xfEMtBtEK+F0ghZ1sB22VjTWingnhwYhpmLbRNXRdsZabnNc93s
wZXvev3O/PqIqOYoHXDav4A0mgZ8yEGCI9STxktbK5/JfMaSk9ku2s0e3CamGNn80qdWshoCjAhs
qEf7r4XJ0Ma7+3FFkrGXaZdSYF6Q2SWZyL60BF1utV1/gKsFy0I7ckIE8267ULq59v34dwnJiR/v
8gp0GOZ5fXwhbYlckzXtAUC1AzIKN9H8UKCU5bUGPMuMVR8u0cm3yP8BDcMYHUzTI9MiLTL+xa3G
nSK1R5ayGkLwD1e55/S0bEr+bL8MmuItSH8PAOztcLJ/iBsREdSDhMGE5IINTff2Ddg3FjevfXJq
+TElKokkOoXr23+fKd+Xv7Pe1lUeYYZ/zo4pl67JzL0Jtxr2eillTlh/vmpSuyOqqihYKtOpNiNm
Yk1ki5m5lxidtKpWVW305e7sYuRREtIyIxqqqTfvhZ5+sxCbpq1y2u84lUFjYY0oDNYTj9quESkx
yCBXpqg9xAVMkCEdms/XUyLY4d1J+B7T85O+dF02WwAfCYz55XiVL2MjeNmZj8kDUX8dXAr+fCot
60PE9UoPonvTEWDKcjHihkB54vExuH3kCYFC7xXz6xHelvljfrJ5AipYhl4OErWDtRhz9Rjm0OHs
6vpvXaaRk7aIXsXNgODq5cFrSekUQhwyE6g9pWSBDZgzfDtpWpvIyn25DEuadvMQ/FWnJJ+AOVl+
KAE3pCkfqWCScb5+fxL9vYtQ+CTv0N3cCdUPyN+ILyxZ/56mkVaUtwjWVo6s/AkxkM7lOiDzzvqQ
Y5X5UlvK+y13Xc1Tr0CSmDtPUUUoYWcW/gNYNhbathXiVg3tlrmxoFOaRwUVVr0rgZ0BGjQdokl0
ND9bBmzy1dvi0jT+zfwG9CsQ7TW16MyGtMaDFi6QngrPGv1cj8TzzdcVGLlAK9GYCsDfcTiTS4XJ
9FjxkrqwLLouWlEUp1HvhlkBXwCXMcwOVVy760qM/ZjogxLHDHQZa4GyLM7FoUNK9yPIbbFAPNN0
aqoocgXYx4QAZUnxUpeI2jlKC5RTin8vPPKBvdFprEdn+O51MrtRNOm1NY7aBTAbBYbx7cMnUV5z
EXYXZItH5lIAZdsH/GcUCkQAhriPSJrwPHPOkTIsjE6i2u7TOJLYFzlWuhyyOIYOgOM0PD0QrHQ6
IL5EJA3MDnIqv3xJAXOcTv8k8Ek0MNPaxqa/+HfCwzzIvOPay75jSUT/+i8J9Axyvp0jj/dKpnHa
PyUUS+GFNQVtI5EhNL+PVC1gqyhB6aG540YVcyYhqecg9B1MNmYgzg6z9pZOE4KLSsKLJvMJo0Vh
zGssYALeKmLySu6FKbQEXe9KCfmrt5vJSqitY2mkBdmwCEm8Z0v6aCcBvTK2XM8K0d3kIlPGtzWe
djr5VdlO2CpcuaqMS6eOQhM/d3Nwzn2IcKuEJTYGuOskL4pBl7lnbHCWDakbdvcvr7ykfiin+VHz
Wc+cnbYrci0H/KTKKR9PTHkoCiU1oE2Bj0hZFUFGHhUcgfMoccWBmAYAAogSOd4y7byU6Q/Nbc2B
CYL5nRw/2Ityz263QMpxVjl6IzdRUxrDhJIjPlG9eDEfEDn0AJ4xXq0lkLOIoxDrDmKCOCvYbYbG
Ht5/+RAEzTnMA4bBdnVEw05fIXa+9yK5QZLvJXrH7/nxuQA3cG4HIkAZ5/+T3AQ/ZOGgHLZv76c5
6IZ0gKWInLG7or6v/aWyuXkxu9oHrtqgPTD6wDd/8JHS9DeGLieOv9wTbft4CX4DGffdKwUse3Tu
Z/DCkTdEhEuPPSS9CIZT/T8qdw0dg3uN5FHdZWExvahB1KiX4aXs8gYk0HYYpzs9HJHlQBbfHUbf
Im1saUuj/pRE5CMoJqbEVKf/vEUucojJ0zvJPGzhJpyTpxayjiMrLcSxKm8I7t4Gh46BN/vX1Fe+
7ik4RDHsjEcculNA5W4EfTgUlKiWhykNwRy6mvwwZoIHTbbeTeeIMA8N3SxK/asheQdN2XrwskU8
FpupA05QuasnjAs6K6wiEo+AiBe/EKH36o7eQtF9HAoLjXuMpH7l9HKxbNUgfdLeZoy5TlZ9NfME
apTZ28HVGjZ7CfrsrXMNmfMieGZmyvUtvV4U9P40cH7buYSeq9ZpOuPumqxnQR4LRIz4UZDBdccW
P2vmw9B5aRL+aO9RWe6xIYaZ22d0mQ4qimvxuWlrUaeUKOXYavvDXQkqi/OCCLNtrK/r0meMS5N9
VcQHD2ziZrNO9KOrW7xJWaIBWOwwF2lsZD7DZdaya4F75SDGtwRTI3h+UDP6jGZAeLQQxIer2ddu
U9WmFNErFPJbUDmigpk3CiMX5cc+2K/oHzVasy6Qmjfqn7RVNaH76DWphOxOYpmYw1785j9RLEKf
2VcnUAouEgkwREKL1Yii722EYYSpvO/HIjcGWRPdrE+bY8lDhcG+AzD1IJX+VuPqYNYhw+8KZyx3
djfqYWVdUWIxFKNSel0iHFWIB88AL6YSwQEvAIfPfobU7UCXDEUvKusR5Os8Y06qWaM91IEMohdU
/tSYpjykR5frN+KQfnKhe8UfnBLlLikunnk2wgHt9OcDN98f56twz66iJEH8zVYoCyBHfwxdfpjo
Kmh+ONIw5TA3atD6YjlV5UHekedwwuDdMAu9guz+/bTed0C7L1LRKknTe+HcuX+KYwE9/l2zDzvB
3+Gaq4JTTASbTqXvlH/ut0df+EN9wY++GKESSyCWkGyHmYrIhsY/+wCJh57PlUIpy0gQKgheTEke
4tccwn1wGG+oSybBZpoTa4afRkaLXDh8I700gFT7YCd6Ljpb7MAf+RmaeJ4VTPJmhGjtLnYQYDcI
3p3FlcIceacIxLPmwTrOItHctnxaKXnlqVHt9bfi4xll41f0q0pd5hGUA4m77QFimQctQWU+d+Zb
dYbgMC8Q8yvm8Mo2SLQC6II8//PBty9gsF3jD2aE01e+Fu0EZS4menhLYb9+PQm6YGOyzyJpZCTe
N0JWbAOYivZxyZ+aiMVE1EiYz1apcsaGIw/DuCppQeUcrI7nktPgBaFYTGWknXDvW0IxdWLfa/rv
z+/n+8S9WM2hcDil0glY9dYSNwlM0kHBItZwEXFpS0moywrqaNuBgIKO/qPVWewl/iJQ1605FuMC
v/+YXHFQ03gKXZpIWHrhq9ntcI7VvddItsnlgtM9VlsZkq7TF+lv0zGyJ7WbvUnP5hcR3Pdi7+ma
ebbvq272Snz13ap1GOmsOF69BNpWq9YuFuJgdpph9jgUNl43kmwm2T+Y+8O7nr3k6cUjjWgG4+G+
OI9pzuqhbSsfzxwB/q+VLjwYBOZbP1YqtiHi2zfDeDZX3tAxtGj8nmxXpxnslR0tEvLhFpyxIayk
qmrmY3MBaNyMxPE0ICG+oTqBWgulSdU7GhYWFQ10uXCtJLu6sUI63zxsdCXv8Xqya4/BXhljFniw
/kNSBlmgF7HPyWoGPRlClKc+pnuazvGZlA4+dh5McX9rVqXnk+dr30WX3JCaiezSOKaiBwMZlS+R
eyykwCDE3FQLbw/T6A2/Zmr8ROHeH9zzTv1rd4R+7+VvQb7BhEZ6JEC5u/1urepkW1qNyaa6/Ho/
n7Etzbd91UQ8NShdS+M6+NFTnyOyRg4boxithNZcD/ZfM86VUVeqGwvBd9GaG+bWtoh7SMzkMS2O
tPusWEZMcYNYVwAyEETa11ohU85dVSU8JiBm7aPSFtCZiNE+NcyISuODWNWuUJxyswr7OoZu23Uc
3QawS6bsaPo1XmwoRVzGnzBMSLdz7mB1gFOfIsvjDnkFE3cIFbaYA0lQPDARLUH6XEdiksAnXZFy
2ODuUO2LPKONyvzb37TlekTjkpwwmlP48aJb1zmgRv/ph0tfU8d4PggEFjI9pRkw95AFupP5woD3
awYSlZSjztGoDuyAg+Giy1RuUuyTJz8Zg7+Kgv9vVOrK87Cz83FhXTNIPVHmD5PIF9KwQkYMQRB1
4WVHSUGVheQORXBzZndKeSZqDMaOQZUL2HlsvzXOBcuBPolUcsb0bEdQhgRJ7p1amGrrVINKTp9T
eiwaP+Szmy8O5uX4GPhACqwiC+OJL0qLmgnwhJDtGNCqcBv3/uWdhy7KiEeqZGSBwSzPyP7Q1aG5
snhQyp+087H0qHzrWpKDm6KO1g4+stx7uAZ4MoAS2eB3zSMbC1cm0BGUwEe0WHnkVc6PzBVWMJzd
RJ9g120yEsjZ2Bsd2Ks9V+IAUzAyQL8C61FyPYvq1+ZYLpo/CbIYQgdMKzYqLSP8adavTUBWn709
eVaLSOY8pNOkQbCuwRIq4Rnr/HYXbdOGYARCPhHZB49obIbshaVi0vsS1qQCfouVA1HKw5Vzng1D
oe+mxcpruiA9fetpVBXuLQTnnL6vpJMR72IlY1P34Y4Jtb12lttstoSDP32NC/WVoDnY7gYWyj90
iiERkea7rufXosWS7kPjasvO9areFPfoM+gVP2Qj2eQ7JXy3yQWjzxLpvn/EddWPNvT3awvTqVJc
nCs4Gmj1jVRl1AnA/M6dj6RHakoEEG3ypcYoHW9YtRWTPE10wgqi7cysijfmKlKUsZ6csfQQYzDj
JgPsfH4x1EOFuEwY7bSEqSwdD5McQ3OqzJc33zPs/H9IbIHVZKz9dtYlinvZjNxwSoul6J5mQpox
ZwW+ppknuMZMSZbNlct2D/FXg2X7kKyqDKuR07R54YnxhyMFanAscWmxymKgPwHDZv3De1GtnGgi
0Uhspji0is8B3Fat4ONVxM/3bqjjb71NeWySAKlPkTliK6YABX7dC52PRcD5m0MLZRRpopXpIkYD
YTSL40bVDGqBbWGv7bu9ATaJoxw1gDGRXpJa5QcGqrnHMKVvNrVajZmOT/PSFfcjHody8LQS0UkT
rnc6gF4Uz2uOdqYd5cfABY9NWz+0t3dfxQdVLJ+vf2k1SknS6I7LOTHxXfC0lePTwtbvj6eRiAvl
mttZs0qGifO8faDWnwQrwFW7AXBjllz+Yia7re320Vy1Kb6umBSfIoGAjUZcIyFeYgXSHZN8/wal
CeKqrr/phpWNaQFX2Wh2Zk29WlP92HuRZIHib5u+KJv5zS3RBV6ojZythO+sBms3R5vTFWgdiZIO
/Y9FDla/Toc+ZRh0Otv34POcdvThBTJCwOd++jejc2eODiZeUJlWLDjcxv+wgCYucqKqWeZqLq6w
fELtODAcoZDoZEyJewAMxn+SzmYLZRgyY/0uU2aXNPvLezcZyTmI8llqRRTHiIPyucPRHtyEv88U
yAsSArPxbX3TmoXJV7PoUVspVKL/JcRYbcEJitoM5hjhwbf7QGczf9EL6j5TtzKaUurCWi/RXgSF
SO7snrtRKOyljhiZNFpx47YEEKPyOfWY9Q+oFEisjhtLq93tjhxKiSAZsxmvUCLIL7PTazey0+Qe
YlyKsI6n9NO34Jovt+XkDM4Mv1xI8z8h6V1eWnGUZ3uWxNB5QEPfw8ZL2QKD85lKmFV7CWB/rvGi
D4KdsW06aJILB710fcYHtU5+ERharDWDl3k8tsjKuOWfIYRDBf/qF2YgysBwAcKsCipCHRpdb50E
sMcBvfaEPtYHm9N1m5UcOP69TvUVqn44VaOqPmsmevjZqsgVXdIrAl3+PIhl7Mumu31njGe/6BBv
2CCGALYBowDbC0o2KA8shtluJWlDtuRMh1AieSm0mj2G3/vMLjsH2gxcVTuaeeshvsYalofviEex
3jOFBhOzLOuG2FLm+R/YyvmMq4IUjS14fwyywJ/h45PijPhZnU+ngrsJoR6b+mAAmdMTvo8VkpIz
9Sqj0BjrRCoBJZMBCgOtt+qKbwn+99BoDQudJsLLHeP1DFllzvjspDdRC5kgWJwhbb3CMOYeef6c
rT9Z6UHGx1vgyVbmtCEdQlZ11jhD9mU48PF7+Ny7qsJdFGiNfUCZtLGZgKmeKTvdPadqwbs6qS0T
31OF6sn+dFwJTogI3A1cKN9gxiT9nEh5wwlOckRzzJUBM6Hjau5CRcFeQ6lzDsPFOgvYsNVW49eb
u2S4LYj5WJniocsnVTFPaKHbMRckD7nzKV7uO4iIB/jpfVx/Q0cMPNrKu5z8CzoHSOd7G0LtOFiV
dTSOUfcS9e//OAnyFRYrtzG9NY8QwN83VfwI70pl63iC7F4GS/mRqcWokEmZvaidsV+flZlgD1lr
7zRoMp4+jOvjkoWoh5Xhr3Fh0am4/V5pqsf464cHgN020Ku2WRmQdOVExyrNHKJH+P8V6dh82grX
pDyIkSpY0MgHOzLfFwW8AumRGWTgNSIYwLN6OvPiMpBYESRDC2rMsTFPuwQxKFlNDl4kpLk1kHBv
WqduCOJpgsCqomkwhEovumzLexCmPfa0opgrHOkKYoVCnQqXb2nA+SSIzEnvi3tptDqI4ZRMyzYE
ZeA/NJmO+B/0Wc8rDSFBITOQQDDkgr2hgWRDBj0MwLYP2OEv4VSgbQOsnbx/e+ZylxWC2JD3y0Ks
JY0OHuLS8BNHYjwQw8wNAQoxeblz77yzHUfJpzaPeWSFVHwM2mEASGTLuY2ECfRkV4sj7svviANq
70FxDxKRj4Bx+Fccvkm7QTCnYFpwu3WisqM0hBqIoutCEDigyA7oYuYnic+S9sGjJzxWedWyPOZr
I8OOJ0iLWJ8+ZXPm4w10MhDVTp4BPuBvB6x1CmsZ84hheXWfVbLbDjO8jtGb42Ly0XHRx6svN71P
0Zv91gS5NHkazkTppIY9omgNUktGto1EXV+pGdzcjneKKSnrnOO3qrckJbdtkb/pDOWpA2kJU3xN
8WkeheLeKOe+jSNzI078pXHemA53rseAIYXPRRDb/9Wl0hyHhyMBCp1MT3GRyoHzGunP2y9pAp61
CVCblvJbOPHExhlX+6edfX1FpxcDkU7SLovngQ0ysjjt0sylha/tGlhlUwOrcjdT6xUhjK5P4hk1
THqhEfppc9pK7uNu213IggTNw6Y5e8Ip7gV66ykhWpeR0KXYrOioNf5Eq0amXlCNSPUAlBIeKukY
QOfi9357ghMlRgPDnYoXxQnwad1f/16s4RkYDxlMwkhVIiEUlN/MESZsrhkjFl8sfTwZvlofEeUY
XUcXtzelUsfxXWQI215glUozeg+o7P/KFn2M2gbfxsL/73nnMDQdVZjme/0J5xbTPMuw4Y0uzaqS
NfzNgU8tbdfIy7sYC1m7os0TFOeXvWBSrX+YRn9kixkeRHpIU8LKmeixUD8vxpGo9Dmmpm6fd/Yh
kGNvXz3olQqxEhdLaxY99cXDJzAJumpQL+XEJAYu4Yf8r22pxM5rX8w6qH+RncnPoRU12ODGAf9S
+lO30FgM48azfznh/gQUldc/8V7yJ/+Y31YPr+whN4/tYVdVTHe20G86oE8q4SrMPUAQXe7RE6Jf
MGAByIsqL689f4XACVCTTtovw5uzzRETti2oQUy1tO6mWABzlqnPAPt6PIlx3d/5WMcI2DGfwwSb
rCsrCdnqlB/8jGRMZQYxwSsQgBbSU+TWOmdZ1Wdg5QAtKL+7Uc3hGqpVSwwBWdly5fIzoC1BJazv
pAdcaOkiGUzgW/bRiY7CtTqkqhjwv+W2MjjHyy/yKJxxyCo3lsc2Wh9H6yoTVKnA+vRNdBfxmjmY
D+Ynx/sfwoBfDw0bBBRRp8ixRLlIUU0Cd1chm/g2tkft5qNt7SsBzfnIur5nchEF7GFSIJHJRWAv
ifjEiEWtKys6E8bjmM/8+thx2QsUrdJfa5FhpvY/CtPC4xyx0/27pXEqt9wLAiWkYlQ52a54MnWX
gbj08NDBikSfck85Ai6oN8egnioxjS7OStwKpBt+O6WiUOej2GRdE+NaKGt6MHq9pj9xBM1+8P4A
PLExKkAIJIr/hS06cQTLtZ6BM2h+g34r+NZHaP4Lq9dOmtr1Z+3XsKKFLKGR8GOujkV54aRI58ky
sSIptaBdozTXWvPeX0+vkkLCt3UCySGt3TGWzrof7G/q4ncP7hNVBI/j68FZYn2QMDPfjIXu8K2C
te3sdIgO5tJzgKvv5WhCXeXB8j2bjukCgNDehoxIrdFv1S/MtEKCMynHBrODP5+r6Fr1VtRf702K
QgOS53ec5xbECmExOiqOZOwQhDgJn2OQCXA3kLzLFCmCG6TOpoaOTWsWHwYhK5q7qVDS4J9Mc/53
oEzkPZKYQQO0m1/Zjd7CHQqjpaUrfGLSuT+AhnnWsepvRV2LBMUchCJd0DuWxTZBl00c7CXg2HGn
RzaXJoaml0PynqDd61Z1orlB8gW1SI9F6dkqhRBjjFZOKP3QApErXQ68rZyRUYWpyYrjO4Hx9dSe
VxMCRDlMZEsvpwZvR/BhE+6Ve44LHUOdiYly2mIO9fR8/Ahc4vl0SICwZeffJpHUNZkbtIqV2kwB
oEEy9AFb3wephZxSKY38heB1AtNu1XXnM9nDKK1fNFgN3gbTUtenFGmrDDRsTaztel29dvyBzNnu
RJxmFHqRTgItskPC4xosfS28nTR0NYK5yEpRoxGRrmI+Xl8b7K0yQEs3THs64tJeDA4BBwcHIeIs
hZPhPqFMVLOa6MBmBUOPbCzn69PSmc7FjG7Q79XyBzKJl+0FfsWZ1tb7gtvw7JQlmmxq0f/u0Bya
37i4GKFLRzkbAdFKSicGtnEWJEyPnL9c7DlN2RzmNwCmwkjDqI3niffz1Iwl58+mcStXjJmbaUIq
CtpnF4J7BAAQABGi4EfWBURPvNHbF3I0zSsn66rcNAh5JOEwutVLO5jxcCVurBqQ/DuFpwa6Fd5U
9AwpWftlUvWU/JHfsjREKiWobsnL3SbWEn7uhO3Qlrlv0ORm8gNlRIdf7O/iU52ie7q6M9G+7+FT
5myVnRrAq5jpPcoH7CsGBJWrGnmBoZ0ucKVdNQq7dJOfcpS5MAO+s3ckC3edQc6GsY9eWhfaYYZZ
/VRGUXu70vasG9mUzq3NQgKZovWYFmL81DD1qXLaKyMHFNun7nIGKxVvLIREYV3xZgXAW7xoUk0t
zBuIijUCFwQeIw8ZD3PZET4/YfkvKEmLn9rPPhov6D0PWTxHzel3EikBCIiknmqCumqpVsNBg8Y/
ZRruDdt7E8A/EXlaBcUON68pCsd3/TarLfox/CfjVSQrne7RtlX0oCX2branQEln7FXLqmVm418K
53I3L6HSlJU6+H/pdz3otrOIRi1xoMusUELbJYeW6GkKBydfHP1FH2C3QcOjo8Jc2Z6tYsZxKav5
Xyo+XHFlvR5MCirIfFrakotanf0nFvWO42T10pGcc7BIoPodU303kskfmM0X1RhiwQ8rzNVbqo57
etWVYVWd20iH1yI0bWW6X4e0QMI+eFCwMzYTInhj/2sKxdrrJk8JhaJ2vrBrDlsl7O1e4E5glRFh
RWXvjzNcfwNPhiEnZSghMAavh+tE0sOaksS3LtA6ho/DuT+hbFUjQpmre6AjHNo/WdERjbQIij5r
NQd5mGHBEvJ8233yqVgUBXTlJw5wL4aQd1gtGcfWQKjHr7Fom5d8Hl8O9DVHsV3WGBGoIeFDgK1p
OiGYY6f4/qZdQsCpgUPCauZ/3lt/OojVn8luWSfFFgZk7cCxvh38JTKoD0gtOZxqaot4eTsZTZE3
TAp8JyhWdRhlhSpuVBs42loRYaqj6p/ewk2WWv6ORcAa2TKHDEElV28Ybp2w5jF7six4Espg422F
CwBcmRdDr25zTAv34mMA2HezBF9Zckem0GVh/fZ6LOQ7POkukZ/TvARo2JWTyXU4xlL8WRGJ8CVw
9wh4MoHgkHnwHjK3BaHftD53WWdrrbP5vZe1A4ZFIT5SRpwoWARXeZ6pNGFXWQqI9IIrnXcNx97H
ymGA2Fp1sn1xln9ZBgINc2PWpfd3tD64t1MCX0ZxwJ+BrADUE2EEIurwrOh2KeR/VX8VaEXe3ZBP
Ii+uLvVXbbphi9TJOr7p0nQpBl4etNX6sErxdz271FlsYqPJGJJOOYEMhLXXnVJWCKhuUKMWLrRx
YlfeScznOX6u4qowZRGDMbM+HTM2znYoJvkA3FMVFC1vEi3HEElAEBGCZ/KJi3hc+NQxjrty/TQK
3cFe/DzoFPhVVGUJpvexP/O26n8MXJeI0p90XSOP7R2x87a2VHhHjyNKCSWNNJazywNoM52VXJt2
mDyIhcAr2roYGYQlZRZHmDeFO2SRsIUR5CcbZKhG4rAeb6OeIYWqTpfzEnO6rkhIomf/GTMUP5v6
NrlD7XoiuCulFEDf7WcOf0ScYgPIdASjKpmy+MiMBf7ZSybUuILB9QdDwu609VafPgxi+q7nMqRX
REF2T0098HiAkbKq+yEst1NVTK9U/8h8IpQWuzlZl5kIe9rBL79VpFl0OZr8rT9XfBpwcVFgPHIW
+NpjgKpKbjg9E6CKytRYP+lFKqq0mUTX6PjpKWEEt9NFqcLCThoHBAQDiCwVJWnvHVmECKI5W2u7
vHbr9ROhG/CF0fCN7VYr4Wi245eqxPNMctr/PwZMZtFSmWFlaSpCpkcQnc5HxJnjjo8QTeDfr9Pz
JdUTBZC6SQN6eTufn9mmvhHbanpRugEJZCV1SmZSUeK/FUPFd/ZWqChUKbIqWYqlLNtiwHNVfN1y
TR09An8rfeIqv+I1husiPnzeoUvIzKoJdJHlS7NpxtsMPcPSnAej3hFX65ASKBH8OpeEVGOpMJd8
e6XYnsoUjky4Jb2qh0eC6hvZbF1QwMXojT5GrAn0v6M5j5VgBG8TahYf9Dp9KToWxrge9RGODAZf
msfSfzszb9tDDJSrYCBuPz8o0XJ3n/l+B7BZM5fZ/4p6xgTxYCQEOjsoiGE6KaOanC33vUfVlDAU
hBAs/cTi+FXuFnBDeY/EZbtWERdjEkKWqZP6CvEcYrbBMa4bSjk8u1Px49DpNT5o+359cOJO3Zuh
BEkeBizD2x0BG7eLVR7CYlRXsAFZkntaHuFiTUWv9asdRBVtjRtSiwdhOsXKM3/7pF3PwXcZNhZS
keYvQf2trMtO9qaPsGT4ar/WYZmT703bkLKyiBTo2b+DEvgqCGK6Pjg3V9dpsJqf67oD0itzwAew
a6uCUJvpH7JaX7ZGsZTBr9jvvkDU0EhhCsS1qu/IWnPVMHIdXpfCVaIl3p0Djsfi/Jo6o40f2iBr
SYxPj3kdPwlS9gq+o014UwIbVNSieL61vgH2k/V0dNZtNRbB/gsyRUU4/Ck0OFjp1Tg8FpGKjlBo
Q1ViKMgLj8qbs8eywMp8kzye1iAX3Si4Br5OdCEhQ2SCPxSB1YnNzfGbWIKXw9v1XnX9PLmU5TUS
sZ2LL50EqombBPfcuzyA5pLeZaj1jZJsfhRZwM8z7RwJcyOw2d5gEgEyuUvJjv0xeXYpRiTGU7ex
pQYtI7ytZmpPXwZyxSn5Mffa1oemkR1eNyVqEO3DWUu1KP6WhmefEpHZxf1LROZvtl2LgqZrBMiM
mgpT7BI1HU5gB8rwHyt7C+jmCre4GYBoX+uQFk8IlLGo+YgBJbjzcy+1zzOzIPp9Y7DRBN4HuofM
wapkB39KjwPWoWgCwh7AbQzYK7Ioz0O/v1sOnh80UtndmRhISROuJjTT5tI9xrufvcS2HDSjOK/I
1ZZefU47/uyLD2vZmffdNdPfRVTsHG+0SgUOjhDqoT9zmuE6POn9DDHgP9TmdDFagzek8gNWUSo0
dZQIav7GLr92Ok74OfcXcs1w3WFxnIJIS9/w+dkqhlaZrIWZ2l8aPfxDREaDwAeOx6mKokyZK5dA
yHlfrVzS/gQraimXu+aZ728lR4aCTZlVUyNcZE+VhtvmLQSBhBIAbBNB435S+abpV2WLgEZ1tS7F
CI8mUqQ1D+lBUYpLG1rAl+HeFp+znCztl66MJtj0YAugqrJ7htRM6+egmwVyALLdkHkyQugXegCi
bkabGH0bF05Lx/fg2gx6VMSFXENnRiSdmEKGvYt5RqD/Cs883h7dCNrp6wyaRamqkzh+dIJQQPNo
Wao3vlsk9zOOCLFmgILZgJyBHXGO/zNdU7ncufwZoAgWI2ae5B0ff6QbIzgERTEuFcsUc4fldl1c
HF1kL9zziaTAG/A2l6l8btMX0J6zIfwICusoHMc/W8NvQCr3U0CKiqnK10A5nlIdWik7ZXLeH+Ir
uPYm8u18QFtBxzf0QtcQtHzn/9RZ6TW5oce5JbDxjvkTDExTuJmUVn0IA2h/nrAe5lUPLVvkmFof
MjzhDRTEZEF7J3Q5MYXHqAfJURtyVsGFB6SMQeh1LJa4/lV3y5EAcXi7pEzVebSXZ9AGNG88MPmv
Qe5tLzCWzt9WBuMwSoKBet5+z3j4Xid/fSSbN5u1n5HXGJ6WH6zWnO7IAs+W6Ti5lGbm1vIMswk0
M90HRCEMGodsfwLQYlxaQijMYxJNob6rcFjOzLGaL6yFZzCIh/odenoAgE6xvvQByR4wr5pHH7WM
XSivguIVfu0vSQZ+9alVed4AxxfKs6vBKVbKXqV9sx6xJKK0vHy7RYTMQGUdbDm+UaGt1v+rPnVt
oO/vO51XnX8y9n83fhqcJidSjoQMmlD2Qj8mqsReQEPaDUYLjISH2QchkN6WliXF6RAxQ8pTVPMq
IWb5fhQmY6398Y7XNsWqN5gMzxCGeQAbIfBbY8Q0OrKlQsWu7A8PNa7g03uf9XznXir8UHqhWMPv
7Os81q3twE4Do/vZAJZEQTK1LQTvdYPKUTlhl3I0r7I3GcVYt3SvaEqqkMZFSGu1TRUJGi7u8rmC
EnZsbfi4LmGuLsNlHnKM61F5JJiHmyAZQfE3U0l2zUPhjEkkEw7PncE6xHRGDgapXqbx5Gf3f3iK
1zXzX0pngoKVzZQgHiwKZSlfkkRz7V+japWR4k02BP/G5AMWViN/7hPpupqfXKa8AMtf8I4kGqPV
44Y3XPHBMgl6/gQP5g2v7BcAvgq/8cSPIGf0gNxMM/4Ja5K06pauWk6MLIszZdWZ3XZgkf6Vh5c+
HNRcCjFlRiPR1CUmSov594ZTzXxEUELK3Du/QVlPn/LUp/5Bejt85K/djyDMEK+7lSD8Lt0lc+BS
cK6+deEoNKs0G1QFyO22YKNDifAREuKRQPd6c0rvCoTowd43/0NWP6YJATZHX3xlZL/1AzIyeUjV
d7nfP2bfpVPPBnrYl0+gOmMwGnr58m2K77iVknei5H7q0e96XojubTUPHt0tF6ehlxyO2+WrOH5u
mFtHdctSaPetpPPLRgCxq0dGBBm1Avep26pkSnIH1Qz1csLCGZFsfP3Cb6pVi1VlH6CbtyM+/p6D
zMyGZ9VFoz/krWLtQAoVinvBzWmOcnIIzJ4wrLdSC1Umx6rb6dSEZEkPdJLao1G8FNoW9vYSs1fc
eA7kINhaeZ8kPxRHl12YeqZkm+zaiVJAL46H3l0gp3XxVWkuoiOT6ag4+OcFy+vmH7byeXWUQqZc
VwvmYxtnhoBZHW/HDbAJ73Nywme6uDOo409k2DNyOWzPLlYn0rxsjNtWbOzjh37STSroS6LE97/f
tnyen2IphWq51vkFqMp7LhnTieNQeeq0dKY9zae6Zzja0AChIDKcMJFlAG94bOVsvPfe/f4db6Dr
sF+ciuIELspbf4JDjrU0aPut/aLlZwAW4hMjwXjHB5jJ/M36LDglJTpD8Q3fSVfGkv0I+h8JttQ+
o9jVqrrVs3HFbO6xAJuwfXnUIsNJFBKc4wwRDR1fYdQ2O8O2Xb9ainOVvU5F18llPYYJE8+F+47U
cLuYhBWCyd4Y4zuqdQV1NX0q+uxvekefvJ4VvCFVthwQ3TimDz4wHcqxMbybSsBxrhD1p06csLKW
QFDiO8csVKgv4hH3gRTSlujFWBOz8hCC49yRN3BsqOlBt79WyKvfMcg1YBaZFs5uKSc7GqzeFBby
f2V+6C6b/qVm18GEWL9p3b3ac9cNRsh6A6DihH0j+1Yjmq/s5vItqY1Av3pG9edcvHW6DIuQOmU6
pRhc9ScF4jDeD3ch5z8PBSH+aOlC0BN4LJAEM6ADNMxPWzD+vlFYyvfrpi75cfJq9iuZT0trThWT
bnGa5ZXiDYJIZqRQDnAjJwv2RPe6QOoO1nebsM9+ea7Lt1v+YDSkmCEyqE6SU35Ng2j5/yXtZNb9
wUTNS+ei4EwoxJKvhFG2VqRQy7n2MaiIcI9w5m9pnq7/I50nf/XqauJp4kYATDfHu2O5dA5EkKLw
ZIbJbm79m8Kev9RsLwpOzudb9X0u2l/fti5eOI+yykX7JQZFwti2hjzSVTPTpzDitoadWg7wJFEW
fkN8/43v4m9Y7o62I9C1uQGBnXnoUDbzc8kOJEXDRtvjVNTDL1hb5mGbGyPFU2fE+RN3/jeZuszs
7DEOIW3iUthNe9XIm6Q0dQ2HqEDVtr4wb0TGZd8VAomY0VwfgxOCxds6bCBY/F1Id+regJb5tLni
cw1vOXwFEyKw7JMcvc+MspErB5YJ2yjUOL8QMyYjVt7Xl2+6xptqkdJiSyiEpdT+vKwquxa/JMaY
dKqZGomx8mW67/F4auyiDmo49vDGwpEnTzUCBYV8VZcMBmo9EvViCPF9f9/pFIaHH86PSrPMzF6q
oMa1nZ7tIUAoHC9cWkvqcTKIHELA09JL/BGBgIybv2W49816u0CveVHGO7kr9HP+xgQzDg1AN0Ve
F1aGv+2qLuI0tPUSb5x4KGjJb1C7ZTAFnJD7jVpco+sGDx6889sM0M6GFkroWUrjDk46MfAWf/C2
leh8TVdhzmeYq5Sn+zBdB/zLdB+5+zdBHkAIrbuunPlyHq2YeC40a7sMq0q64EyA/BTAEMsk2Cld
FKTXucxdduyfwI9JHrbpimjhcMglyd89D1zIRYSfSADWH/YVdQ4lI7woINAIi3dcQp4GBeLGip9F
RjyN/AkOEfZZFweHdstmPQuV0ND5XtvcU+p6nmnIxwz1cP8dh8VYEoOqSDff3vUlel7qODMyDbiG
a9+gd8e5jxwSxtdFyfRMNFUOZuisP9UhOEXOq+mHI97DHFl9d+fKgXgp32jp/5I6fcNjsLpmE2vm
pHv5pWBqoIxk1XWjZ+YsbetqJqS4xotJBGUQyCO19DM42w8/f/UOD5j5lKI07gl3IgaeLGth0wG1
Te51JhRstsvNmIMIVsndcK5bSW7pJsEweRScfRUvTr0gTzYN3/uMmKzjWBsssfyyG8FUe/JxwBhg
r3SBMbsso5uRuf5bntI1QBza54DNBO0/gB/4tW5lg0ktoG2sTm+dCV2ipZ58BJ/0NwikXv4wB3oH
F5m5VGmpiqpMxTUdqtRnNce3voPFPknkkDlIPWvO/LyhE2NEjVC6flvMzzs8Ur4pdkWVgV3FXGDm
R8940PYJue4ravRN3fSVbv9lQscXCrAn1YqRg7mL/SuIL9Oj2e6DeKibt3bK3I5RFR5nrFJ7uDAv
F3IAI8w0BsWhQrwbmkrjHEkTnYq/gJce9WyagzbbmeRulP3OAxwf2ywGSkldHMZtF8vacegEgHEz
ItGPcsPRc/i04VKsDE5mLbhtMpU4uCJalEeqUkKQZoH0ZMa+tg2hpr5h7Xu9Pls9e8JEQDhCco8n
OkoczH4yMLoPxxF2E6W1nK/frEdY9MCTC+xidPwhazU9mOdszu8F9IHRZDVm5hBVEX3kh6vCmpMP
B5/mOJNkHFQ3QIXWnFB2SQM1/HK6SBHflfQNGiOCVA44KKkQcDunh8l1rmxB69VUGojfKDpAtJ+p
WHAOkOb6qb0vyrWB6HNxm/Xm/OHAHya05Z4/f9ANw8jDAjg9rFRj8+oTTuGC2Vk/7GXHaNCynYPR
m/ZyHqVGGuajYXATzvo1+lrzeZC5civIglBrorhmHOT4AG36qu3MADjazKGRmwxfy6we4pawD0FY
0hMcN9CEK6r+AOvnPCpYIC6VOzmx/1LVMFlemRR2HpWHTtcs3NFZTLEz+uIdZyNp3selIMe7TBNE
NBlQVMbe6re36SBTo4kSaD8cExpl5RXgDpmV51QzDjalDyc4lfo9PCzPFbt88DWiJtTgD5/zvsRp
ZjzgJ7OXo6d+DgUeP0Dy7UvNUBI0qDDQAYXkoYdVwSael3ytquIG+DLG/Sf0dfyLP8oe3Cj2fs9S
U2nitG+W13FFTMsCny5UmiqZQsyPtf7HRJQFO0JvAKspiqjrMjOV84iDRaX5wgb92LcR0R5ls379
DdZisB/vPIODv4MMgvtgKiorDpRXYDd+D8+kVJQXeQh0PDvnJI6Kn0qp0MegcYf9sRwWe4Sh01Sf
Z5e/jW0ygInYRQr9GbZa2hgA9t8tCJURAcwUrxV0nLkVuR3Bw/ibXKARuKXZPX/ytxw53o0Bub/p
l+uAN80mgkJkqIQlo/R0sx2g8/BRlPlt4IDcK2Zx8Oc/dl+Oaythcm0/JgcmNY1+c22z74yNf3LQ
fhobdP/LCV/omtU3rFDYL8/T6zmXhLfCNsM/HKHXm+wH+sWDD+V5RbZKgNud9IoS2S5VfhCqGrbO
/DOSA76DEF1ky7J4tf2+aZ8H5LSUGI7M7va5spr131VsrrS6BC6BeFXyw1D6nJmVpOCz7tje308C
tw9BiaHRCFLKhxVuaxCiLvdWHncHlo/Lpne6UFIfJDZM04h5r4NdA6ayvwiq9bZbvylaZbx5qH+J
t4JQvG5Z9oj3O4XFUQi/vMfOJnJeTRTB4f1Zih1d/ZUaHnCtZQogqAQ9zVXpVyG++aQpEvv++0dm
5+ndGfHMXTq3zhp/X1jZ/iLjr2l5RCFlLUo9dpQpJTmXd3p83CWy4ALOTzb3xT+7tSm0lzQ2N8dY
abZBUArdNojfJLKO6e0wzzfyzJE1eZHHdDBJWxtDC38XPOhUxB7Vpw20Qz4WcJBRymJoA1do6jY7
VIhbUVGt8Vyo6iNU2G0TRsPWWViTVzG7MN5tC9+ddw0kOoNWIBtQHzu+ylnUueOHS8op2PMG9SfU
oq6nZ2y8FDWMfLqT9RSJ4plkP8Xk63Ck3FI2x3aPxh3BxVQNrUm6EpWukTzHd17Nx3n/2iD7rjZz
QKjabyYsoXMZnvmYn8GTvvhEqZ7lvwYBj3ILIOsYJ4X93+gI5LQycADHyqb3ZhiLQ3kZRXe52DEn
xZKMx+42x2dTFwVLsSLBPYW45IiK15riZrUlPG5RztRci05euxP+/s/dA3N7NIEaXwEHnr/w8f9+
1RCQ7FhB9pOx+JHoMj4HM6i5W2Ym9jhD9SB9RR479bWgwn9EkGDkILvx5psP36ZF88rifLqAmlh8
6nZ8y5PfiM1WwWT05aaxJMwnzQD4g+8pj+km9ldzWocO+Cxcls7LqyMynGnROZ6QNrk8++UH+quj
wG8HVpZkcxfUueC11sL2Kc8z4Tgjs9Ys5Tdjadn9lOA6haIQV6C3ChXXZTQ0J4irGSiylecjpfjP
v+PluM66AyKIBbm+Dyi4avJ8M3HDbu9vymdu9B04GP8vPgYfhcOIUTrD+PBPvwhls4W65R2W24pc
YDR4MwBv/wD2aEVz4Gp4IcEWRRwy66qMk82HgI92Uewh03ltERSZ/z8hyJuXitVy8mSWQt5iKNxa
BJ9dy5hJVtbCmhRjvmKJ4lZ+BV0pIHytmuvQfjBYmaLHBlh5/HYIW62WoYoWHk4R6QNjDeVrGUCv
Si0CB+FqYVQg0vBWXQl+BKi9vpWNkJG9dtjPgyHujsY5X2roIpZHebfBMhapBvdXmT/u+wr7LYIM
5fBkxHWZEsrRpEKTc/wKOKZ+dqwY5v10Xo1+ymWyxd9nM87pg4yTIKbQuWN+lZXqlSwinXCTUm95
AkkNkT6PcxpFDZDFthaWWI/sEUBmzJTeNmkjyS70CcIe1Nh4oGYYP3O8dIl4D4B/q3+b4nWBINyG
hcaPmFv6smBHXT6nwNr4pqKRSGEWkTiBSMQxqdR1XGsn/6vlAiK6rcm7l/kVU+DlX0smMMczKuBs
O5e1NTzpBaBp9zcF8dgcLgDNW303JZGx1a3bCY6WlhOeVNNvr8kFXA66C2Tg2qQ3v9+IKToA0wzJ
pPlR5qlVogJ3/B7rRWdO/jl15gEHDKgoV8ESW2yf2PCdQhXp+zPp0INzF+7SmUGU4KElHoGEnbK2
mudC8aUkC0vWfeL5r2fd96QrFXm46qghWP5vJH+2tssu4zbMxUWS1pBx+w533ZQwp3JTbZmUJy/d
Beil0h9i26L/lFqFMqzFn0NSN+4gcU65l8I6f5JFRugoVHm6gygAz4kzQt4LPxD8ssuiNsVFJChT
onuCvkt52PedlZ9pVjQ/H1k0+Znr2BV1hqR5BZIQyXSyYkegQxFNVI+TMVR21D+iMY/IbS0tc0fU
1tymuJFuU7B8QJCD0IH5sn1PtSfI6tiLcQiGHnyCfh56OI6zwXIFirRMu4JCXy777/szZQt2A2yx
D3SwhVxwGONWGF9HAlXV6V+e/0Ruvktt5XIRNFBRjMDbAXTzznqSD7/CfOFRH/TWzY9XEkSB/Xxu
m+uU0xIR5kyrvvhi9r2t3/hmbww4Ly8WtAGv/8RlzKmx8maUclkFnCQp6itjaWZ9JTtAE9gNjerS
tSjSLfS6Ule3BHeEqJ+cML/F6qbML/UWx4LRyp/WoooBAbVR1A+JN0dImvzmfRC+tgUO9UOxrN0f
dNXPRnLYfjND42DpOfu2oHycgOeD9u5k5vwFpGV3HJxOx67DruI7UJveR5AbaHn8ZoHwHUFAvVb8
nO/YAT4INqiN0qfaAQQgGgE/uVK5EnTq3eTAlpHKHIdg/UYNEANKcO2xdNieWvZXCG16IT+5tusm
ulBO0zodbGPgEPPXAhPia/oCqx5VYaVKinJJRilkLedsBXJhSiqmccuNna3O2EiJhYUxef6fC9q6
GOqY0jnwaHMBDfntlJUH9s0RDwdWe8gQoBUlENd8MCCsM7aBJRRtKdy6WD2RDLJsmkyKfA4OHhYB
zUYs5vQuWCn3nIFL5pdOe5q1iHmWjyN0v4LKspRCLMMe2egACoHUOgnpBpE3dh9tV6E07UWOFs2v
zLU4hsgc+yHdELL/o1j7ynGRxNIeaYDSpreoafgZmViTM1lc/SOc6nuAGhBzJj4UUIYnFk64S9DF
yOHP/3u7jW0jBYsmb7cGxDCYbQezrqtRSZ8duJTfvsQiCLQkGMXOcFAfCxi7Gl8EUn/ejadbvEtu
KYJxMrc0jjli2ny++vter9ecAw8Myu8zSCAS/4Vl0YsU9jKZ0OEVnk0wv1Tquj8nBIRBWKutDt1i
C/wYVBs0FEF8c149y59euulTbEj6RL+8a1xl6/2Ogn5sA9ycDcepG96rnOIq1Veg5sMLmhbolDED
dlAuwY5dFiHwrMgyTK/zItzfSi4PWYCsCpZfFHr3c5Kvg0h6FdmaUklEcNJRJAtl8eOw7m7drKKO
IOr0JA4OwoK60ynynU7XXIZGuK5MOLA/wSwBGGRX8SXaRaxlVyE6jbjoHjeKfjMiFaK5ntoLb1fH
pXkPDagCJH+K2FscqHhbBJpXiX128Ivn7lZQIyS1+dskhCdeP9y2irA9xkQJz2EX9UUAL+kXKvDo
V2xW2JoGMIPN6EmgJ0ukBCV68Jyg+WAt2LxCrdaP7/OeTmOielQ3JH65UhFCYrvWDaefRabw5bdx
eYZsxjtKGkRWggrpM2bdFba7yZ4VdRX7toiD19VEvGKdHSJDXuiZ50Sr7rVghGOpBnNSA0SRLgq4
ITyc9j8GJyIWLZ1WUa2B1iOAY6FdGHfqPmnSQhwuGJtSS/YbvgYtEDUuKfFIdoGY4uJx+v5M1bWV
w5/c8wircpZUBHfeHJgQfLi8xzSaodF7Iy7VX9gp/a0O7NzXE16zChhxsf8dvesuqf1he17mG2Nx
BtRD3Q39aU/bfY1ReEhWPcQELhrRQNybjOoOHxaAR5JVG5bDcS/P87nTu6g5WCYCBYkv3a6xiBzK
0HmFeZFlrSL2MKQoTfBq9H266TWhhadzo3C0ILJzdmewkmx62eyT/XG+rU0kM6GfUMELznTv8Wz6
+z5ZpQ0slsTOiv7D8tT/XPb3wAeXqCX9iBYYX5gOa7bhmxmhbbVxoxd7CDcNfT9R1YktOJVEH3zm
8d2WwFLEiQh5ctBIo6VKCLGYQIJMQKefYOvbkuHV3+KM3FT8ztEiRBUS3FWjGZGl8W+bfjLFMo2A
Zq1/v/OKoMCNX2SgMGBFFH22RMPBtivJpu9dDpaIT4v4FREclj+V6K36ReBRgPKM15Lm6cU+M5Q1
Z/7H9zejs+aFqmJfCPzcxNRmiJS5JsK7NGw5YC+qEtakhvgSa/wtXv1QDpMnPL1DkMQ5lw0PmWod
IUBoisxXpPR+e1IhffIdCUOYZyVDQCzlRi4Wt09xg7o47YWcC0EwQEpeuzXOpvJOHpbdtwVTWOUt
KYRb38IJ50YEZV48NYKtv04IklMOfoAEAi24N4vptVreNrdLvgzrXjT2VYnvJaObgVvtWRLSWLBW
l0hF7vyk4HhNOcEfDi5aatUkXShRZKR6obWCpvSoVCDIyrSrROwUG/2jmTDSbesLxe9JwW2ze8uk
rlJ3UEan70GPtyJYg78c18aHwqX9wTPobil0JEWWGh4+JnQRG2tkrdiZBT5jOfBauLrxiFImSHOb
4PlE+FpcvF8M3HttmWbV0o5P3xUdRsWdM2Ba7CjFdD1VCDTqmIatfoKySZ0M5ZbyJ1y9fsJxDaqB
FpbX43+YaWLZnF+B++0L/3n9JNnM6bT8t9hxqhL9xYxahYtTHGk+E0MHbFmVzE37lGOQMxuZr6rs
pSo7LW+XIjzZTr1oeZZbRB1eObCrMvSOaUU77qow7mOw0zJuPB6z6BJENDS/geHfhEUVeAp5Ipes
PWYsr85Sn2bco50P0WKq6H7PLI0WHGokAegsJuIjPcXHnUKZPytdxXZgGFXnE/DRkKZdCpTjHSmp
yr8ilLiTXPmWKbsedYPiXSYG5ade3CgSDGh8bDbWMhlHmbVfo3rrzR4lSZppFerOANk+Gn1GLX8C
W2j4UfaIO/uD7SKa+jJgqFHZTYOYsCiUZneyIQGf/o/q76T5eyw+l77I5BhGEGIVVp4B9fZaD39O
PkUT9LqsjhUGlR2aw3B9NRueZ2Ui3YaNwgGatpm2ftiS/8d3nfq1vdSI9ICB5euaKgAQ/EB1wI04
iSl3o7xD66PJFJS1+4IcieNZV5wdk62QpiRl3JyMgZj7G/t23sP0xF70imEuqZS94u0FfFjC39Xh
B6sbtP/+2ERK3nr0Y+rYHzlzftJC4veY1e21JsnfBxTvY6rXbGxW4GykA8/St30gTSEkbNs0Y69L
PbspK3FILbHX9DXHRw57YM589/WmP+jeM1EOsW4P9bnlUdbXb+P6GQzdohFHI6YrilL7cVIhtCbd
+zMnsGpMt+HD7esvlbXdSS0ZU6lz5LpiglRsg6Enwk1mTx50lPJMzrsGxlKYb5IoY820rPG4+8Sj
b5moq1H1X7GxakNq1PloturPo5087h1+AAfS6Rup6zGzGSGAdGiIBSaM4VCg5s3WntaXTGZfw4Hi
f30iNUxbQ075rb4MC0vfEKOGH+obIFBWX/lkYuZpczmwb93j1g3dkE++ceyJ3v1up45myTWdpHxM
OE2MKC8/w0149TvxWQO4mVzrLqwFetv+pm6qQ9Tw5+Iof55Y2e/T6aMYvgqj/MjgIsnqgJGrLi5x
xk+Hcf2YJfzadhHwRhwJ2HGL9K/cpJ4DOerAsaFUZmDpJb4/J9Rss5fCEo83OneDc+IVkCXATs+o
vBjwn9R6HDxuAAC3achR/JMSrG2amAMjMMbiKdJ1htZxqaZ50Woj6SrgOhVI7RxMFzGxP8+v753Q
VPr6Pyv48o5AA7iAgVg0Mt2BxyKbmYP6IypvnIJziJFHzt6Po2PJbYgTQTC9+DvkAvpbRo42jJnW
9AjvQphkavlBHlSufc+7sLhk228ZobStIGu7eqCUhsLEpoaDBOIbSvg3AD58LJ0ynwi+XhH4GgnO
5RjihG4qPy1SBv8qL6AfwoLmmHrZNUsHW+Li6oRDjK+hdXXomxHraWIbhyO6zAhLS6YlVJjovlOz
E6igM+mcUZK36s5mfN/4emhuvzMgv9KBWqCEh7qPiNECC6cnEbavLq379swQV1Lf8ryT3rmPA13Y
+tGbRgRiCLZ2mJCYYuGGNkwa7kZAEwSL2Coa351lvWj5MAlNZ/dCtdnDHP0D9jCTqkn7Vo/45Jcd
yrdMi6csVzZKufGmjLd58+v23ubXNche5ngKqgG37q5dtkEna1dInrLeY7/ZK7LbIMTiLIeGT5H8
ISb7lRtPBPxqZgZx116lUsuPK1H6MDh4uYaU7qybuoBGITfYnEdH9VwtotyA/5kTjVk2FDCynHxP
ySfAdDeWL9WUQqez2OcoUFyHH83l6Fmv3ZNl7dykUeVka1rTqgWdMMdQMQ8OiX2QT3hIH3ywEp1i
BA4aVFYRNEJGVI7jt6kLFp+m21Ag8zq9C0nDsysRQYNmdFG+76GQ0/Em/uVLSLYC2wqWY/BzTJQo
NYscXpNguvE3wWpbqF8QT0/McPw9A8mp0efCa3BNwA+7MKxR+k30ANbH1acmEeT9/ngXPnFCtPt1
po3qhap/Z/jhGkBkdW/zl3vutwbS+D9DY0W4jTJNTcj+ns6wG0AOjlZHUqk1ymEOnxMtKO5OQT3P
eStdHC7cIDaOmL0lpRnjDOTVyUH2LVSZQD65QFOZID/hHm8aQMAsMc9J7YvslcuF317jwgkeXEWT
cdkWTRb4JqERim4BkTllG3OECKojLi5B5f/QDzVrmsEoeq3rvJxrAGCF83fy1UPvi1ZrXpIcSfsc
Ih0M2FWoE/w8ftdaqf+lRlXRcULkJacAvNmI5/VKi1RKCLSo1Ap9ccOqvKwXWWwYRlur8uCS1TAq
oP6Tqplk5NtgJL4ZGj/TAKiyfkpiCBVkMf9vhgECp/czZdSCkLGhIitwccVdCo60Tkhpu0SiC1OQ
cL3uwrDyzkYEPqlBdMO/S8q6wqfGLCMRO0ufO5yBSYPEPBaMPyw6SJ1IMr4h8XAOjbV6w5xs6bIy
3vgq8aVq90QPwhnhhbNAl/OEX97mi0OWurOGwhnCYWDubi+VQQgGr1i1tJMBR4ecRD4sT7lbJoqP
rbCLrfyNtwKI7re4LKMdsP1sR8NXXic0GtCy11Fc5QgWrW71DcOoO8mXENTlxI1oeGtrtSzOfhiu
RIMahwVqs3RQizu3dx5nUwqA+wuovqMf/VzQW458bWdYAjfkQTXTDDQ5uSD/KcKALub+AuMzmuFC
R9DIIm6tmrSEwDoyllLURNdiXIsxcmb4ezgygL7SnWrr7EYvHY2T/anenOGBs5nrsgn8Qg6QOkUz
AIkjiHzFIsb5fF7pvQUg8r+R2Ve5DZATFUBiD9kRejEA7ZAS0QqsYvRrSIVuU08s7j64S+ZbOtAC
zR6dUjJTN1rnxjRO0xvfJVUX3HlWyTxRpUGJcJ3MKBS8PvYrbcGW1xQ9J6U0UWpKOZmw/pty1R+N
NZ+dKkkoBAN+UMc0ShK4sdOW8qcLQj3jfzmcgycOMJEgbPrL71Ydi4QA7Dn9ZshrXH3sCYotun4X
roSrLp6k1L3F3cilZWN9dP2vY0zv7CnA6ARuHCXIXkcfizOfbot9f98ac6+A0VCkdqp1OY4ymYCN
uEvkkBBylCeD432ozrXxIeqQv/iexLJA/+QfV/u/NkoazPKHFDH8C0kBYcpgiAG8UHCYgYpenTe4
jlnPJHPHZ+VaJ5iIXVKt+RksPzb1M1E4vZgHznxp2sHeZg/B0nDBeoyLVQ4y2u9jxoACLcvNLH1V
mSolZ/puhnn1GI7BlT1IFpHUTCrCVoE84w5V8lWTLqdwb38Drjgxkx9QBJkHRi3jS1piYTXWszvE
VX7zDgfENxmb2UKHKZ6kKIWgOGiH+dtH5H/CqA33/ZdYYufLA2PvBtkp19nw5xW0NFey3aBz+a+y
FtPkGnsH4fi9iNbvNLdIeUyOr7Efbzw2n4a+UYigk4BzRjVo4CDC170wMN3ZDP6eh1vUVjGglh06
D7+Goc1X/c9+FeDUo3ptqbe6NUBkeb16/EzmZkmktvcxqT1dzuN27PyU/myKO8JdM9ZZzApJnSDz
RKBIZGcslVOgbpMHqQNhLfUQaYLAUD6LnBvBCNr6GV6Vr5TVXRPQZgrNrZOl7sJDzndoLOSGs4l9
CmAV9xcIqQk6RHzXzKgH2+/4gZmi4sTpyjPwtff5+zqZ4jrKg0LwSf2lcFPYsEBSmYafZpRYfFAP
V9V+VwC08MUDtNSlDdEXPcwRtc8zgmsEeqDmlIlVtwkq895Bx2lfK6H7WGGEFHPVGLr550gOCxHz
xIOcA9D8MtGNCJpSvF4Iwmbs9RucLZ59SsapDAtACFRb2bXlEYiwvdlYoK7PrdEqxmr7zyaGZg0k
QVqlS6KPMJ/TVV9u8K5ocSNaKaS1oAK1Yx2Soyn2Azy5qliG6kUiF9nlQbuFs2KKvyXJ7C0jMIG6
IISlK3zKuY5ZIEI5HsCWUc9IdX9F93u+siW4CKN32SD+QnPjjhCELVNnsFNkT7lX6g8zZhnDLCYc
aLSRdygNFrBWc6WML9HMi5EqbhoEiSL0yY9hr0js6VhpGNxsn79GHhcWsv0mRhre/JmqZUl3fS1E
VE76SfpTmg9MtN9mEDNgKgdRpt0+vvtX0nb5GrLHkZNVyuVf4Ie2yTbAXNEBh8BuDTy/ftbPKcG1
DCP2a72RafSwNkrQgwfCw9W+Cx1XUmeZj6AnesQhehKeh97cmyoNsV3H/Xa8SWHF4w96sjxoM+lP
0pEcUJGJrsauGokfYce3/LF2rTuUH7b1J5y6t3S/TOl+RWgP3xC6Ey2V84UgE8RHqa/BzCb0T4sH
cbF2w8b+GSUayUt982ybyC1q2zBPAmTGaFB8OnqBa+1l18nN0TCkFI+bCdv7lmuXRF4HivMTF2Su
Q/G0Gvo1GPCuQE3Xozfy2I3vUe5SyzpSfG2+IOyenoRjsncXPdDrjyzLGXBoBSu83Ukw2S/CDRQy
hbuvM8dUDB1F4FlVMUg8JpP3GvqQ18LPJFZ1lBee39ndIGVRU3m3XD6/jJ/afKhYqkUr1yrrowQy
tGJx9PwczrcSmZaPkx3I3zxwFRtyrAPooFcEe9SmfK229YHyF/9Hu2zZCSfptedrxm9KrX3qrjBI
mfpZztLx3yIDdbItMLFQmzq6kLzaHBA0p5lMVioSxW4RNRxGEACfSHUNA5dYPJnTnXfwKfpzy0LP
KF/IX7R9R6FksDZry4xgAh7x1aQF3+aWpZi6c1GYJczwEN4TBH62Jzh80gS5PRuREQLnwZpu270B
0pyVXUoxeED0GXNVhif/0A4Bp2zz2KbibnP3LXyjU9+S+xjB1XRNeWlvPeEoP49aCOlCV2fFkmPC
KhvHpqZxpcM3LqRzvSEzLKf71mqW6n7r75SAFylNa3kxTvpOYHeQeIndR6vpvYXLp6zSi+HroJu8
ATG0B/kzwXYT8DAob31fQrupWHCGTPXecx7KJ1bhLHH+wKGrV7QpX25Z1qSAUge4HWg5YmsLMBDY
trSMiheE4LbASPF24T/I/TciJ/Smwx+05RhBEZA2iOHYvJk0W9+gNIRJK97Rv0Qr6Ia4PsBB5xKO
Q5JCjKXiUhttN+cKDmCGZlB1H34+K6VKHqXAVs+uPLu8vpVaCfgu/j8xHpkkS8RFaBoyGBNTLj9L
SQV94SdzlaKtYqkUahNI0ILYJWLkXIcMoXW5fe4Qbp5ZZZD24RXaj/2oIaMsCD2aqlq3qqr58xvy
RSymYYuyyVRBxEkYbyzAZJbZ3B7ZhGoCs6hNz+/wx2cXXWGrbP/ETqZKZ7wLTVMaHY0hg2eBSzdC
gEpZvsOFAZlsk/svkmRtS9M62Mbx8tfHvth197vNRQONaVzWxQUvVmbFaUZ1kh+vqv7O492n9kfK
rZIxn8d46k0GZ5szQlyMwp22YwmwrsVpP4PEhOs8CKkFTiRK4kOtu4Y6i8KJmjLvWnFqZrF3Apih
GdWQLqq7NSGwyInxXaWKxhHLZFQ8U8O2+svOnDw3vLeRgo058Dem6+/UOHKL5hV4lfe/40vOpsVI
3Lj691SsPfKYImXEH+6AfRxjbDO8zJr6XYMSefrGi9++MOQzpLUnJm1xm0OC0GyMEddJkBSQa61U
zpBSRjC3cmwAF0zpyNSAWQr05MsAyLBeWrSa+8kq42+MKm1tHEAOg1ydx0nQuZRczJTFq0JgJnUi
xK9TlFEbodzvAh6Az+UDYgXXsqNXfo/Tze5jLPoqbuJOV74CLp6Qq6jaEfsRIEAXFPVBg+2KHQXR
ywoIu0XZzQQPDismdOvCdh8mI8RrhaecWY/VRXAbD8jy5bQf4+0YT6maJfgRmWbn3sp9bAcTxtMH
MOzaq/2cvcli8CvGgGqymlLbux1+MwFf5IKnekKikYeuyhh8r/SPezIZDoIbO6vcFpO3/P+PZv9L
CKqWBEy0EHmXl23xEnI/weGY6jCTsFM0ZJQVpZn8tAVNHlwwiGSO/RfdxuydMc9WYJf4YdZbVAUs
PA+TB2aNXzcc2i2/uXfzCB2cva2Xz7wpKHM0LxSAfUqCxCeaSNy2fYD7xuhINy7WWDJoJQRbqrmY
43cIKvmCHXeLsogfCPr5W439KLHmPxK4nJgPQou4vj6f71y358dV8xXZJX323GlyNQwM1cW4DZVJ
rbivIFYGHpNlQhUyWnOgdq4JMJnjalj2P6dGYsjVzHO/gFFEWcCJYdbRkT1OOvWT0JorY6L8DUf/
p9z/RHrnvugYr1l5jh0xyyeG0g3iAz46Aoxa2+Y/4lcZvbOE5TMNf3I2sTk3UEM0+K6T4zBz+iHp
P2ffKEofiq4HtiBpBtsj4jSknsC4ySiiW7gmZJCSP4oIDpFzSp6lEcKwK9R0YiNyfBnyxr/nx1WZ
Q84QURcpbIEXucdI/yEjHyFfskXGbGT/XF5crbO3PQ5jyDjZu4oaIq4mifTTyKmGMJc5UW/y0CCm
uF4A9cWYTzogl4MmtZX4NXIy2qbbzWh3lfvcDbQXkon0Pw/+rDZoDkViWemCUkxHuQlcdpOztJTG
XcRKIDHJhx3hqS13s7Zmr2hWPB2bEqv5xD77G0oJ6sSFQ49RThdnL2+L7hIcLQh++qDdmbvHw1Rg
NTi4XSXPubn+F4miraPcqnCPklwgyrOpsOaAiLGHX3fjSh2/ME6yTQmj+9L2yh7JSblDaU1f6+hW
5CJqnKKomP7WXsKslFbVktBaL9ZhglREKFR92m6msmSp0i5BdwxxLMhjY/LgM8KF/djhH2kldOjh
Kv4MGBaCRqzGMbGVjU7NhXP2Jp6F02DSroN4s+tdi4+c1HobeJcZ7k5xYaiY4KuEITYlJ0quYmvE
tNqyv+Tu7T0nKuabQ1TrRb6CIkxasyehxZLCI/vHk0Fq3CYSIzX6ZHqGCDMfNjzS+S8d1QMdBciy
X/YwRYENJ0QMi3s5n2gGof3GsW4WISQGhNdWhfLSU/VSiQqU/chA30MNM/DsjFsx2exJxbh6HDmN
9jBpoDkOjZ5F2085aF21wuD8gVp6d8p8bvo0JmgTOpOAzoo2AB1DjKC0VT1ADSK+GOFWPrmFHxPy
IwM0ucwYPk4dtSy/lQyOkxGvy6arUTl9WaMnD2knetXl4sMfISc6k+aitUgz+wJnqMkItSxPViNS
HKMKon3+Wj+p5nm0WRHtSM7poUNGauR7eY0leF8bC4BY5GGBVD6dYMv6oX2PFUBjwG60rV/dKkpO
vpJNNWjaQVV59GIWXi4w9dl5+SSuPUzaiunLZKwta1e3QwQReI+vuzJKDFP2bo4tHhS/edgu34gV
STnkh/lW09f9b1q8+cdCsX/i9OuiXJA9yvuKVMGHeBw507e1iaLqHxB3iqYADWcX6Ff126Qhph4K
TWeSryjHX7WsZ8ShvYZG0fJFM28Nn9Y8Dio1oMeupw5Ze19gMnASjaoAOBFpgrZnxOleUo/JMwCQ
oNtKv9EyM1zjt/o3fQ2xA1EsZhEgWak9DmbnylZ72Y4EaNoXQJziFQfYgsTjsewKkVzzGmS7x3JA
nFlCPNT65Bqjo8rH5JLns46Jigua3sjeCnGOryasCgyd09ztNR4A+hV7GKM6QpHzUUWPyX+aLZUR
jJhD7dK5MITKRDDVGR41IVGWFVckO/J7VHG7lXRTehds50/a7w3qKUtD8ZBn0nk7IXPNV39crVER
/QUPrAWAZPFgf1hJoAnOE1RRUdZ925C2niIioVqJq0d32k1qQSxkim5mcEuxERkqhFtqnV5/kRSp
2gmGZeo2nRBky+uyqJ4q9uLmAiWRcXcDXqmaC+1+ZblVuJ0IjJU3GmI12Y+lkYbXAXuHOTEpnu8c
uKfpJwAiAqTiuaX9UJL/ml1xLRpxza/2hFmLIoNLljXP76NVMGr64lkcahUe9H3l/bb3oufwOsPG
S+bjKnVnw9YErHXB4tr8LH1VcarodBVUza1lEbMa05nYhtTUJA3GXhSfXxnCahdvvJDSDSgIzkFA
CFqEdK9yqvzYi+1kFJKEa5mkts+5d0/0WUAXcrUoBAninbBztnEyugRw7m3Siz5dmRktveJzcIbK
Ah3bBBir3QRqNDeXqc7BBnjOXMONEPccF31qAgQkE+jLg6oRqw+v4lyRTSA27DYosrNELL7Jb8FD
G0wsiE2Xseo2NmEeM1JvH5dsHfV/WHqsBuM2/vbXOMtE5UU2voUwW+OJwSGcasdlFxLdvcLgsgYF
fyZh0nCXHItHy0v+1GYi9yN19RP78kEvZDhYpwGXaBfT4wASDi4xP+XlmCQgEfZONQe+E0zmkDmN
elNeE61AzvVIz+joUAknjrfTs8xrsukRGcxHe5Ow1X3bhxL07wMAW8fNhKuiYzTXDAtE5ybKE6k0
0K9Jr9fJxj6CBLh5SPlKtb2fLylnBKidlHjpIDNvyTpa/OICiG0k4aHFt/T5EKQfxzm3OdL9WqcE
p39XdXW4CEFTIn871EXp2O9OF61ZuolUHxXzIShkQj+46al9jDyEb2FUeFv/aEQrc+cVVj1EtkZ/
DS57CtzbUtux/QEsyYVofHZHdWGfCNNE+96Tdq6nY7ZccigEdq+1DIPY9opGNm1w9lQVZJ7hlTaO
gLeaR/rIVypjRrfqds6ZKAfiRk7qIqa0n2FbX9TTUhQglm5Nd23FNOFR5vp/D1Tt00fZ6cpkw7Uh
eS/OPM/ATFK+Edcn+XFCfB4RE+5wjkZOxg4+i0NgCR400rqsUTbkMvlxPuIEafvNBFbSDDWwvMw3
ImaLZpB+jojSeVBjPmzIMqfhfeSpOtBRzVQ+doZX+j7fPwU+6/60LLc0K//cl8b15b4lgFmGyMwK
dFM/kBJhCueo1AS9KxoIwQkfmbnHSQaC0M4TE9tQv8Q/9mtVStE7+pl2zTiCq+RFxgPaROQGiMT3
24QOLvBVZ0mnbwRF3j/hrD1rQm8ni5qUYAtTWTSRm/K9E6p+5BpPLeDSeSIBrH6ArZ5y3gzcBhzV
4nZMUTtafKI8UxIpJm2fxnhcOtlNgM+iFqmtOkhcQW64NP/MNJbqnKdvUDS8gHYD4KW7ZKiyg2HZ
H/KWTTcEYRndT+kGJ+tGZhrHCZb+PQauxBWhbl99h9cBiSGUrAWR+EiFesCwz4hHFDIFGH10M0ok
P+cttTT/zltzjZrMsjKjvCgJ0WWcjgRHjcHRtXPwugDyqg6UNlgOoh2KA+S3oDwESu9T2gcSZR9z
BWpN8SNOtQd06kZVGRZY4n++o2HCva8SBBYWQ3q7jLiVrK3NwwZPnb5wvfWr4CAle8OeeZxva5Jv
JRUSFxRZh72PLuqkcVx/XgFCKgSfgzwxSPdc479qmFRqjfLV+aNRKh9IJdKPvpdqkFeI7KYHUuvT
bLKXMVHwusN+yRflJ4X5MT9ZQlayjsH3rwusxAyuUihlGEgf/YLfEAhwusD1WMhO4vGgwSuT061J
3j0AS2uYN/9wOtm2u78EzI3JFtTg5KcVXWGPVO8h4kGqvNkq9N+gMy9rXQ8EzAkAjEsS6GULOFrk
zzwvaEE29cSasY4vwIEZbEbx1lib7UZDnxlpZDtxXVuHymJTQ4JysNBDfvKJSOpvY1KADbRztpFj
vwmb6bd6ToBuFF80ODRxkLQ0G5uRIXo/8yS0ObeTxEdfkfbG/VRZ67MRWUG/qcTDd7p/WFmdvWWD
PCL9kD+Q+/D6Ey+DgY8hwxY8g22tH0W/ybC9wn8FgKUJ2P7LcIh7mLH+EYcPwOU7GsINseh1MuzZ
KhfL9UnITvi6+L0JhNKqHqLnDF/PB7vQRPyGSMSapJy5P2WPKDxhNcNFLUhBqA/WG44t8wPjQ8j4
Nmn9eSCwzDjhBlD0Qvrvy7POURAN9uGqGuPS50vNJHrx7+BXXo7J7duHA6Bhc1jlGdF+bNUUZANg
uJIqrkFBEQumybARWljOcvHnJFZm/359mXi49CT4aJAEBiV8PzRHf3YYn8NEpWpQWRSA20lLUZrt
y5/3uTTnA2BncJAnPQtY/iaZerlwV13SzmJ9bbv+UXZq6gufkFG0wnJ0rwtWisUfqA5P9uWBkacU
6GAS74wzapT0gQ9DWyhJcAirgEK7TEZUbZONVcOX4TPoJemX2xfFDI+r1dkRNaSFHKEbg1S79jdf
+J72XrlAq3/s+pvSmfDUM0nXYWMQxu6Sy5bFPatfsB3y660AhrXrnbGvaHl6QvziwMP8+X4bhOkL
l1678CWUmoQfdumXKI86mqDeEub1/KseIGWUwuzEWOMBML0r9m0Ul1UuxB9OXJnjyKKli/S6KPHj
w2l7kCQHOCKdOVkpWPqEkgqfPa7Zr/qsRBjNDR4uP6gXzRyAIcESIv1mXkF3w9i6mnQjuEluXUCG
Uf/ZwAbeenhAKZhat7WR3wviP9QpdNGHf3ZTG/EERyuG6aCDhuWycXo9D9OUKkO0V225rF71m0pF
hx1/G7KZvCVQU6BPajSg2+2YsybmWu5lPQSCZz0Kr0xJ42TIxrAaNEmCKgkGUeDTlgX84oN4HCDA
LB+zZm/hrXlAvBBX4rwFzU/SrYtzQKfxL5KCjX8T9QRxRiogFWdnmEpLbLjqbRE1174tQpCMUueb
qjqakoeh9rHMh2qfRV18ntadMC0dd253qw4+rhjj9YkQacLUQb4BPyqX15Y5wpqAQSv/MweStpHs
ryXgLyh49FG40L7KEUlWfEThGebg590aQ9xTgQvlDOykaFOklZE5J2jTwC5qbnq9DXGjs9Jlcwkk
/tPd31Q5LvqbflyoSSPZ8LSPAR73BjVZyp63N2vzzA9HSnfYSVgeyjKkTOfX9WpZz0RHwnT7aZRp
Ja1o9/krQUbtdNPceWQz9t/57f+IzK6lQr+ou2qtrk2jpC5ePo6A+rRs4fU1xLqc2TZ2nGJGn+tL
23H8x8fzH0vH7jPG2Wf/QKxS3TRivOWo6htShUsLn+TAaEYAKwuMNV8qlp5A5dD1GiF2d6Q/7L2A
B7yImrQ02vlAR9Hw9nu8c6+Q9OhYqpbBQxJA5RPCqGTbh8p/dzksGymu5GvJyzdm+4/hBI9Iax6j
MphBCcQheaR8sq8NPb1ZtXPqXIz6LD/9lER3sL5+HRGYk4nQ5ZqK7eSfwMognWGNB5JzVAR+JtLq
ZUYEH7qTofWrAS4m5W3/xwEfbOxsCtJIuXDI1hwSTWtj2xYJGNIjP3x2crv7EYqb7G8bbHL8IKnq
5KjnTFePr5NQAd5q+pW7qvjD67ZIebTCbLLWEqso3GknMT5w1/bf/NLFkoXSkegFJZxBI7tVG8ZW
mG+LKvkeTc1Ezy9n0t3vht+cvgpGPOCaLsCvz2AulAqXmsC+RYgujIP80p4ca43WdUeMPtqZMMe4
oqKkqmfusGMir7QtT06ENPLHPg4pXwiQTK1SV3GmrZ0aiOxFxTNDx+xNW7tUS6g2wSClrV6MT3eo
gLVqvocm0RfOgKKeYXG/pbSOuhgvVYsPNKU2DFk5XQH204qH7uqCk5l6wY1qI+4m4AqLi5vNENl7
shf/jf7r0cuyw/+XHZQJN3B14e1P7dBGOtvvdbjGQVKl0KtcrFpRcni5DB9hZOv8kerF3kLnK+6Y
kcXZwe3q2r89fY4WPmz/RaIoAh+FagWoG/jujyAYqZG+/Uf4CDtm0+BrHPiu4guSDF8vHiHSP1Km
cI/gh/aSa4fUWFxfg2QiXm+Hq5jeG+kJ9a5eu7odA53rYqoqK2z6LjIuY2ZxtDdaA9R6FdkBnYId
ZQuRdBWEiD/YjIwaQBwU7QQDvzUc8oyFiVsk0aptc1s4UPfcQgKoK57B+S3r8bu3SGecJLtHkvoG
scXYi/LUB9Dct0Tn359MRrxzs5R/H5FvIjoXj53ZZ83cvv0bJOUcUGqhkFLoVG2uiaayotEVlkEM
zfsQu5yhqj5/a3aFHOCbQqmgAJnQGiUQUs5dzFxAtoUGepIrVxZrriNJCCFUAT7nBqLDo8+04RcK
9yvRG9AUPGmS8ENCQjWetMheyQVl43+sYi/JqpFPs0CLU7KHLPD1QCmkyA8jVT5sE/qsta45ieYx
C/L8w1dBqeklTNXegmhlwdewIGyj2Fdp8RQxkVAg9Cx7TUzmHO+xVEkt+MFRxgO9pawEdWJUUsdx
3HCDa5JX1w6/tqsX1PLVzMg2c5+sSmh7Ptnf8q5m+kPSphhVcMa6XhUA/Iv02wLyQMq2XEzJ5b8s
zezNoZ7PXW8nM+tAsxWCtMRlCnnqKQ6k/PpTB8HpdZAWPXtKl+SWlT2agdjmQ8Cefr8N/YjvpIGm
c9Ydl5+sTaEbTmzUkYPP1GJNXTtclP52q1kZX9RlPEyDdrRqdLx9rBIZ/0q/pYTDUZYC3b8JR6wy
xofMO/fbEZfkwuWsHPiA4kV1F0Hch64c8bTiVNYK8uEhOlNpmSNIX9/97zFt9vHNlryDH5ocFb4F
VuOpHY/xslVPYLcYn/xRJao0/Ft6rDA2qIPLoM7G00w3QwIYhBXBjV643bcNhbE19aVgm5tDtEx/
8onlmaPVYdZBwN+gq3SjlV1MqgKiliAzJOg5VkfQMADuyoPXATqwnsNsIVNEnayTjrBjOO/RFX3g
Cj0WUfssglugiUUxwOaI3px3K9YJKtV3WL0ehTtZrwdTXY1Mrig1VmtT/3zVUk+F/UeK5NkytjMC
gr3y8sWKilFp/s47cJpxi3+ayy+h7blyayjR4gteQMYTogzSzRe7CPqWUrhhJxmpNmv1foNwPaCa
pLC4zw3K/HjgBsGFbqD9jLcp/XKBE07QZ9WMyFvi3py6l+zUrjYHzFrgFriFqIuNIP8rStRboETg
JsMM0Xq9hxMH3Pd8IWhGYGq6vz8bOzhVufDlzqEqc64R/Qluncv0UqVMkmlnbMh7dRkLmvATFvbC
Cz+wRUXHCI/vpz39EK0CJOsCYGscKRJT7U2B66BjwQfgn/0oKVmJr9L5zjwLcmZxC1MPUJyhzdAM
FjX2ir0EL8gze92Hne0mK1NMBuf9lI9Ljn6/tKi3BPH0xsl2YAa3YlDIse8KMXplezNa7SSkUPO9
gtDqJA4LHWHX6kp4dwF1zwi6j5pJgwE8SUMVDioqDCSJ+t2/Sszrua4D4tXtz3BScc5mfNUDQRYI
Gwp0b9M7BJQvaLS01MvPSCxXBDNp2bPDskv8eFP5xpZb8slP8iauGO8Oaq/RNni0I32cIfO9bmSz
fJuwr9VWoLOjY1I2D/uxyJzmm4xhskVsRZCGI35JoWeJlEuSOtRYAvtgERw3G2bXGdFscPB/X55L
FKVCdowYQdKx9KCWXTC7SIOtvU0LWeMYZSvBzD7xC5J/+B3Km5MreqsCUpvCXJL/hdde+QUq4ivQ
oxq0w9hp90IibNxpe0LtjydTBE49DQUOQ1sNrHRqfRJ07yoPC3e/UxWVkacocfkJehrzrI3uEiKm
6zI2HyBWJjaMGB3yqWkMuDgp4EcxDH5of678DkHBYsOfBKtYEFJLTX5KMt1xV/yGXehCGeKnnECE
tFIfywGo8yhzE3TwVsPgUZ0C4ZgF8jydHEmsWgIP73/p6hHx7EWs3YwRZUCZc6nIv4Gxb+bHCfhK
AHK72p/WyTCAeJkywcTZT6IVRjN4QrMT7+vHNhN1BwYf44Ef9DZA5fnwcOoLc51BGn4S8fN3RhoO
mNoc7jiNZqFLHqEJ31gKaHJBiHmrLCuz9ooivJUm31ky24R1TX7YIstiuu6r+AYeS9AFWXxxVYBH
ziGKAx5ZOKcq14cUisaxcJPbO8jPw7UE2hXptDis2g/HO9TUNDKLHNpl4gRuzLgyRNx0RxBgH5Hk
RB/JEViCvG9NPL0lkYlM3jYj2fCy0hMaYF9tXjQ8XM4GJuuyue58K9f2A4nKxajrk2ZFS1/NpYx1
6IZDQrsEbhs2R6DkvOhBL3vgscTp/qoFi4OnmaoX2DoPdENe75UPazQdpdbRvAKBevSHIflFJVrP
eh6sZn8d3cSrxexxaMLm9jBWyr27W5hd3/qATX6sdGB54Mg8dkpXL5upHKRkJn8u80A+2D+hUC0+
CCjBoN7gQyrOVPlGw6tKzkBjZ/9cGg7bd0hnd8wYfqGkVE0D5VckNRKTUlWw5zjO9jm8uNmy96s/
FhTY0z2Lvd3IHE0dpue5DYgvmiNW3XayKSffmG8vjTxN97n0nyS+/7njPJSogLftZLrwXJe7pe60
QkILNrJh8u7TAt4I99rXadzSkfVNVca1vzPTnnpDqq6c/yfrPnIxw75zuIMXrMsyD75qAGtMlxqb
bI3mdDB8XKvFwZlzcGEVHAppeXWv0vI4Ye3ntb5xxNdm4/Yi0M+CrGFWcQ6tQpbPv+fDFwS1mG/s
/SV7EJSbmqIyhdAn8Gz3GUMzzYD4PlygCXbGLiE5etTbLxhd+cOTBdLWzS+LSSddEQ7H43pv+zBd
33xrMHLLInXXeFxXQxgClFSHzqUXYfwquNXJVQ11D/PHF/CBJBJgu+disfP26Tx42KxhIuhEy6w3
7TusRbBSLNqyUZTcygJ0sJoI+LrmzUzBhEX9GXWQdDmZBMfKja0jLIMKnRU2VguK33zDRU6pVxLC
ffdrMzDRYF1o2QRpdIaNnzj9awFuY5qb+GU/hS19253hLoc9H2n0gySMUK0YR6kjy7HOq8/uJxcb
sMd6WiqaDuOURejJehZSBaCMIMZSqZUZucAVgGzvwi/+VfWsgg1GYUyaY6NIy3/5lCSA+zbkPlAC
HzBK4Hxav/jjo+2hgQwnb5IhNmFJF0pLSbkoiv29SQRdwvmeSURAnIxzpjy3+kSkQPMrb6xuqqsx
ctH2o+fJk3M+EvUkjPYd0xWY8ysiTTHLr4k36Nr2W8r4/WPOJgPL2DMAwpVs06UKLRHI5Cv00DHM
twwJ79jkSFI8t3tvZ2k4NJP+1DLVfMHaqXhBHzA1YNzNEpHog6WT8Vjw+3B+GVMTwBiJTIgz3t+Q
LKFccKXkZP1m7+J7cGL58FSItOxgI2pPeSlwUfK0FGO8pW0Lb5xzNos17hx79gQ/GWCiCOYSux+y
KOUktnND7MdOs3dcGL3TwyN6UAIl/8/jmkTDObsLx8B2xqLgfzGujvMtyEOggFAZdgkLzRFEsdug
xuGPfYAGNtcOPlfWEaBCmXLjNSUeeghtn/tbbTnLxWWSiWR5V/m1zAmrQ0rWChWh3XlmVhSqXdPH
AYeXFA4RpD+N6eBgwTEhmDwsJj4pi7CbQCqHRZF+MMhPtzwYH/A5nAkXvG+jIE6pz5fwJ7gLE2Yo
otxc9owNlI+cImmmD+vE5SPHSP2Nihdz95ylHwfdI8T8AtcCjzqYb0Uptk+UvD7JSe18Xvt9yrID
7HcvSKqddb9IaejGsuo9ue8eKZtpy244MTwoxXCwfeHaKmwQQfcY8aW8fztcqrbx8iu5ew3ZUIif
NDtrfztB/OoBACr9hR2+yJRkDSsTjaoULHe7R5zu3JE5NoKQ9iceJtkvp9e4+AM7VSRo1B8YjG3o
f4yZrKaanX6T7+OVw3NFlkaHD5ZH/fVR045mYf9kYgFPy7Gz+EpAygZ/2wopRWAIOoOFe/IF70rv
NwUso0pbfPdgE3m38uneUGsTnhgDq0F1ns3PMK6CcI5rl+Jxw4HqolXiYJAes/SMaxDILzQBHqFM
C8vUMUE0tDotVwV+chf3r1dvo1kygy20MGkdbpV3o2OrKjkTyt9Izgt3sChoT6XOgHyZRs05Av2F
10BJ40XXzd25qWuoxIf39+fY/JmYqZl0pIZGRhth2ppobs1b1G+d8D+tj9OB5ycwALMsPyFEP53k
eBLYqBbekYtwusvCibDd5/tf7+heXLz6YL8AXlqjLCO5xOOhqYrYQyIiFXc0HsgvdTaow7XHrboo
tNAEoZHz4Pd7d74rGLMT44SdA90Dh/Mt/ntEcsVJgyfpxHYxoPi3JP663MKTmsXbYTd2sH219waz
l1kbZX8NpzqaXUaUIYjM2ApVaKRUO9Fsv8rBI9Cav8RACnUYDF176Xcu6KXMlZrEM4JJGmTCDT9K
4o5aU7AIap3SGVsyO7/tkyvYhOqK2iSJBwPu5Zmbwo4mQNa+zsOwbC9o64lMtw4m5DB+kuapHxJN
h4zrx9pPgADcPIKpvVsCyt0YP/KXdMUuvM8J6rbPtpXxnARTp5sdhdkd+iHDNS1w1CrMvbjrQXt1
MadJsRNjhijak4XKzp6OJdH22jfULoJhLQymmLWRRmYewJ8RBHGPP1CUiKkUtnNa1q9IJ5cdakcd
w05vT1ZxGOqkmOlS4gH65dhKIHFWxsk6nRDoIWYqzt9Cm71XUvFGVwi64dYdQjftbkA8E8OkFnQu
VWlrzY3/AaVraapw++cPPGQYtLSsFeIlPWnBWvKumKNSseSWqUCHJm/4urw7+7hrLaWaEk+E/0xv
NbUVawIWIDF0y3LQhfVzHxx9wZebT3U3LRKsBWsof7bxIMZ1gmPTAFIIxm2IlFKys+u6PRe/F6Sv
+a9NjX4JdicEQPwupffBVasEkPR+2Osca054ceuyHuNWxVlNx6S2UqZZAuXYC5Hve4zdqytNXehc
Tz6/wEcv2aAJkLJGjQy37zeTF+Oz3IqxmX9+8dh6IolCUXomJlH4PzFaJ7Ot2xjA5+1lkwrzLQuP
Nod9qaa0CrkJ6HgLf4w4BN3IUy0wQ958Ts0+CE2k2ku8nEn/cGDEnXLwgFPHZdl1E0HazRNeOwDE
8ycP65NeLTPn2+0fZYbgChvZqi5ggEsWPioPBMrbcj3UTbjyINs4gHPUgiad+tGQe2di4xxo+nly
H30+lL7uxSxAZUkgsfQxptKJ/PjmaF9LiizYim29S5dBGQEdXnKjaMCj3Cwm6aK+7HhryNlv2orK
Qpdk1ScpWaLood3Ndz5p8Uf0Y6xHbNT7296LiXsqbnidBZqotTtZ0WiFkW7/rTegBBf5bBXxuRaq
hVGFIqpzUQ455X85o6hbHx4HPsbK3ciyPJOnnc+98BngXBkBIcdQRQMhzD7hwrhtJWF/eIW5vYO9
zlL+QJB/RWuGDCYib2W56bpvD/07LMek4EFJ9XNNlbKAG8rlThGzT1ZMqCrb/dm6D25B2boMil1I
MyhaodS3EVEhZD0kADrO9AuWfda8Mfra8FrPpUW7Lj4t0X6FH66CQtTtCOw0r7LDIalqpIXf1FNT
ohdIFQ5X3BPl+68DPeybICcJUnuzbuC+DwyMbhwuzGZC5GPBgMnYKowAot6qv/0Lrb5S1A6h18Ei
WhZ/ckByF9QoIduCDo+ge8yS8pDqttg05BS9Fx8NOtpunEUtb8P/bxAI0yNLDmf+J7DCwYJdT3UF
fCUWuE3kL5EP5t7GqaTlpS5OgrrJZ2Q5C8j+6eBYcieR6yozQbMIfvSGzEybTW0oF0fdfWmqUEB5
Zl7h7Bh/muZURT29RYOrqeP9GR29NpWH5Yet/WSaFVkXkUNADw7PDtZcXiKDoMbAjgJH1+BKG1gK
pueDYsIr1lLmrZER0uckNUzUcam6jk94soVJp1Xk7ncj5lBNQi1JCYeqs4ceSVGGgLo1F7NdSthp
olNGObaiLOiJRgrwxsE9gLQ0H3gH9+KT6htmwyCpux0J6cK4liVMIM3ri3mL3J2L/Qg3Ko/cmq0K
qK525EuYZnWcozxE6Rw2EbCMmJFhOngFHwut371530ubu0IqjOdtj6ch+mZcGC5wxktfwhxmakU2
VXqCtcNjLgdLlmxr3n7ay6Ye2OB/aKMmS2lats4J36TOtBhv/wHZ+vy4TEZCqdYu49TbcMyFa+aO
mMTiO9KANSsM8Tm3QAeFAjsJBYBGtfWQSEe6jTHJrl+zXIuU85MOM05W1cq119Y31SjUocpByub2
KWZWuThrIE6Mu6gHmc/+ep3XXv5zMDUTmSx55RRZ8GoS2g2cLb4REhw48+h6tEUsKXnDim/zLrT6
MnP29s7S7e19JSpJkHH5OEEPZ76T67LTTbRj6ZVOERwkwiT2BKKNGPY6DhNMhxtpL4CJZx7TXk+W
UaN8RejFG45oLIz+LtRBsDr7950M14FpNIH6ClzNc4JEEP8Csn0AB5P23TFbGCKNA8TDUJAMFLh+
S6qy6UZd23MaZZLujOYW5VfnRPdfyLTXsKlYm8jq+0mrKUDQQgHayX2XrUpIiwxQniemsVn64CIb
aL8lCtCrPiHmVq+Ml3pL1ebUV5SHgWIuHYzIALg5wjiBfEM0//zEZnpmAb6Ps0wfZdkf+eOC8bTD
YLTvUNp92mjPvhrThui1b8o5hbluNuqfBgl3FTze1DUHBTW8sSI0sKk5ufiACvhvfaPLjRgzFe40
7Z2u9Vo49q1N23J49BeMH4Ojoey/Mr8IxVY7cfcOcS0p/PvHruUKYlWStO0kK0y2Kz+gknrKvIPO
1zaJOZa19XukWTHTEV//BVLzGIFqHU73vcYiOD4ebBVz976HwiBIkzmUZma34HEwLFAWtDsMIt++
Q+j023j+gz0aKHRgDg0EINTbHUOB2yAupqe224o9H71s9LQ7t7pCKDDNB0obNRCH2Jstaapz00zj
UKDUwPMEXoov1EEG7iCVldM9ST/AkVYJmVUvt+ibktcu+7e0Iv6GBSf4rjyxaXp0UFmpo8rWjLNO
jPTslcsEy97f/18yPRWB0F/IMo9qLLT56QCL4ns3skIlhcv1jz2Fk4bkf18iaN52vluPQLeNi2xg
nbUzGwZN3z8F3Ssa4UxvgjQyUQ462tLT2zDlQWKkYhcfEYLDZ8DPipgtFoPKEZBjJRcP5qfRbD/Y
Zw+kz3+UkNoMwnHQiIo0mY2dguRoh5ul7pp3xy9SuC89pnN79xPorHSxQ6Nsp/qxNMBRcop8ratT
5qEWzfTDLYBAyRsAV9jmsQ9AEvjOa2t0Pvr7LBvagAzQvvxp+4KejnAMtSVORiK/95Xg0NJ4KK/Q
7UE7X8a8YgjwB4G9SmiUYonOSdlJfxEuhv5VT4ZKftHEqxtazYUKwPC/tq6wdXGad+Dq4k+DsTXm
jhZLzvKN/QhX7k170eTuzBSvasAUPAlIrythhhakiMwOvfCj7IenpmdjzMnpi5WTtHiZ7bF2kLZk
B/YO/UoczB6H8En5kX6Jes99A8dlhBylFjOrskkzyZc+1q7cyCvXDIECprkKD23VEz//cYSdnHA8
Z93exOnaXjSC30rhhUvynEiIQ5gJUNqudk+0E3I15bnc4oAnSPSE1BDOvZu7M5pgzcWlL48+zvzZ
DclrVDB0X/U3uNr9DTx5OwvrjO/h7lK0LtLtSJ9xPcbJx0ElL9ZWdyxn/J1rvs3OJusJtcRt5F6v
g6VuRRFzMnG4fBavwfxMPhSeLylJfiY7Pn3nhYMZPLiiC0DvjqnG7C4HmVwV9D99E7iB+icUIjNz
4oZextJUstDagAAERancGWh/1lvt4y3uDt6gfv5bIus0EjSjcHv8j86LQniHRvmTKNijnKUiKIEI
a3uJjuF4tXlYQmGL7ZEExJoOjo3cFGfgIT7/dirqpn5jy+mc2wVOgbk8oeWKsT0OPINfW9g7lAxL
2PljELDeyx8DsZpAI6hVsbgrrpQsn3qfUGVvAJ9USBcKY2RJwI+1IwDPeNCmWCKHlIMB2AGR7aQO
N3a/IWqSPjkfElxVb84KEon08t8RLL2EvkYjaITqNIVTxLNFVVq9AIVqENgO4mcfPVa4HzMQYZVo
LFCiuy3nTGz80b9hY8WdV9dbCwFOfqXxzH4uZn5IPOi2wCVgO0g3BxCWdfqXasYNhA2bTJaBfX9X
9qJ5zwxa0HXpExGxgCT/2qj0kfH4+U7GPjccZtYXyu/XmxKsiUpdybV246QaLbLb5f47KeTr7izg
oZfnp/ZRvy2KQ3FYDBaDFDgfMgdefE9Z4cE3tPBvnFNkOy6SdeJzXb6krGwf5ICEhLS3ylg39RGc
3Bvyi3CzohCrcw3zQo53EGNiS8ix25fXImjAoP/cmTyvUXGa7r/26pD39EeR5HrTaMSs/DbPgR1p
d4wXAXQsPtVYx+V6G7VYLtZvVkNLk1SGd8hJasvnx6Tf332XRWMIzjK3wl+s/4m7cN7DeGPJ+y7y
iZwQK5fMcuEE32yZVA3ACU8t7RZ6vrcOCTjNCf+TIYIAM/MJjlGT/3GA6naKyDPDqm64urbu2vLA
NyBmUOgDTE3QIq9862Lk+xhfCjqdSSuOWLaJDqfHRLr5zCm67lZPuq99B1msfFGwx+j5ZuZ+0VyR
gUh47f+JUOdwcoKNuTDUws+NBD6/Ml2sc5fnlYTLFw9CzpgUiQxkBY+b3qHkN6HkwaMl0L8+PS8B
OSnlOHTdTR8aINfrN+Jj1fpRGNiodDrbm6zpykUy7PHq1SgGQRN1giDVlMpyMVwiW/sChqtWqBMe
znLQrHwf/n4ncq3Zv1lCSwHCeqw9joVCiqRMB5A3TkaOx0mUbLHuTlqvmMnuLuCU6EX15cxoQTfv
VdNAZTFozDgMzsWuIVgnVkzy3rW6Owko/U3dJZ5gZX4lvj15c/Kfw4grQevH2vJ/siRr5Vrx0cCg
TIiJDshf4BBJxWhyt8kqfOz0sp6lE6Jr5Y9jojNcSNhxI5kyxhJl5XEp3wHfxooyK2RTwuAR+2LN
eEapHxeOx2i09yMs9lCuPvz4hKG8VJ8mPFLEO/CLwjsZ0gvVMKEtVU/RNUgVs+pSvY+VuQmjYcrr
a8BFMQHJHaNBnV790PXsExXME3M0++JhOhD3e5L+KPH4s2wlFlAW0GCADPrCB4ATvF5qAfwEqarA
DVOQbHiuNkeYhAOaDP1qCjOFmGhH9GLNTukDTdJXcVZLTFopUB6mt0PtdOg+A5fII/ZCmI3QTtp7
0a2zc+dm11y2wcBIf9ACslQe2awHqPxKlZdt8qphD1a6KFNfsnkvdTitCpbJi4HKFLQHRZylDsgL
pag9IINaSGjkJB3LaB3IIeghQ6KnuIf2VC4arfn0xEjBd7EywdHQfl4VijwhDisErC7cSJAWNBGG
EOHuoiVKd55CyLFjDNFqreTSl+kEVYo4vAyXzCpMAWvyea2narI16/VfBclCaKqakKK9KDZt4++g
gOeKFwE5YAgNbfBtMb9YDUEEpl8kCEMPQ3DsSUV2ep+VMoNaEt77I6BPzv7SEFea03poW7qe1nMP
E5QmUb2eI733OKx7e6aSEPNOzbTdR6mwAG0WaByDLuVWid5xlaAB0HZjIZ1t4q1umZ7g/wXgH9RF
nD6LNbYVHtnWQYshxoVyzGymupRSaZbPwNkTXtHCxQFEoqe+YnevjsyA0EX2teXof6E/BNFUqj54
LShxgavQy0A1PtuRBm4pSF+R6gbcGOLx3ZcWBaRoLZ2HmU+Zoah9/G1EuLiLpWeKKXbJyEeT3S3M
HaCxZq2TJQZ8f0yn66EWweUsPP83bis8BB3Qs6EHbkoaUEAWqACqWY7f9r7wO9oz0TDKKF0HBiC0
5vNfpJ6zDlD2Uc1s3bzE9Q1/OaVdYEyYFdchqPCyIQgmaJJvBcoif/NOFk7zSRPazVCtIazh44f6
oAHu/os9F6qQPJlR1L4JXZVBYTYzkR9p4aFuSr8DCSB4Bjm3dbTqdFnGBmcaL+ZFGFOZBKwmYM/A
R4FzIoeb73WDzPHzgjeiPY1Gnr7Ndy78Ugfal/pDTZfq72BVpf/uOc+Eh0TrtWB7nCTTNDabf7Hf
0jlyICpf667KVR3eO9yjAc9amlKk+2Wu610bXQqURIMQeYRSIoZgTfLECD0BwiimF6Z/5xGNfUUW
1GioxkGuMMwyXv6KSqwkyoM3Pj6BvLktReZbdPeoT5a6OktUKxqo9kDioVpCunc8ZcqrY0LbqVyu
zQgEWVqdaBchvCeBsreZ9B/7bFYCyGyFUzyV3zCoHSWDcGkMcARYP0Td/g2nwmwh/+1cModVecCD
ocajhOmiqIrI5X7OFQrlMfbnVRWCqCyZ5Igig8JwYMG3JjDQXvyxYV6vrOO2bNl1m/CbCCuHVvtg
dpnvEnkYglvDThHIPyu7+CDJBsvG1yCqQbgj+MrEELL+ol+/nQuHcYkfW6PqIFTz3Wl9P0G01kTo
awXpGs+OkbIVaEVg4p6Dbm4lfWX3KXa3BxbK7Tu0zqPMuFfbypDW+ndIWa8iSIKzh7ZA1qnPKgUa
z6LfWBTcSBEYaoQScE6akMtC3Ir7ZFiom4lMLvCiVP3exs2RCq1W+jdDsGIscIoTKiym60bD2/91
2bCSOb96kq6Pj0c4YSQKD5H9/he82P1sVoTv/rXkOnf6gLRJv+WFi0tr7SO8pjpYk8xXwZu0rqWC
dYBPzczMxa7q7yNdFJRlxiYm+1b8zk07jnGVh86/E+pJHlcz1aH9PW+Yk2cBJeUVH5w8VZcd5slt
NoHnOy75Ol4Vdhp5VNPYDIFWXQX595Z3RndsOMXNV6id02RNJ+GCePE+p6t26qBKjKxnAexv1R00
qYEdoIYx7KXJoouigU0QR3fflV8119u5GC/T+a0c851CR1Cy/4eEYRMkaVpX0ncLlH5/aUUz3Akb
QBZvlU+zYBfcN38Rf2rbxWylPqsmEUqQghHQqFdp6V0VI3/CbYuGZUstGM7vixbtseNjnHBp9M2l
w90JB1IBqoPpkhWnK+d05eDurbCRtLF+GNCIY9hS9B2Ec+JZ8YVj7ckwJXtjaCnzuVRRh9Xl64Rz
8nPBrFFnV1eJLXsonWzB+oEiVSc3BzNtr//QkGfojF7dNvj4cVgMwrY6+lkSGJg6COTorySSKQWZ
QJz6FdB2JBAMKB4vkMiQbM3jZZNp9ETc/aPMVdfJULj3zOQgcILdAiPz+6+aFqaGMUbayF+Afntl
NubfCAY1g2wJ7598bPHr+pM41eJ6V2CWFV0ucwT8by+4kVow8STj/6VdiaB4GN33aThCENjR04eh
gsGhPG2h4W+xAsj15pYb9LKCSpK2BlcxVFIBEZE+lq5pMsn9QgcOb1c1BrDM0HGGDa8QdnU1HLf4
e0fYyOCTDtJRe2B3ZR/QCd+Mnw3Uxdm0VCIIz2m+dT+7oFiOTitx0x0ZBqk8gRgFIExcVC5U1fZa
aLR7NdSYCUaHosYo+W8DB9PkfUlHDxS+6VoDHljr4ULQ0m7o5Ay+HOifsmqZmkowgQS8YAz6xHdm
I2kkXY67cPK6+2U5RdPJAbbyACN6zJP730XeWgkw6tYsBBk4Mg65EAG8Y+EGPZncciOPrsRgQoTO
X8DIzpbD1g1UhJ4DSdQAqwKpuPu/4urf4/skcC2uzT74CBeGIuqF5DW0gWXQxfLIsnaflZiwHhDe
6SuhOCMeRqcmgU8UnL+fvvkyDz1o/uPp81k9zMRj0rzeZwYnSFIkWfpT4N9F05wfX8Usu0t1sHlY
MadUVHgU3eU+3Ady0mUUY482jaPFhTne1RK73ftun4RL6Q1Y3TqGRCpz9B/xLRmZc8j7woufXB2i
smjT5o1jae0DrCLEDMPq6eoj9Lu6+CJHf/4UZyigUY3HpHobQrnzVzT7dAJl+exAravZwkde9igC
bE9XrKTanwTTRblIXcJ7tmGtfG6rwOELZOE4Qoj4MHVYTUjvHdetRvtLgnEKL86N+raOe1pOu4Va
4FjYkw18N98sTMNaccdh6WUyjiCaN+S0odBmv9Y/OO4mbkiHnqAL1W/tsr0ZuiCE8zTht3QMoDeQ
qTJe9SQSTn5E+sUT6EgGHoRVz+pN+W4FZIJtDD+kcC2RtbyhXL6jsyU6whLCGwUJyIljOY9akBTs
EYJNDfquNhi35MLSgDp64faj1868zvIaycZlLvlWCZWYExRVyz5a7rA68viDtukIeXYLwBc/S4oG
Y7u0YB9cXw4t/H1c4JJ7TCeqLXcxJkY+Ko3ah40VPcXW1Fkriy90e5zBqMMwhrJ9DctvdTV8gya5
A5AjutKeVDKNTd6zFj84xc3zdyKwJjSl3/pUijHc/utdqDSwlR7B7B/g8Y6hMMouSISk7EhEQQ/D
N/qyAZ+H56qzEvKXtd5HpIaxCa/0nepCeSE5hRrYYMe2NcPebQ0R2CqR3GdPhVfito9PxG0zK5Cm
tQzPhTcNrOnjn8R/vYHrWdWyeHai/TSYiWhqzyjvm67qqhi/7m5YRlHXGu6IwfMxIBl8NzgDycWu
aQ3+0D5Hmv/kMOc91i6xLQIk63gOla+NKzxQqDkXfinKisgjRjCRrm5Qe+Ccl25XpwhDYBhIKSPl
ovBen4uJuthV0BvKlzsjG3UpAvFJJZEhvckYucXC2SyaQJ6MEI7KXzKCy2fP+kGy+T8xhqwE2dg2
gHAsgJ4cVBLUGsLlCuVywBS3NHFQ3cC0DJHmv07DwTJjP4+vFN+2rEdKEqwldJD6MtUU5nyH1V99
6geA2Lu9wybbJ0QakbHgxE6H9pDFySSaIIAHvixanmXRB/KxncNx4nRvQlxCBcla3+N8DKMoEFnM
sCKQ9S97D7JQ+fmfTUsPgWw853pYTnhy7GTIbeH72MVXNb5UcbtzCe2SeRPo70hhnMbeginEm/pS
gFyFPGxWkPIlG7Ksctnm0sXUOII+iYKjmqPIMRFupQ/uK2dfr9Od+qlOmSbWNu/PxslUfoySjAGb
G3guCauDqPOCQB0Dzl4EEECLj2UFCKdX3k6SHe/yJdUvmVVH+gGVPehA4UF6IVlyBqXXLyAWUpUS
MVdUR+7ZzQQQ8OblUoWS1I3sMww8223q80xBi3PruyCLMvyfX620GwK8cgE5q9ah2GBiGzUrApG0
AB5HHOfsu7ZYRcQfsisyfH4MaP+vpLySKs2KuPBPYnThw012aS0MB2pMJAjeDo7IdIQwfrMcSSAs
xKoGf2rDqZxpomTK72eJTCZg7fOsdJPXCfT+/X1BoTeVA6tGjB1t7vzTj5ISsBL3Nv1x3ha3DHvd
qJ5NThP9QCWG9okcMyaMsrrcARP0YI4AXDpi8V5HQ2t6r4z4WHUOauet00REAwnMetbVlT+eT9x+
54BmnDu5GYb8uY8gfe3EqtJwP9K67D96TYS0St/9vi8dYzZzmdV3BQczM7e9yh9a1IEFPeLn24Nb
9v5VuMoU4yxWabulTRQlBbqmRvyfCuZPSAS++qNiDJr/nZI8zdYB0uoz4e3N0rixm0gvyOD/GYpJ
1X9GGhWFKBH3pBXbQDXYRybuhEomxwHqut+dhd8f/+XSDQ9ZFBKFi3xeLY9yNLuhCfhypFCMQFOJ
vTLGXnoQWpJQbHV6ZZ0WdKZZedLlH44s915ng+aD5OoO5Tn67IWpw+xqhS5Y5TL2Rv7sNkvkeiyu
MbnR+38lN5JKuzL7muhyAsXdBfEaSjpaSlU7BKTv9fiHvtBxd43EnxstXqFk5SNp/aJkGBRQ5Kff
vImRwUDmJlv+mHy4JcM6nmL6NKEPm8FIx4uI6GQp5ROs+D9/5NPOEM5Fon9eLS6ExFAGh4ABPsDv
BL2dWxYxa2sNFcDUkQFt1y3SP74RB8DDTQZh3QA/ojRdWvL6Qdr124gfk6OFFhHLlEBX6fkZaDRp
yYGvPpaZOciOd18pLdA7zZ9gRgiSYEvW9H4VXriZGy+7sQP7hLKdex0cVxnL0l0FmVWIGcd6KO/y
a99rg7ooJQXA02AYRN82a7XwuKmfPsJoN+qpRp2tmM0Nn9MBjaDIQaK0aEhk21ckbMs1e5pjxmuU
rDBuM8Wz17BcXepAHwa84wRfYj5GZSUKYQEpekcLaUxak/LFGBpg4eep5jLYodKX4HTrR+buQMuX
uE600uwnZnYfl8gJyNWZG6iC5vsNvJsbqMyKUAE2UQ+JkvurcdBHN5n79XoVXzWyXmPvYH3QyabM
JMy39ZGm5jFZq8zfXx7cZLUa1dKQb/3q66Zsnkq5NHKbBR8aRaCi8XLFrfCK5NNYtI1zgyf3IHtY
j5mMrpqPkT5zUCBM4jqWuvhmn10X18PVh+DikFQV/wFT+5ZP+tTHUi7ukdlFUIAQFAaULMVcd1Sr
V470VtTRnG9GfASWYjx65y4zK9VtxCX1DGZyuDoMDOwvfkwRSmVvvjaLkRTpMF9k684DpEDiXlxs
De9APAmbwnFPGqE/FOfMp9wU+0chARO+iFMJGkq1HrJi6Ac4pt/zVLTUVCOCRtvb4h0IAweT4Hgt
Nx9f/eEHBbdv7mcICWsNmgyZUH4vf+vjiwLAM5rtiafQc6y6cXneEamhTiBeYRbpn/bUpzTAn/jD
Dhng74ROQBKMrd4LQIp8NFwkL1ajOdQRWD18jPnnflzHdWWvJBZ0a1CAyrxSDtA8UZfrlrbAMl5v
XHKJ+GcTlvBVxFz/sDYOrAFCdWpmGsq2PNeVSx9Z6sjO6v+W2xX/Ch5uwAyw1SqLHhyuxzmqJSWx
EwWlTIQ6uM+KNw8aw8orWb17v1fs2rV8MjgCbDg3s4W4M72NmraDxDUK6ebbmyjBcgP/rVmkvl/z
VXxHptFuB9sDFPfNFJre/qIUia8EVJf+4o5/17psvO5lGvvxiOAjUn5e7EEe7ExbhOMG60Jsid+d
aTR/ToDc9ri4agduMqIdz/v3ub9pUlrTARmTW0kPkekPGczgNVEYHoqArZ9oUfkswn/fvCQGf1mC
8Sr85Dgz5Rlvv820wcX58n44o6jR/8IKsKkLUnVLk5E8Ljx/jrTxydK4qOvJFT0MrBzkDpeJqmVO
qJ5wialTKhjBUKE3ONSCSeT8lvZnntB+F11VyumJe1Kq8GZ9eB8JjCoIyOMy864vrvp3KMwkR/On
aS6FKAve2fFJTcqzcnG5xuUG8d2vRC4S7BWxxZkxdOGZyIN3zxUFopg1ZGyo0NunD7zhZ9vBFtfg
UZLr1jM1x7j7KqblZoO64A6TPyTAZ/UMv4IihxbZRowJ9LlXL9ssjQ1ocK2S4FOb0KaI3Hia+ZI9
HjjIzOzFZlJegfxjW2OF1/29tYBOI4I4MY5icGLHSyRwS+xwvwBlV9e0slg3c6GVSVetTSNrUqDb
36ud4yuLgfTjyTkCZvLYc/xPRroO9wHqV8jwpknqbDBK2Y+d6gaFxtrtEtOGt9MAm4osF/mNVC3O
TDYme7uHBEtBI/KS8fJDmxQjGO/AcivaJUfUbTPwF1yOc+a4Boa8ITM5ltENtrMTPYuKyMfldVcU
dCY5OeV9IQGpW/sMeegDNfWM7KJMtYA04xLagkR004ZqjigJCYGk5Skn2b+d5pDwPrS0lbx1MY+m
0cIDjjPfZEPAA4DJL0+IoJgmZxDkGt/2ILWFrmtj5RP9TWm6gUR+HCa5e/5dMiGL/n53U3eh16W1
uaXRaFam1vxeZvPoyPhk4COTBVMou2PHnPAPP7aISkQKMLkqMht6rqdHUIpMt2z4WShNQwKIORzA
D3xakL10l9XpIDTHK1Xu1TyzJh1AhFn4ifeTOzOh54tE428mZyPvkyrBqg1tcrq/Ii3VmV6fqTgy
gIwWc8OuZ5nMCfteslBxMCe4ivfMZzxqIGkWQ5Zp5m1szfL9tPs9ep9x29Nm+VwroIKO1uBdJ2Sl
ztFDLjJvQsyVsSDAPl9NuAXGz0CBTRmiORQYSZnJOarJ8Uc9EblgwuWAXFbgIoBf4tuJBIOROO6r
gRHaQ1VT1gOlJe6cJlZW/Z6unJt5y7tDh/OxJbfYWTZ17pZG+TtL5aJC0UdFlsd87UPsN8XwW939
2AgnDg46eDu6VbXnC5HYL8XNsh6ITU+eijViGT5Ny9qwHc/ciRlqzUcFrtZjWGBZjjoHoVIhRgJ/
eerTeaBo5bDluvQ/8/jOX14G0VF/Yv5Kj1bs1duP2SBDC2GXHToKAClKJXcKPb19AD910pVGSvhI
cjdq1VU4JCKDRB4mrlfOzKWTF8j6uANVF2FP9VpfuHFnbXcZyifBi2ORlUKUtzMk0MtyWUQ/0Zf2
3TKU/wlFXzcpW1VlMT3W/6PPSO/mAHvEUVp806oqCeFdBGPPnBFjnUYYRXUIPksUE5yb8EFlllrY
YcpBqxMVGkDMqYBTLBjHpfTIINlfExeZuiRhww4IcAGxnQ7SNzFJzU4afTOuwL9vNp8ASiLLzOVZ
37iOLExMyrRpStjymiLqi+qUZ+gM0MboEG7AqL1vsmqX8fRm9dWfv4Hk+3Q+KAttwAefH5VKLApD
bKulW7tyn4vcu6vF5m3of/xXRqdBpOcN1NwybXr4RwXzLQOV1YJKJtfmeMmPzFGZpgkfrWdtkH9Q
fRmJ5gFxpr1Xg3dA/ACdrRng2WZHFWcrbrgNYwF38f7DCCCQeBYHqvy8NdJnbP65z9BnlCkKf4kS
+SOwSaoRGWr1MimsDG2yjBznhRZMGiGeTVobEdf5N9Zru4LeTDtb9RY47yn9qZ6ZwK2gqvgXss8f
k/KQwSeMBkHi+tf+GZ/Iswtc5UjgZbzpspHXzfjnyttJB1ett4+2QVrNZR8OvfdAEz53MYk6FnZW
b280z9m2TsSsaMJcx1J0Y7U4wmlhhIYtJ3VCwyrGR8W5th+xOte4heH2l9vONXv2WI3aiBl7a5p/
p5Bi0JldnkasO8AOvkU5IPgu8gQvy/E/acfWY8EoWWXwkJNE3Blk9IwSRLk6jpF2czBLABE/GR/G
19/EZOFodJ6G+WCvlQ7hxjXmBTNeaEdZt76MwI12II0q7+rRJmKFWw/DlMCTfyKVg/pCQ7Y+959Q
qG0zF/1lUxyT6Os/IK8kC+vsFXPQxR4pPY4F6KbVVdZ7Ha+sUDwKNuWf4cgyk+ys6t5WMiI6wU72
8xXItTevdPPfZk8v4OF8+pGn5vstGNGgzynYUzfUvHUxa5VRUat1VIAa3OzGg+jnOzIdLLy3I6hP
Wo/z2jFAq1C2ofhf9/tzAQ7u8JHCwNvwoxOFZSxrJ2Osr7xyIrhVV0/3a9YCgo5+34iGXfzxKlBK
50RSXaAQTHH8siz6Jgo7v6exyOrty4ieilCjoJ8JMHyjuEjbODV5E+be53WiA2GFU+2+21aeF8p/
LQhwbOjB19aUJ+rny1nzoCeDL7/ScZZWFHK8M70S6H/Z4Kw8RLeWzO9ON7qBwKy67eGOvLqAwyvE
tr2XeIoFya982ljWJ9yivDRAKXjqDa2VAxFN8/RyUMzgvidwERDa2e4SQHx/FxS3pXtdr2IjPz8P
tlHjEXbfKnYk9tdWXxDBC39G8893w4A9KFIvc3Rxw30nrvP/o052RJ9LWQY4kZdqzW9RDG5BrJNp
vhiHMu/bqzqzYJthy07J/SlFU/OL6+p/tBollcwgyuyEO7AnLyvuX0of+cxGWEezfXoGtKU5eHkK
UWz5iqCggBJgQuU2VkOUii2MzQdPs8HF2dSac0zXFWMpZSOGLJ8jdmhokVf0MEdpE8rb2Zad61OF
CsAHp0iTzq9McxsdJvlHXmRD+ezyeV3wdpwchUoVCqlSOK/iqj7HYv5w3b/EhJfpY4BW5gsrWwpp
VNwoln0Hp8LQrvXiWh5d8aQK84uapCtA4J2UCZZf1ELcICB4sBucnAsa85nV5q0vqnbcAnwdbN3I
CkQvGTnGaeN+N9hwH5WKEmB1/ljgMRNS0uxezbUh5pRhON3YnFuAagbnBlH1YEbZzym0ljdtShct
OWhkle7uzWZax8OTPfeMjKSM9JBpOu7aVXlfKJxS/YJYqwm9ZaIIgGChdxO+SW5hfTijP08Yy5R/
rPXVSfjNIuHpmPksBAUfkplV7MjfHcEB0HiuKUod6dpP901QWbfkgauScO7aQi9O3CJNsStagWW9
egPMYxHXNaPHWnU8al5VmWppAAuzIF87l9KgouUdGfgrqT5bBrlZyLtsG0LyuY+wdQklp+MhrfX+
0akP1AjSBoocR1w6/uZ1VhJBUvHUj8WUZrhYRiA4CRZXqADhMGdkZpNhejjkUjdvd7+rIdNshjGp
FChQkBgcvlBw/OTVjD1QQM2MjUtYcfKCUrSyZy2vdOb1aXpXFQT893QccXbTvuI9HO30UWstaM5Y
5rVnwkf66N38sZoWeXuDjK/oSmYvdc3aD8lbg4rkWLYoenOF0XcOru4A7XPgyqAzyydE0h5TmOpQ
T8gOvQP8sBntKhY8JY+ch8gI9f4wrGS3emjC9n2ICyyp+LngGdBXe+bjseOXnUE5ERePPQGYjnX9
JBYUv40kXOdggIewyhVhw3FKr/IVnTlN9KoVQTFaLyd8SWX3WEoy5Cyd71kfO5fy8KMnikHY+axd
27gcycqhG13gbo5KJvACfP+A+Kksl/geHBfSDcHK4k8yA3aYE+quuYDgaJJPPl6Mzs+Z1wjZ9RaU
btimKs3/5gImLa80ueyY/lU9w5Kuonoqoyg+OCxufDOmOK5bCU2oy3yH2TIfq/Ien7N3aCuycK/A
XFIS0CNBcIiQRBmsb/5hePvz+sGIE5FkK+uG7pTkt+gN8Hb7UWJHa8q+H57OJa5iw0JdFfojRncr
D0Dd02drLh0YKx4iepr+29OhY0iuIDHCXoWduFqYwV56EJocpGIMtRbnHqWFKraw/JmMHujZTJPU
oZIOLZ3RxNURiJPxvxVWA0KlTBFyMltcNsbNCnC/FWZCsw65ek4UEtgluALuuj1hCAVAOaMUF86y
385SWa124T1ed2FVk760tVoRP8QiyQvLhATJQx3IziG7QECdEUi070C/zG3Qhv6Bt4VBBZvS5wcE
LjiZtgij74zy6UIFvvcwYEagdTRn8U1A1o5ZG8NdrdKYtPAEtsox/Q5io3/1Y/DcPPsZgLCGCV4B
eEOWbLxg2gD+f/fMQ+uJEdYJDagfHHQLjjoM8oxk0UhTF57I4HXxrElEDjpt4t4Ja8XuAiPyjdmu
xKsGoM7kbi0kinkfkwKGbjYp83OxRBCJ56UrCrNKqEzX00SL0w/lbnUrgsFxhLVzUrGeYXcJ5ZSf
CKS7MQvtPqwXQ814gAM4Ja79u9vBroNnb6rDjn46DHmGdvt/dt3RMQuVQvdbiTXJhCtACtUztK8X
cCpmQsUCmzpauC4qNQg8ldNW6SnpGOZFMG+P+8cJjfjuVvPnW6mzdL8mxpQJ7G2RIpT7GuGZGGvy
5CvplMoVzLQWBaHnEKTcAGLI6DMdh5MP+Bspb937sSR5Jb/xb73TEvT7CZjO/YwiAeNEcVl5UCWv
WeqolnDL66pDprDONH195PkWnS7xdm094rNvqjWa+XuZkduzPyHw3FFEMVPzHwuMqzD+9UkUltaX
ysHDrfrJdRAaEdp9LhPBPE910g5zp2C58zA+AEmR3o4NXHE7Qwh5KFnGhnF4AB0DBcGpAAlAjFQt
7i7pal5DshgXNzcveXqO5r7azRLPxdYVsAuejS2y6DHyAPRG6dG0PFOab7kruus/yWTBO0gFs44T
irURGrTtf8y1KoBCqVqAQxdYo7eGuMNXgz9XwvUXTCryIchwb4p6Iu/KqPsDb/lUUSEpgj05qKMQ
kWMBWgCM7qg6BvwDlPTmQ/WDi7P4ajBlIVfd1L2/bYCflZt7HMd6SauAJ9juLWnnMaTK3pnt00TT
6EDpamUaWm6jbM3hHTciOONrHuQdpSfJsyZIJzwdUMIIai++2H/scFgkz47kqsEZqdgUH2LmnQ7E
/LMaG8yLC/TpNaWDV/irrIYpkHyYDxf4/4jRKTmgdObkk7wxjl3xjPzntJGTtvovLtacYcLGhOLX
EnAuYEF20K2KyKFfvWJ3k2mHJnq5lb0NC8QJnt3puMVny+L6HQyHH+YygoYNZrlcJ5lac9M7yR8H
XamHiaLoJzabD/sD8h7T1neHgS3qsqHHMKnMEhCsDp9zA2dDPFMiXI0QDtM7QK1cFjqk9yFVvsOb
qzuYKiHj64S/Z26kU3g35qxtEY3Hg3RNw7WACXi5EXz3PcaOvE9lFSyYMRejH9H5XrHCAvzojBur
hA/tsFp8cVe73c8C7UZI5LjRFDKgWznKIS+08sdTw492XkxmghcHwjZIalDuGE/Tb88yAtKMVv7B
IIdL3JCajZco+PzVVIV9WE1+J74O/vzVVPe29vWQOIoEdtVFqrx1x6rpY+D7NjdmbbjSKm/GmM2w
A+SB3NGlmGATfiHKFE1cj5sVpaBtpBxg+rFQGCn/1YdhltSGxpHcj1ifNAqR7IqBj4oMfyRDsT35
wA0CXAHPJRIzuu2ISPCyRCxtfwnpt/cNchBuxVQGeJbABy4z7hLgkHMRL9cWheC8yAW+jrBafnZ0
TM3WzPoCpqKDT1nq7qSE/SqeB8uS0zZgHEg9YyZFJlL9i2zrHvIsuegrZJehqa9w1gaGWGxbaF4K
o2wsW9UhWz3NA3Y2EstqOZFPxWu0SsYdOY6wC9jhTtsZgL5uBInu7CRGV/clrYrbNfFsMKtOYQFw
TNFswnH4tCcTxuMZRWD8uvlasAmjV+2aqmh9G+k9ZoFdCgXFCgP/olBu/TwfK3YQGVWe448nEAt0
jxkkeym3uOMHlVxO51qwPj/v7ROi0fk2LiveOpsCNc6Fu8yvJCzrApeWksPh1Ny5HcrHyEyaSvZT
HZWmEsKWBnhDBLoz6jUcPOsfEeeHFb5jhj7k1NtdTIWo1ocXj9vTU6wOTv3fVITdLp8fLf2xg0dV
gzMNPUAZPTBx690A1it66+r2VNoqKM18jyPjTcT/gxTrG7672xTtVfm8zrdnEhNu7Dbrs+Fz7VQx
xDwph67tL2cX2BI5vsgoaGnLMcrkhNlkWuFD3DnMpuiENH/L930DFxi8ESShNzRxE4gSfFfqsLF5
K+ik9NMG0LtX3NUe9JN2OQbrKHP8ueTbTJWHxMDb5DNaoDw2jvDI8dIsgkCOcORmWLOdFeDjYlDY
Ouox1vmsL14V7VcNMcXIcj3oUAS8C0lAjUVy1p7/afh1Kjex31NjO3vfsnukOjXbSALSTiRRPnOm
cqzFOBIwiQkN2OzSvu754/61IZE0+Sw7EF2cWCN2QKVIDUmHyRu9oHspb4WRpHixnfgd3/TakdXZ
kjoF+IYUmCmQeEcA1mWhiy+rnhomYR54CtcdjG/iG6kjsm+Zuwfek37uOWQCME2RximCleFhykOH
DZsstcuYGcOA9EkJKdnKk7M2cKCWEpNFwTa/kKU6PyVilK0rUSeKZ0pYC1TX21AFvBvPLXnkuYDC
M3E/Xc0J4vewgQhK13i4pry1dFcvv9FdMpx7i+GVXGa4WfCvK5BKEl1egh8Cf74QMCWNJZGDAf00
E5DoIkvCIRI+IFzNv5tyQ12tuyec8im5mdBzWmE6lps0RW9Zw2WmAWnSkXotu3ALTAc9TBRAVWM5
+u38soZMwKpUbevissEwXQNyUGMZ0I17117rLjvSgL+/hB3FV8iffJymemXWBgnSTFG99T9sBaPo
jYm3fR0YDdLkW0NGkHaxh7/l/O8+pTmNRcQw6cFa61vck/ThTETeqD8jm1+QKLnplj3hd7ijfVzq
4+v8QLIAZYatOjkaBk5wH4qPkuxGBboKBNpXM0WruGo44C934zpGCpXuA+emuJufMaNRgUNQgBAI
1P/aiXDTyOaHV0igZxPbiEIpU9kdGVORhUGGW/77Hk/sC7drW01VS6htOc8PvZU6zrUEw+bvInIK
NFtCLV7fa5n7E2Lk3ZTxwZd5b1DDLexhyEO22LGgEa+QZnGDFHdji8rO0nE03BFnBQIOmfFb1jq6
wgqVwZMhyuTUWab0ps94T5DTKg22tcaoEYet77lsLbFmrlYn1ck+0aBelSxF91CLr6wKI4lGZCKf
PyS05v9XyID3y6lyL61fYcpG6Ju+ZRYVAcDxZlgOuqvSjgoiIB4Q0Gf32wLSCPeHvAuBaAIlfket
PFRs2OrhDYkqq93HVM+Hwtmdq4434CwzQnYL46m3Hwpc7sPOoLMg4adVpli/CIUcMMCDjoFO4LwS
Kx/wMXuavQ3GAf+0hj91f9uxa5v+i07BzdgBYhce35zhfGYo1ufyEHXQuFSG1D0dyy4AVH+mfmK5
NQZF4f9jV9b+VSahIf9JzaWn83+U2CE5nHPfiGfYqxC2i7vggmK13bq3iUuo98yOC8eUcf+NZUED
minQnlUa8pZ+0Ha7WLH645uNuV69cqNX8aijW5bIgnx2Xk0/0BQwTGmqB863X+biLYHc88T6Iz+0
BKbgUtNSHwJBlHq4SZkXMB0QFGdNm5j6eXklgUAsc+ZA+LvuPltVzQEiElVbnl+2pIcZn7js4+mz
/38+1kZpNETg2qnNwSrIUXY/9OAKfNTtQyHu25egTX6feDFcR61LYKYsUKGCTmSkjWZcNbUUL19v
uNhAFWkUtXzSWbz7tZI/OPD+qx39cCNIMklicv+AVW6l+DWEKxgbREhaW+BNWCj/r/yvBqeB6Rbi
qTFBD+CxhyC1K08UpQ1RtfjFnMHthcgqjV1HZapyrUm7cyfJRjxbU+2Bb1QjRjM8SK5njR0lCjEE
021dLNcYX/kPfG5vm0c2+T49WkOKX+aU6d9yDpX4d5cocmseAy+7e4ygliGfPInAIPBf6I/2RbpL
iy//OcxNw53fooKzrRsdSRmAh9mSaFlQk09fBmPBQi0AVwt4qbUgG3A6q1Epz+cP6Iu/xMakPuQ2
9khfq2TjgoXCzmqqLuVCGTH50s0dqhD4fQ4TOSnxZs+ZIMy2XcV44J5eQily8+TlNk/BU77cx1Lz
CmsE/RGWwubX4zMIet/e9IXs15u+Yw3n+VH35MRY5I54DAIva0iN7TpHrSg1wA+r7m0Hwm7+mts2
LdP8ejLsmdhYn7dY5j8BzSFPFinL68G2jHy2ZBT2uCEBneJHEg22/yui74Bkgv2HCEi++WOHlkv3
VPZ3zk4VXmir0GnyIZxlcj/an5ipXtMpwI4g/riDEY9eKBa9GUWhaQzwdE8GCHX1z0566i5UaJ6N
Wk0VpQZkneb4Msm7KdzYdAW+9ffYO7cG/YhAkD2vqLSmoS5rbJrSTeJOHzBJbjnD6TcFeRnQFmUa
ihgtpfzyFrkwJv/7X+SeM5rA/ESTJyt003PH7yeVMUCNOmJzxV9BQSCeq/zmBUQS4X0nKP1M+6xJ
WbTqO4zvNmi96I6JT9DAV8ZgahwesGKAHueuEHQSPEz8d5l+hWzHSmdbWMKP2Y9fZzZ2kriIYoLc
EJTtU/Db5g7AooTPC4TnaS4dMD2cetKt/Ojno8V3Mc7X57rrUQSsbNMz3OhwY5bVy2JpftgcVcSR
feGOsWOWY/7su0cjdYaZ1LaHLrACHAgtCJQa7ew/iNsXyrEmfNLILvul1K3dabPy30VlacisHwne
ua/SME197BUiN9+mf4WGWQE27+8LSqf7zTxpbLhfIBmtSmHlrGl88Kb/JVkXcwjxOXmzYS65X3AZ
bCBmZzQeDjQBg+qx+IxSo2DCCQ2Z2yLInUPEVjEKcoedd64kobhG9OoCEjaUbjw22edV5WAkyR5a
+qPq0VaKQwiC+TaPcTYTS2tqZ7tCnhCcJAz6LWLUyELNYsquqZv7EdeXxKFxOOGcYlPujnv4dJcq
zhM0Z/ffYKAx+sMbc0ZEJnD1t7VuBqzuV7XGVdDQtKekWdV55C4t6PxFEF+2IJzIcG1J3cF0fErB
q27KKlmEaoJPLcjd3W2x0JfY/wZa7VQC0kgKJ9IQf0Fcvm3ZqK2kjjogaS1aJOxNUHGdjQ4F3rgS
+uUWEaGj6sL9Xx0p6Rb4Fklc2+a7WciEmZtHv0KI44n267x9NqQLW+EtnrfM+eS6Yfse65gPwMiH
+xzI/2z9i23cHWD5D/IebxZ5X7EQt1TaEIinxp1EV33yrXHxbTkEscDGZRdpCmsfLeX5GLdGNFZH
tcjGUGWFHO/vCvA5whyChiZlH0Y/aLoiAn3eXj8BRxkAdxLIEK8Z2DmpoRj7uqaoKkq6j/ErlTwN
64fYZzwJcdBVs4jQ9B6Hg44FVPi3/UwquTI1JTjX1PShxGqCkxuIPk9z4Fa8r98WY1SU8YDa2q14
rr4Rvde00fN/9BkzL1jcV/+tPo2FiBh+qaHNVxFiOP3CnfWU3IRPMgqrcAU3ZqPtCI3aAaMGdxIt
RbOoIdSjosEViyiQ/Ft+tGvLGzmaXiAQjVRXLtVgZLK29gPDGZHQpQyvUN+vAfGPvwr+sczmdxwA
QNMCfa7Syabfyq1h3BtzlQzzTWPASFHRia33104n10gDB8UCha65f/ipcr1vW5ie4Zo4lAoEWg0A
NbQGv4iKkf/CB6O2iezcJ7Gyv+7GGWpoSCaDTrtJktexgnVXgItfuPuTD2aYqSvWjPwfeHRul1td
IWATwTATxeNRMyZLMkfvX6exzedPqzN3GNAL28X7bp75RK3EGVqdQgXDWQS95pNVqc4WJ7E2fU6L
vyrz0sxlGK/HUDO67XlQrFzC7nG2TF7Gloyw/Cacxfjl3bNrNgRm16xZu4HsHHZIXgP3+I8ub8js
KIhmvl674EXlqr3qkx0JRwHwg4ttDC+424qEK1bJ33Epsq3bOsK3gy8HzJwJCyOrHlZntyjFBsEO
LXxqQvnEsrM5+DzQQSJZXXN5zN+6ikUQd6v01Wm7t6HJKLm4Y12S3WJhV3i9RHGGloyGhgZ5YXK2
y2ETJFZK/OkIrEYzah7+br4ki06Q3a8j3Agb/tYt+P1Bc9cvWRNUErLQFuvQ6x3818eNAnYKPWWg
MEbFlh7e3OOe95F6oIbrpM9aeN7UT7WSgTPRru0Xx7BY6PVJngEQqn05I+kRob3JgQ9SMXzMh/Fq
5mGJz6supocQcaiMcZH1qsUDC5gt/2eO7yBBZ9YHA9EcBv/lbULfdIo9D3mgQgdcZZiv2cIJ3amZ
kVukwlHX6MUDCAAYzCul6+X1wdcnQGbIyb3gBvpmb46P/1zOyvE5eoK5X0aJytFUn0PGXtPYvP+W
6MZRWO03Ia/lfO/pTRhBD9Vt/GM9dhNa3Hzin2RQc/A3YZlsT/9eCDpUb4J2MnPqKJf1wKN8vWKq
G7tJHsKLkpDtt/E9JL4yTY8lCDlyzPynPNCYdOWjLD0IBYFZ6WBdffcrN76QZplmb1pCX7ty4vtJ
lq3GetMUP2LGKckPtHZQN83AxtWSAJHGhZBbNiJLrRC9+nZiqPWzqBYhozoK/YTbvwuj+uzL3STU
jU2KjA6/3GJCAVKshrKPzVtEPYihtOA+H9LOUNHDShiyxC2sxnMmOI63p/jT9REjKpflj+1l8r0g
epacF21ijy4JMXgXal8u6hdRWEnoRTMkjMxl6DFlR36rxloYUo7Zr53SwmX1SAbLh8ZpcEsqmHkJ
KLJsaOKwe09165e2oYsIb3tHPf+4ETXIFD8DlCyQU0meaU1MIeUv9cYdFVqDkFr3jEA6ezZ3lU0x
7EmzYbNoBeQkfBRk7XWAugzrDb0lEK/bV2jRzF5TfnGtnNxRaL/HC8Js08COZ3M78H8lclYwR9O/
afzdjQaNpVoyCHGvPuANJVW9hFt6ECeM6vKATyaro3y2GB/5jrppPDMjtlFxM0BD4fpuOXjJBas/
P8WX/rnIof/yAEU7CSjAAz1Re5daCQ3fFPnaeJxFqr+4Gfilmo34CxnkrPdCC/WnT7Q1XY9XHVhE
2KMXfyi+kL+Ip5rLw1ZqzdN/WW+wKwLGSfu5nclkUyA3tKEmiCi+QJdmp7hHtM480SWd7yFECKiN
7Mk3UqOJ3+GvhUK5zplaVT9e5aiSsN79J9iRy6bvBoVbQSsYyP7wCBJQtKOPZY/S1bcOAdpLdNCo
qs3T73+0bKmIQQBk2go2bNBUH6sTL4lL4teUrT5qQ9HxlZmSulUc3hwdG3GtLjnnQaupfnuRS3Sm
ELgYb8eaGMUcv/kns6w2mz2PA4DElsjnYTjhtTxd/1N4tMn0lY7y1Di0MjMBRBuPtwYoT5Z5FXTe
FCZ0FWCH4aEKHf741tNUdbyuCXz3GE2DY799vHOTse7UuFURHJ0Tu5tKB3A/1zUTuD2yPt/bxJS3
WS/eWqyexvyEExlcjsotrBnnOcxw3I7G68wMxXHLe6YoJfBR6SUQ2YuJ0pcYaG6/6/5TNwYnEjAC
mfz0s0vrYMqw61Y5MkkXkLhi+Fz1NoCB0d2usaXLNq3RaenHeHFfGiq3Y++bg0nwP6187dgfewCp
iKcwMzsSJxF4ul/zoclxBJkkrJQrTKtMrk5Rr7UYPHMxPAm6RA2U5eU+wgMh++vJ5PwFNHAWX2oh
boGC5W8Mk7i40HFDrM1eVhxusjWNxySh0PxoFmB1vqbTcHHP/AppCaAxq26oOPRtMg+upwcwYXSl
hfuXHLEod0HarRjY6XSeCYaYhJKW5B5b4oDnLORzJkL5fXVQb7gG8dxukiHetPcdh47kQnjrxGDc
wCjr6OAAxC98swJ9q5wtaifjJ3k/kH6rk6pBdcUY56mvytl4KC078dYeNfKS0cnA+7u33TPf4Qpx
vsXkSLFT8/fvEt7eZHEU27MiVYLOO6na4YTLGAeq+yNI1dzO0wqF9hI4vSGz3gvzb/SiEUc+7EII
Uhyd44wm67GtunTq1ch480cjCDLImPOS+yR5pMRMu0+cujkPLJIhaGw6atavPOfgeVaGBjJDp8XP
0ZbVBNiimGTYIbkck723IyNiQ3B/qXyMW/XZJYe9VBn1w6COZvav3tEvZHrl5qM25SFMiM4icWAf
tck7gbkWq4EV9dvOU/GzbbMOs6rdOh5GGFwsFvRNOIqbCQElJysuDhIQSZ+BDB6JV5cE7jIv7Plt
CN9jRBqhw/rTsFXXx7cWrlzeme25zLdaJzDvTCDlKdS2k/OUlSD2kt7HYwAIDFpYxCRrEzt/un2C
JGn39ddVNcYBURjmNpAjKt+2lNqRri8Ug+Jp0q+bz5ffWWg2vt1FuPGAxsoQTXVVFO/VGDCAuySX
SxKg9KF0rnWHOUfzESgUM1mlrv15k9DFyKrorIcYfu1IDnI/bSi1KctbiJUxV9ZGkjG61kg/038T
n9/tyWUQLtVUEcFxk+b+yC3KHjzXSGMaobLX26ioUxJ5icMU9cASst9375RHNi9m5ZHcQmjgZHTQ
fYhwrE9onbxu48Yl0FXG3g90ntZ2wP/ITJcNXrLhYOV5XBNenGXYgNBhevctFxOnP7o4+OtCnLhX
IN4tJx1rJVHLrxMrRCPyrDR7Qr/wlgyAqC8C8sjxP6bne6gLsMjjBqUaUFvoK6VcrkApmUB5bf9u
gHqJSXWgg8dgO6dmXLZRWtsAp1y+bVXZpVF2lt19gTywG1eZhxzcV83U9gy2ik6ze7p0jSUoqPg+
PKvj3NbVrYef+3KrKjtbW16pywBgMxB2plqdmN3IZ2OSmAn419eQ/zjxoulcmj3XWBXGE1ZSsnax
qzY5EIvVBMnhwFYQwBSN4M9kPaVGM+NRtKzIEYVHQKQ8AX5GaJ+Vizp8A4Nkr0U71hBpzQM4eYsJ
5I2mOuiTlUnuXglZ4Zxb5aj+M9g6ldsXWNVd7oBEZTLeEdOtIU+J8zOvPA4oy13iVP3CCRFaw+sm
Sy849oc6ePM3TXB50yPPhy+w/NQpSg0yEvMSjRw15oVAXBXq/Vh7OV2SroXaA4zSgwcd0wGxQWA1
nczEHF8d21xFcDcCOD5feLlOzgaeP3cHQKYvVrVfj2spjYd5AVHfe/RqCK1Ko/78DLYvsVhtfI3w
RjniZ5uxK5tNDq4Oh/TjmdqKQoSfs/tcqWDd7S/R8XWP6kMNc/UkJGdWEvm5x4MzGj/JUiKzS842
uQNsmEZWVAyLaVeNt5hQ7nr/A7dn2alma2PnIM7VgseZSasng8E/jxnmH9YARsbG+kAaapLSKicy
jZz4lqz/ESdhTJmP5VFLJNgEDPxFNMWf41gLT8pY/yCzfQZI0kcc5nH7McoLYdZVm91kz0HFMNRj
t9yeCup/a/1HhHskrKnwgvA7NyofuTPqBi/+//7p2eSCzqGjmCxgP0snfxTKUPPX8vJk1t5LBDUu
x3uZ7fwFhdPEpWkPNTQPuMFFsQx3bJn/So+D+CnTQwHHf3t6qKQQo/rzhFEWqhKB+xB9xefnG2th
23i7Diir62ICB/MypEPSlNB3qgta82SJzC5ZifU11kGx5uSMtxfkWMab+zAfpHvqmLGlfoMZQeYT
t+EqbSAdps0PkxXk5dUxk0zYK9CV0/31OzmJhO26CTQJvTGsWZzFmcSRrfWBaoQOAyXEynshYdxD
QoymLSOtG7W8FNBaAITDez+zXGxmEYodUcGJRSYpPUCDrt4mWXHEjGOF+0cRMmn9bnCfgb3YwIlg
7zMaKIe40T1tjpdzyx+JIdoHK7IRqyMdv3DNPjS0NZIX/Yn3ievaOFAAH0vTzEg0QULxvQLvDdgS
ejTYyPvqDcfoNZE6koOeMQVjwjwtDoEwV2RJrnT3S1iSVdrAnLai4qA8CMtOZif2OxR1wYBndrGE
/df6tMeAubuaJlPM5i6gbjy4cVi5C+/kguVrdPUtG2V3kOgxmehwnoazxcQlYaglDAljY3CwVFWt
n1nXqMQsPDfjKG53qf0MCnUL7CUBfzrUgfG/wYaglYY1m4NTAwOJw/wWCwM+0MzgZXhjpCwWZTny
W7fwVUY1b5uKvXRZMSRlqIh1lZPSQn3FRppJkyNojGDK1iOUYAMC4yllXLsPDM4tISUravvZDESi
LD50luPEgJt+zsMfXXb5dLHGA1jvflzJ3WyJsRBfIMPL4NkfWLH7c2hosm7cRYse1Eekvl/FBKHY
Wle6TX+OVc6EcNjwK8fr0kLRq5Uh21Bt0T+Ze04kQQUDmUUuQymVqs6Ch4x98rUlJfOZvqtDitIs
Atj67RILHnXI5K48J9WfryJ3b2n+BNQrNPMk+uqgJw2OG8v/n9mdWyEp0ot2JGY/CMmBHfX7fxZ6
HafkmeurfIigjWNWI1Jm7P3X0BMwOvVA/Etx9ACz/dK59iOnvIcvK3YfnFcaTr9d94mMKCC0Ab4H
b2QeQTHc+62IWtWcfnPhgHLcCi3yuR1Ol3DlnT4+Xw49MzRstPoagYHQwjJ5RIJZJTtHkjI6wrOM
7YSt0sXrQ/rot3VuXYVZFYq5AHsgfZOx+u1YWD9lxJHxKIRnGZSH6/d87j1jixXAiFMGczqOk2gt
pe7q6wy5cTg5g1bmJF94Zp8g0lYRr4UkHyfSYqbJuR8mRnny2ECuNfvqvOLIo+f3j9BV2uFJIft+
qcB+kTlOzZiduR3JNTwPzEie2u92+dtODiv1iuHnxQr2h6psLk593JkcqUkYjcJKvT39o1iMORot
xqsWsrc/cVklfOvMm/1s9P1mPIbMXyL8NfI5PRFWxCiDI5KwEshXQVHvyLdVAGzjGtSuINDWTyom
t6UXdmkGf9akeBXK4xvRmnioiuCiiJmbv0/mhPl7zSmU/NQozInZM+7oWAXIM8Ibcau3fOT6yEGZ
G+1MdZQ8+lgEVbEW7RKqn8B/osCDjE5gLPz3IpqFhtg/BHawzfJJk26LhsGcFPrGCHziWvQgGIf5
NxV9vpTA7MrqCL3vM6T9nHuGXnxFz5ZSTz2sZkUWT0hjOwEU68bJBuI36AtkuFsn8Er7ynn81ACF
B/5C5YyNGd8lv09GDM58yLfjIZRQrDQXPwbj9iWd4wO8gDYuk38X4vuJxQjRu9rIG0wQ/Hxr5B9x
AKJrLoQl19yUJ0ji+jPaRApW6/YeLa6hLJWXrBS+lsqfLx1vHcp1btfbRGyopNYa5iG9CNDLLLY7
IXoOyidA1HzSUH3+2rNgkqmTQI+ss0ULKlNRxBuEpqeR1K7iQzEuODzRslVyw0GiLFdvr0ob6m9r
DsU+GQ58plbivCKCqDo54ux0t7VOs9WhGARSgxfuOUZWESgKSB3wlSKW3cIWSyfM13TOlcAcmwCD
5Gq45ePcee6BUd/YpSaMvggZ1nBZStYe7DiQhPJVRuk/igq2y8zIGysRfW5A0ivwHHUYrsYyhdU4
mQgisr5lWpHYyP8zCQQ479H+bdbEssAaaGfKyGMssLHXUCZtmwFIASyvYphqSO3XFImpLs8xfXD0
PnhGqoxUaQKFLZ7EH8Zo09oP4Vq4vVFGWF2903uTl5xoKD577ulHTfFIC53bWxClSnEyf8CSNAmd
AFsi/h/P48heDDnF0yWGsaddFj3HlPKKDuln5nn4tx5RetApyUfF4fdzf8jOmztgtVawVQkQ+ViP
hPd/Q0z3+X/LqOIexM8BIc99mQ6rO1KYx05nT0J3NSlehHWb/++aWD4O7zB5sEflk7P3xMAl8SvZ
tnBuVICEipCtsE+j1fNmgxIhOjBLkFTiehs/F0kBtfMRPtWBFQRsdhr6TvwKtTcUDV/AXz7vUZ0T
IXVc2IpWIjMbwv73uEkubOfCemYpVx0+YkyqisXLK+SMqoJc79C1uCAf3EnoCpvyaa6/w6CRUsKQ
kPJlw3Qjf+e0J0pigx4t4OMd6BDFUL6g4rdfQWr3IG4uPz1hDZ2q7ZiF4lO4SsZsXIvbxAHnL7c5
ZTB8Z6gDu1ArIflW/v8z4i9rn5bDEe3BrlQYZQx2atn0Ylm260vFbDpjHyMEE89XYLqD+vNqnu+b
9Soqq48Y38GNce+ceSq9K+0ic86XbQUrC+1xkcXr0VipGflozr5KTWD+OuuLig+F+urLGo1urWjM
io2qZMaLWlRcMi5zkP5Jz5N8qorvobVjklV/Ej2NpjZ0+hDrf9/cW7PPZloz4EfFK8xiVkKvDKhD
QpBuKq8n7rcVll4rL7BINyDgZJPPIbM4NPfd/IvM6WGIChRg2PjmBmh+k3w0FY7Bd/CmYRWzsTT5
UFQJWVonqRcHNKW6RGUxu5fPKr+q4EeXnHPEgKap0JKkWV9jbr9lS97KjPq34ivO0DZEsNoWl2YY
c//jEKdi+BCpRSxInBv5IuzmbVWVdZUwIRy5PeDX0fhYKjmYNGIXrZCAbTmheLFMHDcbsWEuti4C
vU6fjmt2rPJcfNbTAHgjtZZhBJSSrP6O2Tbhd5moC8Qm5OrgT/lAlfJz4xPhw5hopEpgxzirlJVf
LK5dMo07srk34JKm1Yy1AiUdCp9elFdXtK46vlWr9xN1rHBRkcHAtFc0Yy5s0RUycnv6nL13reCI
p8pVeEMs/kiODXwIcZxzTGhKJfwad5+e8JKMSFo6awq2Ol7jDQkSSZWbg5WAOVhsT2YXVsaJQ86f
muOt1/5oGkkpve5rpvyynp9b0yWQwpynkluTOYRkhzn8sIY2LJS94+7XRSo7afsjHIcjAYSLK8t9
qmoW548xROTW0Hfo9qFtGUyXhdhoZMJghIlyp3x0ogl8LSavx693gf8zugZrmLFo91T8u0TE16a5
kWFzrilILCKpTsVxOG6sC2RWbvyiMGakxXURgP57pgxd2SP1BVIuERt6V77aAsu83iR7bXEFf1pp
NIq0XEgF7vYGvBER8CrM2tKUx8A69fztE78OGxl+nqTysCru5UuH7yWLevXe74qiwGij+fxpELl+
TRidnn3lvQrIbvARNJhgwcgw9hWWJUh8QcFifsVRBMXHpaud70Ds9C71i3KhjDWdBuGF9mQkq8eC
ufwzZQZnUGZL9dtSuzd7bbgztu14ZTVj8zmuGUWp+JT2MwdxIWGZ1+BFTaJJ05uDkaKykhFuOr/F
fbbPr6DALLdDOyKjx6bIRgVSXwrXhtiZbLTMCTmR8KrFzc4JtzQvru3GASYIhFhAhQctTMkiicQa
xtRLN4ijQrqnbL7DV8K+V9eDDoIslk53IYQLu4vI7SdOl0AAVCJtNzPp9nNInxmr1gXDeUJEsgho
UFXfJRun+Fucn6DGoo5KC//771BtqIT5o/7fDyJT0jMWfjxJIAfOwYU6/AYCSu2DqV78YnWGWMJO
GQKwS2v0FcaUKklCJML7ur58PR+z6Vfy00juGCAHZDhda2N4Eq3MHqZIhGPzb6IvRQYmxxGzrbd9
oAwA/oQWAssRz6xtypHSUc82T/At1DyR9WX7RP3+1MKCwUp7EQeqb7gBaPclwJB12OgjlqZ6gtrz
Og5Sqn0f/E992fwEGCfoLU9jV9IUUlXujHoUJbwBQljMM8/YdtOLMo6ExWWKqqRrcWtzmKnTZuye
wADuPAyuRLpUS0pOIAFikRPobVFuC1wLqgQfTVnpAElEyh8nQX3b1n8ietnNV8I7nCUpp/ZaKmhC
Y4j7micNF2hXrBdfamwDNC7M648YZHUywWQjpex6HHhdbnlSiwPwjFfCFYB8HbKhnH7eoFoLTVUi
w1h+WnNUdjhoRKmbzCE3QcFVgeCkfduzHk3XUA/TBbPk6/cQ4DGkP5LsY2ePlNQbPQBfvJkB/pge
Z3MYTf9JyqesV/cJc58kNuO0+UQ5NvmVsF+AO8C78zNpl5xgSN0dJN/CzwmOkktKcM+bpD4HNlq3
UsIeGRS3lxrPOEl1UAQXI5Fc8NCbVJHQi+mu/PZcvbhTGeJSkjpbNQBzSJKnTuvLahqmIYDz7Qxw
pzUwIMGWSaelcQFFF49NOA07Fbwi1PwPPOzGfjXK+B8DxiM7M3QPvckivobQyPtKZ7u9Jaia5HeT
cO0PCnk3UyvsarBZn/ZZtvpkYMWZi7q6mHFL2tL298rMOlDfKCPBvR3XvZZF6ZANJfURChD8PN7L
gu7ipJ4nHgyLYwVbZ6vTyjI17OVl9tNkmvO4dSHC21YoB9Df8AnNStp7QaZXEQj7o+WpUwevqB52
vihEmNtlQIf9bYae4+e0en8fApsp7bEQINp2q33cSc3bo4a5Qidm4g+6dh6eoMWfsTpS/86WuYWf
cGnd6Ez/xvSju4C8DL2qM7OoDHZXpllzAJMR4npi8/gyvl+Cr32uiOp9q0PI2lFN77JQRNnv4qRJ
dU48W7jPOdsY5tCNA9yY4mQ2AZIr5E8stiPvU+X4MJlUj1aUmfHbNOhu9peAFAGAq+RaQTpzoFge
a23v+Va1SblcrrWnDqdWiCvanWAw1y4rbnzE7h3LI/3E0bBNmIkZzQCgBxWBbpDHqDlnAgVasmH5
qDddGgB2anBenE1Spwkxhjyaz7erG52ZyCBuo9sU/Vy8cb8kGmf8ibnzMDlzCNuNrbm9ibfKXdCY
pWzJ76yq8bbjQ5npqQ0Giw00RkYb8L1RaabxzgQBK6mmVvMt/VMOdHP/zaeBH+JcMkpK60Wh736B
6VZQrhkKi7X8fsbISe8ewXucrj6cQ6GGaTt6ebT9zaf0ffttZyhGlt0yPOJD2AYZsf58FEjU+hUH
vgYJLHPGFvpC1A1VlMWskql/jhcMcvqv5pIPzzyz4FWhjJ3BSw4Dw78mxNHwf4SykiNg6x2u+lNg
UOfCwNTRAiVSvRqrxsF+29n4xANaFM7B3BQF4NMyAYDpYSQm9Z5/z8G5d1+YjtfOPVhlF2+O/0dZ
X8TBa8EEmYRSGhtZZtSMoWXMBH3xr9OkDoDpQv0T0xztKj1GBXGdoi738jP6OquDyWkSla+wTPwL
jQl647In165FlV0LvJ8w3Iky0Gek1Z0gCHE8w+c+llECJaC5TItxKDDEVS7x3fDrgWvusEBmMCyk
0ZalTvY+1LsKKEB+sP/gcNzCsn+pyjP58f0/IcwxvRBySIK3q1xasRQvtKEOu0Y0kucWZNgLo8GQ
xzDq+28I6RXw8ubZRTYrn8L6U/HRFWTnF7d/NrXam+cbmE/lRS9L2Imlh+CXv8RZFWmiTwss29yX
xrxW3Awa9DawSZY98MTiFFSYnlMCh9Vsg8gFfcekEIMKIOwjVgwu4G/5GM5TipYYNMo4miBvoL+D
xcvvJmSv5nhnL8Dwjp+qj02vLZVyEa0Brwsc0Nt4vnj3FYK9/73yCwv9S2OUOlmGX0TFXezQ54Sd
z/i9kdWIQ6KpRekHO5UiCGM1xX+3r/1gdAHoJr8Xh9EqQcHPhgG41ODb/9CXsDVGyFK2OVgNJ4Pw
XIeO9czf9+YbE7Np6eNTaGuKessBIjS+8IuK9CbZbvwjUMFRp747WcApQZ2NekFfV3x8pcp4EUMV
mCX9CGvEabaIQSjnUBij29aN1VQGOFHVw51L3Ej1svQMpIlyRkKDGbLEdFOKf54xvjnkXG2VFy7L
a+b7dR+gaMLkh9wlNAdejXGxv644O5qcMuDNoKV7VcSMb1bKPZ/UiWhouOLFAJtJlB2hzwZYHzgA
MM6GRdWs5ctHR1Mg65U18dPRBcPyUyW3ICVpMBqn7Uq+/YY6uWU9AWhcTD8pBFRVEgCOEDUQR1gI
J2vLLIuDhBvav30tUklffp1yaTiu7nBonON3VKrQH1U81Ie365BI0lDiiyyZO/NhM30R1hw6uJyQ
lk+/W4BKeR+fah1NDXJkvU7oYQh8qJrP202UdraGpYbFSXf9qsQYuExqKrB0z487LbsbbREuHXir
YlSuboRZeDZb7Ke3lZtgaWq08FEyTea5N7urzQAHl9cyyFbBfVGAVrEne4vkJVLwgCQRXHwdu31U
n13abWNlzGLr4HtJhT447Dq4qwbKRhWjPUx9wvOTT1Y26x4bFAmrdGpTxCHg5Rk4heGh8aUxg2ME
zIR9Mzes/Q7u1t3B+abnBHBY3FgwZdlDC3hx1zQ3UCXo/uDKQtYN/7Hdn23PPfFCk0uHC8oKdPqt
jBN1OxLd0VdFBMlHD7/79CluYp3uU0WcSXDj0xn3xK+XINY6DA+4bbRtAxl+GAhb6gBRWqhcsm7b
JVel2Y3leLetsy1Lq+FDnrTykf7IORYPx2PmvTNdIQC6FeANaBbOqtFBHreqpieLc0yvpAb8aL0M
Ga3k1Z6WA8lutfbhEduLhFUE7Mlf9YB+d/RPnQ2US6KaNS9JTj2W2LFYsQjuBOM3Foc90I/12T2W
85+lENTJtu0xhHxNNjtjjGCnN6Sny0IZWO2H0zqeru/89WyYVIskontE+9rI9YvKG+N15EqlKzRK
+CREsIiLuLmutCIcKlomiXzQdmu95nGtfsKv/pN4YqAbYBUFTLtGFRl9CmLz1gCB1A+z6yNJ5otf
uOFAfCyK2vjWwt5w4vUkd+JV5aaso/tzmWOfACA6N7LZCHNQo+ZDvKBqVaZCZQUIS/V2rCJNmnGP
4uwYdRaNGOD0iPC9ox87jpnMXJm/bCEKwPrOfKCemb/YkSmBxaF+C0N0F537YljaNx1yryApmXFo
GIzcdojyE3SkGwCz8iWjhPM/VY5dagzKNhw9g778DrX1rLPpFPJBWc7z9PqlKIMJD6Q0N3C4L7IT
A7v9nA25Ed/Y3CfVrHwWOTNaoL17GCUS+07L24q17YVWNJ0wGwQHseYH5zYS0nc0q6UK3p+ddoTM
l+1l1d5Qmn6wWlqjl0JCNR1fCPIMXDu4bJgMp1z2yV6ilddVrdTlKH4XeRk88sSXHXAmYB8ZWiul
apHk74ofIX4uOWPUI1ZX4Ktxc+DsDC+xV8KbSGtvJUcQs2ZBN7kjN6nXqjsYAJ4Qz22uz4wlYZLA
YpPvh/cU14TOzD42cKqFUsbEQ9EOUBXsc2hbqLRtZPRNDYzomSm63s0C7p3btSBJ6PNIEN8QuFMW
Vrv0wicmB1H/SKQ1/p9ef3AIQkn2gNvzEDwpxWAFqMmzXXlQTq7qDhK95N0QhOT7aAdV2anM3pSP
WLe534pkivqkqHeRs+gVzI7MN+iOwvnhIjdN08oPFK5uKMq3NxBwtetwuI9a63sr7L1H8oUNXvS7
MeJHFmdHRj7ObZGVxg0C/WKBJgdef0O+HR4gkC+LAmQZcNRhihhPzT2Oy+7/GbUN+JlFBFVOnim8
JH2QAP4R714uEESxgkH6GeF/Tg5CdchOTUTQKcdpO4hbuE5HqZpSRB3nmHuT0kuIO7ALDIkZD2ok
Hn4xsT43ryKO9V+hGVoh+FvFk7R1GNqGjXcJEfJECZ2uSbOX50xBj/S8YBSVIbq/TwVoJ/zT7V7z
HkL4337DNAz9dDEP1z6aw6UD0OGbFwrx0KmBo0iQMd7C8pdnBl6C0nHYjFrL2kFlkuM8ruHvsLjr
ga+C5dv+p6vDON7a8/KymX1qUQgnVrcNLUc97qYsfaS/2fEhmFSA2LZ+fubDxA41lFe+PobOguVV
0kvR/TGv5e2ZLvppHBD4WFLojCTSWGH50dcO7N7UCudteORbwYfGmVmIt0JhR2emyn+oz1SSVYR6
gytCevRgK1S51BXXwZ7jWujCNatZuD/JMTRpboweqdBMy0aO5wT6D9rcoLlPQM51UUQmYQh3FQcu
rtQd1Jp5OxSCAMhPUnsafE/TFC/bFbNkfVn6MKkfVSl8aio5WoB3Ije/uv5iyAZWdnLTiCYfnEA8
IMqfYWlM/uGKFXya/WDbug5XKyhC6wWggSlAWFCWrO8a9pLxOqbBLpMdD96z+cDPOvUs3sH+okmN
JvUB/i3k7rm9uW+QDEGKENmrLkiv1XlagQmOKs0F7g0ZtkvdhpC89h5E68p0GXIJ5JOQEjV3uA50
v8bKRVe/w9UGjwP4zby6tkk8dXetM7k5HViuK74ekYFcruhtMcIsUrm1YCgNOccOpfbtkHePhKYP
Ou5sZcsIBaAzqB67hdoYFHWMQLk5vKXJUnPYoJ62J1ZcGPwSXEDj+jcVX6Epm6MaqT/6gtzLyoT8
uhhh7upnMTO8XjV8NWSXY+LVigiOKVhTYneGtcJJoqZvoCQ4jRdM0ZULzeB4aVi3qMLcTnctdhRI
EiJAyWdAcoWkOj9BwA0+UH741iQlZ0s7u59YjItGOXX85QABmWZGjH5ywxQPqFDTA0Gewg/JdTX8
4vBn2zk+aBcv9OjHhRed4eu3eWVsA2K3KRDqqpqFAGxpIH9bRZq6W0+ddloUcz5lVR+/Lk9BRKii
V65d8FiEoTWnevcxE0Lh5qbVbCLhtrJD8PJ8eahzpsa7mCNtzQh8Gh7UcXR+KSm9RLZZkULhPDeY
FEEORzYm7WqUUi7SbAmwIp5d4u32vkXOcHxo6Tq4TCMgs13wgnp9oUF1S5urB7M7d1/GF64LhUjO
lMZGCvFGWEIj3esWWCvE/1YQtJG4tUbhaZbCC5mxtw5uGSXoaB2lS2OnzTwmaub06egzmZ+SBAYy
dTX32svi9qfcXXnZEhX3wDN4z9rGz8kXPONrqt8VnM96hg6w0C4jO9KUQIysQOM4ZAJGCi4LJf1K
ILDZCoh8t3WGJ+Xc5fbtKwvHQ2f0s+2A08Pr5xvrYfy02I+N3zQ71ZIfKa2RbLVK6gqnmIqNVzsL
1fN2K/DPQGhUMz9dW6gYgW0Zn2f7+FAXvMbAL1fuyGnJliZF/a/W5U/l8f6VwCSBYgCCp5MeJS9C
2Nu6bKU1uTJU3T+fifdJQbdnSJNEJ/Ks1n3qnQFwnMGfVjYCTfIKthaJuB5McRbRxenzJ/T6S2+D
p6vMGbgWtUUkM9huKHRtG42B2Q47Y6Wsmq6gY+yIUALxjY5duXLp3YAHfU1HR0pi8GHv9DeAwfWK
yIZjZbiPsXe1v31V4gS/ZgAjvsUzT2p1jVEE4f8vkxWZZNYJj32wBm540g61//qbCjWldwTxkToD
/CnzGOotKYSkvZkQiDFvGcYm0Uo1YIQXZNiNwIgT/jhJbBpkBM5pmJ2HZZsFRYyZkvltPfqVJI0C
NkbM1J8E1kj/t92g/JthGYpCuIbAsT+yd7pRVUoR6PgOXxsum+xWzYBcL9FuoNw8In7d8MOfaEWV
d/PARj7KnfuVc+RDikggH6aV0FlwQOE8h4VlO3PFjvoLgtukKOyN21GWIknuEpOlDx58SNg+i4My
k9EbxlO29BgVAXTtNd/G7e+TxzTm7/VpKwCfh/LyiuL3m0etvBgZvBXBCH2zizNp+5409b5NlUur
xoHNbSUqUvzaoBUCJDAXqCJnQZ04aYxhVlk7zDhCECo7uHyQK8EDmO4qEFesdOOIVwgBGltsQ5VT
YhYYs5XCHO7PqMvPI93I7LB2w4XE3Wmz5CmPEekoL2DLao7Y/QCaBW4HsKGtaW/WsZxLQv5flyQG
vNvP1NYbixVxlo73iHkjMv8Cy4jMYxIwp2Af/ANjWyyiDrqDjkq4V2HMPWIEpzgSCnapCGP5WWbc
UDP5sa9rPw9oXDytgSxritTf2Ln7YWQH2+rSBz11KBV4Q9b1VhvrCaqTDyg8S33Bu4xJXwHG/MoA
N574X3sDCxoQLmYBnM89QBDYFSC6U55JYIXVVtVoMiJu06P/HCGuJqKYVxsScKeMJLtBobV88nGl
KVYIp228lQTrIJWOxi+5s4rTzk/t5x8qn0mWgnl8PKVX+UUPGazP4u3racB8qT+KykOKQX6RCHWi
asLwGsO1euK3TQpZ67hijRw3pxF5zzaZn5N1LezbtbA9P74ZI2DVkAgJRePa4F9gmFTotmhEPNiP
GxffoD4qy9Ve9pBnWyp0x9XfB2teilERhjm52vRM696RhtrtwsywdFLxCXeZ2AEb1ukPqlEUxzDZ
lFoUu1OPyxHUYrJ4lQZg9mdgklYI7tLzuNpjqszFxMfXbNHu64Zcu2pj1hGJwfwjulBuZSepN4H6
jkTcR2mSkpH3E6TBrlsfLQ710vyGg7QrnBC5TyWh5g4RnH/g1oJ8qCfitpeBsE/vATucSxFS52RT
bydIsHbxH/Z/iQ9D70/M+i3FpHAIxqKufw0+rMyzhFmZlKCOO9ZWtXEKekkZH1b2wSU9G3F62XHo
5CRhMnaiaRKwT4tnsFgU7YFgBd41r6mzQ94GYz5LNWGvSQnuKPaX1NOFsgu1mVzmD0IqrALR9SIE
/C2M1elsOQ5aysoOz28SHjAeb+kTTEcxhXhdJbZvYAXoVWIRlzYyfq1z/DiD8oW6/yIaynfzgFUq
SMbfW9mEOxRSPBL9QRs7MF9z/4RKAPbJEcZY6FB5btSAFc3BnKJ2uvTdLqq4gVoCv8cpSZ8pY/Z6
3vXYpV5YM/X9v7FXJgN+VSMkVRUVA2VzEXU9HeCm2HEXPOwTzXIC1LA+Sj688WdXFajbQuLTm+VI
3kS3/6zE0nKrtId6iwK2f2x65j1taTPvacE1MQp3yceAekBTYTU8s2DETsYks2fORqYUssh8nsPH
g1PP+pTWdbNcizVysBiYzuh1CcY1KZsGlQu4lCl7dzfle+Z3gSyFY2Inz8PhIgzdYPAxo/b9nWDE
wavYds/xU1mAPpEBXZSuEKVh/tWuNxqzWa662eRXJW2OmoqI4aNrMMBfAfD81lFuaSzVwk+sPn4A
ZQgENyc/v1VDVPEU8Hng+AXTJNPpoVnmILPpzoajQJcfTpR1JAJiKLya5yyY9qYWCzyTahLYzGLr
b1HSQuhuR4smcp0ae3xEW8FCwx4JidvZLnggteAjyzefv+L/TWergulNuBcUZ/YJJMMMGXkLqW88
MEgnqqK9+zxaD4fkJPkQPKuTft2k1osemcropMJk3D1VSN1a5ZJMeXq0msQfkdB24HMFdH+zmah5
ZVCbavNJP1VXyypaniXt88o48EQyW+MWJbMJ/Xe218bXNr3og7Y/a74a542/GfVINnO8hNHPuNOT
3RXYCNqfxf4RRWqonWgQKNkjJ6d2OXFWKr7YowmcfK27TwWVxBIhxdobegfE2/dlqVabftuiRBxi
ZnnSDnu/mjeUefTSCVcqgpSclTVY8DS7oTI0+8wDL7wyfG4wO14cyUMRbbqh+O4X8wboHnhzEWaC
wCITa6xAVRFxMFoB1+kXT67Jj/NwM4wkoz9LyCkp7tJTVmSJLpaRN1jH9u6/sy1fVcccnk5xCMnB
SRyJPTmGgYJKPKhetFRfGjmAR3w/33632RoZDjqkaiQrOquB/PA4Z1dCkPj/lgPnc+Go3nWwjDsl
NXWlMOW1IxJrk8LMszytmhYr1P1kfr6614zyG9S1SaTN55+HE57v2C7SyswprEXwEgOZE/gSu1hx
WosFIiL3PHeBvuQCEE7r7AvQfbCibrxQ7cLKqgu0YIANgzRfm56XNIENgr6PEq+XuNIzpvXH44mg
S+wZ5FzKuD7ZOHkRafCPyCtUFOWCHw0R3/A5O+ZzEZJzpGvG9atqQrFgpn8jOzejMQEqG4fmuIVO
JXTpCqesuVOfbVmZ9n+p7hh+TjZ9xSOwyy5OTN0ly4Wy+H8nOHCaUbVzhRJHU9btmvyb+HgsmQcm
AzbVrcPy5Hm4oja4U/b7/WWkyYLMJIL7HxSQ8zmJ6/8GzY0N32iJzXdjcSqKN37kRzCsKWlt+tF0
xHQMLCRkNoaw1NSARxE6C3lEkjHtwKfkOHmGv/MfVoJKx0Re4DztgpnsfIXvKhlHPydySfsMpO1d
cDN+Y4mpxwtS5xBajTfZSwHJImmGROZX2CEgBCEPAI0fGtB25WeiW6+VA1L6wdcXaY+OVncz5Bg7
rc/Ul7Q/bkqtZHpHW0hjFniAcoJQsgihx/FHo2iHNOEDjlen84D/jPXcGKoLf7SUgo4S/x9n4FPo
pjrsx0l9elg34JgkJpk3FIikWA6CiKvVsDCR9zDoGh5NPniGU61FVSJcqNY6Kn71ymEVl3eI89gf
mgL7AVQZwPo8vyDigwot5AWFoM/DKlO+Bh/NIV13Kdy3Fhaic6dgt3CQk3TakyMtYZcLT1Xi9UQ/
Q269UtYBChtlOSwU4hIk3k8LM3rZT1VYfN72EUfD/+cZxpm18z0bziUEtMqWygkk52rFPnqdNStV
9ANFisgeolRQwxmE6Vodeg8+tidoRXbR/9EdSTymdsqryXpJ1gnb4BaDHFCneA8CG61egcTUMsvk
LYYJsqIbPUljeyH50AXpMXeUZit0+2R3+L+KtGD1MwYIMTYGrCb69J9YWdAffe03H5wGzwM1vRmW
4+3GOxyv7NALEZoGlOdm4sCp5vexV74TO3syKx3zairNb5L87+3RpHSyB0Nkj/BDPV5w+AokcYkK
DoZ5akrIccE0e1D4xfp6pfSdDhv6k/772RqK5lZTJyJRNdLOKEYUzWmPyfhTs+ttdFLi5Ccc+zEI
7wmceX35udBS4eBk5ajHMepkgwq0lVbhWw460PIl36DSN7M4OA38guOWxfqoauPzk790LYqzEPd4
ZuMqM1miS706yNnhVlMM/2FYS1KfUACSQpLzAx7PFJVBQq9OcVkhLimC8/PaqBpvAPJUFZv2TTP/
Q1r6Zn+rkIVkJPv3nfB5GSULFsJ/wwZZbFDWWaFdqIAizeuVo99HBm5JufYgbe7t0Xa2Llb04sBQ
LsxsgZdJM8M3GZzd3PKWRANSwxNW3A+I00QqaJYI4n2X89rRM8xJFrGLIvBPs5YTNOQ5EuhP6kIi
J03vQ2xk0jQQBa90EgbQ0tJhg6eAUJ09rwXQ9gTbT8LQLjp9xTwgtJc4/YBEf0wm8CsXmXnlKymN
bvo6KD3ULLKLWcU2DFKA3SGeL6zThSIKiE9sbdi8C7nCL8yMsR/p9vurY+IP64sHIIHpWq7MXsZl
X0q9qIWr7akvAsalrWEHbdjFZ7/KlQaG5vNl0y2gWruMyKzs8/RvN9l/IMTlERH1wpkSGHgo9XUP
HPTjMGUqngRaQo8kxmrbw11wjAgAOwlH/ppAg7uNIfP/oZ0HYPUUanLKG7Z4NfPWELSiwE169AJg
tH2e7LFQg3NpGYuyT6uvt2wFaEm1dJydAy75ggD1iRfI6TQlKQinQsG63KgRax2GQnz/Qsn2MDsz
xK+K5YQsF7FuEfaa1qENyT7mMzhOOVVWF1lZzURWavtY4RdkBGIcrLq/Dz9caOrErNTmSyjzlLMb
pWqwxRHkPJ+IwGOBmthG7GJQhMuDVr2zgtWVhwGDAzMbFxol9G7OdHIfWHdf8EB5WlhxBTxEZpsi
aGKNHUmjpHjuqVBVo9RvZdQRlM6Z5dAj27fJxiGq+FmZ0EaxRWs0jBjUZmAx06Gv341sVYMR4xTl
3O/5U5+31J/6XJf/jbASuy9oyRy2dZ02ebbIPdP8LeiPgOG8ZshOq8xDhO/c5iapk96od7qosm+W
BdkYVfYqnYEnilWcw2KjJaniq6T/pCl1M+qKztRhc4TnCA52HYAfDcgdnSup4QCpjomc4K5tmY4d
oOhsN7INq4eMC4wHbRrYyq7qN7vwJTcH8fdcju5mWf3uDg82Lf+F7dpZgYhPnLZoqSZ7Xw3hSYkH
iCirogE12KOynhb3vmSKSR9hBAxOSVkiwhVlsgYvtYSFiPB1TtAePalhnishvzj0qUi/NGt2NoKM
uLUdVxfQZm4m2/RCFQa7DDk8HJOB9FNngwYTOKHk/ZCCBdgQdrNP0Yge0y4QJQ0STuk8lZxkKCgN
c74dSiuNIDM4Ag3SEHUBDlKR13LlUCkiRRfrsYKpgga8me6vI26nDsHIWYgaFyRiVU1GycGCe6bV
3gI8OKfoSEEQSLOhF3uQjs1Jk6dMu/wCvhWyeso5oh+WsOKvXdjixtjg3DuJLsDsYwWQnmTn6CYS
arRqwqkhDJNKMm13a07qXd56Bgkf+seUWQ/cDITltPb8E1DhmOkZHwxmlUs6gLQMGkkNlbaVx5aj
Sv3M7D0ExhfoAoJmONndVFxrFtVE+8hVP7Ta+btKkD1XrK5eA5sdoFF+5k/GaSg9CcOsOMLLaVZL
U/ELwqvELNqIbCXRvdTzgMwI0SJ4g+EcqKkST0XgenFvWGDNVzQbUM5wf5RONapnrunpO7mQ1BxU
J5L8jWl82zjT/s4OEfjEmNSiywhsfEsND05kVx8JhtVnNv2clhB0oBwbCueIm/nXSNQpi/VG5W+E
BDzNK65lld1tX3NugYggQz4nteRDK+irpgzCZPSEyxhSzP2StggGy9XOa4nYvTNZ7kxgFJXYg4sv
QUshKQiQbmEBxqsKTOI4sHVFE2oZ9EPpr5kPXQKBKIwVLmFWrVn/UA/15gj+kmOt//1Km1JO/X4h
emTe2A562fdQ4jC0D1rtg+H/gSdOSsqWM6nynXzs8DQU09AsX6mFiHQf5BEhXpL+xIigB6WxgrOp
5pTRBubZ6TB+CTz0orVJgKVK+tGiGIll6Q0aS6hP6SJWyxmDhJNTyhTldEwcgTZ5HYYVA1n97VcZ
00MD0OA4/iBnxf534kNeF6mLnwvx6SJrd2AdCMPltF9kgi0MzP4I8XYOnHW4CYI82CvZP3GbVrLD
uGVl5N1Cefmd8KynbZhEdiecK/ZV1BtpSJArZmVwOagZ4HUZiLNO0ZLvVsfy3xqTBdKPNPIoGvL7
17pJHZJFU/RAIf28MSVH6ygtkWgLSh05IPp/6c6sPI9mDVRBLfQSLgwcqHbH8PDzG4gGy7Iu7i2k
KuWGfD7xQhUCco0nrA9OvBdCV0I9Hw+ABlRGFF2R2NlqXTz46EdKxLslzj/rNn0b3TuAN60wHzbR
kFViA4V4HeuJS7j29qg6ydzrUySdvvz/mZFpPn+PqGrbvCrHwFrZu+G5UjA8dZmcC0gfHKIEm5on
LjxapP6d7T5xLvHqlpxdk3AGJCo71QDWPEpr8/AOadI/8WwI/0+3GbhHSBUPNMqlKPAr268b0SNk
qh3/hdNbp3kwqDXIzdQYg3yW/v/31NDuj8rdD4YCnXunuGJH45VvI9MtBi0Qgl8cNh6IWTxU4WuS
vAM/ohKypW1jnDSjJI+UrOY1PhBkShWIgcspU6tzpO3RFMRP5caiQUSArB8MqUeakuJcyDGVaK1V
hVpKKq5sActJ6R6IB5f+iqmb9FDDmRtqlMmc+Nad036wxnFQ6TcAD692PROseWan3qveozy9XAoS
0w2fD+d2tXkITZLVKUQfd4y+8wXlajFhXfFvGzqOHBxq2ps2htXbhsHkt/sCk8kzK1fYc/PJqC86
b2J2+QPFYfbUxTChTvXx4AnK8kblmw+/0StCeZO7lHP0RXoKWreldegUriUcGQCuro/dH9/RYMZj
R2b563Qlmm1y+GyJcMWKvcgVB7bwit9Z3n89Uh6N59ENqoVPd/STh0dy4bijY807DuGGsNyPvEho
nOL1cjU8LeDs4Rrm7JWKux4Io3tDF0S391WBO42dwEfcIsdjDjKFiE1p9VQhupy29s9CZHqWVIS/
djgUMDVpZqF1wIkZiXjLETA9axzLmXIMpt4NK9M49TD24n5BHauyU6KEAB26z0E6rBkxJRO5n5Pl
QPhoJJIkXiadRkm+W9jvufTVyBObzTiIB3fS8Cd4sOGwBliU0RXy7PnaLbPuR5XqdwyZ+95iTHWH
TwMSnSeTAyMuDfmTJtP9t9l2MVbltlmeIXsfdQpbINzDjVILKFQ1N1/Ehe0O6zt2PKNc191baxul
kfvmElcUTbQA1p2fmAenN7Lp0+i+PWVKhlDWXNO8YGT36pE0ga3X6B5VD39ZxuMrinmTdbPvKZ5L
hDL/q+JP67OphfDyjEFQ5cUVVceCC4YWu964Pnnz8MnPWo++KX4DsK6yfPAvFlkjLKYLnvEuoi2x
Tslgy5R5k/bKlJLjasF+/KLxEg7YLJMnqLyuzuc16DI8+5/UhBW3JSYZ9YtOTW/ATI6/ZWUVjVLx
YZIgcCTLOYV41XbQLxhtwwZ/o38lUjBRLdw5L6QA5ElTJXmJkCn9QY+Dj6bJzKkTchsUHgNLiUJ1
vL1+exSc738avfDsaFGtq+U3oFmPoeOLNo8Oy3eGJLacz5zWDxYvEfiPGAgwhOF5fyyRvp1bbfBy
c8XkolKDJUF+wX7Cq+6qi4Hv4kg5nC2KGnmYRUtPgG8A+ySWuCqNc4NGIcia5vqj3N9yyryIuA4k
7j4YDieoKZb5YzAayLsGtyW0MV55ktjBzh4jaRwEhZhQKYvcp51d/HqVVmWBLHxZqeOwFCZcgzz2
vaxj6vWjhP1k0g8hy5dfqxR7OgF64MQArFjfH4+325yxuDyxN8qXpR4loN69GtfO4j/PtEgNPOZG
pfkStsDkxngZ+v5gDxJ2B17zsqr8kqZc5scUhHWKCuPl4XAgjBNbZkS43C0LNw6PHHHqrJTXo6Y6
Pbjf4KYuU5Hc72N7KqrnTbHwRn7IcL6KVKJ7l3UlvXofXw0+WrJQRDn30kZ2duRksVc+NMvEHkPl
tb/ia27NCcgjVM8Eh77KLDAz8zCdLAIN6Nuj8JqdMnDVP90Wz7O8FVbTDzqgu6Si4FUo3dbPvgzP
2jlXdWaSjtRwCc4uSI0yAei3A7cnCab7ChSsfwNotm7HEgHp1/lDo41gneS78x+ArrWTp9Vh/O2v
nbU9uZ6pbNOenY6WXijqRpaoStKCTPnwQ8TwsKWx0jZbGSB28HRhPV68IHkZu8uXFbAUAGByN1RG
KxYaK+z94eaF9xeGyJp0mB6WjJyk5gzl1sQqjawbBe28KVT+ef0IAlIWyjGRvROKAS3dO6DHQQxv
aRS7576P+40YRsDzrS+09FIv1dL8CfGHJ83dQRjeXUvKjWpMyZgiomPDF4CF9H9AqWckneqLUG5W
Zx//cqgQTZjuNjAWoYyUjN6RDl4wXUHX4BLoc5AAbwXY29plZvZ+k6ZSFyrtLmOIFsd3MVo7KPz3
O2LvC32BwCQrGpeZgQuMHkdV/GYab5MLIRVuDfFRJ6Pd+gwsO5EHOG6nSpwRceA4Q6cxMomPJX3O
pTT10ODEnKe7TYRuPYkhZ11bNoaiPlRQ9Ndx2bNd7TJFc3yotD3JgHz0AaUFPjfMhkcdiHBM1n5H
XlcEK3Rt0q9P+El89Q+7Am25jC0BmtDAq8PRJgbniHPnVG5FY/tvE4CtgjcthB3+sZVntAMccOM4
85MKcIGdMv2WXt8FDNtwLrpWPjSJQTvKsbxS4LiYzJwfJfNnH1wTmmX4TbaT2iJ5LwPfWsoroPqo
TFKgob1MZTsm/nfZJkH1Q8P0V1XfYQ+0spv87+PCwgQ9ah5OqPR7UTlkrdJobF7I62AgrpoP5fZM
/2U9MRu+dhYcL1SoQewRL+V8u/ZNAToFAqW5tKEby3LGi6fAeHNWmaAku7BUhWm92C2zHZGHNaec
6JEw+W6GZWyicMesRDA4u8SI2ae51uE5f2QrSSCjJrgDVzInSPeg4Cp7I0LpbnmNo6hd1nQvBm+F
8UHEH+pT9OMRoQun0UM7Uj+3XwQCM0HPomPOu/iWUjepXlJkn7r34i1TPXtYaa+RcBy3j2bKvPz9
jjyRqTq3LUyr46AE7HokF1pTRgtZc3XTQl6e9wmrHayy2gfWlTUWtROwXoZxIekKbfKySHiu6TcR
Kd9bdwHzuPr6tf1HfuQEBaFNpSg8qOJikWjFKQ/oGUprFkXMnGAsZ1koheFYvnI1jYl82813w1ij
F9qTIdG+RkqMNZ1RopfVuJ52hM/uvwBeusJ9/ZM/zh7AzquBECf9ayegk9qPimdYGI9HeJUFbulD
BU1fIuOWvh1Ov2HZqfBxhq0WRz19rNacOjz97otU1RftjTEBezr+W0RJmN5rFREjoAol6rg68m2W
LJFWP6tBi3mkq9nfBGo5UejJYBNeYTMvVtFM9+YC0mi3C6bLQa7UWU5v0JL0VhClzGIeQk9/n1AP
QYSuUIvgj3VFJxZ5stZd1aixmGiVh9CfVF1KiVSH4uFg3/wBt81VwCgq0cVJr0U6Z9smqAdMLE5r
EFysljedonm3t9OIEFeEm743HX/gwHDniuFBd7TLaxd5AplwlbJIm/lmU1jchEvRmZtZnOr1wd/x
iZanxoKlgkQBe+mvyP07iKJrF75tK5o6SZs7Pq4g21+qdtzbdeRCe1Wg0z4OFo3nH/jUOe1kxEik
CxDJtEtJhQk5zT5Fe7Yr5YrVqizNRpKYotvj6/XDqOJMHsMMeOLyFq5wqN8+xi9nIWyJFg+TDsJZ
CpS+ZOsZMr1IoiBUxn4ZranOqerwRyOOuJ6m7vndNAvCHhbbWjMUJllY8xi0LFWclC4gK4d1V2Ah
n0G+Onj3A3tvyR/CrjzBvYw3AuZDbaHfDKRdYyuCAhO0+QapwdMsefVnxsufUBzvlozQI+VzN2AY
UUC5suuHWpko3pcQKPmo20uVWnEvou2M6/rJn69lM197xOTSnAX8QDWENnr5mkcEMavVCj8Im0Yr
Fnh4+eUBFxaxVsvIjGz28mNIu18o16gXQzNFoaP+mvFcmWNBHWjkjCKZsyVA2AYNWv4wEUPHuviu
M31VW0xGYGxbQkCXzCacUmwDSaiOUv6xXvGQXfSf8NOId2Nh6hwHyhziFnyETN1+qnFKvBgIxQZD
5mkU3780/Tj+wTwTLX05BPk+nUVYpcfXkLEr/XmMHrVYjImZdi/ck+aBWfEakHxXSg5F5bayQstq
NsGcOHB2zyruCdOC4k0LXVulNr+3yjtl2jQAPDZav1w4GL7X3GN8ZlalDo720QWJJWp/AAUzkxH4
T9/QmUyI8mbM7KL/yCYxwx212l1qgFdqzjaTsLWtoHwK+LtPkEVGnf3CN1qkpFb4JQoCK6Pppllj
XuMOZBguPSzEc1GjtlgujfRlAEIdUldhjjPYxhmL51bxpaJ+eqLkugQo3a5ft4Lh4Xwgb0y8MF4W
c71r1gfjFiOxdXKVMvxx4ZCq+KhCWmnKMTn3sVJeFMYkD8zmp8jreiA9Dv6XpGr+SMkKHdrILMeA
dItoUU4BrFV70j+dE6Cp5d0CAv9tkSIJ47V/vfWkJqxz8dYXJ2hQr+eQ/bgESJeXCyfIIjhfKyNf
+Vjzy/Vc5MUDkhXX1+5ile7u+jGdD/fcJjyR2K5XuMG2RtsWIGx8p0Tv4sah/r/fite2M88IKi1w
+TsPU6HCjGOLk07ZCh9Zn5U8if/9X5o6giRrGCn9AhbISVGRX4TA/U52JzuQMnryFa3D4Lt4bmUw
Z+4xxiJwqwO3y8fZcBv/vHzMKO9Yy3ATXxWaS2R4FSTBNy3q6ODBZnicaXWiQN68r1h+j6QTJQqP
LO7AOWhtDIknFjSt4BHEuXigo/J8LOLG5T3Y1aQWAdqIG3Teueke6Y7yxkavr0AU6T8E9cZ6ERhc
AAySCJb8AMCpNdGCdVrbc311gwex6oOGfJK1otOgcEMjs9UKI5gUl/gd7enUA121+LNjNHeP0374
lA7nkuilRXXXKjHY5yr/n4EQtksW7C39bFVarpG6Od/Z80TXsYdxTEI06/Yc3kzvGsiSmpl8L7a0
28gbG6FYugPwhqiVvzzfaAgQ50vUOExTnLjb5VmPulz56vumz33oaS/aVq9DoRSBa/Mc4+GVgNB/
LCuLlo3GcMyTvdBNeo+TzYea+CTauQRTkNW09R1xbV1nDNwAL7bjQUWFwMTKFtJI367nSPyDrjt+
M8yeI3l6qjbcvjLlfvEVFgCEWMI1eSVO71+J3HjlUZK929BTtucR6PmAJNTYFUc+rZBd8ZKnojBZ
xK2Jt4R4MSyUUBiCmEdMHpeRREBpO25tGRCg9DCPtMCqzbh7OKFGIqIJKe1ywDN1otSOsOsHeMgy
bo5nFl/ryiXO/Moi0QcB/yv4AyMZ/2TB5D6Qu/kRuW/cBCoN28t+94Nu5fdOXKMi4iJTiccgmnxu
uX3W01P6jLZ4zPPptchUj/TcDSWpaY/uIiF6wLJ9Evh/thFhCFIQYIieto4/5dCIGv7X9QLBhJyA
gj4XFSeWVCCHsECS0J4lrUmNpk2u4T+eNeZdYJEqS3dcNsQ0sFAfbLUjgqhXp6VgoB9m2/rCBF6d
Mw5DIN03nK+ytRlVFsG/zv6hiZRwx3Rc+L24vj3CYF2lszHwsdbsii0iqclP86fhLnVLAq6071UF
q69+MaaPbrDpdfVE8ttkxnKunTj27Vp3LbkpAWj4Rni7h20C40zNsCeYO6yikokLr7PM12ayIP9A
qU8Yz4p/yrMp/+1seQr2cd/OtxirWGCcIjhzhgP9Zg5CiYG7tc8I9RPYrzM6+4tsM72AhdGJS2k2
T+pOr3UmwAEoDe2/G6HyK3fYV96iBwEjoPOf863POUhU3u+eOxI0C4v499mugNyQZWzGPk48JuUd
zYpGm40QOKyMcfrabsjFSQirGHVKwnBxemo99TdXG/21pcd0MsjdE5sHsKwjm83cGlkgbNIIKWzJ
fnop6TroOoE8v3eb5uKetU/xrcsbnbR0VX0GGjruVqtIuiWOdD/11PK63fYq9Pz+7oxwYKeaVVQ6
g4k2hDPvUaZ4IVdnvuGKfqUK8Q5+vr2/hp0VoNhu6CdeCWGcKjf3KcI0bFugRrQ/caYoSU/G5Glt
6s2cvCQ3kw5cAzY53N5vjZXWIYOhryghVs/MxzmHD++xOjLe4NVgdFvh2uEWiT1CUilf+m8bbWBw
pS3z9KkkW/lgQpfCr2cy5VFtamSBC6zpmbM4GjLoK7D+vxtKkH93pVpg4N+Zks2/H90Bz5UpRhEA
uNCZGmobHfyh89gxRQcROdN/I6qMBJ5iCdug41J8IYunCOqtb5soqmweBJUv0rlw4wpuJDuKldv5
7ikoh43v6p2g50r7zBHDrFw3TVbFzRZJq4fU18NLt6PfMmT5mXOZAasBtQn3ZZaoZmbfFdtEj2uV
l8XLwsMau3HzbxCPE9d+r1F8v505REQ1ph+bqVoClijwVSBXQBHjWSAkv4y8RHLuKOU8mAg3lGDy
jioH55l3WJyt+gonwRlQcBZ09aLIRbA1uJfSIrtW2S3kX+ecRuueViBlPpxY6wtDXXAt9ZpoAKAt
WxSvMe0Fg7fHg9dpy3cT2Lkg0mnZ76BKKmwuXSD/KzfdEHl3G8Bxf7awnNBhba4zebP56Lm38ecX
i/wSCZ2dOua+78yf5o06oJxVocOAaF4IwrdwrRzuchqYTOE40LAX7gja0xgy6LioRC5nD2B07Tvi
usVqQMu3pnZuqXYrcFfXOf0zizO0zl2cBQuvqORYIr6m2H72ow/kPJQO679f2VsGSl/lJISHQtpE
su3v35JiLLl12KuCujkswAs9zkKCVtSgyGUl2x3m2RzDNgHBRUqYipBoJNPiVY9GHT4suvmL96nw
necR5L3VLLz9pTaBGuUen5FMgTNOHm9X4wSlvzFBaLKMWxviOYGaggZDkONtFTaTl7P+YIGzT3ke
C8fPbwOQ/UQdWyPisTjonlrHA/D8nGyTBQacBD/qmTwQk0BWCq/FhEShhml4I0G5ch3ggZpWkEER
f366DS/b/v72ccbE1L91RK3gAOtcpgikKl7esci6wMk2hK8XM7VrG1asmQQKa+5s+pxotax727cz
MkSS+6HlncydR/BiUIm0EVFJjdx1oHyimqeWAPUbdZEoT2NRqc+20evQtkir7pA9vKfCIoxqDQyO
KfZIFbzhzidfeaHt3T/JozSwRKaCPqsf4rxzBnqMfK+EFisXuzHEvmCfLgc5cjHVG1onwGctTvD2
M5E6WVN4nOxiYsm2h4nbiTkNIXuRppOB70SyCSDcuWyYXJ4kKrwwnkxyrGQ1nec3WDDjGFDBUVf7
wUP6Zcc4kA2uZ+UFYrivwVNExbevXDGbt9G6WTkJL4DvR+BgD/X6rHZSxYPFP/DtDUYfDrkI2uKQ
LEo4JUnggtZkfZe3Wqq+nP1YkHJIvVfrnF+K1lToGhtDgcKRwY4FGgHtrPDKu7OWW2Zw7GBcui0v
5+Xq3DcjbmQq8mZ/TpubORXcebUOORHG6prL4vf54Xz2WB74QkbTyvhrfsI0YHwt72NSL9KEw29L
2vLa0jPME6iKZsN0ndWURB5s27sBVPjwn1REAm5rp0n8XbPGBFJ2RHp4l9wYx4CVoDuIFzmrxHHN
PD0QeD9DReoakG6PL6Be9/fmgQOqjwVtmlhNhTq9vcLG5R6m/jIwwKafKnA+u6+O9lIrFpOFbx9v
nkFgksHQIBZcFvj0ugNufRjXMukgd2S+yUCE/4eXKrEaaUv/kj5FEr3ZlqSxFZ+XmDyQvMflgNX2
UiCtFrSyHUslY2IHc8g2YEJ2VvpEUF9MWgY46nVLAopLE2SwoVtu4tIJeTVOWWbMREsdBhDZwVG8
f1tzXfres4W68N2Rn3gKhHCaTRvurfx0BeiLViyW9aEMnPjAMzwYCCLnPwCS2G+kJIxxfjAhGjE/
AwMOzQmvCOg5rr5F1W7CNuAQjivxnNGwN0bRILWwvcvU18Sv3td2XJjmnjOYfJtDIwqKNk65FXJG
s8+vwX68S1zn19srbZYL6cmam1qdYX8EYgJRRYJ0lxWk8ue9mCVHH82AnvDnsNPypaqgY7FCHtk5
dNlAlDgDBzI+hML7fffXUNkTzJ6HKfut/FNkR5U9yX+uIk9tjLmDLQE5rzZVf6PVgkGBS7QbxCnZ
XrPmstS5aaxIdpN9rU3N1Lui1b94IyauvupRQuZijFWl8j1uQZ/LcwpQ1HpvcSdfux5vUdOIjrak
TBZ29BNRg/O1ud1jeBzyzXhuXh/kExIV/VVQIBzTkXk5FTKGeaQsaa9jY20tEogkKDk2F44Qf0d4
6/V0/uBxz9U3NgHi5YKwOyVR4eFSn6MA7ImQQ4OlZLiw92q1Zqwzthl5qFi18ztT7sSrDjlu6M+P
swdtaCBGxZAf783VjVW4AyiA0qDk1roPNhnFmIWejIfwRTu6vRw2fZiquclN6TvaiFATCy6cOFZd
cVRjZaszKkrr/Ve1LuWRsCh/9DNFPdfCr4Wy1j7BWwSqFBKDk3GQzIRJExfSjso7jTrH6K7vv28S
njhScpmfVz/xj50wTKsyOS6u9NOgnHqgpQ0vtLfaRX5hhdYAmKzZbLtEniF5qOqyFaokAELYyZwF
hw240CyMGxzMC1BnyS95OhMsnagoIJKiqsU+VhRvxGIg/AzPqPCAabeOGS6ffj3HN/6x6N6cBOU4
fXrmhkFODk3FlEXesqjtecZ8RXPft+mYbHyubcEmXAfizyvOv0e59TnxFu78kfauhHmhWqMwMyIn
k/I8laL2T4YeVAHcZtQ6CR3+DNkJo/qw37NmCJpcLppfObzc0PEdcBvYyWgKfjLcyjCex1dS5eNY
c6zhjCgFxR9SYj2VsCKAIjis90IWi0OLIz9E9GEZo41+N4ETAQTgECuUSqzUh/Pj13oGVctjH9WO
Te97GLkFhuSHlQ9y7gusqGv73GBYIiGHYu3dgTif9Jwlo0egJC5eD2fPLEik2NvzZkq9leSadXHe
qMGqkEteeDnrgojgCrKb96i8q1PBfo/ZMEIMD3UR/s8KLgNIJ6HGYDAmud6pgRba0DnY0VLI9uEs
XyqcpIcTKAUPcxVkrAL9bq2KZ89uD9lxZikVIeLdTiSad3xj5lyISRgYsM0wm0UcSTx1QdHDxZoD
0gjY61VgKwjL6i4CC+ZkCVDW/IJCnwH2lbJjHZ408vx3Nx4B3pbaVYeZHxvRDM+Rie/2PbWCG/BJ
DODTlV/D850k3v5GNRaU/usJVroi2/cUYgaWVO+ez4KJ5WypN8hhfiRxBvLWbzPq8D4jNeWN+xzf
NLtMnfVB0MmR4FyJ07XMmwgj4O2J0uiKC6mVVeOACFkLp4XmrRTMmi2DD90G1WpjsjvrF0Mi4VJk
kgDT/vsIlQvP8xBj1zvmGLZKSI4n7dMIw7/2ApKYiYXmxjDCt/B3OiBNd6WkD22Bw0/9jVFX21Wd
vh59WCHcFsE7kVHIrIE+18ttBpU6kr/uR/uK6eB38LMd8t8pEFdyj7hA2Bzk1ed3h5fUSSBKbTD3
ZdICFEkxMXPcE2M2FaOwA2M8ej35qrfq0bhb8mYzJAt2ethlVxnMsrQrmFukVTPfS55zaX361OP4
yNTiE3ALujTko+6/51f99x4zBSxC4A86/ibpwdxqPyQTSYZatzYbm0JObpPre71FespmpfJ0Vxq8
d2ClM6JfvJJHZPYbSWo0oJUvEG3YgXhVGWjzTcCGNE2flFTRbNj0XcJ3ah7EzOAHpK4Tizxeaag2
pYwXaE61Mdi0b2MADDVNfygqvISd32gocCfu/DfhmSOhgdo87Ok8bO/GNWNQfwllwao2iKIhUgxo
AO+NOfQwNL+7LTEChYZLifARM1Ef35W9pLuN1rYLtNpwhxoyDM3PAqKkVAjGtBdO+GRpGpWQvSQ/
hSodEA36uREIdMm8hoje6qygKAHfhQtF2yt7I2ESo9Tpv7sdFrw1JzsN4l6aEaMAdPBu1eNKi2yM
6jz941HIz/YnpBYG+5T6KnFM2G+Wh1c8n5iwub/HwUa/qBjrecHupGdq7b1/TcqBVeLZKRtbjb3i
fggSOHrI5ytJv1oqWbZUefXjsUzfwT4mh9vda9/i2tNw/CnAgpLNhEo0aKiIaKcVT2yVh9UKx1sX
TOAqaGGFn2d2DisQISAH5DNlj2I8JXFxu20bFHUSHBtztLbN8oIHiPBZMZKKQeZ3HxCP9mgtLScL
N19C79z7LoixLcMsWgtLbGvHqz47I1xcpWyFO/d6uSYgZ/I26fwL+q0yehrpXKFmz7Vo8+2EVXkb
U633pOatg0PPVTulihVE831L9FRUB/0pvCu8jyw/r5xpwNa31DRCE3UpM7jx1wzyyFkJ6XmRRYcJ
GJWrZvSK6jq11/nrYPA8rBcQoogxBo1F4bKtsksRo38Gqe66XxdswRea01GafiJQiXMpaqQkqZ9k
pem02lC8CZmgF6u77TY+ZoDLpAqUUJVP/pX8j5/1f7jkj2NvRuNJTlGat8AjZKm4mAFvu2ICjKr1
aYC3sh9yHEry8lTSuuPxznGgFjrPPEyzCQ+heoZHUNM3m6ypaRqQEnRMPSdeIwmdK/i4n2o4SW5h
aj6/v3kjBasgbIeIDi6zQeqTPHM8N7jBiSRVbZWrBte3lh/uQD2uETQhnq+JvCLw46zRSt6lznCZ
bj/pmd1kvru5qpEgjIhDufAqWV0pcZwpw83VpWvuPHSw/laVB9odwPvQp3dopBdbQvqE25rYk2+k
brwCvKbXh+mz3ZE8nx8Vo1Ji5909BAxFG5ySP/oESuzZ/CxSjQcQH+YAytmpCqsUqezeWA4FPkcc
7Pd4NAOONg50CxwUcclX8k2DL22b29yPI24+PTShcQu8f3+XU8sipla8S27Hx/tpb0w4nItbtxOo
lEXy6ZwM3jbN1FjiDTPpBOb8L/VhP+lVsXFHbjgq7BC8VAxcGBkNHQJPYJbxiYFusOOOXh3CzudF
0DkhJ5vDfuOtsa3H+rcHm6QVaF/2FDpCPNNi4q6mMmC6HIQAl0Sdy0VazURUqxjQ0/vqaRtBhea7
VWgJC2mjs78pBR2W2+7yJjwjXm/JOh3P2dp4JQI2moieRx5nFV8tZYQZZtRhnR31Y4ibMCjOaQhd
RCOMyjpZE0qKARwRZ/8neHUbxiz1khHwCaFAVPBEn31y+Mw1m75AO6lZ5ITtQuaiN8HpvInx7bNc
N2o8drd2A78zXdh6Gj1XQ9hCoqPNf2c/C6Pggf64QDM8SFifmtHuWVjgEvKKlH5vUXGw8lkv39Uf
ZcOrLGd4XewXC73hvJYlO6/XgAK88f8qz30WNVoo40pt4U7cMiBexNg9Zp6+KCojgdsausrpDk5P
NAxYrUmaBjC70bh+5TDXA5QAaVuCXaZnf99gji0BekDjz75SacMR0rYUJRvYOkPiWKN/v0+WSlC9
C8KkUg1IkDBErAekIePbeREqYp2fPrWGXFyRE9oSKbsdSHG/yX8lIyBX9FCQXby7/CZX3paHOmWJ
ouGsscP4kkrcbZo005xfGJdI5fTBOZCYDZ0lwcFLTR8imXDnuvgVolPYVPDkp6OResoLZTBuei3t
USylpNn0cnIDukwNhj4xrJoq3o7QtO2TJ7HzKqjMq5ZqaBj7uAhCejuShNPsu3sTHSlL3IRhnAb1
3v/ilhSkTouTYZj3fv5cPWIqnWsdIoxEpyhs1geaaJDbr2zpHZOe1idGnUyrnmkhIwLM+3CBffKh
kUn07BUxXoIMvs9eCEKswu7TuGDNw9SAKLbkpSP04QxxgIqrUt+r/XRAbh9rZV11LK9d0R8PWPaY
Cn9XrcBBpLqonRhC3VLeh2+oHDO6uhvE+EVWmBmQnlM2X13fsFEx2HaB/QjQvg2+jHSthQB7SzLa
hjOKHW6WO00CBGUqB1TxQqbaj7556VVy3p88AmzCGJWL2CV9HBcdWqYO7mH65MMSccIfN0uIQ35S
rEMqcSCoJjIU5B3BkQ6lzsz6FuW9jGhO+V7fy0ihoQtfXvwk7IsSFQm5pQwWqzwyazXaGala9MhY
CC6dfyOG9/+OVw4p3ip2EJFDsb8J6lOcon4ohO2jjUo63sbVJ7j1lJPdG4zH+UDyv7Qro13tOc0C
1Vpj5yawkIhD7N0KxWnWtQtEEEGj7TG7urP9pNCkPBquQ477iT5e79/Is/1uBCjfkuwV4DPfkCG1
y0SpNTWKksM9AMkp6xpNruonkicXGh0GSAyXHAeCU3m4ULcSN8Oa7whqYNYgAF56MAV7hKvApZS1
blj81UFOdZTp2Oi/0C9Qi7XhjA19/h1illIzgUN8fsTB6Mvk/nXWgj45ctLjoXjJufgw3EM+Zpnk
pESt0LNqtfBCRvIjjIP4Y8wBHqRPab+bQ0aDJblfyvGZNzwJryZX6XHh0mVzSMm5GljVWorxGE2R
79L5VyluO56BlBipTksHkNVzSzAIsKYBOPWohxIvciTPXA3yKCktUDV7f/ambbV4l1A3Mh6xBFAa
8K5sFfqEmL51MH1n6fGz+bGJ2wHf6ok1WhCESaP3uh0YKV8qmyEUW5vwrUPZaxbRjkpsJpmr2LlA
hEvJ2ELdtWu0tPT/YzHBRCsT03zc8EBJdJTuCCbynGCE0SnGqksgn7oxACa9+rHZHXR8n2iu/Nof
hRovtOtEdlKv5ycpsi+M/gayN9ZpNAfgAKFTNR96gXyPDbnx04wyG+S6fM61KmBm1ChdZVwrfcU/
EHwa6QB4W2OJnIPSKCAFFq8xg2gIeLxH4Bq2aE/DrYQc5f9WOsuG+5GrWSqsJOpSuVT2tiWd57Mw
zlHFVzQ3LsQO1FNyD5+s7xmqWlhMwRo3F877zK4GLruzR7kDo5zYmA7j3FVZctVur2KqvPOpA9eO
2tkwWb7BGnXCkepO7h6oGXBvRO2cshw+RchSxJG07/1J9sCck4ExWpeeLnXZjhV7x/EjaiChX6gb
lyme19YvRJOEUDiGFb4+3JANvaSaPbgLnxOJYv/xC70AMe6zY777Nvi9QqMejBtQzjGUHd+/omyY
6QMrwLCz/VuGtATZuuTxMrR/DiZR1M29ylGaWJNOXDFuIN+X1jMM7hvtfj999NK3ECzruX9E7oTk
RH1TOP8beT4Sr4R7lwRDp75QIkTkPsJROAA2y3S6RObfI9GuVULd1PYOtIQNrPhjQrK/LO9klpfy
mPxBhiX5f1Z6KXpqxL2PRtBA+aORVsiA06j8Fyt9wGChkE3EVI1fylLGZZ99r92abPDTsZAw9XCQ
zXmVaS1oKOvW6cbr7hSdRjJCmjHL076mwao3hOdmcjaNC67P1QzVcCp+pJ49b2PyKwyQG5WnP4MK
yeAXXaYXY3BC7fpR3ci+8pPLYfv4QaeNH+f0yLaQT0nCin1oPVQrK9fSj06TsE1On+z3a1gW5QGt
qHQ+ouI8wyE/P5ta2BcCEfAnyGU2NWoQ7eiRvc+YcoXqGGRbQY7xHUgWIG6saE+46OKwWOhhllzm
kp1J8gnZtwcrzbYnK0v0uNuVHfjbqlyfvjya0NiVSqafus/hEMI7WgMW3cpFxYWPQK4zVTIfIvrY
xLnvYwvasZnZ+Z2smWGL/QbYqolvmDofPI598zYRxVhEaIUPR0TacCuxABLOBNBvVoeExMrQijoe
ll0xTy/3uxqsU101nQ6sD13ltOfqdOXrUsmxHFetdYOTGkpCP37W0snSZlWzuYwvWIYXeB7MASjK
v+rH3oi/AWRtKvu2jaJaZ5PSsWIgmEYjFDBCn46g5hKcv/p+s58iO3Pm98othPHg7N6wQCv562eB
Smwyv9s/bX4KUv32ZllL1ummfoWQ4k6JLS3/aoZWeUWnV39ZIT20+fQGE96zV8L7sH1Rpbqwj4A5
M9swP4P6WJZrHCukpVlqS6WB02q//kUfrhHXS9+0I0QYrRFpw/vmxg1zBVVdez1mFUW8XQfbVFcb
ID7z2BQ1aoNiR8YaEgMwnVzCE1S28zDf97aIOUULzsA4uMYFlBgPQocX6cR8vJiOba4ZfQhnyMFy
E+H/j/o9z7JB0Z4MMaFTebvQsJIcAe/KWhKD1rbx3l2jBnJgqXlUtIkxFfIZ9ccon4JUkW7YnA/3
qJpIDitU6QBXNQ9nFM3HtPYnazP6Q1oJVQcH+osM/lfPEIZa0PeAim3IZUSXkeM3UiH2ni2kZ/Hh
Go0BeSW7y7xm62EzaMopUZGL3vYoZ2giUQPdHGG4r7cJSu40gr/0RcUaujRC7EkXHxOmoK6ErCJ7
HzoOVN+Kc1oqgUUlEDy8B/kzonlkkhAOh3j2gbUzWads+KbfuZUoxnOVwycoN7s1rF2itSOM+IDr
gs9nCyIX7bXfrx3Bjh7ysyYgS2Z2dA3H7aHJYqi1AfYRKxczOL5y0KJQuU/55cGrtoB9N2f27krc
DnYgazC00I0YOCYf/9ZNbvR4Nt98PFdFzcItS+1MTu6z1nLZvDjI+n04MVSNExQL/jaekVMAyyRx
kvSM3HsEpEP4jWiWnARm6hZ3TcISWMPj+nUWKIAqjHRVqONXyHWGL8Y/kwCEKRaBOrZ5cvTAjdPT
fyRY2hHCuQKq5s0X+9LnXpdemLZIsmoVzPNApWRLwit1EZcnKayKx3TM883AEDKfbR1lE92fb9Qw
nCi7tV3X0Aja2cpOREcoTeHw3aXqf+Vxb6UOTVZj9lIK5zD1GbWzt4o458RU0iSnk9DTq9xPieSL
zKlSqeB2b+e/okVo9vn9QLoS6HMSThWWLnPgq2+/PF3+PVsBTR5fyfiC5ghsuKInPrS5rqmTEEMH
DhN72GMM/VlPRPafdf7efiB7ZVF0s9IYMZBmh+oMjkVMcXjSk4U38GBi7rdxZni4nzPVKOjJpgYb
+XX0hs4LbqnlnqV9zYvdP3no94jT5/DTexPCRnueDsQKfdCf/W+QNUiFdy4FwwAlfUpypVDrBl8a
eU+mve7ghjPmVJIeRnbC2r51lTmX/K0veztJVQGJibF8XfQ/j8KPseWrK3NiDypqOZiaMBftfMj/
3UXJMF5gl0Oq4hsLRNCIvTgGpWI67l75WywQ9zpcId9JCn1GMho6MJEQuF+9/a0DbVWT21E+bG2V
g5CYjEcDTN05kW1dzq9ZW9Iq8/zJy8FiItO3FP+axrCV3HtdAGecbaAmY0Cuhreawig6YQtqAVNg
/AByTdyBbvuO0+e6yt7Dg36s/ZESe2uRARABOPsT+jVGBlcCYmeVL25DJiBLCF4JgdVPXqrg2anX
EdCQBk0DzTUwmggtmOAuEj4wJAbrgD44i8N08xyIHW5GHzM9Hp0U6SlGrzcy2zdPvhMonreJSmRH
grvgRVDgU+/t7Bnp+80mgAv6MJDzlQoqHQLp/Ir8D6hIDs599pWZrztrGYiusQxX37We2kPY1ryo
Wsa+Wc68zwbWBs4QRLSBOQAG0vDt/NZLQ4gK0IK2tianfvi4V+jygXYOmSIndlmIOPnfuY3fBacv
4jBXdylmrnAAAIKlRgjudgCuYHQ983//qQ3lH3UgzdgQsrxTvQOqeU7HSpWZNgoF8/gqxkh++2Ue
++Rn2egAa60OP8Jjb/8gsSOStGMWLEOb+JTIK76gZQIPyEab/Cx5hz3T/r8PDF16QdfaqkKQczQw
KlCu2KyhZECfDX+/zqz87ImEunAJ/U5tUM25KeP4zKlhGpSaq/FsJJNkmjOTdZSGemrNHjk+JsfQ
SXeDlYW7CSWOCJsC7Ak65YoWdP7QKAqgHw4iaM/mh4Sot1JCTueDILoSmpOvox+wQnmBJECgyuup
ltPjE8oYkqPw7FBmhqTumu350cwU6dJOzdAmncjMbncV3+Lqm+5s4jzKftefs+e84oa92OuOORbO
lc5XVt1ofujEPzGQljiUdRsDwblzauvNgCltr1vjz1Zli/MDyKteHDcn6UtXHOVvA7k57InHkzmV
z5qmahNBo2AewaMEps5FgcQzMVjGa/sLo6TNjIaXlHcsnMeLt7k644aQ1aCITHHhOv3nZv/93jE7
WzOXBbi/crjADHC/I5wBbwA8nhGtJuZjjtjLgJYM3y52enkV6cKjHKSTf/I8LzccriOglrL+xHxf
g53NnlTyJbHqPppRpZKmn6YUxpDcJ2e6BQ8tripggIeTAgxv77TgFv3td1C+W6aqMPV6R7iJZMZJ
eEy17lvR1tZYc2P/6qrN1LAtcwm5sZkcLkJ6l/zlyFHnGDD9J2RgAw1OGLnw6n51ypj8VQdH2HDC
iUZu0nl4uSCR15MBs6DStsdvvkwXoSrTRNHNu6yjnsRij7z8DyoaXlwntT9Yoyi1IKpTcmoVo1k3
/aWdVJFSeMNOmfw44RgKLYQFUbe/5u2y/f6msIzZUeEAwihzeBe65LYHKi/VyZ+Du00TTi7uUk4T
cwxTC2upDnDeCIL4ZbQeNVvJxgaFsEeULkHdJGLd2TpWI2niFRQfOfwAFin0gBl2vUjok3HYmXZb
x/GPDWDDNdJz9yC9eCwzcFbpFT66ASMgPxyBwNl9E0pabq1hIDd4gQ+vAzemKEEOzLhB0vMzgpyk
CNF210BUCh8EzoMR74g26WecEuNfSBwhsTcsDeXh82+/az+8rmQsYulbkLwMLMSBVMcEfP06J/vu
ZPYqZZxmaHJZ5HKUHO6G80bcKkLT1Az7SrKPoB1zCfkLiKx2ocneNb+VzAccqiKCzu+/y4I66TNZ
dTkESZnB/bkFUlFhcfRH9cBtI+TSO8ZxRivmQOnQ2I8m9Yx+f9S8/enhjtTLpA3rZz/g/uky6AdX
sGqw1WKkyrZmJQXiNKNFSUX0OrPnCyrx01ljr5KyU+3jcdZy/LWtsWPgGr1TEpXafQD3l7iXqJ8M
rLJq7iWj4l2NSI3aXT4uATNIBLQ7OzCGEYYWJS8dLq61Cd6XWkX5UblQ5Z4lN18D+c0DrGM/Rt+Y
4QUrBtCjLtTUNMeKxNDCChqghAbvusZG8Cc9tGfESkFA518kbNwjaSwMYjDF/YYVOyP7NX6ujxNS
sCz9y/5x18BTGeXf7BD0uqtyOTYxt5+eXxmBNnPOkTEkd/5glbcqm6YsAqCBtCK3i9MCSlwCQfBE
REnU7LzN/tlUioWrfwmrbD1wG4MJIJrOfhIckxLrOAlVeiracMGdLvESwkp36blTkFyZjeX2yOLj
9/nKNfN39dggrNqL+LoF6T2NpaQHdHRLwe6SMt/qejE2RaV87wb0DATFXNwEH/DERBl1y/TJpUlo
U22f7OFe8R2+X90IgBjlOm1GsHKuvxf9rHq94gN09dxz+Oxx6hmQb3JJ9+cHBXgsQDCYG3uvUERm
0FR56TY9GUwjBeH/24DrjVTg8am1wkn/6U6OtnfxCio8vAETeNlypIdZ7hP/GULPD3g7odhtRXSH
YKp2FSHF7iv9efqhIXCyLbP8FdtLO/Iwu/uAA3CDqEvhqzWTdhQHuSs+0hsuNXeA2CUDLVidt8Xo
kBXK4XJVG707STDzlCYJlNvQmAcBqlXqB8BqCPh7Pvdoei4HLhOyrMc2zgi7iDWvG4+7DLlBIVg1
8FlBm76HiMloQFkFQh6XmKkUwdPpTiMVziiknFe5bgjjTHnNcs7wazqeito7mSnusEAVc8ciJqHI
7wMsw1Dak9bxLwPW2qm2wdIoByw/Is+0VDJQgt3knpSMN/OaMd/mf9QvC9mBWabZiydFviHQrXR9
wUj5g4/K8JGMgMmCLkxBUU/V8yKQu3oq4Z+JzyzdSZIWB/dlG1qqVB+9PN7vMSerdsC/X7N38pXr
JC07ynkMDJScKENrzyBrifbmU6G0Zw5AUSBygfdQsO2VZxzoPQaFKWcGfu+fveLLaInLYXRZvcVA
6lzPNNpTU2aS9ZmYvxnAmrBPydELxUkABsMIn04g6RI2KCHs4RxRnMrhseRq0/RICtvPkL597302
CyMEUZOcVAzrBHPVls7VRYDg+6Dv7Nm6UoKJ0j69TvuMB7vg8Z4viftvTg7Dn170jYYz39usB3Cz
eBRn14MqYu2U46T5Am+N0P1oTtU1+qzpuqZuZwFwQwMgEjLyAlsas8dqII9KjICvLI9R6dEcNsQf
1BnwcS0ApkaPtX/ZN9YbeFp9oN4oa5VknHmBcWghITNWluxf2PkGsXHkj5NhcIARKvCitM2LeZlM
tDkmQqaI6ZSgt6rL2bT6IKUmL91BFGYgemvhUsN/MnrrNHc969KZ522iuEXxmsOrVEzzvzCzWUaP
VyUNDbzbgfsZZ1A5z6xFUhIo0k6T4dBf1NmWpYaRwEhNeYgWGVkKzdy0cnfl8JPumd1p9Wlbf0Tk
d8pScHnL/T0PNqHQ4DqAO13e/L8Q97CYcFJ9afxHvgdX1H0dmu6oubsYmskri3miONPPBLQLtrGa
bNwISq0bWbWsn5HC1yg0xCVpisK0GMSX7dz3+x8+9TpL0/YoyMnef6Y+CzW/9AxvlxymIIzy1fMD
38hvOA7NESrehhtjDggI6flCzLYZhVB56/tz9oBbovlUb7FWD86DXB02kc19PHeojkJLQ6lleDDh
f6S45SHnoPjhwZNDL2XtJI1mDIDLsQntVZ2JtBtYZTJHmnamBY8qnjRqvhSgnMnGfCF6YnbpVVI+
BeCWnbwVavQogvbpnw/EXksUfRfffAKy7oNwU9TOlx6FDERJ/yz2NGzr3FZ4OT/rtYdIwACUb15t
YonAWukjJ4/XRX2ownHVGuZ04VgJB11dQL4UAqvfWidWPvu+HID/muIx3WV6bJ0duu6z+eq6gOTX
GhZt2BAGOgUSZ6m2ejzCG9gOy1F+xyVvPyAXgEh38HWERm4ErHwFq4ofPlFrRm5S+dsUc57TTvUR
2ZoHeVWYY1qK5lDRPBj4U4SH5qBovnv/SO0ERfoIIPve0ag1x4EIINckAdSHuW3QSWgw9IrTr0Id
UPJZcZZ1e2aJjMmeJ0y6aCGg6LKR4KYZ8RB5NjJwGSRlZHHf62a9EL4BR7riTCQB5tanxL91IMYp
p9+6Y7fFcOq4eGJljKLmvm2JeWH46YIMJBUfAUrtQ/BhC991mJvH4VKsFl/oAiFvD6wkoa65vkjd
nw169FkVENs0/PCzHQxm/2Zm2VjcRDO0cs+AjHpG2Jh0eZCfH3WAyPxs+5bgLa/PAo6igzUn80G5
r3MlSXj33IaXK/0NSILzmrd+Vz1VQ9YLUFDhuTa6b0f4eiRPZa/WUz9ncztVedRUOxvF3wmb8pwR
fsWhy2BvVLUK/iMJbt1+XrWQYOGtr9fKVWopaiphBlS43awUJ7b9ve+yXAWw4+UYqhhFZG6yWUUV
UfjdC/5P8itFLIaDTKTcZiGOieCVNYndr8RcdgSiSpTTG71jF1AASD0LCnKXTA67ktupR1rhnPfc
f0xyMu1BMOltKPH2SrWtttLugR0v1J6ABamiUZnF5lGph1FNnn6bKKUrKEG62P2eYgv8DQ5LBMUH
P/4x6phIsn5mfwn5g47otrxIixEkBIS+fXlA0SqYi2pAh6xMJRauDcyuueNkpK8zvFCn7CDFuB9s
mo+uEvboqCSPUM/qeLNfBn8BxnRscv1nLVLhkpiWYVpW+eahaRrdRFNSANjsTqDoCX80tjIMMGQv
ck2rExO2V0KCksgYZWlbw/zQSdvCRWai9jMl5oNnjRDUdMBFchxXxuU7g2UM/wIK/2ihc6uEC+WV
jkHQQ5wFlAn0ICCbXAgWjPfWI8KrnEfkmPToFvo9+F/rQ+kpinvbAsEgyZZUEhZO5+/AHA0cyIr8
UL+eJa658mtqHHjvfT+1AgMXudfVoILvY1EYUkpHaBmCAKF3D9X9HyKR6BKL3cBkO0NPJNjHAzX7
+Wb+zJB1NDRKMCmdhWxhiDy0SNLLGCJFH+gXsr2D8CDVOxxHY5Nn9UT59Ig+mUkh4B6wssJFSsST
iF+yUAOqUc+oUmwnwoLSpY6CzCycraS4+Qxkb+qj+YztAcewBPKuYCKf64IiSbBQmHIj21McD4S5
7pI3Pe/2/RwfJDgR1EUAQv0YWtW0RZsF135xfOGATaW47NOgYL3eK8rU0A+IKv5XAdutc7Dgbnoy
XXbXYl6lu+C1sQG3Q8Rgn0Dc4p500FHEiB//x2058vQFB1P9JMMFCI1KcFBATxr2gtu8NpbUsEGW
4U4bnYiVHqFzOHt1v6xvUF79+gFWXzsxuDijowWN3+rsXqiIdA0TUD6pNDxGc0ID1FYBfhl87USz
1Ug6yl0ozxAiXlUZItRS3x17XWAsPjt++++6NG0+KDlRoDMa9GCwP7zVqTZguZG3mPBoxAKXcf8c
QGdE/p29lUG6DMrSTl7uE+PC5+S2mv/R9M1kcmgOcxJmujZGeW+MztZAQKC+IO+IWsTVnwFJgBH1
JWioJ/4AlQH48b1PCuHdqd/5MAyB0VNxTDNsYch5BGLHv6NDm9uTDnr/MIsuKe0135/wP+HaIfJQ
IMTEWc+bZmTgRQYH8ZYgNE9/Hzt/R1j9l9e+TftBO3sW7oTZsMmzHAwFyMaILq6oqpZ5Z94UDg+O
HtW4pD0dZACmUB8PWLlLTDHFUJLkkryErh06xQr+KKIZWz/nc0/1nuYtnvz+mKosz1+zI7B1WOdb
H519YC8GEfETtB841NsCqDrUUyKBDurZmQ4CaGt2BIHW4G6+SdRws+kqgrJfddkNs8n/7oLapwf4
C9lxf7l3x8Nxl+vxMv6+rC03Wrfkb+lgJWvF1+WNJ42AXIKN8CxJfIS1FqgqT+M6a7vVnwzsPdyj
tGGN+LDg7I8hwO7i9MWFzn55W8uX8ymxbme4YMz+SXZIpmATpvc4pHiuHpRvUuZeKf9g9Al7JnFk
LM6wIPmjK29U2/kwsPchvG9irshJoE4zkYJNtLBp5ruG06xNWN5BuXr6ShZB3DwMqX4WVjQLNXHt
Qmo+4/jbAwL+W6ln4EhXJ0+D8YLc6LAGBgxLwhgyplDbv7YkSIj+L6osrsItTRfc+LuZr3CSUTi9
8f2TthOLpylb1ibNnXPVd4WmuJdBrUDnEMHt55/oK/v8BD/BGMQU74lgq8k9Aw/zfzAXIqnxHseK
dhsuJVDK+ji9HmTnxVr0m7Brj3i5w8+E3Ipi3cEjoLC7XAsGhzXIXLdqK2AsNGinA+whwoNIH0VA
U3ytZ0wvQ6W+UU+FYQ0uiLeRP7PsOaETZx4mNHMbxJepUOy3yXHC7/hGCXYLdjBsyD43mVDZR00h
ZXcv6j0qTszP558mnbRsh+EbQhnldVWEuQ0NdZZNfXxMCN+PlWmMoU4liEbeHAlnJhxRTojjezkp
Jt2g/bcSQ+IBKzb2n2/lnqnx584Ma+9kUZcuA8fNVsOof5dRuoYHNhkH7+uRFK5Llfb3yWh3FdZU
ypBHiQFNzHbzniZ+UiV6w2TcGoUdhVlMq0OU16MBueCSoeAABtHPddixQT9KttpjSdxrQPyh7miZ
kNEivXmcTlSgz/qbNFAD6WhMLbQHRGzrcOxUWH0cA7fokrxh83yoUaHxrmfJUr1KqD21WlWeyNao
auKaNYzVIAWQW/dNPUKN9h4OZEVr+Xu5gE8C+SIl05GwywzkEAJZZ3GxerkL/d5+H8rO0feJQv75
BxNHWWpLbXLiWSUD1PZC4K3dqb40knCPhexoINbeiRzUvsxxosnrjKDkNCVEt8BCKb3aOkqgsos0
iLqdAjzynFYjrO3TNF0vFA8JnxExIO+xQYg3nLliXrzLuvAhrhZlI+QAHjrSQexWkwIrDBn9kEp9
fG7DvciBJi0AiB+wzOuB38a9+b9Fmn+AXwTmutS9iwmYyMzjek+4KGw8Omi62vt3M8ft60fpV1Tg
ku6NsL8zq7DbsLhwnuoIV9EcomKCfMqaCnsd3p8ZkIrX+zaGrcQXXcfDEJy4yWN4tMaxYGN39r74
1ctNYF7lXn2WhLyconhquEf5Tp14wkvxjfwV7SkmR4hvc9Z44D2eU901bPmb+HSQvFO36x4DnXE2
nL7CLiiYNNwnjIKAzQhXZI0NTKVrT0dCxr8AWrv0IPMTX2qLU+il9UJxXu5ALX9pJ9pYq6JcyX9q
PQ1P60H8Q8zoyh7JhFeQVxNs+AMsSHikJMrqxvIOcLZ52ZL1W2eQtHJ1OVtdLNFuHHfn/diUWaO6
dKlKIJRE1ngpxG3ld5vJWMY7fKdeeOUk+RlIFrDixbx38QjpVT4hehrHOT3yr5gvmz6gXc11G1hS
eJ/rDzryWFUp5W/o7TptLxE6uzeMINzARkaXzGZpw2yu4Yf6lDyHdoQYAx0UdAP7KdlvtL2e89Bg
+ScAeucnkwTYHKhc8lZH3FKYNBeT1GW0G/E3UGfNqyizWF95vrjIwIK472cdFBrzYCMFvsIGwbC1
eYQw1kZZuW+iV9FG0tlD0spAWVz75HyQeTDaBWJ18Pni4SASHb9pGGiArQfE4FKuu3je9FvLC4pa
GEPNbnHM1NO+xz+TAsFpKFTs5mLZgvbyoDjfzsWY+lTgl0gUPxb95bijiLlqxqeFXqpmWTh67yOE
WvtNqwVpQlzu/id/QOfy+k2OzrgtMhzzVmQ/3xX6rBPPdFNlMP0KJh1sxROBayatJ2nh4ne87IkU
aFU/Imb1z1zzqiEMv6TH8yc9Mi+BJahUAc8rb7mbPveUbL7n9f0jY+K++quFwKG++cSAkf2+Aucc
M1AqkxHGU0JB5kkfwdm7H6bJmrgET1yTLFsVOf8XsbzbLxvyr/SAgu+dDkU5KSIZxM1b9Nk/6wvS
DNyQGC6IV+QRTz2CAHAMB50XWVz6f3FZ5wY2izB5rCMNN0X3APy6FGFwp0QcQ/awjktWRS9+5y3t
TnrqYkbKosykTHniuVywVxu2diu1XDXlA4AiDyLvdT/0UW80bDA65ALjTh6yVn5/zZN3tmr8GsM2
rvW51Jc6lqmfXLenIExkdG4O9Ysb9AIC23C66/4SXw5PuimO7fsZkSl21zBL85F1xCQ3RjWUCNBy
0GyefLUOQkJ18d49XbpcGmORZhHK0Y5paQVliNmygPfh5vOrgg+yJkQ23oOmx6ouwZGgPRieOqSs
izqCsEkUWR4zOzKmqBjt+6HuX7oyCL/BpMrKJGYEtxQMfCjGIYrK7VGmGRLiML+SyJlH3yd0n5ay
A7nNIzmrKUcIShw5SkpoYLHEqrH0OClnC8Rwc3odOLvwnEtgpzFT4YYBdTbKTyD4l05JLcjaXZ+s
MjAap7BZOtQA8SkYvNZx8xnThmZl4w3h7ik2jpp7EIlW/PH0EqtAZ9q7KdBMr3sHC5LXh+/6BXsK
jZHyTzb9VRkPaih45lNqwDCy+JEFOXaHpcu83MogIiKUYce/A9tL6N3nFR1v8HkECX99xEatWosk
Mlh99h8QT5yqz+co/t4zCk5uQJAWlUt8OdY3s9AsTd6AxDotLXtmC4kfovqfxpzF0L6xLUfLTbHp
pLW1x6QofpSOqdlEFokb09B8N8i87oJt+R3TNctL35dXXyUwttu/yZRNdYXQozzC2wq3xmA/fmdz
5WAI6HOHSlfClSmBDI4i6M7kePj7kBSVk+aJcywrsSU8Vx5WcSSo7/Du6Cz85DXI9vGZGDKAfZS0
MA==
`protect end_protected
