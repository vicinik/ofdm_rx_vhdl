
use work.LogDualisPack.all;

architecture Rtl of CoarseAlignment is
begin	
end architecture;
