-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
e5UnfV2yRC9OtYu+rRcP8U8kgBdwF2IcNmlFhf4c94GNf34NnunIfORrhgfgULP4zfX3pA6zeSAE
eymvLxfBM9voy6IovjPNLKMabKovp308tFxrul2RWnTNrHSUStRIcjF0ZysRp8d8dBC1v0ERtmai
HoNI5z+hLYNlsytFsDktdjr2hL3V0mB3T3q8lO1tP0NEb5NMa2LA5avcJqZTqBrP/qEla97ICZ28
6DKthRJLXXDnSN438Sv6damySAqoNcyyUf1Iw8chPgyUhNgCylgWJxWfhpa3NY36ILjcCHATj1Tf
5Pr4F4wMRtrTQ+thTSiRBpSZGAM7xsRb/YwB7A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 53376)
`protect data_block
DtnDqE0q6KggoHY2h8ryuYz1EuYqBKSZqSnty7F3+M4z/VUmGka3E3VEg6dKIBfvtcKsHfBIsSzY
Atxx/i5qo16FOwb+kBmlon8oVxYFlm1G+r3++RszI3OrW4ffEs5p6wE9d3WUHo/KNlT622xkJCd9
TQPmp3LaxufOwEcKC7QXjk9QMDTuo2Z4aYLOW2SaUxkrUWLpccTxdjumuYmhxIPW7Z/8OTEVRb4b
VNK0fxIro0I+zyox/fEDYuMT9Mj3HPyiCOMbk3sb++dPO/lOzkZ8f0XsAwp0t3rp3XM02uqRckqj
5ja0TI2IyPMbbxL0TrtltIzVcHte5JjgqiEdfW1UQF3FG+sb91KXFRaSSEKFdM1CvdJauU++4iDD
/uWMFt0+KWDphtj5svZr822STYoajXGePxG5LewsvFWfGbASuY96kJKhp4uVg/cLAUdeaPM/WExG
RK58yPRsSvbOYpwI3ivjfTcOroUQvMTJ0yQIENDkDdEMqdP+wCAD1Rgyp0AX5RMPlVk0LgjMqChg
XziXa+xjuDc9unWHZZQiIJGtIGN+PNllrli9HfhZdadMLI72/s+rfDOARBSIPQDVMiL79ePPj1Bx
x760r3oumPANo7jHzp1SwgN9/2CVwJNrZBLhCCAc7HU49YrZHaPYPGuxvDIfKINT+u5gwO4KzIiw
vJZZooJP8GYFHYp3tNvjlSrVfuyz/U5oRfXmxvRCPv9NSD+4nO4leh/oMrAqWHIj94djY5s05QRe
QiCYNb17Qz9TEXhPUnnHTlvDIcJ8j09pJlYRdp3oRDG5obkQVU8DTuOw3IdLTSKQOwy1lrefGhia
7ZPVZ6ax1PJzSTU9LwfVLCIi6MIReU7IyeNIUiy0TX2ldaj6yz7fMTmnmbA2Gpk+OEKdQbQwKRXp
duxIkLb04vLTekfXlphwzKMSnUpnCE/+MHfp6HXNfSTX6umKAp1vT0gcnv/eJlvjrQl/wsJDw5UY
0ZSPzJUNkoyxTdn1bi8Telcl+p1TkWrAQ9EsKd4GiqTSG6ELbk4rCN2mmxYwGembCQvmdrb+UelM
Ax+l+A32guhJXCgSMTm+/UOE2chYYNXTieez8yRHYdQOPUOWRvsrs8S03HctwHrLGD/UNkOuNQoN
vE0c0fwJUA15w/DPSKzsDEq6oDQZpVvIT7WC+W++78/nKqzVNvqtppc6lTbV5ZcHCxNkkMjPIQs9
cG/NHzonepCYWo2LsIZmkI0wm8TIel+ormpXz7+3CR4sb02pilRztCrCr/vecpYI8SGsdnUZSd1t
jrVEvo06jWXVdWZGmLJj2OsE/s0rVbOKFCamiL7e5s11RlRJnzTLe0MQMOZ7T4hcq/ACJSicD2rS
Ugg+B/isbzrf0eUC3Dd8Gwq1wxaNSbZUyv+z9YSDlepROunCL9DAO6HcInYCKjkoSBdJ1w/SC7i9
0IsJ1BDCrPxzDBquggT2akpfbMl4KenRek/FWFOYGFS6yWMPUsHK6ip3vZUGD71w4RDKXzsLzc2U
MTG/0WkGqSSa9nRtW6d9dRMJvZjc53HKcRxIs9QGxavt5J5w/qyzlOI2l0DXd9a9AISk6wL2UPTu
HRCp0TCytW3vJtOU/aY6hf02w/sOG4EWwlKkL8VQYu+Q0iEd/rJdUzcOH70zRA6VTXxMUtTfoV52
9Kim6MyCS9rxDhr+o3aKWbluq7drV3887v3jSxMEN9L4iFkdU2qg9IH/L56MAmUjqqXic5/LImcE
iKjzTNbLoO90qqqYDKeMTE84NP2P2XrM3JSzaji9YzLRCACmEeh/WZps/8JxLDpiHsJMQ4AjIiTv
kNU7Zjjfc8wtEfIyEg2lVntYti5mzN/rUcIILO/HdvZEropxB6/ObF1Q308gX2tn7tjEJSVoiREn
ZYArATORD3z4FK6Vq+xV6Qgpvj6Zu9zrKQhYk6xBX/+sR6+GCRGzbkCduRgZL30Kvqpfz5NUK/yn
2f7+okyWVXKrorIMn1uKLfH7ZJ5XxOeX+I6SP0UkQUjZ2u32tq9MLsA7CKH0nwoLSUr3s+bR9U5J
tK2V73rlpD6DZl4Kp9+ekDV8+RTbatdZbVV5AmuQyANljITDi4bA6NkeLBVD/G1hH4bil7jISRml
6BgymhXoGtHIFkZrmQeWjloXsnx5DtEJZ8P95Yk4uLB33EVJ3h9zPDAmGOxDqcWLrKQkFUs2U/BZ
x+PJ9PvMn9Tr1PJSnfyqDOJYFTnP9Lha+quuAOUbMwxw35JMy6mI2h7h4OO/VekeUNeYbcQfyoPc
wXdS538EgScQwODwqd2flv/f40LeJkPYNa+/a62FWOzcClAcAbqQnMLpkn1GTd9ugk1SH/hz2CJQ
Rav49zHBhRLPySo5LNieQLqTwXAq5Y/xuY5hv+U+w00LXEN0w1kZV2B4JApjhZVqlSijOWf8p935
/hnwcBhF46FxKQxnmVJBBjrKLxfChPFn0gdUFYiwV9/NrIHwpQwRRcATBAmN4h3vnZ8g1OajJn0B
gR07eww7HJEhNdjO5jRotCfo6NXVMt9hKwTMO0bjrFa+R+Gn5hKFGIbr5xo5Ah0LNr7P2PuH2ZhF
JRw+0bLBtqA0d+0OwnqEf2k6c6jpxcpOvZAmnK8Mqs3o+bk5QIUHmxwTfY5sQ9OTAB446/TCIg+a
KAQiv7b6TwvYr4Me8Ti7wJDzytQ40RD8GB5cqhRYw/gAXmV2qGpkWeK8sM8VwmM300Rv0RAQPe/h
nZxXxVcTeDNuMcgRbyKT6ibkdSuU10v0slCDfK7q8NPFJHl+RoLNgb6yUM8rl/CqM/rUCezVg4Yk
xU2CtkziPcZZmEdpjWPYg5slxObKqdPJaNq2/6DIg8NiO5LKGFfGICRK5+TJHX0qB29v05J3t/BC
OP8ecR/t2tnx4B/jNh5WXfpa8MmYkji1jbw07aUvh6wus2GwRk1Vpo2aXMw+CypIHdbB0YV62Ajc
qlTaQSZBmxSfKNCYBZjdhzwsiV5c/vAsEyYsiCB24WDQCQKHGzGLes0dvRAtVbtEZKiXyqcHO7Tg
VtqIKskYf1SFIrVgZIBYHOCwN8VGjbt8aO2Xf5/42Y/MDmFaL2raWN/G1tJDqYH4VO1QJub0OWFe
IwxkrG6Fob0B7LqfNrFyJZhhj5FnZCNWFKD8ZbojJFpTM0hx7a3sZJgnLVCNdhS1Y6HgxC3XFL/q
36RZN3+Y1EYxEZ+Mx8Uva9EPqldghYRYOFbFli9uv5U/XO8n/12wXZBS1h8FlqwtWs27ssNBIKxs
QKAacxNeWv1z45PA6I4pyjvexco9NOVqg6KkHpeAdX73WY0oVqbOXaiQBDksFJN2CVYC3bhLE+nY
QAHnlb2KNyYYnEthLbM0NV7uNVC6MAFVMbhXDSujijXvv8dgcHXGhd9DJzle3z6HrCWwQn9QNlZQ
NjHX0gkE56C+Wcf6vuKsQTmEkHi9bW/VR/0JKb8O0eF0wI4iGRP5iuFgg1NSSiyI/yjFsDuttjxl
r7IEIsetYTnlK9MLecrf9booS9cpsSrjXxCTxNDYDeHyuJSFxwFCRi1V3cNQZYpdiznOdYURgCXO
Z3zpoCyOInfm9303tEJDR9K/3qTzHML34DPqoJYJR72tCOinRSK0JF5MTFUxaL+T1stz9ZJkdSS7
C1dJ7RjIY2prFxn0Vo3KwOZi2XK8Ogyh2BnpoMU9mPG3FXeplQd6Qrmosz7vVI0JpUn23m16ELVQ
niKe38VjH5iJYuTZq+QUD7QSlcfBFF17pAdn497D5gKKiKg8CtpvevFEF/61K9mfYsfOVRhNnJYB
GZ7FUx0YrAEhtCky1kQZ7Ff03sEdjbkkvvw821WHQqcA5svuUv0T0QR7dfAwonbfQTnAu6Nn22t0
1Gvz9HEBOEuPRy2AY0l+dFe6hEwdPY56XDvTmNmQwdvV/XGdO4lli6VMkEezlMM+kP8UhisT63Yn
pNNlYHdxwOyFvj3a4Cwl18abIFBHcpMCpKdJpg0xf5wqTM7Ix/HD4MYXyrNBI/tn2NxlM4pv3U1q
ynDjksKpa9P9bVDnsaVi8TL0zEoP46X0K5dYBy/hl58Ox94G5WpPP/40k6OZM+aXszIk2wSCah2a
73hDbm2NugDRLR0262BAmuT5SUa9lce2X1yGnlZwpFljWUxGgo2570faTNNawKKesJFIveUdGmcW
6nxhyW9BQ3nUBOWnvIwIkHUVG648UZV06Npr05Dw0xAff0YxrTX/Oo9qN1JglYXzxlg0sA+ojGBB
60nl9lRck/eIRWX2S8l9qcJ9FQLCRArjMD7PVk3TkzwIg6OvVlBYbo4MIRT9UC6rscAy/7heKejN
i/nVi9HJpGnyx/gLniZziLy5CMvMqADxQZSM+M3QLc1om3+lTuHpHVcvpAiceERhQb1DT5pZh0pR
BAoYRSl9vCQTn3lXobknBG+3IcHvvxAO0uiGlscFsz5ftmjjjPaBDpPfSNihvB1r7m4uBQ4ajz6I
Y+c4Apn8CMqoK1iQu8xURdLNBMWXeF9tYKcMdqx2oVccnZd+e+zyEM8Onlp1aRaox2OZt+unJp91
2JoBw7l/Y5QZDhD/xQRzg1V1VgIshjxHJqFgKjmJfymk83BninFaPycvGEwIwY6SE+EH1N+e2SXe
ySKS0oVuYeZt88esmuIGodWERaBotvg5KiqWqWbLHlGkc9W+ii6ISuiDJVZ9WcMaNMtFL9Q1v8+g
dOPPl0MQi/fN7pky670tKfctQCEGaC4ab9fr/QoM2OisGORXvEjpMVxkLTGPUhPmd/wFZ4qphhOJ
+eBxbPROuvvapMJggtyCbrZkCG8JhhTglp86lrlN7xuA9cu/jAsoPmdnPlinhWggu6yG984oHnQs
DC98t3BIMefdA1GEVeSelpOo0Ly36f5oWBK2DcCzpnXcmuVK7DUoTsMF7167lVlzjT8JDHQO7MPd
unHU7ty/VCHY0laLDTYAhXM1sJHsLC2hOJ4+nL0OUa9rFgMii+fSlTecGsF5+sEbYHevff9oiMZR
PMilzrCjsRseu7MMwTa18vYj9ey1t6Ho7T8eFAN8eeBSUC0O55JznBlHSy9owezHgLlHytGOOUEw
ckuT5Xzq/MGvis3lS9C8Ut5jrIBP3CToPrRsL51b127mm5LkLo+qDd6t0b1UjeQcu+0AHs03EQFM
b6hSlv2d6QovIcsZxhEbB3l5Jdm9dFT5rtfhrg1G3Uu+4Zz3RpIHvtDb0ttF2CHC2d8uyDDu8SgY
UrHRVvkdO4h9BoL0gV8j2CWHt8mkVIl89FMWqkbNoCQI3MR6oHfpMRiF6MwlipPp63SwLzP2D2uf
UYjL8+M10jD6HpBL60alvu+90iT3wIRHYZU0iepwqEsMP6sbSyECj+iLc+LS8PkkCSZm5kGH/LUv
iR+JxSUF0v5rnQHJb+2XMlvNnP21u4dwm72r5ewPy7PkHutJLTzggG19O08QCcnShkKDZVZ1ylpO
QARHDabOC/XG4S7cZBd/yq/7jP5+iKPHjZnCjxVZ4U9ahMVbugJbnFNVJNio+i/nR0KP/wKdA0pC
WYvMOtNHHNbcHvHqcj8M0jQSru8U2y+lf6YN351W3e+gWWXV/wGJVvw6J6YB7nnjAe9rs/a9b0Si
Q4sOcXSR+9M1Evj76wARF4OmKNfXR74HuwJBxXk4KpnfR4OCN1/mp8fq6IHrMCbkV/rUQJcnXOYy
pywIcB/QZuZHMBTkjb4AcYZYo/Cj1/JGPeubMvfAkbJeeR0DqZwJDRgYXpxLA3VQiv8AG+vLY18I
UEvvo17FIMrIpwE3Piisy325c8Ej4SHl6oCV1/AHRYKQ5liy4EQkSr6wBgAVeXN4WfDtqaYP7HMc
okk6ik4jLYmOAUCelnDQbOON8piIsx3fWMBwkjXeN/KNLJDKyo/apxjmUYs/Bvo3Xu9cjFKLTs7U
X3rIrgypEGbYydXrhyZbck5SQdP//n98GCMIftO1fuuPtN0O3w2BdFIUQke+DloCvkfzmWef4dYM
ZsFKdWQ1bUJSmSZTYbYVtRfDfK5XUDI8UZwi3i2twMcv3EjlLrblD4GLxC4IMv+GTP1FKU1CX8/C
j3SEVgZtIsugylDA4R9QKROT6v6BWqKgl2HcgpDZDzd78+AM+Q68tbSeXOQI0c6ZY7PvqIyIqeYT
zN6e6wE8gjvvKu7o+mCAqt4veepi0c2EoC1liQOBLJ1WIPZoHJyeJesVpzyshTLIcJYOiSXoMUAD
JokLwCb+vuojAM+4AtrBoMbjrXpx/Aj7Q4hqDQYzQ3nn2D2saBrjYCoFwjUrwkjS3Cizi8ujBbeS
Ipj5XFgzXs4m+vdRXjQ6yLajLvSu594g8HeZPhQT8LlTHPxrmCz78BJVSPBV8wO61dOH8Q2J7n5U
xavdZqnXBe292e8tYviDxkdq9IvF/qrTcIVlqVO7ka2ycHtJTtBo+DkFVmIom8W0zK5pjyPimINc
5eZgjqWbTTrYsNn8nyaVtwGixAuWPoxRaRDwuXcXhBBbC7kSqS9ls5PfLmdb8jDVnS5u5lTX1IsZ
Hl52F1YZ9aOJMTDroQ0jduQoWLMzAFW7qv7QT4RA6ePzt7lS2SQEQhUZ8PzGCj+XAYUq5GouHwV2
gGNEJgtMwW5TAJpNDiPqDIG/mxqih7rANKMcHsSXGnXATdkoGrk17ubcqYG/HFUStdoxbDZYjl/I
9y6i0/tW5XajLLGsmG3wPEGqoC3xP6qqWgB9lkI9Kvpb42fKcb6DDLvx9cUP2N3e25PdiogsdNYX
/+AWaDRy4zMhvKa3JZKaKRAsTVIWydYRDqpw+1+4NVRMP1y9aggqgsnnT4AulX17LBzhHwLPMrbW
YTh3AxmrxNuBmFpCNcyqbUZsZxGvV+yElHRuWSB0E/8uq3mQDbjG1gjsC376NPiARjYidHDp9WJi
zVa6Lk9MR+BexJ9RQtM6kXe/6Mfvvru51Nw/QDzT7yoYP5QNsqN0uh10cLcSmruW4RyAfu6or6xq
kjcGX7iKPe+NA1k+hyyacapu7BTmpWQCi/nl3iJT06boKup6o2i0KXP9TErcvYZit804EAW4uV6x
Wtywz1zMYt1ZxbsPNE8cFVaF342/5hHFfFa3YluD6yrP9HYc1Ngi8pqyfqk/QOxuTAPbMJpTGC5H
grGdC4oRXOxjZftGwh2VhLuSTol1CkKOY9Ba0AE1rAheLwGTR0YDuijlB64VlMDOkaDqQPKUWOdW
2Ino+WmR6CVeXKOPamVNChErKBDL3RzPQgfs3YsH1t4dkiqt9H+N1sFMDIu5Vz+KBw7xm8FXk1Sx
q2SCpvOLrvV5dKI0jjVAJ0JaVnv7D06HzTtPlOF6JOVmtcvEC0F4/0pSqFUO0uQOtmzhKyVo/UJs
oy1cBXdFqcbozV0MwLSJHRspDlxjDNE6rllqSqsUz+UmGPkO1TcFp5XUvNPtDxLfJtGLgSnue5jq
9kL4J/rCFWtV6I1JaKj/V6gLbJySaHpEHgiftorcnTslnC+rG3QYtNUDTjAcEMdDcZrScQzClfrq
zIzcVlnR6Vt2TVZPgzsbGZZQwd+H49WAhLO0t6Oh/S/CG0IVPgdVgHJzcVioGSpjknzuLqqbfNI6
CeILFKGObMtMM7Gp16+oC217lB3KKyMI7MmPA3EMpsRLXKC/daTMw6iRB87zxg/JG3T36ln9t4tx
fgwihfkV8TqSgZDHu8vrMzyjHIxb7Us13P0fUJq5BUZL6q2P2nCEltoLzce+Jve3pcRsUJC3kXYz
Quk9vvesPTGvLzfxL0t3Z/LMDOy26bD3HCGtPi/3nAQy9e+pww4IYFIP6iWUi24F8fJWcysypbaR
u+evu7LBjz4HW+gnGR0DvhvnMwoTQS9LWw76hhaM1I4yLJxgmpSmfSC0WtCx+RLwzDxL74/intcD
PMDKxlGiAh7CUl9lYEU+Wbg3H8Jwg9gNhwcJSMndu8RiD9QBJRqV/wSRlbcubczarVf77UVCvKgv
A6YRuxr89saX2yGiOXho7n8htXKktVoLwUrFXR/eiiVJXJXntoJ36Poo/Z2W046uWDf7leHlYhrh
nuxiaCm61ggSMWplOMIoG1s15SR6OjKuPQxKdcxfu4W5KTTX1fjhTIk2RlJMDI6fBUXO10qP4puJ
Wc7e9jbD2rwzJoEqdDtvuLbBaoXrpCT4rmDqCjViy9Q6bTbUnR9HB85n3DZGwme96+f3CkVoKG+/
Yn+mrsJN6AD03Aa4dL8JBvAIe3QA6cUoKA0oe/UP78SMGlNirazkwXPTtP6uNBeKZCsQKv5KdGge
G0hqBbkoKtXrmCSDOvt1WMrfn2V8ISbdhY2CFZodnZhfcQ8xWhalhA7Git5Xo6xvz3m952j84Qj9
+vlWiC9CQR9F0kSD50iHSX5LcABWqe9RiNZLFN9DPmh5b4Gzc33KbkhRcJqqGhbGicliuxHvCd55
kOqlGR2ApwKq5lD+9Q3kIipSry27NuiNEeW5iPlYMX4XTK6XLQSXN0zepWfG5wy9W33BIrjJn1Vb
xHbeJ4XKhOA7aRdWWTIkGia07KojUy1P8t9RRUaiCzyNZHx0TDf2IzNxqv8q5W57bO582WuS8Pfr
J6htXuEqS4lSeBf2uA/ySEVhj0xstf2yfv+R+qggBT6AfYfOZ2M/YEYw2KuWMUTVGhBs0LcvPEh1
KNRI/hkNDwArRKzSM1TIVS/CaYIqpxi5rjn3WRC/nbJndS7whRLGmg1E1t3fThgiGdq65gtBlTow
JEqva7qbhyQBVGt/AOIZUtrys/EtG3niZ81REqx02IBLQoUu/58HA2ukdsd5FtcOVjiK0mHDBJqV
NWUQFxMxPxQkaqBkNwM9yUADF3bTQW/+LfPynczkYUtI6uAvx2ejShVaZaud36eddNtHX74A9PNo
lNq5n/kKZeePkzCRxLbBJLoJAbaaaznM3tq6OHdWxS0PclEi9IZUeSmStSaO5PXhJ5syuvpE5iW7
6G6S08yt0ix+ZyKdUb3V0WV3ow/vuGJlkYsX5Po4WmeLCPotQGPdDvYMCzafi5DTOnJQvcZQDxQU
tcsHMQbXLMkYXnXQLj9aTCzBe4Znnc/tYZ0WF0EOCypz79ElQcuFz2McQt188AU4zqGDdNklj8Eo
LS0GSc8Rp51cbvQEXCtHVpuo0/nOrdROpeBMiH8TwQLMdk4nZczg34tPwBGKjRjh4a1e9XdmeH76
fx0vzXGugN+t8JHlEVLMXlcrXy7JoBFLKYdGv/iv16K2s+cxFEcuEyujSKtn9zXTth1XDV7PXcMy
4xmAPCybqkk8YrwP0Qgngih/Tq6OqGNjFL4by3T3P4lH6DuECPoWSPMUu7yN9bPhFnAsbH3g2xQE
U3LF18I/ng199alSYCp39OWkWNKk47lk7P3DsWK4aR8i04592C8iuBnlO3ApVbgW7ksh4gSz4Jdy
ZNuAel7u/c7ZK2qzCjywPFmyx+WZFvPtF52EGPfcpsNEAblXvo7M3pyKf+ytDeXaUncXNuzOgHJH
pi9/yB2XEHHHyRVb3khf7EEK2sSF4z6vUk5N8r5BSaLF/+FTNZqXN4KLriLqn7hlR7sA45aKuCP1
upkZWgwmJwc5mhkAJuCBTLLdl1cMtWPytRqMWCs5Mq+ow9juMG16vEElJcu0BbQ7Rf7m+abuvN1E
5G9lkje3vBcRdAT9j3nm/iJVrRSMtiNeoXR8mM+9quXs/g5htCYPIPTlTMWGeBmvek8AbUm40SYr
8SPijD9RD2OMJmtaXTA+4juHidMYUXBdghBakqvfjRAZ1u4tXnRJ+SLGh3D3yC8BzV2FSeSMxBGI
hEoujcs4Csz+59O7Mvdst6ej/KOlENeXHTpozUKoxyf7lz9ZmRXWv3CPXWWSUbH302F3nbyV4VIg
yaIXpjd2re6FqEVDzR6CLXuiufPqxYUmRv8e8/HVt6NkGpQl39zAGD+ZDzk3xrcPbcR/De1SI9FY
hjK0Qy0Rh90PVN4hM+GZ9TAbXy/+AdlRp+O0k+Xpa671DGa8+/KLnBW/ZTpI9f5TMwf/AH+jt7Fk
d03emPdtNbxsHh26/NQPeHaDqYyoA0tr1vSEPB7GqLKnE/wyUVW52+vaoVrx1K1JSF/sBhbDgTvF
MkzmuLDJoc+uI77RMGu70WqOuZI9IxNlb5K0rW4Qj+lmZOuK4736TLBQXE5AqjdgOtWAVow/dkdz
wOrzjSJdm/SSOnNmFMhqKla29vsrq9H6NvignY3a61pypGZnhjSL5JpltTK8UN7nhzl3u9s0R6Qn
8UqwqTI7/EzI/eeNcMZmiTgYHAsTGicGmFkzYj1CJslosk9yZwLQr4/wP7Je/VLoVDbb+93+UKk1
9YtuJJt1FgsLP74uZMEm+BFB88rBgNV4KJmwXACbx6Y4kbwkrCyoHpmChqbRTFVhTMj49kozyKC/
p02xFPKY9Rd2gmxKB7P4sY72VjwEHa2AC89+HRPM4n17FIVNmPTaGihhTukcbk0MQlBK4Xu7rB0Q
7lByT3E9Gz++AQpzVrgSDfR4zXA9oi2Q7mus/7tcFJ3GI8B4RTnpzYlZm9ZUyx9+1RCOQD3TvM2j
qaEddvqBBpgqLwhB4DfyBbQgDkHVzZqFhXXPyFd5UPwSFZG5BssikI66OtT6FA5DevC9CdjagKHs
LgS5+71WDx0i86EA6KE6Mz075grzrDmPyvUk0rMzDbZiCr+CkzCrpbh1W6kR1R/RalVL7BTXYYIf
LvGzcHQvncP7hoVCX3neb6C6RM0SIFmCXRYetLIR3X1YdrIBZoHukU1jaChsvqT3XeaEkHxe6Ya3
bfqQsETsVPzg2GOJ1Oai5TnTvMdUYWkNkdSGXCLi3WygYyxN9pXNn6nEYtTmIqgHeSZxX5lac/J8
Uonm97gFGHUrYDyqEElboxNIHb/UzS8uBvZ/LHSEiYUt469aynWvPFPLNhQVCiIrJ73o/Ti/xRA/
KRGKV/ZRcmO4ykDtjBAqa7uzR6dSCbqumvgdd09giGQNLKhh+wjZAZMqu/D6LeUwM5mLUoqezXkF
hrvJxZheBHzCDI2Ed66Y/1mlpydkQKgKJHr8TMzxj3BQcAi4Su8IEOgiYXIC22Quy6YPhtrC0L8w
GPbyPmiwOq+i5SYx+eiU5dQbt/Oqb9PnICceJnJcztxDtqHXRjf9bPZGDZHrg7fsyqHJkr5byNRk
wtctcP1OAtQPPxWQcHkzcwga4V6VNX1vOwRKJAeJw7Sey4XZy5H2tIlfWhCsJJLX5zIH6V269Tq0
eoHDx4/LhLj8T5tYMiryRZpiA8MLxz4iKqdPdnf4PbygBkSzYhDmXd972zeUoubys52Jj4dxQ+wS
4UOm7dutoGTXo7FZLa1UjYEkwGiy4tvXVXd+evP6+l6AXuWls9jKzDBZCNZkT77iXY5AwqAj7aVd
J/eN3C5NuR2f8bgoaqck41wh9rYUearcYJ1Mr51xgn96tbNGBHIYJfQVlZbnNIR4PoZxQnLk09By
7fLxo0l4Tc+iCzieE0UBzqf4M2FGgXXeO9fkRPENUPH6Zz2a1tVwc6FgCDwEeisTXQ60r1ILgKLx
tFDu4UULATfBC8NysCEEHTq6Yj306wBW6i7Les7Y0dUZwFLC/ONoHziUX17buNFufYQRy/sUbNlG
b9I/OHM0tDHNHc7TATqIA47uJq1XmDF2Bx3rOhHnzExqtWi5anDLV5IK7vsGRRM5Ecoc8U47g8Gi
vluA97fc5GbDTVxH7phFTsXxsf1P4NX9ctiCSJsPmVwjJqqyqYvKDDjoLPtIbDmg3xeKq32hmqEU
cRnXmsOzC/0e8Y8ZpIvRi/ptZtTAxJ0JQWlF7PvS5E0Sh6OF4cj6NnAi78vEBpWCmDZ+SixtUauq
Mwa60jRiRHwZL6T9x7e+5gMlIQktk6s2nYZHBqcGdtwPmTFzyglCgMpJj+DHEOLCwVb6nWVAMCUl
poPyZ75dbzRfwX68PKec5wed020/KsoQIN/Wv4bGtMOdHhdIf1cLACl1cz8vecMl8rxveeqAtuVB
qGUbpTxgsc4VgtOKo+v5+ygpNeOT82dWH1pN38Qaw6rv9BRXEAeO8R+9U6S1KKMomPPHKOzjWjP4
DCimIvXgmqDDsxCsOqlLETQyNac+tDnz3BvVg03Gn5uXrnroErEDk+VmE17iVhI8eP/ZC8zZxOEU
kvhx+9WgicT6vNF1ni3fM66xQ+DshP1Z0pvtHIesZG/ocoCai5fCvWnB/DwVZvlIngadIVniMPzV
1HbchtLN7cYdU4lk2gZer0db4oB9IHMLROo1JQO+gSz3+r9x5jmzK6+HXlIKAWesypO6lMuIuoiC
fHqtDCb2bDlmU4b8LXgW9CjpHX+l6KbAh/mNcfC8PTk1byVjIYfbLzAG+2i2s56DCRsWqg/7I0wG
5s2mt9SToLpcQdyaMU/CIl+NOf9FaYOW2k51rj14iKXaRdcSmNlM9+6/x3/IssbKfaUq8UH8T3mM
X04ixQk4GmfS1K5iacQzvQjxWqoyA3PhtKOS/dfRJNBtorwvuJ7bgXdldfRoBEIo10oxvcVVaJ+J
rAlef/B1c30se+dPFK5xyyPtBXCMMexGIuAdzopy54Y+TAOx5LSjAvgaHFS2E6nnoPov9QvgawqQ
A8++Ydub0Z1a64aIaGTsbxgdzW2Waarwy8Gdwi1kGF6Ebv7hTgDw5KMvao9Y/lrNVkOKocIoE8Rl
PhfJEwUJD6UBPoFRoybR1HLCKefUgNnyHMfeMo9h4S7tX2hF6Ub/1wHrPibnLut/SkPAHKVp4eht
aANpQLoUv9tSf7vekbdhNJ0NtTP0e/97CR2trUgahcZjLQhg3bZeSAmV3ofpvjey5KGsy1MpQDVY
zNoKSO7bzTfVT/gpYlr0e7d+CoyNn2Jt2Lezm3KYrQtLEtenFQarVfLmRXI1JoL4J14t1mrIY265
eEgmQPnpY295bq1zmeRRYfLB5OrYLgJR/uguCDU+5JWFOTqqh4SKSHDigsavhPufGIWhI2AMsOWT
5tJE09wGeAkxqZrHLk8roQ6vncSNgkoo26i8s0sEk/9PBTyU1hIzMj30lsYneOp1G79YmISJe7q0
d8yMCwcEWQpko25e7Kjb4QOo5C3un8CNKHp8U1s/sMP/hZN4pqibuRzBZbKso8KF92PWq+XXjXnY
EWNk/ACsbv1QTGyx8s4wxegbMXJkvRGz902OxVqiliWY+y8vej3Kn2saw/6WN8n8iIs7fMGLDtLA
5uiCn/l7rV3dMzg6iK5v5E3IG8gftkVD1LwUlzne4OpmDNHH8LndhCdT0PQKXNC37A8JaH98oV29
Ow/IAVMY+RMRvv+Xg2m+T7gd2agrv2qaIMwoWGi5x0e6qWNPdVpP8xNhbUL3YHox58SAUjmHNhW6
RAm1/QXeUd/CPOr3+/S61XFWFX+IflN1He+Kcxjk53kpaRg8kzxdaNk4hFAIpZrhIhOBxFd94rzO
nZTH7boSU0+bn7duzKiDWmxrtqmyjuwfA6K7ynPr/Ez8gLXzJ6S1+1MeA8Jk35brOBKSK0+F9eYu
z6IFjQ0TbwWhdX2x6B9Utl7ZGl5xGvKyiliWakW6R3imO6kyTQzjSujWSYbRjGdCfESmj0g4b33A
GkVWCaAo28QaQx+yPZpckh6B5qr/nNneyPgiIe1/7pVTtRg/RM8WSrSBEcVI9GL6pbtZ25tb28aA
hbYWmFvctZN2qwIUIpGm+UW+mMKzVuO3cPCsK9EnCpzFC3NM/5QfFCmVadDf5HMzE/atRcP+xgc0
ntGk3tNMqct+KiY0xouSjztJqe1FOpoNeO7lznTdv5zXhyRYUwTVOn9/uzo3qdWkhaHLasgyJDok
k+DMcMyXdBy2Bvf0VDWD+j98SE78YldXPFlwBqi8NlGBkhqpzwqTDkAE6Q8k3NW9IThiY072gtry
ptfJlYWxim1rHIFzkXLIC8ZOcOeVinNxuLEcVK5qyLXJQeVkJXSLYyVbJUWSFaWS2DkNiKigDiJP
h0Evpuxi2d6l1X4A4Vm/XUIBqXBrWbEoj1GGNNSiSS4YqQ4PBvGwUdaDlY+FKAUUxFX5X9JvqGzN
sWbNpV1GgUn4N3nSclBHXEJWdk06zmhroqGglNVo/U92fweOY0Dbxu2726fYW6n8Cw1J9GdfPfcw
sY0KpQNYW+60kHsKeRbmtK6y9BM4E4nnS03uGTddF578sqeofGTwTieO2XH7WJ31GzsbfeuhFcrG
UjB19vyFYdd0INbnrmVAOfLolYWfE+tXcsfAhXkedcbNRNKCEa6e8LbA5C2UrLD9OL3cvizrNJ00
0tDfhNJFFesw+fyd7wOckC1kLSU+WuIMc8ljR06TpCsCQkDOd6+KZVN7XSQVCDu9xMSBYGS4aBDN
OD1967uWjIRB9NWcma3grkj2C+2S4lBXkdMWGN9peHHM76x7Ci3sKo+JOO8JTmc5PkCjN4XC+eha
7T6vcVCid64EgkLtr8KUxWubTyyGJritj4HvJ9bvcgY9DWFbKawpKK1IK83TMlFusB3iA2zDNgLX
sXhejkb40Ft8otjma3eCUgyl0TmJAtqZcM3Y2I/NAnE8G6HUXoIMT0cNIDUSIWox73owKxHHukz8
KBlbCUKPt1KXdhwauH5BfhhQVvMKgbcJgjHGXJmq8ZwV9YjkyITUvDI+WN4aANy6QUz0kklv6iq1
Q/ElXeFOIAjx9XNs3dIu3LxMt2Ac6za/G6gG9EAhUs7Ld7dujvpYUZu8bchV5/De9wEML+hr1PYM
3d3nqGlJJz5sPq15L00Hg/4wxHoSBCohtPaiDeTDWmbtKVgEnK7Qf/TBa7djoDShfGMJ68d0nXA9
56yj9ppG7tkhZ+8zlMuw7VS9t7p7qVJX9zXzUqFMqgYw/GzVvndFCB/vY6TYk8c6imwMwiyZ4Vph
wMDGVfXrnVfnqw/oKeFPAFUIeATsal10ZWLUGWlolGiR6xPNLJ7059pq2DfbKTp/rfGWoqpxmcNn
d2kBmWuNw9evgr8urHWENbD4/AaywvK1KqQakuzRQH2BVYoRvQkEPXI5w0PjRMX3BT1fOzI7f381
MgU5xSBk/p9tPIsf9sgH/JG4I2Adl/jgJg5R9D6bjGkq8SEV61QuZrD0/CLMRc2I520whNN3c6tF
d/O9NSzo2o/2Vqb0Idofh93PE/tzNLp187ftGt2KeizU+qEW0dEGEchaHcL0mjV1d4BiV3IrSg3k
BWWfzwIGXyufGBVaQvVRf/5ZXJ2mUZ/fNB37teEUAvdUnVVGPjwLQ2hho4aErgdTxlEEVUXz99Cn
gEGjVLEx7mcXXePWPgypJNa6POrtPvWcufGVnHVMtj9a5h9QPAgnhU4OU9RDs54xEpD5hl7rLPew
qmXx6+UKWv1PcLHxAUSNLJsg5ujsm+i4VxKfsdOw3hDEkOrIUTCsBFy6GQk8E6O5xOQ+Q4EZ7rJX
u4pieQT4sggkId0taJ+g1JQg7oF1+bGU9A1+/mBQHKgI8cRponVsMsAV9mFPppf2fpaa9TZ/Wl70
E+RSNpBeUWl+zdcRmZGeOmhhTnQ5UXY0ZOAR7UGbn1XSjXKLwyeEy//1R6kGRWgLtRw+xlo/eq6c
OkqYicnRSC4ZIbLjjCjdkokWBtPozvnnV/sK/nYrnid+ecFK/xBfuR3eakhg8RkCtGi70EwH7cG7
KI1+7rLnRBbCLl9Y40SCQuRHotLW4Cjp7fC3McjAMSwmaaZ9on9rvSbQ7APWV9InNT2MS/UFenPf
SmLDLSAUq4DL/T/8ZnZydyXdxPnMpsnhBZSSDS5bn750sOZ6j4otUhQyaSnD9jXWtrNWKPDAyi1r
zWH3H/oyQNGrAft8B3WGAhFBD3SjfKoaG62SvjnFO52LL7/UhcuYGOPT9eS9O1EIXRtu9ZkDfHmS
f8oKkMV20RhvqZeyufCan9mYIosmqwtsP6srcbmHkRALDxOQV+iHEezigT+Ql1S1u/L95iqi5xCP
GhC5sL+DCaQnvwIJcyc/9pMgSvu6ycXef7r12vmlaJC454Uwe4YjaAc+QrFc3AkVAZCiIfDRvgjX
e/8jG4lx8qzVqLWUV/6y+kmpn6lCIJdxAupS1P3QzjtcqROLnq1T9+7t3QE4BCUIgmZdOnwOZ9iW
nMfuppx/BC719zTKewt6xzA77ODmkMVYrFmausISWcXQLLjMO9k2QZcW532MsJCibRWUYdMPYgqp
VUsUyiEEA1Qa6QXZqC9MPtm+AXnzj8fAv0XXcTi/rTq5uIx45wrN2BrA9FbiCIBjDrDAllmZ5yxw
2D7xinaIODm0JFrlxVkO56NB8UvbMWxv37a4KI8imorSy0bVoyByuQbTUxrD2Ny67XhHb6NLyN6T
u0vIBGsTU8agyej1/RncrkZAmqvhRo2e0xQVVLFr1FM0mq11hhkroWge5+p5Y3mxAR9hzikuWuld
MpKBuRyuQYTV3SZOpXgbScvSkxx6e32ksNbjVEpJxnHYRTJoPlueDhzaTHrfnQX6LVDi8c43Hw2Q
jnpq8k6KSmeAjdzPrqcTnn9YoahxkixQFOmSsE3JJY1piAGIcOI/K0oyU5aHJCgON7AfdJhLW170
cloaup4UtM8d5RRC+zgQboZzctVpnge74WKCzG2mNF1lROpy/AQq23HhRC/eWvSeJikOEso5QgAz
xUBnGoPD0SQYlP0WUO8J3CfoD/fxBvIKpQI4t9SbsnZ+/a9XBOgZVAI+9LM4ufoG4ZiKTT6JBTh8
oOAm2a88uszA8qBGMrt//VxLQoycpBUvg+jOXnOGA4uRq8ntgVUMN8R/xWbXWqAoe6bJa7MJzVLQ
csLIKHBqnB4d3NRqe6q216SMMQirLSRw7iJi41Cq7ztVb27W8eaFV6+t+m0ELvjHu9s1RdZpMZuq
ytH687LqDYFZvastIV2+pGCH8h6m989tOifbZJGj0YZdqzTMrtMqWGPWyIBJ1kBqMx6UMmeVldVy
aqM5FASl+UoGmGrRwmtquxi/5+ZSrBK2kXXNfeD+v7JZL38WVNCTkSFOFaAlvGSiM97WzsrsPvxb
eGrpndAe+sALyr+tA6DdmTto2HVw16Q43zhIK4QTeXmuYxUTYk3TuQtRuuhkd8cpVwYG4HAUN/2h
k0SdWOUApq2npnnCLvM7qiJ+Jad10+tis6NAb3ThKN8teuSg5PdsZEpdC3VOfiwoRo84vi5XGWmM
ek1UZvvetQsvuWKiQKdp9JWBjqdF6XwIBRP2QoowBfbLlXhlsAqgIfxDgADWUQvuoxxhqmDmF9WS
qGKq1PvD1BcdaxF0oE6PQKHHhCHLCTT6yhDsyrGKCMj/vaDryI7BFKD25/sQx0Y9t60bbwVQrryK
AY1NmeQ8szDJjXRFrU/XowFv5PNG2fI2NDTUZ1PypV5g6xjF9nupsSw+tLoFV+5YyeutH7Scwo7n
nWuZtORGPKGGHgcksNb3qWju/JfSa6O7LhlmIaeSaevMKPPfe95lX0eM+g7BZG45Tb2BQ3A5AKZY
Tq9IRkbIIBZbTvFJ9XfIWEsNfXmR7a5rfoF9tJgewvhUlnXxcyJX+MDELs714xIOU5QmDgZFtrh4
v5ShTQYKu4HLyj5v/JJfCYFgh7PmJvJHm01J21MkWduqVXO4LtE+FvcV+LnDTvQDqWmttWLHbFnT
jfEaBN/Fq+/ypCDf4CC2gRagS43vRWna6z5mdJHWLlMHPf+0NnT65FSA57tu3QoVANqd55WL7lSO
Cd42hRwOfJb15cwI2wTR0M/cRpvRZVGfX1o3tFdVz5W6wKcH+82aIz2LKyKIGdyskMrcwSgXCrDY
AANMkoFrqjlGeqXjXt/dKG9jBqWidQ8/KZ8Ko9znVgrCXaaQluWVfXyMkUL3a5yP2Ojas0Zizmku
KuGIcB3EllnCRSglLB1c8abUELn4HM0bNEa/QGzTPrB6LkUVItkBUGEJhq6CSw1ZXmuDIZUpMMcB
DlVigCJgILwcUbNhmZ0INGjsZMgJPUylnmmuaUlVV6d3c0zhh7jhOsO4nORbY/d+Fd9v26COzDVE
IbH2vteSBgenxvWecZtJ/FKrhlTiiER/kunvmhZKdJPSKJbrRVsQuWtkmiczRQcVkP1NyEEdsc8g
KSKPi617Rd7mBKRHtTR1yO3JsSyoOXJBWIpShYXYwXZfzdEcmzw9qI3tDVEvCeuayRz1mypweyI2
xFcXnBNFIXNOMPhsA19JHIiJC0a1oHAOIhBxm+yqI7hbGJU8kFVCAx5U09cARs4SZY+Qq1+Z+2yZ
Xrh199z0wkK8yu0LV9Gb41xB5SJH7vm2gN5LNZVEAeLMm2T8slcAJTeqm1Uz6uStrpapHNVLCEDR
AdMCuYxwS9QIV1tEQfQtGiN2deZ3kl4jkYIGVJgfoEb0DOTcj2yGF/7QcrA870aS8VSlsMVAkVKc
/Nt7bmCuPRWHEAz+eXxN/f8Qe0qe7LaBYc2sHjxzuetJJPtSwBw0l1oUFyQ+uvGY7i9jv3amTm+F
eIZG1QvQjj2Wq4XZ7XqMZQAXUUB4myltPNbhefeGcmNsijXkRQKp4Zer2ulX1L5oRd1f4+NWnJZj
dk+hgk+44CPdRmyTtEzwbXbe1wEL5tnM08PxdyXhqv4NfJwcs8Mts4FX22xbW6JxqwZ0xQatBYuy
JBo7lkAYCcum+ndL/APY+UBXM2AVjNcyexSE14KlT7X14VyZ63de1jVchKeXsjUmdfF1MAQCQJPU
aHS/OL9XcOU+sD+QjggKojt60DrMYGZ47hZoMz5vPVS/Cr7DkOusuvrn9glYbYzsZfdhBEb++Jji
X7NqOUgDLNRbHCi9HDfptQHEZX+TyOZNkVEYOVF5mHG7lUXIM4r+Ta1XIosJDUKV52Dc7GlKOItn
Ti8EzObXkcoYAccpEsGMP9eVmo1E6EFPNqZ0x83hTCps+pAsXUVz25lwKSnfVlgylQ5WZSpvL1DN
x4ggyV3zOkjHsJbk2RkQlPoRDh61Skb+xHxmlkt3TJx1hILFNOGPAUozCD/LZ+JrQuBSqCoENJOk
nDFxcVHKHl2Ap0Fr6XFSj3qt/cyfGwaYQDL+rgrK9Jb3ZXiZkSCU9ZTuu8SHNfqm2A+SlL3N2GDA
ZbvAqTx1l3jPVRQJdYHq7KqCc3i4XNaM+GXE+WLJSkO+Fw2hLR5QTF8pUiEemN5xpFXb3yqZzxjB
CO2/0sVSN2DJ/4dc98lGFNkBS98qzjgbn71SLhq+qtiVxfI4ah/6x1eQwRkyIfE0G1tAhY5eQ+Mg
rvGSUvNJMnSH5zQEMyzVWhB/yHfxfENoG9vAyU8QabTzEjGRaCNqyvKD5sM/scxlzN5OGmFe4Ts6
wFJCn2QJ7aUwDxVJj53EnQB7z9cZ9xKFmvi1mv7Mvqs4zNt/GiUVeYAf/nrnR1dIyk3VsK4AJXDf
CEt6LgQXzHLLEaJhuFEDI7P/Yz5gFuB+LzhuqcDtVq3NnHfuwrLkEJVuaG7CCxjQYPQ79Ou444CE
24n8MTgFrtQgcXyULHrfIMCMs7zoRFqDqN8M2IEkflnavQEnPScZIjOXiGQAFs8C6B1WfgsKa5ic
qb9dxfqBwKfDDYHiyaWKyKQDXidhIb9vdc9AWe1LpHDSrBOA9WOJ1z4ilcexOLKxG6X0Y1iU3U67
RwIaDzdkO5iJyJ/hGNiyVXjMubNBQwo+KPmakME7r1jci8OP1GRytF5mJQwbxa+LAhjBrQm6dDqx
eW4PCzZ3zGqZ2ks1aZBkZxWlBMNA7XiYuTYbjEkrC5fEBDq/CkUpvQcQqYGD/AIF/Car4KcjPOcP
RRGvGIumFBdVZ+0ZAFEGz7xSOP3Qmsq893UwvTPA+M5iME03BbEsrBdmnypk8l2D8tsSDK67xnjF
YmLITPaxjvK5lg5JuT3zNU7yWyXebmf7q3WhmwMddrNMdcEYewGepjnVl79YeVv/9+fQfVa3iUbP
83PjERU6SPZ5nWbqCoLJb5rI18UDZh/WrTmtMzbD/zWhGTb03kasCbkidbQSN5Wu3aK/NjaXbgbe
U/3YhdCmRIFnYmAwlYHNxk8I/MEss6kKmAaaaBTnQyR9bcm2c7DYbCJVLroGrleFW4lz2PHxZITC
+4r/Mu7Pn1ochAFlgoj5ZOxWVMNKk7wRRUYzIlf4kcyU1ACDwlAfBJrqJc7vHvMCaJU5Sn9ReC2H
yotLCO25pZur+jopzXyISuzzlKGNChYeU9citz/CufLujhID/BJp6yO3vY54Xe0CxLjlIBs+Av+M
YGF+X8NjIz6uNWOBs7ikFHHz7QZW6O/JmahNDrbY9Txqxiuo12pPbcF6T5EQpycAhWZ4Gr4Uul9p
gVFiznyP0tz9OJZAHHpqid1O7pybBPJ+KWwph9dqLvXNM7tF/z5B4aLqNZnbg33JMD4+FHNN+bf0
aOC86zsncDqvQLcp71+v2orAFqlMVj7d3rsSrIUN+ZQLN/hnTSXmTqwCK3aDj2tTJApLQCAi4Tqv
bjtBuZhsiGs0vk1MOJt93+px5Ikbfj3HXkRx8la+d7dicKsHrBNuGYxccNm6j3maqIQOaDgN0ptq
4DkD5UJEX6ZY4kd7/FCXmrASkziS+uvQxG/gKXXXlRmpk5dWP9c8PVd/hDXbOu3bLhc/HIyVwL5v
fULJDzp1PwE4I+tSuAnz3QaJ3K3iODL0aMp0j++wDAd96v8OEv5kuDO3Kbz7cIXoaKNPZt3QRvA3
bSHiaO+CmsN4dEDLaPH77lhi8w52eQVkrZDDMyXaJmBmzwMfvAVv/hudfeceK8DICvwxIfSlpEQF
11I3krk8nqX2T4Vlk1rAtyskfj2jkPtSO35DxoDpQqOVD8Z6ZcUFwOl0fQ6HUjYA3SfxNyolLXu6
b1IoOEquAe2Jbr1EsRRoQsTRWDfd9lKSMhDysyZVHyHRoQOHvBvzcT45hlxEqvT2Yb4jZzBrIvc3
xSHN+wrS7cVKQuxb1daMXnLUcmO0j/1h2k4BN6IgOigz+E/5bnNg2o/uRcVEwVRErdUFtA1N+DqG
WJRLnEgGj5meJMHadbp43CZhA5OR39XXlEL+OW2UpXWzsiOndrR/U0MQnnmX5nLQ5IicpIlJnJVG
NaZM1XFFJBqZakgbiaZ9gXZhruhR+zf7z47CIlAIor9YHYYu7o1EfTN2uaoePFSeZGwXm/VvTALM
bw7P9lBAZ+f9sLLT8QbqD778kboMHdJRXxTgX0z3oLntC9O8L7btj9dGLIX964ovtBVUN9kiZl5h
rpf72jfpNmYXIOGo2IGo/VftJKibiGNScSGuNl9geAREVJBOjI0NT32KXIPGfW6xJ157BN+P0g/d
ne/Bf5/OezPTz87ydRXy1lnU9bc32TWUOP+Wi9jYZ0iMZRlPudbFqeGOw5wBpl3pXlcW03sP2zd0
z8vXrIQImL8sicLRmbj3I3/hLGVyva0FQH5XV/GRmLj3WxJbLzGkof5kdYTNEyD9BCQ/cGDV6hCt
HTYAEZ+C/IuMiHgd4tcfgmLBAkyWSorf4jBQEzUbD9IdQ3QnaCKn58LNKt89wkdjWP94yxIVhDhY
3DpcyPD4XiKz8RODKtFViagAmSkTDYUU5iUT1SX4ze4m1q8Ci1i9HX6uGlGuGdNwtcGf2VaRetpI
qp5UpQsMt019GT1av4JRjvjI7uF8+szmadU85xvADQHp5J0X4bb4q2ShcJ0oBAknbW2WGDjYyKfj
C7/t12zWpLh1wUslNf6nu0q+baq29SEf4X6jAsWRO3iUUFI1fBiiDi8YxUrgBhFiVEKpicsWhJ6J
st9qlja2NY2Q0cqKVADdSNqUMbtvUJ0+dTWTLjeXo615c1RZZyfr+lWwvfPmMcKF2e7UubllItsn
QzHr9iYP1lVg8rxARI9jcIHtXQd+ZSka1HLne7Eb8WZxX5DmDrdcWcJ1Mhpvi52IfflFDmZCfI9z
nNX5NFPhcu4ThFGlBXB0j8HAEKITKEFUxoPjAZq/jRdbqIqgm5g5lzAqoP/NQ9P/ntq3h/RCkKXp
RQNEyz6iZ92f1bSEc02vZcGGnXYmZfWRfMhTuRw2ASYurlNF/COGElGnMUrAgg71zcZwnO4/0rSb
fer/647KwwdhkRIZYDUpYRH9kkPjRg59pxj+WF9dU50qbMOjlF50/nyALkUjt/sKDblV3CDzR4sk
zcQnLkMa8POOTxBWleNCoIb8b+ty8QPdAO/w+9SIYmw5vGnCA2RrPjhhygMlXemiVtpOn2roX+Xc
SG4UciTo3jkCeBLb+wtxQRE2OB/d2Weaz9givf+74wLzVH+UVmUcC7Bopor00ehv76igKkDj9gbm
QmyIDrbocRpLN+VUZycPtU2ggg8Z6SdhIpfU/zLw99DFdfY54ULPKkXlWMIrTJvZHhzT9I5WoiO0
rd3Ha7+FoUO+3P8m23Y3gbN3OQ4acLKwJyVKeInarmqaR2FhpWYg/vwiCa5ZIwcgzA2RcWfbHvYb
Ggu1O6XDhbuDEDnByCuoGnBNd4WHSPhUgdm0u4dIYgEzqNEMCtA2EZHP6LsSPeeOOTS8zDAHEk85
OMByTVO/6HvKL2UnKaWyVvGQQkRq3Dv/pnmFRs9pvK3EGr1Wv/fFJ5c62lseFFGn9pPcI7SAV7Nd
1KeFf5qKvRC7T6xZObX7btO3YbZoIRV/wpBu4OwpOFn1xOkpvpcvcpziVs++cN661fRwMrh46iO1
YVDkY9ok9XJx02s8v8v+APL08rmTTADFQOxyd7zTfSI8FPCqS6SJ4e/KkmZvU6JATWaJ6GOhaAvR
YnPJDmRF6wW6kgcQBJ8670iVIEKENtOAIPOQSXInto1YLRTBGCTDEh1OCEsFEz2TT9tPUWuey9OA
hdAdeV0EHJGrLsBxLfkeBjejDl0fBXCbHojcFT+1djh0IUB5iTV9EgSWhJRMU+kpMHIDEVha92Jg
Biwo3Asp4b/FwVGpORy24w0l+oCHtVdaKnsOw2/P6hvyHde0JXFkeTzk6/uz7WZhZz5xYB+o3ND7
AYrZmNh2y2HM7Sx+6pqA1aeKjaH6B3Csnxt8iPbC53hiygxvfsrN+PXTyqrQKghBOH6HAaEs0xFb
Elkf5xWC5FPOssz/UXfyKTxjQGb/iXqxOi/+M2Fw/QVvcaIC2pKjPe6nql8UIrmTe/fG8ZDB8Cms
bfWmy28mZ1l3EZT33Gd3GTLvm4S+oDPtLh+NDG7lzOcWcLqRVzEIDY0Op+JiZTVpsKCkO4NzfDr2
QNClZ+4hpIyKUQLRoEq6Ydlk2dutIOz/9igld6fK8hFLmlCvMGBLbhakYDT19/EY+/khTCsCzzN0
aAC+kMjIz7iDo9gy5w7BOjsE1/iX5MV+RBxwW7rfUZvppV5ocO1umOWhQp4sG5MeSfp0YnjGUxES
0jkTveLIOssaP7LQo49fGTndqwBV0ozcSf3cApWdT53PFvaLL59NRrd+c+UbiG8LfM6eNXP6P3XM
Z5S1QeRQ2G4LwHWgl2e0PAOHqHMTJaK4m0ccbVteeq3ghjD3WbI7udn5PX4Y0+PVj78tei9xZRQK
q6IXiZQX5NU/1G2iOr7atwl7ACC+7Sw206+7VUiBkDoV62vhELl6bCb3Yjp4QTWS/PWBDVuhcS9G
TQuchYfhJbYLCbOl5DzjKmKjvPbWLj+JXjnwzE/A1wjS1Z+c4jnhntvWBWVLid6ZMULSaVFyE6u6
XpQj9Pfk9zfAvCOpaG+/lAiYQftZqVZzMu95uD9KJ+KF6mk9AWx4r0SABP/nvqBap6euwrD4Sr+o
8UmoHiFbba7muQBcTKiv6tCEMkWqV9DjtYv4tddHhWFSuaO1uGahoKzMdEp2jdcOLcrxftusO4BZ
FxPvsrhdDo7KTjSKGOxgjpMfi///av1f/cTiwVmg+CycLH4jxtSrwCB9BUvzm/mtlJH/C8t1Gm/i
ll6VvYN6O7hUHTVub9713fUO6FStk2yBGqfDbnqNM9jJz+nyexf//lNLoZKw8jEHMqUWO8uu6BgY
9+rP/arRuPkQ2CAAMzGq92yp0y3TOHwV7+C5Ft6eNZKzG3ohK5/FgH3VUsVa3uRz6C0sm8ttPoK0
+1gZfZr7kxo5Bro5s7BBUyj77+WHTWTotSsztt+Mh+PDA/6Ok8jHLkiaeeddtKqwdSbIAojqgrlC
PsmdGN9HZDNAPUIaK7OUiHrAukeKOLEKAu1RFw6+xh85H8E57cZEoA1EAlhR1u7HlC69PY99QGgP
K0RBhbBrZMFkl+D4dWubAJu7h4iG+I2Vlv5Q1RREo2fTVKB08EThArHNsH1dmGJMVK/VGRJcbRck
SnFt25ba7DakLaPRYK7zO6Snh4gtD1LJZ4ZteVr72fcFHvFxTpgr1kyZLNwdww2MFIfAaQ8tuKEh
fs0FDWwaGfGk0tFP8iJg3O7Y8AU76uP3IYYMVDA9SZzKaMIeJaWFm93PCI+inejJ4Ov8wiDVpWec
ogcYjbXnV7ZA7ScWTD0rLncc2FwPcjXN4DnSWb0ZPlvW+4aB4e6pn8JhuVOlo6jvFKdpxU0JzViK
AU2v8y/Fj68WG3fiL83RINftolrIC0Fe0gn08bSLjziY85yGEUhCDJa0t9l4nJLSPJEde2BoQ9GP
zMMos/fOS7KUJ1D2BDkLDtZlU9mqHSivRZkXg08s93+hfVTuWrhVaZsfCfaukKCtFK/e/F9dzMoH
Eeypz9V0Xymkx5ZsUTkajvLrF2iO+NH8KNnrXe7fU7l7IqYk3Ug10GUxuGdfq+uVLsqzq+UKF7XZ
KX44KzOP4efJicCWiUOpKedtMI1pLuj26o6qDlc7G/p/fnyqFPemxjc+QO9c4x92FqWar0fkfCLK
IJP+giAq6Blp84qKZx+DowtkP24ge9DVI3EIuAXLV9sZhURDHh55C2iSHndtjM5UO0w/DBLaBgUh
qFqWLvPHpFx2QgSJeJ+s13XD4gN89gl9Vn9lZBLzkjqR8t7PvaWgA7P7p4ewzxqaprZEsIKiuaer
8cjriIJ0cjICYr5QJnnR9jSHE+wHG64g7RrACBP8ErJZxPl8CCtqUn0XVMHyDGqLeu/JCBs9OrP4
oAfheYlCuDE3ihXPNyJCxM6mwpQLpM1cP3CwH3h3G/ifgsJjkcWqawgxhnH5G/O7J4ye07ZBcruS
Mf3t1aThdOMqJdnXipMMkf6cgi3k0dj5sWDmsrT3MyWdWpwhRIw8ybfLCndkFvkt7i44yUD2P7//
S97BsMWKqDk2uAxyAup99Q4CDS1pHIFrN2OHRWpUfNeSEwxc6+SRIahiqoGBITTguUjt+sFtHJa6
VXeVJ8X9KYXCDMMuxWrPqrERJwaKx7/cWqjYUEm+cUABiMnNXkyrDq18Cedt/e5pSyPiBnmWKhio
8kesezypEvQ6YzBSe0NUXtPAcETsRcXr3ZMYvV2DWwtQ9X5N3Iuyor5sVlK/L9eL6Jp6bOVrBLWM
PoWWEDXb/lJK1VnISZ80MZj/K7QqiF8f5Ik2eLJrV0QAPc6IRWafr27jPDRUo94ZXunIkgVEzfao
NSXM4bqPIWaETzn/vG8EQzqYosbAVnycoqvPgrkxLsDVae28WwRBAkWSvQIuncI/5T2hrzXsNWJT
zQ4U6uVvA5OpBkNXrofZOk6z9JiKJm6ujiu37eMn1Ee/V1vryzmkBhni0lInLFWIupalyACSSCKl
rrcXaiQuf7qQK222I76WqZfMvd1pV0UtYDZdHynP9EquWZ9l5Qgbukz3kej6jeh7Pr0KltcZarg/
vHqdMMlsuItcVVjt166SIDIjrXHBdrCtwuRazu4OOIukembqKNdo/MPRc3jEkk4ZeHPGrvlZA/ay
3RyxSEcP/w5EgUueYel0xIaRZTmK/fBOorqh8lQfFx7ZghhbUm3Hkrzc0SvVyHnu7+6aocHXrhLC
Tiuy3tzQbsk8Ramho/Ny3xc+HLpSXBIxgy+13wdu59yFsOJWiMZyZvuG87hQNcPzKeAdyt7PHVwq
xDNdu9e/KTZvexujAyYcdQTnw3KpbY8phZ7tmer5wr7S1i5Qhjb9PPFTpzMJtBBhHEznKLSdVdBs
OIVj3h81XNfE00HRny/kNdwytlB0nHXpHe5KL8MOwCTMRfsLMTRa1vzZZ39myMV9QBWg3MO2cWCs
1GfKDRRSm13gAgGlcv1O2Xsp79e/rktZOWGsydtW3UOZ6JTBaONzqZEkgTg1QfCcwSWMdyv59ofB
4whwaCzhdW1+vxkAZAHHrignUEFPfsJJGg3CPiJcfZv42JBejuzfyhBsXs+ZWf2mVQ5FaEVS4oCL
qZPG+pK9AI2yy/kdnLlRZfOvfmUkogBE6Rrz4gQpKkF8avzvOt+M/gGa73jQxQlDlLa/RqRDhBpF
YFGs7GX14woGafKIcaBf0xwTmGG37RT1gkwkNrx4bRgZQrO3WbdfNKf77zGn7cphfE7Xt8HJd2MX
lIm/kuKESqCo36NzVOi/824v3Y/Q2skE8y6W529mjtlUu/1yZd896pu+nlURGYjM3kiVLQbidD4o
7ZoIwrKBwehJ99vpyxjGuD6iQtJBTOBwIL05wV2WJUsK0RpDi6xCinPv8kNSgoktCxU2PPsMKdbw
4KYN5zhpXdORo48Vh98sKo2bZ4vRJqicpOvBAWBR4qnUx9emW4omSDz44PRvpv5WvWQlzGLzKpYF
bVK82UrISfSV8MI7aDPO1SXC5JAJPQUzZHb1eYoP/w/ssL2i17oNojknpy7aPKU6bJAe0GbUHbWD
fAlUEKGilO5AzgLNhoTE7Fqr058INoQgRCWa+UT/1A+5P0GmpeUROCnmH1PN448PGYNxuKIIGzcm
nqjsuLWGDff9433VrjcMu+s/LyuduSED11yMWdVvlkpztta8USDkfMvrmfgmyyDKle5rh3ZFYqoF
45IxA6tJOMlyUuEnm0XS4Wz48hWjF8pcQluTLmObSU04uRW2/4TfGYP3TVppfiFjumTEAdtRxViX
q7mbhkhon1AduBi5aD0V0KH9Uz3tUbhUA4Hn0jAfe43HTRYm/mTidN6RAPoKi8iQ54wbbBiA1+7H
VFvLK9THJt5iI/JJeMeoE3uKivBb6iudbMM46xyAWcnpslSjtqaCHZ55F+bA8wph6Sx1BVjU0KmN
WY+UTEI+zY4yaOfEwszO9wI3vkex0sLmNatPyjKlEUyifMf9IIIZ5+xDPUafHe+9g+MOl44XB3n0
tvetSyYl8mCVDT58NHaj9HORxfriB92kZA0qGe5EQoOvDfMstaEWFxeMh+3ZHWuzrEzT2BImgdiW
exAftkrJWBANm8R3pEFLLt2BAjzF1w7WtgmSBeO03bdmJCBjn4TXA9IWJwYiO6muGCMAuMT4JuOO
D3Cw4Dp8LD3jXNC5BClIe5Umd++rJvTaQA0ev8GVEnCTFGlfvd2ulxdG1CSkkkWtUCpb8+4ciTK4
IXPV7HZjqix0hWiCn9YQuoAhryN2UomTWIPxH1jhPJIjqxyyKsiW4cq8UGpwQ7wPMW/qblKRRCC+
vI+Dm5qzUEoW/FV9SnVIEHPW8MD0i4MWZidH2OfbINDrPqdafg7uOy2xtl/hD/DamgD4+qXK3b8a
pNlHPFhicjCKNU0B8z1Wz+7RbZ52qWp1sYtCTemdPjnCTABnrMqB6aooNLlV8gaTiIWlPKDwWV9C
+xdpm6jScP2IVjlqNOJF2x+VnAq0IUWsEklfbEkUx8qRBXjoStilyBRPJD1e+S5ZFII0fEOLE03O
oN01+PM1FK6wMoY6XTBWihdi7HXfloWBNgKgQMWhs3mN3oKP5JBRaKAKvvr5T5v8rGsZl8Oh07SY
cF9xC3kF2K0pW3EVY8TclDzP/aKg7E5FcIYmGZ3Tn5T0XdsT/o0OWDjYxWkmDeOE2zTeShQ2YL1R
JMLRa32HHIf1wzg25lVv+RrfoMR9osBJd/2yRYEaM5WY9Kn1v7jeF2jyqixFFy9jv9IXVjJ3lNDW
V1Zk0A9JFt/hWc86hwCsMg4XhjIpAwoeyWsR0LXnvKvRsM3NPWX+w7aOBvyRapKqU4+uQVobysOv
lbTjZWq4MTaB5msXVlj5vQv0vIGYUGAqGV0OPxZafJhoDZ5zS6WnArn1GLYKofnpDH/58Xuc1+r2
JxM3DqFEDsgjOJPLJ5wATa5LR0ug+6jZR3SdtD7OcjLjBuCbZT9PZXmNTmgHKplQbG5pjr0cSI0O
xpyVWliVUi1j5vQet+5jhf1DPTMTG+ExZcVz4crkdUtm8F8Sk3GPU0zFAel/8VrGhGk+vRDu5YCM
6qvNXizl0Lqx1z9Ltmd4t4genkHQxHMQMcqAseZ8SZsV86fzw8FTf2czBohmqlDEC2Ui/zR01Dn/
+lBBhuh0ztMSAaSYrbFQ+P+q6oh1oR6EQyEkjrI2f40EI22RYwLPpnV5r1aNgZzVGWtONRZ5sGE7
9ph5nVsONpOWh5D0bNlEdi7xL+kjQN5hCvHXc8L6rnw9lotfG+FURKdTLlUulFYoMqR3sbkCU2BG
9dsjV8eukMs2ZlmrfupO74OBnE4c3Q1f6Yoepb0IN1U+6NUo++zwVhjSDTrIZNN20lP0+Xi/xHHf
k2s55rerkYyTrrfDY1m27TFG9QhoPiorQYFCITfXsPFCBAX4ypD4cbB127hnAyo+tnd7nRQMYDNv
vSFObd9rel6wSv2RIhFN/fT2VDVlS/9VRbFFIzRaX0NDNhcm0RYEuqr/91C8+UkQljrS3E2Sk3lb
8G3GLH5wt3BCxLlaMFZQRbaodzBRCVkYWSjslXnwemd46FCTf60yNBG0glDTtRrwsvBsToLxpuVD
akwlqGhGGR2DXsDZFABFBhEmVvb4xZY1DFlEF1+kF5ksfFQJtONwQKCZ0NgN7E1IWMZ2eoEI8ZoY
5AI4W9xP+/E0cBQ0tzJUg+8WG7XYptmcpDJKTWCGuuVTPOSR+OhShzpUr1NUipY3T87gJ9kAekLJ
Zn77Wp2mUk2krsNg5XCWNkyGByFp190BFAu0vYnJc09sbh8C1hBR8iaHV9xU13QPuU6la21UINKv
7kRp0elmgrHzdTkeFBOArgemFvYVotLpYbqbSeXbgX+OIB4tAcsYdAhf+ANbxTMU4aeorHK+Nncb
vDX7aHfgyDcpuygl3l0l92iv4Ea5d8GAMbqeCQcd3yXCYwIKQnwoLaY9jhTYqnNmNjKITIBlh5zS
PLCZCHPrFLKOrHpoasp1hAkBCnrewzKjWzAXGV5lBSEbs1Rf2ERORA9ruK+6uGhDgKsMAlH+hVrE
T8Ernc9jUlO2//tJ0zw9+lN3hv8f810oXQfT+4exY7q5GA+K01gTEIU3jvGPrXJCfpxQoEHzMBlk
UzcJGNEr7x+2N5zcPBHgKl1eszmdzKa0oD+hBUHX3O3mtd8+B1cBHbRcYZtptLOVouy4ENKpdWOK
sr7bqIFjLRu4/yforpHDJwMr7FbjQnzqaRonrDou0LSMzDovgehRqsrSWIUp40g+w1uTaoGimZE1
gT2gMbx77xbabiTBWCDJMt2S+Q9UXbpzBkHWnXyx6pGhvi/WRTvglUyqv0nVhlb9my0QOBwFg7aS
JGtqvVHKJ6GUASP9npuDNqXSAu5GeQtPxGJz7g/C5TwMCTaEaPmHK/IwxxA1ltuBwk0lo0nIMXJx
jqD0IfjI7jnBwJET6Gchtmnis7oKws88Bqx5On/RLJgCjxN0jeRZZpAcoFwojQ+ax3B7woIcOxXU
1Crl4h9WQEEYEu+wlANux/WVnr4dDgKQiooBxBAkQEGmDh9Lji/fk72qo495/dmz3GRLyv61FaUT
c6GxX1++DKHwoxUsvmPTyI1lzb/rA/CCNmikr+yDe+QZ/S+m7v4/ccdnehBc4EIgc9bzf4YCIDon
qP+lbiizBSYkvKc+behAOtp7mWrREzR/2oBRZgLFxWIBXsi33Wn4GEIJfQVQ1osT91Y9LwrOLTsE
Ndj2vQOsVhronuoXy0ajUBY6xxV9NPEaxF+6aNXPiRHNaflh24PIucnrNpoCuHfYp15FIa8fVqXz
iQY7Mm6kjIDA3mSKvnWl3TaU7ZeJWoc4GjPOtTe7QQS9ZNGf8IL2PsTza6RBNrODJHvKTOP5ktEA
/FUEYfNspRpQB5FPvKnaJ4yE9CR9PdfXTBXtfDdE/EEz80dlovpmF2yByNh/Gsv0BjqxAZu0MowB
R33uTcfLnNAYkhG1YZRj2tGj1qMh41Jp+0q59oIgyXoNXSSPJJMWygs6Ge6mico3+Z6FXJhAo6iV
8yt87mpdi8fvDVECWOpivdxe1CRciu0n7R7i8wqs8nKplVbdBseqCwVibJeUQjpAU7qHvbnHifPr
gj1IV0yTTsuS5xcXBb1FtSkqaBP8XMERrGJEUG/kVxB8OmWimXclJ1IjAGFmUBo6+OX0W0x+MPh8
l6ZUI/sgSdryZ7Jn/xFcVCDdmk6TRnKmTCBytayDMmibCduW5EdXjOto7Su/3lU31RSHlc43DSQ8
O+5nuBZXYX58pfEd02TFwAU08NHCGI0JvGiEFxWvzkX+RR+MDe7eltqW7FzEuy6ar/6kz5wdQdZj
wdkIsE4Fx3/WnNHBV8w7z9SeOh1/3B+WFtmt7vca7+SfkTYSlJfQ2poxIz7ZekPr3gRS+F6ZH2xX
f4Z6PkRb70T2p0GqxuJW1wEttArIflCsyqJpZ9yeCiMMUn7iXwE5zfuGl8OP9cr//PyEFOAMFGpH
VZ0Yk/o+jxF/xaT5oc6aj0mFPiKLJwEwwq1A/Mz+7xN5P5051ooH512+dr6XHHX9cBsh5RQSq6/z
5jlsdaJeajL2OdKnwtBno2Ha+RnXxy+8ETFspk7oXeVHFGgrmNJuWbg4SzOMpUNvqYzpriLAoxSU
MXnWK1Sp/dOSbH/jxgn4UbBoOyofqY2feuJ16l3nE6XGPmoAu8w1Esdfb4zA31Wg3Inv9tToeH9T
hxOF5ydAAeUOmYbo/jJv9c0MFMtlo0pNYBvrIwNrnR1BhGcHNhoors/txeERMDHLp5EmjF8yDYEX
KVS235vmdsELPH3nz7NsLg2rVE10f6Ci54e02GdrZjK4wVsL6UYteLf/Ag0M4c5VYwcNm0NNPeVO
RDcBgvOYEo4w0+oTBfna73vVuVPxBlIrh3CCDataRpTBu6baVwtDzWD7hjKszAZfG2Wn5qyndfhN
Hq525gyKaJuybPtQNJNCMJh2IPtfk3EUjhZkL2H8lQ1w5RQnc5Oq3fQlqn78l4twcj94cX6lEW7B
a8W81kU5CLyK8f4XFj0jCbJriCAc8YCQlE3Q+NiCo6+LDc4D4DpRGPFhbHkBccWNwWdhBskJtBYg
xV3oiX6xY7tdeYSWi/zioiyTTHbUJ723m68cYGfiWm2WYrt8lIU7gAgJo+12UM4Qzdo/ZgY6xORw
ZANe+01QtGm5jbBAE8oyV0Tw6q30qktbyD2EaUwyeVYyqjgYgXhbh/RbzfXaMU+pQzsLSW+jDlH0
RCIhnAy2ZDTnLhtrZN56pY+egtMZ2H7cxjl2laYt/u+Yrhf9b+pX+vqQ/IroFRDDxtwXbliXXJeA
N5EbINEyKg8ZYP0d2zjg0ka+V+YUHxUNp8axgVUE6jckwy+0+Ax0hpHhhMm+U0AEC6UofUtFvvlh
CcCzyU3jDBg4oOskHLUPB9tS8WlClyOJ0/47m8Q70RZ0Sjrk2pRF8uDRtgudck/VU8DF06qyeodz
lA8PNmpqYZAGejRGX3eRguLoZFDoH9ZjFyht2mIrYzwt0sTnLuHEjsk0/quj7XuAkw07Roz4OfDS
MhS/gyQqNYMirZU/8JOBlOft2/HmDTnGuqQ3Qt3tfpzm47fGX86M9PhPesPDa1XAsDu4HKXKF6Bp
Hh9IKTPrSG/lbv8OSsofo1N5dUU1mi5iD8gp/uv64At6HkJp2m++EteojI8Z8hbuupJpnIF6Qslb
0xMLTeo/kZ60SCSlaIOnuh3ewmN1OmtSug55E/t1UdABpupns0ZtPwqX1Gv+/Hk66xagnoWwF701
j8ar2hLp/z35gdK1wwDkkfh0zCFVVGXspdBFcfDO6iYRAFHZKSgaSF1MZ8DoRBJuqpChBohoqIDx
zjVD7l+u6dbVR5+5Qr7Y0X0H2DyHDJCfOwmXOKoGSEVz421hbwDsuDSnyhIUwSNyaucati39Phcu
oEKX94vw46rVlbzKdq1tUouUfVAOmzNCxW0uLKfqWM/pSs7Ntr477rbx+JIbAfCNb6/b2+e6yx23
gwIdIZL9wFTsy1xV5WsYUN77c3SvjSc846tMgby3lcotJJ2hizglVVYUNw+Z7oMxxmI9FxyY46jo
umIh4WhGnjAzInS+BIPaq51VeB3n3NsZtekocDLkf9TCJqhbaquVdiTTgn6J7LgXySY4Hev75Jl8
lSMY8z04QbTsX1ADTuTNj8unrP/lZzcAv1PxXltxhwZqvSZB1Td9+cs+tXJ/2DvOy8+oaZSuslfU
xkfFfKk3pSsiePb9FLLtXsQhJ9XlKhLc019SRSb1NLxNeAEh5Q6g3vZlU79WtuBATolTnsTva+bu
QaZZSrn6FqPXq+puo2ULHgYkTPtJkYLvE2Qfkb6lQpymKoIm8IhQEkdnjg+57lhjx80z6vrWtIEk
9hAV0IQKUh3Jxd+AnYpUWH7/n20I12476+i6yfVgAFxFQjwQ+NeQw7MvErHMaI7TrnoBWpRNZqMB
xFEHt91elVvA+YkSQsWacDAUrbsuczchiW3Ev+EGKpUOQPJfXrf2/9CVPR8veYD1ihDQxSMZdicX
Op3H760/UsU9tVVshuoMXxOaN+2u3Q2ZandqTzT/SGBwR1166+fH0vzYG8xsUqCxxLABBm87di4h
WnD+eZPPpS+4FXT6eP7yuvszZxeXDxCZmPZAPhRL3XOlyTMGdOwCkVbD2qLq6pjslQPUrEaqKcfT
sUSEmxnY+BeXhcrvY11mhcBBCtYOD545+HUa8l8zyK+dnfFIL9B/93jsu973RYOzHX1bjRRplQz/
ElqimeOUuphAtjA2RaVwjtYhAKrQus54oeSnFnAkJ3WE41yRESwINUNGoZ+5VchdmmMRm+MLr+ro
qXbZCRGTQVaNS59a966TA/x3cbuAbH0OU8yDbUclC3LtDPA0j5PGKFURTISPYAlSdO/vfbNNHYw1
RkkVZuwOihezZEmSvPQw3IyU3b9RB1Kmz/cPipgzXhJuVov+rPvqlgEgx1DopkQsDbaYFU9ztrmO
sZLWsSFR2KrZdBdJ/+egZFlxxwVNJafrtNSYIf+r4LevpstdULaQDs/be124fFwFtsMRDwlddnrZ
OJdPd1FT+rHdFLbZejQRdY1ejtFVDMC7/CJQb2CL+KB/jf6LAjNYQ5unqe0MBIfSbER63dO5qOO+
UE5THhUI4ddM8OS1xVpcbTg1sr1CFeqbcdQTrRGEbJ0V9KJqH8lcVO/V/2AtN31a9imPwX3ZM5WG
lVmbyFC9g0T3FjvLAoKZHPIjY97WCHPi4bQmOYBZgmsgjCLu/s+5xVzNp8lsKClckRv44iEsq5Qp
CUCHLsI/a6hguw+vbPSCZpFatmiY5TDSx/D8z6ALJzkj3ckKg1EAHOWvoiMzGtiR1K0lx+CeBBuB
TNF1eSiY5OcMRfyQ1SuTHrQZ/uX1874Lq4k7UGh6wHv6WLHn14ZV+r23V6GlMSWaG/Ze1FuX59Ue
NAGWb8Llv+Hj63v1UttOK7LbrMaU1+PFMOAZvS8RdwM8SwrDmP3FoqAX2sZJNVRKXiWYE2vhbBZ+
JlCGfeCPPNfl8nQMr/C3BWXaILl/9udESo5LwB+0bER1F7GdkUipTITBycWcqzak1lTwfu+6NZ6X
dOuby38gW8id1TL8wFTolP5KgZqZ3qASxKcHA1udS7mUgmcqu9Si3BDvzdeTli+2IAcl9Y7JXaCQ
5/Em65n/5WuCXmsOXCdJbMUvVw1uvTO2M9Eag1sd0pQ8dw39+m4oRsZ1YQkxv9lm/vpFcTOA1lDA
6ElMg4AK5ww1jZw0mwJ+2fzwRC6j/kXVwFUJsy+k/d/V9O+Mb2EnUGENe02bkfgr+QPHU/Gt7IXp
5SQIaodmj8ihEPDscdF/jHXHmFcvQlA1aoswUHX7jqniBoP+NAg7er7C3dRSRBQCnDCuwaWDCXmF
mTK2KJEx2ksEijMuv59Dy5DgM4Y9QJ7L+8uubTTQ8Cw7xKw8g9Kxo4LbwpN8rJBi4BG7ZUkrE8yJ
3wpqA99TwrNBEc7FL68Onez/BZm4MWrSYqQ1aG94gzddhijfp2nZgO5YYRPAk/ngNq2fFeA18TSz
mCbV0EI8tZecLxawWNomLlBWrbYggQ2P1tt3/kCybjt6cJhOKTrmVGE7UfPAtswAYisSNiGLZ0ZF
4VPDAiN2VxVS/gPcuc/MF2vqjZjbS8g8sKKnuG29ExiHVFjS15n68VPpotxb5D1aoh9inycqMdpH
0sEmt1i5fIVg5f2fCKmHjIiG0LOlXxBMcp82tvONYt5z08D0F/q/f1+Pf4Wkxv2BE6B6d4vw2iCF
kP4rExk6tB4L4KbxXfP9TGKvwvEOLoJNbO2qJS4w2C1BvoF/SLZV6K6F7n3U3babGcQXiPQvhsX4
R9GQOk/yVMwBx3PMKv36+L6vjuUibTBOam8kPRGdh4eUjMCGDlHqsdmNiBBn6UUpCmNHU7HWabPZ
RK26bMjNzl6o5eRKzI42fE0G7M2Q1lIx0RKPvm7WCas4X6GczMt09yM1+57r2yTmBdPjLSWb4J4W
N66922KxEg5NAHiDQdYbRantPoXpG2PvaEdelgPEhSd0ZDmb8ua4Ow4MQ6GqiYA7TPPtyQL+w9Jk
fBzu872GcR3OCk/xMj0PbghziA41BrkPigJ8mVwGPMlFVMxWmE2iH0sdsDwnibqg46flZO+iWLzS
OSddkuNxrcsE4XVndGH0ZXb/L8kjJXQEkWPtU4sFTqphOrwz32/xPkPDebSrgc4IRH3qjOC5x43l
b9++vo5oHtSCnXQNqVRDCPXXhZwR+IvcOn2+IZZhjG0Kz7zrmR9CKr8d/1UwPRPY3X0LJZcT5fzn
2C681Li/kt+EkhVEDafQIsFpBQ+7i/pI5qpAzck20IbBDvCogXp3NIzS1Jv3M/sL807VQ/WuZZ2i
dhX8N7eDSpfM3RIn4QeJ45xN/CA8PO03eS96OU297s2TYWvt5miAWuqdJy8sGKM7++5c0I/pjvw2
cfJ69h6JQDly1X6BeWxCqdYlBeZL7c3i5uFktrgbAGRmP5tteYypyDUelRKrC5pCmftKp9+h0r7o
6XcSBfZTjWfT2AbXvbOyN017Bxsua4Zcq0i6HkkHbjJhNg5usOELx9xSNVOuiKzrfz5o1MhqkXS6
7+ZQ4f4ETFAHtmVkGbaUaOv3bSJD4MtiVNJRVIDo7nomQK9xSiRmbyUgh/9QcUiiYh8REoP4sc4q
eTL9+MtCR3ljJ/gec+q9IFj2ixGCdZpEG0yQQjLQloWJqnCAS9sV9+FPdeFQieOeqrYHBJWiUlbw
DDDc8scadb0Tu5/GP+j53vm0IEXnhaE5An9G9LPcIhgSBNw+Vq7PA/zxU+ZYJY+nIUjUtEjI1l2W
sI/Gfyou1tUraJ0wc/Z0oNWEB6rPcqIdtqmOSa7iIK9imwN7LoNa9riBwX6lKQ8qgH2Lay5y+/G/
PBaP1LC5j7ptTVKk3TdfqIY4bUKqPD8PKgc8/Fma4f5c4wkXPvZeWSA/vThNkUeBC8X5ffHBkl9M
5VaIzrVdDN5MDufGwmoOWPBav8DTH+5s0uzlRHjx9ZmlhX2B2srpTLewdcpwhHQHt5yNW6pbcBWS
8BytsjixWFC5ELQkzVmjkb8rO7LpGYalVgZ7B7pY1ybHrcz7EWBpwd/5Qcz8QzFz127ghPVLDseT
qQdwskSSCK9z89X0XeDI5jYyYWIBLzLIt42ZSxZXi4f7hYoPA0iz1xzRW3z7O3o9UnWTlQvWMR9Q
lGCMCrOZWEnxJcZnxTCxgUhfPo6T8b8qtzhfiH4EiggUb7Z3dR7C+gM3i6qeMgawvMeOQtHtp0B/
UFHEUDsNbnJfpnyOAm+51452h5tnFFa4Wl+Uc+zC0/AYB9LJjQR/exzL9TVTzRoqykRXlCR+eGhV
aYW5PIOcnshm/tN1albJ8zPd+FLH5FxlyNdb/A1C3ufQ/+R4NyML/Mkf8+60ZvSRzc9OZD9dKB1F
6sVLYSt475xFFv6ptHFenA+R97GPH1eX0/jvUnitQRLu/hRGn2/HFUycSX/h1yrRYBEAqjnm1egY
yWrGJUYussCUmJpd4VquLCGi5GRU7hTlcA3u/WYZQcdvJwiWduzcvQn+0Qhb0e4uvag+twaeIW/F
57962By07C0zA71V6zXe/jd2fcYxCdIXZXqyw1NWVA00CZQN4lvI7iK9hTKMxk15z7p99Q/XCoB5
gVQvu3HqJNDOwACYxPIWRI4SSh1cxKLhhIX+SmZqJH7tmlww7thsToNtNJvvIGj1FXgYvErWVl5C
axp8Q5+0KU+WKsr4JUMdShW8Q2Yk4+Fak4ole0oYyusAtOT2eEEWz0PjldoS4yJN84jsFkydFYP/
m4iJv5TEeeI23X6x3zFQbeSvJEAuAkzsyr9Kl16BTVh+pjZN401WpGLdBHbir+pGyNCSjTMbujPa
63FQ0OZztRz9fGi37pCJwAysRFKtVAnyUi/SqYk5mXJevf2az8Pmc6Cq5UhEk+wUyP3sssWKo5yk
YlFz1+410DDwcebnj7MRNJItlQbP/wS5zP8+JBmaCEHKvJR8/qHGPt+agdh27WRUVT42xelzaRTW
I3gskqMhTbn9xMblv/w+k9izn6ezg21AMsui5TTw4AVelZ8lKeoF+d4aUpctatOZADbV+t/MHxoB
UliA0KUji32CQROA8aYTooe7Pss5ADb/UL7Syym03V3COi4CJlBkrg89wPQnIPsxhTwr5f6Nga9z
Ibd9e8zJMdk5aWtUW9Zw4160BsfFMKnwVxZW5UR/Sn1SI7Sr0a3y4415lKf1Cng80dAD/lBlCpym
DlfcmlRIvH4zZh+ooa4SeA9KHVrM5xQyc6It2UOldHIjN/ws6CUZ6mQ2NeEuNAYfvafzK4sLguxP
QjKlD+05diFAEFK3AGuABeaxUgTFpYG4+Sw8Yzfy6N+aDOF/D1wrl2eeV5AdBbu9cTpvbHGdkiyX
QeOmGloQYsfq3dRs0LoDlt5sLM8sxvzxNK84Sg0Eujw1bvUHNKczHCvntHXOUFaNum38Imtle8HO
72jWRLwFxsBGK8MfwNEB5/PnaEBEbdwB/Fefj8XI4c5fsk+CC+mTYb5zQLuOTlia8jKd/nLSWKnu
+flTMz9YbOQgAwFCLzo1BNX/mlDYBryaqDhLtRyE2QkYpYpoxHxynYTynV9pSkrIXcOO9pJVgqQi
CCMSW6a5oXdWJFJte6wnTd4/YvfAtdt/V25cd84qvAtyf7crB6wMTJRIB+Sb2os3MFjdegnGVtMn
Hy6uXYE9mUBjDRD0MS3SEsWBt2J19kjs2QdTFD8tV5U358fanTOpDh8lW8KPymqwZmfehCdU8vf5
Qi5p08oJ/m8Zmbw/8Kt7fm4QWG2Q8ykgx1nhOwgqT66LZUW/C61PqYDN9ex6Ly3mpuny06uDYkCs
Hkj4b44q4a5qfMSZUTjliDDuV3gb6zcqR4LfmF4ryt6HYjXPAVU1YVnub9FsmzYD84rghZiGHsJK
BLXxJOHmkLVbZx/ED8dbT4sEsnRgretnypNTJGzPglB+7L5hmLc3xAT73Lr0DXaq6QnuNONyPfUp
tvLhYwmSTBUJgCMOaLaNm5bnFx7NnjfFJgBcEBFKG8byz8gdrW8OZHXC3wikuYVbpUKsrfyz/njj
00NWSfxlyNlLiIXDVmZJ/whITM9sz71Biw+Hxi3sqyaRMe/K1s4eb4L7FahB+HMt4DjVGvlb5KO7
SwWmIEQdqZCow3zTe1Ny9DP8v1bKdHFVnl9ROsoaHj2L35XBWd6KKWk1J6A6HV3F8IZud69gwB5a
AmNLjiwcz16vy/VD4YSq3H3d159CpcpI5mzMkfxfI5gv0Gs98kZ+s+JY8tGZSGYeHB8BEv9ig3xV
2D38LHXOOeywZsaLnWkoaeb2cuoWdy+aHgNt+A0pF6m9XJug73STIPGvt5nnEm0Ce3zNXXi0aH+V
yDaT8DngTuiBpKzZ93J2KTe/fh5f0fBwZmJx4pYy6XTzm+ngVUE+MUAQ/WPS7+zb4/t0TjQY361h
0KTx8JfMAZiOBD1/d3tH9GlWDg8oWeA97ScVxruZv+Qsuzjt6yZ3O6pBRP2HJ+8ufe4h7GlOsHe6
0LtJiSiufEpZ7jJFjZvLa/RPz5a6/eQbjuhpLQ138yedm+t7aGPv9pMBx5o0xZiFXPownnlSkoU6
nxg00z2CCwngTQ91zLXOuxGSz/y7kmYFNp5Q3tQ/CTEkExvUCMWYvkEzF0YnFlLNW6mnrdnhYPTp
8Q8aH0uFJPPb2fpRR0glrAlCl5f6uXEdATH90IJB1qTuP2HHfvZ7r6b6Jjp2CFuDO7isZV/hnvx7
5y6tafPYaSODLiAXS43CAvstd6EMGo8+VrqLI/fo6RdQLqKgWw/lc+P1zs1rbXje2//A/r3D2TbI
VUaJksxnqredf1ldIeXpYs9tVmyMiQR7E7kToxt3BNR4E9jZtn/TnTzE+l9d6RiWbh4am+KJuEFu
Kwv0/6lzU+ZpQV+w5l+6tC6LE60mWQGgNlqdPdOHZ6BeTQo6B2OlRF4fKRtoPb8zacwdKBs7l2yb
ALImixsfvVuCmLBbl9zvCDRfownEa+m85mU1LRsBYpaj/SPDalj2XfuF5RDQgoUnSPbysIYoH3E3
fvvHei58gCeEV+OwrAf99DoRO2yJuaAQhhxPOPpHyiwWxkKAwvKO804VNabEYOOK9FCKbkOHqSTq
SJZ/S6bf59ZCEMLhX40U3ENSVwBsQSJRg9SD10uhuztg2IUPNhax8tuR2WPJnYJTeTNeLILdZCSQ
SrJnglkbgB7e9AOmJirv/Opx+S5W6wjnCxJE5yXsoOvyGZUWvd1SOulAXl1NA4Y6cmGLl8ya7aLh
d9d11s+y0jqedT658f3aFjyiwVOT9O+axLWIWcRDT44mD5mPJyHrhGz4UZMThdpHFQGD/AB3lXCi
PTAKBfBb6P3ZWYnj736YzwEeMF8b1hsVwX4371BD1RbANM2K5QjlDbPi2ctYuo0+5SAdM2nhJ5gO
mgnDWKpZkpamSPs9GUdaHsfPK5H0WYJlHsfwsJ8ih5BxtipGBrIjRe+rLIe6vjx7JL0QjoQNQ0Q0
SJqm7qRSd4mHghrE4x2SSd3J/Vzdcu48/FneHB0brCXcJpY8m9MNZXxNG4PYrB54HSgG8RN3UPxr
dyUX7OKlHLHEVALnX90lx2ljV6BNldv/yMmN2LKVQ758fyzwo4nBvwF2K6kFskb3cYe9On+qkkfG
MfzS1kYI2cJ7ZOuguY3TnCu1Spr+ocbPCHihDr3ds5hSUet5Oo41IsvHKcmN8rZXWwyt4bhPIOD7
qUVjQOtMz8XN8PpAkKbbVV8sUZCgS5piJr34km4QiY3OWzWyNCt2LBGWn9YdSIrgCS7zrspmn4Wd
g7aTHEkEWTAr2Nnb0d6PEpxOTVXPp4efTFKAndULYoV9GqI/7eSPGVq18uoNf1LCM2rvKnwIMNuJ
OsIGwcRcJy34Zm6xquPsjX/HMmYyKz4IpP5UawHcfZcVBybtFPsrnrLcHWoszi98j6DaBpph82DB
yM6GR9US/Kg7fuGaqAvvvOOK6NJ/kh9f83y6RmdcsrYLLHLQ/jyLpTk6jgaNfsJ99A7DGJbI/EzP
OJJ7/Vfcwv9Ckrqshe9dgLD88UYuTtwq3w3CXwsZSORSbVFfIYnuqSmJKq3ZWK3aQHnSKtaBKCP4
z6bwjaJjYZ3NXVhEnMGTNQNYrKkkkeyqTzPibNluLngj9YwfCBm0x9fe57h2S1mng/NucZntDlTR
NnIiOxQZFIfN727/26aoXWV51Fl/DPJ09UUt9yTHhe9OZFtDujJjHG2KBAYLYIyPMfvA5jzAaMCt
99calJhONbSgesuQBfZfjS2gMSjAMUJfaTcLp9jeKytBBWoTcJw98TUTBSgtD5ZIUBMY54RlOlaX
uJmMzqKgEQPiEUYM0Z+Dlz4aIgWLPcEjQ1KNtV77/Bhu4C/fgVJ42V946ThuKAySxOzsMngXT9e8
rHE/SBhM3P0xuK4VJFJ6wEU40KqVEomk8ipvjT24uqP801YI3SgSWayaGUU4o9ZiJLaLtrDEX5yk
tMX0i0iz0rUV/2ZNyMaLZqD/OqJuoLVm1Wp2XeaGuE5U6WRZnuytQKIGU2G5r5EkGJj3WGxJxUvZ
So7G4+CiKrPb8WsAg6Klax9Guzi9y367m9dqwfaT1F2A+8Mx2Y79WHh+fu/kEpq4LSjgym9WWba3
EhOlRdyH7mfDok/9hitKEnHAw41wQS8bDyTIZNgWks1naqzIL7/+kTgd6wHarzBS0YPmzT6JoPCT
RiBp6ROHLqebcz+2oxTH9Rcypy1zUh/cm/uhaDv3qlMaGCArgIeUKyg52heuwWvlN0npV1858o7l
Vsfd4qTewTkny+UAczQULxcudW1ZQxrf96Be95Epk92PJCNivguTSDnNFomxy1vVZFZ9Pvmk4kig
dR2ndnBoqRPJTwLyOZTLcGUmU4EXBZHMkoutf65Cgf2Fq+owlkp/nhYQoT+MXaIL07LPpnGlElg0
XS1kO+W0yG3ipOHSEdLecdmCLNPUPzpz9nVnR6OpMastxu9SJ+JFvgi0n7QusKZbSWdtYkWynowf
3EOxb1gLnCsfbSS9Z8teJ2hya98+LV68+pc/BD0ioAHRF8RwvPBmgwl2+EBFo6tBi38SdADEpG2D
ukYRF+0MtFYg4m3yuQs+/jjiT8hP0vIw/n5Xp78wer79uFcYJYsmx4yGR1eGAys/RRaG2p1m+X4X
4BpdEAYgU1t8n8tKMH2/vZwZQpVpnTxrfax012AnI3gffpntC8T3Z5kLTYgY0cLaoY99lToagFoB
2ZBjjuj0q5gLQtSYjwUmjNELIbdXbHYpTb2N83Q78apkGfvIxbC0Kl2Bze695Oqd9mO4ADkT/B+p
BSeDDDdkmCvJl9Uya9Ti+RsLm6n1plbw86ivcM50c4MdanyNzTkMslOSEr64K7ij7WaT/9e8ul2H
6elr4OhkUVJ9PDq9pE5UxxIknCeDOUkZ9sW0EN+2Tu/vXEtS3bpk5d/g7h2rB7ewtgtHtT2iRi61
Dxpju1aL7T2TlTB3gdyznNVvK/Vg+Ul0OJs0kbnxI5mLgMSJe1U91A8bgWjL8Kur1Xf04NEq1Exc
4ziibmW3bn5qzo37y1hIiDH/+eKLaqpe6Vws/XCf9HoNtDtqpbgzOgDdMnUaINCvUAT8Ko+kxVDX
o8xod3+kstklBXPRfk95GARuUhLW4a7makZLIqVjdFe+qEj4B0Ja1svfhJsmXwP3oskEBEQPIJIc
oVRMjkynf7tus6mwmJ06DRftRuo3uxP9Uwuu3sNpqOmOhrgXihUJW0VWSziT3xOMiEmo2jS7mlbS
RMtXxdP+fi6xMj/9xse6grRGHkSWoR0GEFAsg1WDxl6YFlcxOG/z6aTmv5BA7KIRFZalIcCaG+TC
3IIqoli3xV6NoGi0vE0+RtfKbQoqWckAaFGa2Ld2cuHPbGqArGgsGZU5jllMQG3HCQXFVOVBwpEm
erM40MN3XgWbeukqvQnPpe9kgQM52VeWldE7etTF9fnYN5PvEaOH0cvLS94EVq33LsM05wfktYX4
7JiKLo2AA5yT5dgAi9fNrfAPa7cao7TLujx0ChPHhwoN1owC2cGGvX3XeeedJanGuBZsNh3od2wa
FdN6mXkXl2j5q4zzxVQ9b3TMjZ/zS26E9XtvYdfEUQl4A+UrDHqGIicbOfgYi2HNvo9MZ7KHtscc
ouxBkTosiQ2azo+ttrGNqNBNU17xNr2jE8vXSAAjztfg9udijBAFbIWR8O7KhvKqB/1QYT02Y6BH
pgh1yH6ToCgvw/J5uV/exx1h1aus0/y8A1ZqacxL5wB2bHh1iRAXjMQdLC0LvvRWR0k9RsrzrL3l
z9T6CeFtf091LgcEdq+bvVI+qNA3lVHlKcQ4oCs7XVT5TfJRl7OeqBidpDi6MyjdFDAPOBiKAGa4
zims0On7I9v4dHVvFYE4BlorvrxC+5+ZmdLY+FAWKxXld0S7K1HdKlLLpG/KwfgffLNQ60lfH3o/
Xyg8Z3f0sr339wXopdX9EzwRyrbOPz5wBx9WBHPpwjyrYt+VmI4JPkyPqs84rKwr7SuXI/xzFLRO
HD6zJNkbYTMQOL0YnwKzu5QkryA31FSwQA4AVRIqwlKTIrv5VStA+KPS+dG5lD4Xga2n7Uddpua5
rAKdF9UnvUbqCxxTazt7flHs8zOi382PWdjbD/2eYvifGN6US4CAtWOeZir8zaduazWqXzWgPebv
3VPh7GBO6/mv5qYE4//zZgt+XbJRuuleQEwjrSmpoSxKdNHuIIiPLSMoDBhFDVNBvtfisRKkoQj2
sGNdt+/Qwqpg01BpRNVK+X5MmN2apIOkj6dQMPp7Foz20yuf3hUS2Y9/s1o3Gw/eplX8Z7WpUMnz
N9Qw2IdviAhjyyavBICGGTQCkG9Z24S3ZMkC+aj7zfd/fBwiat3gc0yuOgoc93lxNsRK2aIdLvOJ
IK9X/pJkX3jY4XIbskg8CJsjlOviFXUYgU/sO5Mj235ihib3rrwKlzQ5jd509N1PNviEdDLy/FU5
gAaIeYlxjNKewlAOwWpLXQpN66zbKK8/dHfnO7vI6YMYy0KjsxRa/hoYSaS/3RcdYrqMbAVxMslb
Nfl7PD8gBq1e/hfA/r+KMyN5Iu83lGiWL5cjXcIMhWOq9XMrTYq7wIZxP33lY+taYvC0vIr8ZpD+
UDE+jdgkhWjA0Fv6tdJd++CnyOyNYdVrBGeTGvKyLDlA0C/O1UaeFmFw2oGOoTqwm1/awy0f1M3W
DIEIB5Z9J7VLzdUbezSqw+/YoFzVMTVpHAOPX8vUy9pKbEUOmWJpqewspCZhQRkPb5ZFiHtuXu7B
YUOzlAa+MwpD9Iw693Y9Ka/DcXfe3ZSdz83xd4+W96m3XXubGiQo88GWcYPhM6lR5bFNckrzj7Kc
c253D/7lS3WZGgI41uB73IxKW+Jo0uC+n63TF1FS/2PgtHk1aEU7Wn4KrTjE29KEhrLuE1z5ZBV2
9WFG5V4tq5nvxjsQPT/o+YqwSSAOs9UmTV7dQysFbQCgzIl92VqaQTfRqP5ufow2X1H+loJ4jb85
rdHwn42H8AmC5PB3lepGpMSAqIjL7EMChFjZIwVqq0Upg2qsNkno67866wwKI0b4767upcvNHtqr
2PzQG7faT4gpwdDpSXB5fvUs1LTjL5qDfwXjftOgJbuljoOb0NdlP7CRpD0hhyiOIDaiQK1Yv/y9
Xz/eTb/hmGWm/tTh0lJy0CkW4bsUzwC3mGu6u5A12s0QyAuMgWPqd0qjvo/vgjYUYbf7bk6bV4sD
MEXumyATxaoDTHQS7qyRWw5NCb2GT1KZSS25g9eA1XJiYPER94ToNt5/iYaxtvLQW6y6Mlkul4gu
KSIpLruOTDWAS9VqBit8srjt3bF2wrlKugNlBjXkqKDuFkb9qNnvCJ+f/BNJ3rWWovrmhiUoRJaJ
R3PFnkddKmm6QIyVRIeFe6VhQaZziCzqTviwSUX4fvYgg1KR7MmB45Zqdg1n+QjJSRMy6P3Sg6OC
H2XKut0g5Pw6FSJtUT/B3BGgDtAPvYWxRawhj3ledeAItMwR7B2GHxcrSazmmy9shyX5nC/SMzfi
D9rHGvH8hXC+UNxUlIU4Hque+WRUiJ3lzWgKpWPLi+n0TG+5DIt8lNJdBpWIDtKfxmZiUdez6aK9
NSAsvqVfd/5k2Ep5kLTX+XchUVGJy7pZPumclkiFQAsSKZH91GYnlxFu1PBGVBAxQeSsVr6H8+2N
F7tsj2f+1oC69E5xeWNBrhrSPQkpTwyWWKu1PSsJjD+CDMB0woosKnviU2mqIIy0dyjS5PbI0Vwj
lTEelDLPHp7Wr0Rbg5eHpYXFw9G7Z0oOJTZ4OMzm87vfL7SZaD5ipReQoLY6geUXk3pLaRCdgBnu
CLSPqK6MLZAO1UV8BbWXXZ9SUdXV04UIFB66THfdJrPpCijrJKFPjOs+98Um9hKP1gA8DWDtotVb
h1c5Q9suvnlelQOY5cGOzql/YN/u4DttqJx55pNwPfDsNxPsFXlcwt/WWrzEdMpjtgRAM8V5HyIf
igXyHpGDobl+H4t1h9r2GBEWLDUENLOqlT+jXYKtwGNzN2SHNonxQw0iutCcmeXlBLHJ52GShzRP
V5jyFdyDwE7EiE0NbMi1F2gIfUzm2EnsCtPh6PsmwHukwbM8nAXCdHKgGF96shsGYq+sXILDj8dI
AwobHUH34IVB/2FoNRfuxMWQhL/XwLcTldEcyLFj2ubB6mQ7M5NzJnvGP2ayNzTccMaQ2+ekA9En
iQkJFvt9ulVJ0+7VqLTEi8EmVL+/PLKIbW6G0tQJhYPPfHs80XFUWv1YJQPgtNQjgnjK+KqA92IH
NL49MlkRnvWz/q92YgjRul1YLy+qbo+6aoFKKNTMbf8K2TT1+fmAVZnF0ucRQPGtTKZ9WRAF5Ozj
0yGc2u1OFd1VgLVoeRA+aOXzCVpFaqICEj4pW90XqB+33UZxf+JXcK70JQM/8PsNciiqL1pa3Uc2
JjENns//pHLTP1ncBzu0w//7LUkOCzb4xsjIS6zt4oB3Emty1YlSU9/d4+tu1pXWMwiFRFIK0qdV
ejjgrU+eYumLGd4OZm9O8mKzAZXrnBN9utT2Zp3xLJ5eMarZeqfDe7VSLF/FxEEEL4LTM+IQyb0t
YG0+SVv3uFPKwh0bP5SeLSG2dMzRQOH4eWXteP2+teDetdrZaAXr7JwXErXRUeIBM9A55Ly2X7S8
zrl1iaeI6pTX3QB0eMQPD3LSp9bf/nhB1Dzh4pWwg2yZJRKvMGn6mZPNGtugkZYX6F039t53dIfA
29tXkkFtTcyDCQCluzaTBVoBrAptyVyTpueD5Fm7j8ujzIt1WQE5AvSX9C2kuP0I4CPd6A8z1TTt
jDBfLzoxJaGlUQ7WJmowlhuNyxCm0ULttfhq8Sdd3vMznT0OiybLJUS8fG0l8c1uu+5XbdvxL0eU
JxyHCoQ/LTqehEr1M3rWeR3FKxANyESi9T0iB4ycfqNY8nDB1UPYqRW/LpEXdxCJFxNQZcdlwmQ4
Wk/3939lto26Fd/vEzUGDpsLmQpXj7eOqC7LL3B7r6GCbeGP5Wv+Fr0CAEWX9okqd24RJURHYdrh
3Qum4H1VnLPbBX+GUMqKVupbSwcj9Q/fbcNtNoxX5l8ixvhQyfcxRvx2Mljihq8G9x+Qjl4FnAeo
FpEJbANLGlsY4Tooa9pXAVVe0Pl+ukIaOMj2I04h+LE7zbRElT3jJB+46CNnLNowyQUW/XftZmVl
XstaN4a8jdJ4TvpXhWz59g8p9DCUxw6LcIf56EJcCpKvIFMoGjlma486ZY87rqA+tTZCZiM1xEJ4
rkN12ArHY25HiaFB/l24n7gHG35hus+/kIlqSyLp4W903uqi+m8FfYW2C5K5TpMBg1GTEBqFXC9N
BLM8ZAkdYlljZH752IoyGEPgZqdUDlFvQWbQbFGSC66CuAyY3kpDV7hxrSq//hsoetTiVvSFPgBO
9vexyNZ4a9Po0yTS6C0ZAd0V3M4t2dPSTaM9mpv1eUu7V2R/+kzWxgMgFjjNIFcOmjbuZpH8jBXS
PBJK4oJ/zbk1UfJp0S+a5SfTxtA4zgyoXAOffgy0aV+8u2Dgp6zp2ue4tvCAiR1hMnaWFtA1r8Hf
sLn6wGDIjFvX6uq6tY3JTUyAKiFdpj/ye1idUZ+X/HteXlHqzjpnTGZo6mq1SW8M2mCFJTq6VT/C
ASN57G9PzqfZEVmMwaRbEi/01DMW5qAkXOm/3XRipWa0rar2hueEgh/0ZHD4ZPWAHTysr0S8pOdE
pdSxT/+8N7tPnq2LMr59Fib4lTrQQTt9ViwR3O7Kq4PK40PgFrwbiuPTalFlHYD4PVMY2EGwtsWw
Hga+lFtzA3pZWWxoFHcb3ZyHqvlru9RAh8P8PGCdcNo8oy0zFg8UL9kNzIhNclvgzjDv64L06gU7
mmQZ6cuhONLx3HIQ/NuY16UZTsMS7v1W6M04nz6iYLkpYqaR+VRNgZ4MeEauE8iBYp0BK2Cc67fG
Vn54MTUHxzMuHZZyVwmAYolcEhLzaV1tFUsuPhhksnHKQBaV3+MGGL24F2REceiWyr902RLOmezI
Pn3DVc/FPDJwT0nrVlpekAYSyNlSpV23saVfI45Ii+cQxWPNEXjnnIMIaa9JGcyhd4xVDzeX9/M1
af+EliPMiLjtvNf0CWWV3QX5uIOmZqNxdAuwpS4H4DfDqIje0ZZPxgkmxz3nVYh+7j92+XGLrQfH
WDvhbX91oAijX51L+5B6iCbLzerUQIi6O1yRMw3RqR1KT8C8Ub1rLKNTMvVRAMyN7j6H6RfH+BfN
XYn8tULMRkeL6q1J7V8xbbdM5fVC3XaSHwgtq2Mb0Zj9fD/2xTMdCQvn4Q7tN2glpQHGCVoJvAyQ
GW/D1yPoreEmnKRr5sIwGA+5ueWnO1eksQtifX+qKFAz7qKbPxcMJX9qst/FmYIBRMfTmfPb6yPV
wbq7s3BLOhx/N5/LVXNswZE/1zxqoBrNHJj/H5hwSrg2SMHpzZZ0pztl9y/BfbEq1FO+qNURCxe8
WRcfq3RfNu7PZC59d1npI5l3YRDl6Dr0wF64ZSiW4EJzlYrte3nkJCe7E/zlFDaxH5USqgiDzc2m
eWSFHa3u4KuqtoBYwk31aV0Fzg9NsZQNMNmqR6eSHkuJpVlhLYFZr3JWY295uI+JwFJzeJEcMT+U
MOZw+3rduDjPv3LA2Hw6f4ohqbg8rzjcoze+qmI2p16ad2M9KAUwCwSxg7wzgBxz0XIn6KYC9kaO
sAgUkQC6z/Jf8csp5IvvrdgSist/apeEEc3uUVP43gApLJWg8QWsOmqMubhMN5wYb9reEGJsqC+p
8iJF69R+uqj3bmT4RUF7uPCPXzDInJFpN3C0Ns4oTKWSZ8AEN9L+qsmky2rmRlaYmw/vw+jeRK87
fYBzNmcLxrQIKWTzuEl0qxkK7LxrkFSwAEffqy0+GT0Hmc3UIlKcqA0Hw5C6snC71C2as/Ph1jeE
RD573xdlLNepCcuO0C6x2AflbW1Qq/hjHCpBjXow98RuVpIJ5JOKXsRy/O3VvoXWH89bOj37Er6O
zP9x5r6gNuaHNfH4BR8Q58K8K/BAwImWq2r4173ZhHMlCUiUZU2M6JIH68KEuvJpjib3LKYgXrZE
YMA2+3G6FA9xnfABH54SU2qZLyXYZYChxcBPwax2wuXZEggDrUCH+VbJUv50NV9ylk3P0N3omrlB
p5MoTtZIMzln7ove4+Dz/igOMBZvY17Z9LezId4yKygsI+YbOad6fADjYilSmKClBiF2LgHfKktt
sJssh8QzgSgzdmpXfo8dFwbZxs7zTDl7iHnWi2xMKQxL0YgxwZNyvmySyb6CYX6ipGx7717jFdNn
Q3dj+EWi484CJLyzM61T9UccAEIx9yab1kONfJL89TGe9ITX6w/6KAc9bFeT8ztnjDjjja+fUGLA
BXWDAP1gs8wEqqVhsMgxfjQFQZ5ZQ2P/haJ5+pCkbZmBJmn5SYNcNVxMKU3m+yNTIlbOPIrnGt5S
2v47XAJuklqAArv2nf7UpHB9c2Eh/bnh70o/H3xHy8IPByvsUGhxtwqWp6Kgvwu28QkQWJ9cIeVb
TRx7jiCDGrLAjOM1Z+lbE00cv7sn6Hu+BH5AfYpYiI8dPYHv8omtEVrXm8ThLaN5SqN2xv67WKyL
11VH6zuggimmdfpql2Dfv/zDKbMg846QJ7xb+6V6Uhp2w1gN51QiVhQqBQJdOznwE0ox6Lw2AOLX
5ssG27Av4MGy6Y5EdbxS/DzDAtdrX4bn9n/ufW2VyyJgggyVTxD8YGT+uiB0d3n4ihIBtnqvE0Ky
iPkr+BLDSqjm8U9BIn3QwvU1V9qWz7W3riscAgcuHcuRqtz7u27Aoeo1EiG9BqWZrtC9IbKHdCVo
V77ei957qfBUaul93c5zFi2++gAZ+kM72S1kpHvVuiK/3+jlvZcRbWjr/28vmle1hBxFIBjvN5R/
/eZ5uYz9QTS9WK2hEE3WLixK+C5t/8UlrNunttvr/X77M4rOO+i245rAMkF0cdPZ9AabPvLJrSQZ
H+t7XP24jsapIToh20Wct8NxBP7TQ/jki/qn6nVY6A+m229RlKZRiA2AfaKtvCnSnpG72lFkefdu
79elcjL4Jjli5p7Ae5LFDHhVaIrcNNszQ6gHLCrX9q32WAUEuYpefqoTZbZfSGLD5BNZ8c/2Oi+m
nDEN2uZ7qWSPKn8MulIpRBOUnBTRHDHUNjW6Dy7P4XJvlSXHN9mhCqfb0EhPnPgocroNpxT3apoa
WwDWEj5caZ16kM+0hBR+13t1bh8Di1HOOVo97UFqmDXKFbyPLkMsJ7ygJJZu/E34GHleHJMQwBwU
6GB7Bm3wJZE7kvxudj69S3jMOpBMrpPwNe3XQ0mpDgrOiO8eTOg/ragoXYLNEhrW1tEil/F0kAzn
f3o8suOh6oZ1Pq3iidFBqmtDU+pcUJLk3SC/bUjtw7Jy152jT45I4oJbW+Car3EmLYV2weAlmdrI
dTZz/nAUy7hSIfe5s84TiAdax+wHuVUUzkwcqKWuxqNk2ek5myZq+m+SKDzwrHLXOjfmwy/Ms4hU
AwoAVFe+7h33qiQB1UyYQTvgorLqoi3niefXCAg75ctv7NRMvIC+gBbMdB7IOLDAWDgW3vUVhpuw
/+68RrV3HiwqasSPmpdO5hBkdAYf87pZnzVapXVNXPfGIgZT9ZB7jwsEe466Vihtgxg73f5CZQHx
+6f9oXKc/SOGk1o9HbB3Y7iMWxJQuROnQgcYXEiziFUB6+2UTrWs/8RSp0VsXlgIaFFJmUUhHgt7
1ywyIiiVJPjt/0R4E303Gf1ETf7oMLRd0KUfqiRIK2dSlXU3EfUwp3mB/UZuDMe6eJ5lvAwf05Ux
r1vYrxxlgQWgM6bmh9LgDpP1s+hiKih07DMRPsza5QHSVR9wzBVh7KKilItP+PN4n6hTM1lPpBvC
igX194246mWSCEqcfqFq8cVMtgreN1HOYTN8hPDdEV3ISGcHdJ/iCttK2Ehk76zRI6+zXSTH3tWr
JS/18HL5pgb9kfx+f7wd6tB9KPQHJTV9iq/jUVzGvPbiXDmQgRwvMrQ4/uPRKFNsPzfkVccLoJ5A
tK+Eb0IHI3kWte+rMLo6qVHOBzdfqiyaHiY3I68arq+yhFiR2wnOCO887uxK4PWrnJuycPISq069
TrkMwSdmw5vXlOQXjnx+joRl2jViF/nF0jiSTpGDmPGuI209B/mKfIHNep4T/k4p9ud8QiWLW5yn
q2h+RPXFgytxgEVlNhNMzUWj2/+yLgecoJMPhLdIljV9F2Bx2xJQVd8YAerGdUMWO2hep79jUHsN
hzybjTpicPkc+PdhdiwA6TZmn/1n6wOxEmB74hopd4H468LgAYzDsgRjW+14T4CqZ1ngLvJOT8GN
aW5meSnkwrGFvUUQiakHE1gdPjY/Dm+nMPmkOe7Z1MP3SkNrz6Pu0dloYVcePetr84nrwjiWaEpl
gmYncZ5StGi19T7iAle43TSpjqX5ad55ZznJFS+60IB2VJ+sEGUCu5L9v0vEJD/OB1LFrA83i/Gv
GcyFV8am8MTQVkIeBH5bAnmWJhp2wtRqFS2/aLYgTo9oUZez8SZOojAWR+WZwfX+arfCKhY/Lrre
rQHWOr1Xx6GCFUjbRjiQUUDAEm55d0HLFuYDQsMKo97xjg3CVwkOetT8IG/XecueP5rfvgy8Uh+/
+rqa86ofbAV9rsXPPUB+YcBs5EqDDc2jDGqlWrXmrhOOJlIQAalGbdSdIPFVtFxzp1mA8GR0JPKy
vl9QI6+MTuBGALPDlJKWbgAszLuncHv5QN+/7/y5IQAfG6Jyro4kEYH4z8GjVOACaUETVF7FjamY
MG9vFx5RcKPFOoaEyo+ZfhtXqDIW9Tn5usHc4Gs9pAFaYCmgmxdmIv+rLdzmGRprMV8AbLNq/76d
c7RWtYTGQsV526HDBa/yvHPlvxycYEgiR+826Qcvchmg5ljoTgjJpXtADcXZI41zbvGpw4tE+0Aa
qUWg9wD0qt4/2Du1Q0ipNgKgtm96u4DaEXUyS7Cno33dxYrajEeVMujEJ6a/Hg2wIHLKAJCmIyb4
9XXAWkyhogHXXx3e4ALMdyoTlx18QR7pALgCZ9DSfXOt+Qdjh9LqjPe9xLtLNaqTNMo2UrmFBbS+
CpoEas21TmLdxzSNsqezAAR9DAXe2PYj1Sm/ENJOqmaBE/duxwVsPDWEBgGPSKXwyhGF2WbK3b1S
fkgaFmixpU0/YMA4SfvV4Ij1aCXPGbaaKJKtTCIvZS54CTeJkuvCN1H9sICyyr4GtEP94crqs3ZA
TXydMjGHvsQtgnE+5nPB3WWUYRI0/ukbEC7Mhutk/2cNVINk55tUGigEIbKncNoaFDeMyzkBubgx
9btmihgPz4zhCMpWVDOS0rInUvY9OaDOGlDd+1WGlcmfXlwu9HnLWGfAXZeDlV6HwZDJZIedfZ83
rnhSzJBX6d/n3H8QZNtTZ6SqqL4T6jnwsCSZD1LqdCfXwVB0iSbA68sYskeAeYpnIEFM7QCJSJMb
3XUEuM9CZ3aIXq8K3/Kr6xLMJExYCU5IxjWZBLpTp+RomIDKwf4yU4htzvluNAPcaTCFRRqxkhPW
UZxx/WRlSZYmGYS2YlYahULgNESrAqxp0vH9oJUWD5FM73FoiHDJvV8AtByN91j1s1OQdykX36UY
L5iCIuGNrxMPbZmMY5t8YknkqFvXVyEosqBft1oQOvPTU6Q43jVPXgcDbY6tiX3UcdtNObDcK7JO
P1ExTjO5Nzd0DAtjtYN84lJCDey/WxF1jjymRm7hBeJ61Qzb8Lylho6JMR2KmTJ1YRF7Mu+vxzqs
MggdL+KpIq1JYkKQ6LgnU3GnrNdJbGwGRwXqFlVF5TulipAP1vhbaeulkwJJqOt1/LA3jxBj9wdk
MKs0jz3RGjTSiJplMJH944Z9x9M4RqEqikYamLS0JSxiCavxtQ2LyoJ40rnj3UwXuB2h2SStDg2T
nyqNHsSVw+NKig5jfo/AFz5SHnUZ/Ip46xoQUhvqG84g7tAArgUP2yt6hUroeLb4St2WPfArZGWY
/IyQEB3cmlSvrk7AojJNoForhWRQurb83QLWx65roo0bebG3is07jnf8XGrAseU9H6xM6GssU9oi
cO+fYhdl/kTky7Bgk9DN3m7sQYuvnzNpZv5zvM0qh7cf+k+HTS0loOToG28qwSszoXjYIbrk0tvo
rf6rq6hf9aoz/f/Bz48Q+f+llwk9IxOoHL3laJci9o5XeTXJ+M1w5IQcPY35jSDSVFQRlnXe+qXk
nyD8F/kqZROIbPwiikgjFuN3jkC7P3bsav3t2LFDDyk5a2iPN1mXi/x+ExeAYKTz8pEjvyKhq4zX
Cid0Y7H01jTfaKjCVNeD4ULTCn7sO/O4kWqi/iepcEvePMHE6UbkTWv6vPOi0R3VIFkAhzEAtqT0
TBEE11i5pajXMSqTosrP3vdshjEAn2FZgG1M2cN5LwNGjAUew2i/N/M9CkWaaC9ddK7yN9BvMOo+
QrrAqCGNvQxv7oXrQYCKQTPnj7+O/Fl+hEOQNX+FIxxIqlGZ9swHxQE05oM2CbuJ+uO/ZYgdZGlM
jxJxffDR5LSThNWJWUqSInIL+lswE+/jAg/5GvuR/Q4zO0np40ULetvXd4ZKbLLGnVaf+9CAGuh6
JwUqncCoLZ59bO5yfd8pfFWaI4pN2Rx6LN6DPD33rhwgkA/2D/jQfNoD09VLVhWEKpS+Jx1vkQK5
87iR5B4HsC2ygXmDfSxiYzkYf9ZPE3muj5tWUTT9veWvbbQVTd7o3UXyqRl7d09DVZGWNfooO63B
FCZ/K8QsrdOHifl+Y+Hn5aHXSK+Pqr7jyg16wokI+FiXiGLy3QpSu0mZbUKiauT2cggSgkqYTjnw
30A5Xxufa0XRZR+66Ns6onjReeDol/59avIMjtwBnMmJg09LrI4hftt2hwf1uTPg0AUYglLZRy8N
CsF/aljLtYKSUXUXUgil9wLSZ5ru54kNfs2jy1fqdcFnPM/15SG8C0GTjJcky4eQoPzcYbeUo0uh
2xrJBkT4KcRmNdvDzcTdVuIXddWxdJxTFCqGuBZssr9VRPwNvfLDw5zmme0Il/lAZMRsU9dF+hwQ
xqbrDbUy2fpDMomBMDsyNijtm2lPk9zvVmjFzqBx4Cp0qkPvC9lAvvEIaWGuM+ZtPZZZFg7Vl2Uc
NIKp2cegKsu5pI2ExtnsLrgKfnM6M9upfC60eclyyY+7O1sYl0UkCL06GpWRAYIqxNeCLtVUrDst
ZAKTs/V+PfgHLxxbXioNDWRA8UpdeiYL3Q/DgikA+tUP69jgGK3U25RxkSh383IGuX1sgsraWhIB
HCVqs3mbmHykZuHvD7eIlRrntRz3z0lyJYuZQNEkv/MbAChEkd5Y4QftMMNXt1/PA5ySrs4m08v7
g+GTPm9+xUKkga+0NUl7h0HE263jpL7JF4XH76SVQdt7ky95OOv8abFttV6sAQWvJOgrIYsRm7q6
ezHaFFFIWHhBHiv/OhE9/1E6CRDrrRZGXz5r5dX+NJAakQo0W5DuSpTlP0IPArvioxLEUQsHu5mW
7N5bd6NltKQm3WnLglfml3bFximBaUYZJZVhgSMW3UbDt+7rhFXbfZ4CAykUhCDNjy+dedETDLUb
sdAR5kLzK0mnMAJLTWGTNYNbFYZRkDoGVYH+b3PLPANUcRvsqViHmL8CdBpELLwV4eTsYTP/jEYh
CQxhlJET63BjkU8jDE0sphaCTApwEi88MB2m5ju9vFS9MX4olB7inQfIhbebTzKGQLhGVQPuqs9b
m4/u3zOa5hgmbtyDuQbeW8IdvB10DdugOGzGVu7JssBLgkF75xorGuAyYQLrGZ4O3/eENPRtzIZ7
1Oxnxe6hU701znAwqt7sqhVMGdX9fN5+s3Y8FJ0RnTgled9rCRPWbadTLBZSWu1tFQgxeqdptXvQ
qnQ+38eZtM8ZLUm/g/Im0uQV8aUyN9UtC4ojMJxazpo8biO40zn+8frA7qsb4B+6Uisb4NT6ivZN
B9ZM1cRZwVIf+igQExld7wkx6mr74EktrYOUw+mqy1Ah7Vam5327Szu4x/1e+O41vBiptb16eE7g
cNSLxDJFxrPx64OqpABk/db4Q48Y/iljWykGEBlSUWH3QOihNXsgkHMtIMtSWjbwlM4JJii0uQPD
I2c91liEOsvz2CjB2juV+BLIhS7fnunWK7wTR78gqVfM+oJmrKGgspeDsWy7h1A9z+rhH7GBKuYr
KVqtbQhibMeY79kjT6iWYosrpekXXjh/zetY93ygUqfBSFedUdwD4VzOUt1QQwNFQ3pj0F7hTBAR
PJ0zbjJGwDm74sBDZSVNv3qAQiV+kDvS/FDcn2y1ncpop3mOn3EkZJtPvwgD+clsTrPWC0W9aslw
4/jF6q622a2iBvZ5JUpyeNfzA1TAb6fcCmBg6ucGVnfY35q27mpXotJBlim6Y7qQ0JtTvX98OQ0S
pcNj+i+EOBpHD8eqCF5TshE/KF95RWODvUG1CdrUgaSJjfh+FwgaiBvknm6ZvodTEEJIu1n4JxHo
YtuQoG7xGwDzCgabBDqJ8a9NUj9KtdGUw7VwHKcxwkLrDhse8HF9XdBQIG7xV+3Zp3xx+CSL6Tqe
cyBZ0rRh/rGtEG2ssWtUKMs7aXo5K5YVd0WEGoCq7JjMF7OeAbJqNVEcFK6DOPzq2lJjrVowq4bN
9eLUhVq2ZGNEglUHDnp+k+dwoi+4EbGK2kV5AbEF4JP2n+Hnt4bvJ615JfmzpmlCs7b1hEeQROQR
FoIP9s+SNXOCaDF9my9SyB4bK5/szlmq/gQmctu+AL0JRsoYnmMwi6wQw9QwUBTpTNcQMBy82EiB
3eJJjduOgWsY2qemZA1K2njLISrUbwjZYh0ZBVVmrOq0lHd29uGo892HQE3nlnnEeF8NTzdZ/ztb
Vhsj0LWGv06Hg3F8/Y1Ycw49UYuNNREbxVGnGwaRLpoK85WuHog6c+8PFdGL/+IR+uUEmi6KhWiG
hCisJexNnj7y8XI5/b6OzeaGT/tjJVrQT2hD0PlI3YJdbCbZNCqh4Wri9VMVSDw/FmrDE7wpoZUs
3NU3UDbFEFJ/R/px3Nl4C1rmJk8vC8y34dKW2qbqjeXPDPTgcnLi3S2GYDRCqUZI7fDpGOCeNaN0
VVAvNBKryGb1D1QduzaKhyj/vk5wRiXRUdB113YBESNj1Ujs80gXVhi25VhhaH7JFD6HTw4w5M1V
ptRYOzwRz/0yR8H5KndEKzbfP+9yypOpJg96rISS8I8jR5gxLnZvd5wOKO0oJj/tRALtilgsARpo
9GzbQzhZDpzK13SaVofsybl77nA0DVqlyV7pO9FpZ33SpvBkaKtmYmWiF7srOdrFPCx3Ca6+6inh
k8Tyx59foGKPWMFDWJm8zAj04rR0FvmH2wSPGfDAIC0SDWcZAP7Ol6eeEbKONEjW1QAVBGVbZt/2
6Q+Ft3H4+xJdiHNB06y0VVyErT0uTh7Lfiyu1rTjeGmoNkc2LKYQZdjrNM7sA/qBCIJOFfeXzyIQ
mXaF+6Rc8Ob0SkandjC0BxvpgiiKoSixR+GV9HY+81vbrd8tS2DbrpUB14gbDvsgOjvLXa1pmO5p
xGWaPM+gO0QTu1qLdQNFY8ouUiC5h32T12vvM1JzNJ1eO166s/dKNYbojHY1Fq0D01XqSKjD0P+i
cVOoyk4ZZ/p+biu5JeRjzKV2ya2gJ7C7lB3ryJ9iOOuX+m4rDS2N9L0YxA/5grdEuS8iIsV0DZTD
ixhSFdW+qa63ImaX/Bb+5Cv3ksI961uTUe9N2/VVoRyAewHZEhpVCEHxIAVFn7N75JhyMYPhAQkI
L/jigcAKQGToie8uhjzfjAgeQC0asadxE8w320RSKJOf8KuTpBOZKJwWQ/wBokV7tO3vgk+Hi2vN
yWAdGCE9GE3cn8/FfniMr9jiRFlqKRG6gQ61XRHWyT9Crce2VI92jTY1xuCnmcDrBVyUi3GBNw0/
27W0us18FyBc4vzMzyBo5jg9UMp2diwG2Hec4r0hh1NFSDsvEVXIMBA4SceolSVrVZnYz9xPUVyq
KFhQKhBhrviLT92ZTpIoUwd3rcW7KVZEqjdSEZBUtuPfVWS8pXHhbvwEG30x7F+5If+VDtNgKtcB
Ovj2mUSPOzYRmdzmUokmy7vSQ4z6jCxBvLribTbs6Zxg4MPyaUHIegx9IVn43/BwXJp/mFCwZGVc
9D1OFbwdeMnlgTWjwXbTRO+m2Cvi2AMniAJ65JDqQMnx0MSrMncDUIXKIpYz6kWvifPhBEI8U2u5
H1S0crWlFKCmOH6lcL+Oilc9muubjX3hcB4f6vANFL9HtdMzMcRRcbXj0My7bWRiJD4Y1zTQH7mc
inla5R4eZeZSLiz4DSORF9a1FktvyOdcOaKex6pAxFCY3Vweb1Nu07OvgNfBwB7lUg348Cavy3UD
sPfZLjGl0Kwt3hcTF27YJ87HedMjWsZUk9vPHAhnCQWO4hQ1X9+xOJWkJFuKYgwweWuKfe6Rf3bb
ZtISKlxtBbcgzuYY1fdG7UOx2xTRq4fvjCl3iyvnrxq4xftUbLJqpQwwlHTzzRL+u1APy8R53aeE
avV7GFtRQDxPJ9jcM58EypuWTsJlUB+eF9aIHSNiLdAXQsWsm3q+GYamAVWKX1HFhRTefXTmp5YD
M34reLWdhgPXX531Xld/TVYSRBqPCM4iRVbh40T5AdEGvALtCUDOx9szj+fiLknbIwCmvE731PI9
HeIcujRF+wshVOHUev/pdH1xMWJJcsdVLErDoJ/UmLZ4Vq3ehHl2zInGOzSNrhHeR10MwygXYigr
RWdgfEsMxr+2/G92lHcRQGE5vllb9WOt7VDldIJT/6wGNt01itHY2DHQGtR5DfWDGjZ2u0dhJssd
Ob3Rj0tvwVuPvoJxQ6myPyrO8yB6bbuYdqmuvgOBWkkdon61GfIvgxRmhnY8wybkrDrRDRjKX4Y0
di5yCNM/qN5RuKZzhf4VNcWmDaqTS3H72DUZjY27cM6NUWVeoZ3AlXmULl3Ow4ZNquOLPaj47U87
dMrSY8ut9d0K+DFQD6S4HQX0jyULzt3WnfxElYk2v8kW1FeFYAKPY/ApUgfYpO1KaAF4bbpOwPw0
8ysaRo7oYgU82EiEWfSskB6o5Gd7gDG1UFIaiCaxdrMwMTd+nv8meB225Wdx1hgL5MfobNHl0ua5
jGpGbmwywBhMyuG5tFXbGz9cFrdT/4bK9+CvnyOxen7UBL8IVQZRm6R9W+RMni3zIdjt48Ewsdoa
ku6ghX3jvI2LvhKpxmZFN7yowlOVzwKdGL90qqGer8jcNi74H6ivFlFrqnviKjEvvZVfeTnFkFXc
S9ZJr2HKOhGZLcjiQfKmI1r7JG/286cB/gsmkEwpsLd/GNlqI6qOLjl2oCMPxHUSo3dA/DF7K6Zs
kkX4BWI0LJs2R5bR3wC3zPfL6jN3VFe26MnCr6ehcbFgYbLfU9ilGl8Tq5PI+9rAxKb/7E/KEcIo
Ld1iAZ74CyLnU2N0rLJONU6wgtF1Sfyuq7N2V3zfN8wwTNKrf21WApwX75ueF1MSlI2rjCMpCNuu
NiJ0mU5fsi0uJPBGncKQO2wZSQfeT3Mig8KtV8YeX5f6tiPnHrr4kp3kwdFZe00xmx0jjKIB+6FC
glzXFwFMQsz0tNuPaBgRreDV+l4xmv36xaY6liU2ZRaIAEIG7qxqyFcLL8JP70flj8LRhZXsgfbY
JZignMtIPwwpYb3V4ZCDxWr+9Zfcf9Fc0kF86VpsfRS5b9baCahGRK7xgY64QK6NQH8+c4E883xZ
IULtzir5LrTr/whPKPwMICB7lPasLTWrXoiPqM8TfU4S882VP5JnHVpRQtLz40myMoAWVFQU24WH
yeEFHheiGcozPAms5IYtEuyIAT5IRB0bDeD8lBebEXJnNbVHHRNbgYWJRpyXes4xt9dIHZxhFnK7
tBDTjToDHBr44W1VlrDIDCWBGMTtW0yO3u05gJdh8RqlMRpqqFPJGj5vQ6ZUhZLbDUwsBVLrqa11
Pfm2gSVHTIoKw19EiUPYjhGrfcoJm8QrKEh9mtOHVIQ166+MRJU6I2mmXaTFDSBZnTovajUL2xPD
DSuFxoA3yRdDDgP3qEWHMK9Em43mDWxhemgcEuQafIqOQuUdgGKQELBs/Rm6Q/p1xyDE1Hv6/1PP
hAYbribYDPoGbeY6DrsNbXhUQ6vsZVzN2sCZ1k+Psoh9ZI4kFbqjPQT4GdM0MmxT3Nib+hgfyhsj
HMaMm0WgOUbWJlQJZ7bBpkywJ9nxTm4zM7h5x04JfwgZxYY7zO2QZyxXgHQxKwRoSAXR+71WbOaB
rMsy2HuDNnU/q7kqDlCA+9vpOq0U2AXKiRiJMvdGMeNO1cw00ZOcBGyTiZZ1eyU6rDmQtPJroC53
j6Xk+3FuAO8DnVkov8okuQeCoBmNJuy32Oij1kQTyB/VtJ8CWi4s79bA0KUV9xUuoP5va73wTLbr
n0/8j6q9nulNqiomWqiAflLOlw4ClSCaI+1TQa6Q1if0sR6PjM6c8PUfGSZ+U4w0wUWi1zU44Pfl
2Lw/wu5UmU11R0lnD/b34e11MiY31EjxN75gLx9PkaFwCziBVD8DHZocwkzg0iB+S0UJTj+pfv7K
kV00J2XVxL/AO6DT+10ztpOv1uoKeVfltQjcg9v5m86B8njfhLBJWDu8RkDWzL0xrZO06cu/Vpmb
8KWNbCfzWTgePGOmqLs2qmiJZ6MOSwNnuussZ2Y4XY9i9MaY++eexu79F7ng3exJbpjgmw4b3AA0
e871gv7MZc+ggHFWJO5x4WYjVuw6X9TIVHkE+DCyzH+AwnOOu08XoYuDnQclHHzp7HINr8iSFMEv
OWByFXv7fDsCBacY4lZAoGh7mOQwhkRSZgQwFQIq/w/q285OG+e+9ysEL+WdRBrmtY/Jkljea2jL
wWzgDajT6f+jAn6UKkBPFveMJIr9uexjWINOFA0A+G1/GEW8KCUGNv1xnSODkf2HeucG/NedG7lQ
Adb5fMVZBbtgGL4H/P9IZuFebIBw+IpIn+Odg3XiAwNxtMCUNAVBL0ozxkMXSQ6EvsahvdShEbdu
SpoXWtMSJ84/R+rgiO2yRqi5vSXvJP28KfYW5bi+C7ifdCylbU/y7hFrpmnPov8eVHgcXJs53kGT
7KschYVmdgEDeiDdv35H+clYCeKOLqXmfqdHRYpOXV4cZVdIdWQcIuMAngX8/UgQU2NJdS2mHT4X
X/HU9g4iwBzmnIvm55jvf7CegHQPRdg0mFbsjQoiwrckKzYuJvTc45GUcvALfuqpS/4yV2U2yMB3
1inMA8zc1FL7WW+hibWcIxNqTTR42rvfq0Y4DUIUOApU8ZnDOereU160dJ6zVOr/kdLpnFva8Few
i/qZkBaVS0du00oxe5suVgl+zcFYAeJfV7BA9of/PeKSFBpV4nOwQ5oOaWygl9K9pTAfgiJLjxOC
inSfcrzhSykDTg/yy0P8CJcJfcL7WhRKopmC2cUYY5I8bMDk+9C2HJNb6WHblC+dXrWRJbxs0fcO
H3DrtmTzSvX6iXDFb4Wdbht5tZkk241/Io7KH3gWDMXXi+KV7S2hW2ApV8u6SR4fNzkpcCSGSdJ6
iov7/KJ8SlCACRyQ4NE2s7Z7UVSrCWvKh8O3p16FqVVjNS/ySbWLXoYs5kOcUag8WEvUqs7Uxm1k
pjz5bLu0p6iJfKe6IBeYxcykxNYTOu06/rCp/exsKwIawy5q0c3XcSuW00Zvqbbe8rvewONRSInt
4fHjD5TfQObMIlQf0gWu+rjNPRZkftJ3rywE2T4PkC3FLnwmtJoJtNlTOOl8OfSTn/eO+hTcj3pV
61Nw2+b7YnOK0f3VJbDvdNN3g1OhRzo8d+1HnN3ZTwVgj2uIgR97BafavIi/4+KUl2/9JBUok51w
jU0om2iyrhU9rjZTxnCgYP57qMrYcOsi7Ozc2bTxMoDPzeChK724zIRrLq8TALHoOifQdOrA8SOP
UWNrXKHE55zQuKmK1M6Nyi8eMOTAu/4YPazpWJHnv2L4Mm11tFQfoQ7tTcDgve6Hegxj4yJjcwAS
MrPMzcTxj4nO0fbUR+L8D0SoVz4iFyBY9A5UmmAa8aJrRB8Lm4WQ/DHvBaq51uMn0ccWagy5zIAY
4f5OZViWxmC8bR58VCvqQlzOifr3Mh4hMuBRwin6rCy+qda4ggnm6/m+tm7iYGFC5XN0FkD5NSKN
ELFQ3jF/3uzMf687AiHWdbAcRTx8ZbnRRry6wF+GheF1WrmydPqFey+tbFteK4rSTLobOGaumwpV
opOpn5GHCE9Y/BaUVD9+6tzW13Kq+X84Sgqflq1aRISgi8DqMjwOKrxglO3E7GbUJnzNsFLhcsug
aNNExBMgJ57jLwxoXkc7eGcPbFbsq4VmAuW3oVTi/RF/a6+BWq4VHMaS6fKRTq6w+bI2hWVhfLeF
LaqGD/ls/ag0GzRdv92QaqRu5q40jlA0nsciSTfjmBHoRQwBCMmBWrwXPQ4hnq8rmscYwLhacRff
rrJCu6FtGVTf3B3NyZc6lEuDbxZQf5vSCVxF4oh6opOeSIWowdKifnHD86UGZoYmlRR346Iv34PK
yxpcqzf+BExA3NsDi5GbrRWa8US4hJNjreC85D74BghzcJ9FYxVi4wPCHC9eeptfenIewCycR3Wm
Lt1x2AXkpXl7gIe6SnDYFiNN24akwij0utNIV6Z+RzD69tGsr5IwZL1tpGWNjr+ygrP0DkrvsFNV
8hzXPueb860FbkaBGbX85lqXfU+kTQwiD4XGe2VcaTRhEoApYUCwHkH2kFjTY7t3lRzLZoLG7fTn
VJOHNkOvrLRAVZoV41rhcE6URk65dj780CNR0WCG72Nr9kzqfT8tNyRwMntBuXVgBdG85U31NXJX
8hc6IeBRnfp5OhAhu/LpNdM4whrGmq+fldjcBmwp3WJ3E0TU7jVMaslHz1Gh4nCcK6V7J3i4re8M
C2mpUY3U5tEtPudFldCofROBqOToJFWQe/nA3Uy+SqE8sfZz2mWji0NIVyV+WScHqNK+J72YSfRQ
/lhb4Uu0s4xTMsg7JpYvQVkyC5UyBg3EixsytHNJjcXMKk4Q6ReWLzh26BRnpQwTaQNOZXF1bIq8
SLDtbTQrTG0qW7gToIwgMwprQ7nvXivh2bYbEhAgWoMtsByeQ7nrcwjxcncExFOVGjdq8qAmGtKv
2MVwGoUNfdzvxXPlUbVPlu/UoVQvEiW7ZGjYZ4I2y5kE8qtvq9DqSHGWAMPWTUo6kbh7gGaPWjkc
pwYJQ9WmlkuzGVw/Peko0HgxJ9EBynwKcjjCFFiPsRePtHfUcBgi8K2BgoiRp52B4lni0lsmoeyU
TAdEqIni+6alATWmwD0lG3CHX5OecsUk0CQV4PtQ0jBL6ON/FlsqONKXACyIrBBhJslJVC6WmXjJ
Y1LE4xVXVafm6GLXO0CS4qPeTBtaauuHPg+0WnsbxI4GgdMOE53LhKvLAKbDD/v3ErocOHm+FDHK
yczFuxgBfTYUX3qxu7d//HjQW1R186CNdl9PpImftZ1vZ+gQID62HDqL2JjGSJp5wKpz8osjQ6qN
w7PicZkNfzB/mi+ZcOrs3qNe7IKTNN0Q7LJoYxZtXeoelwbdVHh6Z7mwOtLTL2sZv219muZ8CiTI
q1bD2ryitjzq8A+QAqNja/lfMYi/M0U9liGG/9ua8ENr/aLkYPV2SHmTTLmX+GrEuRROn1LifZ/N
WnHwN4mPfqXthSzy+1LUPERYJxSdn+qKcmraK8rGqbfKXOqQ1Pt18QR5qP7Fo88PE/DfLJa5aAl/
00tQYmzPQXG72DGWs8fQaGpCHQIazwz8a4mRcZE+H6MFHMWAG8F/RAQX8dp3qP8wUVtbAqorIsAA
L64+y7dhoUHNTWPxJIzzR7oVdSiAHt3Wc7PaUpG39m5xMD6LaBuKqsIp6ue+/u0J8+xLIbHgtn2t
0xZCU5TzZyaEEnw4WqEp7LbSgs2fBdnHI5/CObAuOF7ekb+Pc96ndOtDTDq/grCwfnYZTYNtaVJH
qdF7frI7Uwkserb2+3xNVZN86WbjBk9Ad5xGdeugTG64EhtzJPK+lQK15yH2KmvYOt6V1l6U9kEV
xPJqSNq8JElUAXSwkie+HMLpOi8J92WSxHWYcwLOF8wpxxuJSZzFdEqM6MpAfllXDEkzAnu8EmH7
OrMooYsprgCeSeG5FM289iO/4d+klAyUGNt1fE05IvhAWWlzg4FMtlji7lFPZOjpe2Wif3nWKCnw
hhbXfsaTISZ7jp1iTHsRLSr5XR/ezRUA70PhfUgI3KtiyXatfyHAAR24QmbX7qhNqRWZqbsVITHV
zGdzmEbzXGGWMCESmajTEN7WyFkA4XH6TU/ZZlvfbuXdn6A4PIjO3YYIc7IwhUcDIwiE+svV3ZJp
Q0JKAkfckxsYG9cWSao6zz5T852lD39MyRGEAE7v2DzTNDtpBy8fjdeJzDXJOML+hs5EVG96XG5s
VQtH2oQWDAaHfN5XgHTOvxvM5tnJAbZfJAPaGYfZnUZiUB/PcFyKwv9tOumTisYvLmtOSbE/eMNP
6PBO/xnzem9F0X/h7j6gC2B4DcAzFJTpW3AY6PI7GK+FHLhtFjyU/0e0aVlK+/IQ1/bMe7arSFx2
3wwo/vb+UUxvE0H7pGXtziVg4zZwFUtz41uKYblN9utVpUklpma+/nad+pjg5BG65B10QK7bO2Ab
cTyt+j7Cvt6BIutgFSfcBpjzPMdDFsB60rsjqjQHPTHf3667Kkm3SxRBqT9/NMRgnYLAqT6xVaYm
butFNQ/ldhrqTxNX1MJFzE4piUtbFRKPcdGPGfZCR4Z+XnklmutUWuVk5UAf0xn/idJ8iPS68rJ5
IfJuZipI/mA/RotA4N3bR2jukXAsV5ihoKyMg0iA/3IE+6H1mKFh3HAdkRcByoDyrTGEmlwSA2A7
4dgrkiEi43sVuKK38fyTAtC0c/0k7pUaI8v3h6LjDNwUKFJneaijmFO4qVM+iZy/VTHc3dsUvkTA
yNNZ8ZY5UU5tFggyz0NoRW/KCLwGjgHb48RxrrhqTI0tmRfi02upZUi1IlaDYxBrbxhpkVr1GQsp
4GBaNlyZ8Dx9hfBpL5dZJYNgroi/gqxCKMxqdPCO6VPNyWOZZvUCFQq/TjZvlzTdYkPkhN9yHXrK
sw4ABrT1M/G7RULhBVndgIbTCO4+uziDTqXIahirhej0aec7UnMayRqcMwFXkrsEWkitXpCOkrQg
etoNdJbuwlWv7t0AainR+uRYYs/cShF0En3VPvD9BtPzJtBos8lTZ22+QVmiMqeQeErYJfZ+8fOy
lwj3ZRNc2ifF3A/ehDcuSJEfSpWqsFrgN6qVzs15Ef8/0KCLxJHm52olozkzJuXp4dRCSa/B20xH
37kjNxVZvgwm0KM8tc+lURJAVqEU8SXTgvQP4yezht+UxjgB0GEsyr6GYvoF/yZK7hh7E3sGU+hK
RZ3YikBjtY+csQRgLv/tLkKB0AtCSI4mjUR1CfvHl1S5wLf3Eh79PwGDHEDdcFAUvPg6eU9LkYTy
Rlywr+3OX9OYnbjch1zz73UE3neFYycFfyDLDoyQbwdtXwsWJbSwrqoB1BTC9DQ40Wrv+f78kEkK
FhkVI/Pqtm40mzB1LqfWYwA7zHJIZ8u/wr/F49LZbn2G+iEe6t6l6bLCILM93QMvfzgdIpBQNObe
bWsE+dJHRzSq9ULxwcwe8UmIJgzCcsc7Y4fse8yNxCV8RkXeUfOD/hVf6RiLvb3BiSgq8RPo2Gnq
8Rt/vYR9H50Hdr30puVF/6yPF6nCcNxZj7hSUd9eT7eOKP56h4qBIbCKTUGaMmI5FuRhIhdTwAIp
ityPqX5UeU2YlEBAKOKSlMRk0L1ERGXVEpbVYi70UfaUUf/NhhJ8qyjvnDDGVyL8Thoj95WDFqkl
khh/YmhLPl6McPErmlbGgvWZwKVFZVFCrs424KbxkmmXkwQ6TIIgZPGebwblZtGtlW/YsZDsImpM
LAUvvLVetdWr6CAFKPJgWT1GDEq/EwSuIfdDlVix2O5dCJbxR2iToezdS07B/+X3spwB6gmauf7c
WOdooprwC5tHc+EhJka0fGW12TgzAidM9VlFt1kK5ck7Se18AMqss5bRhiReNX2e+V4nnOxSm18V
qQRpa7CRy5NkbrSi+ZibbPjCvi6BSC1JPeemJQowbrvyqa0TpPO3/Qa+0WpGEo4c66uvnaYbqlEg
eOPxvdduGTcSmghrdzA6vsltbze+nmMrMPXw9MD8qx6ULVr69H07GyHPDih2bCR98jRHMhNrY95x
+11dNLAIjgVy3ZS3bqDTghYd44Z5DXw604nTRwgkSAIsifPz/e1GR2JQdLUTjqDX9r8lRdk6lqUR
FUg1qbgLkQVpyy27IjHGiekm09Y5AnfHpoBjHfnLlWEjT6Yo+pb9NSsS6Df7/OeAJirubumC9Dwg
w0zvSYUmddbhHiSsr3E3EnCC82H/c73xnQPi0AhO07dGjRwOaXXxqIg879L6zz7JidAbL0DsYdrD
jBWutu0KLhveGWXHFhljSAkwN5azVaae5mhLhSGM5bmI+NI1ULNRyrvSmDEuiC3cHRh44YGQzYYl
NwQNnCuJ4udm7QzHc3xV+dglsyZU+AKEn8Od49Q6TDcnQA3eAGUQUJUOiPVPRZTNGozQzJMUTmPk
HDQhRkXJCcd/dyOuzOTgqU6VOpaoBUefbpPaOM+jJw36Xwf+A/x9HkyjZM0PZY0X2dmBKxszONwG
gWYDdDLkWlAourYhfDujeI8IfIxHYL5JHHQJNI0ukLMCbEGxCrIp6GUk0JizCi4zvxNBnBOdHzMP
PVnyls+9KdYT8m8tlnOC8DVonAXuL2bavPJHxmJqUYltr6+hYBUyQeql39SLx/Q8u+yXAUr7X9fw
wjrCp/eYhNUm/hjsNV0kP3HFwVZBoyYKlqehFwYMVwAN5+mCDavkYN842/UyVFMxf0V0c+xdAtf3
rKFSMSAPdwZq48nGdyyBi/HjE2uuc9+/Np65wmBHM0YzbdY9qN2hNdEI7laTILYNHi7+yS2hg/BD
fDBUZO3ggC7Q+Ngm3JRTQKzQ+O7OUejRS1AdYdkthjvXYyNXnkw011hl9c1AE0N4tMk+8h1vdVRy
UmzQ1UXrwbRyYH9tdHAS18qoL8Cq/z4nfHNWiXcCr7RkMLEFQRZNMOxrLTPp7mAznniaXmrnQhz9
xR1/46FT0aYNd+HYDoiH5Mj/dlttTQkxbbhO01no1cZZSy79B1QXzuhtrvJPQB0QRgqDt7VicQ64
yvPZYY0GObZ7+cZriAw0LV90tshthJ0F5uJC3mbCsSMXpeYjpma6FDUzaYCAxHiyMzDu5W6l3Qtr
r1TSK2GeWg3i42ryoorqKFAk6HsaqTdYymPIHtjXlkRN+9RSaaYanF+FbUGqgIJWEQ4y/w/5rczj
vZVtS/OsCHzSpxs41gMUpCBIgykHi00Q5neXepJ9xmSMiGRG0VSyDwJ766ZqhxOvPVkKZVihLySX
F9IvNSRGvkNsq/PSDT6GaSP2ytpHplFTkMHhiiMPI0o6r72RO8kZKkknL/tunT3bTIG/gZcgzkPM
9QfkDUz0FiK/Grynjy9oaLZQP2cb7a25K+kFqCTyQ2lOl7Wy5F1+W9z15Kj4tnnkUz5KsvmLdOe0
HQ7QFq7Sx19Yl+JtMnsziA9PP028HGP9y6/XLT5phvw/EcBGEacn8vUC5reYuME1CR7J1wZJF47Z
XlSvogXclxcd5FfLn4FPPmAsMQRMsSYRoLRzLdvx+XYX6VkAp58QzIWtjC+7hGFt6Wt0p4z5I/s9
bTCDdn5J3bLk68muV81x44icKmSGOo8uFbS3udPlkKeOJdZtF4pfn1g63i6l8v46gZk8DgId3d2q
x/SN/bUgAwm2TLVTZtPDvo0Zqn/HUPJ4vSFUdqlpx9RJHaNX54AD9dNSESz980xn1ruJMs5+sf2H
YX/dqV0vrLwY4p0Iibvs+ZsKkekqsc3ONXZv3FCPRxrWD46lOQ+sdgOcr7m/sUmJVIi3e8j0miOu
vMyNEl88zfdo5dkGvVlj+a4jrYgv5g0NEhrGRAM3VBrtooCKH5vP9Gq6nfhur8hqjOdzw4aK5Qgg
xoIATO8I97uZ2GR2oGUhfa8Fs0BPXFh23WoJK2bop9/+Cv9Lf1fdeCbG+a7+F1LIthp8sjr56Fmh
HHrx0iFSqbz1FdWOz0EflGlM+9n8FA+8pj5bjW3XrWl+l9pichRcksxfWWMgjQsMRTOOYJVUfH4V
oOee6UYN4WsLTzoCtC5h9/ub5FQIVDamMXyYqfX8RrHfq9F+5Au8QsCZkKQdfW9YWxZT+npFGU+P
UXbP6fRT8/RPfuHgfSk2I2p25h0B6DHvCpqBzjNzAmPryAnJjFGVPIGlcnlLzy4nEZtlB/5OHaM7
vtkRNDfXGropb+qSE0kkdl+pdU9Y0hNof0mKZuzublvCYSM6rLDz5ivMag1Gt3RR35eJf9Avlegc
Mn0O6mruqNueiGKzHnzsjPKZKhimKGm3RNudpegw57skjVz1VpgAVEsCWZ4rVbguTXMBhonSnJLa
+yoeMsDUzqqRZDwU4hGgJMaorvF9Skf8dCZJPjvnLf/YxbZIjy3jw60CI7vLvReGR5gbQHehy9UL
QbxGd8w8b22BpKeL34c0M4Jv7PqgFSfdaIjxHU2rUpl2952B8qMbLKJFLZpitMz8pvmFAWR603JA
aYNcOWdoht1Q4uaDr5myteVLLEHyWr/WMwEjQ4pKTM3OPdq8R1Uzf9h9HbdsiSgWgt8NiFmbUVqf
XWj46ZRKx9K85WBHHBe9FrGPF8BBiOOJjHmGnCujmxO/tREzxmAgNct9d7XWGptCECM/lF34YF1m
+JTiT7uYjIOX7NWt2QAa15d4/K1Cup+Srr+KH78yuSW6yA4MqJDT5ea4g40n4hrZgaSBeznbpDp6
daStrAZph1OtK623yhD0VnQZA4rrQeh136ZDQE6i9LJp5YrOFhREYfAeSccDT7w9iGuyCkXcRxGh
6TvTvErvYga9OMEkapKdp3CR3SqLkuQMBhFWWKnFxJGKgH/jQlh9ixYQU+3+zP388ZbDBCjHKfp5
uiieTLUI0rvyYTl44oijd/qpUY46SUEBlN2viv/4PjfIZ7dyad19kr4eryMtxTZ67WLP/v5L7kfB
yLAickcuUbs1EeFt8Ld8TD0LFTzy5H/8ya0s6QcakqI+m8Lr9guru5I6tUihKy9k9Q4kVQ8tbFjv
ljisskDNbRmX6hvTUMVSNGUW7ycfRWYqtidXGuP4aaZXTy6ZRi1nz1RuBW2eY27GluGEwHfmQCV+
XPMoP1Q8tJvTUJhbLq9IJPusq9wY5nppeZUYyUbxBwNcXwJdoOCFjttJsQu2YFG9j+m/i4zQ//Ka
YqdS2IGTo8GQSQRNAUXOOo9V3pWehNlzBaQ/y84DaIxNnaOwr+SG7XhQ5dLuKKrJKiC5mh1f0ksl
/QFLrCqsCKVexfyKE2G1n3XguSnEo7TMiSDm7+YgQpQnRrUm2jcJu3ZvM7BrNy+wUkAGDoqeCC7D
YjpPCYvt52PWB7q7CY6wwlwy9Yg55GG08dkRglEZ6zDDc1NamYTgV/BOYPni7hEKGigcQS+w+LSx
Ru15mn9kNZEbeWu+Omgw/cNPvWC8L08XipgKMWkail/09b8KyYXUwcv1DMxa1VZIckGAKJGVCu44
mzafjKJqTfJNQlXJR0jEToWz1Oua+5Wb2zzHTyMZjDtfvkZ0W2EWNpqQoYJC8ZuE0rOlGi2BrPYV
JO4lxXWyX+BbR8P14rd0TU9ONEACGAI++73wFtdcj7i7n1KyFkpqYgBUcrGYQ5jmkxFzASWy6uT+
zmspxSF1875Q1qD5Njzi1G5grEy1GNkxh+sGYEzfyP1QLPcm/hCRDGJp86HvzADRTlTQM7g6qlSl
5d4MJZ4u1HLVmJnuyrkSNxmTIlG6lAkY6RthC9jrz8ql58HbWskZyx69snJBZYG10KlxpfOmfxWS
N9MP3+bd9yzxDEP1sVgyNFNa9LqCukOT3XBeEhI6kOqvJm8JHs4yYyOgej1vn4g0N4uXl9tFApia
7DfSgO93HprQ4JG23i5XSSJiUgl8yN6P1+CZwFtARy8XzXpuCZ8GcuvS0vY36gdLPSNUo6/exu4N
uv8NZt8BlQtX3cSLzr/CWIRBOjLayTt9SGHsP4POUFlxn/G24DLR8r31kXy/0mhxNZEA7VnfgVKq
M9LNE6IHTJpMJYXF15wlB7daUSVT4ccgsROe0p4NuTe06l1/tVRe0rLWWe8CgIHlLunxXdwtRZTZ
6ael37nB1c5fTc3NqGxpiXJ8pOl9LzvIuX0u1uLt6381JXl6j1d01M8k/t66ekfmvsnW5TqChlCZ
qd/XL+NmURJSKIOw0FzajBbD+MC9WjAu/21HXXTqgfy+OviQUE1MOZc2q74Z6a7854ulwdHhJ+fY
KKEymiRWEPsGA4B5Qjys6dFCR7H2ajRhULfskJtBmbLsHOk0srL3LLpGMQh78vykLfN+EssbUC2R
2HJ1LCo6D3SdKoWAAlGEJaHg3Vke41zKVsAr6PN0hdkI3Y9fdbWsbYCJodw4FQVVeTJwX3ogb9K/
uRVU4Cogz3XUQUqPY/FivVJOvtpz3Ys5Sqa1q5bR9c5rsNlZIqn6gcUkIk9AGr6DlVTfTAGx2Zre
HXpTdMdJPqq15ROkIcoehdFDYX3G+LAjqual5etaennsusKxbWbOBopM/1mg2lGvFI7itVVNsFOh
XdNvb5rzUAfR6H8Nep0BLAnIc+BKm5Mq/WnbcBilOu2bndouWYHKIiK6wlYcYhYOR3qkKVq/JsDd
/yeOaxY/2795Ke2ROqfX4O0VgRJ1mm3hUIj5mxQ0QvbhOTRplE1QRNkceJ6kvica1Yf61AsKQQHM
NfeiQxhtovaX0uizRUruTlM7mGWUlqe8t5Vl8xhLQLXHJNwSxy6imRDr5zNkM+F0ZPSTlTClDUk8
hEPD9Kk5D+vlQH0jE7zLNoKq1qywjObIrsXEFJtVic2Ujpqbfx5r6sVfMmGrBbHbwtKit+fM/dh8
52raXrJQ0uHM+yVqIw7BMbSY5lZ6AiXyQ0RmkBJhhrtmaqBTAOWxSExMmgdCOypfvLfFMH6pP0Jg
H7P7KuDOOHkeyJUZucjqi0Bey9wHOxWgksA6sLJcbxDObn55/Z1EFdeYzcfystYocaNJJstNcNjX
/gV7qlsrpCzU4DHn0vqFGK8hTcD9co/tCKjSGMSR4/fi5/nRsp+u5bZwAoEHlymqn29IW1bwi8P4
lO515XKI6n0rZPlq+rnbEslqnJUJT/q9W8V2rUg3ugpvb7Sl9efa2gI+A9dAGCfIhK7HSO89d0sl
jldHM6guLAiSkkaA3y4rKSoePM4cdi2mKSBaEFfO4neSJrMRKib0qNFZv+f5pbqW/XPieHDJtzT/
a+mWkykDXRLbFhA3ccOZS8jYBEVo7631FbXLx4vo3K+6znMg2x1T5/CbloM2JymwcLSjx7FPFC71
HWd2X5DW0eJa8a3V0dpz9jXUjVrZEIm2n5SXBJz9DZXqlpP05788XUEs/WjaSkyt3DxFfO+UnIps
QCsNp1k4Z2HLT5JA/sq46KcGM1XRx/0kw1BhczUdLsHr7Wu66wIk1vX7cfCNIXZYWYDLs+IaA8cu
1fR5YJmZ3cTTjNC3kCU6ZiJhG72KNFH0PNygb9sW2m6eBbH/SbKHh16zC42ZS7mU43Y7i74LHTud
wkB1HGXvJVhR4dCo5Bd7KxocxRoxYvQPFv8cPd05ozZiiqo+00QIrZrj+GWF7lfdPnh0iKFEjEBq
ceDvHQ0l1saq8OlmCXa2AzKBdyGHtT28FGKGtx1mD8+8b1RK+f9KjHANDELqyDAuVUmrw9gAoJK3
np+WDLpD4ydVRqbtJ2ZRprU7DvyKwRhJ0EzgDSSXp5awNbg5OAlcVVcAPAjOvpVOw2RQ0NXIt5Yh
xmdIE4NG0I4coEbYqaykG4cLvjoHOvxvyI7RJU0rvRCpYWHmRJC4nXl6ut0sJnfmgtTxdK/pGghg
AgKa1/e36/aqGsaFMIPkjFn6JVK+Unpup5qAlVgtRAgknCLJXkPn/8Dif4pEevhCQL/VNU9FSySG
tGMpiVkkiYFf1Kp/lg02QIyY/vaCGRpD/MLZUyzklEP2klirHiSQ0q1C25g8Dc4lZggIvWVGChRd
Gyy7SUKLfqEmGWpzNnaFc5GeAe1sTW10dHTOghx02iMhuOBB6w+wLxGXQXydO3KbQWVxOEOgfRTe
BGiY+qd/E6qJFrijKwjs3rwHJ37v9a+93kVeZmmQn/iLblX3/UtkfGmWbhPfh/8sxG0dEmm7H6Gw
+WAmf3VIQEhm7ljT+5vrXSqe3bjbV0XlZc2HSh4zUebKFjShZEKAwbN/MbE26wXYdDYOHlpgCSQF
gUSjvIAPRABX358oyAcR2RrOwa1cVRpxe7cnmmayz42xTwI5FG7ANOkUNB1nmEWrAXJfTMqZWwfY
DeukAGOIrDHg8QTFwpU4iMCsh/KbaVZ+oLhrjruETeSc0YKz4a8J4zZ3RQIHkk9evkqfcdnb+WDF
/NEib+HH0I4TPdBPxYelEhpz7LSe3X20Oa4zy9kqq+chc+9mw+LxRlPF24u2QspuYqQWT6LY/KoN
2fJucPzUZI70J6L0zL443Ah4TUuXMzfUlKTiM6Fg7nJXcm8t3YzD78EnT0Yy/atEuo305LFpfVUC
BgpjWf1BAPP4bOQ9GRczs3fedOq65lLGj1Il1Xoqsq2ZwNDxsDRzzsmd3mvACUj//3PO4xSXf3vl
V62mj5XTLS5GH0D0ZKWxrz7TKo3KIF9Sbj+XM4FHbenKTpbBBSYkPv6bghnzsHAm3W4AdfUhTj9H
0D2rpVQ7zAEbyz45yU9EK1d5A8t50ZF3XZ25MFzk+YaZJ8phjXZjSGdaWQsw3P0K7TrPO/vlGPUF
B8wJwsDwZilM9exk2wMsCzjV8xyxxyofKkeAI6PQwQLJLp841h4bLAigODPAmPYH9N4gcsVVIrR5
uJmvPVn/fPWX5C4BwiVW/EMBn+1kF6pyitBDTwzGpFIhg61xNUmGiLMZtVe2Hq+5AeIg1At7ag1W
wyXPbYkzaHMgIVCUAJ2YXCJZWv6bAwG1S5MqvmZgWGEmUl9FP5zUtzWfwgDVALwH32y1B7Av973O
YT+vgzsWaZTeUbdcHo1QiVhpDqqJqqSWJqjkGiCOCi2tKukzEHgtfwrG1pBg7jQQ//uLxW12A2Po
l0sJ1pdbLxNUMUSRs3HU0bs/n3+a/pbYglJtPgfg6vgDoXvh1htl5qdGCjzGR+jCB3j/Vi9J0Zqz
TDWeJ4Qiqj98kU6oaPh/Paa5jx3/QaJl0UwUsHEHRvCGXARJpyTZrZUk4+Oh/wv4NnXNRd4MKFTl
vLZrRS/LVkP/aXeAqyhCvvwyboe3sHtaLfmdNQP8mbfH3R8uE0FIuEtQkKb7kf5a8Fv7TAJwCqCC
G1vUaXcDoArQATdhc3Uz5LsiQ7oPL/ixZTJl2OQCgSriG8e+VMrdEjBydwekXi5kJwFFwOeo6qM1
sGcgfdCg+FBE6vWMhFzkvaVbp5526HXo16m8VHJbXJDzsjm7U821ub8eoJ22Qbl68fw1ahPHReuW
cydOlFAEXslGKYJfMQ5sgw2/MXP4zX0Dne+0PKxSFSHvFGXHH1Huo1kDIYqvPBQ8qcy9aNSpnriK
iEA9rojiOnx3AM2nKjCYxMxwyPZjajuqgw0JPx4JTto9mRHGF7bRR0k0PeLFV4ibQTkKfCI09t+t
yxi7h9IFvzX1S6hcTa2/lnALb1ExYPeE
`protect end_protected
