-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K6A00vcvro+YWz2eXpqZbe8fPV/yfR/CP8J62Fru1nKsLPHr0zrNhMJxfLDNfjUhpi5/4KJU+EeZ
RJ6FVREH0FMBwBrHrcqr7pP3DexwC64l7nEQU5ujmiqIrE/g4kAoRm3V/13/3HryMHDv2nWwuyqn
JpfI1+5KLEYwSzCeGlSw3C7WZZrjvuANvnQ07jsPYZ6EjUrOHrZOD8Oniduyto5uPC9HpHE52kIq
VgPRq+QsXJjymnhdu6wsbNjYAAyAfjZApN1M5xIKwW76ap3whEGhjEkLATd870I5m4VCrwM+8JLK
JWgnr/qyAsXb4UoNsk97Y6aibNRaAsaosQ7hYw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 90624)
`protect data_block
ddtJCQuDx4sXbVEaqZK5husnHMzKE4sEYbwFJ4/CxiWzP1ngARszF71sYCuNFmuiw+tNKfjxJuiu
Kv0ButemF9MXtJiUhyaygq4aq9Yszu3waJK2fdSYsuYVxo+iApW9FTYz9FtJd/KsPRWhg5YcBTe8
IbJhQK4asuKF8Mcs/nLbSZOyqVqo9T/HSfli9ouHApIq31f12tcEl1ie5/jiKHEEK7Da32s+HQXH
qb0+vXAJAjCuFIVXI7pYNjB6ZwKyJCDQBlkFQ74Dc7k1KPj2gPSF/eqhdCJrNgU7ynaJ8Q198hkv
wj+PO5MMy2eb/N9YFwLbNMhirKDtpAmoj3JClX+TeV6eJFkJxgCQRN1pDhV15ZMXQrnMJyDIBIF1
R8bkgnovpmX3iVBZZjOn2NaKRDjXZXCE8osl2d9pWM6imSkHQZhGcZkhToFu5NNpCX8WYbKF0Zkm
0kkviuJTJyl272ZgRio7PrpdH9chAfYzgOY2ZXcGGVGqfS0F8KaSoDUmMsdyrlXDLbvZO87W7C6t
ajSin3E8OTzexPTkxy5y7BSAeF10mIFBpLfZ+HZHpB1uGCgdeC2tXOSB9yCeRTkEyuUEQ5JB36hf
UpatvfoKv5rH2yxOr1DgO7sjNyPphuFdGQgV0adrriuAgJgrKfGzWMxve3YdTx6XZnEBVmEAbV1T
yn1nx3aesM47TyAmwE+D00+UaKYBvCh2MufeEFa5kjmx6b9Cuq4D9e4lwLlJevKihRQIfmT40KvW
QrY2r1WSi1RYYwI9kHLOWrz9WopU7Es8sGDiLOUck6G3Y1jpnTL9iZtFO17FSrWQWzMFYFzizVhJ
F4L1gDNiQH9XKAHkNT50nEfmXZz+P4n3DdECamgmZXp1vGic13TmeIyQ7oYVp1rxBziyj6963Nwp
xeFjw3mlyoiXkgS4f5bh04VbJ7j3ncdBRY6430YICXvbnv292Ky7Z2BhUzx/mz38y5ndIHXau5lz
svSFCmNArtBS9Rjec0jh7pZPX58CPLNQWlI3n6m6aHWiTIJsT7oE2ChPWhI5tUmkqstaJu2qa06W
cZnnuM83QtLA9orYfcJvhmQVytN/yJ2V+p1U+h2yM8NbaTLO+7DS8E8LOqZ8E1e63mmIh/HpHyfZ
1JfQ53yab1r8mXC4DtUp8C5oYGovC08ql4wXilLm8/ODPQ4c37/GIA7+Ivi9YW+qihdrutrvFNSs
M4KpCK26otkyM3sEgckTAB0QSvjzyuQjJd6GZa9X7XsX1Hz6W53L9J8aofi+TeVrIsZOsZYuoNd3
/lyVG9UeCqYzqA5T1nlAbdbzJaGU5u77XcxvWFYH6aE60SM5iMHn1XYXf8pbH2iUDgcgv30Uw8oT
RYfrIdBT7dLXBVknwORR2fFmcka7qshBzY5XCBBYMqBQqBSzvkLb4F8rJQaqWPc/dIXX7fwbIsoe
lQGdtvDfUlJnKlkKkYzAMVZT4dLRHvfXx1AEAcdhHas2sqL47jxUZqgJePWAtirWWQZ67PAOBKnh
GiVvb48yO4eXSyD1/VW3zLyt6qDnomI0eOtz2SF8U+Ph+ACsaznNZ4JVMzNwdlLNKq+74MmsUg78
5kqpYxOAp0dXv5YMffXV9rKBgBtbFcrjRnfrzOZQz2rR8LpA5RsyRIadNbYaUvgrMdRX4iYLHjrs
xQvKSUmKbsQJVmYo+rkNAmkch74HiZTOCnOMp8Ljq2Vh9KNi+MRyuVT5PAqhx/GOdgl7T8xQAL9v
262yaMI8v4T7mXynrpR4RE5TrXM89loSf7D/j7Lai1CqoyuqiG9sHjLExh/sQUWJfGrhB/HhO00c
kCQ21pgfSigTCtL7NmrZG5VEZ6pUseUTvrU9CtrI1aar7suvpnROlCPCcBOSU7c9Bgq/ROybnBkU
Kz5yW2aOTxupd63rGtTylOwYNMq7DRhK84uoiIHKFOwpXLAujJz9ZtR6TGKbcgsQ9kbNWCbFiMu0
NKVi5s4SsHQIQwYsuCyQ1R4L0ibljl8Sqgty3EAthDTXyhfobxQx7vDSr0dfz9nPUHsLOH20q/F3
c02e2DqMdAy3g0BW18XPF/buC/Pu/CNG8H+DC2bTfh5dYGXFGxGQwtzQrVQv3JoQgd3DPL3Q0Pf9
AOLDps8JOvByiuJhhSIOJ9cX873bgSxbOCB88x0csZr6BO8YDh4xCBlR6D+Jrw7rX36YC8INEkJU
nsgM48GVZyRodO2gZy79k0gxqDVKxpMlB77BuTEzhbFb6se0A3PKOslUIb//AP4WlbWmbB4rFzim
zlHMhQwq6Hu2oN3bnKHXnwcaEb15mMQMCaBcxIZhrbZ1/shf6oknbGYOA/AVQdspZdTRrc97scYd
xPmPmIiZJBU+p51biimoHAN6G4w2Rqau0oq2pbxPfElCm0HWvjiJv48HQwliipbkRXwh1xgt5+1/
xzvICFQhz9Y7n9vdLJ1Of94z91cvXB5f0y33MLW8mYGan/Qk4xRuhHEBujDW5VWYioezFcnfTb48
1qa4XP99FfRtonAl5/f4aMX0qR8OwealRFpplBY9fZ8u5SYvBqVO3+vZTJ3tnbClYS7RS1QqqO8w
UexHCBxKQhDV5oJiR7pX+waIB0BDHLNB5jmp+F0cw8BnVxrMiSS4OWdfItMFRDUjGP94HDMw8aBM
8iI+3ADby5un9A6l+3RYJ9536b2dfu/C8uAOJLq8fzOfeLp87DIovV6YgJbK310WUlIjMb/ZmiaP
iy6cozQF8Y4cy666Mvp7D6R0Eg7fs9X+x6zBMHoySId+5Xg3tUlcwrKK3TDceruqs7P/p36spyyT
0baD4MGZoXQoHB86cDkzzNEbLKuMglS2G2lQ50UjiQ/nKM3M+u7KPaTe3AEp1gnNrkn3Q9xSk7Sb
I3xQWI2avbHhov6lzJ/hYRi4yhJQPDzt12I1UGlfd7NLVHwIkJBYFhOlj6liGgqfp155xywUyPGV
GAtcoUGo+BqyaGVxR0ohLWzymT/2ru3tW5YXAzKsS1Y9CxL2/1OSO+YLSQoCU8Lh4+/UwLuDhKAl
v5Gn6lQrGHekUWDVqpvKoO1DoKlzvmhJIKMA79lpQDLMRTF00PHpkXNrEcqdabbE815Yfx0xkm9H
ocyja1M9MnVcDMgiyXwJico5Gm+0bThIQYXwtLvGgurNJA2sH6VumG6MTM6hCPaaM91Avgg3kg11
tJZ8uMpMCB2RnDLVZfeJA4zXxGh7j37B5cxt218rFUMqq0TOt//zxC8ZmVlPoC71UL1IyFxWRwu+
hsD0pKr3uRypshSeUn0LTtIL9Dd7s1fBSKsLGTS6vy8LqKN7PXV/rRmUS6XFm7fi2sHu4E5BoLMd
hxfCZoJQPVircqOmPZhWlD/5N6xp/1jf3HuU/YwPIW8tTc3jhsoRFn0aTgNd/aWz5IPY6fJaAlIc
1axd+ix9/mrOuB+cFr0SnBHpV5dRd0/LT6SCGZweVeIoQvnAvlkfLQM5eBELOopFoHQ/9kYSJuQp
E1daUleh+SI8oJE2r2sNZPg+1JWP7Ovak1VfWjMgVypJtaGKaDmAzMeyia38gQMDb3tEc4jhczf4
zgq56RvhkqMsWwEQi66ufPyHkdbKeJmAukl204/VVrJp9XJbqGfJTgnsRpVKqTe/U5gYhf8ctbfe
Uj9PTjnCeIB7A4JYKOzu15wevsrngwh5g4/FLplJrhJZixkioc129SHyFmx0lfQ4O75NE0Z0UUC/
1vPsyFkvwwGR13/xQKfxFQGvOGne6rWAFa4sr2BvPH6g0AldoowpVs4Efy2oWy2LqpQsUPBxVv0G
nC5EzRWm0RZQcDVAYXKdDK7l8yoGxKXpd7SkpIAd7+rVoCHOaGV6xEvIdxk5988J/iA9Y5nwsVLS
abY/VmstVnTFpShCfSbG0xwpNVTmrg3dqYQfNfr7LgOvefQPcvSTmdm7COwB3VrHbUSZFaXFuRqW
RICMoMXN/SSnlLYOdn5M12sC++0f/W8tPL7cFd8q2Vx5A+r/dvRRXgXvZRogiisBR5Q7lch2SkD+
Op4DeRF1uC5e4aposdtLSWlycyebACQ2dED73L48m7YGK6m0Nke8yFU/a440JbxCGpCpxeTbdZ4l
66yn26GGpRT/+IuON0GsOuBmYUi7I+TpeFIzKynuI1KLi/Q1cndkDeqboWuVqMc+6pzEDzxlZZaF
MzgEc0orlioZxbh1Ze/b6abIUKDefSDBuZdDheqgvvqNwUz4ziYGMVLygmGilXeVqPIWCGzqATu3
rjwdnoGyq+djZsytsyjb5DU2QQByuJeSqepL7JE1h4fZ0J07atQ8wAcrBlKZowo4gEkEWaoUkM9G
HP1WHKWtCu3q32kxkH5E7awmMdTPllHpb5f4joM8vvHLYAS3fzlJk3nGSR/5829cPI7T4apbOA0j
z7HVjWmdgI+LJ5ctS8NaF2aiC7FJvj0r565OIDPerJEWNWLi7V1sDlG4tSnMpKHfcgFB5NCoElBe
hkhQagH8/R+3YSG6KmRx37mIgRln4St6sqSnbLpqpu2HZkGDl3n6Y2sI8XTH+XNvFQK8NdYOI7Wa
ZOKZx0r9+SPCB0cACb3LjGI3/l0NvlActeuOlA/OGSyA9vNo3elWDxaQ13mjWoKZBHdXH76OoAyz
Hd6ZgywNKPKQgjRSGMKGyWh/qJYDd0cJdz/Ne/rWVoARcJaAVKIoOsMHZdAhxkGb5Qwo/zUMmNY/
RxSsk8bBSW7ebQQfVSr3Lt3Wfkk+1PhU5E/dRuJaiTyh8X9j6YWAO+UVTjBMXLcTH4MyLo7Hk6Lg
8x4gz7fkieaXiBsuXuHP+paOBc4zMriYLHGx8p66NC3nbeGaO9s3zNFCDs7loHVFVrv8NlcELf3Q
sG7ZWVykt2JoUq/nVpZE1kLmWvliWNWv4mRSJp6F2Bxa/tc+2DNhS9IuGwYKTQIHdiqAetwiKj46
eMYEhBsaG9JwIqvduQ1KONb/1mEVuNVPyWupHxPp/L4840QifzlVicZndOD1BVegQ6pV6ajDAKrO
RcmUU98KkhbvTxhRf7rbPhbiLE0yeX4wy7T+5iKgFcvHwSSHDRKa3kPE/UCYcOGsc/dL7fZYlFEM
ep65uzO9DlD3ZClvh6LZSsytvvbrNS9z0qW7GjMFUJRj8m+5dJqOZSJ9KE+pDs07IYZmNZ3F7qyh
OU3QtoskWX/a9k5t6/71iVfFbea2W6ThI8vV7nR++cDf3BdKDCjOT8wR/5dSeLe01NL+vKkDEmL3
qwNfc0qfYXHzBtei4kFvhNvfTIJVB5882J8GTcwEftR/hbhVUXq4681BGtmYrrQNfM3TrDQX99Vj
eVUBXYiTtzrCgCHJEwYlbmnOIsPJvyELgSjInL3DsuQUC1u9rg43xN3aXzr1ALx2C5+Pbmkkjd/r
wBNtZuoo8fqd+Fd5j51LR/SoVLunhJIu5txW8sZT+Mz5PMDweHvSzcyjD7ZN1MjlNGJFiGgjX0uY
jwHNWnM4r1Z2GMnYBVDFrfEXkOcCn1cJnNeUm4ubYz4zQKQttte4oWJShGd1PQdWRH/3mPk/8kGp
PJpBccO/NMzmpz+OcUPsrQXUAeVLPcbUZgLRwz7oqOHjVrxgM9HBCp4yKEoPrFArXnzWfSZu4bYH
VEd7QG4xMbbU4mxsSpWuTy6c1fu+/fkucot/Rr40WWd8fj6qzyTxWi8tn894Z89knV09XHddqyG3
r4Xzz7G/lQVaqPe88DTpG8JAUrBl/QkEvJgpfEW27z1aWHCnJExyJffDcomIMJuuWqtwlt/BX2GL
v0qEISGnikmDNwLkoe1PdXpUvSTtE/BPTljJhykeXNy5vbjNcNmp7Kv5ixXj8YqWaZuPmtuNxWjm
hVeQLBreKDMmNeMkFuSc6ZJsIDfBgKJ7k/SOcje+nkFXmChtuNBIb9Gg3Vt4i0pkmGJhNXrrgFkP
RwKhBDSpO4a2vYlT676t1rOifk/z4pDldYp4J5QCOU2haxYC1TLr74APc97zJoOnI5my3f4vsgmF
7WrVCH7B89xGiivoertSSBXiWAajAXFy2TOKUyc+e+pAENygCGEyzWZzs21rWFEUskusry6FQ28t
of3++pM01nzZTyzZJW9Km961twgXRh5UrN3BRHLKSJiiw6cBl7vQLMBRbzZU+o+ZFcLef75742eJ
8wv3NOMW1QKsPQmKcbS0qEgtTfDnnmpvtVuo5WZkGgsdHmKeRUvixSKLXVXR3kqETD9Py1+/DdEt
ekjwJtZUCS/6tIRqETn61+a14L7+HOypZoLhBQ7sICeoPMqT1Mdq5wJBNXvlF5dZ7YQZZOjbLrB6
y+Dbqb51dQcf/Bmar1MzIcT11ZY4OpD/DYZ57ZcJ9GJrK3EZDJ3H1rUh6rLTTXUC8V+hg8nFZhmg
WCvMzPQ7HTGYg7e/klvuYp4XSFns42LWaABCLFqcqz4cED6ZtVbJU8Z6WxHu/p3+7ypS4hD5yEYl
hMsqLKHP/MIcbr/Odwvdb8olEVkVW0GmHgsceTZp4Sno6DsvZFrGtWfjGl1w8Po2N3WE346SJOKO
qX2T4peYpIxDeQ7lyLIwPEQ6RQdeiU23vaA7pYbXWNNLNNI8TfbmNILNCpELtIO1yCy5iTVGpBIv
5G57BJ0dtStD5arcc979mLkKk7OizLcDsCN92D+Gl4gITz382hau0AVEtoAC0Q4vZ+aC0HM8kHOQ
H2UUR6HGl8iJeTBEi09qp4ai8pzU4UqH+AEbU2lDE0SBsYONVfhfMHdL5VPM7SEaZrd6yMujN91g
ajOpA1k8MmXFfNXXrm97e71bqyTvGbow9rgrvUkFVV3qD4RxRiEDBsS2RsQbn9FMClv1Odl3H9uQ
c2o6n5EyzDRHDG5TIqdO33muDj401SNfU3CsNeVckFhZRAINqUny5BowFOT5CuVR0q/W2rzvS7Fo
N/Er2PVG2Ikj5z+dmq8fR2D/VSpx9kM4dDh2p+2N8f4kr2nfNpk05Na8pCvxjqiPZHKyEEw9WUP1
VWQLW/MedE9L4CNjv/JbTlmGsA0ZKoq7qwwXtbvAOJMZJf0pyj1QbAc+NOYC9JL3a5R5ZtipTorR
Xa57/H+BVnC7tv5/aXgqRm1zLAMTKxSdldwcQ6Z6+mkX+42wk+l7esAxT3J8y3Kak3nWMY6+VP1c
6SrXqrJsPWZu4Q5dUFBs4KDMxLaILxAxdWvGkKx1mbxhgavXlW9SRs7pGuqIkmRix3bfV2bsbM/5
nurNsGuQ7VM9oVMWG2gkkjOGcQ8jTbeeHESTP3YUAaLUwPRWkjyjoMPzPi7RYtbB9sQslq9kOcm/
qPLN/he8idyuONWCRe4x8VAb8+0ZamqdYt2e1v+UmBH4/nfDXB0vgUobnNds/auvyIGQTadQ5Cfz
5YjLq/KXEI8r7XZUhkkOC3zoSwIS5iTBOqQPEdMsYNm5xG5GVAp0jiB5IyAfKBRCNRU8e0RrkoVK
4R9tSK7smghCuV5wbwyheWCzhv2hyojgK3UY9jL3kiUvEuS9vRZ2Zs0bW0cOg+iS3fmcj4DV0/D4
PEi4z+vnuCtez2APJGvARnQGTgjebOqKebV0fd7lxT9qxOeOBLRSPIg2/EcqOf+KIaNy7Ty8mYNp
wRpOj5kxOwhAdGd0nnCR38iYhEouMbo8s1GtT4k/lgnFMotnXCfYfOkYgl2t0Uj40UqEnRMrcrFl
UTFfxNX1/JXUoGo8QwYDhPHjjgzKRDaxuepXSV5fV+7luyfHMFAe8p91lRVIrEqlfuu1yDo5YOn3
Wtq0xkY6Ic8Eg/GhzNQbG668o2qFUHH63eU7GURHhUolw8737nWTEsIVLw1B40uRHzLg34WeO9Wm
4NaX2cLNsKkHPHg5P84xRmLmY0FLH9IA7b4rirZ76ftYTJA1IR4c1G9brZXfXm0N9ZoiVsf87P6k
DBqz6E2FhSnMnkr4/5WZsbOQZG1VVb+EEc3yaWILVfG5URl7TnqO8CDkFddRKQnDliem6MLwVK70
uZBWANHDtjFebP0CY8wBkFu6KKXC5OMgmohT4DhyeO9VzlOrn21xwkajec7Itf0MQRjGmOSbd731
QL6TCbQoJmQLwvxndS0EKynJ5QTLyKuAJoHQCxh0+vS0zr1l8i+2gHiZQQNPBqypXLzbkN/YOV5O
qiZuHYg/fHD87/i3AbB7bbKGZytp+h7VCbnr/8JtoYQSPf5Gc23lFos/Bs2DMSdLDZSoUaztKNme
jGoPTx4S1jfA4MisY1rcj4HKdxJbt4PK4lZzim0VdD9AEDYuGyMtTWgR88QpE1IjXW6eySKWcoU3
2l4ifSCVYWel7jxHHfepfi0JZoUqIPHEAkuaqyi4TVVZ6PhikiUMb2ZvzIgP28s+j+w+P82u6IRO
ZitmGYSDWt6QoYBzo2vp1zNi7MiTZfpHEF810oEBvT6SRuVvnZ0pW8C3C5JNJNims9HPy1f/VI04
1sfwp9wtavrw9tRK6RYWLz5xnb2jKMhdz4gWHkAIClx7TnoDxll0emaHiKAWWi1701wv85egsIlS
BLNN/ewDmla0mkggFo4LrfLEZF1tud8rvR9L7E+7jVtvqtJADMFgT5TTlbrYqhU7TVU5KTXxtShi
0Hr967mJ1yg5cy3IsWLsMrKvwLfTMp7WlsTbX6uPQczdLEMedKPnLWEMG61JYN9HPHkX/aga3417
018lnEtC7MdOYKc0mXuodYT+eoH9RzWzcH3RBqoQFrtvq528kQjwxLu7klFuqz6CJL3t55nTVq4K
20EPtB8RW5U8rE9CMEUM0/EBHrw6MSzJTO5pOVPHm+jLYAg0a8gVVtaNLMj8zcqoHVUyGvgK/6dN
jhIVQLU3xPSrSvbI8H4pygHgclsyZs88BQxjCzndpirWtolNgplo+2RWlrEofupG7ArleE6ldvoq
kKJ3PQQn1UBakIFlGFfk+VZ+ab5a6KxIXDQtrzVV9DZO4UcKgP4SPaNxqeZnQjx9bkpE5W/05Q+k
faIoikhFYVkMl+xJn1WVTfl4lxiTbQam7+lm/X6Pgg8cZ5/Nm65hSbUBcepNtjdPT+KmAEs9zZyf
2svs63S1/U7YiG5+g/XQdKLLct1SoA3YOcN4vCu+I89Z2giZL6o6Q72CcGCQl33Pu+xTMuYavetE
I5id0HlrxRbeCpSZb/wnJiMY0bP++2Zr1084UKbVbPIMMYthj7QbRnvYfsn/xG48nBHxefAUzL6Y
l8LDYOa82UHH3mMaEzkhemad0ka0DgUtvr2l0aHicSktl5wx03DHTlCrn5XEs/QR7ZQWid2pgDTg
D3a9APiwRlUG2EVdjm/AVNk7aAWptaHqL42+YxKtrt8gI/fKEswzl0jFEFeRPerRPMmkUeIPJawP
pGxIJbRe5l193nrA7nYxpmipJx/fo38rIXE8aXHp9JjaPO0GOtPF7jekquWEoNrdOpb17y8yV/Dt
MRblMGgyt4eP0UTxPmVaPXoBvYThkdJEZZiTUiImIZr6we//zYeYXVBcBcvVtrW4bNP54uipQevO
V/e900c5vyQTlBIn/PzIGPRnRJqPF4njDQU9GVE+s09rYz7PZqU0KqQPuxkzXQRTG+YW/HhCMdiz
n8guy9C+qxfVbSLXJ2NUfrtoRBblO2+nE56Ck5IsBO2r6Bd0+9/aHjeUIaUyvyOPRxXAkzLiZopE
nHSXu+H+WTQnyUfSzRtxh5yvZH2/xT4ctjhU1jbM9WSB5WMxso+zN8aeuEDCm4EtO01jXPf2QrdM
JMnvOSwqRP4FK6EP18yzc4Y214XhJxqiaCRPhpoCJPjuGY2SC4IGsWVZvutRWApFxyxZAdr4IW+2
E7+v+Wqa1tPY7snbVO4v4t6iSqd4MUTNGqj2JVhwWGAnebt+B2CEgE7Igo+RQnfNqd4j+47YYadN
ZCU+3edejRP36uaD7azfA9H2s8i6mO7P0HBleRmv6M1i3xS1oqnWnsKWwN0kRhuppZap96/J+9th
PiJCZfGHM8olKMzMdzOqZMTVQ7LOFJufkgNvusqvkuLSHjAftInprZh2YmcpxyAop3Kz9zzSLMaR
5uORqj6bI3ocy08X7r7CoeG0B0FM2omhiIz4l6GMTDI/x1GN/Nlxov5WfLvIjWXOpRJr28Vf1jw+
9dsz+o0JUrujbdX8cd4plrQy26ZC42gK1BKJk0xwTGx8ZMMaK425OXuLLwhIx6jHMNS7F7pWrzvS
A0YfDDvPKiqal+8dIGIBLKU5KkaZ03OETURHTE3Lg6W7SCuRcZ4HItep2vR3C892S9JX5khcoWKf
ZvjzAjwMFPNvBZmsBf0zMQ1KSNLhatXSI2bRr2NlwIo+qkJU+C06+eGg2pJBgxjD3dfJUddMtE9C
J7cXCLsHqvLuL0Xd/ctXwq7Weoe7GxuJe+06MF7zGggPzbyoXDXfngwF5f8yffCjyFGUzqj71p/a
ak/FWhlyEyFVYGDi67D3PQaGWLuAnqCgOYweSRtOX1z5KivCGe2KDCGU3HB0H5kDhLz+qLCBWtQX
EmmHXrMEA8YzKdb8PHw4T/EMnq/gJPvoKF0YhVqRQNPBAW9GepSlZIh2AqwPFbJWLa3mfzFfUl8f
VNfmOw38sQhLKgDttQqRNDjxhKJ0WQX4/fQegzCvGJSFadYcNniXsQ7oVfKdMmieX/irpBcewJIa
+EQL9MRtj6LqcSD6WiNuTq912J47e65SjAuLo/x5rH3QjHxIDQifIKph/oeIlCvDRRvv4Vntowew
RHoVERy+c7oy2DbimHYy8/W0ZgMaubRPSm4gopnRauzWgo1Ujd4kVrpvrXDj2y7AQFZbk39l+7AB
HBlW5b4M3IuJhow6OhhRJPG+7jvxjCIIHU0R2wXt50xmNsCebI+fFBLXSwtSDLaHghSpP+zjoLke
CcyUUnqPDrQMyax7F1/mE7g8QCKs4aUrPoyGwaLq+fs/fSXyGSVPqJuBGbisupf1wtEvfMujegFJ
X5384qqI83ZeNETP1JOJCHBxo7sZulLy98+MoAw7jsTJu9tE3qyFSFlx60BPp1RXd7rRV0MfsEiP
MmbaXokP+9yFcONWr24QkUbC/5AELtc3+IYVlb71JH5JcCcbWGt0JQw1Fh49UyJTz4td6YdYiU1D
Ux38EC+8i8zjCtluSyZv5RaUOSPYZjxg9yyeQM4QT6tYCIya7Iml1IW5YWW02zRFr22tfCqdfPNK
hUkAz+DxRDg4qCj5NjfpYYzYjMYBlvs1TQDHKy/Dyy03qcPkWp6V1dGZYAUNmQ1CkbeVhswI3Zid
pRqhXK7iiiTGuK4HstZvMfKwLlvDo7eU9VOAYk8dykbpZ/p7w/94NIjxwsbQy6VUokA2liLrzOUk
ex+wCdHEzk66lez9D3nT0n+zopoU6UM8Gh4ZRItqrhpVamOdfgCqSNISosm4HJ94dWEX6KYgqzOt
t6BA24hfX2AvH3lf4jX/usZ5Sidkvcx/Us9j+keUCz9ZiPB9I0pfLnjpl0kUh3irOG8out6m7VGb
Xwn5GtpwGVqj36HYvyybJuOl6588qg3gAUOs08LqoZYZuPZmbCb+/PxBkvXnNFU35XcVrukULpqm
uJIal9UWwgg8Q0PBiHxWavmtS+5wSg0Z7Ap/owaUxIMO1XhA5WcdCidPEKZJ0LbdABAaYKUdyF/E
eqILM88Za6dt+onoibnQk/8AVNJq1NlOyuD2l4kVXHZExJS3Tkkgb0bQUgh7Z7/9eodlSdf5qS8g
LyYlSUJDB/bzbt4/zzaGYz50OooaXovQrbKK6cvfTQjZqw2BFiUOQtkM+cegccWLY3b1Wcyw5EOU
r4ubjB07RJMiZHbBOgue6Yv/m5QtWTwKjn8wyr6L6VFcEQSajG/XAgOx344mOKLNTcGJU3E6Qh+I
ngy0LGpw/x1k1HD616+qaklT7Oengv9Rd1hlw+dix+cKyrDDbFL+HyfcJ2zJnQIWxPc6U3tifef/
OzTbctqEv6F9kv1NG7qG10jcxOt0NiXjhu776t2SlqGBzSvcbZfPgik+mP/nUUIvZsheNFbE1hjH
Z7Kge/hi442ka/FFx8sLlcHH+FK+gO4PGVqtR7BRVu3YVNy1BCpfK9yb1kBaA0ZDpVfP4rWmaSii
Olqs22+SjqdSC1HwK3ZrqoJgn1Z1UW+muH71BB7McrakkVh+d/YXetdLj0qgnrz00+3sxCrsUIO+
iGTmj3laRutydBTG2Z2jCsEzAjZKOfhWJ78UYEjYWlL/aiRbpj4I7Ch6J0YVzcYBzx/yKVVI8nmY
VTtCJTYFlFBpCAH0s5RUTBl1tGJ1RceqdUG37C2e9bF0Y3+vUbVEgsGsou+uK8+zTAQDbzFjb7c+
ngEWsRwl2v57P/vpK79GY6PbrevJcYz/KE4qNdFOhEEcms2FGeH85ZRYWxzhsrb4n6vTJNoHV0fo
9/mSJbcaUgXaolvBrx8QDdxwUYMKfC2yEDPW40Zs06UpPUNq6UkyeBpGzzFEksCE/y0H+OSxmMPV
SfqoPiQO+i0h5CowbG5UnCrTc1/GOmTqi9KlXj00rIP53of6gahwvrFqhf7vkBLHF5LwrfjXWLQi
68ySGQRqrLLP3Vv0tGnbchqOa1fYmTnatRvfZ59orTPLlNMTDwusG9huMr7xX9tV0YIi1QHgpjbF
r7prCC673aJZGsaB/5MtoHuE55i1NspNNDR5knpjmh2cbS/sDO3sHDOd7b2rcBV6S5o16IZdbuqu
Fw2mVFlAg+P/ALutTcc8jX5DcyOnEp0CMYSzw3KlTVNiG/1Z0pnK04sUgW6qOR7he6N4fstgMaOG
Ha4oFJH20K75MB+nZOQ0AnxIQoSxgwhANzZSIcm8b7aDkxACTldS4vASTaVhyqVPldu7irZwxOaG
9XFF2yeqbaDQ3YHbVJy+RiphPcNDb3dCgCCKoeShdTBKiv0z6coOzS3WFVrTlshuDZSwUmcRWFGv
swnrJWX7xB6BF6Rru2s1ToPAMc5zHV49EB/smPPX7etOv08eOsI32MA/YtPUhnwBHpvYaZ2WipOf
MzbgkNcpCpdo8rSJcP6Sxed4z5r0b6qSJL+/v2YREt1UCroKln07hO8tFhieuMvHUNaAXKl2XR6T
k2XZt1oUokaD4lKXQemFXV2O3sNq2w/fNYJn49j1deGuBztZ9JJH3IX129EM7ZRYxvRzeHqThRCu
rJc3uNNTLpBMPRm6SCOTLGS1wgJ0LMqB3oWLk1VaAd1QcpoomWv9Pn1K1uztkLSzOKVgurrijAD9
hxchYDf41NHYzB7/EiZBXWFS8QAiWupnO9Ug7zLlaniOQPSwC88pg8EgebWcCJq+Dx60iUZNlira
sx+qCNYb5JgMksNVa2M8LvW2C+TsFjT0uGdkcfzE2c7+EzraI5Duq7RbI06IstaTRK3zgfiVLrgK
SeXLTe8xYGX+iSWSi6hAcTaRHEyol8tAr6UZWWjCZyOzghHNqlPoRWa0l2cx+20FTnP2j3QqwzI0
9FmNuFVxYhP8cvWmZsb3PFb8VJnmdeygu6F4rFaB5sHQypAMyUFZpqX1eO5vgGkhD++5lEtdlATR
ivdVk+FgIC0EjwHoysfGdOdOUbtSosWjU2XPYOOF/vVCTf6jlEuqdW08y3zKHg9NstIhpGqAAu7v
PuWwRWAqWq14g9JzbA2zj/9yXbi8bQOSiwqIg9o1t05bISWS458U5lqDM+z7xCfxj/KvZmPSkKkq
XhFgcl31qRKcqKRcNIio2g0R+/S5QI9aEUJpPXmAovTUSyDOLjtT5AQ0okGkzn5spalu7HN24N8M
eMT69jGEyr4GI3juz5JU/PJ2vpsIEZ1fYg8gHv+/6D3HfCZ3G5hlPsMw0JTTJWsNjUrknfAxYA7I
W/6oep447VhO/w/JGl3QJawtT4aEcsUkgXDjIgaH66oJfIeJez+W6XbaQW8GB7ylJX4J8//B3y1W
ntHyz1mgfDaLBGJz06zXXFsk4A3WnQ8LXW4raWQV/n4WiojVjJmyJnxdOFBIcZivjACm2/0Un1sM
N2v9Ru8XnZVfZWLr0RMn1NG7fXTMdPt+LWJO628SVqwh4Ey7aXYvWW1nRqHZFP+OdY+2589X5ZgG
zwvhO585CJP69EbDPifvbLb3qYxuLP8jnk7fR41fxj9cknrnZKWfaLvMG0cFx3An8ZXCR4+CwaBp
tf0bh2j54TshPNdcZUVkFx4qgQ26l/uW8Q1JWLz92VHmnd8cbSzzkOvSBHY1IesmOI54BRVHwYZk
gHOMAbmKL3/c9iaf87DY9uR/qBIijNyKSrHOpZDh4Yz5vmSSLScOPg18ym9jD5C1h0TYdaN9x1fy
SZnKnU7N+ujNnHyeNNLaeIF4IHsmxXSN3W0Vnx3e7Ue7H2y7c6ipjEaGYVZx32Y+Jy7Lgy9IQ82Q
IPYYXjpO4Yfz82uJwBplSmG0/15aorFdaFPPIUrXHoj+HW4/kWMXUd1D8BVCU27POras+S9c8dGa
0GlmZESrjpSr27XunloEfkziBMv1/3PgFaeQSwUjT13T4LrUEouEmE1uT8eiDPUcJjbh3LmWpReZ
hj0lsoYm77aNDiKOGYhIQiXEl7rZG/iJ139meAa/z/rrxfZDxSPteqQFJg56PiDz6Atj02c0Kiz8
ll3E6qEBDKQTl/B/54dk6ULuOJH9tIYUY+uHRln6T0b/RREKiPolFaUydHBRhPYrZrLV1Q10U2JQ
9qED6LO4Bx/WoYZc4r5ADEwOhxPtELmDF74Dp7HvLsJTxabmeX5vIf25hJa8kJRj1UbDI6zPeio+
UqNSdoeOPZGaALiWBdcPNkLZl9fRmvtPdVJ9hbDojnoygX2XkY1d9biTDhm2yVmOzR0hGCneGvGo
+qX/NG/iuI5JWz9yn7h80YYZxdKZdLpzXTix3+fCVWec6R1n1SGdT3naZ9qwjLWS5Qx3M4kerykM
Rpc3sv7lDEcUfNwYrH0h1IEmp7JqO4h3GaNxM8wzW+Km8xyIuoh/LrceSqbP00afHd92JK2QhN7A
kW0sWif+948ad6Ko2oYcIaLSfFVCYLMLemhe3bonhGXS41zmJflPmuO1qjQkIrvhHJBzE/ZrMduL
YWIq1hWY0a7RjB4P7TG/X0stDZRVTCQZixhTxqAk4mIclv7tbCDxgmZlG4GIFv0eq59mOWqsH/B+
/uleMTQtP1Npq0Y+atCjffEUMzPbQRRse5UV0sSYymCa1oWKL/oNx5Kx5fE2gcgqGYUFPksCtoz7
wTWJd6uqFcSJ8YP38aij/k3i0k0cqDwWMdks8k5aqAJtud48D79q3qpKSg+lzGLLWkwosT919XFo
lTUoC0qEE5I9cukyCqkyHs0SIW10rrgWSnJFyQK5FTTJQZe/Cb9xcg/JJXYgoVcoHU8Ug6WDEoCn
2mmdILJNodihQBxNKUZt0OVDHUfXEf2zF/U5i4lyLDNyY48EV/4jLvZNUHEv2Eo4p55PDYhIAmiw
fcS+eX98txsYMHbN1avLkHAVnH7I5w5fFBPlSlszw67MtG5O3ZAaoys8K0Ltki4G+FHpra3toayX
z4pCIXlgMsleEFgVfuCiAw5uit/tQeGqi3cFGmZejHSYAE0wVVpdOCRjs/1HXoFdnjJOa4vqEtmj
2c44UusZSVGRlcdcYIh3e4OaUmvLuDucqapt5QIDqjKdNDZd2l+UuMAedEZWoSdXGgDjoO0mTCCm
TC+rksWSc4mct+GKrP8i2VwE8sHj0JX0zds6fHMbjQ75xap+2UPOQgTS0g6gdvznHWkFnK6RNyuR
LOhRVgh3VBaLWcCkXqPws4foRk5n0Goq1JDXko76Q/XhM35JH04J2souMiYKk/UNJfUMEqRkWvdI
Eifk6kz8KezD+P6H0r5G47ZC2Aa2rT4gZbDNNZW3m0bpwItnXmFGLxpaqfEpo/skZxyOCUdVgsPa
2gaqmS07zrMiiANg/3GDFxEaNmTlcKDa8s3lV7kxExjZkqvfGoBL00V688HDa65MpmZoHo7FcGR4
EDcnTRA0zgK43eplv0MHc9tbT0TJkQDd5gslbjqSE9bFB01v9e7u7rA1X21CX210pthmXkWHng99
oG+8avPpRCnBxgZ3XuO+Qcg9Vk0AS6JxDH4IPDthXqqckSARgAEz9OGCwNDV11Bm3B5kf2s/6YcY
35yZGeNZtODOTugHqQN1DbRcVAWNen5afqP4BWEv5zk1zgBSpE4ygtLYt34ZUr7Tr9W5djZWYHG0
nDlQsozRU079AO90GQBbaWDr2tgfLTZMpR6xbeCD3/ihNFtLajQTyjWk9F19JuMUAWJAYuv6z4fN
gXY7PzOs72WxaXiawLKhAsgznwkHyO61R6D6ZcOZ09Km1y/FN6n7DaykihzqEo0OJ+RW/Npi27+t
gNAycR39HfaWbcly3Aoscu/IgQoigH+NNNO3tTw/0Rk9ihJAfFvKf9dn6hCrAIW3EKHsJNG0d8vK
2uCzqph/c1HPp7zYnrKRqrVWvlDoYp4pNOBBuyc1dwuKTLskJBgERNPerlpLXL679DJlPSd8UnUx
/tJ3pupW2B/6D7ZgP4fD+QuRoEolfshFew9wupsk+K2RqP0r9WWUgj0+tFX95cAi2anwQFOdGnHY
YMqvKcneU8Qw2eZ1H0vKoXzE6N6OHUvoNAz8hbfq/Tz12rb31kZRj+AM5ZuVARE6jH97zodzZN+A
cMZQy0eDHzqlEEEznt+Tky0kaNSwyvSlNpigHyxQVn6S6BXHRyXCwtaj2lH83lIiJZjZYVtZ5bO0
YzDLN9GFaBHbY1mvfmbv2tXY4GqBd7d5ichVyR8axh4TjS4j5O0ALFSIMLZ9lpmZq6dDYAL649bp
SSfA1SQcxOT8QGDikSWd7kWhHezWEvg9tPxZF7RbzT+zcsBiCFQyL10i3J+YdNbiCBS5RJ+7U4BS
iLcjskhleTdu9HeGsBqb3KpWY3flq+qzUaB9flZG9FPdi5pKGz8L6woS1C5VODNShoYMHv51ISvB
0/vqiEpo6i5uRUW/ii5TFrATHSj7aHR0lmS3Gnms648vr+eilhWc/PbdXjfZtHaCFtlr4mvgQ+9w
rSIOQ4pUaKZ2d7HNk4OnZu7E1Zx6X0q0dYmOonl3WCvVK8RMBKFvaLAVcGJUJyGOyNtX9bj18zm+
2+oGg3geRuQuT/rbhWjcYbah882ga8FCA+O5ytEXP57TgMrRlyA1SlctbDaE0W43XJtWS3wSDcMT
rWXX0LS6KPTC+xC/arCKBEUHlzOLstWANQ5ev/8PV2jebXhpy50pW5Pb9kXg/1eoN9BULhX0ojNo
SxZaOkuOXVPQfVVmOVsnL+FXBe8PxXuQnRo61sW0MsUCyqFe7TCFRbHxPuI+tU7r1mRsu39QZmYS
mgGLlT3I6X+H32uNcSEpwY9LCgk3tEK79V+2V0EbKAvhJB/x4Kfb12Q89ET4XMF7QytWEYL81MG+
7HYuriLUO2oXsb/IR5qxoHNbG3pxBJI20h0Ybz3+M88iAwSsQpq8H4Wo6AbVMHNms7vMJZbYArs8
tZaJpy9QFqBqPsrYPi2jD84nDBnfsEUFhx31LHJtKZ4U1D5GQPGOBUcvEe8LPGfMl4UDauLyI+Zy
Ou6X5hbeddRlBzZKGrN2fxxiFKKuAHIiNdPZzdG2Bf7ruVW9NI4sHBEtry1+rJIE8nvf9LO8jBmi
zQGM7f18AwKmAvleONhp4g6IlxuBQuT7pyDuk5EgLuWAgC94X/DL6dgQlcG/ZOAZIsBiwHqTwrXy
36xd64pZqM6BxF5X/u1r8yTeMQhKIt+5/jXNDD+kw8+gy94wuxo/dGqQFjRucZNTouFSZwHv4Cdg
/ecR8IULGrSW94UQ4VSb9kICLFKHKyV4ltyAFAfXtM+XNKRHJYJFPTlxSoHkhqKXFTxZdO2OSBRr
kqCOrAbWMCzcSdNgpLXTIkub7TsAaTEbKCN3v0uD8ZzaKc+czYd2X9TSWrU8nbeXZ2PcGRFNDyC4
XdXTErLfRAcB/vsRl5JLlX2pdqcmFnEWz5w0q3E7hpAtELbmAzUvYH1benXzZR/455L4CtG3Bf+7
7o7lnuu2fk+qW9GODagTl9MuxJmrctA6YlgaNK4wwl8XIxJny02SKB50mDwKFvAklqVLHQSYMXIT
Dm652FongkDgqIt0Q4DUZ3DS7nk2s9k4vmj3KUgGCJZ9m7fRKy5yf8PWnIds6gwBF9+kxFIqlSaz
X8lZl8FXqhgq2lNU1+6FgeJ/x0pB9NaUu1q6EHMhsr29Gvr8htjn0e5b6UnLvKE9XwtVAb75zHc9
hjMbI31m5ZfmR1oBTJrjVfymVy466ZucCpCRR4zqBvD32FFhoZf51RYYz+PRDih4+cjomrWa9B5U
ufer2naEyYG+394y8+AjtNdJzGrBEaD4K77GOFJDxWU2BFG06bpKVAf78ZHUAa9TbFByiV5gvV19
FKGjdSNllLQwcbSF1ojiJbmR4xZsle/M4DvzDmtc2nhPL8rrjEfViETh6jNVVPnPZtBGv8Qdrh/S
n/zxNhc8fZVIUKAfJpa7W8qZQvxida5Tn7/HoVArcVvb/5RzjRnE8oPARGgnjbIu5bXvlrX/XGCZ
Cm4Y07L0ABVzEtrS6iPS6/zNWLcjS4LdYH1uzuhSOi8cCAuHVXjTpr3OlRa98+pUpbcpjD0/MEOp
tAvtf8Ba/LLj55a28B0Mz3DY3mn7c3WKJsUIoQUqKi8jQVlCHjJkTSQNuNXAKSQ0eYuQUhlkbvtO
4sxMEN5chFtAiiVq8NYppjxHz6wADxTFaWasqMy5wO5kKi1+QC2DQTNINQMIVLlQgD0M18Dqay92
n5f4G/dzf0Hon5cWbOxfY6RfT3Xvc7o7ZNUNqbCEoRjsJSPZ0LY9ZCj8iGGpP1XU41/O5luqa/qE
vrLtf8AEYlqWiUGnc98IyCX64Ko7UbBabSP+AWeRMKUmcgWjxwDl4v0w5uhbv0O2hC/l3RtZT6aL
MzI0bCIdUHvuOO9v3puzQwBd3mk4yUDXBfYM23Cgmuv8EJ4/TlyoEU4BQMHTaCqWGGJLff1b7fB7
E2/oR9S8uQYzBBeGf5D2y69NguSCOinghSzK7kMPOEK8YZf+MX5Rmnwl2Cotr/rjJSy3WaY06k32
mj99divDWLn4NH0h+dzRRTul1xmauwTF9iTnXv4viF54mDG1K4Fc3B4y7ZBjRLyAIBY6WDqvZAmc
Ub2YUjcthTCGh28sONs/BpW2LEWm6SZaawtP+UNl7ohJquhL4Z1Z55C+bkjW5Yn8QUaP0VYWf0Sm
0cNdbbjxBmIgo5eARm/wekYwND9oTXezVR2EbC8PtGml+JBnpyHhusjyrvISNlI6xxYaFHOSaq2c
+enfDxGFlg40hHTL69HK7VzqPS0vK+Ah46LFogaCoIZXb4ylW0uIevn+PHG6ACaaRE7TXaO1OBLT
aaSFEm59Wuv1zNAc3pUyIbx6c+jSUzqo3VjReEDt/IqQs3eizG3T+5AdcGsWcLu22bDmHP0I96lV
DU1QoMEEsQ3NKlrXibxbKUsCCnbzVpQUzXu1wKYlccodvBtLQwhoIhvr/dTqnwb56bgZXorS0D8e
OcZjn7uHf1DNo9O6JefiMbafWLxVEWwxCCatnGGcOGtFoQPkQiuNS5hzeLhEVIy7crtJtWWrX17v
6HloMbqVcPZjJM95+tu3vL/9Lkpz8RPEU2c0GcfFOiOAdelkX+fBwrzEgTdf8QzXNMuy7mz7tDvA
UqKNTCi63t4eS9RCn9aljWIS9K81daBktGA13RN15KRZ5UaC4/DqKvV0LaDOFJ0e/Pgx+s22ZqPq
1/55n8RXDVrMfiv2g2nv7Sx+Ze+e2zeuMExbUd3je9cGOzBmJ2SLarYs8Po4pNwVER/Hlti3PD9z
sBFduLXFIYie9S7c/dGQ+xnSE+/HftE2Zje3M0J+t0P3wA9MuSSE72jKV4gzSt6JV8d3LfcSZvMF
ecnIcgmFuctN+O5pho5Jgm99nMaP+605Rd5R25+42R5/wn3T6aNn+kNVivHx0EsrSomhFawhesSy
OH9MXLLiDpTu8oEE0DAGSPg2rA/fpkC2hVzMdXZS41/WnOvnrgcMJzZaJPBUCxCOSBrvQSztiUS9
pHajC89KpzNSYi84tWTSnyg99d6YH2X3wJjN4J2u2IcBmGRT+W4MD3cVCaSaiRv2970OsammkmlY
aMu3QYnP/hU2j2r9ICkNm5+rxIS1C+zKL49lO3o6p7rBBJ9sG6nTiyfmnXsBP6JDPHpKOYJs7zgg
hUOAHvQ7kAAXzX+4AGq+kicln5sLSuQpEpk0nEDUjPvOV033NeqnFIvdNkhFUgXHiBM6+ScH0lPR
LLswB2ZVkYV2r+IqMLkwT4UTVZTmumSBlYM7VtQHhYgyAKiIepOpL13UQUmIJKAFjQXgVSO+8vM/
0B4Sb2Dmk7yp7s/0jh6XV1lfvuLDSjYAmcBXJdXnW5+CumWTnQvRVhK8nLbBrbav+WPQT1c3ppDY
PP5Et+NFDZ6qPD7gpTNujZ/mngQId06tXc5GWQoC6TFN6Rc5WWyZfv2K7vNROgpVUrTFYJdIa/6p
yt+PEyOEV+0Wm3oEvkPRTKZYv3wDFICNRd+xyTGatTtevtKXq+XdUySNCVGwhMCXp7f950Yc7Ra/
E5JbjhpEmEt0+eZk5c8ev2QxLAqKl6w5YGUjwJybKavbrkC2c2Js8G39Lm6fmPehzrv+VoqPL56g
fGcgDhkzhAyg2y/5f3JFbJK0CMqFe9JZvPvBsVBL6vF9p0zpj2ARRFm3azYrx+J+oWLLhoreZJX0
DP5Se4DdjjJFQaJBuofjR4k9Oc1sKSjXQ4qD1E20mrnsMgLh4aSzMOz1IHTcKm7/Pdrwm9gvMIjZ
DiyLHsxHfl8zx2TChZyuTDxd8o6J1O1X6jrgu69jD0qqzxGyJa3eqi/ZmAcBv9Mvs+h39XBiYsye
woRf6eH8P2xdof6mC8wiV4eWS3aWiI4fyltytVooCrIRE7tVaM6UcbragthiBP2RDFUXPR8kQiy3
RTHkQ8v83knnAkxY8PZ2/8uJIcj5Pu+DZQOs3U3FM2+hDEiLsgbnsv/inRkHkSxDvKqR6Bpy8pSQ
Ez7BEWYsaLnP/HQW3tgZPL4UGcJTIv7gpQVAdzOLTLiyAJZRCTDjWqOeLqPZmJceitksSO9tx0xy
2/jy6kaU/WArgnF3syejmkdzcm1SZ35VktvHeBnONgpp0ccn5QYdOfYxa+bYQfyes170z/umQg3p
pSHQJjQDswB7xqGVYXAF/frisApC7G/ssPvKd5MLAJGD138sZNptw+iFWQS+dI6cygwjxNL5g2Zj
FzeA4OxKQ5SOI/f+7aJhgNSTg1MMB1FJZ0wMzJmgJL9a5AXxeaWHUXBxyI4PuiMHORM8hfx/6LtB
bRytbOom6Wac7fIXZ4uVTSH2nsLmLkGcYIxbZ8B0Daeq2t7JG52sgXdCxkLVxc92vjuavqQsjt1Q
u2DoERoAnLkhQ4wY7GifNs4jWx+wpQT6lOj9BwTpVEjhpLLC2anz8xm6OIRWSKLBRy/IHWGg9OUq
ceZnZ8ZcPYQHaY7Bwf9yKlDZVtQ3KyXbjX1I4MC3Sdv0cVpDAVbaEU5+gNkExwO6nR0pBQvAJITy
CRKVeVtFP7bEFLxyUXQKCaJtKHV479hXaNQq9B2ilqxPO4d72F/LNanlvdlDIywrh+QSIWFwqHAL
yBfP26n9O9pcHSHkk/bhPPTHDUFDZNEXI7clJql9s10y5BT0MkAZaMyiB68lxOgWDliL9mR2f6Ql
D7cybPnfpEE72sRujH0GMdIj5KzkQ1qKLYvMxvY8bgE4+bCsv4ScDgVfUXnh6DmQwEncxxs384kT
gBh1K7mUQu4KoPNL4W6oy2aNAGO/lH5fcZ4j+BHCd0a/o3oi+iqU10St9sGYhaDxosjCc2+/PPcj
b+q2unb6iPeXy5WfVxcuIliI6hYWT9LbNFQnYWz/pwWdSF+pmTYMbkThM9ZJiG6bcxOqr+Qaw2RP
WNjOCdJoXcX107HB6CJtaCE/TZbO9kGyI7iD3GzUWRDpzTmpTjHHVSYoWLdrrznr8JwL7DXe3DZg
pOguThX9B8bt7M1vPXAxusiFxDvQGABiHghZtx6rNIUlZwrtXW1pPZlVQhqvkhkU/x5QbPXhsoH0
SGl0NlMNgrGrTBKv4nPkcYQo3z2lfPpqtKl6UbCaWkcyR77oqexJhwAWaIIdKsrCIOwKyk54qn7x
b57affzfIhDHMK5GIjdiUdBISw2VQDrlu05dKwPEt6nY9JLbrxrXB7X3gsLBRDKDMxwh70LdOvKN
Xyi2+kCQkGSYvR1pdP5Bivpsbrj5s4K+HKOFZIJhC0wILSQRhEEgtB0JhVt7dFpoQHgG5UuXjKcf
cJp1F9xiErumIzQRO+OiAqrvpPXujWDw/vSC8Rz9dDywtA6YO0XKf2fmPSq2FBFSbrAVZLNF+hwL
LSgowmKK+3OUqfbR64JlzKSyS4bgrb4eN2iWFryFBNBR7+KUSk9AqmW+eyQowBY9/tZNWk3Ij7Q/
iFpniiJw++KgCBO9dnPtZ+1gAa55rNdOtSl2hLxAZcuXQ6jKFgh/pmc8SaAm0JzI7jEpbR9A2nAj
3e8OiATcHvMPi8deYwMY1WVKHc4NG2JG0EAW4fGtX27m3Mkcda3Ei+kicYYKswv4CaIKQhnkQzm0
5k5FRw1zlbpOeFS+Pi5uKgeMAN7e37VqZbBPi+fcJIno8SyxEMUGYpUd2frGwJ4XalP+A35NvCQO
AEi4laaV+8szEeO8XMAAtT8vxeXpM35j2sPf28EFaGqBCwipwBWcKtyWKYrk5yl7uG74it5PdPvJ
HHWeZUStTqAoV39nhz7rFPq6f7ZyB5G5Jcfc4fCzXqEX0p0wabcw+ApkAPd3oRrOGAdjbzwYaac8
X/PH689gEvZ6Con7cfU9054sZAXrRStcmHEzUZzLUXNO9mhCcq3CBni5mbxwxrFgZNmdRsgREt4M
L+lqFCMhhnBlbFJA7rQDzK/eaJl1OLAN6fGBDSe63ViDdBrxs/it9tE0oy5BJAgt8t4to1L7xYEN
z9Z3SQdMGol5jy0CwT84AZG+caJZ0ubAWXlr6KCB5y9CP4YNKGDOx4099L39T+By6tZy1CHlP4sp
B83tEJz8e5wCoV6/Iw4ulVb+mTke1gzHpaA0zzpdWF6Zj3Srszkzsj913q0XFhOx2IRg919gQnqW
kro6oPkg7bJMM9f1rrJIlm/hHNPcOrf8YaScRqOP78t2fbVwaBXFMevpVtXbEuMy6eDy9tVQlrQO
98aoU/qdCC0aESpRuFuQgt+aiaOw3biN8pd5ILQwyITU/834G1rK/zXMOYnfLYqmWTHqkq9Z12an
KgPH7fFWCXiNuE2XoSVQ3rTBmulzaWuyCFlotm1s/j3fNwxGUZX6qhWQtbBmZI/NGLlX4berTrDS
hmpkMbwc7hVCQbg24RgYpH1aX94w4dmfNWkgVBcETEvkXYsyW3OvMRa/FbfxZR09CBMIiLZKgnBp
56y7C/OrxmLwoc4EAfMX2Yt0baOjeBE43w/nvrO+OyIs/VkmnfVEQ6jNvCGw8zLEAHd+4mGFh7mC
2t0GjHhp70H9ZJ23Lwkwk1LsfMo+hUqSk3VP9TNW6E8TZ1E1g3GYa98hMImkzEeWKCDQTw764Og+
BAw+E+WSWJK1ej1BjJOA6hrgK68CG9VuP/ElH3lFowd/1OYsGPaqimrOQN/Z9TSE1l2P15i3aaDv
ty7DtmQr3QXK+DXusc5cEtYyPd2vtRyhy/gSCBON2TBdr1xNonq/rs7LeoLnLImwnXhUCgvU+Mmg
OG03XwPmcq5Ujbc3uaaU4XGCz67h6YT3oWi0W05CSDua3hAmhpfJtCdep1eSkTVFptT3Y9PGbD4U
ho/f327oijq3ZpkVW2c+zFTSAohsGIq1feu4zlh9PidfvmnhJXPZS34QlgG7OH3d5jd38ZJZq3Vg
AxuI6wnufea+dBIKWpVLFF0jhqleexwwXxGC2Mfi2ABR16M6EUArSC1U99D9S74H8oOshFBSx4BG
W9Qwijz1I2Isxz68U7JQZcG4O05dORUct6HJrpQVXJgzM/zCXm6yxjaJyUFbafiZJbb/iwXU6l82
DFBuJ+i259a8Ug3XelqtG1vYtSOX9+N3/NJpiH918nhec76CqpRv/T5eL5VP70fRZ5Pvv4O5hu5T
wRAvrPyu35sU1BJkEtJchBHxx9ldxOuThtDEGhbzL5EWKfWrGaWU1fxZ1flnjOs/YSsPlFikP7rr
KxOeRD8BKi6f75mGax0mbmMIW7c328NEaCbDrxRSDaeKI0W33vlG/ZG2iC/3oGOIAP6kV7uhLMud
4YBGHzSNLZno5Hsi9iYBRAcd1Hl45UYjMUB8GCK897RKjKQnwxmfJvoQIM7OIRla7/XrGvL5cCC9
QXPoYMyhwcaQUOPwHpPqXhT4+Y0bZeK7HGwD8uccrlfmWiMk0fpyDEA2vnaLnXMObkvYe+d3AdWZ
Ie+PKCj7qkrLiUPUBGTVMyLfvKQeIgB2uFl08HcEW05/9ioyrIvp6cAgyCSB5feDjJLuDTc4jww+
tTjggYJo909WSETupc1/o7XBjpW3D0ryRyESHfT47ZmZeYDinoRylpejuVN7VTSACe08bycdTPqz
X32xbwVbLbVedkQ9yDOr0qGTZ2RNIgYNb5qBFzUREiI2AOAjLlol2CRjVtRXYxFepgyjijkRFrfj
WgteWeHbR50v5loK7+CRMPXeFS7exXH0pewSFOHnrRVDn9MVdjNLHdRZbIa1uYAZqB4zoxXtB6fy
Cdbsfits7X6vvMxtOYKpH4MtxDrt/+ZTVXYsVBvuDTB6lmD8L3lTYnKKeJAZDLH1DB6ujqHpiydR
Lxlx8t3tpiVO0FueXXAs7HIZVUWNYde1fzMlbLqGFb29KCFVzWAj+J3cRugbRK9tDh40s7nLAWUC
oK83NHCePM+rrurLWtjRW55Wf+GrvpUKqyoVSlSIWOg+gy1C4U1MCt/I8EKL8AYxf7FbQuu4wzXv
NYdIE39Spu6ngBcqRkENL/s31wOh7RHYlYQ5GgVt5/aZRlF3kpPW88ewYvW5CYWeMcXCYYpL++j2
82A6U/PzKXw6XTHmtOrjrInR/inE1Z2PwOMvbYJ2cagqdIIFDwLIsdi1AIZ5XNzJs/VHZyNT7DvO
5rvzJHbppHEhsi2Fy+bainOC8WtERcYaHVc3/Y+bUZjQqPwH3Mbh6SVQgoGFmn/F9rt+t9ckvOFl
UHbNNfn33h0J4EL53kuFyAdiP2dYFpfVm6auS+W0VBtjukjjKTMaMPTcGMn6SVLYA4PokoW6umlN
iQj9DTt0gNxCjJyMsFODsdmlP6cukTENS8KcDqTC7fpA70OQzKclqGARKE0NpcI/Hv3PKw9FBzKL
r1INoPTVKjKhgxvHQ/D0BxWxOJTtYH8BPIbZz11wrfP60X7UROpl/A7xpy5mrkvDTDJCI2KsYNDG
2Vjdxo2J+/WEWaeW01XP25Xen6I+ZSaRwQhAYg+Fngc/Kgimc2Xd21ZNYxRHI2j0QtULlXLkZdDN
YqPaqYlEV8noATwajZr2iJb9NiHLHO52IVMR64BmFNX2B5rLU1CfWvmZEBOvflxpXky3KMzQExBN
B/xGAESt/Qikg+0cH0jBtKTLo4IkBsnpC7EhFaX/xOSMufyYLXKywM6x93xj8fEg/QftlrBoIP8O
D4JeJeXc3wP8SHmR+edAOQrZS+LeuZNqkECsgz4c4+08QSKI6h4VgukhErTzl0X5rWEI3Jh1vk90
CzvegJnvKWTJdzLnkJTaM7MvNq7vcUKNcgLBTxNjxvWDmpGv24RbfIvtBOFPUAW5jLcndV9nNtiA
nYGboBaDpLemmm1+2pnXnyV6iJgu7xDqhlvllgvLdouWb3O8Mp0zhQUg/OdDtoK8lK+HmXqiD2Y0
aApMd6fmpA0kF+cKZpB4nHryZplQnCigMm8PAptsxKqCW/4URgmAiygL4QeSkz55oTcvYWgFq23l
6xiXmw01caLdYKVS2VaPNoamXAC3sNKp0t6z7HWtBKYuHfOpGLmZF/vblYRDNhPVhY1dRNS+ukLX
HksnUsoFcJPm9YxSPHWNUBT9lwcuI4+YsI7QP2IJZxJugsB67QIMN9Ky/B++kjbW656YGaH4L2Ov
uqv9pnplxO3ThLbeTcFCM0FBGPKAJFha3ijxN+YM5X/jy92DZnX8uJaBdEHxrXkvnUAz3E7jhOXX
gIQN6sYKPYNG0Ki/i0qLiCSROa5MoWDIeRRJmGrtjwY1lgb64A9a5bCjeINi0MQh2HpMBCvHmRVJ
aWNeWfd7uH+40weuufLyjf/0NJBSBS8yzsdqlCCGTGyP9PQrRsXju2VOi3Im6Syh1OkEDwckqpRi
QIRHnYuChGq/W991ZNGSu8RhS1InkbhT4fFY4MXCp6MYfbkEgtouufcQG0Iv76W0MNGTZiRB3nEO
226bez5qzoslbPa8YYQN3WlgSjOxqqK7l0P42UkyW3A7DwYSbrysnpD7g414W2UO9UfbqYtz7cye
J/Lq/SU0RmNJx4YUrLnETNjnjrF0tKnu50TLqyw6ZflKVY4Uo0VeuP/CeRYyUWp+KrzqbHcBREvV
zZDCcd0H0/nDFENicJOQG+C071uALbA0c68id7W9CwC6K4xKTbY9tmjDzhn5lvjZbziKyiQ260KO
FGg8iiIOS8z3VLLbGonYTkZV62rZu+UfM58GgaNuv3pfurCX5fdweCpG0QwQJk57g/rUpJD660nD
N3WKydWKsxOQLYx1mghExK+FdYs8C1gwAK5QMWzVPQKRNV6QHbL/M43xeej5qO6A+xkw9GDLKgTv
1twJQgtO/8rEgHatSN04zfLP/bQRZbZhX0ficoJ4E+JYSNUIS52kihFCkbpQ8dGyQYmm0LRTNzDr
0HW1IycWBYu6bWS/febCoYaKiF3cZhkJXSv6Cj3MGjqNWzjLz7ghGGEhyousdEnUJGA9u8q1mGKS
AmyAxUGxV3LU4yLxMZRdytZ7u6MZntKJjkISPeeE7TpUiJuOY6tJB1Yhb/ELY72KFgfbSwosXkKr
H5C3XwQEdTtkvx55o7cISc97VHN8/EECC0KQDBkjhCAoMNEV6sMOtXBgeJGLKRCl6MfAFcgErhDA
Nvu5gZACxjf6+tLor97AjacvGww0MMgNbjr7qfaPYgDZ2t7UKJtZdEsiMQ1MVZJWEIjk8ZUivz56
xMhLxx9XhrFOWfQhzMvr0NZ2S/AYHikzA5zWz1uQdc6fuv5VX2pbJOZdz/Odkpd1oAJEdO8U2w4d
KP3+dfkmtPeX3SJnDvq1A0c4oC+xfHtPPREUxEQGmi0VcrYUAM02obDjY3P5CCnLtYZxB1C7Cy0z
QJ8WlcuYTlzzVMldL3Tl97Nv+64xtozMAWIzIFZHEeIihOwfPLaDvF2SlMrTIGoHyx6sx+ZA6xI6
JW4ZQWOjFIMyNOQS7NOUnGxR82/02cbW4ssU9Orrj3z3CWQGYs+zYuzdBYIz2lv7nFuPbLOwI2m/
QJeSo10wL69YY/QmfWO1QXVO6jX8FBUa0IEQw5titePmOnvG1/fdt6LapY+EJc7qSQxRLb+WwbMB
0et3ryGaOyIy0kDriBP9e7kXBI1r+/Ko+Zw54+//VE6/34QufJgPbLy/3qLQzmLIQfjRy7pMl29x
rYyOR2yYSroK4uzxGgnGxfZPZ9CfXt2g1R+rcCQd8/LIkZ2p0Fuu/P4zRz3eQMZ5B31ldMoydOeG
0kgku6temErfxx3kEglVQgpP3sAKAWG1mk859Gntl2O5dFw5OZtf3ucPY14yZaK0nLgaKEKfB90+
WXWOUBzn7KtxPhCklnEgfuWGO8bkiJE+IdEkJYAGrhQeXNYM9JQos+KU+K8qejP6L3PkbKLIS1PB
X9WERd7JMkpds2PdQdaUWUoweDdZxvJICrDeJwL9XOO1ECBhE/Ot/Ku8M+K4akjKsNK2lL3dwd9O
spS//dvBLyhdGa82PZhPmOtgg23d+fFxJu0PFCY7REmnTiE7doqkKmnv/tOp9JZqHKPD1NqA5Xev
zsf9fps3za4eyLqmJii5TMl2cchqtkyrs6dYVmNudmFYYqG/8255r50F+GWzI2edlmAjACx4LV2g
jpB7Q7EnHYJ6qDkkUH1XCjgoBcrlYnD1WMNjYq2DhU3ba/5n744GS66vAeGS/2h2bLSRAax9sE+Z
t11+Usv/H+YGY3Ikp2wSgnMQGWJpncD5dCCqyDVGIULINeD/MMVsmk3z7Uxe6BK2FEX9LN4IjfHy
zydzp3kNtYSh/WhUzLKbSgQSgzzVfUewIzzMY5bbFzWkk6BXcxYw6V4zEm2sIsTo8GB5LGNb88RY
1f4Pj8fa/Rne4fAVwwsOGIOoY8DCHO2tRNWFJd7yDb725n97IaKurUjrBAH7+p7aZ4e+iBnzxZ/8
J4RdWdHlcB2+p+g3nxHb5NBbOgPPhNZqd/YdxchTpmnYWdxUZdKG1mxyWYk5xDLqPsyZx4W955Oh
OeihLlDpQVtJisJBV3KX3GdhnT6dHDOrfE3a8ccH3teF//+kgNEzFFmIUj7cKUKi1Q1kwLtqGFRq
xlqCgl/KamH8AoHhzETCwi0hCA9Fmg6bTMq++h5lYTRbE/UtLbeqt8mM+vp6zZ0r8pHyxSZQpO23
MU+Ic1FCgcjswP60sDJSIWOZI2dR397Nh4DfXDSd49x+SHpMfA8Astr1//KDCi2FHz8vhjGD3yrz
KQMVc7iCv6y8SjWHdK+eW3OLaj7Wln4qoX+yq/P3skxOwTk7LYVBY+lpRInwo1lrqdVi4tgAsazG
68qJaxvbJAP1xZJqsNV2JDXHK94xt0TysJvuQ/aZbjQCXQDXynl3j9sg6gB8zcUVRczC0ewPQ4WA
UdQ0WTntIjTTCLkS4GDH1s/JsP40Ejf1fyxhHo89esOjZOCB3GJSpZHxh7hU3jrYhxbJKc2KiyB9
P5kK8ssKzW5WtEU8pwCDNdW/9Bi6rWBWoR8E++jjOMb/28cClCDvvTX4rQ7JcUVBniRmahhdgRkM
13MpfkK51FnGRggSoqVvGsMHGoV3VlSi1NNZ+/MKKTBN1nRi2aeZlkPy8+M+A35DST0L7rmHFHxp
i1xjTWFdE179xrTQS9zXsEb7I6XTJHYbJs9To00h4m6nkvnWyTugfuMStXtVcwvgDX0gWRz1gdR+
CMwhD1D6ewC/fmkQc9wdwrwnD+Tfwo9ub+JEkXHSrjOc5EhEO2hc+X6jLVZtRs4Z9NouS/3Zs5vN
2kwMumZljW65nO9lUXaXy0TLAVMqUfduqSqG1rsHVd3PaYrmZup4iH9p91BHaUSSUJXpGXTkOXJG
nzDGBeA5YcnRzecwEBOc+FSgVwdtsFSnMGFZOxp47+Gs5cNiAYOgUSgyTmZQBZ82NICKPf3VdpBS
qnscRSjz26I5UD7gfuuqsPxgU1HX/hx6v+o5RBKvmAVPvu0oWiR2ADUB75JMlLR2YKKS7nX3j12t
QZG7hY5BAht7r6kwScE+LIEW+pxEkj493mrs841ad0s5DD4+r7VAJWDiGTkaS11RF0m3+fUBKy2E
EHWnIWJp+0FfzOUXnRKbk0PAMYg8C8AF0UWI91p++tMBmch83hxgia1Eo6E2wcecur/XNWYAqdDj
XHC1YonvERP/rUxmJdctg2Zc1DAx1MZzPaJwEX8avhfRbmwm2kNt5kKnTgN5aqM9zXMHl1MpF45L
klPfwZ3POzOQUsDvamRUnjHBE4ionCwVOzPRq2qAglDkzm8x1HiYNbPVqa27mJyCusZohoMsMhBO
QWwliNp3xcNNnEDZw43fw2oP5TJomOn22+5ojPVEs39w0RTeHuPgSgFfphoIT8mcBMZ45S95hktb
YxlTsDDm3i3coVY/aMz67j0xiSuFKSx2istTUhJl+2r/JboGvKNVJujSO1eaQL/Dubd88j2JT0gv
8xNCT2tr5JzJFvyRDTpXBfBF0ytYzwPAFjTWtLFXJU2Xv4HXJyfK7/92EghmkuXd0sJdgqP18kwT
RKrfZaDcnv7Z/k43CocU0FvZVPRIBIiRjuJFIMVS+EZqjfnVeryDzQDzknL4xe7FuMA4OJ3hwXuV
ehPX4FzAmvYeN3JfGoPrRAU5BkFWSEJgYxPxSrbcbsGDxGPSqgQhtTkKNV0XuT7jyUN/ym1GBx1a
GjSYKaGMvFa+qW2omnmtnGUykGajrHrhHFrWdZZRudkIa6P7tidG9gf3z+E34y5JCXrTAXvh0Neq
6Yauy+DCMYOVXnL07M2xh0vkyMg9EBpoBYUBMZIzN/qq1IRpmjB4Pw6omD9yrDLH5qvGcvmmZND8
MeX6DmobcauY9IMkIE4oxj70PG7ROB68obumaQJp8eV+KTaO8e0cQSOadxEnbxKhUkPmNp2z7scn
MnOGPUCByXSg04xGhBzFP9G6YGsHf3mEdzZA7Dt2BJUU20r8hhL64I7//Cwws7bO9ZltmW9Rkeyl
L3XJLYQbEPgO12CwK61tHwGLvIWGOHyQm+UeAiUQJLAmxOI8+e7OajhnQrMWKQy4QfskkSCR8I1s
vftxigSHUWo4RHisMiZlejhWP0FnsgN+8RjqZcmyJpz/jwDqrN060N1w2BkC9UNsvBxL8x/M7zXm
UtcuVKZSuUnbH1BbR/daTI/B02HRku8KN19jlW/wokf1X2mmp0k/eEoMeQ0iKuOMzDcCnSvJNJTN
G8hLkMIlBWJB84fJB3rhOrdJ82erXDVa5LJqzH85CQw4Sf9/iGIxq1oQ2SqjJNYhMtTgQWsZUYtP
ck1o+5FCheuq932eASiBKuy0znknBnhvDiMsv6oDpqq7A9epfgQsTUi0nKi7SPIF8NYl+XM+jqr1
+gWokF/GVS1MJM81bEsmVN78Rkx1IA+83Aatdim7sxUkLeyJrduzXVJS2qyeZ5DzvpwfM6tIdTyy
PRWMayhpkZdmzcF7aPL1JSSyogdekrtO0ibpf4Zb0pTbESZqVtyoD0m4Z++WrNJep2s++JsQBCF5
BiNkgEx83AMqlMpyELSA8jekMzr5l9m9nm1YULu8bkLyTJDt4pVduW28LmvZ2wm8jbXxWLdQQIIJ
lOpAYlVVVC1oLDiH+O0HVbCU32DZ4xAxFjaTQH34BxD5wjMLi0HlleL4tlNaYNG+iQaQkCfj7X0a
xN9299FR/2XZwYMQcGSSY5vmiK0D5TH9L5WcZTpT99q4J87/GYd/nFAtd0hoslaot4gyVqhrkVIz
pi+GYIWe1JoMt8jTpt8bpSHTXqBo+7+4iwciXkS1JJrLA3SL4+FdrsMAQaGQ/OpdcpOzAa2RGoXn
aflAdxbgc6RQv4+mI+xe1ZuthdRYXJvHl/ZJ0y9nbcdh/EvxFiWki6c8c/YfF5H9wR/MxxxWPEsQ
MFzQYaTlDxDLwgxxNtvJNmKpD/YW5Rm+ZPlsrLh/Qzsii72ehK4IfYsQCnbmtyCqKgknJdIiMnJ8
/bCiOKGY+2+edzisTeWVRrksUIUz444l7EE8koOuwuCq1MZP5j64vO903mMueK/mgbX8qaOJa8ED
b0FTlxnyar7uevLViiwcOznNVsG9HXH31YKKk/IXGdn4u+LYtffR/Xe+04ZiZMPjVZN7eNS4ygC+
M/EfyQwUdXCp/rBm8d716ELrfPB5XiqlYL1PA5UNMMFJCTGk1nqudd/R/gzRstHr6JQrQ9PxCiFJ
VkL/T2J8/8ahsKNOKfRhvk/vkG6nqd40HNziOLn3VPRuyolMcZI6FsqnF5a4PbRZ7iaGApliQLZ2
npkhCuKupMaVK7/ril7pydtn38CYWtA8AI0nCO1Yg6s5SMY+HWtscH1uWCU5VSz8AiIc0979kLiQ
5qXItNAoo/jT+hk70iQ/5PwuTylWyHxUpmzFXIZTEg8gxYpxZNR+ovhWIC/5jCfAf9ZSUKq+8grw
ob8mtgHWV4xcz1wWiHADAsq6DDuExxvgopyHy5p0+pgNAtJgmuLRbgInk/zbfhItNRfkE/FdI1EM
AIMnehzkZrgPeXTuGXQ2HnjZtq66wyl2G4/7sPPyMvvCrXsikEidfsx7jnwhLcP/w/lLphc20ppY
tPZj1a3w4nwBVSq2k+bQDKmWKxmvjnxaoeN1zzs33Q6xQXnoUS9rOzNSvORTgCDOmWi289uSmYAE
3P/Qks+j2gE+nCcHi80RxtprMENLY/JP2K+3kWs+u7xBMdfP/tqmGasVYCb7kQtqG0o1C97aFvua
R3dsKb+QNQ42KeSf/YnyuQG57FaFdgdatdTH51k0t4qjhnBMrWB5M6dL/7yuGmWZcL5siLXY/E4Q
8iJ/XSlAEVqqJyuUzMK6HY+u6Zg9A56+85rD64XfVUNTNb7RT3opYN81qkC9fQd2/zVIFeiRLe/2
LySPsPDAX1T0z1XJPM8pHtjc5PrbhD2hd1uSLfAk1LiBNnvWZysXDd87Ehg42QbR8/oWe0+cww6j
nnlEapbj4Rjon5YFLvTJ4rDnGaqB376I/liihZVKuMTIuuJJF+B07bcFD0DZOSnFcwgTGE1zXf7B
FrgCYMvVi3+pz1C4XgyRFrR+UpiZuEftNcz3Ys+9L/vOvKU1vUiGNVByt5pahhHF1TPio7uOzOlE
aqrmVYF39qtOKO+1R9FhiN3qn5J1hyzevaKJGRZor3ldguJITqje91tmX5OKdSutDve2avBAIrLc
2tKHDQyNOTtnAUGN/gJ1lYNe1x7WJW/O4X5LBzQAmZE/LhlfjFQWcJqhwhcPwPTHvoS0PHFmnvRx
dynumGwJi0ZeE41iSTHk1DcVy7wETZSEfwVwzTIBGmAokcp0Q/dKEvBYA+HjYQa51YPDHcp9IUVZ
ycEZd7DqQ7Z4LCMVZuzmweC+h/xpVKyPLSauGQ8SSRpZnvkfs79CKR1ahxypFGUH6YFIiB7gkoMX
BPaneuQm19n3qk9+/LMc83vpFngV9HYsUApDjgFtkR+tBHXy1KxshjqyLw68JChpMwvtxDLVGFB5
yGs6QV6zdMxX92zkv8Kw7jzngayt5m6JGNLmGxvTthOBihzYsiIkjyWLmfgB4itLoakPGD4Wapz3
pItky8LrQc4CXRdSGBS36xkbApGtVB2d/tW5mpR5HYUR2RNoMrjqeliU4zoWYQ5OCxhENYLPn0/d
4nPdJV5JPRmmUGTjv/W8JZMi/aZA8FDrPel8dUoBOSTTn1jvlUh3BMjJ2GPPMOHsREIbPvcjZO38
/UwIcfBKLC7fFixVrXZUA5OqdjY6J2zxaULz5DF7vd45ULIIHb3Dbyc66Ewm3X9Ao7K8//PFB4Dk
S6g1Q895ZPKE1eYu5zFuTlkxdCxbaBjyvS1pn0A2TKi1dH3ABxADeKAzNKRjt7bN5WKYtuHaCgZ3
WB7SFTwBj7eUlvtBD4XWnN0PLA1j5qsYS30vtUG+VaAOeGgVhS6ruXWhvu3Z1xurXfbaM5bccMah
Fcg4Mf3GH19njG57nnUh5PJF+hT+YdjeaQFRY/VYkDV2C/sN6IvM9E7RTkbK80U7CKbWaF+hUvfV
kHNnhBdAaEEfs6ty2pDZj2dTKSF97RzJCCEbWJuX9QnTP4lvZOd5q7qHUjUeQVAvA/Zr3EXtGvU5
arA8rG4ucmGk4rxq55n8wMQsOamqo5wbR8pRmRKgs8qAoArHP8GbuMK9OYZ99x+wfSZNDF8cHmJX
pFvOVBKb6CpSXazyI97xZB3WsqtduCL8C0MzLXUDZIRLXLVtXN4Y4p6VMqTXBGRnorODBE6HRobf
giJ3bwT36UE10rZY4D3tdvGmCHBKctI69Bw7cTuZfVC7mns3r26PjDRsw4bBiNK216mFgTlmqWJy
oslCnUpqHfsenT+OgTE+Hrqi+zQR6jp7p5Yhis4VuQU0NXr/lucmP/hs0jhULqmOJblzFmM10MNk
FHuHsjf29GwgKWgayK/JA/0MLL7BQV3G+w9TawWmuVvQV3rvruzm2idCBb4A3jEPrQoAzoMycvgA
zCd2AFvqFM5f0h2fVgP/HKX098pfXibXIXzpFXfWQ7ESAVjcIiwDnJD7i+Yz2uMFsNgtFyQL2rAb
gSe+o8oz+U1BqFRcGpt/hWkRStTSoRZHLmEv5UILR47B6Gm2CR98N+9gk7yTTp4IJ52lp2nQ01PQ
sobwUI4gxkQcDRfkDHByXbRhTTkWrCJcpa1G4bP3mutlrudIkN1BlUq49UU/SRsd9gzUURRgbNwu
UXrt+TsVZcNhtHOZEuE1+deLwU3maU8KLJskBp0R5WCLuxMrtH/EtQQViodOgxNWnuCxIpOl6nZv
mydpVDBfkqJDt9fEA1aArkHOvslKlx4jgrRXzmzB42VExLuylheeXMXnNiF+bGP2UTnok4ZVh37X
N1hQT+pq+0Y3WtZIzgk7ckzBaTvZ9DHbVppixGqgAMsmAIVwKCWOccF1BiQvPPS0liMqMOL9Wpjc
0ygI6Q/NxuVbfSi/bYD+kt6t3WHglFgR4Cf3xc3k+14ZumfWK3sMnvhVYquCsjvp/qTTepSCgHDf
kaicARzfY0/BySQjyCR/xcsxgUeLrfLm/zVBn6rY7WegjAtLBKIwzANyb09QYy54gKH+QDIWl3fv
DItZUdPKRsfmFNqdjKHc+zomqLqTGUbS0ItzR/ginZsOD5fgKspR0giFblA0LoW5zQZFMq8s4SwF
GxVhHvxRZJdS/X0O+phngUq4mGDHQc8g3I6lWzGYO+1lZgAKHbrldwBFBHWXUf3JhtAMfVC5+bvf
PxlkcpnrcGQ43hLg0qFfndxlEOPJiwBKth76zWtt0w8ZS0Tlg5dF1kowSzYjgN3od6gjisb1Mbfo
rFRp7EkC/2s125mCxAHFO++2S3mVTgLJoxHDgX5mlVULP8Fvf/3oCjXWcKAkxJ0JK7XArG+kIReN
87nsYOyVcq376A5XiZsXMgMCo6eCVteyQ1GEP/E04DyC5c5XgnabPCtaUpiMKyZbucd1yGtzNM29
mltca/KwEwnqxgTnfnn+SO/WjuKLKe3SabqS46936RqG47SELieb6Bp222ZuZ9DnZZFetrHAmBN6
POmBxMHD+ceKm8PeLsKunUN4UF3wL05r4T0z1ZqVmNCtKGeErWAB7s1dgqSKgitTC7IJpgXRceWA
/F8TvX07nCjXP82LmwMMGg2UkRhRjLdzBg7lvNMyoPyUzxGF2dahbK8UPyGNScElOYwCkm58SeMQ
O2R198fKpYZn04dKKVLSu0T+ns0m4Xt8JzQNNE6XaBvVoBNirrI1i1dCw/QxnGFvTmaSuUwBZ7TS
+uy7gvXicYNkpply8Po1vh226gdndbeobYs1YR74stqX0bQJZIeu7+1b3s4q7JxdleMNzQ3zrOrn
mcmWPHLf5JgACOVEvFZSFI8HkaSEHrHcI+FNlqhXTAXXCwjdLdN0j4Xym90zi8joS193Kqwt8c9G
OPOo+os0g4QOV20TQKSgXq0BK6nGK7sq0CSrcXBK2Io7n7hwr3+bM3701nuvrTDRv8OWRrOsVK1h
IuFXOwYJEk5qnZ2hIvpEgfi10X7eUSGlVq+3ZHseqoKWCM1C8acbrXt5PRUTUS/kM4PVM4Dk3deg
EhzIWh/qCyysgbb2e6HT0rLKotRD531exNUIb6WsLfg0AWHpHtSksHVJSRTqe9tHsnqOG7JDMA8O
PbPguI2sBjxpTCIqj/Xej2DDMefjeGGQm5OK3oVaqGhvLUpl6+z+Gm/j6K8UnhrWw9A0Vzci0Aed
GD7xH6b9MsbWQxhBgLhWN60/FFfXhqHn6EvZjQYvMnd0eWofj3iODQaRne3Y8g+55VUWif182bkP
+hdO5Ze8qYuLmhNg+mc6ZFZJxI7PCsnil+YkjvrweII4pWHuPafJbbZB9u2lcwkAKe/zwQqfjxSC
6J8ZOnBd+0DPJ3aRUyleQukfCPuyHtHa4pRObXEN18fjMB0SNegxuKrOTw4kpU7z4rfe8GlePpVp
0b9+F1kT//r2vaWlv5YFwSrYpNI/QyOCy5bVwe4pLmwi4C+Xx52T67AYWR4NN6w/4b8wdubKXnN8
8brR4LW0tRUNLAmfRUPMH5KRXqF9FQrhNBHeQ4ioStb1ZixEyHtRSJGrvAOzlC7uLzwKClzn/IL1
w8bk9QGdE97yiWP4we+yHtm0tKXvWd05RlbTXJyRsL3vn+UVbraNG//Xajy7NfYHCfsNOkMW68NZ
5KpcxZoip3uPpXW8qxQo2KjqQFEm41VstpP8yz59UcMXTfeVLYafSUHA1vmE0b6H1gUe8N3biOm1
+u2DVpseRqfgmVGPq2IGZyYgKdcQsuNW+Wutov2466i1hH74SoIGMXVs+mr6Ta13up1Ce99iJLpc
x6+v2OynYiA8hHvdNsr9W/83nMa7UeU97PWmufdvCxlK0Z8YCBVJzvpYqM22IbAHpKcfCHFe4BpA
pHqsMbnyZJ3RcVVh2NIrnL+F9OFPhrijOkOopogpyp4U/oPyA/SDe7JNoq9A0JCOXHRitq6VJZ7T
ff/m7CsWuuYmEJ92XX0MxzXIpDQxHrbq9P6Z39IziX1NrW57SzM3MGOy3FgASKMiZmnIxeik+jlJ
5CvxOFTsMmgpDGdPTfvyMImGgXedYliv821htBQts/kOtGRgGnPDgPxacMNMAERSc7H5JFcrEprk
6mk/jz14fp3dzSDWvupVSTW+12FAkJHWdkohjVZ5UvHPi95yAfWF252Mh7ypc3c5qVUULPVXtEeV
0zid5t5KPutrEdE8eRW5pYPWYJKCYo0evecX+bUARCE7o8NokQFyTSmhq0pbgITaywU/WQeSzbqt
z1gJS/b/4d4k9zWbGMKJDY+4VYs2IAsy1xuKmp/xo+zqY7H/+xxhnXDSe8wn2TtZDwl/hOSjNmh+
oz6CEdXihL+gOp2mW1nzp54ZVx52/MsIAqO1JgwHeiNrgvzTi4C5hVK0KiaP8vO3hCUV3Sz+C1R1
KBMqxCJVjklRwLcZ4Z3bkk5MxT3FB3rNXiysYWCfQKwtyb3izvtp+k45ZSmpfu4oYkceH0vTY4QD
k5eKkEgi57QYb4VBgk+qFV7d7xS0wPn7iQD3onKXvuTEwa9B/WQFytryLzg5zIwe3Rs+wY4NtbUC
A1gAX357921kwy56GL4Acg19Is8eTyGQ3CPXRQuhF+oaGqlu58Ntq56ShSeU5Njkg+gfdTCpqUEw
EhUWdE/2+nG/Q4d3MIGsPhxPEc/BSPynmGPjZQTojMIIoBrw0Si2vtZSGdMKSeAY71se3UwxaYMl
EUTJWsRgKe/41pNgTdxm6sweYDYiVYUtWxi4OZS2wpSB/kGifEwdjgMknQsmL7XRsi0RjWHsXmc5
RFsW9SxIt63XUXHM+TPOEpkc7ltopUcCYmJmc1MYg0f0k4xXc23TqK1Vq/DqozaamVKjhP32vA3X
fEEDbV/zstGi76n+McenhPxFicjrMnwP1/qLiPZirTWrkr6oRn+xS50n7++gjZPw2d5YBa1emZ72
fqGeLZO/Qm/SPhgy1dkpyiZc2wm4IqfND5ISPKiPNJJIjvajdI9UkXZaKL3L8bzHELCQs748xQP3
D5JWDBG54QSogmF6jVuk2LEh23MVGxl8IPdwGj3Aq8QFoe3eU2MqHl9x4Fe4NXYOL858K9WUXdc9
8nTpuHhg8JUVuRolKlvXuDfeY6N76FPFCxgSCPYhFPZM3y2XgunzlKZ/ANN1twc7InelWnWQmqdv
H+SFIUVlswUxJZ+7i6TT7EJ+aP4N1YI9ZCpcnTaqBZ6XMIcp6fGEY2T/aH8KU591RghlrHJnuKg+
I5prWzVpLwJYtkpqp1w3JQTAIgrNE4VWz1ws3SJhusUVNqRvaLfdV11dDD1clzoRFYm9Q5iVOtuB
pMNdwAtNC9zzWOE/aEiC7SiD8Y4eFh4TysClm3SlTsaPT//pSu7znG8dO7BlpDy12Xx1O0m9C88b
xN4G4GeC1pjBpp6wCtE7/ODNQiQnzszNYzIbZnq+XkGp6x6sAu8AY3ML0hxPsONZKcOvn0elJRuy
sfK5F/mkpVESpfHsizIL9ZEdcOS5fow3JDHi4k5GkweitFeuJZDh2mt0WPFtv8UGoVV5MyLVeiNd
DNKT9obc23+GCUcmLU5r/5EucnHzJ0JE/xKfmG/RHLgh62LXXyINVRqejPk/aY3f6eK70lwCsgFc
PbEOaZMsg3NUdBxoem5uW2+Y7jNqPSV3MDfm8iAzhZqAacnCadlZxBrRJ8D1gI9uxnBaqaXGkVNq
dwK0lS3Z6FbnPKtMswb+OnGbhDryEmTXsHBl3b7WncE/jNBUFhjiTLzD2mEMH1cNp2Jj2y5chtzE
0/JGKd4S9H4STtZTWjUSuxOU71vAST4c/by/B77NJo4QoqNEOCk6SDjF1v8llK0f8obRCVBSgcB5
2qKA3xaR0PoHSdQxff4oii2fSFj2NRzxmb1WYkzqL73ix0GXgZNeA8fch4FuL0WOAejplnQT1KPj
Lh2XYrd8QXaS22niKHU7V8E+wLr6hlYAqUWUCs1ea/hzH3L/gZ/wljo9k0fd/t66F+beEGUNIc2d
vf5Yf13iz6wcNW2j69IwCKXmUtQGcjlwtFXvet1Q46ZK8oheymyxs++JXn+1W3NjT5mV31ihdTtz
l22sj5JWTnt4k0kCXD7bma3WksOEiEn7P8QudCgqNeQDGXfaW1p6hF2mw6fv58Tr2bc5g8gmlw+d
sleEmPlPCiRFZZGIelc3EnxtMEhP+vyi4YqzRi1LjbTgk/xXSrQMVS7fPDUhO46b8yYGUvU3kw0/
PLon41Jp1Z3I0wml8g/ivUFSS52AAWqEZyxlB6QcjoAowVipN4Hbdnwjedl0HHtO2DI5IkjwnPjo
4EFk1x/aqPCmpquuVKC/7VO/pGjHtGey1MDzCp0U3BOwog6CqwPP+AVEzHRer02m9QHzFORul0ae
ETDbNUQIVeW3lO78UZBmJnaSWMb+zbyP8HSMHkwbNOxTYybvUiBjtxh40NGRXKDXc9KPwblN+Fsc
Cb0zD8Kv+WjOPA5uaKG9qkO9dwmS9X/z/zgy+9EVlgihp12IRYqn4nd2NHwFAtEPhDqXC0hKXHVR
tMVnylzS3VEWjm7yxsj4Q2NrlzO3F31l312ZO15Q1kBjxGtYPIccWnU8a5zT22b38NyDc8PNdnYh
qi10Ama4PJ2KyERZpM5e9rWVbQs9/lCu/K3j0o6liuZ+axds2GwHRXoyJq8P/c91SPKhLCUVJ/rK
nURYwVazh/wvqLIh4f7rtu1gni7LGZN/io8v2V6NWDaiF5489dwuIavqFxTNhgJ38tBJSyR9+ngW
ArzZuj2tZmdfB9ocjF7sKHmeVpPhxBA1n3T1QNh40TJQP1/mVn508O65vcRe5e1GgfY8vFkTbwDj
OEsEld4QbQtKGwiGK0ruTjMyHWM9w2OL1IJXvVRMoh7eung82Cs2YNNwP4Tq4MxmzcEaXbRjgrs0
F5u5001fddZsjbm+K2mkR7lPdyD7ScWazyaaJLve0Jnht3gyyb89iyGKOxQ0Q+bwomh9uBOU9XIX
MG7RhFsT3hqPp52nZ1PyMZ+PaPaII/xuqCWHsXZ9qhw8A5ySJgEhyeIqKfqoFZYcIiHokp651pBf
R0xbVECrMN+Dzgo2DQKGDQZLzsofVxR37cgFU3egAn0wSLBb4dS9pjnSF8TcmdOkptiZ2gqfjZtq
EpRdF+fqZ+ZJMhNWF+7Ip4XUeaOFTKtwdLYN91pPxVs4keIr7+szwB4RzFmooyJ568xsnNxZNldz
fySkhcNEb/RP8swa76YWWEYOUhUvbe/34k8x77Lnt1TE36TYfLW/b75EmxT4rYI25BMQ99DuXepw
w4GBeMxVvPjT5Af4q6fKQtqUPRijF2qUMy8YeNUDvEx/yy4lA8xNqkXRbRU34NOLHwkyOY/0Klli
tEoOTzfUH/GwE3VnCo0bO9i7bZhZ8b4u9EN1528gKWByFqOEUeG4CAV+T1tsZwdKS7mf0gcYkerl
Cc+ajIYUTsLL14BW3BQNJHQCrgHeOVXof/pB0be31mjry5LJ5VLWR+BeDo6XCjGgTrZ4LKHo4eBa
+Nl+59HcekS/awPoQJSwDGyBmSTJyIxm9Ls5dueGBV0WiwCGMnGEqTG/nf+nYfn9YFEA0Nj7b7+m
p7RJumCPpTIdp+BnG/Y3lUuaq8FWECy96sz1qpV+qgDfJLeiwrY8WZj6qUDx6BR4JOLSW0CXeUn4
5T59WPsQcNZBXySN2rfW09i2TEmOZ9OogbhDng8ARwegqWA9J7FsmML1mHKvW4hgUEjNghrmkBAo
9E1rIKjIdWqSfkH/Yfv+fwa2Xsjb47UKzUehXDpmX9ywVW9KmTKda1rxRpL8CGnub8Y7wet5CilR
sFFu3h7KC2SJvChc+IJmFv2QFHnx8yDzcbi/u57LW7MMtv/VjXPAMm1U0wTgBo7sc0BDcRLvxl+w
7V+MIgRliuen47qb/S71mPiTT582EN858D8KBRiPukmUjun9ZwYbTl54pCGN1A7OEi7SX9Fxyz+d
BZYfvHaDmqVn0mxEgidH2mHGGQ9s19GMwPqnsK0ESI+rAPq538I6JEpsLF5pspJzbEQIzxDM8Y+r
UFzhCPs3pqpxwNpUoqq040YKWE5rG4F91VaRcl1F7shwtLFezRWSx+QJmXsuOOLjw+Rmex3xrlhG
yFkn8WF1Al3KUPfnoGB6vIAt5qWI6LkZw7u315feFvBcz1QERPyo7Slxp4kMORFRARS1mwiDz7yp
T7sqzDHFIdW1hvxGiq+PO71muWUG7omjdZRBn/iODoJCRoIYCSY0CildAQiMpIC8Zm5Ivx7TL+OB
XkuFH4GOazU7hSt5kG8N7WglumKNx4gIVJi6BhOpKlwv0qG+YMPO1eKp32vhx5b6Hn5r5gboAKN/
SPXC2UfZK3152bGJXRxdBn5ZP8CL+pWDYOsoW/KSBxFUj0JqTmrQav8V4dChGsFXfTWBWdGG9V3a
UVdN77AUgH/KL0yy7+x40E+Mo3Ro+n6RY09LB/AykI8Rp2hrxAmhWmSXLLuJwkLUtxToJUM2RtG4
e4E9Z+SVzmoKzOHjZmhm/u83tt2kLi1shJpHbUsL3z6yBaaj+70bEUm6UtOoNlD8y/vNqQTmPafk
mO6vpFfpUeUMINccHHf8lxIYR61hOVjWiC9BgEcr9YDpK81zwD10suQWJLGjMQVCKYuBQTZLRepi
iBvjz02Asaq5WB6ZzSRjDmc+qkO/9bUQhYiG0KwSTdXr9ux4MdyROuoCeucLlyJDZQVqg0l+GG4U
LLt5DOIH78KDm06/lF/UfaMe6RPlxtSTSfTAQdxDFFai4w7wXNs+5SaurBq+rTY2QT3vGIZQl8pf
xprvFR9vOG1/yPAlqLt09dFT0mYC1wOIC0f5GmJTKIiqsJ/a02B8N4IQ7lW+WhPlUl3TL9VbQyWE
yxKPMAgjrP2NSoxL0psRoHAdgrnti93MGBa+j0//ZLRktiM/FGRwUxs6ruixr1GdeU5f+l6H59fv
eD6aTZOa35B9QK5DI1klJLHEv51CNhLUOEcwWoNCg4SZkIR2rJaDVh85UlM0Jch/FE3OajFHSxH9
lofRo/TKLFlQ4BYZPphON0TiqH3r8ak/z9MQO3MbtBHX7y5qL6LuEa44s/682BZ+lP/9/H1Wlcib
4umY8UTsAEiGjLA7PEINj+kOncMk7rcW76575wfrS2wD44vr0bkHdnOnt/ditrzESaCEa+Me3yh9
sA5yZidDCX71QYrigBmIbUngfgHZLW9+DkG2UIkTExRgRZXeGrujGidXtuhEU4IINGo1NZScGmyg
vsJBtzKsoE1RFi3qurhLzqJx9Ru9A+qORVJKLyF6rvLDGAxqWa9A0ZQu51JLvmhtWUgSQ1DOFPN5
O/DYWROEynD+GjjE1EyEiD/lXDYwMpySh9jnI3jUJAwyyjAmT6YaDgvdEHnpQRpsHPnpXFvF6IR0
fU+D2VvRyzu75IRpVk+Wv1hZFhbLZQYEdDZ/gK5V/l8pC2Samfm84Gb8x57wmsj1oGXdhtozEqBn
rsCIvj2xXzY1FkGeQPwvxV6bpVIoPI0d3W6M1UQ4dm7fMo7LfFsJ5qlYglYNpKlFjdgX35JspXKr
mNWZYpwHkI0IH9+D8J5SJfc/py7qn7nN1i+kDRrX4aKHPpLKUXOx9RUvKHxVwTXIo4cBeJzxf/Fi
ArDzd33VJncLo99GbihgdDduuIgsHzVbr4khVcTZCGgWG+cP/wGWTQRai7oxRMYKPF2nyw5Wbwo2
+9ZUbC6gL02L8tixJLvqIRHOq1zdIyhcrCJg6C7jUD0EZK4TC5No/EunUeiAnwu0pTgtikNBnRYm
sEKa+G6TeNJik7qoEN7a9OuOZjvE6Y+y/vhqfwMRGTTogDUTeksEetGf61Pe7z/exjmF/wJZC7kV
eB5n3Zso5r1aeNRQbe6A1soxlOSVF+nHsA8QJkFO4zh6qPT4VcYVoD/AlWivBbP+lXy/cGc1VJYK
dizRikjne0i9j7Bmu6A7K93DhrwN1eBnvjVcXYb2fUu+bfV90dhd5x8vEAV3riwYEvEmSaK03q7s
Xq17bKkpi/Ms2AV0DcrFGyhG0Nbx5d0GX+Vmc1f1/OUEwnuGLbMLJF8q27n45kA7PuoNYEDtgBjz
MT0r+UkCo6gbw/97yVF6SlOz5khNighgOqWprOpo7qh9396WHahykuba+2WhngpN/GPK7GNF0Q9u
KU+purAJCnpK0qelXQoS8JDbim1q5qCcmntl053eSnPjURWmeqX/daR5K4LGRl90WyakoWx2Trp+
7Jwc5HGxc9XbE7+1jMN9U0ZE9m3zjCg0qpvkMRCjq3LTjvpqbErQdCqGthCjNSj5hMzx3MQYQqrG
3dalU6L5ThVxGlwtOvPwoQoH2G/LMPuzrqyXFfmGH0V/rSJTXJF43G+OsOhW5vxrGk3PgJoVKsdO
/qWMl44mnPr9mBXiQCYbnxJ2DLFeXci/bsM3DhlFxeFVvFcqDiS2usMRnqIdXdmzTWOwSyMOvy5a
Pe8eOId4lpgiUujFRKjP8SHBFsgRacCI95fz24/xADrhdlSfV+3MUcOIHtUIM4kJNxrXkFl74Qbv
hVhTnbAANTslwVrJpd1NnOYxYu4ul/Ane8f2dVNFYC8dxjLfnKjBRt8p2GbLHYrBaOSYA2iWITrX
mG610P+N/LlS1UW234TL/Kbv8eXenyM8o5TvT4humWUPcrU0DGV92KDr086Xrx9IG326AXz1twvF
GQ9MypXG4c7tUx8U9015wrY00oRgtz7qEAiAC3n34HhEliTRYj2Wr5rsSL1ky4eeFDgMyzKpg2jD
r1UknAICTjC6BQ5hASC9bcIGO0m8H6c1NAJVzK7cxPUW7c7xGYIGOykHzME6/FaloxefAdfXenlI
M+sDO+wbxCLjaYNpK0Ii0Xe3x4eryCWvgvvxnTcXousVfq4EkvWtRu0xZf836BRr+ukdKI0R6Zja
xB13ZwBWwgnyj4SPZ5UVP6U7qz+zva2KUhP4q7DZoOakG/ilDgwfQwhNKNTUxRoaRF39/YpUgQ/Q
bxnzple2zqmxZKHm3oFNZyiRbxkQqRRAePvy+TJFBToXVr7rl6AQNLvJSLe3StbHobuBEN5fJWJM
pJvyCrUBXh+r+ylr6OSx2mK32BM7NGFPuZZyCPfsQ1k2L9T1ZZRGExSInT9SAgLsGcQHNVnLlJyI
UMRUYPWnluf+5g3cmxg0cv/uv2/GSScee9rtZmI/Q+QBTEPgDgJwzrZFAcq7I4WaYCJLr6aOimSs
Kl5EGdARLevmySRBTs6wM65lR4Y5HCsV9Ebk4z7zGSKD6zwm3z3U5hsEvWE5/74WxwUwdn7UhsHw
r5BPeQ8zUzqh90U+vsXqExSybzmPpGNxAiJX+2mxe3SrkAtMDIST7CHKonlRCWYfjg62zaUDAnxS
0V/NfbrpoomhXClBe6Fr0KMOpKpQuYM39EA97e9HbCKx7loYnCU+p7E/OfXRmkYnKQPMmf1vfilB
XWHzY+K1Q1pHlbPS9pXa9cKtzM6O+qNuIpa8I+71se80L0O+12NBhaPt1PufnOIIViB/ZvNEOQi3
6VMAhhwbvDQp2GOy9aFDqxb9Igc9i/IHzbJDRdaeP7dx8OOd8Co58zYfamQGF4MvupFeLrcScI00
E9oVpMMYjYlFZXEvgdcmDOPomVD/KsrGeNKV1MqgJ0FcVi7fiqqF3tn1FnS3aXSuYPOCagMA2aak
Hzl0uzBXSt9x+OEX9uQ5lf2XmCnQ+vYpiXCryLVKl0et9rNJifj6u0+I69gJ8OJcTA9YBnjewJwX
mo9/2wzY8s6sHEd6T9rRtAPatYtCPMyAm6WVVhTE8l32xZAZYChYEnM1heE38kIdKx9q2kzrP5Bn
THNjCAXWF3plIXm5g2IRY0LGTG17xJ2+3Qt+9pbIJVUQ9wNdRN8A2NSF7YSjN+aro4BAI1LYHfpZ
M+pVw0un6yXezGjA2EKt1x/YtGGS+YQaVJI29h456aeZsxO+g5O/A4SPpQUbcGbVE5pV8iYAWWhE
r4gIxFZvBV/53IFNsK5yjXQGeUgZWUpA6igAZDM8D7Q8G0ih4CaSGHY+Omln/Y6x3nIh9zmgMj4N
ZudGenL55GN+MQ5j9f0hPuTfQHT1RBXaNx3HkKuE47MxFK45+8+OULhlAfQGsEisgjQwY9qIIv/s
Fq0bOryF0Do9oQ/8TctYLiFm9ssbWKrc+zM22E9nZb8s3R4f4jsaxslvM0EX766WVb3zlLOV8HgU
AK7VDMCqfWHZRbVPn/c+GEi/Zf0EKowY98kZOFs303gz3iWNwNtWJQXh+KsGv3gbKgvNvG5DAhln
CvsnMUzi4OGNBIhzcqMIaYvkoRZ/k38KNLp5Sumeq+EvbsyeF4SJts/9Q2OJCBSC2tClH3HLmwA/
cplBQCkyOj3rvUDD4WbA2C6Calf3YtfBqwp0GAzZyT1AiJzztSEhUTu3hYUIhhp3sIjxMfERaZfG
uqMnUmPQxO0XuVsYbjyRLiTIhMSFtNIXZkA9Fmkujrm9Qgfu5VjD/DTm7dL5NQ9iGpG3gIN2VVI/
rsAx8ojOj4a/mhgykWZ83bF5sPiYvnrnRz7Ya5DXeDH4bb1yB/w8P7pICIPU9TEwkbqRMYO2BOt2
0oVDPQt5zRy6ackbLaBCYy8ypTfQeyeyP7tIj4zgwjR0jq78+TjdBomxeGi9q6h/1kwm69aq5nSl
sjBL/Ahxd7/O4LRQ18VuaxGcvX8hHSm3KEqyelGQM90LfDkLOwRm3D5g0+wJ/6RABX1ipi0aG2jH
CpDR+gg7xa7XwJYBZ7C2gilULmupmeesiuppLFiNZHJxt5HtSK6UqqmA05qYvLlBjl9rUEkC/y5s
D5PlswIgirfFs6ASGoGDvXvzJ3gziocldZLUY0zWE++RVhBvYsAD7hRQZzvREJpVdhcj27noBEar
Qek2WtWILwL1cw/D3zWc3tNFADkENQcZitGLJ6twR4O8dcajKKBBVk6URYjzvhDWqvBzzmT0NOzQ
Ms+e8KCCWIA0IyC52SzAwwMGtCfPqE+ubySQD/XzFxcBXFRmWKr4W5jn1sLMclyTtb6bIeemI4tC
2ExjzoJ2DGjy5Lx3+hiKnsDwiDxUhM3OQUQ3bjbbBQTmzuXi2MLnivNMND21CmdDJuozZ4MSawXK
yrY6BKM439ioxOHlN8hZlRO9mArz7i8+6vbMbi6t69lv10MN6u2ISOWsNzZwhz6z2TlZFnVR+dqD
90XIR/txAI2xCsJ0HHSudE2QH0gqPLBDKPPQOyxnwYKZqmEXASe+ooaX4goFQ/X2E/nUEss6rwD1
Dn+QBDf4cRRntVZC6Cc78OTTl+lPJiONCSka2d+6XXpVcMGS/NSMqbvBFVK99gXinRUXJXpf4w6C
LGtClT5PFFRjPlzWtPrzVhbDu4xQjEaw3k7ZRCj675yWjOH0Y5sKgnHL3dKLDfD2QOizoyAoUVJ0
2IpVE/LsI21n9BQLtwhtKV/ecUzESb75NDPtLfCdlErrIQkSAv1yOafgyBoNrsgbq6CUCGsrls9q
SsoX6S3Vs51cLDj2LFwod9Xt5j9e/FNxgUWXySEQjea8zt4StY6NsgaH89jKEheYyeLWD6hgRaYB
Uje3l6cKd+ZZFGz5BRb/4k3Ttv6xaZji/Nt39AJDaRtGme663CF9LlEBzHs4fLN1EJ/b2MI/dmt5
auiX8sj6AfLgX0eBbqeD8sqQoiM7xQuNNzTK9nnwMpy0pbQ3oav8iKHdjhBdp91HLGrhqCVFUQkq
LUfCEMyPJokRQPxiI5WsTwz7YThPFXHUoPMRvUt1nRVz/I5F2tuAXP71VQDwpNGxF/x0SyqF3up7
DwJ9Tlm1Zi+gT3e1fH24NzGkayuJllf5roMR8gP9BfnCym4bU35T3f/LRNtEczujKzabPatcKdk2
U64RjJO9GI6BRL30uxHf4YXE8xST5eVyYqjcZUX15LVelNaO91WRcbJyAgDTGRdhMDXTlv9ImFwN
R6WUa+Z0WRCx0B1T7L8Xdls6/RA5hy/B4J6c6buUaM8Ljhe5i9tuRJJsvzsiYsaP6sH7wpKE/AFe
thv9e3iGzoY5fpAJx15rEw2p1HwQSW87C95HjGzN/JvCSL49X7pJxTnwLcK2XNn+ims0aEqzxJEj
lJYElsp+xmGgcwoNsppbbqHSN/7RQu599yL/WogwvBmGCj2Fzf0FB+Iy61NMT5aUAvaiFtW3TC2f
7tXSPZFSFB3rSYW2ggAnrOxsRZ1zZTy03vhI5X0strJ0UX/TkKO4duaMLvgn9Yo7XVTrGTziZWll
3hbSin3ixKJH/ccWiL9GiRxuhRQTYWNI8d6Gutm10ufbbnHp2OG1vYUh5IJ7MOeg+elktNp3tUCL
BVYGSoPoGSR6N96OHH9ygZQ1W6fo38GCZRJEJi0y1DOSYpSXCKdORCiKIw7keCN3njjD+VgLrqYt
SyeLd+nk9SmNC6pJ1aPKgCUo+ZkRcRw3nam1ARZr4yViL7o6sj1IaxaEiEobK0DOrCeE4crEzI2o
cgIvo30LwQWumXBeQpsfNCWRty5Fmen4STtZxP9UKLCDe8BxnD9ZL1JlvySB7S1hh09vtzl4ASZA
HKpa7k7TTWM+qGv8/sXVAJ5CWfigRENvL3HsC2KyENKhCfHGAlPCD0XZcv3sm+D6QFRt7Vd4DCBf
MOeASoeGDuF0+VoBHHGeFED1Pc8Yl8N29gRa5WHHInCw+QCLXX0yF8JhsPw6cKiKHfAFyU8Eee2x
dBOMKpNSaNPJZuz03CMjyQYzuUII9j1t+77Jp2ChOkTil5UGnfa9YWml1fXH6aBiVU5wa80vPKTu
Yc7pADRf0QFH3pDIyZBG79KlOdFohsHZAIHcH7iilD6VRDGYX3WMTJgNsb4228Axa5GCd4RofUCE
boBW5HjUoZqR/IbHootqtzuoZ2keRb27wGU8EWTBVIn7HE34pT+fES3y8cIQt7z3uD/rsrA8I4Uu
5JOim8POMTy+tDi0hiHlVEiflSS9FRdmHLemE3e2DBiTZjLC7ljPBUMb8hCAK+CA/XLtwWUkNUHw
QBzV3gQSSoB8lR0COYGTDo0B1J+GCvpTstJwioxH4PKS6b4daSb+ymnYgXZu5c0xozjVymGYJMuY
Kx3+wAwK0t4De/DSu19xTGOY/4PzdhUT2vXxVeIfICrMumIgP8VZY90I1C9ozVXbS3p72O59G2Ok
ZcWrB25vUrpjoXWCNjWoct9lMMCWNG2LidkYJdY7kixnVd1u+/UxaVgekMVxGJpbUHh5o0O6KSl6
v+2GX27Ieb9ieEQAnIe33Dlsp3AJJc7E0YE+8O4QEbO57UT8hWmuRD8XalDgVZKrpLxji+hTsVuQ
EiARktER0pSYAsnVXRDs0xRUpdg5yQY+22YotDZzd5TcA15Q55fmRsEexTe6zvnruGrTOSM1xvfk
OatrDl3xBKa1l1VbVu3kcloohUyLdkfUCpAfNLpM89RZQUNyhXqv8Yu29ou5qghf/0oR+NAnddG9
e+d0aXNn0fE12FQXtVTTpL2XlZh0IiImcVNt+DcpCAG9wCyW8iRZTiZ75xVaT1ecFdLbkvEx9vBf
qvtxKvdOWOXQBTadvZVqQ5lMAcTEaCIsMCPftZ8Vj/Lz+pEI1YeB4hgXmPH7MGWTxi6a+Vym+cXc
yanoxGaRmHXoWJ5JesDufVR3OcYIrxomrTTGSKPBpaJar4lrasleAyHD1SMcZxP25ALrioYi2q8h
hZuZ6yTJlcEIpFHuNG7kVFdHt0kBszns4QyZEkAa+A7HRd/NCIaVvDPcUoPi8lvPCfa7R5Cx3g3b
f7x7qxhJuMgcC4dZLchyCZPACHNaXSftdu6utgjByGYp5Tocv5L6Woy7n5w80zsiKXrNr6XjBqT0
5m6LeuYvu8GorFCOYtM26yGirL2LNaLpfSxqsZIlkCog2nvJKC6jUYk0RwU19ZzP79sCxQwWggbi
V260O8oQ0XMV3dPs3us4xWWBsQ5gq7JOqw/aIbhTLTDrNLj+m8PDTz1N4ZrzWcSH4N9SFpmgaZP+
lC4UAYJdKd75GYk4EGwIP6SnElHHebAD+O1oVUL+P0JzLxtWfhVSO+uLC9b5r6+DxqAH6ZzPFCML
fagvxV4izYa5A6o36XYOGl4dwXKC1plP7cCdHtln4Ji8qv+ceZnLYu5KGGct/oq0QwCUDVSWpciR
/licP6ePPpsJRFgoNCbFwBeIMCYZfjD/drtOoC1fTC+Petdi8nme2d0GiLBzAxk0IUlZAZtVy8++
qJoAVXbOXZhAPvaGVvRUANF5CN238xhAnAwhsanENWzCz8TPFHbmAGV3Ew7CoHVZFncIftDh9GlK
8QQZeZ5uufh4Y+qtVwqDvvite6Vd1R1aVSh5S4RoHamZGKqofZBzq2FfzbuJ9toYAxw2HFLYJI+x
LJ1OlYpqqCN4P44iuRlHD7x5MKSXQTpsmeedjrAIdvZKJTdYCKackqLDLl1yfPHuidIPLS9V6olJ
+MLMqw4pG16QywhuXvjpmaQ5BCqcY5ow1gGcaWi8Nkh+eDgjgWf6GqpLBtcHwYJT8vwh/BT9bt4x
S6sUmUQTFAw4SIluXCTTW92VoaKeq6FKxWQNP/wzy57UBR8utVGCRJhmlJObBjwtR/L7ap9Fgt6K
S50cPAipxJRdE1Nfe/VOolBG8xipj1E3JKG797nQZzk3Ppj8ATE7TitjZBqCy/vQU0/mZ5J9qzKs
lhd/XB3wm7Renp/m2/g6zuhQSR5Ax50voM3dNP8nOcG1vgUU3eHASyEfifqK6suGdG6W66Ulw8Ki
HuWIcivvHDy+NvfF51QNc45szK55YYgNhY7T/uZvPNdQeAqXtW06TPMf3ifXCDIsiXVrSTzORgj2
ZZE8/itbgVf+WQCHxmXn2pWys3dzp30fIkHLKInkhmPBad/lISGLXUsnU23MmQDqzHNto94ah2rc
5F4KuBLRsjvIKUExByt8OprdDD0wNWSIHYwqAsooExdB8JsdkAysnXV9VVNWve53fUuJHnGaBJ8E
nrd/MXGMiSxEy3ldzfysEbdR4ykX78criVadHDdzjnSZ9xGMFDwq6JE8H8UPpW1CgF47zGKPKYIu
BGiU4Te2/J22LrcrcW+BI8ak4csEW0Kj+cTthNQaXXK22y/JrQLvHQ3Vr8Yz9BOwGzQAPaiHciOq
8E8mPMtvsp4li80M+QE068aWLPB2S/sXiFMhk8kkfO8PmnT4wmWNy9hMy+5O2qDyUy26c+x/1dv0
LK5oRQMY/TumLZjAsiApL6pG2n+hq3h3JPMespgq0br49vYfMpkgoOx0nWGdQF44CDibgTEOD6W+
EzYTqdbaUvtScLQ5Afxn0QszVV+IBUu+QCwNDYM/xpG7C0AlbObwKVZfhoqVhKzz6KGo+9dSsPh+
J1l31ba4Dq3jbJpQo2OgUHhdYYH7+SjUP0ZI0y6MouBVyxHSNQxtqwCMGH/iZHNooznFfveVWbII
lnen1ieuMU2oqGl8IQFAkHQB4/Yk8RvqnwK8Zq7wbZ1vavQY0E5HoWrOsiGL9w7SiOdjEGeffRKM
aNwh/e15pctHvpXJaPHnKaB2DAb+VwM7Ple+4zATjv7i8srQ4/DV5OD5+vt+fvAwBmW1iVje0PAD
9kIt6eRL+yDqdHYaDjjT67OYTI4fCaGl0qm1Jnzlq7D2AvDjvRV+rrOOb+unwfti1fCrbOv6VQqS
TzjIJrY8ayXFxCkVh7mX4MuAjJO3rDpPlBswuLYpahZMadDcGOjB5LiGu85lFbZrJiC09Xtk2tBp
C3gdgjBBuZFcWDnNe0D5Rw8nG+HVeYL9xXU660Sm60anFMwx8SHLjEJumuHNMSuBu+8KYLJGrsL8
EDDI0iAnEV3mq49iDjXVYaTYaBi4RPg7SLFcGHX+Xr1hGtQxeCTAWBZ3nRrQTIdTuUlJmC9Q1SH0
WFSKhmbmFwU+PbT8NEtdvaKu3lvC6nIl+VXeR3efsCbKgm7rsc133msoTI7h1zMmWRVJ3V7+ngJd
z7JBBa3IwTCLw7fxFaInlQ01unF3w0vZ+va9pSpYIVyGBnLyFrvS/ZsOi/r6EGizTkPK0wOAq0GO
5pHoebH72WwwJtJyCr5rYva7YWylKVjviFXTOG9F1RGwPu1pLaNJKwVB62NuSJ8+r1gLrjfRioJ6
5akb3txmPc7bQERI0FtgQKj8A0a38VALZ+ejMjmBoS7IyVUZO+k478LL6S618my5SU1jjTCSxMzn
do/x/A8aswcSziUjSIbY/ukAxFEdgtHp1eVla8YQNzIKLV9qAGynSqgVa81epnfgo6r5w4+ptCCI
lasf7kD5GC/5kJZc70fz9dpJX378LIX6FeHNTanuinq3Oob4AwnU2VntksebK569TayunyYPDXOt
BQW+Iuspi4bBAU1tnG5JoDaMZPCI9FVXs4bDsN+KiNNE8Vh1xmaV46OabwvD02G09KooodZqTpXI
N1gxulgaNmXPdO6XwQOL0nRt2/IOhnSb52eG+7tVgh1ew7sf4gnJyVuXSIpfGkozUQynvbCvEqd5
Ej1MBIkqT6bvT8QxcG9RRtLHbn7XTDJQuL9g3RW9XwA3KszEsJvA9XlRWJhqCQdWFNJYju9rsG0+
MIYfq/od8fwEDNGQ6t/oqY+SfIx08S1YeTe3MyuydyQ9r3nJgzsxjX4U2bdyVptzpvAV39kgGqtX
XXMOabHHUSHc5LB2ZwEqrfLHxRuwlT6X7pwIHoH4oQ9Vizysywf7FBKbFuTcJTF/VJRzUyI22mq7
t/EXxjHYw99gZmZqUdwdOM3pED6HnU2HBOYZ2BlzOvwSdHWcjXFZrlRNEN8dlO8phh94Atanv7Ir
0MTWSAWGR/H5aw8YtyKt79UKrf6eSTh1L6kjtwWwr/a1mhNFsj7MWr8WNB4PTDENh0CZSqHOs5RO
nj7qGRzYEsfQXPd6w7FFUHJP3Z6MCT4VKWyeXk2Gw7kERVjk4oiOSQNP8qBMrenKZxLE/HoOOSlW
LHllWCT2DaeYa5yUaXObHJKEuxo2d8ZfEUJuxhWlmgFX8sJMCN8TYGXeOgdnYrVTsOjHdxgXRKCo
J0P0JcOyskibdOo2sCUmojh8HUqvQWrm9WLe8lAckzO9AT7ampNxIFb2i2Kne276cHal+cPSVtkb
jWzpf+A5BNpN0iF+tzvDRmz6u22mSYqjXxLh5G6J00Vy13+l/jCbatdszU/dfij5L2wLkA4Kpj8l
q7jiEs5xDtzDU3efkrHeoibzNdvN+4VSaTbYRd7uUZchHoZ2JcAOhIso8OGFNb4wAyWwuv980sdo
D2UxpvaJUCL9M0k8dmLZMT12wsoq/+RC/WoF5sj2jCPfBRjBn7qhOptLl2Sd5lvFsyhhZ1rsmUFz
s5cR7fY46PnyvrWPX0b4FDNHQZP6+wpmRJIwI/UzBJ7Y4U/1O6d0FbJzkxnNbBac8N/DH3tkCzN2
SN4Fw7jDalUUJK4N8Ac1S3J3bJAYT+R6RmHpC4PM5iRcTs1xL9c/6d0SLSezV9vLNB16b6fhyy8D
SlbeYyCDnRBIN2AcSnQEvGd3Y2oITq8+YRSj9Tse9F9RBC09kG3R28gWLPhMSl+Met97BCeQvA0L
0ZdYbz7Pk+k8LU8u3s3QehU/P7wksLFOQOmWwLFNVSYfs8PPkbiEejfkgccE9WGkz1O+UwZSdL1y
teGiu3br4PCFU9mJEqXs7zsK60FN1lkxAmUeRQJHeh7gD5wPThbXnXcVtg3szk/wAgj44YgLSUDl
LcETXH3Ni6iM+HwsNtvaLJ0tdyVa0GwBSF5997WVtuPa1+iVAl7DbaT/QNEvwRLkgzeC7H+QWTvl
+sDKJlBeI6MjXLImg6yrkyLKVLHMBAQnBEZa0OxXc8qLRyvhx4wNy1bhuNfWKEDRaQ45YbK7H59X
2HpnV9wqEHRSZJjhWXirh6BBZZkJZPDIyCfHpKw/EJ6E2iZZ3T57aq/K7JvlbEwV2NbdGBGJpZwC
Tx7pvNc0iZndmMwUUf5eNURUOBh/HbOw+wLcD9lrdlbI2nOgNJg9/PD7D5PZOYh65gO6PBkbFkHd
v2HGV1omo5VhqDjP2fb4UT33dSaUdvLnAaZ9jEJPYLGO7XqLu0xiKFlvMn/PiFSeIG7fdllsfUxP
EGkY6a64R428/5aiawGPtBvx2S5jQgzF1N58e/khx9qbDc6lPuZCbEDtrkTV8zZxWxnzNI5VlEfz
NNrJ496dyHJedR/e/FbZXsVZ8+bUx/jT2i+fgr2qicr7kNLkYOtr6BV+VivhNj3UrBW6NzpILp8Z
OGuY8W7Yke/hVNZkZCvX2oDeIJAhugJTv4dXe9GrlWDzSwRl9paDdWfZ16QqT2Zn1ijNApT4OwCh
J2kcalVgqa7VZo8OWU5qq81lS0mTRjMccRMLtw7uGM1cvxFB+qS4uecKjFCI9phF+2xp7Bspaiqk
DkOtfX5IFFf342W5Dl1rLnm42OkYCQH9sxVGQLJn+ebsTrGgONxnNcjuecXxduQJmsqV8BfiWRK6
Ry47bTChup2n3XE0B0i4hn8NMZmgdBxs6ekDISc8M57lZZ4FVNZKYywRJ2swp4KlCLgyG/c1vW9c
S6VdE+0vJvttieoWkAQjrHaD9593BLVksudE9bHaDPWEj7vm0j06Zymg1FNbV3hV2ae9VgLY7cQm
4AB2h8ZXlR9kjPjv0dAFd1/7E7wX83cwBxzBFFGkCmOcb+3hwjpABZgodpdZ9dDrmtnQux8soQoG
ikYsSehp7iIxHyh2PTUiyJV1GYC4qgkbEmhYkyqLNsv9fF1LOKHwAkaIK+fRpkiMJjPQ3C8bIOve
hoF133saG32eu35krJ21A/Y59UyqDtABfqwNpNhJGTfnilMPujK3uM9POAjQ+szbso8+gvtlxo1n
GTNao+cfwZJ9IQzzXROxsRenR4hDWukePEQB9dV6bWPLDs4KrR/7lJs3OZ6ckoTMx0Nsb4gkWbrI
NP5403U6LY9YAfJ2EbTRExrZZQf7ycDu5/BQ7rf/4F9ueOgJbKG5/CfwMb1mVAzMz76Fe4vVHBwR
yHgWKr+k+GIcEsAKl0iDEyKqM4O142KyIEH9B+IyubTRMbVE+A9+6fr9iYUWBA9Cn8QOb4PMUHvF
aJHLOCggxfF4f/K1GGNvtdt3yqHoAIHjqkzTg79bGbRFCbCmWPD2Ow44yi3adkPlcZ+GpicS0O6O
BAsJ/2UZnKtynBBwdAESCmH1dpS/s3OG1bHbpb4GVpHiqbtb96OJAfTFWs2keUrBoYZlzcmFqRsc
I4yvyj6vvK1appGvVFcHZ7LmjTACjhAPqw78wPdtHkS3pQib6NUxVPonyCF+w7GBnJGbgMXRtkWn
lYwKwVTcmT+ErgDnoHWjnbOXzqV6mIC0jmcdMKaGzxp0TePd0vlfd0GSbvmNCP6kuEUz9zAcKba6
kXe1OpvWNBnWFBD/UhboCnWZ26goaH0FS2MSW39l2rhO68oM2tfIQqc0gZzfU3AJ28vHbRxmwn1k
ekr5xac5yE2/GijErKgEqRUdHI+wU70L7kUKypXAk/ueO1ObiLvJLmoock9z6OkoOsPqlWafg3P/
lWiFd2H/441If+WhKgI4pDakK9ekdyc+lsWb6ubaK5i672snd8ej95qnNqZJYajKNX3xvHT0aaah
m9fhSEj2LdhV5+Yku4eOH5XQJ7hbL4Z+toQDHYKGdn6RHWCW7ndShvPtqD7pdiTCUx50Cz3Sw7Mw
G2cgVSe6FH5Y5wYalUBrrguqMKcdSy3PKOPo0A2aGRh396TMiPoa2E0fngCbJVj7ZBzdkm3cGOyR
OVdCl1vnyZkwwQx1sbtSqrlZUL2vWYwYbMoPIYY5nIzRsUuK0Mkcq7K/Ob4PCEaO7Ys03sg4AKV7
NE0C6e6uvJ97QuNyVkHZu+uthHSni89S/6qOoe/FUOvHcSEURWbtFmc82T2NzzEnknefgUsTVHD6
5FIuVUnzVujYODY37S2qtZ/jcwvwmdEN2m9AQESzgaSuh2X4SYnSRx71iqMY+6HxmtTn+qyyz77l
jBs85u61xuYXVbAAoFgdxU6HhlyM/NhNfkBoQNqHrZPdD5/QJK8NrFvEwfOrvy6/8uOqgasM9idW
n8yRbWoylkSWZTqZnO5bhPVouAcUgCMk2ItxMlRq+SYgFzzh1pxniRLsk6idvm5EG3wRtbFI0/eq
Ddkfv5qZJF05JyqlcDNMy4pVf1k/Xk8ggmi+qUyqR6+UvYNE4mdLaKKmRtSqAUSWvgAyzqro+25v
5p0OrYpaEJHuhveiiiq/4XmTsmA+ReuxNigzHXn8+E7e5wnG4Ib9eeMUWVzBJAUtjzlY3WkUuijh
rvel3JnLOtlbxnxI6pRlovMj8WtBXi41Z5QweN9C3aHLY9CBoezZdxWj3JEarzr/mkB3dyFlfHH2
7D3bVmxBPFMjmIW53m326gaSbIZ4ajUn/fYgbvwc/Q6IuJhCgJrL1QE34heXstCe6+sviz408hJt
FO2j0KrUgEpmyzELi8mMbjfXLCa3fpCBBdkxW2Mm5QPa6UORg7Z3lRg2/r/gJDcAHTk1muc7jgE7
Gi8W40fAZW3qv6fuBDkj3EJQGFZP3SMGs6r+5LpHmUAY4JYX6M6oYSW7cQZgntnQ9/BG+RQqvUDC
FqFsUHvzzKdh7ux9F5eeCaHC1IabR7VLUYXjhTdijQWRBH8H9i/dcc4EE9RmW9jzo8Uv5zRCZHCO
lD2m5fg3uXit7Q71RgVH9f3Lo2D4yPumhmFBTvZfvSArOz6lp7V8Tc22EDuQZ0zmbdXLLLUbIbAG
LzaRcJ/PCjlOf4D53zWjY/7FUZNOaB/7ZInM5RUoWBd456AJlhepR7/jR33kMAC0dC4ujsRDVwtW
8X23yhl0D4/f/zcve8NhXu1v4oQ3FD6nNRmhyMPSFaDzT2WnW2Lm3DAvN1JJibtLni/o6cXRuleC
KAIHo2kakQOB7rlJnO5S6v76QuOjaFHXY72ilfJUEiFv4WsmIBQL5c2ak7a6qhJOEklsE4moi7h/
FqjjbtoL4BBolGRsPVKmostdtU1z+xQv/rC0CG1Wr4nSLuvMmXdMINevlte5ctSnDoJ5fq4NLyKF
VzW7M8WcMtj+7+qjjcJritjRVwQ5Q3sEJxKvqvunRCkM5VinDb7wlNsF31v9St/4POL9E8mrU/4s
lQtK1TS1t+zrXcykjNIch7oGM6zzOV11T6e0YUqMCyaNVVZIHFwGF6P2uhSL8+MDkU+UA+K6DYtS
iWCkV87f1E6f11xb3n9AzY04hmiCK3M6jhCqy3CR4zDWhxRvv8KTb5jUcpRkutoMgu+lbKs3kFOB
cfUOv3oLFmynn3arY/JJI/ulcVUzHKruxV1UNlgeeg4yDptAukatHH3y8H/UZUXzePv3SgrbWG28
FtImsNCVuzkV1j7XQXr6IKemmOh5JkMinoGhJKwdJt6h0kFUX3zvBn4qPWXjlmMbCfAxScs2HQJa
9cm7fR/VAaLQXV9z5KC8QZq56NOxyClHFiI/a3nRK8M0yQxMYCtkqgWmz4tqkxxsE+WYlPUTTZ3m
taIuLJLpaxL68wvLwEzPXhXxyowUgU7pT6LYXiLMhWIh+tdgfOtdAU5ULyN0NIpzZ0T2ch0fzi1T
sw3Ums932LGM4sCjDYURsC+uWBIUfP0fs7Zk0m12n+olm2q4j4MXqEfPr3lyqd7jFhx0H99fXeEa
QOoBL9Hda/NEcQJgBb7rSp1x6VwILdQXTBB1HCzlD7Mw7hL6vrV0XQXdijdcn27mTQtuxy39jP+O
H7/AWM58bqVKCx84ZXMJWpBNoXwMOcpV7EJ8W+kqhymy4RiyezgFhhHs7D95a7uFLaxBXmlDJFAf
s4nCIsNV8HIFAhPP6yjYMbquiyxxV59FQed3xOMCEnINe7mPYXADe9mHrbUqw81f5LjQ0W27RwRG
4hGoOVMzh6wMIHwSYXc/2/NUastj4BYFYJza04lMpK1Sx41cpoHjchZz7iHHzAJguCYTE9dGT494
jkRwdY/Eqpgt9yj7l1wr5+bVv5ko7R5VeT4rNuyyfhAYPLpUbzX6e9uBkzqBidea/awUGTNoOfL3
W9LbGbAyXnY55xqB9aS1PqPNrHigauDQTgN0Y97our7JBXMO1oYUIkfivlaGSp5zoPnkA4fB0vZt
gvAjzklQMfyRr/NC2D7zox1XIR331ZKOltdfjpFzipKdntC1NGRcESHQ0nJoGFboK37ZQaz0Iq1A
noma9gr4OuDsqNUc4pH4f69d8zVtzAiQZDBEta3/KuH1MTceJVKkuT8Bcx/exbMouNTpbyr53vma
JgonlGsgBbWJG1/851p3zazRVDY5dMd18Oor6P1TZ7EsLIpGKboRFTRGbEvHrRbgejXo6jA8xw/t
jBRvkkAesG+jTvL5K5ITBhfVnArc4f+QYVwcaF05/4XwdLrzaz9TookqzdRBOyFO3hGX9Po22qJa
xlTVkx2Wr3lnWo6C5oxFV/YFk0akVSsXs79NoJe1mSVDmebMY3xaEpjGFfSdHVTp20UF6xsX14uF
+fc263o4MxY44QWfSrFnoBCvZSo7yUUT6LwFu7+bockK0ZJjOLoDVQshVwTIDqLIQESHTDpY1xMF
UrQ2BhrHX1cFzlWvQop/PzsDdlZpVVNoywzdlVPg9XGerENZhTy5oWWuWGVrXcUX7KEBmIlty0Rh
7mZ80BvOgXrWwPU5IMOWQ4VR7aBuwV85eQOnepD/3izFkWeZCTOv0LRYo0ceG32rClrYo3sY2sWH
tyA7RfKKU5QZViOjZWBr9j0DlR8zNyYUF0+JnPnFBXpNw32bij9GmgMxF3Zl+AatN3Gx7U/LnRgo
1ZPuWwBIdH/f43LGEeRX6yD7NE1PTH99YYVXY48ZNmPtCV0bdVv/6uPLSeNQXWSuT+7+zT0rwQdD
+kgyIXygL8e0/rM+ry/dCOf1607T3P+MSc+Qez9tTCjp9Ecx52F/cUeepvE8GsLh/c/29D1TRNqa
tuk6ERLdDkSt4AKg45MCS5BueVgLLb3zCI+4TJ6jNoWFB/mIipDPr35dWeCzJmxY8hnd6i/K3Dp4
vi9qbClOBvxI2VWX1mGO0+MbksOZx86awVRjVQ6DmQnTcxzrex32Fz3cbKnnrFRm1Q+D1AB03jT6
5huCmkBCIutXE4M4pcyDnpfgrxxgybpi6lDml+UzqFtNkEX8jINCyPX4odKJEdNS2KoGTMapyxWw
3c9fAT0c3ajSqPZQM72ZJALZIwxDT2wpm0odZf5Zvh1yKhI38ecqtE3LPfvTxg46yKdowO4nUHHf
2AttWLz3iu5hiDCGTGEG2nZytcAW/Av6xBPjmm/azy+hbcyirQQs0SSMEpO6J+hjzovech8lRbHI
OoQZFULKVRkYJEjgSZF6tNGklm0rGvuruUBTKwFb4x9M8OwKKLyX1qQhKtaE0s9dR6mLHlFuLGtt
uK9SaYWpvAWSuubrmBoUnbw8fGN+fs5hTkabA/fcxPZalqyreiQ4HhRDEm4BJDeEVInvYhygYtv0
51Izs1QBggFt9pj85K0Yg7tvSgOEVBxDGWRROTuwSfZ5ZLdcEcMF49utjX7PaKFkgNgSBn1UgfnW
trx3njyBg37IH5o/J4ywENKWf8efprwNfJUn21IQoirig597kH4e6iqBXkWxWeSqeLWb6aaNrUZS
R8pcIstKCna5yRBVBLgRJnIgDQjnIjZ/Db/v3fZRYklrFxzZQtEveSER0Pwb76ufYYFTcDvjpLyG
ZQTF7iFLI1MocFxVXeEQmb8ML/MDiJd1DADefEflaQ9124/2hASq77xVkJMczen+wGIQeCyKMiSv
ceIFX2BKICd60PzVwxLeCCVtzRaZikq+PakTdQ5Suty0mt5WxznDmbBop3pHF/EH7XzO0WCTQDF4
PU8mBokeB0Csqhh99WBnA8xaXXnji43syzfji3QxXFKcz9VKJn2DcpildU1LYw/SwsKxd+xYrbCG
0rjm/eoFeG3BRGU91J5ZImDf4DlqVuiqTMU3s2wy4KePScYsAalvR6nOUi3OOKvnmTdnLeWIKLu9
K2Prx9cEBFO3ssKeVLcWl3JgmOVwglqsEXJ7NM8C1J09rdIqfFGvzwW1q9gtM1IUdhnlCTPo8q2S
5c9AlqjyY4qJvXv7G33Q+L0pMCGaG7Qn5+xiv+Pu8HMd/dmRZPbhFEtVFdTgi4o4+7aqhruizbRr
Md6dE55Z8xNk0WktMOkZrfrsLZNs+EYKX+BX2I075l+HIw7Xo5y50gH+NjXjerEI8O6eHXfzQGGW
b2QvpicT8Ny3vPzfngTy3ddVJpGGiHLgA0YK1IjwtpI5gohDsQk25xNAbNIDXQuVyT3IHX7cGO+y
M1Z/y2SL1Bnbz+sPBBk+C+Kw7D3Wu4Ijr0DEZC5XmPYER7m2WfrM9VRFTeIs8FGHLnCYLwOFXYuE
qlgqY4fDV2Zy4vfJ5Ki4E4NsIWChzUJ6bmY8+nVpWI30hxdZArOaOt6KRnMwoiqSuzjhcT4sH/Yn
6VJ4uXHPiRsuGucaz485q1FA2cQZJiK9tbEzbl2PcWxaJRSKIH55mJXdwd50qhQVeyJFKj/Gk/G2
s4rfA+ljS7BA/4br6+F/VexSFQkay/d5ASmwK/CAKGk+cwkxYjo53lN5QhzDAHd45yf9BcEZg+wA
41pKukyfGlkccTtvcJUYfwE4bCt9wBWy/0K1U8A+2aUYTsshPHulBBskC69JpT1MVNWbjFxcXQMJ
72MJn2vo1a+GJX8fvAM3Vkjnl8hA0Tpa+hHQRYfuKFNBm/aGQXdYjHvznHNsRycF0e0GILW7KzCt
T6m8izS8h6ILd+/AgrOTJB/nUK9539vf5F65ye5yJ/Kbl/FzS6uW6hZO20/NG+eTeELFb8PDyS04
E1oencvSKwjGdmyj+XNbGVlbXtXIKOMggy6W12a+8ie2lN+9pfZv86+RLaPbXWK/FBr4gtC46n/O
+/NUq4qRFDHiUBinXhsPnzWS1CrSXQK/yJq0AsEYWXV9v8oucNYnKXR1Tin8gdjWV2/ketvfPTLW
/PxOPtNn+7csP6tKNI0amyGL+o+l7yN3YGXLF+GNQWPf4HtrZu/Sxihtyw2FgJ8HeEyqvPDJDrG8
00TTil8Ad3Msb8MNFUFaJCPCJEukl1YJ1UjMSVRYwYZQargpEQW0b7REh19paFYsxErku+s7+qGH
Zu0NTRzO+ALSGfz7axg7xj4i6QHFKwoc/uDS+05/LNSEyQvIFeLsB7Rupg1K2HQKE0pC659FNH+N
tFeMPpaBkXFN0+EWWXJMKIgMCY+IXLXal0i8Yx7P1CPBiK2MA/3VO8LxCRWqc7A1YH0vUpM1fgDc
AlMF5NpTjLPA4pG4w7RcqaTp/9Sfn1iYK9dgfCHtG+KF6ehwO83eWEGn4OmpUQtqwnULLM4lMBVy
436GUnKs3pEPSQ0UjqFLlW+9rDB29y7xs6XiLB7B4tEA6FD6ZUCflMp2kFieJSeZA2UOXQRWPceV
dLaIFKGhUm47PTnc9LBF+JKvCqsGCY2RcNT7gYMZguy/TLeV+q2O0eo7A2L2ZiuKgtWPgHEhKcwz
yQDK+OSlHFo7QOdZtq8piFJkQnmfsL7fvNsqWKDMB07IX27TtfMVDJyP1+nHgqebkRXUtu3RlKl4
wEHsZE763mLObApvaRpGUFjguud0jeEKz6pOVGXldarMINgq5MihAHbV539NSZmeQJXvkYMYj7Yl
b9yzPlN6TiUoY0C6DZvY4+pfrEw9B2Y3HDQxbg+ICb3XsZYZDDDBxi3r/0e2rgclnEaW8OtD3uTm
+AtNwOezDD0UXfvdvnSRDzEcYXcFB4xFLq65FoX2T8r0fFqSjS+C74S8ggdpVwCDiMElegRhbcLk
sCq6Zzk0DIetgOGq0m5ofB7KWGuJgLdWzRUSI0HtL1w6HlEZrCHODimVkTIbP17pu0GV44MKg68t
K+lyXPtdn8lRqQVbCJibHcFO50wbylxs4KP4prKFPi3chjQ2yx8wS/PfV1xVoZ1h2cTPiyu7qyJH
iPSJLs47+juSWiC/HsDBliINDkgEBcuaifJ2EWFlCLNdvWjSJnWhi7BYNNQUZ7zy0bYy9BwrovyO
tWYQnxz8Gj2GGnXbWfn+178vpyETZOUZsEyifYdtNL20kLM0u3hkGU6bGOPo+miQAdkYkZyNsPGi
cEbmYsvBfd1FFEB4HzKcJNbV+kqr/9m3QF9XBmGK9jdTZHQ2Eb7fj4ejmI/Du1hGqHTFS3hutSiP
1PtnPp9s9krWKbnOtZR3O86xt2HKtKzlR5vp62aeXqwljxUcGe/bOT61bhzfOyKBb35PQBkZIHWq
aNdp6HunbvSBkEl7CBzewmW+dnN25CRsoI7rV4yFnTsgi78pfaKDtII6qPlxxlzlX7rurQc6m6eE
5x6WMtQBlBbJitck7Q9bxTwthgk718ojVsWqI51Q2c6YBWs5HR+i2ANnseyiZnab9qwN3Cn/09Oi
mhe43wJxay1hw+dcEiCOnhB9qOxfphvrAMddBQvHeFSkQPF/phJ9J7Ql40Go7lqTSGrflec6ibt5
L0gaFZO5vTOeMKnPOernM4mh2fRLJ2s959Xhs9hDMouNkwP1TuU8ina3OVBHl0tdYctW8kYaPrqR
z301n5TuGArPjsCe7WeB7eIvCEArIN1vJZfMEWsLrtJWm+FnvFoP/eMMGXbxC3Wc7btgL1tiASZu
0bI49xSZ712Q49wbMFtPRL5KGCh/KSBNHTeQ0X3Ll6eDmiJleWZWhI0pRcoiWWm914qbh2Xb8riT
IliiHi8RibM6+Ls9huIAZkFMTBVGLV/2BG+vzy0PJq6KO0Tw+oURz0DnLMsVXyBgAv3kUAHIDxxj
sxAZuvEe+baLRGjH0QQrdH7jVlF1z9FRKyVgv80kappUtVB81BL/gV1QovhEYHkGVp3fi8FNIe3x
PZQNewQs7IyFYfgmv+YHJb69mABYKXTYoM+vjbcxH2F88qC/qYyvfVT3deYtJgxbUas+i78C67/z
PrwGMdtj/VIbuAQrg1RVZ+IbqevuF/DYDucT1PvrLO7PCuKlEWKJucKUsj2UH1EDPfAQym0/PmxC
qqnT5Gxaho9/lxSZrQA7dW5EENj1ZXMZFwzY54LeFKxaW3DD4sbmTfbWLqAafjC+lfE5ef+CGRcg
Ju5ibQnz3iQAKEE/cf64vi8oc06fNHc2jfJuD5yuySEnoI2ByddlyrXMr8wio+hLDdyrZ4C+0yrJ
T77jtFKNxiJn+/nDxkhHMrW8p6s+AR1mnXVCk8IoLOnEauOfetOagIJ2Roj7q/pTyQvGZYjRSdu3
AWAD+r8y21ZsQNc4HJM7Gzk/5SVLE7TPw0thGqUaP2ulJbXt/9ul8D+cR0Lki1y2t3Xz51O/2AcF
+uvkhvervjf0ECzgvBZ/N0/1RxBBlswfS32CgxrSnnpQdcpUhVTuaSwYxzd9AQ9IYWcjYcX46Ita
AHIIdAxsoxVKaUI8Ao+E4cH/5ToGTM9WyK0pN2w5pEFBxxUr8OQENBxj9Mg2uEgyNRb+BJyUCMjt
K3MiPolVf3oOqVZgaenRVeP67mQAtIddpv65sJ+VuQniF/AaewEXjyErweCtg0oM7r1OKSo5vHit
OG2H5UmdFgtJQ7LCz9n1uVJYca3KcVj3kLGSUJGL0pmtXlje47npIE/PIIZ9/Pj6vGNO3f+OoY0A
kF4YkUCzJsiU0VASkrJ7RQcT+SpPL2Y6PtDGgGv2FtIiGQdO4TV0O7D4EdAEuAkMXPEkIUXnqt/J
LodWf1HsiTokIsXcl1wC43SbP90iQGr+YQJTcGQY5iWw9g11tEmLwaseQRqncQJD1o1JtFWBgqCq
fjXwCCXBJ8rFI8oYDUqgklahMVyQVSOs69syDb5jrS9ogZFzVAWBu/liipzol+2nMXNtlr+0pjeh
CDX6m5gz2kBnDTfHrTrIClRkbPw75znzSjCon3TzwsCEZTVTWRVOVCS6cH8+RPYv+coEtz01cVRs
zNVHoqeWAvxpe0Hd+6Hfud+mKd7D9IGRkrijQ6dcSnbpU05glTLWMa+SMqLUFORsZ/r45XusS5gD
0epN8/ul1XOSQ1ESzVordrfQXz4C66ArVdsefS1gwdHOKrJ+ivyubIE1dAFJcXWJgWiHG1gQyEWa
Q6g7CUMItJLUgqdCrRO45ohrKv+S9z50vk2imc7wPynoIryhura4ZzeMAmgLxCZaPogwjve1m/vp
BiuZZKWvGTBztMVRBoLyvw++F5ezRq1UC6puJvFPY1y1qhmMt4p/2LOPHF68109x1eGB1J1iwqrK
ryIFUeCGLwcsyZT7cg05BBQvABMDHIIugRPCo7BmXE2p2gSlMTTxNVliTyLAVfL9zllFXJ1nHzuH
QvpoqgFganS1XEscZ3xIjrXOSLL2SNYh5ZB2cIx6TlfKhX/yUjftKc8sRs1uNE790vkDuGQuGePe
XmC/sDtWWiw/6fPgaZ70qfn0cCf7ITBRzUw30J2bbIYykBxYGboke6YCFtdzeGInXt/HAPn4HZ87
B8Oocz4ZTyh5I1ALwgG2qAONXbbP7HczzppS7vKynNEQu2VMxMQPha8p9TyIa2vl4/iYnbhvRJWi
5mTD/GzQKwFC//M0A8kBlYimfb7yA2/pa4Z+sWJlk6CmbiaOm+J3qQqHS1ctxqOem1IfVnsU8nv5
Dg6NSIpqhIiA4awhOS93wfk/bWx5g8stg4ahUWkgD6o6a/LlBBV2ncBsvZA+cOLz0trQVEvfRs8n
5q5mqQGvusdTXlGOAHY0bol1KTtjvDtgxg0uXd/1i5e+/sGKNflWzMZEEOJmBke6GQ/WQ5zAAmbE
K7nJLqpKVfQDm+XhOtV4/8EjKXkD0b0jQL2Qa7CT7KymO8FEZH3ddJpML5QBve14pnQYGYu7Pe4Z
lNj8LAEaOMUSEb++rW0CwQAJMI3xKp+vON3K3gGXAiirzRfMCZHO3geC/yBuroMGzFzA3sfNTd2i
uavhUMVRfV6JkrsJKfGZD/LEZ/Xml+ziUHjSYSU2y6CSJ17wQnQxrf5bhCLrAIbdRpg7iD6H3Ihy
zUye8x6E3FTMK8NAnGH96OaNrR1a/BdDnpjc9z8jxySV+Bn2cHGzFownRvP7PVGIbvy+kdRrf0Le
napxMNKgiqSwj0SOLXn7wYxi0m+EbQGp5CQNET/e6QFMOQciLymCrFcZtWQu3Xbf638SHjtbEkCq
hjlNwj79i4qev3FHnUk3FFabrP01xtM4F7y9Z6Cnr3/JOOc5E5s68h4Xd9eogB+53myrHHerv15H
BanVqkRCiTU1hH2hB+2nNHnMWjWRXQmx3lUuoPC4y/OjXUycYURZnWHTb8KuDXkDEJ72l7N1dfoE
6WIJJfI4GwtZ71XqO5cSVa77oBGdBFK1dS/sX4nnjOfzOt/0h2SYlacCFp6kxB3KYQqsDgBYF4H9
XiCo16RL0OYaXfO491mvHeb4XVVOStLIeX0VU2p5Vh1OqF2GdcNS5n7eh5LUFRLzEb5ml92pkusA
6d52frFp8nWVxY24HhmO+xQvivyVJ5daIiOkU2Da9d9EbXH96Sng2Tg/flB0TI/76/5XjvHiqk/5
KtqEwe6B63oVJKqOXo5ex8pwpkBdhemF/2e/cOgdcg4XF/NyPgnSobv4XFDOxbrT8NV5UK3vjzd1
TZeQhrrYEEnurpACqX76w5dNLPfR6yekWi17ffQnAgHYpIUn61AFrz3MnT7gnCQtbVl/YV6ZKsJl
JXPF9+EupvoG9OHcISWriHnzDLxHD3Y5rqYgYIDGbNuw6FY5ffyk4wRvujD/ANTisx/9eGFatnfM
tsluX+x1xZaDBRtbux8gC483xggjn+Uv97IhWC9fg2d71ex+oxd7lDiUPWm/Bm4J8xm0D2W8w7kd
nF17ML8tCUbydkIvYhvL2iXe9LxQ6gw6TbK4MxMuWjCcJFXSlFS+X80SDwKMJb8hqdS5S3TfdLeQ
iEO4yP+JJxePOr5nel7RQVpDlHwU76zdYrliySS4PyIONg3/X4rGYOjxxVAFGM6NOhokDL7BjNr5
ftgA5mxV/jQAGTvaQad3OFE7dmCJyTan8BI40OtQquGnaJ0PTgbiZFPeFMviI6N7CRRhvM7I0glB
HLQ6Xem0qcWXjqtsdJiR0MoHtypbMlvevAMVwVyhbVPdbFpW6qewEWJgl+9PcmLFjQ587+Lzv7I6
kC4U8Kqxm1AfDATUMzn97g53k8+umcGV0obM2GbHovLYtBRzCLzTJ8yndVKfcekezOU2CFIGnko+
uS/GMroHzOhCUmsvD4b3wvZQXdtwgLA7ftLpAtWRQnr11BYF20SY5ZrtUFub+sg6v8PLhrjG+yw8
Idf5l+qJlt62DGahAi7mx6BtWF9eKkvfQox1ZdCjaBFfK4gG0t9nW9ohIkCTNaXkIIc2RDWB7JVP
kSM1B6MT+x7iJMFiXfsn+FuR85Sh9YEwx0B9Kwn/6lfe7pfIF40MGZYqXNy5h42ZOPv0eiHPLe0V
5w9QMdk5TxjNOiXamQt8fZbBYzLwclwIqBlcdEr/d8H/dIjghCOVfTUJigmq4VzsgbO8OKo2p3+5
X7YSrGepC4uMzXse4XfrCh3enWc/7nGUZZnkjHiwRlyh3KTl8kjGitsGV1n2Z1ciubssW1stLkAN
iii5qkPOn5ghvrQtoFZaonavDvHUoUoJgJN9gMoXl5d9OWeSvhjUC5rNlqyZR5THoZY0m4uU7PiJ
IlsV50jmAf5UFwibLKU3IcMD6M4tvPeuSr4wCGiciO644pIvBdcQmU1VV2y+JcEiN6EUPVnsp5b4
vtj7G2BOZkF0eii8NvcN9fHj9R8yTMMUkWM/KzqpxKNcoGBmdfs2kI9D7awq//9hF4cpMf6caXn7
s887H/Jm/bdXm6vkG93szymH83nh4R/8AbNL5UwEjEVjq+Ne7/qq/y1l9cKRbPLGJDPR/3O/zC+T
vWOlr5cD34TeavvMLwYZmGc5S7YooNSKkfQ00pyU5d40WGreXpD6NpZCSN52urCkNUXNCjw6ubzO
20zNzXO8OEWfgoe0i8yDfAROOsJeeztKVafpn5WIAg2cF3p1z8myMqLMsitMjTV3Uos3/wrV6cE0
jyMM9foFLggrRP2gFmFiEXo92Zsns4GWrvS151Pwgy3WDdks3brnX9x2USdT2/4mSjbKbc7ejpdf
+rU+BqLtnqX+bIP2JQTW7bO6yuOt4tMRv0J4Y3P2FALn5mRJ72M9JwhAuaqBf2Es0KAmFp6zZwwU
TgwDGr90kwzLGooRikJY5ZO7aHi0HpXjkkexrFLtfQ9dcA+Ga1vL31z93BrcmIr75XSBJmlbnB/r
SXAlMO9mDNr19Zp0AAmVdg6NCIRMsSJjHozOl+NoNza6Gl4R4BqZHnoshlGogh8ktN8SIzFX8lz2
BNbqIQP3qep9mTf7Yk2kXI3sq5m9nN8S4zaDCP8I5BTn/8M8cp7ielAjyujqOQ3bHynr3PCZTfRy
OZQLYIQ1jZN6hc3K1TbhTXwiWG5MFs319wrGJ7CEyB2Emp4HQwt5gh3Q1kv10ovwgQv8czzp+r5P
xMIL+BBWP6WGg9gu71c8FkYY3PTEHYs86ktfZPAqQAVqRrsuAY3AkZJnuywXqn7PJ6fB40df7T0q
cZMZ84JIteH+SNnXD4v6zm6V1Lmwtjlr+xhWqi2mRvAC4r1Lzj9F5X31LPDYO09VlnXwOPn2nb8Q
NtIMTDPLfNCdQcTAXgZDehNgzSGMWVcXYmuB/SLkAMrfXbzxhgrI3bXso3pROsxLyvhfq0T5hVvT
+qaGhbPbXOfUS7EdtxAZCJ0162PSMuDHZNjvOflrTF0yNe7tjDQviGoV0E6JuHSfctYiQ6mtWcKi
kAVHMLQau8yy9+0bWQEG+gDymfqbhRybXSugmkTT2PRFjbLejYL86y9hy6N06WO/VMY6aVF4L9M+
DHVLg9NfmQOHL+6ks5G6FwkGaSbHWiq+CH/3/2C8Vw2u1mhLEhSFjtSYu6sGNpg1HKwy1rSBPcHw
+kw+GnP7Jbrmucujd43/5SOYIXwkBAWo+naUt4xba+MYXweiK3+elKvHy/2l0MVW1CQyCsWg7RiJ
rPMkGJQaQXflF6MxyvlQDPSc7cwyyUAFF4tmVardxC+hJnkZj1B/gNr/qb0kRV/uzo5NMGvuUFo3
Bt9ZIkbH0H0ht1RpeCrdQwboZmO+LeQum1dJuj6vR2XdncHEHBotOUdgN2Xxp/R8bxcJu/IeVgdC
50REqOh7ow4xYCdMzYtrKOvGraV/3c5OvTCQWS17Vw5B8YHgfgLeRwT+w77+DznGUNGUX8J9PS+j
N5HOfaDrEPZ0We+61A++FY2QUVbg4taj3KdeDD2iedBm57PY2bSPLCrkfSi0KrsmTu9Y8rfHtVA6
mMG0Cc+ZLQRrCEGR3U+FhyY1d570BZrC/3iEUieYaPOhMuJdg18bQSscJUyBDyAOl38V/1ObK+cd
rauKzhtuJiMR5gTXCDn6VGOHnQlbVFf8UWv5Md9gSGXN7SzpyFuTIPGnW56NzvlFs5MEix6H8kRS
9ZbYq+SUF+a+pk/G5Xd1A9tNphhcXGQQq/7BTaEw72AKK4PRf+c5ngtPGZoIzo5bCjtB4djrLi+D
uYzGZEpu+7c2kMvJ4Nq+Qp0fAxlbSqNhmVekOF+YOE9YzQvXHBRe0nDWKxnAcD6pjfNAv5FYoL22
jsKpPy0oj9BiR2qz7MGLC8VWM2FSr31l58BCLagI5+eM/3GC7XtttQqNfI0AxukLiKxS8X7Hocdv
swTBF8xKmwGPkttDQhnzAqWRXL/Mfjv5cnTa46neLnRZroodtn/LMnHf1xYJ7B4phPU7GGbwZU3I
cZNDvytXqbg3DgfCErsBKSHSag5L/t5vJ9ib7cgJZKSAh8/Y/BOOW2ucz3mg0JcSTqJccS4Ow0tu
mG4whNVpXPYpdiY+ECvN63HH5mpiW79uEqmMiGVbhuWjdGwZQmhazL3YGz/3mNHBudSPsu+SUN58
OkyY+oXQMg6NSx/YQZimTfh6BR72xZay3rBAyl+ATvRzq0WATwt0zCmXjH5GaDEFnKIUPI2eUaoC
OdBqTK/1cKkNbAum9SWOUan+KyznhxCBQTagVLzUplQWRVDME9muZO45DmblDbTz77o6iDidNoYZ
CNyD6OGGNWv27HDtc1AemPCzJvssbaDCKLd1BJQA+avMTbWXzpkIgA3+1g2JU0kvfscZQh0uue1B
WTSt2o+xUFcttQH8dwWhAgGjiSZZqzrFM3SJx+O8oBhY5LrJJSLYIGJQGbpK2qJxK7Ql5TDCk6by
+lEL0A/fWwPkiQSQF0A+eZmWlczrOM0yaYA0TjKEn4Q4VeUqEEVqzelmaLqvE40PQDGcGAs0UG0u
z5yeOL8dhMI0AIM8kdjbBjs91SvWoykoX8o9Hq5KOUFue909t1YiJ/WBz6q3o7d3Bz+I9VESiXM2
luFW+dzwvEwrk8/5Ids1Vsm/72rt/ka/moZv1GBV4G4sfpejADU6S0DZMaBGYo5hYDg4yxVTC2/K
YtipO6OXVe8gI40bDtnZ5LreUA+W49OLl36CPxOUon2xzb4FYss+VxVTwe33IZucxKA+wCqudvGr
zztUwAdds+pKbDiveBS2HmRk3C/aWiW2C0lrk4yDEzIXmyeVJ/2MNBg3YwLIAprhg+UZ/F2k+l1F
Bk57m7MRAyw8IVfWv41cMDQAzklMORZiE7H6QqsaKTRH2rOUOkO6vGFum3/XtfdOtfFcXBglJQ26
JQtZYYM2dpznJDJ/Gb2BMCXHsBS4MckOziousM3i4cZwBVJHUUA1Yv5cXxmnuvC1LBSqCPwaBjqf
p5O65CDSHz11gFy+vRABCqT6Z1ehf2NrmkTnpa7J7OemDsT1QOE/NxgW4hsfYFh9wSGbKsjx67IX
w4K0xkXWIa9VXSCholYP4D7x2skMpag13TxfIfovc4CFhY7JSbGvQIkyfTQQTuvbFpXBdnVHDdGc
JDH76yR4FrtisbnosR1yQ9qZWWNiqQ3O89Vx4KHC1Sriz+UzA3f3sMaLg1LPwWmdr86wmQ6PeSiJ
Slhnf/zfI6DhuXBB5I0/faKhugpBkoea7liWyFZSOO0tYWZqrNF8LofW8jSk6yp5t4sU5hmy78Yy
J7X1u2VITF0rFjiBxo1FrMyVjfoQLiZLaTKohO1ur6GQPjF0prhkuxmrVlbdPg78rKt2QaargHhN
ppi2PYqmvRnKBFvqTL3a49pIGd/RMtbRC+dMMFlJ7iJunntnhk6M4lanLBurrG0CFGeDQyCZFWmq
VzwKXoJu8Zcm6oDnwrXzsegNO46C9IkNxBSm/9u5ZGxjGzXcRMYfT/Yi6jkqK3hOtvbq23tIDyYV
PBl8m61GWKEKGpuzUk+2oEErqPnAfIwj+agc/df8+LQrN8ue26CPGpxlhEkhKR/A+hr1vduWWK6E
hfofjYDVm/HN9MwTMwdAVcv+4h8CK/bDw2497M1IkS91J/Wy5qevl+qBOO+h3qwSw7SQ5i9zckbS
jntF5Brca6qucxrzYs8D6k8UrwmasK1vw2IdScQUg4LPbjZR7GAt3EDusEErAbmImXiPLFDAiNwe
ZVcIaMscn0znC0ZSELverUvmbDW4NWngLO2joTryXehs6AncUBf8GWchyS8MQ09SaSCIhjVyULnF
hd63PrgPWXbEGWAME5i+tkWiBTTRr6jt57kl8SYQSUWKmoVprzsjudFmEbJhdEJn8UX06aFij7yL
ZQnLRSZPLyhes/FZzMgNwXeENFmj4chF8ZDsU1HEqKefdphQdJwkyg+8t87pudSDiCuwYWI41SXK
yzHi/fcAhuGNYbR9HhvPbUrlMMeetHSJ2dTQXNOToYPxhoPu2oJ0qogiPuv0iMYhfJiWt1ZrIMSA
qXzdd0CNeMf8+JNqMrCllp4u2hh1+e4sIqIMllnxtp/E10mBKytyqLdGnQNY6vMSOzQs+LRjRA7I
ydfz3Kv0CgHbj+m69Q1bwXfoZpVgmfw161REiPuAg80Nc3U/V79gpQYIV4EFP4XejTU7zr+ziGxU
rsIEVidraDkK43h8MZXH982f/Qxy0659m8/nyIZagoEdkytcR4weU7hHlpCEjmPYVRUHrHnVQXYV
Wtv6A9cBw5UqzhaKRfkGdzcliZNd4576o39Bl/b926awXjsOdEGcFN+85eDV00/OEaNWJsHp9I1w
9vcK+EMAojyQxbLV+mEoiGj7PzDXjbnlsQBXWIE3fYV8/FTygrFBGphmpoAVNo3Wbpl0zf9F5D8R
Bw3X5gIxNoFMdHOf11xGn0bMAOvJmphpNCYjCXaEEQFgxFKUWWuoo/v2xkHmToIjLvttIYwoNGIL
e/g4nVu78/0dfB2MLjoTUwdclfPqXnXvWRxKoPJR5AZFU2PwN8Re6joKddX9xg2gNwR/A3EZkPze
55KCM6CNwRLWgcTnv09Qg+QLJedtjEf4vdEYQ4yKjcdqT5WBiYfxFSnGcCAc4aX9T2m38SMxdJ5L
k8QZzQeYfv72JslBoYdDnc/5ly3sjL9oOsD5oeNpst8ZO3KK/SNeUDX6eahyGAmx0cxAOKwpEWsI
wOTakpQvV/xvO7+PCOnKpzUZivdKcIvow6ilIH1gWq21e1fMLHSZL2VVyUJ5lkkqyE7RwFP2L19w
Z7vbsbFQDkZRPUJ9abNXZNCRZPdbcW7+q2up/rDD8OBAo+rXTfMiqUvhda/1YZx9YLz4cE4dipUR
YBe4Vv0lYltRUImrE/xqB1nZi+3Kp60k/yOvbMBa4CkR2eBqK0B9UMPIhaYd/IRdfsK97fsEu1oP
nBNg1QYTsHDrYTNo0AhcZVcVg7yQ+qWx4DYKc5rc7/7qHuA6uUmGhxsErna8zZaRmql01O69Lctf
Tekr1GEewzVvklUEbfHDVajBbIMtoQLSFFTdXFcbZ9g5yjiw+95yChGisA1N4O+Gyz7IJ8aPb14z
j7Eumizcap1HbbtltWBkuFNyECigVYieE6TmkDBbqccM1npzgxP8KOR446xFNB105nDnPGVu//Xn
4d2tpRA7+r6AidQX7dHD2ws5NUDizevzoTdS3EQu8MyupggoyFDw0XMVKYMkmZq8m5kT/rmqTWgc
Uq+qFFq0qVhjkkfVuc7JusImCVH1iIsB4mQ6444yRCybMOBtRhqb+RWqg2eTZkKNwEVgRBhpyoz0
wXTOYDcladcepWzeiaBvTMG4dS/tGkbfcYKK/5xrLc4hLGmGkP1TL9vAHGLVUf9kqZ7RpQz27pbC
l0/Gl/uoxxkfDq6mf3e183i7bNp9Z8QWsqdfURZ3joCpgrY9JcjKJCNfanZ+HK0wv/70U60GQtZb
iyacEMOl898f9saktETD/JUwh3GzPMdIikUtKMJZtLSKeIjXIZBnwNG7KQlTOvOvNxpMxBlF9Gqv
uHH2T/4WaFFtJ2DEVYVGMXNXwNTMq4NflSWo5AkOy4aGBc9rH7vRkXaTmxszYHNtET0WVaeO87TD
8r8Lej1ZC8k4WvotQhuAOn8Wk0/QIG0otK1mVrCIEEuYxPal28my18Ia3Y9t28fL2twO/gMKu/h8
BAxm53fD/0+pAFcuYBOHtvhSyKGNT9SbRfFdlz/umMOg85uCrXAsNNZJhVsFBlCe4cEMVNGj20TN
LrKjFt3qpYt0SnSOsFc0EqdSCgOoIGqEnLKX4s+iFMUFmX+z0hz7fQX1sXoEGKRar4C5l4WC8l6e
3PrDFioxYos5hAtrmIhfKnWOavKzBktsFCrZ3P2yq6gcdbULdF67XhLimeyg79HUv8CMZCJFJND0
K6oKk5Z6mpGP6tZ22v81iMgMpyyuLely+uqh6MpCsW4jacyxnxtgjXwthnQ68UxxpbiPxaKmLo4c
HJM8iSkl9tT/Aqrr00GkrEhvjl9/KITo1jDq2TBSb1iVyOQgzaw/PG0haEvuM/iG+EVZqTbquzQG
xxhLsBtBMvwHWJpXF5Pq+7BVmZKIDSOm5YSCX8mmAPc2JZ+CHNnTQXZh2Q9v5CdGmgxBkuIdeNWE
5P0Hlsfv4C6eMBS6YyHNW2PBLuIEh3BjJcSn5DSZgi+bbRODPOivspcCy0UKJPvd5n/HxL8yuMaM
BetHXvybhFdNhF12BSilBkfehREJjOAVB6S5Na/6881Qe9X5+wg8LdKflk0+9XZR5laY2swjp/tA
onCWK0USTNiqI4UIdXEjJYwriIqMvdeo7/EICCmz5KECtQPUiEhJZJAFYdEhhH/99ip3/KXbFuj+
CjZr5WgrgMakK4PD4q8G/DJiWJ55PYOiCY0FKwZi+7Ha9Q0VqXoFFHdgJxvx3yR2zUt23EtmZKav
PPWBWo50iN3qH+CSJVFjjL7BNnucvFWx3VUaZPhpfLqR06n9pKiXywbFps3pPy8Oo4z/dYXaFbOm
kf+7EGap0ED0UE+dujhRvNHGEK2uPMVZ7C7O21NjFkpS7IEmttzYnroar4WgmzinhtpvjmORZI86
ET4YIdK5RTaz9C8KCXODH49tE9UMs/a6SUulwPO1MNnSSzuSmnda1MHyuXQU/Rc5hEhxp/IO9CvN
DGpN8ZXLRJfSPiMOlWNBjz/O8rRI27E/b6FpQetIB8jPv3LL1AkU6RV1P/d/6Mqqzl50lXkeczbh
TSRTd8dzODflDsTfvdqcOBQjx134Z4QPYM9HBkfXPkueOyP1zpd648IlbeJS+zHFq0iPZsTG7PUQ
ePxzWuFOlOi1FfU4flhsVF/c7T8N/O3JiVdVJ3XrsuLTYs/QZCsj367QQ/Oqk/FRndrv7uaxgTD9
WlgFSko8lwBOBJjInTuABeH7mTwzU2crBusYnYA5aluozyW8ikQSsvkjShPMokHnUZjqvc4EQ1mo
9JN1UekuFukgsbCtGP+pp+6rBEAEo6Rs3jV+2WRyfL/PVu1F6sUQTF2d5Wm05xoSXAW+HK+hd66v
yrT6+pwhdWvcx1CF+l3hsrVld0RkHg4aDw+wc3doSd1KauUVakjBkhgX1WNQStkT0XdfT3gD0bBx
Tt/gCb5RHfO7/7qwV3p8AXB1YwtjrMkFjbwsAT8twE7MBEChxmXvPoW8A6CGFw9RDaXJao58j6r0
6ldqDEVEGlewyfD6P4FcxemiDKj0VucgPsdnU6D0X45c3apPjkGI1nduvbJR2VZ6wN1ynu3LBrwj
USJ8fbSs3HzdOxT6fekP2j/R3l1SnWbiYsDIXsmsCBgoW9ZNte45Iyur6NFCbjzgGOJgnYzm8FRo
4W7RhJCgzvGjl/KKYZznN2H95I7JEiYV71cDb+R4EZTtnx0BM5IIQIdt779f//s30ZCPeC1473vF
jA6L1nAvKWF8blVBRgmihaND+DCQDXGnvApl6MOngTCBFOtpW7bxxN42u+wT5MKskZ2bInWNrEX0
eAhX+ddk0fCaBLYc3Ig40kuGYtK9P7KL2T0/iqXtLi0JV8FsFjiTeoeF5AkW5oAGA5XaEA3duDZo
Apt6jQwaNA3o9hB5wRXBNiyxLam3GrYnGi3jYH+B4rD2u4AKJkB8z4X13KxWmlF+bQsbyXlV4vt9
pra6uIo/x29V/Y8wDUPSPDb/P/t7jMrv9BdQo++OM68/puMFe8K7Jy9DEez+Gu/xV/1OdR5WTb6H
T/fhDxC7RHUBoGGCTE+/ce/jS0Th1KwVT+xN8MoZ5gqYFUQUxgRo9bmwQ9raq/0abibs5tIrv9cl
tZY62y2j0tif5l2MDhjdLva8Q3xRAjQ3sMzYQuP6hkjvQYXeBgs1K0+pCum58AZlhuY45Eny7S4h
qF60O0GdjqHvL5IHsP1+SuRvYJ4jAAPEOiwTnhnJpZD5cXu/0A0VblsTigEpzQ7ffJSgitgHQ5/U
qw6wpoLNVy0Lbqi3uAlJEJQxI2AHqQdLpfV2hUwG8HDr4bGHZ8rn7yaSoA1DJBK/LaO+EJtgVXL/
BvsNtXYz35VYnhgN6DXplFxy3xeUsD6J7luGW1MaAa+fWXt4If6RV1JTqIfmhn+MLBjyvuj5cXpI
08ozbmPXPL9Nt8dC7uIJ7XfskcjWtVqubSXCbEi8TJ9D8oSu4Y+EAlZ4yJiSF3RNsX+YFfXfUbVT
jQeMTaiNskZNeYlPev52CGqDEDx0K7fvXpKXosBNqBc+8xxGujYChILfQ5ejZXY1UUkdU4xzq3c6
4yjyK002M8FalQDPZ8smwYmqpGU5LN8IU0y6oFdNMHYglXvDOZTlx1zQu+QPkP/hivGR/ioZ9j0W
i/+x8+6GIAF2ypddI1x0PrnthN45A9oZ5VGZXjWp0jPSuZSBKwipBq7kZ0Jdhm99lqk+HUai12ak
lg443hoCdYRwh93Qag6C49jMk3V+1sp8tWgz5jjN2tEESU+1yU+0+BDFQNqUhORfMLKrspdtRKmV
ZbkCHkJr8seiNAe9gFDXlQxFNCL/xu1wmnt8+SKu2zB7TbEEqyw+8v0a1dPyt77RQdUiDX/d4tpq
s92uy37MOzGhb4JbImbd6lB5DsP5m0I5R16ppefA9WigJs2CVF33Kh11sh1WB90gOw3KV04yWJKP
I/wGigMh9FPuKON5QjiVxHpfkT2h6IbcES1cI5j5iLRtNnHBVyRyOX539Fo3R2zNXmtaHB70r925
swCGZAPxyo7XFcGUhJspKXFYQntXZ73ZyKEs8+qe+Oc/bitZ/1QcCb4Y4pFa1y8S9lCE7HcCNBIR
dJ+BDFahtPcp67L227O1CpLMAZoxPz0NYJMbBq1JS+7YdmSjD7om+i88qOj4IonMHl0XWaHIpgB5
xz4Eavu8zz1ergTy18qZGRDuCuj4A0uFc3vE6RrT7g/ItlGzliGSF9BT0lsxA7Rsj+WS+hiPrgNT
df8+qz5ufvUa6olJ/ovfnSjfQQeDNFOCpW7GVxtKTra3SeDwjvrmQWS1hM9Y9S1eKHtp07AquDKb
sp33CU3RR3Iusc7HPpizf6WdbpcowX5Yzg/CDflpDRbG4wNWamctmGiH2WQEWPOOS4yK02LVt22E
zRCWgEABj76uuSxKzr4pUk4o28MoRY94+8BDMcErDZ189q2HvzHbG+Rzmm/qJVhFVjDeRSwoBqPf
OTNjJ6EeVr6lpc/oPL7yXTIqH7aWmupqdpnbYnYWYEWhO1mA+9nFxrwdSX771IZa46SxNTur4jJs
B2YV0oWjesM6SeAtCv1M3uo/c4PwwiszGp416w4WGCpZxlThYW0sXhQBDL3sGSZLSk1wohZAqIe+
7akeA8wkjahLHqdPNjjA79FglVPUaBshwMXzi+K20KWvGhxpsdUzCUV3aq0hijUSzid1KxzTAVkI
LupUzIjCu73jB/s8kNY0nn3MkJ5xrkNHFOL0dExDfcCoQU+kJflLX+CoBTNfFNsrlzzC02mNmC3I
tvMkMjaR2hlkHxcgNoPhXtTsELuWp7qy3MB5TMJngP3QT4w4RrciABs+zZ1eNlZGZ9kezVFZRldg
o/726i4YAjjbzgVdXp6KFQ84pLF31i2AyVcSjuJygv6x+Ny3lMxp+QnJvZkTiRG/JDkVfvmn2Gf2
EHmEEf/uFkyDCKg/YL+s6ol6pup6PX9L03c5d7hQVwl6FnlxkCib4nR9MJq7EZ+DxfX9ZQnpj/DF
SYm8Kn/s1TSPALE604++SaArURMaC4/KXQ3k5rrEeqp3Pt/g99U0YMRFi/Zh94RP/B0+1U8jKdhW
cMp6wvNTnZAM6/FOHJwS+kZCUJjUIMt1BlwS9nIA5tuy7tJmdte51/xERsN4j9neqw1ziHTMcZTA
FaNLnwe0ztGlsW4JamhFO5D/WPbEDNqUfmt6NDF6f4soCWMVF2W9Cz2rKsMnGqsYBIFYno0hz/Px
6SRyM5DAF+ThE6K4xMFuwRilpCqzHCKc/Un5hTbImNYRxjMiqbH0hobQMxFV8wJSEAlPdfS7qCEW
gfMlYACZjyP71S3ncLXUQy8ZhapNTOanTEE+WcTNZ+nKg16Jf9QZrqiawG34B9eE0BrG1CsbVYsk
9n/ACFkbNncHeou+FSpKHP6BHCIGh6u74o0aI3JSXglgg9PSfOyn5d76WcNilkBzEafuLDqqQ7ZH
9D3TTAaNj6QxZD17DvyP38yrSa99Sy3ar4ktTU+unSFZkT+xCWdl2zEj1iRmBsxy0eJXH+kN8RAG
c158mwUKM1wy+VZ3DkAmNYH1cdfVLrV9zSLF5jHIzWBJKbusKGwev4rNQ8uWZd/xkP0A80T3gWgg
IEo3VM5C8MOds1kbZIISOCMVqtwA1jMhRMF9c7JUEWVuTvkYJDC0Y1ngoCrjFyStlpY9c9pLDQnC
trOlbmDCD/q+E+qh3idJmobvAFQ7OUj7N9S96zG7gJEua/9KPhPqjI/NOjOV8qrtd1EUOm1sICuv
IDcA3ot3dGh4AX/L47npDVOD+xEqByYtRx0l87P1bm9v6mlUVXANOctZOhQqItCfb4D+g1Bc1dHW
7g5EDODYq1tYbSKZEFRofMbV3b28Hdw2cqciUUyDXI9I8pGgUNimYOsv1wLdAA9ZqBllCYmiDQp7
oaC4nesJwl9ndidEO3bUK4x3ClTnYWTAFhUssPr8yCc/rR7YdeE1TpTqfp23TVk260Qfoe2JXr/z
kZSvliCjXlOZ54jxyz6mWwOPDLq8HFf7JDT4tuH7AQwPJUldSCkZ2qL5QpQYB3+HHpPuRvNC1IYN
gtXNp8jsKy/CebF/gYOu2dXT5EWE9CP9pMld9etManH5uqLgR0uWvHYKw+MIlGNUIAFIeBI+AwQQ
11B3tV+/5n2M+bBrmZ0tAL6HF8awvQxwzwQnPxXEVLMum/ejGnxwWjmDJZCCqMP/L096d15Qsh6O
dDCf0DITDAtvp5zzqiGaxCAL7stnb8b3euSjeKSXUaVfi7ssHiFZ7OFEHvNsA4vxB8xxcfaIM0FD
Fla913JAfoaWAhvnfqhVnHYuCh7/mIvZEOKkz20b52hACIAkw47Q8Qdq+gLKv/VlqAnyqfb04/CK
HZU8qOReqKTRcCS+W3/RRvBxqcoF8Nw/WPQ7OBu7F4cBVopwTmFsp9v4qR+1ENO/3kQHnlpFHd2g
JSx640Qg3ObScZUOXqY72yJNhPCxYUWAcsk+PIBFEvd4a3xGRHw0Q7V/COBMSwrOkJJqAhZoMnIJ
A46dlK1qF6SuS28HBLG3/BguYC16JgtQl2YHG8Iqn5k+oN+8h2Tiv/UMulapLGRoJzTtFdeFOJGV
4FpD574LF0XJ0GGxHWyR+TqXS1rGJuxuypHopgm9mfqyl1usitxAeoNmpiMG3LvCzm/zijUB/4XR
EOj/Bjw09ZeLxLLdLeQbHjbWWOuT5ici8CaDYSpMzAFwtEN7BMTarmcyfKP83WjMfzUC836BYGkm
Il8POAPOY2rgTh4T2y8Xo3oRpsxNyh+Cpwa8w9pdo5q9w1IfVXeI3AyzheqpSBdkc4C0DR0OwQKo
VNZCokevzyQ1JFwaMaG4c9v8R1tkcFJeceHhhBad36ZodPsnVj09gYo7eDjL7NctZXFIS8sSd85K
l7Xd7C7gfMyYqMAzpGtDGuImhrUzxJDgd+xUBJYdFrCGrwEX7d8pdA/BEX9B/zIWyMAjGFgFhi83
OSQIIzVmowcyZs2h0QlsIBF7gz8uFGy9eYl/3TZ2Qu6mxulhFeokAmU6IxfejauTtp+BKytJw1+v
pytpP9PpIRgzThNLNup3c7tBVI8A2U89q7HidgyefIgtGtXRpeBYDngrjxmL0mxLARX9sBmK+/qo
cKqwcBs4negH+nBlgu+60jpjzlAGUS3qis6vwPDqmRkVJD67UXggd0BKvYqf0Uxcan5STd8eXihX
Zvh1WUeG2TUVrZP/H/TZBBoqdAikxoYLt7t/YLJ2uhqJ15WltSnbeyFkkBjr8o6Vk2G2JmoeXpY3
O+aH2Ls63ap5Ff3zUX8j61/tYyBX+MFtyvkXY7lWs0n77Yd1ZBIQpKxJYyeDuCOG2gtoErN9EpU0
fufH+osI1tJi0iFWYBN7zKdeLsNWAhjtfTkwttvxjR4IRkyj5rXNuw9b7YHXsMILiQY9tU1y39Ql
OWWBcUJs/sp4czoNxF/f1Etnrf7rK+cmHfit+D0vX4Rus3EMv3+jbr+BC1VcBt+FZsPDmzmoOZul
hrmbKluMLkthDL7QzLnDZSY6kbZePBsU0xhnV44pYs98Qk6hChK+Bobz7jL8CLnAZ7iup+Gc+qZt
+LyABVBWltZzH3Qu533/bGYQctnZhCJUXhoMJftPf4b3f6Z4l9Mh3U4oCOiJob+c1sQ1hNK1NLDV
kjiYrvoM2H1HLMBJuDfUWOfNXxZ6EXnrVcs74p/ZZyOsMSq2iFrWOMszYRTEPMNau8qNB94YSKB4
aIfIJMtTm0VVVW8CmUWgl/DgT4MfTAArx9ucd59qtEs9AjhhsrF/HEbwhfcrmt2CF0XiLX6QUbvg
GcNCGMFufi0TPjbK9xj1TI/kM8b6lQFSkLG2quBSjTHX8zN0lDu3FXAU3qEguoQ7UpECEkr+JPh8
0c6XgGuNkphpIt8856NSc6Z0epLHAJ3PO509bh8Gvf9y7o9HGwv87beVfK4mFE9tDEo0hDhaUFRh
5tcadR1Zq9JTcHSy3a8r4Yz53kbMcWfYy0nmaajUpgd4Q9Q8xVmGzuynfWa/IVRZ9grYeNHYaE7x
S0KLxAtndqFyE+eGJV8+CBvwsTuA9RLSsr0ZQCNNLQrdGfQ/TmkqwQfkwL6wVuwEMqVuog47jhR3
KDoiu6xaxQXDhHvuIUXmEhv57nkUmLtqxPFgpmrAoEwHtRZR0WmSqPR0OYBZfuK3U/nJ+8KAcjG0
4OsPLWzAjM9uOiQusN90r8TzqvP8x5Jh/EUdcNhWeiNHW6XneFAfDk9dk/IVKJLSoP+itNbcR8HP
c/h5er3zBVvyHaURkPU/N+yX/aZJkjsfJyDrnh65lfxJmcpF48oVQq+7DD6dnqUoM/osggZVkdnw
kD6zcVex+T573Uln/MxXYoBGQUxWKIh6ore931l9k8H+eCY64g5ZIo1UpGDP0hlImhAbMua/5ict
QElfrF8CfDygoUOqkkSguNTNF8nSFpOinMJfBb0rT3hJ0J6fqtC8xwPAR3U6yZEC+9VCTDslEgA8
kcMBusLGOg3EfPD2y5PhcHOt4uTrIRRJULbVrmH3ev9+IGXRhngisIXxb42TV7EwoF6CPL4hElEo
nzBdUPcO+67A1wCTja1v9nT88SS1beBMLc0rzIpE2zFnRPjfWcj/HV4CLfjOWC6Ko0tqh/7jEnYn
Q3PIoeILs8XKfb0PuAwH/kLl+H3m/eKJ5CQjkFrJaqryprPZmpSMlcyF4pJxCBaoo7IoqcGWh+1z
y2IomOt8XO1rI5E0kgF1Jw4NZ/iCGwIr1bo3nHvlaVxwBr2/NPsoIrKe4d5X4x9jGVi/TEwGfXjH
FsiSAfpgDBbpCsqZZn8Wl9fysfvbzv/W014ZgtFgcbqFl5+vZxv30CHtGNKwmUaqa37QufMX9avF
udVlbYelGKY+vjRKP7gpzctLKA3awC+vYAgwRMFQJ+geuX+btAOMgyYIPm5NK5AFVI3QwqGaQ5kB
dzqVgIMWNPLCoRs7k4Ui4TtXp7AhsaK5CjGdla+zHlbsxk35j0rBR0mesNrCnCZrgmW0Uu96zj2g
kqAylQV8yXfFnSKMTkxh3mUugnQSQTF1b83VLZBP2pMyDmCd5l7Edur531IUeXTA3jktJP8vr0qp
pqfvbf0lXWrSQfA6J6fsy4rSLP7LnLoUh9CQRXtuuXMKo88JNpUFuQW++C/CQUCkKnZoOyN+MTp6
oKAj7FsKK7DicaHDZ5w2NiWC+WJTyu9nBa8aBBoOQW0NCvh1RuRDdYlHhX5VD2pl29v4DwyFYvmT
3Qv9gS6MiqOdqH6gHcNK4kft8r/x2cOGpxyBDd1te/1U8uu9L8EUUBxfadXQeUkycE2Q66Zeoawl
YBWAHdlGyC9s6pjqCSLGjyS35M9go+IZ5kuKaq9wX+NFP0gk65j2gisWXwImtm464q5TXCiX2ipq
4Zb0r2OtuoSfwStYfZQ4PZ5NUAHnPH9afs+SOd0QyB1bxvzvT5uRPRV0QOKMu3nIsmO23zGPsFO3
ZO8Q3nssh0jl+BHLCDGrsV+h4PAe5xVfkJnfwndxn0LEWr/Y6dXpClj0KxE+v5vhPsht/PSvdzHp
xhUtw69McFIt6IUqIlrZSyErvJBLikQb0DHfSHJPtzFw6r2PW7zbgbH+hUS0dvTSg06OSnVL1FUd
6Uz9xRWBbGAQB241ZuMcwgA0u9DxBl2yX85Ll+esgeS/esiu90dSakarJwaKAFTDMzZh1nWpZ4b4
W1/fp8/vkn03g9d70qgbcQkfom68GMEZOQWnBEURcJdR6IikVHJn/lsDtpmk4IG4nZyp8s/cNXSr
wjW1gSpfBA7DL9xFt/2EE4SsY22GoILOjwbOYjjDYX0Vz4LHA1NsTXu3l9whHdwyQst4REDPVSXm
h66H4L3rJHpGQU7VGZhoG6Vv2l98j0vMUSwR3UYU+gXb8u+MmKHOOLwW89EIBZbp0K72Skv1bWQj
FAre7sZU4DH2VtKxhcDYwa/zGzqRxBNXXcj3iI3KU6F3w0ZJzSfImucdobEh6dP0fyO7gaiDubRx
UYx2Kdpt1ir4QbjV3gwzAisPAIuYNr/HpaClzaG7pS5HoiWaBYC9w5pA7FE2hQAbzAn61/sJlkhz
7uiiQFCg4V1YgV+WpFk4+ng+TvUxp1CiAUth0wvLsHoNm4wIBuSEQ/gu/EeaaA8572GQh4mI0Zz8
QnYywfF7Fwq4TWET+kt2+qxSGtEZXVH0f5ev/O2gVJeMsLwPMdF0PSPQC3RiGbEX0WzCi09amtlE
LtNiXqWE6J/LFhQAJmMnRolHvPsa8fxte605a3SjSgnv5q/kQ9bn7B63ie91wp/+jdyN8zXUwp1P
VeQH09a0HyGXSEf76m1/xU5TXhclzpMkOQQU9prDZoOwwwUnG0H1jAcCztXpeJkxcW9QCo8wJ8BE
uSWl2BVpVhQRf4sU53bugQIq+IgWGhFk6wr3Ku8XTwwzsSOyT2EMXuTaZvGwlJUiiCO3NVdNPo9P
7RRQQxdV3PlSYPP/xO5fkasVul1AQYrJh1jFc+1vPuG1lAIlyq8QpfH1xROmI9kZDrFvBTy+rzab
ful9zcsti4t0fWoA883FRGmnO/OTtvDW3mTgtY7wnZLgTQ5g3MzKGR1lbuqActrnFDHA8eKXkijR
rwf2u3bEVOkE5V0azavjLCphTLR3uHj1zSBa7zN4w1mGr84Iu0t2cl5C2tLHSokZkHr0gYYQ6VCk
Zwafdn8L8JRKGTR3BuB6g+4InPvbOIW1x3PTdsS3o7LM8q7CO/8Z0xUz+D6yLNWxhU1tP+g6uVt4
1oj910EtOi+GGDtk72CgnNvj8AnJkxrmYYBrzxnrw3eHaFpcPToUECU0PEt0ypZTXVSngbXvfVAt
9Wlb3bnjWW2k04pX9vhejv+D1Za+UFQ131Xq9DZjbtbm6tlwEVcbQwLvpgCn3oAWHSEo0vAHNpTs
EBKFNXt5OghjaRhJDpdhB2soC7cU/pGmg/CSfg79AWkGS5NCPf/ikCmSra5u/y/Z82GiDBoEMhIv
mcZOpBjev0qawItVa+UdjCvBdp0efas9ZXiMpgJbcO4JNXkdZ/uVJSFODMT3fEngrI2wWpZVId6m
eJ/Z1qssROR9bxT/KFzaJDtLTy5DjdDEY9UeSPgwwC/XYEEyVnHlQTPM38wIJ9ju5J330YFLotHY
ZOE/ndWWEasG0pfM8l6K+R1YdN3HdLL/CfcDBFX6sq2p5UaBY30pB8OSJu59bwWeHB8R0WRN8fiq
9oJ9QUTJxUwC6W2dEBsfWCQxMcfDafjIezBa8n/k0ZbWjugTHOcIg4cnXhFHZEYv/3tiYctWiD1p
9nxz43NwjfD6w15haP53BQ1t7+h86p/6rHBw8RYqzPa3C42ZHyIXId0pVHeiQS56juF/NqyrEldx
bp0ufvjnLfvwx6a3p3ho3+3vl7qki9rhsmsaKejOVLjWljHtOkN7Zac0Wn/SOLGlPIPACt4aLLCE
SxryeOsRuG3y9Xp8SkIokPyeCz0JnBprlQaRk71accv34yQArZAv2qexjd3vkNCpEoQ/94aH0NBT
JaVUBL7wlv5tpZxsbs6GL2nar8+5DYgr0apBAT6vztmBPd7+eFwEhubuyYSOL3vCq83UYDlqFNWp
Z2HxDrD7CJhqHRKY44l6u0Qx4kIqciTlAoybcAbh2doVVX6RraB2AXPeCNEHfNoK4pk4PnUDMXVA
7ID+j3KWvRtXnjExl/hKUfTYz2/KKUHociX2RsRvsvxjwowOvDCSDgJSY9H/myAw3sDAgtWM+Ea4
2gDWgCWzwcLzI7izNg4X9NdeyS3FY4rVdFbLQ1l7ZqpRDN1wQsiUtGMmFr0wjPqOJL1cT3j9rmRS
Olqaz8EOZorL5fxC/ryuYWabZbKnnLAdHSI+AeasI2PLi7wYl7q8cKclQmPdezfIt1MRF2qzgTuI
cgeBkOtSCc2gN0acSy7JNbxs9koXg9BxyvVggrj8/zQE0B1liJlnkGLTfx/XCctltdJ3yjYW/xpp
SCOu6FC199Oyw1aixZV7nwIb+TCyoCBGMc6uax5s+adLDI+gEWYB4l9ZTy9FXXeYxI78iv/E4YaT
1Y1tKKpvHSp4+oYaA2vRlyTbOo00TWxe/887bCIgufdNCNKBtMwaarLQmbluzaMYWbl+/eqkhRFE
8BZIfg5R05JOxxgshD9spR/IMrpLlVBLteKmXIT5zaiK9Ta8++S2g+39snjWMseH7kEBgLKYq6Xt
0C8/V88jj30RdssfCMBG8kLs4q2KU67IJaAhxBKOHG+xY5ALM9ObNV777AkZ4Q7X5YRPrnLyWn2o
Q7SF7L2CEg4mVWPh5LunbEeJxG/pTSnlwnAZy510WPH0CNOAMSsVwlslGou5tztz4gPHbVAhxUlr
WHVNdd0gkNkDOKimM3E0vLsrf1QZHrUM943JcpfZARVddqM12fnVkexFvuNCquSqcRdiNaMxgvgF
SpaZwBfBdjHL9ey+HhZCA20KRr7gVMy3/gpmeXV5rfzDUYLG/3HFpf19hMu6KbSDskFW7DLnz2Uw
mt9pBpmEBgBxW0cy5x1pKRbGMT6PCvyotPtitVlv1qhnQkZLybuKHe5BLr3nM4AkuLyuG+Ohj/y+
grxQS8F3aBndyp9jH0eWXBmtxQRxCu6FT4HMzJWHg7spe+NihFHhFA7knU1c5JnyjzkoJ3C9ECDj
PFeoFA9kchfYxJhfaiftCxdqtPP8WhUOV4yzUR8PRFNyYlytSpUZcJoEyB/7jl059eOa98aSxD4A
YnpwWy/9e1IlE6qaer2cnxcOI7Kj+Y1T47qvDCoGCk0AnOJYemBYc20CWAYXJVcGwZ3HqYN1x8HL
hLNr5e7/3UIjg2O0fSgceNcblQMPT6Z0Z34U+UM34YtmB4R3AqRivrV4FNI+Q5IPW+RWVgS6JSL0
4OuaNkJyRKv/LPR0tbDzoHpv2uYfOyFn7BH3GNcuoOiiNKzfxMPNlMl5N1ZtwAwSmNxy8zmVZTcq
3xR/uzrdTcD3YYk9+s5RTYgcJbTUICmS3k/Sd8nz0cw3LNXfifHVIAyppht3DUUz0NqeWebWcW1N
qSYQvVA/TwXpe6N22jSOCF6cdqYL0+dy7NM8w0hzOdlUnqNImlxRdOy3qFDWUNthn2fXO9fygqGC
T5cB0GE6BgSEfrjyNT6w0vq8P0Lpjvn4AbboRvwHsYjnz+xXOc9OsBZIsWqyvRymnsrrhH2tYoTN
bK4VSA1Mocsq3fZTQDeHucQtf4JVpk+IkkkoQfFwyLatgCcHClsScTvxfEdTHpP8sHIigElfDdyM
HkbdK1arNLAT8A2jeOzpkb97KFtyq0IKos5vsSSd4Y1gRdiThmfBopeER5EncDQA6hA27StfiV4j
hJK3JKG5Zb5V07gxzq50/FXcqGfckUqe1hTpnVCPgEFMEknB5Kblzo5nmT5dN1u2srR7sd1c42Wc
0eCFlKeSa6f9/09axnwkYR0xbH/yLX6fGUgwARjzIz1ePyLiQoCUdNAbZy4HtVO7ht3odAkg3fdi
H67L7ZN3fIEJ7mksq4ItgtJGaMOjbd6t0wPseo9l7WcFizXvOwVJAbcW43OIqmMfrlfGcnvVUtOo
asYcIGM6BSvXbGh/HJcew2+oE8CiEbhsCdr34yg0Vy56XHkgfirZkIfVaH7LC4+PJNQt/fNtb5XY
vkWhBStuZ3mjcvATRtEadsYEOxNlbeIVkVyEbSlIE9gh6yH2nPpM3JCi60K30ZuSpgCHOAfiU6nr
/nZxjMZoGKgorVeGsKAuckvk+658MN+7OG3Q1VNwE/6qPlIhp5cKXWKW0Yvkq7tgkooU6h0gkMY8
nxXssHpMsqPfryC9uAh8V6sxmXCm/A8RJyI75lpw3PgL2xubyC0wXyhYPZVu0zsvikYfTFOD/5cu
XEjucCtBnKspO7QMYYWDdgzeGP8kd/5xXDbyz2pSrlFtt3H6IhsXmLmzQPBe7jJ4Ss4MQmnFd5P7
emVlNrz2H5BG51DVLK6R1Ailcy73Gc6xkgbs0vluqOkotPQs5S7EwwleXLSqgNbJAVkTH5WzsrD+
4Ktv/syFalEu8RE/DmzmBtOb0eK+GxC3bgGTrAYIfNfuqSDeJ/1fI39bKAJvWoAX36iqOfuRxU/7
Qp0xt3FEcBaO7ixLzdruwZatl1mX4U61h1cuPWMFdKIzorUG+KiICQ+/9oJ8pNGrx0ElAIBDtnvZ
7X1ktl5wzYjQm7h9r6chqyzjMgdXd+IZ7HkMm2RBh9gL9xnJs0KXJ2YZbAtE+9qLjowpoUZDBca/
wp03HJbL5eFGJCOQ1pe9cj8vC+Ep/Z+44LUy/iwbwqRrIoALUw3RjtHPiCun395TM9TlViLB1cYf
8Stn+NX/5lZrbJZjWbaqQ+Xmm0Llju/0XyCuGZwQMA0lxZ/gKnFZffwrVz5qKqxcfXvrGjNnMbvI
EOw2wk/WM8KD7XrJOVhcQX8mQnoEudp4OIMXh/xqhtyvIbG6WrM7n5ETfvgAdmDDKSYRR66+jtY6
RErV/PIDuKTBKRu7UgcrJu43Z7xBYgyIEkvMQxHpRIz9+Ask91Cw3qFbphbPeGco5olbNfn4X+s/
R2IgEFD1oVeNsCfUj+dzWBtZ9DegzMPJxVMFZ/jBbi56buXKklI6S7ABfzpNfZqCwMRvCU7K9D0E
mQ6GLpyjqqU6r7tI8zPwHtVuDeFbHVY848Iw07YHARtOujyGLmeuKMl9nmQZQFkP2DjRemGokfuT
g1QTKonbxUHtvgH6SL5Xbdm/e4kWJTaq2/f2BJiCQ9t3Q5o4wfkAepwkEPYFF2sJiRuMp/2LSfC2
55LedyZypyoYsyuQloD9XpDZndQ4/+lFLwofIgqCxWqJ+905ySIKM0zy1J3ADp/HTxpfrnRKyDAB
f7FC3tp7hPjONAcTlxuvEvwc5vi6Kj7i1wd4hSdet2K12qdZEb44nz5dqEj/j+6jBe6sljnVj8M9
YtZ7Ns4PWy3hXZRRVITFW3dcKIKQ2KBu5UZDjBtY6gJ0CTUSKp6gYRwuqYScKVJIUpjno14XzNnG
gjmwg1SWbu2I7fdm0COsB5ac2cRhSG3HMHE9/6Ot+3rhVxg35s69aYwC/bnuJ4HXFUbJ2g0D66rm
nXR/7nIeqAcRRwFa3aHah814ZQxKnlpSfI7ZPjJSqX7a6SyFTzCcpxAldtfWdIHGQwgRrCKim7g6
qICoa+fgXsx4VM5er+MkE9hkWH78To6jKgkOjkYSd3rKF7n6I72bBhH38t6X7WLZt2OpGYnfgseH
c3wDJ42NXKP1N9hWZJsCqsRBieS4Qr3JYboRXxNJ7sa3S29zY4ToJliFeo5JyP3g9LatzukeEp90
GX+mmCvWazFSCy42n2AMncBoGnOg0psjbK+FNkZ+RTNCPZbm/ZJox4B+NZ1dXtaIneFuFAuOTBpL
WidDMPpttpHyxpcibgjFDUIhkMAPYOoefIJYUe+wJGWVmtv7KNhymqC9+MXVx48/T2DjEu6FYJxv
p5p8svgh9MO76Jpyo12SScoBAMADe6SeODW5GYoZmtj+kZ4W0z1RCxsngP/Coqc99w2foxPM7STX
gBQ9m+ponVHa3kz4YKsw+fDktGeC3U46HqqoxmiXuptwalJuTKHVLyA2tXx/b5kIqVJLdd5iM+5W
TQXCoM6ytnYIEIJKT5Lw69L9E7YngYX9qiskmKpEoJZTMZ1muqQKV34t93XVDwxxfP8WlJOUHQDz
TbbsBT55JVglwAMm0sAg+uAbQFqm77S9aUPmjSElzb9+scePrgV3iUcR8neViwfl+A90Vo3NClB5
aLVxOX/+0JuKSyjMdgUSZ4FRssPwfYYGpNzHV2sEFyCYkOBOmx7RW6fhOxD52nSDYjhEBD1xt4OH
h7ahGqKhdFgaPklYSHmd/Bc/NgDjsghGsAgVd7Ab9u2QRj4xWUcPt+OEqTdxn7LytaTdv75fECu4
Ao0OUK04DwZpKJUswFPPbnB1GBEbiHKvtuH+0H7hAQngr64QW9wBFeXc+MMnoTXDuFaztfjdXowN
y+aZIYpCKn8pbcbS6YM+HCJyY7+FcoM9ePZAouLG281J8wFfJPV9DITqMem0YowfafflC4v8gUKY
mt8alwnO97KanjUIxsUsYh+Ezw1PN6YlnDAPgPpkHJ7BFFSzYfwJdYeh8Pp6Jucgo52RQwt6bNk7
iQCoZWWz5ACxAUvvrFo93sFmEaKCmp6BYg2H2mwsB6K6gpYbetkS/KFSCgLTePXIVA4/mYjKk92l
oegi3K54Ngnusj/RyajX/onlfMorrn041eFQ7cUFNfnSxjH+dOrJARR/4f3Ycu8pFjwclz2hrnik
G0z8vYaCvSK3pgkmw1tima71xIljbjVlFG7Y3Huo0ZRCs3OlW5LN/lRzUD/7Ic1NYG2tlTxFcCxS
Cyec8uLLymxS4CW+VxTiBWOqHjmsC2GFwdGJXa9n2tQUR45rj+Yvj43cXLM/iU0F7+pIgx21eNPj
EoHQd/60a0ZG3JsErmIwqasnKNSIcWDN5XwY+iQMHuBpCFw4s2ImxV27DjLfEoJ58uVbckX2tnv9
RVq6DPio8jdpLNxxplwuT/FFAvALIgCKmUn/nKQWt2x1fEW3W85UlJGG0shElkk2amAIXh9X/YP0
QlGSoaH1+AIwx5jOeIkxKKfVItpnj6Gvbx0RdfMOgHmXc68GWQCf/Yj7gBLcfBa2I0ivf4VgjnDH
zQBn+JZdHU28rv4qXPqRLzMxMVQvOZaRpTXk7SUmAQOiHw7tcvnQbwwRtkBWLc861q0mvA4O/5rF
gXq6b8HOgMElAEIY2upNSlZJSCgojpy4QoLNuXQbww4ugwy55Y1xS03SLq2nfDJB1umk2JZwn6Sq
XEWEs0UOkejlMx9AD3lshDCisLGWvcTLf/1KzoHQV34X6ZH4ODELcyno3EPVfQCn3XV3jaFZrsw7
7QrtqpWe3V/aY6RTkVzvDucJuvSCXWzHxawHvq0nRUamqkSTxzU22vwwJMIptUcdVerKZ0BOpo/Y
hclym4eXEQw0fp50AsFwxifIyiulTE44NaGQZqRv7ynDkL7SXGkSILK1l2psQZi9au/wzfByukYR
DHj7D9vGD5E0m+ZjqbDeM3fnfafS0+7fvPzu1Ra+DsVkOqNyU1GrhdjSvtTJjYwK+5IBToB48xgq
39SO4C/uBK/thiIMLeUpOQsYr3PQHlDjCtPRGfLtAAmAGMdgqHMwK6t7+OInVFz12clGYPacb9Of
4FPPiwK35PdLJ8C10t9hqD1OmNuInkff6mGNggQwGSXn4SPofNvf/jgm1ufLBKFNKpilYiJuZyWG
w/Ynd3cSObj+fqJQk39DqhpObaN+UI3/hYyT0JAQoRrbI3wNj0LjhhCsiqRvPmXu2RSbi/83zFJ0
iWcJooUHGqQiv3HqwQbtwxZd3Tjn2JdKf1g5kWGYk3Lp1K3WQbB1RLYwe7/x2lOIPp0FYvoXJxuG
QZIU+hWMPw2V1dH5Zpxrl9+aVHyzxPNcpiVDV2DrN95ePDxmg7ItRQIhXYjBeIlZr1Sj9p3nDnQB
yKqEVH6Mg6hlIW0SfiQFAhAjwaULBCvA38Zm5DHyG/bw+QfjOwMOG9dsomo4Ikioc7lmb9r8q/+Y
2eUlttjhxmL9Vgrt1ed0Ti+Kl0s3UivyAmBMo0k5Y1UygQx0/Qc7/t1ozJtqRnRQHUFVwXz3+NV6
GQoLHla96TopvwJKg/9liGY/4NGDvdEkGbhdIvpkH1cOHBBMKhKb1prprYVvaOOFNXcE9hxocV6N
daKc8BZsvjce6vM5b0CS1jD5kDwdHIo9vpsGfjQYvluW62pl8vIXO8u/TStLxNYnW44KQzw3ol9U
JZE/BYg7y6kaIGFDIEGz90kZxDbT0MKDGIVcZjzSPsTIEiJgpKoCLjkx5MaeRMIbNJO8vOW44UO7
F/TWussBv3QR29KxLyIkdaA9dOtS4W4Sab7EpwpbN+pqQ6BArH20O5EM4c01bEkDtekZp92ah4+f
iyBeB2ogCVlMnZqhWGeUAWRnI1QTU+uR3kYpIiKejszKsd20ymQC09sKMOoe3VX1BIjChh+oSBcX
gaMXfdLcId/mlmU72biwzRxlnDrbi1kDG/UqdgON3Vl0c3aBVfyWhKsYUpy7TJyIPIw0SrpTE8KY
4BhaSofvki1kILTNsb9X5+w7nrkKC7H/z5aE4KuQ4paMiGfwmDqKxQ5TOACNG779tWLGRm/afJ91
h95UuIFFL4pgBjNYK0NgQeDwxoMHXozYI+q9YDFShZ8u/X/mZCcExeMZK6dZjoV87fKo0Dwcjzl6
c4IB2wQdRYmo/dPPAt653AV7TCjeXVXi1yPmxjoLZFBDrUjexOhVrylYqy9ywkShWX8snySlvV1P
JPIzOfEdiBN9s05/60DgFBCioZ9Vs4q7YI5mxROjN0QLUZ3j06Rtlc8nEhTwf3HRuAmxgWdR30UZ
7S4OYHEms1BeDwTrU12wmrZoMX9m0q2jODyHlZICfFMYijXaZTGIbYhMf1Zih/Yudeg30GCPEAU+
1Jg2H3T6Y8muYtoluNok5uCgaRZ+UoHSRVgcXjHdnhBefjNzionm372HBofTwg+4toHyJBurnH6G
l1MW9OMiD5z8k8lPAWavKs6UrJqSc8lVaK+4jgii9G6zDSQsVzeSpEDdn5nT6yzKMABm1xcAYVmG
3PnHz+PMHehUD33U8b/qO3KMtrC3rfeIUuVTv1MextNK5dUIJwj3NY0+g3EL8pgtMUvm1akqdQ3I
u1GCidZeG7R//9mRwTlcGLanjKYyoGfqBHuqbWi8tyfXAPYEMeiECyTHUeMzap2Ni5L8z5nLlBQ+
JhaqEDF53OXT1zpXSdfVzeWlfG6VyxK5DSbW7u1xJ/EoWw9VVhUxyyXo+aUgMi101RRT+TLCWI2V
aqA27XMKAGyHFZG3VwfszQ/tHPtCONWA9y8R1Uhf4o/ayqdDJo9yMynvhClY+PstWpJOhRRfcylI
UQQfBcOW9UyG0XCeCGFDeXO1bVF/rHRh8kmfSISOfCwEUeGZlz4vqBeQJJXXQWkOnhkRljUeApuV
LX+EyUMO1NlxIZmj4XReujbqDjKeQmQpv046HfJCjmmbdv6SayHbKcM9PzfAfx3CxUAcC1s2dcBf
ec7zEVVlWhYf3g29L6Iov51I+MG/mHqVngvhqiqPKb3BzuErLKlbsuxLpYlkodWcmSN52rAWzQSO
tjLy6drFIDkI79xAf6xy4QgIiW9laEIfAX96o5gew73cUR023+h3lyGb+fUdFmUDzegzAWEYJkPY
J924jTtUidRwg4WRhQDNKkg9QgyLz49vHI0rtltfzy8dbCYt0+0ZECO1xcmfujVAS/OIlwF9lBXw
WIaMya1T9lFJPwsTPlAaJjrcvf5VJS8ShLlifn8kmupW5RItH+5Mj2PNHzAHLGN9KHHaVr1kXeGA
mGB8FvBbMyepWdlsd3E8hmrhsJ28rupzurohVsdUNCEJzaXhdRhh784HRr9fybu5UNdM+ImotPZq
0VK9b86KyTfzOmzxJfR2C2mrHH52vdsdMddIiBB3zjuoaxqOeN9F7Psde8ZKXGG9JyQYjZUnOuwe
EXqz6Zd/HYCU47GHehdO+SrZGVIA9HyFEMFrWbocGkeI7k2Qot4hpDacjp/ypy1yMOpH6R86Ts+2
Vo/4sATFAI/ZNJ2enbN/4kQlglsrFWeNxg3OP1PYqfy29feNpLNI3MwFzjaqPVUt9339oOEu8GhN
5OnKg5Am1Is6atn4PYoRx7EdpY2g3UPHuj7gBl6OExktfM2dSAuzTtfH9Z6Pz9ZjjFEi4S70k/kB
GFBKedtCcOTib0FowI6wlGr6vpfBaQqt+nCiAPgWbrVFGe+oYViBZXJhnZ/4v/9cchGnaXNLyi3F
WiOk0kXoqv9Pa2nrzY1KJbQM/hbDycQCkm16/kI+gmmQaJVO3VFOOOHVnF/DRxKUDl5MsQ+YrtA6
eWfb/xs+5nqwVZhknbjmAbjW9gLa7f2TM4UEnsvMcDgFcvRRFGU79RVVdtG2DR4wpJzfPojdpBrx
8d9fElgmnfJEDUaVPQ2sTb4AsluGpa449/l//TdFx9E3po4OORbXt9EfZs+Qkd2db3FqAXd69M74
Gi8WVp47pwEKK8gz/jkySPC248jzhkauHi1QbLuUh+HZ9J/TAYncVIqgj8V2SYn2RxEIjCqotnZF
JSQzPXnNVO6/Zxjof6/ZyApNdWucLdQLjuS/R/pKs4YabASRmAhi5YYlRHD1CEGRpJP3k5yUVvNe
9WR9LW6jl1JzxizWKaw46NIZdF+MbgH35geHiaYuFMpdInvWbKpCxBAkErN08jkrlmBPJGV8iqMk
jn4XxGnFHtdg4l3nhlSt/SN6C6jaVc3y6sp/WU6gVZfIG6fiKCxfKI1WBkdfSH9iVcspT2G7VO+F
0aPvfTNAUZkVKiFfaPZaneUULffFy/rQZ6QdF8tF/5rHorN/zuNEZYeegNEzvXXj6GexA9VTUDNe
OyDUPpj31nWExQrCHyjb8dTVsSlJUFvjaJxrGy9d0s9sMcPCZvkMsb2P6tXy73lvwsBNC4CIOQJj
DxUDSdPcLfnhj+X29WduaAffYHnMi9zcoxhwlG75juiQoK5XsK8P1Qy4HznhsT/C+9mN5hVNI9Ok
HiSlZ8cnR4n1KAetwP+eHoeLzXC/rQsPHEPMoBoGpX6PZx5Gfsnz+UyT2+lWsbm/fWFTTuybFUvn
15ArmgPdOznf3cW6aF1Q/6zqQzRoEON2yZT/rxOed2BmOQzHKN9RLHwlGU/VlXsfWluQ88YeMQlw
VDXoH28t/50iqn5xwSOqblNQZV/P2EdCYIQFO5BEF8Jv934R2/fHO8S35dJNMV1kkk2gpQHP0oO6
PNJ9OUl3pmA9+CbLRMTisz/xA/ewGCqdvNRo4aYIiAwdYxrBoJzSV/MMuqSZXNZvY5ibbdd8rld4
/xdZX0OWWQLom9VKiD2xziRA1lA8+K51aD50e1ul7zzOb05gd3faqeajSKztoLsrd9khUSbymfYF
URUNn7Y5+JcEVY/gLE0SMMAKGoWvIlDBVs1IxuNfsNexUx9OLJ936i6M/MUx064hhLI9n6faEIEa
zlfzrUhIdjJF27d6fR24jv9F0/hJE8WMwp5Pbg58ztBwac1IbsLeACFgUxGN2oraJgqh8ph2/OQH
ZXnK8C7uqDLz5b9l9I0rB6uBIM0m2uk8YxW4iYgvSHxN1xwMgsQaXvDZJeQfVWEzLfOMiG/0lGfh
hZfpm7k/OQunbX/Ni7g40/CJFe2txshv4NVYzp7r074bc/O5+pIfZvqEb4fn3+ZKSxtMN6xsLtgC
IZQAhNtSnkxiYEEbNaPwSNzs4/zioGW2czyWeXJq4bC/8aGhDKyBtA6tVGZYPEgEC7zrP+q0Z9Tv
9S7m0CWAPVnOF4xX7/lSWB+09mNE2xV7tKtUCtLJx55Zte1UDQ3jkSuPbv9Cj8sjv424bXPop+bl
HafL+u4jvNq7S/4DsZdaS5Xe74Z3abYJnKkFIfbR4nclYLnuw3sJNIwsh2FjqesV93fS1CpP+Dhk
h0x1lKPyQ56KHaAYvZJ8N31iw541EH5G5blEoj1YePyJyhkZHRW+asS2Pd8CANUw85RILntWwT2A
1EHR6lP/Y67ssw41U0RtNSVtjwR46RYcEc9YG9lvCNAJ4KkLjvbXfLyIqhcK/Kp4pUG2sQJTMAfB
s5RIRAixxleV6vn8gjcQPivTo6VJCAs7b6FbJCqP10A+9Pq9YyXFvIoIIc9TdhDYLUTciyJJ1SLp
2pxxmpIHLNHDTeZLijhR/ofydEcjawtWHHv7ytVhBSsEgwNciVnxKwhni3Tdr3UqsgFdMsXX0BIy
VnRH6C1ncNmjG8+2T8wouhxwZJQ2Gm570v/mimrsnV3Pl24cVR/rbEPDej7oJsr3C7g4Vye69eba
/wfdkeh1rjnHJAC4Fq34/YZP3FkTE/5U8FoEi4gCU85A4rfSriDefsNAL7+GJPTQ84f01VjEm849
DwVcL8yH1aghr7SZHKeZSCrKn0A+7sNMdV1qiLSLSfYXhqUWQTLksA9mFKDI+fkSrK/9o2WNWgFN
1b9V9SenwZ42xAQNRM98NUMNsw1+G0D3nDRZT5FNGtS6MlLPE1NZaGViHXGMBkqqWag8RSEDC+gO
aFbKih9VBaF+06gl/WldQr+EM/RyL5DjhkAk53p4CBtrxmwiIEx6+V4A2rIiGeNceodOfBemxOa4
VfJ0mREYPzhYVidvcnRFLYV/ssiBDLfZokRREM2R9MNd+DLB5c38vjQIJTAN6sm8V9HH4jm0TPz6
z3tGqfNKWdDeOxpA2Do+uaUpLIXwo+BCN9cUb77dQz1piHmKJ3w1hBIoSUju861rg/repv7EGPPH
m2MAtJbZ30H4q9AY88DTBcXilrgohwX0J36g0eiMywacJda+NRt2N28yPsZpo/zzFESYVx6vggB2
vY42F04PGJ0RE8yX/oJIhylEjNW4+v0EBs6l7SM5gZQ+dW3QFy6oU0hgkLgjI5bPUxFWcb56GMeJ
js2tclR22Bekl6falLRhQmnti6HttAFOyPxWQcq9XL66hWc2AVePm0h1u+6oW4+72MsRyDQvFoAS
OwAqUQsYOScS/abAtFPD2DoTov2Ai2WGbWeAEhg4YCIDbMJtOqPad3mJjdaxKZlajjZ0ZJB0gVwx
RH/dSyju860FMY8a2ztQHinlHKyh1LXCIb3P1NEYAgKCyFHOAx+OD2oAYKxCCTNJnz9sfvx3rOYu
DWX3zTG1pXXAhyRvC88IFGNrwzLAdrGyvCm6QJgw3fGTyJJSdBeYDHFyFZR55FFfM/Zsgjuot0Gx
IFbPusmfpey+udF29I2O1RUX4PXo3zk7IBZQc30z9Ub3mnRxLzynALWqHaYdpKuk3TXpJacX3yOu
FBYMDvY/myH3wpeNFSRSGYnxsBn0/62YYm+8FCkdo8i4aF366Wr+2NgfueeXQ+sKkv1/uCO6ggAm
zp+8DaoT08K1LfcbDlvhTi3g9+CkCuK0SfWNVVYxAdjvaMVSdy7id0ekhTvKWDzBTTg1Ef9nfq83
xM+VJgy4VbHsZM96Ba6oKSwmtRFwOrczc1nn+waLpbY5RUYjuc/cC1Qj/CM6V1bUXmDPmKFoIdMd
1dIxIbTciYGVOlT/bsVDbaRwB15MoqxF69S6mNbseq1mV+BrN769EOLiioJSmPKp3Njd2EZKoV6S
S2qb44MnsDV+NuezNNirn7TvkemRowo0Bs4lYCiGS7f+sJTOafbqNj1VmQ98MlMFVk4+q6HrPnlc
y1R0uPt4I7lEDyXRB8X/1r18iFRjoZ+RTOy8N53xefFcaUiI3dzchXzcf2AmWnkLzbB8oToo86UX
52OwqJ4YzpCswelkIqRCGot5rUsQ0fUGExKeuOt96DKeJ3ufuw/Dy/HzJkFyNwJV6jucGAODneuB
VPoSr8dOCicZFpk9CFbTr3+4/yUGmb0v0QU5nSuX4W9XYQ98Kfzk8ya505HUlhbNcOd8mGdzVsXO
qi/ZjmbHkcab/sBk3J1ZL4uTFyJ0c0nzrJQ54aP5SlB+HaC3HRcOm3iWC1Or5ZBMsO/dtPq3Umsp
f1xnDLzmgUC9Z6QPXCIde3hmEQPAuXgoQWyudQdeWFJVvk1EXrZhVm+/yxm2Q8nP2dnXdWfdvWjz
t3595WXl1XX5BM0vE0GHmMG1yeJci3nGsqAqZDjLvIayVqDk6r4vavg9accPB5xFsy8VqVNm+H2L
O7aFgYuY8A9j/TzYRo5rI18uBSVvRjNZ6aYME8abXfCNURVsueKTHAsh1eUd1ydvB2tkTjw0B64N
us/zkJ5UhoXjSxo5iUYbnK1/5xpo2z4iL1V98a+cujx7AQd5P2mg+HtKoKhesQjptF6FjrGzyDL2
X8gzGb7Cgz6hHDgO+hz2p5KLx1QSpjGCzWY6rOyhKkEymo8nlABO3FWnHdl99Ve6l6PLn77mW4kl
47zbgz8If41UGR4LOf8tlDqZ/WfUhZq6kKVtfhVwrtiVHhBKa4zRsDDs1cLUUO/zKL0mWLWlW2jT
xzS8LAO3XJ3XLzXr7Jcj5ssUepvv3LgIYfttXfec7xZHETu5eew16PZwmSwynO4HVl9ksIt9e0la
z4x3+R+LaUWSZk5zMuiamgcRtTbgwI7afzCx+S6VABB5KHd7JQO+haC1t0UCcK5Zgh+uU4NDF3jk
MoTb5povQ6YkbMjn6EgTu7y4rWIbYRFd/Q3kg0fCGRgD7cUrHvDe+c8Duti8sNC97o58GHmtb3Y/
NmtFy+DI0fG/LU44JMw+gGWe6UPgtTDVD7JOZ55Y4taGscNB+EQJeXa4SuKckjCZCBNoGTUYBllb
DA3j6PywIZD5+Lhv/Nh96R6Y8xTfZt++yuy82pge1sH7wyu/i/J//5p4Rv/Zcjf4gBXqoVkJX10Y
kI2ZGuYp2eP9m0QJ1AQGOeQgjQZ9IaVvhnZams95Vd4H/4UsqfuS5y77nJMNs4nzr5HIXZ9q8S6G
RROtafQ8fa4dT9Cwj4a9f+zVt61atMfUrllJA7erkZgC1MfNOkI7XlA73htxOmOOf32gju2BlvXM
1io9shDgrDtIcny2IWD5dVbZPsFdWN2/trQx9PWWWZ4FlnICm/DrpmSwuolqvspLAG+ukc92gGgC
qwdwR1Uui/wmjkWK4Ow8w0rVGk8TxGEJyTTH4wqtdo5LEO5KdObLPZ8AhP/jmq2uA2YF52LGqRXT
jqKIGbrhm3bc3zKj8zZph9QloL7FqjCUmwwkjTFyZpMlyrzvbNi3Yf9GUVSzgm4JV30pVXtzDztn
ZP+skE15nQHGpRk7t8zR3LhWSpMeq6M0LxZjOPeNzKtxU5ay3J3oWsKAq+UK0TanBozBP1m5/iP9
/gj6EBXQFhMYALHuJl/Xg69TlCLnL98R5BRfs68pz4rXveo9468sqFTEtc9cReYF/WFaD5tJsI0G
ic0FVOqewG1pvNvVDlUR6gIcFn6M1hAkhlzpJCGouwqNV3sghaydcaHm2r6T35GiCqtlcIpzSbQp
AcgzOLh1xLr9V/i/ctN19NVSr7nNWb2U33DnVduBEko7QG/MoStQcC/sIuSbCdyoeAnjmCGcYDLK
76FS9ZJ2odgfNcnacxBHJeSNxXLjgKHZDj4MiDlHkmyweXy4KYSLLtYOp1gJxFcsTvuRV3xFQyrx
E69eCzF0gK2PDN/nHGl/zOXA6o/ikvAomQspej15kqKXcbpgfuxPUFo0p/k/ekhnkuG5/4GDvCyg
7fSYj2iSe4yEwP5t8+XhG95KUIfhUfc8PFNwnN2DYkkMPdBMFQmQwKkLY/GiBf+le8jq46tf6N2+
jWMkVT0mjLxsxFQQdA7gFQFEpLIz2FyLQr0iYY25Y+sBtt75Tcz+gRFMADs+SRnpBeacuBzUVK8T
cVxL76ODaviQAlkEHB9tKjoZc45HFnsd8Lupru6PoZXmZ37cl5Ks8WEu7opuLu7M2JaNGcFCOlD6
6pSsKC9z8UtXNkrFsTGzYXeQwTRjyeGjaAIdhePdiKbIVnTZ2azw7L0OL4lZp5IY0vBb6aKUm4Aw
usMXBOcXkqVTvX7b11hj3uPcHJ6/+zdVWSyd9C+cnUNBAYl09j/MJ8zWHR+QU3hm+BkuK2xmuDHK
K1Cx4v/hncCa0pnLPHlgOBJTwP2SxQGhKXmZ3BY1jpelK32/8RKo4mYcrjrdLVaR9CPgRFDyjuPa
8KtfjBAx9g5wAwYE04OdIj6GxVVw6SrLXZiqsc8qxY46zyPmGWV9ilGVSx2qsbWUeesf+AJB6GnQ
qVOGqvqepXBP5NQCIrWG6gw9bBksAnqRiIftjGf4llHC6vaFZzUHIAocYbnLjQHN1D5/Kb+nanQH
7pa7PofLNg24tVZjgxyxSvjvGMFH8JU/ZW/3eGx0MpwryQKhjiEgL/SohXnqzbEEMBawcsdQ9wBo
yfkQD+byY/Qf4HKGkI9jpXDKYTOQR6LfdxcuMomJDbhxSpSpQzJlVSXoS9MmDXHanUUDEuWDI5Zn
cF9NCzo53P+ev6Zv9aGd+vHf9iq++WQyxIpGwr+YE18I4WY1f7A7KBbwf5UF/ILIgWmENg6b88XR
CgsXhtWTtv9JachOm1yKcjQ1TbI/rpr3sPE8mRpJFgEHdsq3+E197SqA8lDDp53a3C2m0Se7rOrN
mFCu/RKnG9JommI3va50cGlKwsh9cLSL73pdia70nQA2SeiMwtNbwyvaR5aTTdLEk31aL2llm//F
Y00L7AMiL6kvUB7r/4U2GsWwjvs28fxnauY/kjJ5LZgOBEXI2MpYecfhWB6DsKs4gdy2s0kJl0wc
eQWJaM25XkYo7s9q/ge6p+JSCwEK1RB/ZIfJqEESI0bSYhi5lX+/t7VgvKrwo5U1+sqRbpw6Gply
JdL6/6F3DeB0KT7FVm8FpaiRmzONPvEv5nIMm198iObR9FxteUFRy4JaaC4CH5Q10Pcycy6yCq5F
h5+ege5fqNsW8rxNZ6NhkWLKRymw/brngnbbtpxf7kAEhyyz8d7bZuQYmuPbfICv2QqiEMYzGuj6
Iu/5dWZUFS+plMp7WSSzdsd3kFl1oLpSX3Mt2ZupecMTXJzU7SWRb3vie2LTL36Yv0+qMpE4lTSE
CYaIgCsGNPkhlMag+zKXIl2fjpXs4Ng88aYe09QTgRHzjToNKrZPomuPpVBWmrptz/xnINlFuLoS
CzcgwE6JSwiKuW1gDyrajBXrzP5oycBtsHCv7hq3NtaQw7AofHv41tqToOTfxchXiqYs40SgSkDS
3qEC7ZVC/xVugMkbiIChKgkhdD/e4nipvr+nvzaWyVcpCwpnwha/vs8JdO4k/fRUCBO5s6qcnrEz
vFT/ZlBoh3VFtsbU33zinQgaUMLNX8LNNYfv6M0irjVyVwgPyQaR8tjrc+2dV8nNWg1SNeHaOcq3
09hs3BwD5Vm90206v66YgqvRZkG9UGjSoyDD996Qj+MC8MAdfqVG0UzCTUuLPjSjhfyapJtke6QG
6M5x1s7H5/TEaqQ7V/wAvtyFyj0OoF1EjPv6wbXgHz+owlAvJxaj7FLBH/TkW9GlmO0SlbDuy1bH
T3PnhcDMxbhwZpbQZGtPa9thtX3vhYzBqIBQgyV24tMGMuLxzKh9VptyZMvBXmej4QjTSnePiy/9
muvf6Kzqith3hdG15fVqD4XJDQcmxq7OTOW/oi+Lfu04sZGi7nrj954119uiIBkZvn0M4ITJkI4i
I47takDOaPPHVwFGm+CHp7lr8KbcqV6BtDR7qmqVNGX/mH0GCa4PcVjKCBHzIbmAmcoDpnB2rFU0
++61f6jL/NKL7b21bkJPczOnIVt5ueIiKOFFGugPeEYt+JW/FJ46Lo50HCuCIsXWC3ehQZByq6L8
/Fod+gHRLmgZPooF2W+gA28VwF+3rxoF8k6P5PuAbx/vaGrUHNWhcSIv7PAfdE0spNbbn+qnm82X
E9HS8sMbx81gwR+iBdka4+HLeK2qoNU840fuRHwA2Ryj8S2UH1mdQayj3JRFV1s2oY9FaSd8x1Bh
i4lp9vLJ8rkAPg18ldMrJlpUayyCO8exhR+J2suJX/kwrvE2ubhZHbNBvXbOyPDJ0rISxON8xCF3
UhjzQTW2Y2PLSbDTEYQjWqMKjQF02L27vuK2ir9OA8DHoZ2T0l7xoafKH5n66sNxrBzQeDxlaAZ4
gpysof8itj9FoAg/1B9HkkK6/Crw/cC+v/gpxf1QEJGZztJlnO/Qnz8pORLE7RYOLxRSbWxsOL4j
EpjBw9MBAjtdbCkWp44gaxkduPPrLt+xTVC++LX+SwgKP1lNrNnW7h7Fae5qsmuHxV2sfg4rq/9p
Q20NuEfIlSj1B2BbnhmRROgOdbF81Yz0WLTqag+/vgm4gelAppBYkwckV3S5uhk9MtreCL4xgUTm
CaFxEXLhUvSwMNgVD6uKNv8s+PsnomatrsC0pa/IKzrptbvabYSxMHSDP7sDZN602aH+nv90Aw3P
i7hF6/5eY8HZbvlAHl+MRiJHQpoutmOQQR7pMn3jztb3xq6SzY1MWoinkS2nyQWH7q34T5b0waxP
C9v4f+CWirvRwrD3lf5g/tCc68Vz+n/g18qylWvURdw0PigdCd9BwTw8KVba1zcbLzunGY4vkiaz
N0h8YxPiZzZqv6Xbtu5rpO4U5uWNLsJK5Q/R/3g8FX2k+HxmGLwiG3wEXsWoyX+Ln79iNQo4VoAd
Al6LJuijWvb+rLJJ3WlMuY2w3dlrhp7LdEUgFPYrNAbiCC3/ZOeVGsGJsbHaX0CgCgcm82Ku4mc6
vL7MMLdi/jk6m4IG6oSExXTqXkL72+E5KD6eFtNdRJu5/cl8+guenMZ198EUfDgx+1Fa+En8+zIW
jl9BRTIe2xb9A3uVNeP6aWtd8v5rA20TbcfMVCxdLzExvoeibFgmHV4v56efrLo5kAMt8Ai0GlDB
A/Ip7X7+dSGSToDAGsPIicWYtIsHUF7GQ7o2mVYqxB0xTL4NyBa2HdE9iPWz1qp7fZVBKG/HI4xX
Ul7QiwDUxHAKVk9Cewj6XONdbo/XWJThAALNbXoH6XtadULUsH7yNttNREF40Y6VcRDA/M53ppEn
foGF6H96e3EVOZaQcNKTv6maYKzU3sKSJNHgqjp9TuRLtYvg66WUPu/f6K6q50vh11Lof+fVWj5Z
SoK3ijNSkcT/9yOL+QPN56vtZiLTnJD7kOjJ0mcPnvTAEKspwKAczz+/DWfKXhaXHSQYbWjaAbuC
GHCJ7iRZbysBt5WYZM7o10lnuWgQ9QUUKCUzNKhj4LnlwLWDTV3wSuxLTnP6Vv1/ePoLHJtNULCI
VmOgyocZDzCeAuZQb9pqyi+877OcoLRiP9qgM48qFSNt/TiTm3uTa0cx0Utk75qrSxCCN0ijcPfC
DYk56OE4ndwU60lq5k4Tsv48NeMgjO7DTO/H9XWE77yQtBGIH+/L0YCbhxI1kNqYtsyJna+Cfw/c
ja7tq15k60nunCjyS9BT5Tcbc8ZTKvN4dVe0PNABvSkqKyVrRH6Zva5qrdknPH315fWyB1OVqngq
9GdRdNEwOggQbL1KfKC6swdnTZPZyH0P5yEp+ah4GWADXJEDOl1I8PQX5eBt+ha38eTBMISnHGnj
vxTHbHXW61B1WtQPXbILJ1f3scwI0awDS38ZHbsuwaBiqz1eWvWyW6zRtquH7vWAIC16kGXaViJi
xdM2AhKm0eFoq7FXjHdNBF2/jXeCPQgevrRjGh6OY0asiweqPZjYIQRMKX6ciKM2jHLgQXOJb5gK
D8b79NWIVTstsB7+xDYKNpR9pQSVXD73V5fcg1VuXBmi6TySODeBuK1tM9+93W2gqlRHIyrun7n+
O0vGS5Uj32dNOTEXkOOBMaIudQ7k7czuE8ZIOXv6O+8aKVxidUo/O1g5wfkzX0JVXuHNtK6nB1ne
zxqWbwmHGz8i0yoVWWtKlyUf1AfFs6/k1+D5n+XbzuNHc95u2Za2xknEwq6b6253QfIhGS5uSjqZ
r8EqVaf2PmltQN8MJeduhHMRt1sdJ3vHP0srWKy2By6hiIpi4uNfOyamcGTwb2vuIHWghEp5u9Is
pooV2A2XMy8nkqKBquNiZbgobrgWWw1mlP3StRV0Qh23O4zLhUDiXdfijrVAOs5HtxbGfRdgloEx
oL3nzBww8BsZTul7EH4i8jp2kExm/Uj9fCTezwdi+7QlPsxi0Ifd7UBNI3FmIGlrLOf4Oz3szsjz
kcEhXERpbsTk0af6pfcoLCWt08gb39MkAf0l2Th4plW199Cb7qMi6eFx9NdqXPAVSFUbwyVoGb+s
8ko4IoWA8hkIXmfKD0AEQcxBbAd4EhR5U1DdDYTH+LGYc2IE5aBDr7VXmHkEgykFCR3BIHAhLG5Q
cghNEARUIbVqIqfoeEFxZuWISrkhsWThok19OEVwyWG6llrKc1mX7HiJE7s3xKwFqVxxH7Xbilv9
jhmB875P/wgzgpVOo6aBbc1mnFm13C9g3bZpytIUjxgseaTWh6ZJKTk1KGuGgrCOTmFceC2UmssN
Wi4F+DcM9sBj7hkNAo2OSOnF1oSzeHlu0QCs5lY/Gd1eVO+ydxYPTSX1tFvafBndhgQkCeScWOdT
Uv5Ot0wqPA3FqX1ms+IWjKI3iNjTSyoedegufQtts978ie2OYVrRuoCeLMfAVX/13lv03tzgxlS0
13hyvfnxEuAuisEUJuA7tKeYzDRZxn8+ghAVnTNmdUHTqXSemxxnfuZQTZMQLY4CQr/YARR9MSw2
bEUr0FquZGGpq5l+wNY7WDFc0M0dqOV4XlqsfdRQBmAL87a48aI5qnO6VbkQYIv29vuJg+/PFrKW
zDaqH/5HHJ7jiwtx83y1FAANG2wR6Y1FKeDhvAwGHWtVDc06obOa71coLrbYAX/2rp5U5P2nCUTH
pz2sCveA+eRHUIDfQs361OAJiJP+gFRI+AvKQLoCg8QB3AKPPfb6yFJr3qhMR6NFQ63pOtKGJa6S
c/oA7FvWe6jL+98pGwxXTOn+05aXpVOfXi6O5z/4pdFF/uPKBsZ1PFbhG+8FMhxFUI4IWPBEsLpL
ZJdywRV9I1hamkcWzsKTnHXyWbziHNVtjuy/bx5WisxQArDU2P4AV55vFyscwOzLXFoVA9U6hd9y
QIf0ajM/3ioU5m23YeI3E/zTO2nNRHhwH8YteZuynsgqfoNsCU/nczHeP6TN04LeHIqxqD8thMuf
VIX5jfKqdTdce+Ton3l4se5xVSOQ5k9XxdUKMz3JhEeA70fLJPY+8HQ4DXZdmqN9qimEbeHp0KBh
22Gqj5BYHWV487gq1W1gsSf0NgPNBEbRfo4NwiZgsU2uz3OK3n/5Qrqd6bhx3yaHFzpIQNRIoxhf
fC6wcoqekmg92Si0LNJGZbhz4aATvSUtv2Hun37VkVWgeI6R4zE7cA5X4eeBr8YStKIZE3CgjeD5
Il/twCcATh41XrpZDiw5f5t4l4//hentpAlUxRd5V2gvVuDcs2Wnwf3E/XzlY2PEeyjDhCDoWmaT
bTkb/d6QlWosgbCghgPb1V7nvOTH+kCeoaChptjYYRQJjJKvgiw6jIP48tQDJ23b9IOuSmZHpaDR
Bms6iIF8zktPLVqAFR3uYEjOpjP1jq0qGPKngV9AwA8nYGW89Vulia8BvH5wAT+cL4wVHzgyrqCP
cxAaGbuuq6BUPux8f7B4esAYBjgUJWPlVGRqU9EJtWogYeb/3O9/fxYJXg8yRbVqOp9EgwRrpfQi
tXDdKP/YMvj37UxB3fhZQ/4+Q1ZwbDJyPwFkfHWZIBW3T+GYronHlRyw1We0+pb9c5K9jJ+NbazE
DO+z96vXb+W+9iUuApOoMnJloct53lZLGQIpANwY47PRpkNeRXO+cGdzCboQvjteuAVE7lkO/e/e
IOUHKRYM86wZZP3wjCsRDkgUpcuYARJrCOB501HNyFldiCRRAgDnzMBcLNcUAXoIlerDsTM7YOHD
rgcWRMdCfnOsu9iBp0XnOmaEQRmEWSB6f9M6ng8X7UWNIfEcfAD1qeBpwAuwGzkcMiopNS12LRIB
EQ4637C+VzGeqbDtMEKb3XGosgOCT9wiMnKwb2kurkOEBrq1jBdq1zLLhxb8/sQbB5/BSY8pYReG
5VfbRv3H8j1VUVzqvU7Ioarn+w0prXlX4M8pfcYDcyaNyMozR2J3muavqNiMi1grLTV9eh5lxu0n
UBY3GKDxkcWUNxdheuQnzKx1VlhDJ93Jxq1lbhKr2zc0FE7PlCGQwOhfB66qTjDSWNriJ8nVkO1w
mDaORVgHSLPgeTePstm3o4hxwmUB+po8XawSIZQnr+Iyria4j2mkoAlKAmgMq4Q/VGw3aC0QKDCc
OKHwPZG9n4cvQ4zT0XDfWeykRZ0IsLflnEJr8vGrAeevCzb10+47iYIgbRS50cC1EbvFeU7qyXkl
aC+uQjUaEW1lIbMYFLAyA1EX5Gvv5Zu/aUigTq6cJvue5yY1tJkToGbsimC0mfu+GGn72QVtN3l7
ARsYHW96S39W774nevyYUdm0Fa84gA+FI5Cup0A4nI2Fb6gjaWG2h4gZve3KlQf/jS6i+d6AMjEt
RAq/p0gToAk9IMutNNE7Hw9cHrxdWWS7sLeStDxudK6+MKJsYadHtWNpV9MUMNwfg5TcAh+H8rI4
FzsvqZZ4FoV2tC8PXQes2HhjbNfNvn4mqyibgntyaWYR5XxgKaxewj1XP+DDZ8DH64yapm1Ld0IP
jqJ28ujfPIp/t0LvoDwIH0Db4El6Q6aJJ8IjtJMBNXzRPwCrgRAv802BrTat01dg4wPVeqzGzQ02
jY51BHDOcubJURA3+BkaJwt/nBpbQ+/LbBjkUvYRpSm9V+JGPEM3R129xn1FMRQloqQQMlkuLcnp
7lEgyCNC3IKseePhRGjWdeinZTBA0ncseaCyI4eewGd8DFhEDnp5Sr202758uqhHF+gzeHd2AhWY
fzEbqn5JLDtXjn4jX9dvZhFWOdQAooVFUSaGruqQ4PW0blyk/vt4TsQvzaJbz7bR5SxiSYF62hnR
zJvSGuRxs8J4xwxDSgC+OF8tG15NHL2cukr/XZXhtk/5F6cF+Vvr16tR9S72k+aw46CFpz32cVk5
M4sx8/pP+i7jXS72+tVT0fjFcOfNB2SEhRH++U8xyfegR2+LoC2AUG8Kj6kGYbryHCY2Hl6l2mEG
icIK57QiBjC7sulUjkxNGz/rrpU5Cyi0ZzXvjdrX5nPx6vd8fdeggiKPz15Tw3/etjVnfDC7/LN6
2nAWZx0VPXMpHuBjpI+mAeb2HoWpiOpRAN0+8s6VDyqjegMWEQvXFmhxBVAQibZYjgjMUhqx/fAv
748VLkHsqbVz8mLEzeOjKQnUYmo6sy7BKKLTN6ubA+g69iTLphdXuo+Uvhe9EcYMVMkrF8peo22K
AvaUzzTSlE5aoYxB021JgpeyXLR46VExMkrJ2KMbwgKy+YZE2SPV+v0eOmqIgD2q9C+9+Fv9eySc
2x41q/tL7c6z/sgGzm8xqV1+zSg7Em2kN4peK9Cm7UC4BjqxQqAkZtiegMNFxUO3oHBcPyIakVfe
TriZu2XQ3FX1xPr2sBXHqGOAowJi74LrOJei0NMC+GTMifk/sjxFzBw3XvbphCwSRKtLUylRc8ec
+psXjDX4WYR6i0tJH6fDP4QS197EiDUgTNrGMjoepQSvKW1p48ygza0Qd6NQtm2KebZ/2y525pzF
sTH0SBHynjGAmG9x3cAkvzjLOCd4GnZ8QdEMB57KFEJWaI/tAMH0wYs0CqDNO3unrBdpff4k7Q4i
NlBZTgp2kdK2gkQAIfraWSkaLNeZHNb6ek4uW17M/WP9+x+MgtffSa4ndEDWU9JKYkACRX7O1ry5
MCF60IBZBeCATwhLle4eYt5wT2xYM+tOos5wJcrKXMwwpshAUSJrfCZBYdy0J/ibkGKxYzMG+9c5
h62iWKiybdaQCWLtDqPYqxLsjxIvUrkYHg7UbV6iOBCRpC4iDqUHoG5Xf5EiV4a+mcDhBhlL8Gpc
822oACQ+rdUOjK1A8xazOajmWiZ3ej/WGZme5MA+awKUhciXotinXh+uCgPoXsIE1EI/PPK/G+lT
3JZX4FiiVC2zVbxvONtlMlFznNsCon1eIjNVstmZRTvXZjYoQ7ItOtHet+jDOkGtmGlS0bU2oBRe
lfogQbXVrf3iZX+PQKT/BZ39vi18eQHUjau6Zroa7Gon1ZT99sIUeTYbMri1oSnA0HY5pyOroXqc
pOtPRi8s7FmZaAabqZd96J/8OKf3oT0+rN2gm8RQlF5vTeY1Fx+ZDL/GFrnuRqPQxG/WKXI+In5k
eJD/ar/EvpwX0QOqbzpyS6wZlWsHHhPs7DMvewYaU3fMYHvlhr+v81iEk28SDSgNClb9RTuZb5tO
lm9nF9vx68352aYRsAioce+ctCrCbBsc64krnO2zOXEAHMxa66pdR9LbFxEd32C20+92mLN1uxoP
LjTTpOxXm9brnCxL9oSp5CFoNas9ilCsAEJ9m8UxJH16jVn4gE01edigd3LgZRu2Bq2NR8p8eqoa
S3LAgtHRG9ediPhYhCaEuCUtBvwVRslDx5u4u8EFQPh9YH76hsYKp8CPNhWFnvs3YI2j/e8YTvvB
f4r6vLJjK9uxw0z9uK8CyglE1M4/Ki4SIayQ9v2DKllcYiQ76GKSafGhiuOnEXDmRRnKF8tEOt8J
Jx0+uHLtMOfmrg5Rx6I8vtwayBiAKubpJwUUNbXFvvXPyjpwmzJJe93IGtiEiqZ/IID6JI6Ow5K9
EVqbAqCs/pHSuxL9nOwpDpynayiLlt0Yg+2HKXEgPyckQsBDRDASmKl3sMwNs1Sh6pnqbE/XsXRA
PPRXHBgK3oJGNyXA1RHqqR4K3mtX66wuT786q/xZJWvpH9RpMzDr6d478bSkGLyDzAsCVFgPKqI/
Ug45bO+/HGzcr6CCXCbX/ujM85t1t9paygdK20rGwE6xNigM08F1Ieshjbex6ThefdyMl6//zlW7
eHpJ3rOesN+PIpRSn3eadva5EW+7zvyHrKhOk+0rBh+pAusWoVfly/LUpxQodRL7mJHC1X7Dmr++
FH9xFQ7mSMgke7ap7FmzYCxi66fsIxt6tzE61GHANQ3axIiM7z+Y+UoURXQfNPEQ7LLC2xfFbkmA
btRoArgU9kQuv0iyEOO/yo74Rk5OD9cd77uo8UPXDoFc/jgxeLUWSeEst1RHDmCdocjcx3LMjevT
9Fqvzl7p8PIlaZvua3RntKi5Ssv77bpFtSbp2VO46dB2q+z323T9O/lBfw93WFsxf0lnZvO13Eog
IQ7Rwr5B+55tV4PlGeukcStJVc//rUw4jMCJp/bLDD2znuTGBoeJjsxkiBeQDSE4BfkRvm0y93YO
XSsInd99UNbilNs+vNkMxgQF2IdNoF87gG4+wmj8Rr2v7G17zdFtsteOp7FUxMakO21fs82vZaU5
EFgQz6UQg+sNycsOBBCkxL6DnJ077Qdc4EPZu39lt/O+ZfmO8Ndp4olJHFeA3/ECnBgRlR6bJg1C
UNR6hYQMymppPjeGEr6+AJaaWDPkcBzMaPMa2uvLM65BktYMAY13FW8qA9QfulTfUJOXNqXRoB2f
CERNN563rffhdy0HCcYAiXO6Zy2mu9Datg3cLEkZijLJQ/uSW7Bqo/h6cFJlUB8jLmgO4giCFkct
7YOasX3ee6AiZP/ZCojvcR1rFOh0PBaMA9Uhq6dgAMrzv4tSfnUaJO9E8uOv40QRi5mwnG73o5ua
6Ywv2PPWfJpIQ/IT8/eibk++59sz5JFlvAo/z2sYe2zq3VhVxx2gPMpjVkt9w9mbXqMusJo46z/x
7A3ntvMD1ha1NHiQoXepIYgjbMyttfP+piCtuKy3XoGviXkdvvDqLtEcPZL0PGwBBnEnHord0U93
BNngdAV7TEbEIgHUcH6PZPs8ijLgaWeLxiZHshcreaZj83bplZio1yb8anedAjnO8aCt3dKpMsJq
/28/OvN8vPsF6dZYSFSkp7kx2tu9YxyyVSM35V3nNd6zUEGRTmWkLbUu7KRDe9IpLDYgTh8RlKfg
CuMGjXF7mtyfJ02RDaZQDAQszTtkwK6ErpLFogFe9TM+jbBa46LyBWlRGLB3/A8++bzFnITLMeq/
W7GPXm15+7s1vi/wbzT7cpNmYmLXJK9XWXGYAlFetgTx320BgIKwQ1F2ngMxZGI2lWRcjvk5A0Rh
gVI/LPu6xUSGebg8Rb/MjxhkWmgbY2NKBj4v0B3bcftFpoomPEaWR/BnrTATPrqmiSBklt4vYxtd
/GxaY2l+40AItWKzZaTBpsVZKVlK7RK28IWYX4U9TJUnC6a2+IWb/LMKDCV6ZO++jtBwheZ2cxAw
qOD4NJmW7WtLGeE0S5vhBqJaH/TCamNpu+Ldxn8ZqdWQ3F/cbmFfYsnPuGWOFZ0ziJXAjh75irNp
rVLgdu3LRLkdx8F8nxT/aUd0rRzdyKY1j7p+I3FQCUe2+vr7xBlqiMGOmzP4n6qmNdw5m/si7fem
AIbL2PZOFLUte2XlN1Rl2fdrBO1lDschlD97dsNgrGCl4Q08JMbgJ7VDo2jtsCrdhn5SZZLJYZ8L
PvXiYqcELIzMo/K4YFVyr0+McSYeuYAsgrK4oQyPYq94F19IDOmVNrIVrVcsde/mIAojxVPUKCGl
BWVhJ7FAm+m3NfLMlvMpol8YI85EuF45OZYK6LY+idLdL9wqjF/n8oKRSWkQTgr5kla0FIick4GI
lW2zcQhczNNGYQDJeFdpspdsNocvJYEf+3euNyUUowGeDvXb23pWVCmhA4LtyZ14r6e0hYPLGSr7
Phq3Z/L0gbgiKJvLQxBbCxSYEOqbfS6j1AI9/3L+GZuauKYSLQVnQryyWwP/Xz3TfmGTcJkS7dq+
BKgwDS9skQzZdlOQhYpGCfxqCPGlxGfZbejnFwYliXDxTTnGT4sef8KhYK+5KRVD+Kyb25njKQ2u
yRS1XNLd06OfBnlxytBJe8kbfb19HmGH4w0yZtDuhyKxKotrBmvH2cp3XIsR9aHRkNbRNioIGqfX
NEciXofX4R1DttTiNkjsqnerZjCHrIB/V3QAZ8yM0t0UC9KklzfEgbdpeukdbiBaQ2WLZINz0t6S
/qK8dfWG3XVdgPZ5ZH7FxgGBDjcDm4f1uOM2fBwXiA8xHi4KD0h1S2aHUVN470LBg67PZqnnpIu3
Y5v4nYbc2+8/DZ9yGUo2Bdc7vryCAqz5xhJvMLXZlnolFbs51TgnGAWPdDu/sL6UE96KhQLW/yW2
0Z5DsFh0Pys7V+fAIw9iz5dVQE7G8Vtgh1FFoU0DtOAQMu9YBxjy3ey5pVzt/mwa3YNIISAyc7sN
4cm7QjEGF9cIm1IjECyxavTSGo/MCxXKeQ+AUL0rAWgpyjQKMZmR5otj7bdfbEZKgwg0NCKv852b
+HRtqSJfcI7eAx/gwdvPwIlLjA894vXizehw51QDcZLA+j5kZKkBzeirCdw27NfAzK817aqR/71F
hNoy7SOGZihLJD7JCZ1rMOR/LC0xBcA4d5uiXlSfQ/y2DexhzmxNPSQe3qbS6evoRHh6RMjlgfZ9
XeKhKXRUzc6SCVlQc7h3XfiGxcf5c3i5FYR7SgaBsKmf2QZN5ywQD0FNwhiPQ12jfts3PYU/CEpA
R7blaTX7GEM+tGGd5u77jTKQIxdwhDL1Z1oqe2tlXEosucUat9hCi6hNlRqXvfUsI8oz/GrdmLuE
MAZ6ffrSgVdE0/fl+f4Lk/S8B4rdbPUvzVvh1DJhu6wJRXZCwjAyAncLA2dlsfN2LQbPIgFc6/LM
S6qD6GhkcVX7DIGZe7EdojpBG4kZkY7n1xXMhNNSVypggYU/+uN4VJUtRBwpbSlDSSRXMIeWQT2F
uKVmCP5p4KZa6keqkFJqm7YTvs84m7nyWCFKRhanTq5Lxr8nM55bq2xZTcmKWpZXZCZBUBx9QQ8f
+5i7SXASXJR369wJUJCNCuTuqyMGWVf0QuJRegGwSx4pd2NRNeTGKTOwmT8rrEpybcfu5sqhMP+u
ZMBwZ47Oul/LePrWw7yHSpn2QlJLM+53yy3XvRulFQbQu1KFkvvW8LLL8r2znBXDNJmYlxKHW5Wj
Zij6prahmHXoWDzgVQ0aswSct+M8QqPoGEnOn97cEGo1HOCI/7Is2KqngEAFv1trIBATPG0fJTSg
p7QGkK7SjMB3DPldQCwK5DIF/+uU17mud/QmnyDuILx4JGQDRpaY3rOTdmPhTRFe65hChYH9Ln3U
6DH/c2pS0G9W/JN5h7MMVeCFfcvARFuaJGGNe9IZCAiJbzpPY36f9lZ3a/V1TJKprymvrr873a0D
+lITNeWZiBZVTVMC3kQzkqhYfnAnXO8UATa1Gcf8JK5FcbD22li0FY0cppFKimfl5zmaqdi156jL
YYTXllgsnfCzkYMqc01mDNfJX0e6z9aCSYW7vuFD+zQtyZKGFQXwDDQOwvrIlhBGPMjOCzmxWme3
1H8s0Cu2Guo2INsuVCMFMuj6zh+09K+n+fyV7vGGJE0yM0fdQKwfQ+F/JvqGFr0ilFKqLJzxx8Tr
/luxJriL6baZxDBhOl/O6gWPjjPIyczHsfeoDq3dIfSX41CrcMtxAWIFoFCG+HVzxEGCvJ66BLkA
VP3MGGGUV3UWYu8StPjNSooUW0wePM0/UXzKKUeMsX+DKzlCXQuleaaPnOM8k0T5lw9yEW5qnb3J
qJQU5x/gNmZRfQsBTB0Opk5wue7lPDdLNTF/K1tqsuLtzCCKPwgMgiAEKc7Tc/INE/Nye0LaKuqY
uAbEUSKQfB7yzXeJyl6fxmCpNxtYRcKx7TPMp/XHvNN1BaZo2HcM5OEFi/34ZbtAMZINrCE3rpEO
grNls//sGstXXTNduXEP6fKe4MFa/Itnq9o71J3HC8vRpA+aRdweg/iXjY+dTyJJAu6RCP4yvSg/
JVitvUfWFkIn0CR3CtE5X7KEhE++ffVZej9Vt2GcT9BANEWK9V1+Ka+zYBZl7TdQkVSV2MwLTeNs
Ou1Eu8rZHSC+QgDOvueWXZJyF95eJ/f5DJsyxkh8u+RDgArBy4aFYK3bQ/2wVHR7x2ZBKDGmuN05
lZolQQ5gTTLSqvitMbmuScCl9B1dXxt2Xz2ZlynopUwXlA7XyGJWd6NmEGobfJXDtqRw+i4L4nj9
lrH7wgonscVybP0OG15uLaNiYbqd2sJismCTrIcrkwXT6An98aZBUmcToZr7tcTry0ZDexB4Wlto
qs3eeFbbivEVNG70Q14vJTC9nGZSRPztbF5pEM3qxyKriGXNyCu2+DxdaP+tmt8XHFtBYQ7ZjSVE
pMOEDPTjeXjjOZPVGIXb/27vwqidTweZvcvE9M1nEFLIu1imBO4gJto/e/Q5eA8PEGrEieFRqCni
r75Ncf6Ka7h2DMEaJR29GZEyi54TWTaXPJ44hRnstA9lTjLE+Mglgoc0ZVIqiOgXjRhm+FJxOiTA
cJVcjQffOj8YvK650hDYUXcBjxOkfd1cbgszw7d0IDt+PIFqrLFQ8Y7/VTYt+Wu6KxPzrYlca9XR
LGy5YLAHqQRJmKPbNoS7lGAcFP0f19dP4r5YD0isJV/UQrrBjdpjTTsy7fXbW4EsF1Ea1+D4zVpi
HX0EGHOWRsHYar37VJxpwCOhTMtGt3+qKunJdcmVQ37/CN/NS1SNg1iBhaj1JIAnzWOSi7reCj5s
1pJKeCCpBz+tnPPINl/5dxNMVBgx6PzZRnk6RADgD1ld4VBJcWicmhz322icQrQRkrpQj2hOoNeH
W8gVFRMxvXKspFi3AZbJDwrvPdhy0n5yjoKEr7IYB0ef+iQBF+sak3YyPIlzQAGGCJO3q4fJgW8+
L0uqI6HHPKFEwCaoz+zskI86eYEIUwcW7RtSMNHf2+Tkm0Q/zvA9KOHWWol+37YwppoYvTuiauoI
uZ8NP2cL+A6fx2eDj1Ez6z+zUrdaP0qL9brTZiuF1S7+gVcWlmitLi9xjkIqy6huYHzYYdiGXHXa
citmvcZ/UCkqxCoTwKsGs8waArkj2CnmiOPL7491wx/QLaRexK/pK3nL84U9BlsU1/nsCYFyoDF4
sO/D45saNljm8zkdYi2lhGLrnPUjdJEAkW4mtwEj8S4WjOOt8L21kBJsCNfKWeUvJhf707dDH9Q+
834XwZbDDjrPpRscWYJNoCW7gb8jXSQ7aBt2gaXf9tN6qZ8JdeO+82fL2XkEsFmWcGOdtY71f8Lx
OGv/hny/10a3KxId8RI2TfQuHGpvCu2bDslYSHfBw2xl+ISj4DwgXLdq1t6aekNwnA6o4u5hPKdR
244kCAYnMthhRm6il4vqg2jAnMeoEHl8ArvnFSKvsnaZgisccvzxAmQ10O6mIHfmEebmYDpQkFNz
9sj/cDrcKb68e65+8t6Flzf5SuaYCwGEizUX2nJ/iHEMqWCleW0hLTZVn5igLb3oO+wCaD+iMA1p
xuOKn4nvNQONTxRAZiXvlYknAWRqywW6p7I6C8pmJAYEfkI9KxWWLjD04/4YaAUtWaAYIfmTPmQU
kAxCaxIJgjZMspDOiuReidd/enRkQPK/STe0nqxhqlFxefj9ODkIhOr0xY4pDdupvZHY8xK3VxhH
72qYml+ZNHMNex8CNm8dvRtj2K7p4dwVp/edDfJuaYhUxkRwB7DmpOdAXPOURaPatSAXJVUiUTWJ
NwWCckszmNqKq5F4ekdt0eLHFSR4b0k2hvBrAiboDQsSxDrHKcN2cKIkknoBCLLQEKUo5hHmbfbf
0i2fWPezcRXVm+EQSMTIGs9i75TlPAf8WuM2s3J/RtyWExbFAFvSiYyQGttw2uh9HFcx3rg3lfps
zEMsCF9I/icJkwnucn//9eMkB+qeTpCfwLlrRFkWhiIODjINo5+nd8sfDY7JitB0QpNjoIWnfb42
AtIXgbjNJpjlReMeLi5KBfI8ylO85UeJnBe2lDgiYjwY+602Bna4Va+zJkR3y0VQaPeaB3TUHX6o
A30/aU9hNroVAq9T3bCy5aFwaZtGWV50ft+bA4jTQEMPCK8cR4F63W0uMi4Px4HKzkcmwatXCxX5
RzdiqrZ8zAB728Q7QgDTbwzBVf7ahO+NMjc7eSX1gCoxmzirSoPm58GoqITMPEXcOvJrabexBAY+
O/54Pt/sSlADAYMyr41G+as0A9WT71FBZXPj20x0Ym1Ve7Glet0V2o4cRQqzJHRNTGrqGH1OrSzd
q2rXoUtHu9HFJpf41T6JB6ljWJ3tAv6SQZ4597+bEWry4Fkn03ndsBCv0zKrZSbO47VypOldiTNq
6wJbkn2pVCp47MOGYOfPs1L/UojMB+5I2BQ+yV0O1tQoBe7uHghdwgz6uLJpPvQT0y42xJvzOhNp
n0dXwtlrWeCJlV3hH+LiMwewbutJdzhouBd+IMKVs1X6Se4vnEYkUk75fv27bKKYx9YUaZ8R3R5q
ieU1biyogahCX0nxhM/ZJohssihrQzqJm2dfQP51Xusm9T4ZmiVYqD6NmexeCGu93ZMnjwGgiaWg
5YTiAyyMdUbz+y61pr0/I9agXhl8sHJa1Lk9kzBV9/cLYmtE1sAdO9KzLeH+qX5/GjVLhh3t4XLy
T7w4T9YcJNY6IKo11BOmsCHbeCX9rdmq4avyI9GVyjQ3OQoAuijgXSQ7ggVZsg35RhXKmysnCZMO
NQ7brKY8PpolvtiXAp7anhtKcIBYITqwc0BXkfqKlkLgGucQemPEHJZrCWj5Gc6f83/xNPvXvVbp
OhwclA+dkHb+SCgww/7uGP5KegAdaKmPxa1gEd7WdjgPb0r9Exog8I+j1iWtkTIB6Mf9ZUNm1tRH
o9mklS3iaOPaltM8FErsY7Jn5f+63MH3RMqfOTIkO6jqmCm+DAHi3fEWB/2fyQq8ONkQNq6kcZqb
PZsPmA5cA3mPF8weXvGR1Ei5eEu2mvn6E+ulGGsfDvst7NC6rO8m+y2HSSn8p01v5aOp4zOqoJ81
fObJjzG9HOamYQreKVDWUKYy9mMtjP2J+5NPHbzZN/PZOvqd5/fBNrV4FL0IV/aaka3bD8VHdBxC
CE2ORb3w7DXmoAhgDgIN2zQq/PGD6uUUBmwwGMb36B3gnP5ABLsICnfO8eJuDOh6/+twBRNAtabX
2MR94cXqhim2W8g2zJbdBmxMi3kA3G/Aw2w+fiLPnQA7ePNV/08Wg5jaRkhk+DYjKSLAlqFliGW0
TrlHAxKaOlreUtu6FGZfUqJHV8B5L787NTj+nCE165GWNtkHXl1OEfe9WoApfRF9+USCQhG4rQNy
249fl6U3lQQrX8bGG3BMfhy/pbxbQtH6Yli2Sjkf7hgk3M4MFcWTMxh3vc1FB+uLGl8c+9Jx6qYo
L6JKGZgNEMem+SsNtUh92kXlSWXEk1goPbrRtAsC8I0JpMcDR8FwYak/dasOZOpOCJlIUu4zqurA
OIPgxj5+MNe5CXBQ3gKG5Cie4GE07JlZwo/FypX0Yv5fbOeDt7bbqWp825peGzUYWbfHvdH/KmMM
7U3rlNU2pnIM8JL1FKrStEMtA+w0cRrTLyxiMq2jJqp4d6IqDLFiBjarGXhVISqSjOaHmqfFxdlL
4/kWuvpmLeeEUkh18t72KOkXYgJzWVwNoxSQFU0tP6OfTZ3esfh+mmfn2qpzfdp7MZSggicjzwv4
08h1dEMoEvTmH53ewCXvKuXdVGTQkhEHmzY2E4LwVBFTBH3heWaFG6nHPaJshy3PO343SL4okBUa
Y1tcKvxq/QOynbLjOUXkRBUiGzJdBeAILab3i7WrkEyAKGU2hnWM+f+J104V9vcNezfPgjCAbFQD
F6+CoO7p1S2+i0q4CodHgYjUD3RpR2w/iaHvoJ1ZGyki7TXhGzj+G2M/67FfWltnQ9kY6/ITKmJ3
WY+I/rXyg31gMOzaGcoSe0P1sf50yiI6HMkNyYAucHbbankKS0AJDWGhcaZya9Ku2AKE8L6WrHJK
t7dTscCnYgtlDRELznoKQElt/ZKjA0xNJwDJyR3rL4BjeO7d5jgu6pnkcqFBI4sZB4cp4VAzKQt1
wJBeaRwSdofWxkxBkmiucqkvou/d9TZk3PssJcWUiJynLWq4S2PK3uE9StkMjgvPKwLlAtiLPk3P
5tKRm5MZY7vu250h0eyBGXy6nz1J7NlqpdbmwURS6PqI67yUhSXGJb+VStleRlEnX1TfdY11eZPH
k/XVPG30EXLXEvPnRroFg+O6tcxO9jR69KxP48H+UFY7gYBqm1U+JceYEXg3rYSJikWUTcymWl0P
VcQlBaDbI6KDkKVXbXyWqqho4bVSkcjG+day6zywgruI8UUYVQaW8OVxnssLC7J6G71vSWa4J0FO
kTr56ieFPCYjCmisIXGVti+OvLV/xeuVWumDd33Uza/RvR50rpp7bPZrQ4Ms9+AF7GWdfMOgEJvo
D+h03ypmNjMhgKYO8Gk4h+Hd04RF9eeXnCH3gA/nyGwb7vw3UKsNg/13fxxS7fDwomx78psT2Nyv
GU06cH72aRTAfShVfPvIW68VuOaK3OgoBC40JMnVW5crQP9xeA2tcYcSP3y5CJj/eMhT7GQ5Y2Ar
HJW7EK4cFcS+Vmp+qpJ6zR/9tK7p11M6gjqykhh4b0wDwEz7iIthpgfCO+jBwtnaaNcn5U6+D/Ev
AkcKSEpXAz3YPgnML1ELJ8+SqNxdYjgYB4JwSjP93iD4XL09My44pTM4Xotq1e8RCEgZ3J5CQN+v
hrORnTxZ9RI2DwopLu8qhbNk9aPSE09h4FZKVBfgRL/ws1kUZB88GlPu+bf8OYwgKxPyemBsm2Pc
L6IUM6oB5ZJVlwlGAvqUqHJxrEq/8c/1wuFNXPeEcboqy1g5bN/NyJ7jiBFwlTd944sLWpnx1Cv/
3zZFSqSTaRyI41ACZM6kJJ0fh+FXyQiAL2MC/RI40dVn0bqDTIJs18CEdcO7uMwOtSWAUGa3wi84
Y56O/Wwb+/xenz4vxoBeYsRf59rpIgkwtZdTyf2h9y6EBQOnkARnlIfS83/bSoJ1s2XdrdRkINWZ
vQ46XBRBqfpreP/FlmQMgGDZqAgswp4w9/NAdFVNO3dlxByIjf6+/oy+CyzEKvHdDcqBepq1VoLi
0KRawASebNsO8QaSiKTTrENnqaIKGwlgHDhb7JFsfv9NQk9Shh3nSL93p088JkrvQEl78EMjP0z4
zaW5LZocuN341VNE7G96dUa2ZNzphtzfNQ3l/aWShY+y+AKhaZ3/eCnVSaCGlfkgQwNdOzP3GqXq
o0jly0nQhz63V++r1EyEg73bhpRH+hGcY8mrjLLzAN0/Q1Ox+EwrGdQeXVTKcekxyD4nOkQU3nqO
pDOnbxu9q+ZF1Az+ykzle2YI5HBWdmh8aaAsC3gAFbBB71PAnqI/ZvLm3raNexkrfznZsYToe+ha
GG1QLc5cxoex/91qhdvDuRWZuG3RMfQ2B5JLBq7IH7M8GCUcsYn82E0woLp+IZzLiBBLfOyaBIJT
WG8SbpUlzmMOzUpYF5Mj85D46AWOb0HywfpnFTmgJ8F/TCxg9GccPm45BKaYG3xJ2e7KjQ0B4cqi
1djAHlifez7hk0wvlQhb/rILhw9lE7hqUyKBAwpFRqArUv07XlsA/oFy0W0y0umqZyilNtyfqGDD
8uS8w7zFpM+XdfuDV0hgESFgXEeuUDrhqTaF6rA5C0i3nQ8lE8aJ0XiGSMfgM9zXw02PrJ4/qPw/
undGPIgyvSWY6ACn3WvSrV5CtSrvFzS0vKe3XmWT8XMG+m3Qt3wuxe1XcYjgeJrTkeAeUTm/ar64
v0yQBuybiS/u1cYYLFOW0VmYVzAcIDWDADRIedoGzWXi6OUCXhEXdS8PD1WbFumNhJ/D6CN4ZpYm
C37bJGSlbIw2+jBPIyJSv2GGmLNwD4jBmfSgyepKoRAR2b5oBOsX0PJmhy96F/5Go3Dy13MrH8ga
5oZPWqh6bfg1mOnq/0c8wk+ggqqx5tB+viNiHD3OaWZ1rZlB2yEqUBvYYAdUaHjgUEEF7rDBl/i6
u/c9An6K1ipeikeIFyWW4o3DhvqFzF0W2KIJBfSS6HoV8LhdkEJopmrhR25Wi+rrE+OVjqcIpmzu
/f+Yi9wZDfjq9NNu9oMnjXFIPNJLDmjlyri+hrvhZsMhCPU6IX0FmhOBC/WwqV9Emg7nYq3LS7ZU
LuXXRRbEEUhLb10eQ3XfqEwaG/baeF0yXKGNZdKUwinEbAT/zPDyIicnWtPmqLxBScShJ879HQOF
9qCuaWqx+4MZC4p8MjL2OVbsL7jLUY7Vt/2go9HMWuUnpyh2sa6UOiJvNb1V3knCPLvuK1Jr6H6X
/owzGfcID/Sa7uZiQUb/1+yEy3iMOQuE915J/abK0mpj6cJheq0vGYgt6NYFpcEDd8H8AAj4/ul3
tOIxZfJ+Xw4KKvMn6SUWfAml/w8xu1b0hRdPp4N2TALqeZDYMxDZoXfZJTkejpI9jvH8eWyCPS1F
5Xvgehy++kHwmRx5vIwziypiO12TRKx1VY7j7aIPvuLFgC9OlR1kjny8OVGn7Y/odST4hja1IlYp
D2fB64sMG5yTJ8YX1eszUh1MmEP6xS8Muuxq38DMMpSSoDsNDcqc+RyEdVP2i+6yXrQSheFtZ80c
ZxFzXNX6yHhBOnBD3d4zsRgOeG7NEFlQ3Pnmc0k8A0qJfQZrW1Y+Ohzk+tyB8n7Yhyw+oVa5OrWv
Z8jTxKU9xxggjm80dn/cjfMjvfjGt2nQhdxNyi3fBO+EdEN9YeuzAIGkBPau+gAl5X+beExpBGZ6
Lyjh6NJcLONnSRr8fzJFufqo/G16E/cJheZoE6ou8YG7UOh/kAQS1xN74IMauV8Yqfi5WZf5Xk8q
N0CN/mgjpZrX0dqO8hVhe8Afj/3hPSxlzQ57Cx8Ezf7xG//Hyau+KY+UkHq+bVvTY1uEbtCrGRms
/R3X5OihJxm6iYPrWDavfEDjuzkKtiBB38uZD8xkcOAj6Iq4zvh+jEVOklKdcfU57ArCiVZKR4Hm
GyK9qo3bFYevhpvyAeZR3g494OWHZMkjcmctEqO2T8c5S4OMFmMmENRuEyBQpmhz/sWb/Cut2GQY
DBDFRYIeid4QnzY0htaTiVg9AtzAaQUMdw2Pp8bBP75CpL9rOmviP9dqWuP/k4Yxacpwmke2A0+i
xz3gapP4mDuRY2ZeYfPXEwcrcqnsv/adK2FRXhuOh8CDOHxs3aL6FY12M0P8Wg82sjtZa7RrnObE
kFq4e9wJ/6KyeEzaIGT/zQF1tlNPvQyVGEUgnm9g7S4taY0EgAi+z0qUNeHlNqybiaHytQHpkiSE
drsdTgyuG+vi29Iw/mt/DJ5LZ4AGjX8PiDCErTIXx6S9UXLEjsU7v2B/6FyubLQLOJ7tr0omOVlv
UpSBBH10SSI4IjgULD86dJroRfXFxuJ+nxl/xb21ziEwNHE2TRiYNeAlDjkdpw+/lz+VcMrnGSK6
c1YTXJfuF6IjRVvx/FnZKoQANPsW783KF0SdNDG58S8HGRwJ0w913p6hSWhyE9xvAXQyxAbQYoTU
ZB+LNjZyjYd6y4hwEbkKQLjHF0yRVA7JQ3kvX+sQ7bYUHpzmgHFiDbL+D2Nhp+nzV/tXlXnYhGx1
sFRE7iB37QhEaMaD9UZJSlR81gyv0/IBEH9UHj5LCbwxaXOpsZXHNe3pLliMhBV7G2tjqQp9lR6e
oWK9yrL6NfbXzQaLq8nxKyJrn4P+anC/NsAlvyim3/d3wllU0F/S+qqFu+U8rtsHUH5keATj5Dq1
rE0VYdevLljL5m2YN2lva5MHeaXZpG4cspDyMHf0svO/RufgbZMv3Z5Qub8Qh4qNxXL5Nn3kMTPM
syqGxPeBlsVIzIp+m9HH9FN2xaO6tq0dzawrPkJ0i3MCUC78ctzDckER5U7MaC0TiSCojgih4RCP
XCzf52mmdwCjdyJXgwd9yBii9UBiLjIRjiYcM2LeX2PXzb8FVZqehHJllzLCTv0seR4Ph0immEqi
yyfNnJHJk6VWnwgex8oyE94gO6K3DWtC2ddTFfZ14ppRWyzkOC+2RBXzmSawT4LpDRy5RP9X7yGT
kq7nZYfYWIx+hxxJbFXcRxZVJUzmSE7KpCTmsjmqE9DGx5yM3KaVQhRqaCFaTs1Uj1YM4+nljOL+
IEjDYkBN/CBnVNqeGWpvwKixvkczfnabd0Q59j7HymW2L8TQYY57c6cbwlaZM5bGabSfpUR/GTK0
zFBYrXbrjfTxXz8gxO2Yf/WKxCMIhp0BPbjGMPxuNWterOQHtpkluvmb9C5c95L+PpVQeOzDem32
msQmR21gb+OMZh8q7a9m1whk9rWg0vPZAO0nczMjKapLUx9nzL6TQNV32FqFnOiragaxUdoBTSfK
1Oc7bVAPqiYbQDZLCJM1ympwPFXmGzWo1jIJjL6XvXIzJ2ifuzaczo9IN8SxRXjoauCNOAqT63fN
s1f/JZzETDV3QdEatu8zpphvcdfe1gSn1feJuSx7ABbrgXrtZGojeAGH40n8s7lBT/7/bAjSP9ci
NDFx6u8qqUpoV+igOXzyIfkCRPSeGCrMBterFZrjGkflKSJawPhV7IigjvgjFnrJmO8xe6X2E/yF
QQhEN7dZ4MW9TQ3aF5TQSIfAitzv67dQ0xCOP1V2tmq5rcqNqx/pbT2Qchh1xAyi1ieGeKOH7z4L
pVEsbnDtuunl/ouIA2gRZ8JDyZxZPxccECv6eUbwrNQMWoia1qQM4KbQ0/VsJIHUXtqyZICKvZcP
bti4FRCSs4mFHhvmZdHhmujN+rQgwkrjd5GY+LfozTMP5rLGVUFxTel0OQj/PermhGrXEZ0KHH+6
tHP/MkG2fcsScv9bgkbsdnAz48MEKV8EC2/laR4/M4RORrxGJmp54mw3DbnPCZ6qwC4xadZ61Zme
6+6yk5+VqDbRfaofUGKIoZFs170tCB8UqEndz9OvbGGhIW1DmXniAeB4v9A1ztmBM7npLVUClAZQ
iwaH7Dz4VC5q97rR3zurzCDwGv3oAJkGlIoO1F6eayTGm4FUa0JdH2RmGTRmTA+HtPmrKeLnff1b
Xz79P0pOKhN5AfT+UKDpvGpFc+dO7RbgYXHKxcMCSpefWiMGXFosp3iLh1fR7v33l0Ykw7hvZHyR
ZLzueReXXNtNl3mx/jyAP6uVG20s9RV3YRMiJtETf10GK8WYim4aB71uXwewYlipJTRzWvvDFh1d
dH+w0r4DqpHuZJpKZTO2aW6/La2YrK9ULnrGB83TqbSOrYpBup5d3mn7aARi6MNcWh5o4oYw62eN
1SaBUfnoQ8ZJkHSfB0TjiAqki6ht6hh0u5x5Q25+/kVRbeqk6KJXU5P+J3um5ePxPoFy1+0RY9fG
So+ZeRz4wIA60Y/SNtw979i+ENQbOLX4aO/dtZADyplZLfMTpesSTIWvi4mpFeJeUFO9xKF9xNPD
hzBdz7v6tIdYL55jX2HkEdLN3RRxzYrSyH5isAiIiFokyG2575LXphqcj170ki9rn4otYNO2e1XC
tTVb7eGa/aoaU80D+6wrIzBHwlx6M7gUeNaKCsHeBcMmL2LmEBFsDlA5ZZmGxAdN3zzyPMZmz6hv
gDFGdFovUf1omnMU38DHjauQnIiMG2/92OS3qq3JUDjxLoi6fPf3V7+MlRMHGZxeFOaN8Qjd8wkX
s9j28/3dLMk2YmbkbDqVT4IF7b7au6IFuh6RYKWxAdQlqMlX83I3DRFk7DuM5ArrigRd25NjT3WV
qEGQEDm3+qL1D1FnwXZsH2xNE5kLW49LLJxIqMgQYFeqjJR+HAt2XbRy2Sh3qRTnpk1RCAqAjFcH
4uZIFKot+n7dGRQH9rkUxJsce1k7rzdwJKDRPy/Vfl18cfX++b2HU75Q0MN+yrFpMsQCFAPJwZdR
YCSDt/nNkRfnfhlPs+bbZ13/pwFNReJX8OglWwvGS5jFUYgjVBuPCPFc6N9dYgwUCVv73KPF/TiR
Ss8MM+EtHtwshWeVPYi2LEj9Rzfql/ac8JGoPeNOwaA84GCvCWGwyQtwZNqb6Vtby6h9He+5uisM
DRFtKMTXL/NpMgujHK9PAO42obrwxwYl8zNkfOlwPiNHKojLXEez6RftuqFkAhvc/zR1QVNfBQA9
UXlfAzPOnhcVvD5YHtv5h0hu0S7VQWxh6m9y2tg1iMcHhuk0A0z3cyb3FTovrP8t26IZwLfe9iBx
DyjJ759d4O38ZL2bPKp1+SJom4AestYKCgiJELpflhHNqX4KEn3nEYJaZsC0EiSIzwC7eBw5S9Mx
2KC8ZAG4iIp5bCRo5udgJRLIkmm89ZGDQ5JWP0IAXrF9acs5IV5/EejSwIfDduVAIViLLfAoedio
IG/+DE/9fwsl4H2/jncfDPex+/+3qcGVD3WN2CEtinnD962GcWUk4RQc9a82ly/SrF2ZnvVEgIb4
Yc1I+fnqp1fwZt85Juw1hNDYEy0wo6qZTt9qLwWx15YBKWMuhwlFypPQbc9w2acmzN+tSYeHp8Bz
Xpuyxa7ooBS3Ynqhs93Wkb4EJZM/3mM4gLRf+4ueuk8rujjNlxw4oiQNH4BvgeEI2Co5P6Ua0VoG
1b8n7MspGXlZDQ9c43hLH7p8pEPfxd3+JM79Ml6NASzn5NMUYOgcfx9T95lNoB4zq1ki2la8t4eL
5TOTh/5eLCjQshXfQXQMW4LOfADhNUJGoLJBH6+lM4vdAt+k9GLsd3W0eG6if6FVvgDZh/iZiwpf
+jCJWGvsPPLgxFmuEuNTPe3wPLCvgn25BfBEqETiPbFbcrZsNwuuFKWhcvDVyai6aDFkRCyUSa2K
DPUtuHEHJH2ybWtmWysgOg0sU+ngug7qQB9ALRuBA49rlnhxVwJ4zzGYAbUKSS/RhhHfTwqW35TN
+61T3EYgii7fbf0yn6BCZ8VnFVUhZEwdwxD3bYdzTqFvBT3lqUKfBO3qNwpqbiOh+E5HPVX3JGcG
aQTIufZFxVPvetHkxim9CPWGjlYTftbD8+BdEg5HhKaC8a49j2qTehbssUIZjQmhMXqnVMmWqEey
JZ35pvTSuP2apjJTlDloHOIPKWbYJdwnWkGFoCKRWp8k8PbUV1SwDi+x4gLjLeKeTkQMqAyhLrHg
FltLPlte5IcDAUYADoW8i4cO48GUKa7L6TtAuEhkc/NqOGae2ut/1B0dppXcDSG6bK7+EJZrxpVJ
OxaFKAwLjLMDxiM+07FTftE72vY+jhwl32AkMfk5nWj5oRYy3DI7ELdyQCALEWItjQieW3Pmb20B
CKZwIPx/gvIbqQL21tkWc85uEhUZTXPViB5WUAqhWPB2okeNPYOTL7d3csX0AZnTimi1Il1XLU+s
LBUCWQmxYEtyGoK8faoMIE0RLKER7TmiPhLuyyThMuS/hDblyjUL2n6CuyBvEM7XhlGDIFCJE60L
w8TbExrvgI4T2eflEegibEcrySKKxE92Q75vcGamMUyQBGuMrhhX6fi8t4Yfp+FpDXmr0AlPWifF
fu/QOJnUGN8ilMd6mXsOx4qznM8XhsrGB5RCfVKv1CRAGosb+s56MS+jUXYKij8GXp5JLMFA/KIk
f08GSoE5a+EE/9S2z96lOzEPyzpiMyW+Eo5wqmYNZD/i+sqkPcKxo2qmwdDAsQI8M1qxOaQ9mrHx
cintjvGTWEFOObcdqVYYWVRPMwOVaCy0spUWrhYVXwtgv70sdD1jBPQm8s/yn6FY6BVjYsbVfhPr
TLUOzkU++vrY/8WvWrBMb1zK46K1c6tjz5vkTG51zssvBVtXwJHvaObX7kQ0AMRk5PA/RwEQk5hq
NZYetY5qLNtXZfN7C6/3PDV8IeXyiMBslWtjsgJVmb3DGUrrd2sEonZGjESKhnrDVU5XckL0AK4h
DysRM8wmv1u1N9Fmy44KoiJVb4cD1G6uHVsfWCI1ZcNRqphA/pVrUQ4oV5JCkUNhKUt5bCQzCLay
Aca1KOZCvWD068aftGkaYNYBv3OcOzwjWnFcOmbgKBEgBGTtkb4f0tgeJFqhvjGxGXScQhU4UdAR
pQ3Fd7iVchAROWfkQISZO1O0sMoxmJdBOdGsq0EVisKZqR+ttUhO5vT/k3ohv5FSHdna
`protect end_protected
