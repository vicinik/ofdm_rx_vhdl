-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i9dViWhX5+ur3kltxLr3EfxORuHNuRw/SdPQaN+ed6nsHbbOdcjvVwApzsYfiYWgmpT6QnRxNRpr
GB+4wXlR2N2NyhB99QRbgDUmP58JYPsS//x2IscXInKa7CronWt12LZKdagcAeuZp3qKtIsSG1bQ
i9AXRY9d4zTji/SDYRjrkiCep7zMMR1dcG9yw4M3+zSvUoGEANFSLQ6hLc+QzSZG5LG6axBzbfoT
h/t3HMRIXzxo2EIqPdoVdDdIZeAVLBC6VwH9Hgf4oWzX1c6JpMjrjX7EiOtunIwRtdiIlpBeU3pW
IvFcMmtXWqiqOBU6p1BhIb+Q0pCV+qcXxythkQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
+Dq4zwlLeRFPNjKBfFmYOZG4ZmoCTswTgsmgX59+Rivml0YPpCdf+wsi5s7/Rvff4a4xWqhsTKZW
0t5NOgtwbSKOlihz0Ltcx01C5JysTmFKxpZGCDyQ/v1yMhIkDOpgGxLI+Ygnom/FrB/lsOKuVGuc
2NEQODB/fegZpMKX2Hy08hje5Xm8PZ5vbbRlD50zsVnJnq8R/gfbRKeLG1C1Mm1UxrK5vEu3Iave
bIX//J4eVbfJoSxobkhHk5CbyIHn7aNUvujaoVenGirEJ/RwnDqCs4bQVWfRs+nT1XqVK3UgKkyw
g+bFDqZ3dOhih8gHoffrD+oOGZjGHXQxOHlx2F3rh/mS9hU3AxtF67IOi1c5ie2/SjmIW7hZwDRo
AKPPn1tAhQJTQHa/wODzuQdWY2p1QpvERw18G6kHaMuLY4tP2L/PmeIhgd/7ZMa0IlOoXV4BYx74
dcSEIwfUDfveKgMw5qR8hcbZWoQvQmTevzZRsq86b9jKBZoOiZzhlzl57B4PSqq4+Eo783hrDFMP
D/UV2tdJrKJf/jZvoPVTlDymBTFROmWYp7DNZpUWrYbF++kNZIbwLRGq8SQI5gi2VIa7h2i2sEFW
e5gf7h5kvbpNdXZK5h3KQPy+A+Vm7CkiL3tuqf6OLTVqwdLRJu4sXYNJTHLv/I5JvSZY+RSc8yzM
WM0qPQedCUtMbKaDTcqGCpgjWMu4WL43Ftg5dQhg6JxeqTWO/GP/or0PpywVRxUW7FP92QLaLg8r
qVDAUfzrt/uLWa+GXfu6AUKGGhlUyiOjvWs+0njz7XgQ3edqMZKrDKpnKFpPdoOH2rcKsRr2Ke2B
vNOHUF9Ew6nZhnd9QB77WGQzQopWNcMdyafcvORC86uiCTP5nFLxwydAiPR7LQAxkbZAvA0o/eEu
tENpqwZPJlHkMJFveePCbUYXwLgSmzh79xKn6+SX/9jDL8E6SjY2DXeU48v2m6GdOVQ34ZZ3UG55
6MNisMrQTF7QHb/5wPnvDRZfBua2Kv6/Cf4ZfWsqxsVFC96AObEDcDv3Mu95F4GNvM71wtNdHvMO
Skhx5KBxbfpoAJuBfUaDgMCY6YFr1Ho19OEZbwR2xLup+0m3MmN/7jPdDxksXyyfQX2wPDeSmwKo
KM+Rbo/MV5jnmUyl1h51nHklhPBLPpQ/fIqj1SdDhI3CUjjKq9PWgwjqvOZk9XuUx7GmzDD822uR
kX6FGLIz9erU1RXkAJj6fp6nwota3MWfbnBj2KFHourA+ANPhEvY1LYD3XoJgadQyBLNCQ4GqflT
1zdZ57Zt7bb/r2/6R1axPgA/bLXMfinEGJr5sdoSCCyqJkuGdSVBN4Tr2YW1MJZfpnvJ0omAKglA
wiOypkNm5IMLWjN2eKEtNq5rjKKmGr++buKjlONdR1G/0iarfQswEpBJfnVPwDrpyb5KCgvXmEOX
r29ORcZmPTA8OB9+3KrUWytWCsn1LmYg/WGQoqdftbU+e3Vd8uE2DUEGepIGg8CK9GD+Q4f6a53q
zeJHqsgW43sYtltwYzXQVbsg3fvlcd3NKDQLRj8GJPX0Pj4XrYHYQyMOZ6Xo/VuZakGM3YXL9Vfj
dCxexfR3mmcCuVYF+sMXp47bOwBZxz8EkoIlowSYM33SLGSYflnBaKoijQmgBEPK7ujZ+J60k8Sy
Ove/nyNUc/Z2+c0NJpUVdo+SNQ46SNKZYX9FhZESeBovyI94LuMdO+gvWabl4QXe7kc259wULvVt
5PNY28aKuVW3Z5XRI+hoP7/pJRtLUnsGl1MoxLE2H5yGw6V0UCmiW5+3EZ8Nk/LhGWHvgodu5adH
uDFPHwb8twx6ERsv64ltEVaSdEuHySZmvu6gD0DAGURLwB5YzUjeH0iCLJSWneJkElr53gIv2r6q
KyKDWsvyX1hHrXLkCczr6Aog8hR7tER1Mke+DxwEPmn2qwLoiw7kgleRbYjK0AuGcyR3mazEetKv
C6rlSnrK97kbhA4E6jf6dudTqYWsMdg8GuJG+TDnIS0+P64b4RxeQeyHXACGrjsuY6aQ1042G8ad
+xMT57bJpUgbVd0tkxAggPq1A4IXPidn2P6nlK3a9hjensNHtDxnRbc68i7OeX4Fnz5abQf5QazF
2AGabC/rCz1oa/2qvQ760Y+mhqdfoNZWOE3EOmsmKIJ5vT329qKsd2shbrskEgNPwnwBc0Q1XJQw
J9EXOtDXUfmHdNATKoz3O1RXjXcDJC9zduFCUBFyY+UtXtdZrPNDlj//BCF682h90dHgtjmQHD0Z
KdAqs9CD77iKBaDXzu7m9kMKd4bkCf81uXJRCwZ4waSieesrmmWT2SeObRqPvCdRo1DFquLLsOKN
uYMrrLXqBjmC7MwmIY3pJ4obTKCMDUC1wBPSzQjMEDpF2ca6RG6G5QRC07j9ZK9goMvBCJ5H11aj
5gVDhoAPlXIx8A0wQ+paFFu6avR1IPPNu0p3LNZhFd48/qmqN4gfLnpqnKUUZLVtHlehJ5/MBFjY
NSsR1evq1pFQTW7JZ8YeVu5M+N9ekA7hQWJjUHiQKM1kZTJyiwX9q8XpmlyhDraR/Km0dhxWD80b
Com2OadR5aDI57me/YN/ciqZpVSLYcL3RPWFzQ//trdCRQIUiquROcgXGxmwGthqfSEnrwft0hBG
ezepcYfTsDUTX0zyW5llYhMUCBQu/KBIY9/w/ltOmoae43I5hphBepyszuo9ji5ndBOZDvavcsLB
LVCdhWfTKySC5fxH/C2i9bqSaeSWmvj/mrkc8CepitkHTLjuHRlltZXALFBgUMUfIPAiSDNmS8mz
lSWv0sCXzRdLR3vMpEImRpWvqKM+R1tyNDdaYe0v6pSMamU4YPaetMbFE+dJdAL57oASkOebn5Xq
nV7SqW39ZbA6Wpfw5i+TzcSajnKz5+gTQY3ja10HIFEkPEaWtxr1OvIjOW0GeVSxlo1FNglfw25k
roa7P3sFasbD/+fXlWXFdp5r0pYyQp1Eu2vinUnIEHuJWjz8PQhpc5sqInOxiELKETaOrBjovevs
WYTA0SB1mIIy+/0Na6unU3J8B2AYfZwz5FrOOaDcJ95SZk/SATawX1nm9C6eE1T2OctYGsgpw8vr
bFWnq2J7PmMh1dcn/kSG45dPHfnc/6pwdGgqb24u+WDBsmdBNsY0IU3mozTlo9G1XPkUK7rstPQG
hxg6RGSA5Pp8HWO5tBzOgCeSnb/tvcWZlOs/r750hNFq7w2gyj0DGMrYE3VrDdjcJpR1hHYcY0wI
xROZn0j4fzZu1H4NAnd/BkNt4ADIBBQFilMIxcCJhoZYOb0EaFu9t3fP8RvSIht1e8jpe5JOdNTL
RprZYRB/L+tQOH8mJW1ycSVn2NUvoNwrJn5ceeap947Nn7pZqQK1BOFf3miGRkmXKynmgk8irgtu
xcMsi6MjZQxHUrB9/PcnL1xMR5KP0iUr0EEcBg05lMNUsl21sjjU0kJ20PtYP3YV722E9SzWlmgJ
GByX0R9ZBFznmlb+AdEoB9VqdIjFfApVd18gImbQoK4e7Pz3C/Jxtm/qtjnoYGs/8JxT7gPvFnk0
W5jN22I5EmxNdS2pPx77RgXgl7k+89GLw5RtJFIf4mfTaUipC4AZ9G8MRvY3HwJA4IYW01Ot/XqK
1vL4l4FwXpAug8W2W1xTICdRyRjjToaTcSph+gr44lZ/xq67ROd8x4yakDQFtac+Jj8KC9xU07QG
niSR++tEbLGKN7OwA7RE6oeZnBfRUqN1iXamFd7mWqZru0hbGYM1jfx+Ir8zIOSzUmYdQgdcKW8c
0OINPxONoxp8zPWO0WFicQuR0kxccdEc3ZTyLONF8tCyUDae20yC5rc+GlhdL01wAjV8OnG+KP6I
MvJ7RmLri55JD/93RxEaeoTEp6K5P5sTZ7CvNCYXMEC+h7IK4ry6ekRqTl8CVeVQUyrn7uzHZ3pm
TMnd5tqIeFjqebRc08KYVWfnARTNJcLYUpYy8l0jxXJoVcOEAgyUIUcXUPBMS+TolgJg8RxvQgcw
qKaSe0NFXPqWHeiX1ynSjLb+v5+zHAGhKh4ide/96EU1pPQk5V7OkQ61Nm63riNtZXrZHuQFQLI1
FdinIUbHxbY+79fQg7LptZJdfA63Zaap/1QGmaLj9sTQRpxJHawdsdM5BpgRztfSpn5Ni7mj6Cy0
nTdzLNlR4XCgQBlxGH3hg7vVqiso/rYpcTLXWLjueJBO9GcaTWE44H7Yb4N0GNfp7bjfiw4qncJH
J8L/xJipH+yUgzeu8d94XbLHEZOvCTbPqYEWEBMHqtOj8cXTtBEzbN2a4ETEawyJXOsOKYcrZcyT
l+zoXyZbAHHVZjzPJEVCHXa7JAnj575PhtffPHkEtAm99P5QtyQ7xHh9gqhykD4VQoZCK9Ob0hax
26FmEIMuGKzkuw4yzz8CwAIEDqxk/+030uvlx5Yky95Xo1WnT3Ue4/lk70uJT+G7OhNeQGRmu5la
YaERpySVXwhbc9LwXaIuO56+jpOrusJ9f4R21me0XQyqoNOb/sJyXrVOpUCe6uElOLzd0s01mrt8
Q++v2Dh3ik2TgaYcLwzM7RSrWv4nQE+CmoVibvpEMMWRwiMEwY+Ci2tiStuRoz5dOr2AG3fBDYHg
vlwp6RFyEzMUGO7DW+j9u80+xih1qlGo+dsFpkz/UFA81NnMGu0Gqn5DqyuuOHNJeqXow/KHYYO3
svuwWIkLugqbRM9djWAdrTTqOGyOEYQ7s811I4PllvBNB4KkiZIDOmqcDodRguTZZecryhyiQFtf
YQSFbNuKL0S4w6+4xp6eS7emsZcM2LcCXKIUELoLxiWymqnioPOXHTbAWaP1T9vAx2w/GR33W0o0
SpHnn8nAu6Br17U6b/RJureFa5bKpDA/iW6EDPVhoj1xSDZjtfEfc/CNK+nOXPmGlUgWchfEoPSA
Ny/Xz/s04tCRY3nt/VOrCf4k7iqNRlSFp19PnQhmgQkSfzYURFNe4sHPeh17CW8jcEuMws3e2O6e
qY6xGvILCnF5oIM8GGWU+TIx6tp0j70+u217cS4tyzNTz4wIzfvm+CjO1KI5lSMD+hGjrI+VQv54
WF12e9LdyCCHmjdeYO/046v/b/OcnxHWOcm9cIaK/bLsXcqUaCGoYsdRa0Cf+EjPbiDKc6SYIDMZ
R8ijaXC/4bXQV0LftBJw5NPnHaBMk0sCXKt8jyndr3gJd+Di/rKKekPJur9odUE8pynr0mfpjag9
2jDmiJrDXruMchP1IAlAkCH1JAYoXCgVu1PzMvI46UFEB6hNEeNfQjrAfk23NzDmcLy04pr0TcWG
hKMkTX7X3To2Pp+3f7MxpaR3Ksac1erEoKLII+Yswk4bh/xmlksalKo67EeMtroCbjmT6t0dzx1G
JKgP0k0rDovNbjWIXEn0ZJ/txJh/Akn6AActtSxnBRHrZF+cwrCUvLqPKQXWmHrgynpFy/dsv3bR
riQm9o7/ul+GYmv4Q8YNhAe+PMAePjXwrwYaLC+EXApYRcVGYFhKjSHHUcn7ucjU+urKjq+/XDzM
4A0yM38Po0tOMNRhuQ1Be31LIVOSi7xM1BV4dF9wSI0OVmCaeyhqoJMOk7abIMggIf3fDSe0FRLH
6A6Xx3RD1afDeVN+Zf5SJGCWhcEO8bBbPDBCzDIEMOLdODlYYlStOlQa6Jwi689qF+fpSl+n0RXw
klfuhAv7CTC6h38nLHyprkmR0ixBYKtgIwkplbq+IViS5Iu/tU40eJwGFhYAplchY6L4M/z77stw
tMTdiJYgxbLBNw3ayyVryE925vgVzY4ogvzadkL/orRZHiaGh1cg8RNe7WJZKWq2BecXEp7eCLUr
Qiul+8p8zHHZZimlEeNd5Ok6w2qUq1sPowSzfhr5qDb5RPCYftqxVkS9j71ii/wbliEM6IMf3ehf
W+WItUIorgIChe9FYnz12jqSRJM4904fDWZKG8YDCpZq9G7Xk0Mv4vqfTc+6ht7mbUB/rmVe6wlC
2erGFmox8jIXMfzYDEftwMBiUjgEDfVTFRAdQufOboDm2Z9pR4ZHrb/1l66tN4LGlyjFVScETv5u
k7yXd8GareKZN3+lDeYvAREGZY8w85AeEWikoQ4HvsQWRzTSTLmYqph9m9vVoN7/pjYsqrBfIO8H
I2bL+2P8Zjy4oTlDKTCbSKUGK+ero1P7VU9/Dg0+m4wk2hGqRy0bmK53AWVsNwMWO2vb2C9c89+s
NNPmxz1spykors1xbDA5qNw2f8yDYshDngvufG0/XEtEwF1yfv8vHuy3Gw0gI1q2oovY0kpOFqIb
nXjZe59wkJfLffBEJPuvzUall8EQ22p77ebRSGDpAQTUuBJuYLXrZyPR2S0vyeTxPxOmPI4xEAqS
nu2pXRV7ktItjT6wSDgNjyhQEVWqrzvyi+ftMqazPdpWYSVyA0WnVh14CJC36Bdmkn9ja1tsbBRs
R+pFLVvmCOFBHqC2QeLJh+ZKbPzzEqAiO6beTO8gksZEytlYqNfLu4qM6VahUrEEhHFNMZxuV1nz
ekY/de3B1MXZxkffPgtRkvF5Twi5BCgZpMjUOVtNbR6r2yjBt3lUUuVxMfRLI2ysIlnF5ALR5DLn
UwMEUXPKdCzquLfP/nQJ8MsvBPTnYnPy8Mxuqrzkqpc/STk43Qv+sw1w49rxouBfvFgAI50SddEc
/jn8r7dmhu6IZ/e7OvR3IxKMKTbsLcnDtSc8xpJuVFoMce7+BmEplvxf0D1HTKtGfmLCyfo9O9/O
4JVNm4NqnSxJM3GhMDiSiF1/y5hHU5fItJzE2/P9/mc2dY22zxN4t1w7duGYdhdcC9Cod/Zhr+Uo
4kcwz+WiZQ98rTeFEKb9x5RjDuRevi0N7XA9nt18RN8e3Nl2KQwY/JlLqzc+rEKCmptUglMcZGif
6z21ZqVWOwTfKIm7Ng4R0amt1ovzFaJKhQUn11BAGvG4xA9ZgDZFsdvvPi4dtEzjKVEAS/isE3Jj
uatlf0mahDWqXcCgzVpZyECcqLS7AGNHwQSLoN3Lk4sT14wPCvju+mC+Hu3qcoMSWgBH23mDU9xt
IapQDZ/T+B3NOetSQHuGb5XWwhsvhxU0CeBvdb9VEoKqbYCYoEll9x8J4N66Prc9YEm0hD63wW1b
xVKYkNAbrjAkSIozUCaLsvv1hOh1DSnv9praOtNTMvZ0Tei+w1a6VhtP3iQSP03MYpGuSQDt56zV
Es1B0nX4tHMSKZLH0q7qeHprfMoPyExRYJQbhe/c//If0c+DE9Th9Tf2bJfjntbLVxjbmxFHh609
a2r7GtKf7NIzd36CLSvvbna9FITimsV5VXEPq6fUk4xQPLzrl5zcjIRsqQ6/8sCkCSyUgoLDqBbi
U9dYAle7my3bXFmoVtfcY/Hf12FCMfXZkTWudSt1TUqZnkTX/bfavgSBnusy5KER3uL2BTVF/xNc
GimjPkvbcUAy3Ig5sFZDxyc9BD9Z9arEwEX7HDt4OwYgVz08HFTvggwt+CDNWGpWz/yfLMlcqQ+m
0DF0kO4XfR20dsERDTk9qYz6z0WYBJpROwR/zkz2co+J3O4TaHveBQFLPRgupp5mAcet9be9k6R9
s60YSAW370e6ZutXpbmMhJnL5nXLB3L8+UFfc33hyAPPs/xQmJXhLJTPzz/qkDuR4d5rsDDYNV4t
WtWcap5qumYfvR2AOXinq33nDjPXUBoujN7oSEA+yCdmZSriKUMGnMFE3i9jzqaJM5ADzzTewQIO
dRfUcv107yXmWGfNDsdxN+M/9IBGtmshGThnvpjhFPrAvOKhQHKPfHMaujg6QZA6qEKE4KB+caEd
xiNfp9aDV8mTklEPs8wEN0i7juksMsMYSIprNGryf+/BIIxF+hjgXrxaFAuMJldkKhaii95xhH0l
xiXNueW9G2fRLwVa5kj8bacZGYKlQHCQrmz+ka8wBvyP/YVm2GN8xk1EGqgcrspiINPcsBiHnRVA
RzZBLsPh5RKvPIgOCmGhFaTII3kbc3rF+8JHpGWnO49If5UPbhKgMjxJh1K40RajkU0LMB7jO3FD
vxflkG8uTpkKyY1RFPahKpcS6vfiioQgHwYcsauwSA0NHy+5eZvug4kzsf9W20KC4MxW25KmANMs
xZFD15HXFgUk9hm1KXhGb/x3FEBH+JDdoQJKfI43ZE/n6MHzIxjzxg9G0yqgeYGeY65LjzL6TFUi
9RHl98GKcV4tZQbLZwI7kJA4UA5827/iEz097U6RG0F0VjWQveuAJszrWU7nmRYs8slc4ko3c8rY
aXktHTe33Oz0N0Xf0PXy/V3u3AXafgWzYWKm7t8H9bfwgaNEQK84WOq1F9I2g3krW/WF0ZbhEQbh
44A9Dfml65N9EGVlKdO0d2yAZqnxGzhGbTTyGHQ8KYm0vRcnLxLcqydDBf3B6FgDbftG+soE1m5X
o5aAi92W+IRJvazn9yBCCOlDj/lpwuoV7RciitgPvsg/ddGWYhDLpAtO1MvkrlS3wy+j+o7pETDi
EhDuVlxfT+9ftyB3s5rAIuBoJPpjhH+f7BhTEeIhrdEHXD1bMFAqo94M2W8En2anLk7FBu6A7cHS
en02JISxLnZehEOTGPSGdhIfNgRPE2GFZK6XqS24xB8toyz+Z+8g01tACMOu4HP2ZgewZC0MR21s
jmUN8ljrkZC4FKem6W4y5B1Cp3nEMqPiLGZLiajLwd4wLyPaWGoNGaO0q7HZuId26Ki1dAOi4LCf
W5nW0cwhx8NSrImHvuUBE0rn4IS0LBIKDibWr3uq/RKrJORiStsijUwUebpIC1HKM5VOgonzci+4
+mxoZDFlN9HRWVLobVcL8h0FPDtYpshtCPID9kQx+Y19mNFVAJ++qteTiH81INmlPUap5iSOJvnS
gBoaoMKV0v9auB8iBu8X2PcgXRdqp4j/Q0PEvgPp074XU1kDDrMAHd4V9NUVlbdXH4JAGcGvDlkt
c6ZQMbSUAbKvLtXVevMA5t0zezHqGQg7uPTYLaV7xjnnQeilaIMaosccYQPvAG1SwKVIJEmuqzAX
y1c0/+uMtG/sPHN9ODGNc/icIuajIIhV7DOciaNUeBsFZTxUTiIc2mR6RYTG5sKCvtisSUnN/lJf
+cWDvWKy1v8ako0vPCpdweaqJ3WrMtHdyVgNJCgXm6nbIe2WlD74PYzK4SBNwc9hLcmlXte5w1yw
3RpP9MBdnnTVf6k0k2gvLmJkp82gs/ovk80/xoVZCFwa1/u8yXOseOd33zo1uCV191cRKRpphrZj
M0ydz6jWpn0Vmss9G4W5uvmY/4+1ZCY0Ep/1kkQH0amKhDzHVs81oIpXLeK5rndqiBDFaH8A1YAs
55vgRxnxD8kVHfux8XWL/uQKrtP1WyQSm8lRBIvhcpt2o6QW270dn4IatF834e/VRqMJ17GeYj9l
iseBYcXLFrNE+vj4c0VG6YCG+hHnbTYSDlld0mh+Gvhl4pIBz9BZD3cCXq6BdLPMTIbwud1LevEC
6+oNDSXOTNW94u2om3dMH3kt/cpI1xqu1LuJghDXExXYGq8/ixCI3IuaIV3zMCGfSRTmYZPj4h7N
QTg5KLUmEpFZXcGOzijH2AU9iOmd2GNIy0Xb0dwx+wRWf0V76Fqhvr3wuS/Qt+WasHlUph9rSjyu
PdqYRaM5IbRAmkZk2VZGp2APZs461j9dirDferXlkbYov0snZrTB2fdG/x4VV+W/3zTaHCIhJXBU
v7hk6cZRr2JBzUtAT6HfPcnpXYocoD2ycVCP6bc42y31UKM0OFqYQ75n6bOOhgQOpJLXgdNawNw6
ZXcBhJi1ZFSTZQm/xeqvFvwBP5DBKQVas/y6zRhOkk8EV4C2bbDPeGgc8K5ZQkeYNjZXgEhwLenV
rs9jNsBJZ0WDzr3tZfvdU7b5fMyT3XrIDnhGxfFd/a4mm2AZaGtm7WOcIT5FuR3S+JGcgGCMhOKW
1Xhj/GVXvDVmrnLNtY6Jae64t/Qzjl+XsDLZikVoyamuBYbgNYCtGvD+82g4+ozocw0G8B/shiNT
hj0En14mSxGmDUpN5RQRbWko/Vg9LOFxsuefImFOVXr7fVqiLzfa/8Z1fD47goLwaNgu8P6p30LZ
zvPOZoL4CcFgXLeE0CDYbniIp1qPLSpObbjcxzKxHI5HlxS9Nic4AvVuvN96nhe8iyp4QRycRlRD
Fz8Vvy3l/Q71Obum/pZkGK1gQ9JBCXB5mzuNT8RBnGsKNopxwm5LovxJgjEaJ7fyA2q3hL9Kd91H
zBqn5WFVJujRvvEHwxfMPU448QVjgWU+YBlUz4zLF2ixH9jiXItq6+DbDOriTnOPkQjSPZ5nzsGZ
ByrTvHYNpU+UUOaJT22kF2EVFTj2fBiGRSM/1B+8ZLegJRGK141eShIN0O5Ttij7Mrao2+ergKUv
tVOmiJFtqsoUii+F++AdKzzRe+XYbvd14x4/XjYQoB4sh0hXeBKKsRuJOBlIhrQOHgEn9ZWJF0Tq
4FhpEZaADAyjLbSaeQN0pGdPnWPAXjva3Yb+IQPMXfrv8pALxYN9Hj5w4LCKXbBxr46fX/cZM7GE
TfQVaYhi4LzRzSMb4E19kCAR3wMOzFfRBy9bNmvovOamuRHES2ivr1A4+ZbIwnpPS6K618eyW+t+
PzMz3046sceKL0F/LMvnoEhjcsQTRVJggJtxGM8N9QpWr6ysKJYDg9cx8mIcjWhmBw4WUVJp67rD
qx62v7LpP9wxCWRGeoeYY1+L7FjyOkH0KN/0mDTxqfmWWjDmlupSfWtbkKA4KB4kRXP+1uW+hmWC
G2ZZ7WnX+Q0IPWTbRkKJJmifm9LseqySUYLqViqb1nnPLs9vtkqhTQalDSJwN7GxbVAD+sodeB7k
7AwjjNFXlVL+sY7fmKvX1QlXxT04mOftlmuiTzCI0EsxPTJn5iaVGeQDPMsO179tGDf0ZPXWTP/W
oHyPcpiFG7zvZtwTeEIJ0zdymihX+SwP5GrU+J58egg7Uw0y28hW4+A8dDWbgBquH7HmbL1EXx5S
rCyMWM35wveNFZgTTtSnE5ytKet00wv+yLEvtZ7chci7iqjRZ4NHkgqkGRBAQW586QqnySy5eWTR
6Saha3QFs2WeF5v2Rea7Pd0W7d5jcMOztZcb2wl3nnJE9g1fFvRtzToPitJnjIKxjOBSXVSo6F31
PlIrl7VBWvY71drCl0NrZAnLQYa7k1SiPNeAflaZhDmfZ09d6ZqjxaYh5EdwemV3fgzKifUYjwG2
cL6SZPecQMPGoTH3CUP7+OijozJf7NcndNxBMDSl8f2jhtvVZ6FoD0Ebmv+cbNReYoaOQEjriNWc
oFCaFU8qIKXnK7JruVTD58jFRvCa+gxUEKPSzkLSgC9oJHbnYcNWue5tMsVb3twStIARevWGcad/
wAM4BLJ3eaP/U5orfji8Lg0wONED8BiJGfh8OJrd2UrJj8HWmYHsrrdhLCBwR0QWchHtiIgeqPe3
k3TXmy/uDuRMM727J5ocXsSP3kuzPwN0a3NnaK991U1St5cykameNCY1N2Lch1hGnjUahQ+6r/mz
IiQr/bK6YNY+58X9odLLWZoybLdEPR7EQ2HnQ51OQSVzyZwY9Q3HcshxsA73vWdQCCJQtuQ4udGc
2G+XXAVmm4kVl8eIO4Uv5hKVVZXOZHtD31AnMUcmM1i7ZJvILilOqkzlTmqnBGbkPkq2M/nxPXtF
wjFZdIGO08y24eLvPKEUjAqqM11z1bV7+94JbU+pnU2AO5InRsnEkdmC5G7thQp+4n37/yLkrBje
lQs1dh6O/1By5hMUTHpHmYSAMfKmCN2iA01b6ynnDhD/RmkTpHdIuvzsdMszH96INRNR+xddET6A
2rMkYmqT7hgAWxGuagtA0/OpX9ed6sFhuBIUSrl36KymE9oR0/Mi9MkNnspaRRIuKETIqM9Nb/0s
0+WIwtMObjWc0x5QFbO7sC9eMLQHBLGGgSrkxWNNgZxifncTABI0gQozcWLPcGBfUhHeL+iufwmx
QUBuTwlb2KmNYZ+34NZYUPdvSmapsLGEdntDjAvNHzah/yea0r7LDVjQLmqLJV7dYz5BfFBby5BB
ObtKfHCrANgwqsMRCf8vZDE9uYflWYJQi1mAdF2rHyEkOfB5uLOMsOJwX+6/OIxE4PryAtEgLQZk
DhOnyWsqVwDdVSRM54fgeFxWfLZIAhOYhh73BMPn5dzv9vXo3AeW11pcPegmc5pvsAm+vOLa44d3
UXt+hMh6eeg1xKEinzIQXthK/n8uDuhx31oCnPUpVKEPxHeLvf3qmUqF20SvmClKQFDLcX84HO+1
8ahV20JRpTHs/D7Y8PLmBRFy2F5AY99FtihYy77F4RDe6vRDxb7He3eroAfVSEFmDrZraJ/FaPKu
BHTvesQoBW+UTbb19pldMy7GDrwEIcYOKt/1JpIVqkxaOQUZATDp5euIo/Qkn3bv5dTa8IGTdHqy
t5GNASWv6pNuQh5KyLY6K3IdzeqN/eZ+TJ1L+hQybdgNp4EjZc8DUAJbHfsDzJYJAb5j0TWzf4rL
agBDFKc1TWCOp4g5/M1UGHCcxUc98SZ6XnTp33vkwx4yXHuv+TWkkJWQEokyBnZN3Lhmy9cDk5W/
AaKo30gLkCAce4eeELNR77RUft8VgO0Ey3hksSNY3MXTMKFpGZNXak8G46dWVR2y4zQ0MLihZ0J0
dgF0TpeJE/VntE2vYULOorq8NiLgovMwAWrR5uYN63IYzAF0aTBQ1POikXTP7dqtxb1ye2zPQMXZ
3YeutxPbXCvRf1HhlzNtn8/0cdVoxj4ttcfqTAWkMgDrrl1rr2epIHxqrbhZsaL1ivp2rKTNq2Hx
VRFElzmZiV405GTQCIaazfpeJKvgPgmOhLencMsnRL4RpgTtX5ItIAVkrjt9yyKC178E/LmmcKds
0dugpScVo/zgjwaZ5FjAyFRPhaWuRg9excI1jgem5gjD7JYX5gpvV8C9AnM+gD3d4X4OfIBcNtXK
y32hY0+lKKcCVU9zl6m8JpajAyrbWdSGBWERTi8tlfRp5Z2DiKffEvA6LnaXibuBx15fU7Cb5psn
/5KLK+d73uIYM42izp3QhWtxtOZnWup+h1XiNX+vzseYsMnr+RCiTC7XYEP169H/Vo2V/nTLhSek
zROiE8RC1YgpPqZ4CLNYay8NnJpKZx2Oy2GWzT4uiYdngRama+CS7WZenfCRH6GBjhyzfUwJgUUh
bl5ekwbGEtIZuuXrgYrqUmkHZeeZP+vdE+E5+Hwpjg+5JZgVDci84fneAqZ5KI30njUcKCcCAUFK
++av6/5WoTnBYyDH51CLsjWSm1vHuCQqMPV69Ue4AZHfJuGhKN0pGE31tRbyis15c9VtZoEX+Te9
GnH9B3jdgfCKWkLsGl2ic7Kfna7gJa7vFCluJiwy4AQWIXoxxHVzvYqC8FVn+dfgzrrihp0b48L1
pdUUxz4OCf8zuGajSbR3buUGxneXn7N61ze5uPP4gHyxPuNdJaHxKpD8aJrpbwigxsJAKHBftSO8
mxuK6T4ZrSALxgzfdjS78ZbuJi/0H2K2oUc+CnscGTFj0d6prfpltZdxC1RnIQR7w8bfZ/YNVQmD
haOfC+cFh+JbMXQsF4M1Aiq8ycAp/L1xN37zeerGStMwqZYIfm+o23UUtqOvCt3n7jgfqRdIxoxC
c1WqYSdRcHsxiuQQu73Cbo3K81Jd+A4TtHxfLFSzSoMor1xwp7k2fGwAGoUev00+GBlcRUrfX3xA
quVog1BvEtRVTVcEJ+DXmjaWeOYnblEq/93uHxkswWObBY0eX8uPlZ2HfpHtZ8mhuXoBcv8lZSpG
qD1X5pCFSkTDdNVVFI4sDXGX9FAXvfmDD+fBzx1pfiRaOSHS6YXwlYdkTpXjc5M9jEFFUkIXrOI8
xUv8ajz2PIu9j6aLeCM1GNoXA4nxojb3fLpdKdLyQJjSJ1aTic+9glnCelDcj+nn2ddtIdqp2dfr
S/OkhKJSPR+iJ/qdTPaWx0WCggQbL5TMTi4eruKe6Js7opcToeQnL93hzq6UozeAlWhYk4DJi1ya
rhf34hFhsUPD/LMgloKBF/r3xp02AWHvFj50iiUGcRcI1ywKKHN8npjZHGdApZxv1mqP8ZPTAmRl
rwUOByQL
`protect end_protected
