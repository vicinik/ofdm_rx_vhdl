-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Evp2yMen+eyvIfGdDRgBDOOUTtF1dR6oVRhCgvAFY05ucmY4kq7drZcbgi2unILWX2tyN4j5Squ2
B8LUoHhu7qwYYlht3CiI08QjlzbdkFfd7ObigCSz/SCMoyarL2INmHvKm81T/NNq7fyizZRj0Pj/
yfQ8PwtbwR9Ccl47mbMPxy94ZbVb6XykYMfYCNnUpXbHuZcGP33kdanRpfOrOcaxmtU6sb/9ieRo
BnpQnnUNMDVOGCGnYP6mPanVdW9dVnacrn1iC+18VxvX+PNHowO2NY604004PSkQxo7lqCxhuFK/
OcqrLC+Hejk8japLW+Hb8GIjXGVl3i/29mO1zQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51088)
`protect data_block
knhBIWdDjy0t3tba8cINnl8ptqftzmo063PZ+qcy1iMP7UHE2xAmR0seETQYXgpEhmorzyXpVc6T
8db9Ra4G+zhWLHHJDM3wOg4hKbNiyIdKRn31VmfHT/V4RnrDFPp6bKMCaxBr+n2wUDG6mfqYWf62
uqrJOIwrayuOEPy/zO1Cj2G2dy4FIfq2OmXWgDmYnLdi9flPcQ+hpsG9dw/3262LNuu3ke3S/BNa
VtCbglDT2J3c8cFPwNQEU9VLjGu72yqzwkLBn71FGsEZzegH3ROw87cWFn4NrGcVNogr+a8JTrtW
kp8QS8QgjKlPpEP2fmEjn1SlS8TVbTWXZa61CD25vWU3G5qXOOQK9bIa0icRb3Qv1q+SH8hhaev0
oFl54AtTloWL59Z9qpJvkLRIU2F4NYPmOV4jwtAg9y8O0wmk4tGztS1W7AYQKTJEd24nxZp1G0RR
sKGoVd/DDoIuD9FFowOOOO5pCGmLL/it5pzFnIZ8P9OAyFWlu5oW+ohFweA/HnLolpX+s+rNCnU2
dchPC3D1iqUIMu55M+2vz6QP5dfBY8VgpUs/0dST5PclIo8HpxecBx6cE0L1lG8MqBHtLBCbr9wl
9eoBt8QaEv/3awk1FCq0mjuDMKPUSt+YDBMAtin0quMJf7UKM1c7RwSCjLYudNZDjqzu9cusPK9O
vLEpbT0JGQG+87MTfoqKwZBwg71oAOa3V07vcrondCXufv/HlPTzyu0wXImTK4s8HMS0O8gH61tR
+ZKT4RhhYSoKWi8Bf6ESitLbnDCFOQrlcFPZrpKg8I/yJ0w5IYfDuUNb3Lcky+PMpMcGpDkaZkHv
b9d0xPS9vuwyaanxHbEBakEHQY7fy/CJTG4jphHMUhrpogZcvvEd/8bQ6MzCEtC/KwoS4Ny6pTqJ
RsHbOM6edv/Uh6at9X/tcf1gzuDGSmquwLcmCDMOcOE9nABpOMMbi7P1aKhqYQiKEmDbBU0V65nU
9Qn5kLDG2q763EKaNX1FONbGLjHZGt8GgLNT0RN7hyboiLzf/wNHaZjQCHSZchrxsuWU88VzPiTB
Mg/qgvFzjFWYNJXKukQ71xc7jAfD6iTL5w6N/JTJJ82HTtkZB+6v2okM6g53ypBNDUD23WFHvmcY
BpVvQ57BXCp7QZ3H90YglV0g9g9JlLDgRNqxH87ZrL0YSK/tA6WpPKOV/PglW5tM4KyTFxPt/Hun
EjGRRKoMP9S5LllMYciudl6gCbLJ8XmWrj/B55uRilg3KJ3uEOc+7MeHnqIkyOqF44mBGqQJiob0
uFtKjWHKQK0vlvDYCkWHxy9UosWGvsxeecydlSFyxdZUcXQaJa84/xpDrXRoucTIKqaZWuOVWBci
5sXVzLk1gw03Om89NrZQOUIrjGKB1l9FCI6V6Tioj/I4/yaUcs4qH2YWfEWIN3y5mnAUhhy+WHeZ
dRU8Vo8+ljGxCLZ714PzyXmAxyVuI4ffUZpKAdQAGfdtw0O5IuZvMOV27CTKoilZfX6pYyK/3/me
tyJdd01AYEZT+VBlPOjyh9BVRembWaSssUpRxqQ68TOiOVdU84NF0y9rSIdYyr6F7AXcWAbZd9r6
VW+zUGn5dsoROBq7PIxtR0fMZvDyOyg2DWxNQzASSzKnIYNEfhJ6UdsEcSqdQZ+sOcNuuXFKAnfl
seBQTwBgayO8efJy8DdECVLgdS+qT3eCEDyyPH2xAahaMdxUw6DNgVSuOh9kCNd1SF/P91G70gsb
GJapb/JRAgzSg544Qsj7Ft2W45BD3HXS7RaqgLFCsZcu7INYcGjgciJ9slid5kmU/RfgBjlOrY2n
csSKK0YDqeKO8C29TIpCNAEAKApsptsQ8/Y5dShAy97b+ALJxG1osjM0rOOeATbzFcrn+gIwq7ok
2OArZJzwCZFC0PI7iqrFBlVvKnDjCMpZfdJu6Ej0bmTI1cnMrwNtqwp258qtS4aCfdj3qJQneVGQ
dp2Xw5SqiPpJjogqD5mfwldEsnSbfolkrSxUBa7kdPHGPp8+iBJgsJASzuqTe5D5F6UbTYfjbYOb
yLbbZifaxoRlyIH/6OQ5P4TRxI40dPiNH3knJELZUC5HV/h2tmHkqL+Y+AsTsBl/v7IF5158KCQW
06UpSqPfOqyrvCEtGfe5KBgNkxpvyoSCXgNGjlyMd10dkVIJREdgTSnt3lDXWduyXhl80jTYPAXB
EhBJkUML6afnvytm7X/GjQ9e8pVOOkxmSXSbzFGhIT+ltmVyT1iUm55thoSdvS76JECm6bxWx5JT
3ei1UCw4bQlYsMJ3n9S1fE4RHWTAuqEXE74cat9ZSXO0zqLUajXlbIOogLZb7pYG1NcpCsE5jUq1
L6WndjD/edc5kWg12AZn3jq/nPddp1mjsgLp1HxgRYiPNnguTx68tV+DS7FZvNwP2L8UIHYkK7qP
dlm/1xw45s02kwXWCl3H5XqWapKESrvHubKpxkqa3KDlJwUSKMfltGDIEfLU8L5LzXEc6lQeJA5S
RzhlsWm30KZCkMOl/cVlSk+ut+5xD8qcI7FnOZ437jUZsgJY+LMcTOnhTrc+rNx0GuEsN8poghEY
/Gu0CR9qYSHTAbZB3OmJmaxX5p62KzbI3OZpQlyA/U5TpNiToFtOF1nbv38JdUQ0+iWtdKcLN5hj
QxSbUSZpE7BZeMY9yF/idOUQiBpv0pPw3BBJmpBH7g2CgI2xwwS7MJugD0VF3tCejXmVUKLnGQ+w
grVRuwmdQUwPiQpRTgsonf8ei0tUoKWH4uLUcEOPILY4oQjLlWTvUpNREjrGw/rlTwGyzX0j7bMX
FgYMFjcAnE0HLBMTFiRj5K1IIL1NDYwCEgM8xjwtQCnB1wm12MBOdnrjDhLNhG+vcDnY6qatNOSq
nMaQdOahtKCbqPQuFZnUvmBVL9fbHpbL+ixSy4lXAysii2AnI5Luu9qcGLscTm6Omm1k0DsHpH51
FqTp1dglVgvmR46JALYymN6j+X/FkM8sxt0UcI2S3sUbi+1cayAHfOIrENL+SYUVxQZwvusNR+vN
mglvHXdmljRMxPP/QnhFV0fntD3zwex8GuJhDQ9Lf3WvX1kmld2ryDLxlipx7/cKf9h+xpYhmX3A
iHVy7w91rE+kNyhii6W5LPiWh45Bx0VGUF6L+NJH+mzTX+oPKZfW0oIjYNtDZ9+PFnetF5fYeHao
HaY1W4WC8DFXxQ7/L8vEi/lvd7Dce8IRu70olgXVuVxd2xxn589gcfLCryRIAAncYjMuayzXbI2b
CZ2WNJOKEeXjWFL9GLVBtCA1WF3bNM+Sqm160A++fsdH0JM80rLmxqz9ajs/3RBgglY+6AbRJOAG
QdO5Z4NXE0WNkueroSgHoS7QGpM+z/F6yvU/Q2scLS54h7GWwzK5bJalZEYCzFdzxGzhQSMywKEU
bwO3Uks8638ZeU3QH39Mh6WM8TUUUmaYqSo4MoERtw1eBGfi7Y0lS3nZr+ztCKkFaxYWllO94PeS
GlEFf1DAgWji/j+o7ImYDAkrhGoHsI90cT56+w8Kallo6VWzPaO7yBy3L0/kblIMtpJHkL0H1auC
0/qmUcyQ9rDxlQEeH+uHPTRLfG7QfOG5p0NwRe2gifA6YMeuBY3cBxEC5THwc3nKL0W6mZ+3UM+W
aZfPomzQ/+f1a9Cl0zGmc9HUElqzDyUrjdNvx4GV+fJo2DOwKtxSQdJ9Fod5EursZrgFe8luzPij
fMQGhGuVTwOjRqSI4RnknImf8F9+RGWNksJVShJpzHY36Pxsb8dgurgjbFgnQG1cVgn09m1pOZfm
pntZsPmk2cXGXFFK21z+zeBP54f0J2zIiE+FT1c3TpHFKNSXnZtVEVKauFtkqcsKMSQtoEp1/j5r
pQP6726hXbuOSDhsm/9lNpLkR6RH2cVITpDM3IJrOJPw59VM69eIVjqrfAI3JVqmpOa6MLcm4DHq
kRtVsre8xhYxTQ1ndGNadbbpIeqakc7zKkHyYT0WAyD7J3uT2lFuO0K5ev7Hjw944Y02z8vMSbLR
v+5ARC80q1PrEyWzRLRkUOpLy3QrAdTgnOr+dQQFsoBVVWPGTmNBoSlF8GeYqDWzFWTUjbu9djSI
kGo7sCz76X747U4z/n+oS6MQmIod/x9UH2mFvN5JCencRY3IaxfFN2+LldJ+EemXvHX7bhgmXuYO
9jrunqPeytgXI2mQp9a0in8iQ3NAX4QLQLXLcjByFei7e3mcVeu+t4Xe8rbev8MaSsJ7krQn4xtk
auqFayA64GrI+3xXmc3xY3obCv6yrbHRKsMxzPnXHHMAs2nl9Tk3IxxxnWrY4zjcvpoetrgSwqaz
tSpFwVERffypwOihIHLvzv4kcYmzFrkQDRLsPPxL8UgSnN51I6j3giiubYcxBmukFuRhTQv/4uWp
fbQPVgOqYZ04o7hHbi2tf2lSBOTXE0MMqIVo2vrUyCWUnc2PzUciBKERLAky+sDhVC+1YBJ6+BdI
YbSVg+2v0TLDfkhOAr4Xbv0aPs3xq5AwHoPMnm9ms64k9wBbmX+1QR43HQjOK9bITgxkA+bwmRAk
Wwj8qI2YB8QTfO6/+hsr2q1wsNelBLVBsfE4im1mmWPsPx8nSfiawTWlP/ijxU3XnMW0pulzHuRa
7ONL06ZNZc/0KLCqBs0yhB3Cd/J0LiStDDnqfQeCa7FM1Qm3154Yc5QzR1xKryH9yB9T7r12/fyk
a52U+PdxSQG7kdDGuYPQXzhxV6g2XF7gB4MzNVLX1flIEm6FaRhWu5mmq7R6HA6CY5VdyFgBH0vP
Saza1jtFODMNignE898p1bz/NS3maU9GObuEbWxQRyDNcXuO8CJzkXQG4q0fbqMd2N/wYGtXCyT+
tr4d00anvXF5HI7RKnM9tAlhPnFgNne1q43SpyUvXP1XS7aHutAl4s50V75OcMjkAqfDlnRHgmYT
Wfw1CbsW18FhM9YbhHMszhXNLOXObM7Q4oi5G5GaEbh3N0djTnmwJsq3Edw0U+MBnP1YW/LPxAlr
lU80BQCsXO+CedjoxV5dSwhL4JHSX8t0bZVhKb23XRVlTSs4AXmfEvHka87bNkFlr0sLI2pYA1Ez
iYkd8mLMg/h1HhUgAmp0zsCl/mDLpQPCaRS6LtXiYSLF/f6NKxckQdXAf64fZ2n0mRAW0KHAwC8+
jIDuA60Ec2L1XIeUVW/djx5QfErg252+VhhUCdFxtcRdvc9/HaZq2cf+V8sR5PDPfs7O+puPBdjQ
dYoFF4U/NApEDTIfMxhHKdEN6ewhpyzAsUiJUBBwTcmX79eR4dLOfea3jcLgcLHrAXQ8JR1qIkm9
Y3b9XUpZrpH2eULavf4Ni1qCIgr3nGIjTKOx4l7HoosP7pTsBGi9xcXj9ao1KE28++TrfbrsjIS6
qqjtvOjDbUwkr2qb+v+4BIPV5kKMtUVgzAhM1jKrs6KXxQmglKWpZGNYV9BKUIaL8NiIl/ZzCV7Y
J8DS3770+7L44HbQMmtgE8h2qHvdIusQekHlqJYHgxAkyRAj/o9uh9xoanb5YghyWSKEih5urYFa
XpX0/8ELSNcqvwhfGhZwy3eS4yaXj+vVoGVBtFwrEHrdqPHf8vCsuYAqutK1QNvb9ewgXhLbYZQi
9syBFqRgO6BK35lhMmEXYcrNVqr4xcNCMUwKr4mh80+9vO/3zRwGXpVxFUV/6/zYqrepKb9TY6eU
2wTNBOehgUk3I72z+c7Y/qvMxWbSIAh+LSxHckQ301XvqVgkdfmbcoAYwL4nS7CCufPIOGzFDf7g
PqunxM/FLjXzKy9I9yV9g2kQHijvm+wlwPj+dnRcvfvBfenuqBxAiw3URV7lJRD1dpkfZBsFxXf6
R5aAw+/97YbFGmbhsw+J+DiUBC2xSrcAeC4fHE/N98ZWZv4mA5uXwxzl3/afGenbI+zyMRWJCRm2
pYsCv/yMkdDY96NQPS0/ZOra/jOhzLUTAAreYlmYDtqo5wKTcsA6eXDapjDLksWEaIcAkRI4qyVT
Oyfn6mHTkP7rpexZsV1hjkzAeQ4WEbIUebNerdgPqu9dcEyUB689x7uUPG9C0yjqLOxSUCF9kMSF
ejgsNPR5cR3WPv2RV4njCcG9r5uMC14HDSQ2NIhHCGaiUN3hXUbpm/StuRVD3KREbf6IFLjtYAcj
NAEaWLmiZcE9HlP/ERZyy4PF+sifU7iHBB70OhSbM9iNuasWUi4OEKNBNzDpegxn+TBlum5VEUD/
ctHS4envSvcgwxZPuRJzNV32jbFL8VucXLDvP17sjU1fV5A7DLfAjOmUU7wr6ywI7zBO7z2XWCHL
/AJ1YLg+I57OJoUWfUzdEKbdsmsDARlgR24EvjjMiBrRx5htJt1keFohUAUvk0staL/tqYynhcw3
eAklBgM/mehz148dUBoqP66Rd0Xic0pG8g6v/LeDJmBdoKyr+XENXc0WwyOQlcBSzuSsJOg1+ziz
Zyo7ciXDEkpGDPuc7nTw6UY+aLgogDCTL+YOXzpN9drREHl7fyKrlgHDb21PHuSSCOmkrEXdOqEH
6EYipchoDAKmc7jdf25wKXX0cnBKBMeq3eVae8I/UmtxQmTGk6rEQ9/Iza53KgyhvAO3UGgrdmvM
lgjE+bI98dCFfhy1X8thRL4dDvcvNQAMoZSuHei+L0YRwUVM1Xk+ch5LCVFv31TTrx09T3OcBrz4
awCSZ4Vd9ttznx799bi6ETmadnu57DgtvuXkA+v6meYTO4tDnOl1HW61NVvGsbRe1cGBzlfGg8F1
PswhidK2alrkwxl5r1gSMRjg7RNsnplRvbecPQr6g19EF/hvjzk1dOZ1OoGrebyj4WL3ftwaxofL
+OwnME5QnGmUZCCL7lPs76SeltNis5xN9zAFr6pPgAf2GdSePb29KllRw2tqQ+WOS/JicmTmt7nr
W5M0VeHRDleoNq1KdD0oT/DUdsWGV8o+Vc9Lsd1ZCnugG0nRpxgQ73OCRfKn5OHFOvqS0KzSeExm
ZOuehpZ6PadsJVomqnAh4zihofFURP9hLIILjbGdEvCUuwRHLHk+qZd8ioJFG+usirh8Q4tAdF1P
neJe0deUf677qWXftALesXwrma/JZaTHP0moIUQuB9+fmXDiOz5HEg8ae59JGkQTLL0XNGZvoGkm
TzOfwPA8xW+PudNlNVJdvkPROpTSjR7y+sb2Yevu39fqllBKDR1lTOM8nC4vLVH2xPxi3I3zGcVt
0MKF13yPMRHOC0yDWXRJHMqVekSmlYrdwGzgRlfYROS4jhoL6v8a0f+2dl4Q72VTE1g+PvUdh0NT
GiP8ewLvaSWiWSVkrp5jDyBeZcMvd4q9T5+WGnz56X7BKLfhwnvnczEI0nzHl088dsUsAIbkooS3
hrv1ZKX0mDfGZmeLTzdNb1XZYR4MEOA2gnXtmwJZSrWbwa9O0JZhfHFuHA7qh/GoXVYenu/F1hQK
/QhhrpobnWFpRIjg7H5rvHHRzdJdM3kF0apV7jIqKVszl4kAv0+m5bOwqwud0WRggRViadCLUznd
tV/xVzOnl5AyK+9D5ph4F+TY9eKDhXCZtobU5ppT4vBG4u7n8Fx6XGhl3IaQLqQjuFd0gDdPsED/
fOvAEVLxH46t97NaCWZiTFITJspo9wIfACJ+49gVTBMFRVuSMfFqAgo7sbXD2gAEvmv/sJGlig2A
1fxjgMJIv3+wc8w1Wn/95CsErLQMWzTyZhM0HJRswCSwYJ6eVUOCrtknysIT91c01gvu7fK8S7pC
MjCKou35Wyfc6fkbQyOjtw2WsK0Lp0c06wwfoL8/N2oRTTbJcIFedGpO4Q+5FULkvboquObGSbxM
WONzvFdAqlcqIiqmuT4Q9dng+BDAMwxJGg9SYeO56qvU8YUJIDLZKZlRiJZksHr51v451CiRDkWc
ABUdovUOwd8EE1gn4dJ+uwJ00yYWNt5s9FI6Ia/L34Cb3j9gFMBS2S1dnbppckZm4XoNOcFOWsRC
rzohILGxyDFGqlEVEozaE7wFV6xjNmS5p9rYDgRxbANM0M4LM4oHTx7hjko6AMJr24K74bUckU44
0xuYNAlhNmwOLSCGx0xD1Y/wYuiOy8ivENRqyxc76CAgnxPCHwX6B1MEVQ1sJOcgNAfs+931IKJs
9zMiu8V1AWiPC0HZuXOsBQARwmdHN3B+c2AomqtdHkW2/gjJmaR6i3eE+uJo6FZpqdfpwq/ZKMTf
s4f9VWiBc9J+TE1Xd56ZGliS9FrZ0ye/gIs0nuhm2Fjvew90mCGmayojeksOwSleYKOM6kv1VAOZ
yabpsh1MD3eXVeq826LZBEaSw14Q8JrEk4SdqpW1NkSSHJlSqLb3FpEt1cWLny/Wi7GqbAGJI04z
ti+DAZlV4jy29tZDA4Af/7q00xAl7KLT3HiQA/QvMrwlkjK70hXRP6M8BJnxR3sjmSLZ5LhB7ytH
R6GB+O3nS1zOO2bw3fjSbOiDaN4v17MnADoJXHSHLijPB/u0g2i3sZZxdZ69w07k06yTEy7SJVMg
3BaqtnzKE/CaX9YxSABCgj/r4hEdeUoamzRbc81yvjwVtZLSs4zyIl0n/ir+QcysZ5SUkFOp1xy/
Kl2Ojc8UNRPsMIivtVZxgrrapNRMRRSwcIw9dofGmsttPuaxqPWFsaoQy7XfJGOaEwhyGhOggqaz
xI6+v8etneUtm9YjSEvvrX+i4fNQdBI5MeIhRgf8YSL90VMPHqa8Mu13yflsFeTHGBTLmmKXEm21
YaVsb9iPt8fn63peORs2C8N7GgzPze4UehTg4yBk5NYqdEuZZSN2TpHr0iWcWrPWeJ7rNSdKJlg3
obK3qKJiT9JFT3P+b/AKcMFzpHSRSM17FX2XCIFzUnL01X7fH/1lTdN2rMfz6ePFNjXT9OmGcput
h7GTV+kN5BxOYbyg49acHSSd7oKcDrbsLYfZ6aqw5IgRaCuq6+HoSvdtn6AWcUrT45heEG+8/p0d
w6+6hMIjIil9QXF+gZtDZOXHnVMFClc2wbXq6DFbi5qx6b4Gip1M/TF/VUnJbnGmReKh7rx5D7Wv
Ght4z4O5Im8kAehFuYLu0whl8gxjl1PZb2rgFuynrMcHSnjiKSSTsnbRBXTTvU7u8581/ENV7Jqj
/apt7ULQW6YDTbWObfjCygpuN24BHzetiInr4KB2lpCdTRJsJ6meDZJuqNoscnK2xphgiC/zFjTf
1EDXkRDuN4oEUXPWJPlarUuq9E/PKLsgpwVjPWGUgUcKsoIE+KeX7XMlSDEnXu5sAfzH5yFYnj00
JOUhuEAoPHxCtme9wUxl55fbqhUjLAMys/f12qAUt1ffsZwlhVEjJw5hUcpvXjSWUrwapfkRn/ME
+K6aBkkY5RXCKsOyrzWjnQSb0+WDAu7Aaru3YqtGSONoogXRP036Ly0xy2QE9aD1nvQefI0cSFF6
R/k44WNbItWN/ABHRE1Gcagp8Wu1dzwFh8EJC1ZATWJvCR/y1OmqiyZ1IJ6YNuSxo51eV3WmU4vR
CXBiw6V0XyZU/Z8UU6RjcSV2ZsdyI882gHEGp9j8ENc0S3o99VbiLRyPBW5IC68NK0nFMayURdrN
iKJPqs7XORRvdTsI7Kt+9c/G1JgWopcESKeaysxB0mQScRr3SzcKH2C8ZT3kkTk3AcU1jj/UhLeS
EL8+uxvVcah715cnLt/FIcmm94AG+bZamZyGDIZ4ZdArtazETKnLJY+ADnhG6cGrdvv9OXHBuonA
QELfqLeI9lo06YUzFob30RD006lNw1rNlJ+FdWmH/H+yZUhB9VKCczCh3KWAbZir2QiLch+iprsJ
2IpD0mF/EDY2L8HMhMnSMDvcoy4m84+N4Ao+aiO++7uD38Ar4AAPA1afyYDYWr6vXDgl7fIfmSBF
qpq+q9f2+OP0+g9Rs+Xo0fw0Y84bE8jtbMWLH5FYebZHMPb5TxJE6+bHqsLmRO9dkeBZ1l/hUfW+
Q/z1L+NLPE997NUnrLxwiP0MubpV3jZkNVUopCnXuikKYLnUklz07qyNx8Jfm6lY2EHQvSYPlWPZ
3TxeSHGFx0UXjHlxn/Vra6gBR/QOoTEZThGTMUE4cpGPTy7+ZCftv4tzfrsJq7PEX96SN+QY3/mH
vH2NCEupJEHJgJ2ker9jgefMy9KC1SrsZYK3A0fxAcX8bxkeP6v+knwH9kPPO5/cczJJShklHoYd
MGvLcguZN9+1YJFrx3dLrtFfzNu2i4UStgbvvIkssCCPcfDR1yKoDOxvwoRRCS1NtKMGp4SXy9kx
tZJ/WEa56TSmwldr1J+mTmZ5mRQEw6vs8oUwSKMZ0sxQ1lLHINP+SBDk6xHZaOg05ZuDUh1VFHlK
4ILwD75uHhBdtmn03SuEx/bTdIEiepyUI/gA7rGzkchxCamnT9sbAxZCzX1Vj6R4q9FS/1yfONJu
CEAw1L9lvwsOosOvrDaKX0/8pxK/+y/RWK0fAEObyEW4hFJXOTI/7jx3axIMYZc8KCYF3QvXHu1c
9YlRXSzbGGc1wbSzvMSskMnquu0SEAUkdpDkjnT4eAu8pHJfh/SOYDxEdcYZzY4eU+d0ecWwfvy0
abfUInWXHYL29l0qiv1hYdv38atpGo6QIyIfx/xksdv7Dn+Ui/CDK9REGaHucX9jcI12vqjsW2KS
FtTeodY2W+CePx/B5jIgMhllJ/kgZ1/M192LNlB/ykKapcCtgfiVufM6f0GGGrujUFxO2ASQ7bbM
5RC8UHAm31b1/14dqWOGHC7zX2t0m8VLAkTwwwBAtt+2XzrY5yqE4j3EcUSyJzRCwkOgx//DNHJf
a874o78m658yfnKC/Tt3U8UXZjQmY/IRB4+SIgUzHZmqzb2AJ2BdmqqFnpJUYl3UvlLBAlQNTq5Z
u6V8+LxoeNZf14Ihd+Jg3DoNiFSIOERbAVclopRDOL4ll4rgRMACuhcdHc4zCSkQDUt7oHjZNYYm
4IFzk1i1CQBOCgxA+xC/PaxVOsfChin96wvoAtjtgQmukB75XLOHiKL4wiFkqHiRFl8mZ1/dCrBc
QVuV+0S3EP/tOPSy0hb3Bo+CkEnIgsmnqYGt0X7ahI2T1bRIeXOZ9I37tsktIqQAL3dELA0a5Tl8
eyzlWI+ze1DH/SlQD22QF+yUSpDjBn7hgvE29gTFYPph4zhf1Xu/AbwVTCve9mgo+Qj2WJmj/O0e
1iouieDj7CNRzlhPqPRwvdJWvv3tlC8l5nSX/hx1P5HSdqsa9eM/cDIrFIw81XKPa/yH9bXZRVv9
5L/atBbL8pstoLy6C6XF8+oFpEFtirV0DsuUWjY8e2UjaeRTtssa3U4ROKa4qbIBZdWCURAi4M1S
Q1UxaKxU9+pwfRZDB7LT7yfUmf/lYBW5JwJqAC1MXN/wpv0JH0EQDZnPJBaVqR+6LikzQiXMXlzb
rnhWQHxCOamZiRcZ5kB0CG8NhxC+cz91plAFuf8pOBL+B2vtDtfr1SELChirdszw/ceThQkuqvr5
Ew2jHMZ9Dpte7KWE5rqb977iEL84vLwOvNMbGqBqFDbm+V+0MlINfgUDfZoajEIcn9E323sHBQ38
nYlaUj+dNUe7RkZUbW+tKJdcEQux1Z1chhy5qJ5dZX+CqXy/eeruFTpyRA9hSSgCUNTzoa74JNu1
fbchvG4YjeIocQcIEe/zxSyjyZYI70ycI+NWbQfdN1xS1Fnax7evrC+0UHmowth1YFfyLRH3B+7Y
8MzI52B0dc0MVJIiVyzQp+DlZ0HxGuIBs+Ja2PfN0QumUGvtydR1i8q3ASo1NvhuTJC2YLOZSNCQ
WbXYTZi3QRea6CJLsoG4JLPIUsd9z+eunda57ocrTQmAvuLxEevUihr4T2jn/qe6agO6AucroaR5
Bx50N7XCbHkCT9EwxzRyCaPRP34aKkbNxVC/od61JELKVC9RLOvMSAhB54J9g+zM127h/OHQccfZ
+yP/E2AxTzv0bBjUGOqp1J/zx65WjyyUwXz9ZvRcSPKIDqBp1MNpaM1Ar6UErmr0Jakzr/s/pNuD
FdO7+0IjPViDJywPC3JTVSPXEiMvu/0X52VkIfH2jBIhqjqJA8njw1y0ayE0KYJ2PaKgnEYylQcJ
LILWmDWvDAgddLlB2Tu9ep8+KYs/GS+fUI6lPilFTczLQEBRxQ7jBcsE/LGyNZM7U5EMQiSkxm0L
CTANYhcHox4fxjxd1wqNJ3apB12lBZO01xbBBh7CVnZ5qIeruRjkzjFYlFhiyxBGvLi9Lz5oesor
zWJAPacbOMWfWFqezul8rfZFyLcnhCIcmN4T25bde+3J+GCplw0EiAU08i95Rk/oK6qmmqo7OF+u
7BJGy2dqyga9HRVJlxrAt2WsqK99ek1pQpiIZx0LO5NjrjEDRsRFT2btFrLWanPfhM1s3x4tQTmE
A2C75P3psyLEI+Vo576py2chmvlpYGw5Q+WOhyU6guSnwktIDECIsxc/V20ptm4mIt6051Lu7CO+
u/6/ga6fqrwPwTzErEBPl4QvPdObbjNAZLjmbXaHOfK46V61upyHlxeh0y96kQRtI5aGo6LzqQuB
4A169QtTswvW33pdj1P1PSHNtB1pQspUI8iSdVJTl8sYzlo+8Nq3jijGZlfThy6dlzpSxHDqJJb+
s17qEsb2iDl+7EUqvyUf0jAnHsTulzXmtcWLZIgxlU+JNkff4avijWKp3yeBbl661M7kmn8UXsIw
L7ITARfCrOp8w6rhEvwiiQB7aNh3SJt9xsHgLvGsmastJfdjXaynNZ8FKnlv/lQ9P4dhVUL2/G7I
pWtMyZ0+DI2sqg93D9BMcVSNFcw8W4GqTWgSFF0hkB9mk5qsBF67vFZwhK7WOMCS/gFepIYqq2q7
BFWxpuPOgqK5VfGTswRyb/keHgJCm6/oLmoiFMBZJgfexdWdVCWcwr3JnfFBP39pT7bgl1BxrYRx
cIVjp6T4oC4DaJ/tF2n/8vIiTfTSnF/fA/aet/jfzOmLjYKbNA+dDoNLMapoymVfczPR41pyUfYV
KMaiAlKh4BiRoKwxNzi18nE6gQxEUKsYfGqlNuKzX8Q/SjwTTaAVA7TIx1zkP+HHGL5GLkmYXUDf
U4xDKW7tShEx6fqkKhp2B2WS80BJD64DZ8eQ8tPcFexeZcfbWDipGsC/OPbQiIytrYha3SKBmNVJ
mBEFHaFR4LU3PpPiS2NZ6QlSxEecR5sfJuBGaelDHqTeDlUu5M5rZDQPr+0Jrp+bWsFVdammz79F
ekcrfBGj1+qEik0W8djwc90OXW6XtVNldMzlsnRsYqhg88LQ6K4coXB/J7homh6POQSVVxxoMjN/
IToCy0jCuepUolwQjsGTmlkonRe9SPBZ4X91svLvIphjRcz3ID0ZeJTQRnY2SsrmrSChfex6iTJI
+/1NehNx70I6It0BxjpYdDTLy8QNwFiHJX9Agj+xNpvyOGFMlz7LtpDoW0jqDMJjFRPKS+Am2RyL
ntToiUbsaR62JCFZrJ4Fl+SIPmZyFRxrZqbtsN6LOEQeDyGFSElt6BfwX16aWHFCG00koamf1MfO
fwEV1gKwxR5uNuA7ZVxxOMadwNsdFl2jwxhd73LmQE4sNtVjwYe8C/QT/S3yABuSpeNXfxkj2lZu
LJ1J4FVtPCjOcOEvKxiw1Y5McLrUvKjv3ATS71zAZ6B1EH1bLNtSMf5lLuWWgy6YIDl6hbK1xu3k
assARTac+lXzNPN/7LNAkLrMpXVA8q1x5Jzism5XAMozhuhSJ7brvnnBbuw9GMVb2fvMlOJuUQhv
3LElZO23Mthw0M+J/vVc+wSkMcnsLJeEr4BhY8vMfUoLxJC3JqHAKZZWikb+vLesKVWivSII02c1
OW2LPW1J8jCy7ECUolD+GXxGF0GQSojUX8UHQR6yBUI4tYCTnYk+B8pfoZJVsKTXBhbTVHzID1wL
15OgzokNsCJFkzHrr+qas9brQt+PustkZ/MunNfKBpDGx81X05I5vEK3B9MEqdeDqI5ocSbhKEix
YfHpiGASrqmh2qv7539ZJ+89fA0MxO1NS5pa9qBF45caqLlkdPsaZXETqy7DCPN1gHkZAlRv4nzn
8K0aKTpPnDmtTArd0+SwiNeXPXD1kfC9eeXCTa5z6LrP2kKqsZifZgwkLXTyxlnaX5keXaBqu6MP
wWwVpaz1TZy4jrOxQkMacbdykhd3sd7Pi/EVDCvO192Eb69sTdVD3MulxPDEw1t1hJjJI6xEik7J
307ba18ktZaOLnRlCbMSavPAlOOqclelbqTX9J+UVWOUu3p7SIU9zlyI7nJpaXPJMcEuHkqrkNBf
Kk7sMIj7rswkpouDO3HGYhu5zx+8+PcwaxYA8Lu4lnG67UjvF/iCosBun75+CXJZBe0whAEo81V8
jkOf7iaEykYsfe/8O2Xke0TtDM6ZViYUREPWpRZCxDQQpHEDRMzp6HUxp5dL6SocKyAckFoZ/DUJ
38d3NTl6yBppeVw0/AQGmz59f7241oS535Vmi/MYB/oVAJuNYbxdDBOExn6293kCPK5SYX+mwreQ
1BOmzhJmdjGc0hmSKOzuC+ycd95osVsqbSTMT+Vo7INnVwicRvn0xySjc+VOAmgGOa0rdqE6DDqU
5niaSYw9zBS0ZFIBBA1k8MvxE+0Xls8vfTnPdYJFQchpy7edut1gxwaTgkdaRy+Pq8p1Mws1wPAC
LJmI6Y9ZTvSacxU0yi6FdphM0vwpFANs1oFR/W03Mna936B6yrF2snYh6DrQLvNqfxDHw60/EAgk
kvhk+x6sUYA81ZiQFcNdPkeeVBOZgF+h5weLPxIthf/J2xUD+6xmBg8XF2O+d33eqELSWQrsPjJS
5+Cvz/0kcdKWft0X8ObbHqnCboQDn5jWNZRw0QYlU4F612/gRjEWH1n/rlxtiluQk7A/buYtHcR4
BYyB+LEL8QV2sKyo2Xz47SOhEZ4ZGcqDUnbyGeCfp+wKaPSzKQmD44oYHSODktBKdfWYa5mRgE2l
oThrnReXHn5x3AdS14UW4jysu6xHIWIFC0BJD7j71CvjFDhvaVq6j+63MxJAjmW3tLn2pJUSR8bj
PXV9x/6IGbfthIwxX5zCqUYDSF8wVFFAYKeXYU4QmhAHbpH6537zQD5kLSR3UUCk02hqNv3ItSp5
+96L/cnFFahu/rPMRMig9HZ3TY9pj7jvj5vof9D3GQ0KSlSL2k/3A2uSIWhLEfeVOXYXbyXqwYH4
MBL6/PcmH5UAqc2ekqZMu34g26alIihs0sc3GTh1QvlcykHytpf1/OwFw3m3FjiXNIRbr/lFbyr8
sC6/fEjGk8slyMglzL1IHIFSdAbuz5czTvQvcNbosVIdC5WIAspM/aTWne4kUqDsOlfzVvYzxIez
MosMxpeuVzloO0KmUBoMqzRh8fLBFb3aPN7DqfNMFrKECV3sAHP5/aCzRQz/PkDm1y1cgn5njoMy
OBh3pL3v5UzGwFosAXmfeFB61sHfHZN+DioeAqVJ+CevKn6zWC/meZjkWGM6GRJQ7v7vGtnhTCHm
V74hI/GGbeYz8bJ5Rrx6Od0iVVVgAborEftPfEA6MUIUoSuLOP09GcsezobisL8YuMUuxT37qIr3
IUm5+VPzGcmO+3vaTx/+IH6+1Z5Wbjt6+ln4gLmKQkJowywnBn3LaT5DmALLCgR3lMP8pr4CrhO3
i/5DLx5wYzf/Bokzki5rTIvbv+26ADEzUif8/gSN2uwJ+Pdimwfd1p+7LwWSUaACOZaGM+aUHROK
f81J8bR7qkNFK1/4aBEt8pWsPTJ3QQ4Rii9VGGiA8vnA235mjcVutm/ebpZzVFerpCZL17a/m67Z
VIAM+uVirj4OPckcIyCpS3cX5snsD+ZcdYvlHyjedSHU+at0+hpvfr11sT8NwHSITEYrxKstO+Bo
oh3GkH60lh56OXTRuxWNp3+ZPeRD0wU6nFR4wOcJDaMjSZYZ7zvFcVCxL2eHXuWWLgXX506HYzP6
1ySxooBOxMeOUsELO4rbR7XqeK+6LkD+D8k1J7/cLMixz1ATouqd0A2MfeQS1mZSVLH/ZInyU2m0
+Q8tBmd2IJ3U2Xhc1xueufS0xTBsF/8pCVcCl87GIE03xXaIcbJaSKNoQdiRBhGtaiNSjtPIKbGd
6ly9yNJkWALjEf+Kf06Agw9D+c26qPh7aaX2wCYB3IsHIM2IqQIyu/8nW+Jp+7TZF4ImVh/SpC2E
suvchOWMLScx27tVcEQ8ym/nTjR1W0h9OVkaGqjod/iIMyjtNgO4CUwisbmIfRDchF84Cbw3qrDQ
PqiWc9xWry/K4kMLV7sEMK/rvW7lhB8o4ll/qz7v2UwBQPAEkmIYR9PvgmuLBxSb/n8d3viP1YfN
6UHq//741kcIO8kTQnRNWhhmt1m2hSGjxjdb/FptO/WIkJqxiMlFqsUWsUgZFZ5Hrxo79adQelVG
QiFUqVGevriK45A8wllJkE4ZupRjI0hUavC8hfrRjxeC/eMY50dcxCsMsR608uFIqEu4z4AsSCh7
8WcVBIhSX+2WDJzXHqY+UgzSTjjQdkEQzHTMij4MI25S7588IEv+s+oiTNPORjcoprOLdQ5eUd/H
kGW+WeDxK+2cY8fxXwms/DOJpPBa93085Tma+kX9vB9QR54x/pk2uSorrng28E9klUP0QlH8WK/C
xtff17sprDOTZb188ddT0bBjGPcgplxi+fXURtcp8nFEADzSM5Tr0vR7JZz7v0oVioRQGRppDRZc
iqLxS5mbvqmXLj9Q32S5De0d3lA+ZOO2/ub9hAFniulZRe5D0pcrOapw/ED+gy1NnIPwEp/ec9HR
r8t1aIHhG8t6iUguuEHNd/U22tSzDmY8Hvz0EawO7NVjwzL1sm/FLbmLhxeXn1ekL4LTMQwGniZ+
yXkYZ+TQpTL08fUJ3lnur8aBxWpOu6Sw/IoSFkOUOGc+laBMSkcDi8Y52TiugCTpgnr34o93AgUl
hYGj/MtQfZnpqcTSCIUUzmdMvmK9CxN//b7XPcFVNubZAFHjsDUAnYV1j2ve5djsCiGJMQHTHXcj
Hl/csbCg7yYoQdV2NvK6Igw8FHXahbTdx5RyXiq0JTN3IyTGs++aqUFTRNu+YhScnEWSZBl3QZfs
AcXVriXBivtVDXAgYQfcHdskYe7Dknq/yQA8B8+b0NA4rXbchRsAdkhI08JgLAHJlDs10jAB8ipP
C2H5s9SGopetEQ2YMw10YcAh77m8P+G0b0j0un5uzWpyA+c5jQKGKoKJyfVRuqlcB3bJiotGhqMS
Jb7KfXkbZAdkShUkU5j/EkLxn8xr2mBodbdJOQEGqqkzx0EL3hM3ZzeQ6eHxXAQBH7XvZI5gNN0S
//3XHi/VsXQVFV9KCkcMShCpaUYEfd3LxydCQKzw9C0sJlBcIRSnBp58VG9kYR9pEslDD1Gt0c30
mo9g+GQPzsP/daVZ0OAx5Ugwq6yTwhImuUgJ5PMdfSkMZRIZWkmeEb1r865PbHZGelCg6iTDT37R
EnsKwKZp6xfhskws5dvQWzb599C+hBtmvbhtR0Q2SH2dXPyMgNqanoDmLFuUW4VlA7rjGEj5TXVK
vBtIVctlZk3epaKe4Nvv+oI12i1Bt8AEViDcaPpa2peLc+N6vq0i2SNOsw9kQjD/5mO7c0DTN7+J
f7R5+gOZQhHU2h8JnX9CuRXSP3UBE9/NZzY7ZPTgEIyG5QUkOhfgeWnkAy1Nh+6WZqO9ZTdkCydV
QJP6a2dwRczXI9J4lVV9lCaeyz/LqteEtL3wnR5F8md/auTheJjw0rcnqyTYqboqs2GReoReYuaC
lpbGRuDjTCJIpglQi6RJYNHWzrU91pEHXL3vB112q+io14EdTbQUYKWsqLXtGZSrjKa99YPL7XZo
ELHu0ys/ueXYRCVdiSmDDTMLvmk2fhBhI5WF/PTuYcvOSZ3EtX9qhCKGdAfLT1GnDUrfgWzJizpm
HTZarkK6x5Ew9G4DaaYV52wxWetYEY2WgalKKsXXwuKWjIjf49Rc5gsMdHzPrfSjzuDgmj+SZ1ia
PhhrjQjXdtXObdgkquvBesqyF0A4BTHPBPqIom8t6FH7KycZNT3QjB7GbWR0IujHFOiI2v5REEh1
pudsj/Sxwgyqlz2GZnnO+CvVW/g27AKpAOlmjsSDY0ghKELtIGxsjXMd9IHGVJkQL4jJWLU0R+K+
kLmsmndHEuQcFL3DhDiag4UwweHoudupcHb1/V6xtqtoGuSTzJtKoDRPDr+OV9wNUubSK3PIc6tl
tjcSFx4gTLfi/oa/xah9jWR8cTuN2V2Gjk9DxByZjoZomRP/6INblZeG0omus8eQxtVhKcDyqTmf
gRP3znrfLbcMo7ag4hNuevrZ0GWeeDO3RtMrLY5FhrqB/ridWr754UYryQHDL9NbQyKn4wA2vFuZ
lua++5hvNgLRzKKtn+7Xz3x9XRdxpQDelUU0w+fY12cNG349ilyvcNSAQog7XoI7ONuUb7SMFCvp
BELY8u6/dtVQu6eeCo21+WTLShEyAkpx8FFLGNSflbx6Dem3hNr4vp71Gv8gGS0V9cNRpqwm3YgE
cG1Jlc0nphA9FfnM+p33zD4vVyd8nfrKNc+lWoDRqonGqcAqaPXkhqPoCZ5PphxkzXXTwT9fNqef
CkNRTR4fTiSAY4AnaG27w1zOZ9bzObEkp6SZNBOT9ZkdQF4TupyWuUn2KQi0OIgEetJQuwFb2hSO
bGxZqQnI1GhP5oyvzfGHN6EGQXhN35l46L2uumw/2+2y98KPLVd6DT8D+fEpnhgf5EyDVb4cdnA8
0ol9J909o9Qt0fSeNwwPTJua4pptNNQa2S5RIlL7mlvHALViyzmGmZCV0/h8oviMKTOshGhGDMBv
heeSCPFpLF7qAWNXDpkztX53C1oOhnHffpikbucw4/Ak2xjz+atPaZt8g3ZcfL5w5GaIfKBj03Eo
ybeNbXTelPj1YPIIQTcx6p2QgIa7R5oZAh4IuXclA278f1XPWGGkeouX6T3+e2Tne1KFA3UD92Tu
rGS6lLQvkxffLjGGUFH0Hu4lh1LBbVx1+LnQGqNwI/D7+hXSSxiBIJOajv++tXNE3MSOaYtQcRHG
tI5hcvgmZOaxtnX5g2cFiRuDTaHhtwLWzR8Wl250dSbmeb/gpMljLFqravyFa0/WClxIYR17S0v2
eOMf3z3LA7o8aeat/fFbLsdmL40TkqMPOkesdzp8twL69FxQveJCfrmo0PAynTRnyc2C2h72IELK
WYuEb2PX5vEP8ya5W7SCj/QVVN3MM6EkaLiClv9F0QYU8TzqbJrOJqqIGtIgwuqvk+da1teFWkK3
YekAuyvpEqy3Qvf3rd7mv2RbrO0mt4FU/1c7O1ew/+Mo9nhnU3uzmgV3eXjmsBc52KJEQybsM1f+
A28/xNFDiV475PuIm5/ViZUXgDcmvcoefjEWMWOtwsDx0peLI5dWN5NAblGZOIV5EfTecuSjMKBh
wsv3wg5ybFRHD3ll78uu28CvcCFVwmXaNuVHZUS0G9L+FkUbE4yzuL1rDtO65u3/rNGfwk8zggk2
QE+cvKpSAM89U3ljFn3c1NXCMkg7UpJBJKrG72y/DQZiNrhUdixlL90XTubnLxV+VsmRdJbzBnoB
Mfb6DjZUw2cEFH5hCYfbNssr54m2fdaOCvAap+miakGqy9dRXgCDf3S1/KPXM2kEkWfwB9LJCUtW
PKEpUlsGqL7dFR9HZ9JAe6MjGh8hT5BQFpyzCdUiDSLO8/gEijKfjsypY9o3P3+bB5oFO+abwDXz
8OQ3HxY3gsgeuNYx4Y+PfW8C9stamwqwBwNeb0xuVRDizBiK3EEzc/SlfJBJgvfxZrYPEAy8g3LC
a3aUH3SPfpX7JF4K3/IIpFg4xoBUctGUc3/LVcMfG7D4XuTZdP/HarcD23LlZYigkW4DMSEQ3GET
SOumpUB7oOQ9vQCZyFp/Eg2EP01LltB0F6De03Jio3p5I2p3i+5v3SYwwCU7LOUtC2OFj7S2xuWH
HKI7Iq9u9Rv2EtcC6B91vVYmqJNSd8hghUSnbvFLQR5hZHW4/UY9OmCUbUPx3L1X8ljR4Kp5xwgR
OnrxVuv5VQ/rdZ6NuZchsYuRFbX6R22po3JbVr2sFr/jbeMdJ5f6VBv4LYlfZCYqAaK3BDX8MoVV
MQGlfwO8UnCCTBtOWHiULDJhlf+eczEmt6uHqGe7cx2H7N8N7Xa1YuSEIqLiqwccay0ALi1QC1CJ
rsua9dJ+M0SLWKBtaDKgGgswnaG7S3dr0Xrq+yZY51IntV3FCFLlya0N470ld4X3ZRxZK3wTqrgX
w/UC1XIJ/oJ7u5W9jue2Kf4+4LwLh1QTSgCvHTKAIlAuzqvKYQ+ZwqDTVqbvKqtUoEfzw+7A4gjg
vTyPrRk42xvErAsBrFhzqSTlOYUZRpSxxvIwSS6n7+7hBfDB/xpq4+cqSzi4gLs0ovns8dVhZZ+F
3VuSNo0n410sL1P7RsKR+EaBtIXZYKKv05VlvGH1yazADDbSU5bAtAkDV81HyJWChaHhIDxV5Dmu
Yf6MQR3GQY1ydrj5YhlQanDU/LZDTrOV8BHvxinx4nnNnArnWoalU4JnHBz9tp6bB8uIuRiaZYJV
54KMeVJLbjXt2j4mt7gKsywHlyCCcHjIgsHXuYP9kkFDFBGuztBA+naH6rC2sUtQXFciW+xqOxbn
vV+qdtBQRmnpAYds6TZiVNZKpPkJ06VFhuLvds6np7vqfAVCljk3S1KzhbpLUEzeQgnN2YpZKbrY
iebFZyPYdp8HMyI6ONDCcpWXEPw6V9AxmNChwGCDHZeyucB+79GvJi2k3K2jW1p1CiSsiITGvhIW
W8N2uUIgZGpsg8ZQ7d/dUzu3jFZfNbUwQUObaxBHt6FXcbxU+pY0oEiPLh0JnhsnKUbTfDFzMstL
IJwZHoYMoSi6T7vux5FPOYOKUMd9diXPMWIB1BxJYR/b9p4Hveu9IifsJGhG83JjPIx9hIqOagLe
mMQl4dDk31+XycqCoMEmSJ6BJ04zvrjsI376xnclE/j0D4y7xIDGlc5ce/v9tsl4ypO1s1fDBusR
CHw8RMDFBJW/I6rWYw157BTDPSG3buKbo/piWBfTtqHhoKWNg3tAyHnHNX7Kg5yvAkSFv3hIkXSF
QBEeOZGYPbU6TTrdLHvfbnLiASHY1qWzQ2rv06XoEKNz0e/IX1SvGAE/C8Di9zFhYClwfHCcHFFa
Gl/Hr0x0W9hzGO2xFwNWE0n8KkDR8EzTrcxjxAcr5sS67X7qIxLuV/1AUCMvwk/6nWM4tUHecXXs
1VgT/kNUwbC9/sAwIZ9cnX8xh9STweioJxFeBc+CzUS3h4g8UI5DMJ6+FTkUw0G7baEv87YsCrp9
7BWoy9z81vnrh5gnSEgZd4Agn6PrexAzZFvMuyH9qjT7EPhqZksBgmeZjwXlRH/DcIv49xY8J+2i
/9bi91sWBrpy7gUIraWhVtqFhtbF2DzezW4LzeSWTgulzxTYH0Y64lbKbPySyGxPfN9l+uoqzAt7
GNVe2rpbDnawWMLKiq3HYiUecoD0uTlwJ3DIASgGeRtixinMus78Xt56OMabnzDvg3MnEtFua5tF
r9kQXcwIe48TDk8g4Qyyyhn0DEbwfhNjwTXoR6SSxPsRY8vPpaD1OfQA2BcJWH2uWW4T7mf3BFFE
yLcds5mifP91lS9mde/ulB/zAE3Dpv4J28mWjEpEBxNTZHJjm3l/PM5wv0ATN2OwMfU/NeCOUqeg
AL85XGQ8wrX+sjrjWr45GeQDIXhNDvm9tLbljgaSNXtekjhQsSCDfFzpcacphuINgzcoc9xCLgUs
7zPboLwcoaM7Tp22a7YHLfNYvQJ0qg2rL3lgaWcpxBqTe4gJAnUePekCcj/DSanXfZbKWbimSeGV
hyt1fdOZiWw4F44+3RSaEnwmQoZut7zER8aNsbiY7jSAJN4Y+SfM84vHkXyGNubjzL2CNkI26PI3
GIrjBB+ohKacH7PfpTSh9TNvFkEPWvPcdE8QY7PLHcUQa6QD+jJS19QblmTmkrQERc4XbSoEKH/u
eMm11EMOoayA7R3gBA6Vrft5cWO4e2aPUV/vIFnuK3xYh6DaYxj0a/53wAdrC5its3AoO2QrGx/l
K/KjclkwMvYjTDjjpJV1jLswBNpZgmQMTM/BgpNrr+IFdDw8WoSizrviezqKq4BStnO7oyMB8Djd
2wOM9dZrikS5fqI+7xOrUo0OWlFXK2X1KrT/4h6L3jkunqQC93m0AAr7WmY33ROywjWHvhk8NOHw
kgrGEpaRWzgFr2IHhgCRQclVzrA7f3rPdIrDDmkKuaJsTPZ2pg54M6TEwhjsKpt1Qlirr2GqvN4H
jJROpbfb4+qblloxjDYW2iUOTUSGvL6IRIINOMcIstz4oqx0XQoupqe9aFTmEWi3UIU8ngh9LeAb
GfCOP/F4nI3WgeWru07AnqJsGOkmhYRxLXKRkBxg0hbQ8kvllgBzoC9UXJR3THjtmSfrHiMAo4/y
IbT1rn4pSto+Nuk8vbHSlVW3yLVYIfgKEHN3zoSjR07LRtU2E/1KUwxqaW9EUXkhLeM3XVqKTN8M
3jGYK+W4gQO019/tO/EY9AFo1SY95uZYx/Nal5LWdIXx1O1EK1ez6onMfrk2EuQ48g2kuSiJUjuq
2aE9Ouq3tLJF75pdT/kVyJZfaTABLVS69HmkHWROf7gYxE0xN/cbH6sEGLGRqMu0N5x71EE4jaBS
868jW6GQXZZzW9ElN4pc0s6OvQXlYNRDfAooYZK03Q3xvKeP9DqXsy+OHG2jnlz3lYu+9Ob0jouD
F0zrWkI0+bK0kLAFT5oMA1Ef41JK/5k8bjU7wrRIogs0nV9UJQ8DwcGjMQURStRTrtx9e85QIF4t
jak0/SWiXoDb2ewgsem1HAIUKdqnkyYtpg7elYiK49hd+Tw8A6uJnITVranV4T5Op+UURLmScxCn
h2QSD9/8avqaYjcDrgOw2CubgV8KEALJ78cQt537msHsmiu9EegkZe4x25oQD5sJQN0P43opDyQc
y5BZdBv6MmgRzD+vhTisVFuL0Y39HgiU0SPJ1APUESdP8UR62hFw5FhAHzm7m1yNeZvj0eZG94N3
4PXmiDwgSX5asciyGxiiAwAl5U483nwtayUQ5JkVaMcuFMIkQMKir7J0e2A6jxa0KaXsPILPwBp8
zzZ9GZ2pYByKwrtbiW+60R331hiWA0D9XTEcPW+AcAWQoe8pw0FZqn8b/P12Pv9h1sB3NUCei87r
H2BmsriVi2o8+p0TEyqk+TUY9McQCitdeUlOsAPceCEbIIGcjNjpQPCg9UswymOzmWSG2X0FDryH
uN8VYGLxKzwtRsVXV7WJPyJLGIA4tAq1yrW0Qr8aIBkjX9TeKS2OM7jU2j49XpjRU0SkdJmCBVZi
jOUnq4vryIE3gjLEti2yq7ID4EEumPSgKHBfYrKvbrGlqCO6IN/qCjdJbF0oYMDM+VetAtX8f9dP
2cO86pT4q/cwL/IWwnTNGfJ/YYL4K15sa86cWZDjoomMAY29geGj4HjIMHsyb74+FZFXX5THH76O
Z2kQODWDGR62uKIwsz7i+BXdRV8xQrQsGcPkriVTGQ0y+7X751YtxS3fNa1U+2QvS0aHe4oJYNtS
aOXogOUv+nAFxOW0MxePcQn0ABfcSpoPSwQJU7e/adzXFu2KMkccEPHw5m4uPnEGf+ua/aWe6McK
tJDTv1LqwDAXPFzJa8U/4Rj8JUFnpbMAanc8kqipcVbIxlYLjqK96aWTEq++1nQc4puo950PISKD
kvJsxuAO+/vAV2nAL8cqtOEvDwqRRkrcYodCP88yv/Lt6//xdhXw8qCJRuDYtxXmU+EjCKHEl+nJ
4Jc9TrlJHMCaMIbsMbx0UdSEC4BmFlafv2i/5ZZST8fxPLPcZBuihivuG5SXma4Pl1eLMEnqqmxD
ts9zxzzbIQopHoP8MJW7EkDjY49UINKE0zPlacs7vDmyU3c0QWkMxnUT/IMkTaBzkRv2lIrwZkTP
Unc7jDdrlIavOyyHVYxrgHEECcIZmf4k4gCpG3ek7Iz1Ix4MDn2TcfhRhTAYT0hIX1amZZ13Gqu1
BRBNYl2vEakLiDO3x+YkOnW3hts/xArUllFu1ztfF1ad0tvOfIzuhaF+1Ay7/MctPv1Ecmsknjoo
TQb+XVYwLxXEY1yrYJHCcEVBwrvBa2GLMXUhhuU5qrBMcGlQ/yyQEx3wz0eQyHBsZutVVN1t2vdD
o15en1CetT08y3mCRZPBmV/d0wfzY9zVXE8MwYcbSF/4NJ7R2+biBvqWd4Kd6xvw8nannEzlCXLE
uuLyTEG3JhCNcP7/TH9Ll3dxhfU3jcdKpUesLpgi+U2lm5qQM/puvGRVrytKfAIBmUh9iZUgcRvT
lvNaM7cOc6jumDOmS4/xzd0iBz7K7lJLVTz/lED+kU/L9cdLbAp5z7A7WhnuQmGBL7Jmqtmy3ii7
k83c2yTOPj+DVg1r0nxs3fbViuPvRa5eMx6XW/Z5QWRxWN9Bi83QDC00iTSQkLUUmEPskqMCOSNO
DYgAf23AyHi6oET0qdlRKw0eDfLmatsQIvrAScg36pBBcqtqTuRm/4bm5Y7sNYVs3XAfRoUatxSn
1gdxmKkPOzZ2F/Rl9B36b7jrTSbTB277yp+FUsGFhIFvUc+gCfldxo5mZYvKc4lRo/7kieqH8aLn
NcrXmpLWFLh5JsHzGQAHBvDMcyW9Po/M0nufnnmqaCICX807j72vZMBl6BYrIVCfLuBosb+okDHQ
/myiKpX2O214EU210szw0A655XjFAsrlrbQMQtDMmsEcpvApXWsV2elKcWGtOGY2Ri/06mbM5DF7
VJC31dP8T4D0eUWQhZ6f9itvo1jLKSU27uWKePgIsUswiWgpwbWS06lof1X740he9+56P3c8sw+s
qh41sXqxuxTKX1ZXdbvCp9Sn3icRSeg8mrRj3Zm1xBMkbVJmy81ANrrJ46k8RULGbEHMYyTxX2qC
90g3bGFEO8i0ejcsgXqffnW7UcXfyJc50RtRKhWGAw8yhBzUsCK58HUtRfoymeUXYHHoNOrbbgC7
wqDifqVnRT+VyurNhbD9cXA55GfU2JiQe473H63TzDQb++I93WzyujL6qD47wioSOO90LugaZl4R
OLtXNEOWXPDRDyN88YHkVSbftbL7gxe3xR2DSt1f4sw62DEpRkFhZ5M6ZZnCZlG1WJVmTnEevWk7
EMqoPqnMVuyobW9pKMtIS5f5uEO7+M41jal5w+DRqvTxU1BTbC1kGxFYQIwKqOdxeY3hifaVnVxV
gsXLaNKgJ/ZaIu++Urz2MQkinR3euODU0bcQLKEXvcxyoe5veoaMq+yxI8Nk/igkiXdm2GXq4SVu
pIKd2lUT0x4VaNDT7cULOKnzyziqtLMX89w8ouQv8gwA0ZyCmB7iPrlVq/HFJmQgG85tsr7Z7AMN
J7vlH0OD6FKTncwOAMM+A876dUepQ+3MUJm6joEuTCRJYK+OMiOCHuEr3s1WJCu/hutGSzcLlIpt
u11DN/DCflyTqVP9x66DHh0E80HoLLtgvd+qgGykq6pJA2WwIUWW3JfCHRf0/qcxHx4lUobQ9PA6
V6JzuI9UVXAmxmx//HfMDMxo9RqapLZrMEIir7wrNgmEhC39BCJBN9mHxjbHdzgsZkoDuGvVnIFa
GTXvl5hAtiOdQlJ+8/WgQ3gJ6l5gB2+vutoyAr7My6QtNpdEWpTZ40h5Fh8xEVFa3sP1DPQp+9Mp
frOr0G4uJGq99bbhE7Jd488956z5R1VVKa1SDCEo6891hDIqoPLMna9SAK/zyg/YnFK6ZPtdaAVz
O0m4Rbkf8/HoL4BG5hDSSjaKtbU0/vzjdN7BJoSVUxUBhWepVmFl8l634uolZeRz3NNdbNOoejdW
in2HleHysnbublUAD7kk+On5hmzEckCbgBcclIUanJVaU3obQWs08czH8KfdzREIkqEWG1V2mIsD
IJQ/6qP4wQ7ubKPOmrq332j51RG8sa83xAU/I57PQTmE+h7leQVuYhzz/pIxNiVIIP++RqC7YKA6
yVPngtzwdNFSV4stLZWTGw6YRAhNf6sb1D6EwAD4OLDr7RxC6yicq6hGGulwil1wbufd51ahgUDi
K4f1377zFADEvDYvd3NLBEWQLDphdvIK/uEodD3g3hOXMTDw/f43rP3KrbfTmO9aSBRdfU0uA3U2
e0VKQBLuXUmoT9IELGw5VGVyWOJoYDoomY1UeA+3GLCdJtY9ds3VJPXA0Z2orw+jJ6R8Iwan7t9M
RqwSz9IUirwE6UHaN67KufjBCa9lYO+A5QzXYbLhThyotAJUBrFGSl7ATOvKAYS3eDX7BfBUJ1j7
8/gU+gg5dXBel7HoMzFpxnwJ3B9DTExivjYiYefscCKGXpmqFojRx0NsB0g6z42JVdZNH8+rd4pE
uLAuvhBjb4TM0qeDi1SZbrvcqxHLUqzQWbRu0IYljnR8IYcQC+C+Pv3OFOT8F3pQJjSVWDqVIUaq
LGgso1t0ZXN5jOdOarEAS0kdKYYVVf22NdRM77iWIvRwyjzFPumIy/eFE/s7z136Tq9IlzGbxnBq
lxu49CfAUPYpdJ0crLhN59HPm2u4hPhcjCCLtBw58QLn6Zcz/lt1ia5ddCgJT+HEhh4BknewDuSt
wCIgFZ5q4eq3Ym6nxrmQ53+/ui8b0QmKaE9u1Y5eTR1vUI1i30v2ePLUPywv9+1fiz/PHWUAWU/b
mfhORR0nRgAToTkfdDmS0DgUL28DOhGs3i9Kl4lJeJMWe7HXbOjZ4T/pB+JYaZlDUGaEhAhsXc/a
xmz5MkRo++wclfYQgA4ISJdliUX+wBzcRfdKFoNLAQzMJtlIjXXmY5RmQJ3WEMzKXmSyKqtiaswc
rInuk8rRsMoWWwxnO4xEm7GGnyERapI/T7uflcrnZ9Lks07lttYYSRwr7R4i9wTPSWJo6xHUpgl5
LX8NSbHCtjT23G1cFKOBmqTR3ex+oDL52OTP8+PYGBAdRm3GFlAky+WLFqP7OrQXR76s2vphcUfN
xEP0yFt4HtF4jZLA8IEs8px+vIoeAz7CiKFbO111Vd8ldyPMkiHHIJEqIl3wYhqH4R5NWRGcvywo
0BUYimpLekGZtGIETIXpDPhnLcAWhKfYo4R2ficvf3HhPOHra8JBXlKeHnBMUzqj4297BBY5nMtZ
0XD5xPrjWUi0QOHSSsUQ8RcebzjFbkobQwOqYf8kVCGOKek1RfBPFVHQGXLoiqxwmITGWbtYW1pW
X2T0ZnSzOcA0maknZgy7si15EXDVAHciXKNL6WP0SY+//Bf84ttgXGVl7Jxk23PhaE87ZGWKZFNj
xhVgRHq1HWSDNUqbLaAmgrwOI3dBLdxJEaRoOpRCfpyrxaDz5fsJm6LzP2+sil8i0QeByiWXh41w
vp/8OHvJGpZIXgxDoB+4yzbuPOtaqwb6xyKJcqW6L3BHJTpopPTy9SsBw0qQtak1KeOtm6NuIoZZ
VueC9JKhsgfjCIA820SZtl58tIsEfqI5A7mQlRTdIIXiUtmP1SM2pIbpkyF1JUxexea6zYkzIaJZ
TM49ODT21A4jvwKHVnOpkjq+4/CJ0NbMkTkSZEMDiQjMiazALVqWyUJ2FGkGH+waCJFWGnKr0ltW
D8fIVf5Lz52jhxJ1ULQeNcDBRlAi444rF7wvIP6HICocSmO46O3Ta+kfooZMgvUMofpqHRmwriMJ
dWBo9T9Z4PD3kJXyqOOE5ck2Wm92xKviRsTITXn5xFxtF3ekhkmu6h89YHKl2CqFWhsRDEbcc/Nk
nKj7kmjQd3pKoUSu/d9erz2/y4FxE6eIDoqQ3qgWQ8IADkPV7tDtATlyYJGwA5wEOhguCMPUQkg2
gHLco3MS2Mr7W+l3VnelaLNymTC19Zl2rl9wEHEttdAoPBOLNlQTXrpsmDq14Poba74poILfc7Dd
KF890khqEZZlu4eq0kwToFZukxKT9ClT5S8AZ1Nm9/UDo8Vj/6404v1qmCjUuZkxbzRyddJp3wx/
IosuCyots31+nRvLoWPQlGFYmhzlGLUrrI9LUp0iVsiWpFy6WhdLVUgCkn6SILi2LYcAIkd399B1
ajdh4L8d6Wgtr38PegOamq8WtSC2+IHyHoEQf6ytBZpE3RdvybLEJhNTK6MdKtn2E/DUg3E1xNAo
4FM48ki8glfKgUazEaYyeapH/iKxc0N7sh6zxVw8WOknhivP6J2A12kQwvQZNB3ldhS60zYgyOB7
JU2Fo7NYHnnIcdzh6ai694Ve6L+lze6m4FmVkSGWpS9caW2VB1dcmxH6SMsJ8/PCCexVAXWeZsA3
th+JLiuFzgCZg4p6o/gbbArEmwKFlcop0Jnp0EZbNq9NqM1zzRy7pVzdih4DvJBoROmsGU4Yy1pc
snXHfB2TIwdczbGovWPiXy5/Zgc5ZMV8GN1G3CUr6qcitTMYQfyRYuLVZ8QHhVK6gFNNjBx85Z5Z
J/8ZLz6uuF5OicGCExi3ijM/8cnb3s90CYUBu/YGsme7c3U+1XdXTbm1Cpy48cmVWSz+fC25wKUk
KCb6vWX8BiOhDOzbL/sUfQ0Nx6kf5Yc4DZVlQDcwTcYSp3wOugSyILi32L70csfRJiSSL10ySBLA
T0J2MlXtcsxMNIGgDRqfGWhShL2MHWXHGWLI5zlVmfd/iMsAUCZKR5WD0oMZgA7lWfbE/wfrcr6R
4GamkhFIgLoAqp+W+psQm8LwaTYe+rW/26nlFrz5p7mZ6LCm9cRqfcpsOi0skojk7iwsIblMOJ8k
6u06txOT7e5vURStXIyzoPNwrz0SNzo8U1fOymnbVMAsSR3QHZnQ6LYvMoegc8/A+1hE7zAYrrNg
eGSKOvRelnvgO8AGKRYGXkd/jjAFsLCEckLEIpndR+Zo6uEj238sa/lAB89o6Sem+5QVFH/p+Toq
R4pPc2M5WoMjAuX77MMYK7PgQs7EFHG51UZWVgLij5ZAtejgxYFkf3cvIC3NCSEpdRYXuAh5gR24
vlAainJlTIB0Yb7k94ib2VhLjuGgdVAvkb8ELj/Bl+EDGOw57VEEusowqhWFlRYpy0cQ1xg/c/QN
6uAheGeQXfIJ/7viNlbSQIv4J0Sf8fRr4X2FF3LmL6P4C5OvYs46FH5fdy+s6p9fBPWa8HWZEYUi
UClrptdHy7+mZgMicHS8luLisD7BcMervuFh6unpmDz8Nr20f+jhiag3WExfFBVdgsOJmiLqSEsh
FByR2pMN7K4Q398ZgfzA9jurArMHggS7DtVKI6Lk7V0Rj7QnA4U//IrmF9HwMgdLHy+pvEHzHCTO
3lkyHEwyhFmGj/WboRADwBSYqUs9im51Nywqq1OAcIhpcFNOWhYOMpK0WMifahi+WHPZa3PLkb7G
rqTfacTauVxBITDF6Yx/CaI35BIsUdZLlfzG5JsX/XUSEkZ1a6dO7UiSGH2Js5KLBe/YL9G2PMsx
af7dzwq1bIIJvfIbo1faZbogF8xjYnwEu10lYjgUjuFVNnV0WdJCbEUvmGEclxWVFr3t54VWkJZ/
t47mZia3wsHU7A34a/R4IwqARdxg+lEofzDzL/zrrG+iJy/efzLYoOKTxrXoO9DXmMiZR06HrLgy
vnJWapB6hUcS8J6knAsnRB97fdFkeKTz4wqMsMneAOZC/7G8ktsLqxLg5pZPrtQivvFyXfDA/aG3
1gfhk+VpkeURUI6TJnZzuHJfiEBYyJbS8zTajBKbhkJMD3o8SmpA0KlkjE79xR4qGhjNk4Ivf/xt
JRsxgTX0aiRwDOO3HfiHw2qbLm5bmvI3hnFkleVYwOO8IJCqSP7HCXbU7myDW8z4BVp/qrG+CgdZ
9uZq7xDWr87vSnrwbDJSeTaES6ILRzDTerROvS5dn3eikuKLdr6J/OtQK7b3JZqHmvpOqs6wOUlJ
tc5rB2n3QiTcH0Miqdpff+Dw+TOrlc8jgj9njyMNijWUDD+K7J9mWosc7UeeFfYMo4uPeIERnnp2
44UjWdOSxb6+SGGPYvFDbloXMDsKzhEgpxdpECOn6yDBe2hIeLetHmTnqKWZWsuDZfMrqjyibOGE
6xdvklTAGFnjDRrqQzBhiLr5AvwlfbTqA8KJcWY4YntaTIURieBoZWJmdM1NWvO6gIOo8bVVGRzk
mXKaH2z56VyeXfQbXINEEN/kS0HZ4ntiAdoB1rxCf5oBLBwmribDvJeWXDtbPJYxG/ypo9AAvq9J
pSPFAajgEMNnt0Kvv3s4WALS+IRCIzf0u/WcMFsPcC9rzPmk6PaNgsbjpE+4p5HKxOkAxWybI55i
r5BTjrt+EFfOU45I0NM0kX48AqIbY4bcjD0FSYvzMojdP6Qw3f+k/tgplZ7p4o1azHbo4lb67eNp
XK4c/Wmk9+zh6cf0zlvqZh4tKlxGfZ6GQMlKQK3IcK7eEeLK73cQr7SZZk2KuiWB6Eo+mwdTrFz+
MW9YBl6Yt163Bfx60CJbiAm+Vgc10ea3E4VpQ9dQq0KLoO1hRhWNhVApzWSGw9BywhT8+QuBgX3j
arLYvQTrNXKl+k7tlOe/KCizUO2OSX9Wd8RzhI9NcM6kJWSMcU/GZilb47Tmg8lubC3NBi3u2j9h
bp8QYp9toZBvXBeVCUZqs8s/aPnMSxFVvd8pm7o9/5xaZwSRE+lQYb1jQfbstt/043Nf5ggRRfO8
ccSyTX3pmEeQWnHnl7FaoCwXdAXKz42kkYOrw/Fa+12ARY1nORtJAynE9WRk8IJ9i3s1Hhh7dniC
pA1hR07JYBvTLrjfV510NP0Mw62um3mlKlr8xSaZvC6T3iDayQqbC4sxlBenNDJlSZdxIqKADLAt
8K5kKUo8/cMV7XZKrsv5VpQ/IlvUTaSSO0XpoP6b/ENoWrYSVEVn81CRQthw37yhxsyuLeLTFZtA
uUuoaGd+3Vp0Znp98q9E3Tq0H6VsIVPT6fQIpeiAj4BErLSP+B9WnLYJGMUrv7oNUe8fPK4vJpkf
WRYXMTlp4j0DBUCTxdbu3mT8+sx+kl0y3WDHLUu4DgTEaodKbRKxEhx1bJ6DqK5g1G7cF3LZcY7h
A5nNNfJ6/rLRuVJ0DeS0aE78WwGcqPKr+6OMdSicO1A/yUrhHVHYdWefuVfhMwelcupd+MTU2hty
lJzOCKKXpJ9NXa3qRhQkIidI2M7q6RQ3lCQs33viRJsiIgZmqnyHmY/r+3yrsuBFB8nXzyn4pHlW
nC3aaWaww+PRQhhgSvGEN4Borp+SVSTy9io7ZNISN5E2LVyEr+62DkwNz7s+akcbOQTGq/z6IuNp
ra3Kj6k3gr/5Y6lQgHP2Wnv7W3DgAfT3NwEzgYLl/KtB7Xshey1ZrZ78DGQkQSsd0MmywrsgEnDL
iIh09ha/YDSBd0J4WVMppL5mCk6Z2s+ohLzUru5qcrOf3KX2kM0nhqrViyFY9pYcCx1JtT0wepqt
kwWC1BzIpUUgIjSQCzFw+K+nD9eU8e6C23T4wiMPGI5ExZqBU+miYHz7Ynk0MOUnuOSaNS7hSy/1
nPrz0kbU6VAYPSaCpZO0F8gCmGQscCswA8BPSEyOnukKt4vMbETev9qe/2QnDNUHxZN50GH5ykwu
QRJ/KEZza9ayYKkKDlsvLG19UIm5i1QdpdNb/LTrRN6rradoPbDXg6oOGJS3VNzmzs/tNjOnmNSK
HAnItJ9Ugol8QYC9xB6LJmWTFI06EJTPHhiF3BHbjpz98M1axyVzqL2HZ06LM5DJlpRfv3p3O3Vs
/4h5dGzagiUaEqAuteqjenvxtc5UOaJQ+zx0sjUiaxatpWDpp9r4InrHfhq/vZizJwHE1xRizai3
oWtX1vW5rJPH7xnj0N8HkxxQPZlUrmMCdm7aEyXafQfnFztcHqHUQ4Vyo/8b6dEF2a7HV6580PGn
2Pz1TtlA3I2INWgmSu6n9I6aepOZEVXeK9XIZ4JUIhxaAPg0W3+gk5aK+6dBmDKXIatt//VZwibv
hRiz/YQfTi7kd8KSzjXAPffEZS61xQzSzwNIkx6dJSVxTAG6Shud//nUAZYP7MHUK+T+OW2S5DJV
1m2kEQs3ptQypn8IDbeRjDDuqqqDQQAgC9N+TvobmaALOZ87LsXNdKiFvIPD/Fwd9GUcon4+DofA
ZZPQwEqBHguPv9hSFJlIq//Gp1PQYNK4VrmOHhbTjoNXcn2hKGP/xNJKPk6a/46D9ch7WAagHNL7
vNlyG3PNCe0FtWXCUHv1WWLzygJMf3sUhbEURYxsODrtdHQZaPyv5H4Jx7nXnAgWNw9fZQ5xcA97
FNqoeJ0AyJ5QlOCn7FqzYt0IT484R49lWGM6gD9pR41rC/guPPVWrAAowQAZMr8m8eEj7mF9UxnU
bNmfA6nj8mhcodBDotl2gENe6LZublny5msmGHKg390U50Fd4LaAWcoLNyY0OOrlsEygOTeT1hj8
nm+m7rA0SRV3ndM79NHmbZdCJgXtGj9ySGX1aEIZLw4JgooVudzPJ+qDY5TJSMquDZg+iZ4San39
rMnGlLcSdrJ1g1jWH0WJ8O/uYN0P2odJlnAPVfbNq/o+3dcm7XQ4X80dCbFyaBT3RNUqdFz2Qa9N
B4LJOhVwqw464kvr6msj4my7WlITmRDZ0HXFBZ5NRTqIaPiMdJguaC6YMQZ5Kj7HaU1/vn2ocoRc
o0Xe+qKipsUQsJELY4GmumtfN6uOelqtxKc+XQcyD9DJUUVYEgvTq6U8OgRyg109WK1h7oEaqfc7
A26geGwglnxbqMcVMoetXaIjxD04xBfg4JmEJZmhqACRKKACa+Wy67C8zHqTjPSHriUoQYAvfz6K
E7KCP0IipZ8XpIESvXrn092/IhurweqYjjwa9M6TuUmCgjcvv9YdOa360AdNinf0D+p5XeH7iAEH
P3OSIUNhF5mDaqT5LTuUbZVG49jqvpUSVRFURcP+SOXEv4n4IqLMHH/WnSZdDdcRAxOeAf349viZ
A93vO0B4JKLWtPTuJ/T4hbzWRekhBE8Ym0lFyCSxmsZxu5ZDXPbxWQ5zzHOfYBZ8h/sSSZ/Pa+8J
V2RzpyqCA38xtd/igGv1fy8lyPy+uUgsBbl/V05y+2wl7VeMWBsdwcCsmfgZFbTAJzA9RUy41neA
/Yw9XM7Xqiqxou6I1GlW6R2JIZ2qJsS9w3yB4VvTN3FzxG3ytHjc+0ivhXm6N5027Rt9YSaq/xVx
7wzyHd3nf2n+eu3YzWxaRv+I26L37qKsDOsZYjaBQzSrUrlSkM/uzMUs+Px88eWZJb1M/HCwDJv8
9VKcf249wdWmghtsJuH47HTe0G9ea9JeXMl6diClE3MmebztS23bHif3INzbeaAx5B6tQHYZmcjr
0dxMS3etTR8xDuBXlqIg8zmTfexR7IP1iYMm7qJmu1QWTNCvZo1KsChg5iI4L8LT4T9KmojF6NQ+
FfMpv8cdMSDmZld3RcTjBheU/uALOawmUv0qjdd0UeXkkuxDekAnZglBoH6LdnnklDLXU2GWVelL
8zgdklIJNtBK7r+PqXth/fqOUtEvjuoOuNW7474JjW6+qffoszZODAnSxpNzlQi+e2b2XgO40HzL
gCWv7f6lmg/yqtGOE934Ru+RFLjoLstwyqoMCZcu77VnYATkEd32WF2sZc+qi4keG6wQG/jQtczY
FQQ1ChL+mzN4i7kp7vPVAO10ZhONNx6FHvQaRgIXN1bFBFi/Pk5jYfwQ6BRvWBTd/bCCU0HnUXb9
NYqH+lVjco/NArDHD0weVO3qYgGnmA+IhycZVPuYNGV2/IpklbXpHS7TnJWNQMR16F1hI6k8FKyD
4cTeWTaZovemoQIDSaShb9cO3OwaVGOQep6M5Q0fVo89vVej9lf1SvJX1Hduxby28L6XKq0VDpWO
z1fbikUdU3xDqoGxukWwpKHnCfqQ8SAK2AXygBb+0wRrMIWy6kOfm+MEo3ishIZ58Ct/xYHI3ROH
gfvhON3D1c7ui9tod86gdkZSS+/rfsUVbqnX3vdllJh+NFRsZGamODowJ20Qp6oji9VKJoEgAnso
ttLkYpnZpex+Xfn9uWkKjFdJzLia87fZBluKSjkJKRlZ3ghmDUvxH2HK2uNpCOBGeE1JeiqtuboS
RCgvOUl6dhdnfNmrXAuIH6OC4rZP0AQL3z5ljrF5r9zjijAWxyR4R/svHelNb+NSMrtkugt738WC
k7zueozOW6ehy4YujwpR8ajn1228rpjq7wAX26J6O/8TiorMoTnuQcQ69n7gFTfMbmAHzuQS3K0T
SQ76ZjFFy6NAOCnOCEZv7MSDPTO01h/wAMFrywH7Gz/RYo5gQhE/KnVwPK0+IgpMAZhusUZU6OEt
sIE51zJCNE/a2rA0cFuSau0SdzyXkHV67lXDd5WzpjqyrxiQ1FTlI/1qGocpPi+VHgMuS2cSl8fI
Iu1pBwXJjpXZER1mph1LMQcTQcOzLkXq65YMC/9isAVsW/XyTeeD/f3ks9GFwng2yDtXsAaoYUFm
mZPuaCSntNICm+SO/VtiLbUpJFRChet0TOIG4tSMmU6cXcnFrtJQNS0QJi1MYpyxvDVHUK97mzyi
cBw2vjXz+TD9HnodyToGXkmfDvDEOMvZfZpeftuJm6DpGwFENVA8GY3ViwTaZgB1EOXj8gGDTJVl
z7sM91htv/V5JH2DjhVqZo4EGsNovXNOcXXcKXOstDUferkfNZ3ZMdpSgRubwKuJom9WlX5e5FOY
fqmNKQavxkLGEFqZa11gVni5JP/f3LL5Ib3ae9wtOOq9SiEUl0dc3G7oQUBWdA4nq3PPiLGd5Pg/
PxlYdu3jrOC5sKXNti+6I8dIFsuavhx9KTygMoh/PUciy/eGnFymLe+rktsAIbHbzVIdoEVht+Bi
FR2O5Yph0+xGCxuskKXhltH1rCSRUhpmT7qKGQ6TXtBZY/9CF13dc9FMr+kkzweJ56wIHwO5o6DM
2AG/uHXGPrrtM7uy2ue5/N3cHmfic1suMNB7+5c13+J1QlS9pDMOdUFClMOQXSfaPbKUXUbHPKmF
ft6HADFbcmR/ID5T672rKb/1Gu5DCDrAUdk0+iFqaZP9fK6YkHpMRVHnhm3mdRbXjDQ1wviTwSr1
RKhKhc3jJSinTtnbo8wrySpoLdpCjDe8GP6WTLMb/lKUNVVXp0uWrLwQTSV+K/iLFKRlo+SyTdpj
UMw7k0u7E4psK5S0IWYqaoBRWkOP4ARLFlhjdve/D9e1ZXM0II+1RGFXirTVm74SeEVAUF0KbyEk
pCdscr/XGX4jqTDyQuc9Eas+GtU9Nvnd/VxDky1An9oUWyTKB7zPNd9Su7BxV+8dbvf4WY6Qx9pe
/hrQ5Dqx9J+BbEzJ0q9q+iNlJ51R/zTLppMfqXV0c3JTgfPtZeZnI/5TG24IIezyZbYJboPapDO/
Gdby25X2BobIf4ppo5d5L6rVXlxfmoddXRJmbu7J0xOPIh1g++biuoMLGRyV0jEAR7msSVHwQcjV
AV9UgR01GCYYOYUhnI5GCRJn6mGqqp+lUI7mp/+G/VVMV2FzVFXCCW8nKQcLccNGAQA2Mz215RU6
GWOXNK/0BhZr+5wLTbNBp11HH+Wj/pJ6jIgCtWsEnAIaPKI7ZYktp1A8f5UEWH3bMAbcO3mqr1Na
1lIYS4zIfqQzeoY+yUiF/+UTDErF0OeWjiajPntc0Hq30clLz+ZATbIKmszsx9LP3n8RgOwDttrm
AAvkyqoA4mPD6U+diw+jNagWoyf3t1bGGBzSIGMc6Q5gbS21yt4CBxU5eiBGmM+7au3C5HZYTJVI
W8GMzJbyoa87VQLvPZnk+/cOhavEBIwoARZrCKXXPw3JO6rRYG8qvDGjvsMDgTCVsLgcwkvr2N05
LxY+py0akrT7qBhZLM3nh8XWxSB9Zr30cSYz7aczyeafZPgFTGdkwcAuZH9OdDc7UIqasrE2xjPe
1v2QwfhwCcfHzlmYSWdu1N2YiHvw2cKMq8X2corwSbKAf0kiNV9lCoODF1dzSLzhkhFM8uTDZQSf
v9AjdxhRg462kFar7gTtaLQIgct5cc+2RrzErni1StqtE7KWOzYFX94FNXgRhXRXnuq2q7iGmb1/
M+r1TQ33m9+9NZU5gUD5SO37JJDk8ZCbbAMOe2d++7nPA3hWtdHigk3s+SuQDiK6zdVdAvQfQr5m
iRpeAU4kj5AA5Xt4b9wVdTG7kRGjAA62dPsA3p1f7IQa83V6n55JG1wSAsHQW/FnnzhAyED8Vip9
NUPlRWY2lbfMJMqaD3iG4fb5OXGAhgb+FHb6yF43ozFXKLvHXyIcB2Y1GoUiyBbOsSsOexYXVxi9
L6iST00aXk1TJXEoa44i/xYfTzTvz1aMr3QWIzUoLrb1IHXnz6+adDTrgi3hyytkm9OaZOOAq7NK
2k4gUOsDFc8VCYKZbscwk/5buscUM4D7jYHhFYxrRFKYuKZZB+3jG6ez0a0SiTJe9TTLI/jvxOFR
MoRSmAGHXUSg3zcV0vEKih0SrRJZSyBhTzsvydn1ajrpRL86ZCrs+46I5qzHgmVAyYiKBvrABRL9
oS64mQgaELFGBF/1g5493w3sUgj1gY0NMBI8JSYX7DtuIeRzuxLNFeVaflV5oVT6yIZlNH8TBwh3
ppOjOOLC8PEST7crFCf1aMYkNunM9nm3XSSjDssC3EeOEWrnxv/7XKjxOuxg+bOAvNfos5hXPPS+
nNLP0obZ1G8ZClFjM2/1DnSY1athRX84KWW8zpuO/o6SpFyC49VlCGSQGKJikjzmEE7BEFSpRwyU
/0fJUGxTj0NDT83mG7JfsI5rZDAKGDdTP0/30LR7b4atZY42y3RhCglIwaCV5qLYRuR1oRbd5E3e
FAtlbLPAY0+jQeVOlW5iQszqJeZZR7UMDQQJicurhmVChOKoUMykYzmZeKLKsmmw7aSecUK5TFRC
QbQmcH8UvdUcTP3LOWqaTm9JkMi7zMErskxqaHMQIeI6u/ZDkR4ttCtULP3VIdPCma1YnPdTAi7s
1FzI/JbxnFZoUC8un4ur6PQrAGfKOi2CB6C/Dem692m2hSSkfTDT8sb3HM2vtvL6RnViKe8GP5sL
A6SZ57+2w3jxB3EtlasFyPaHCE7l5ETSGlnD09uoDHCX1PFhrU99VooOjTkzIVgWdMICgFjZxavo
3EVB5BB4R6SAIY38xbSFgK4/UNBvIYodB55NcyfPKvETiLA3uW4bAp5uFTuUae1evZJARvxb9Dlg
Z/o+DKXmENbnHcbPWe1ushpXe3eQF5nFcl8fNE23sNoH7dsq3JMeY/XWu8MsFz1xUchDkgyyDvmN
2mRoM22VHLwgHR/gh7fRrq4+aQn35C4pPALiRwbC3dhPEY/79TDhgbGbQIXJ2+PfZ8zx8YYFDu01
oluZpLTQx5GE9Gxr+vn6O6BOEyu1OOuHhKkVTGcX+73z/ya84Cuwn4Aoxd/WHUvcLL3aAtbXdsWd
tgGpEV4CW7g9rhVLueZdkUz7B3wu/87rUvjAceB8OL08OozKgWeebW8H2tjkvN+mbgiaiRNaasjm
ofjd/Nb9LLXvDfZDROe+Mi7XoDdkZG/H9ApJ+Dq/7/6IO4VLeT/Fl+xuXEMSVcB8PFEnJ5H4AN9/
/4Pbgz5M5P1ayRFU1Wq9Hq52VSQWET3pOYp43XwRZR4LdLHY0fGYH+dIc4iE9bEymdjfwSsf/l27
5Yfk5ZgdBJnc5q/G0KQ5uQas59zf4qKAGBLbpCRUXtZtfMq2tHDIWksgxfYK/iFdNCYhquNZIfRQ
uPJQGbbbSb1vzPerfeE9qkemAb6JITNUk/v+Tk1FAVnfDcFqTRP1ViGfFCdytQjEgVVyKEytTy4g
qbTplp8jnIsGnsPxTQ+sJ4d092hZVhxpiRtc4tGVEdUOmAx7Cd5b5ol/o6WzNO4pRtYL2fJYJ2U1
1uT8MCOjP9LoD5ua8LREC4IsrPXw3nn8yB5CCBPX2+t6jW1kxHZPo3uQ0vZUwqUIb1kHsP2eWxAi
3MxmqYDenZMf3N5YexDhnRAll81k1vZQ+GDhZT2nO15Wn0YSjao+L2Yqtm2GkoTuVKjrOtoPrKdc
PJNadSeWBHj3bLu3KudQXh+tHn0W1e2Gm8z0bX5+ETBLYDK9TvLCcZuLZ4AFvisojKzEnubFn0n6
LDapojEuK8qSIAI7LoEX4Qq7kwUFmAU5H1IZzDuTI2yRXcfCJfUXf8tH+Cxc4GSRBiFnu4UDLiQ7
52vhEgrTbD6lSHp6aVuQCcr1nGDJa4a/nc+7Gl5xu0qp5RCjKFlYykXBnkujgGYXLCidRbJJQrY/
Xu9pcJ6V7woL4aBuJKLgvgmQuSeB7YubW3Kwkryf3nXghdAAqsdf1Ie/riYUIafYVICCZFQDzIW3
mmOUtAIoKTzlN+49VtVgE9b9ReNmfU7nOdzBoqGGs/5jh5r4NixwzvkA2pXImm0mawOedQEPUrRt
EGhxsCqyo6ZmdknWYqeu3UBtr5ujRm4K+XEikrue0iSFVA3PXmSseO/tJ2UQa3zFDUstu8wC+s+6
cYbKMx9h+2OKBRb+YEkciT/cTSD5LcAViqDmF/nwFMdr6MdbzhBbLPV6u1tS0Uv7GHQwghMGtlvr
9rBmffF9cKfD7iKZ1z6uBtLrk+R9sQZm3NGSVpSpmACxxyqmH2C7UA6VFTy71Zy/hx+/MnYIuYFo
yv1bvdQ5PMceA7Iet+SBTvEMi7AYR0p7YTwyGSBQA/H0rqhSPbR7e0Qr1bUk8q5bwEJwT/tMc6Zl
qPkXSm8Rjs4ly/wkX6Ib/7Voi0FPL7X5QXiDNx+m3d6Y352mMMYiwix79yByMaRNSd0KJ55jinqT
ss+QHAgBQ3AM2KPVonkzYywECR7ZXA329DMjJNPAQvV+P4y++nHWD3zOLA+aDxcN+6edAERpTWZy
d7wllJ1yhk1hei85HzYQvHFl8Pwvc9g9/WRZdX8UrcNB3uamzrUrTWizM38aGY9ADAJlTkxODMzY
sWkWtpP/gCOxwnK+OHau0Z9q9tveqs+Zzezi+o0qdXL55FbsSCFb5bJrstcegfu1xyUuDzd4uOq1
Z+K1UQ928yljV3OiQASX6xR9zA6Q/T6dYjyGqO+IUwRylDNXOve+nQV1SNMpnQcbnG6rU8v6v3qS
PUGL0hopP8Nh/aiPXMm9BNQjn8nZqf2SnUJcOObVOwxCAC2406wNxo3uw/Kd/7cd3Uc4J3ASPJ8E
Psk5Hrxm3uWfRv+RlQ9jKB/iriN2+yZmtb1264sck4qOaJZWd46TV4O3zChnfTelN2VLu1OoAsku
WX4kpB3pqJbR58LALflkTdmvtqzF39nTx3aesETmCFSPU5axjehsi0Ns0PHXPxg8HjRQxtyz0M4z
tqER9pGeHTpiVYb02PbKeXpuIeHP/So9t6RPIqbuEj1QVvTaX6nOzs0Ge0sKFyFMK9WUoFpjLra9
xwm/V6a2fIOt2bQloByrYAwy7DYLigtHZKhEz+og8buA+nAVMsD5jb114yGng3HPQXLVpQs25Rxf
Z5mu0KmRp2f3/E0XuSIb9xQ9Ke6qvIYYlH+QcJCtOEF5zVfDfj4Oit+h7ep0Z9OXSBzmTwh0i0zj
nHo1lm+aAC/MF5V52ZXcuHYuYK07nsRyxBjNa19HuAxkDzZBlWwNwt3iq1Q5QPm+tJHv6KpcZCpl
jhQ2cs9BNt2YFTlUHJ1feafSIVaD+xhFwoH5xNrowjufNM4V94Mi2pYGj4IounEvCeFQ0dywGU85
phSOUu/PyEdG70kVvLNsGzWDMgJtlnAbgdUckFjdSjKOrqlsB2zfBDLffY3/XaeWG+OFpM6K8gfo
zBcixnpoQ92Qbs3ehy9P6Aj6hNVupH9GO5NJsFJj9JhrD26PqS7jYG6u3Kj9CfzxhInCviIjG9Vf
MnFjMtm/MzTVpV0O+i9fBL7kkWIcWn+PHx6Za8rLb/DmmVPtWK+bZqg+WthVl0ZZUxbeYjPYLGGl
+v+csqVism3As6/wa+qGzn2S9uC2aB84V1+hwInDQWOmCKeXCZoiv1CnwctNw7ZPI3/4O9gauc10
zSR6DSzjEXPczbwvy55WTZIjrFky16vZshsLQYWqP+bJdTk9XfdgtvAjRPdgF/tVLBhRmCdr409H
HMlBcnh89pwX8EFJ441d3UxVAUYlMjB6jzoFqxGb63asHjvmzcqup52IzA0qMOfzuJVKLfYKXh+J
x/QVwAbhyWLuiNOMmhf/njMezVAz7RUZ8jinlTHNYwf4hw2GSYFb61pJscFhaR5GCl7oVTdX8xks
StcnKX2/5w79fq8yXkEjeS2cdQPglXNXDpNBOf75LkuxlrHsus50o45spHxzJBKQGAK04ef5+f1f
N9g8rDgeRstGoj8l7v2tQfwPjSh1hntKudvbPkv7tOoRdmYnSCHfs+fyRXb2jrUSPYT2QV7J8grF
lzMzN5jQfJ2ekVpjnfXlqUwqKGZuGNl6QWqpwd/3FngECb9RvDOlzbL61cPq6ZuChxBMNlIfDWJm
mjQ2WsoI/Hvawra75kf7+aGuGjjSpt5eQpZWiwbNeuKn2OYQLPrP6X86iO6qeuxgVFyQfWfI30kg
unES2nlvQ0MqclZfWg63P8f0pY3h44j14WDR8quO3eLZv94ImZPSEkLeQluCptVUUzjZ3oBOcJpI
/rFqbBCRfoqXdcoeKFO4xATIoMIJmktN2pKzQunVP3MaVhtZm9i42Rzt3/yDWsF7d0qxiUuTqGnM
tvV71/sQPc85fp+2n38nD7o0d8zei7zeuz50mHI5lkr4z6u3cxWe19Xk9cMrkjZ7i9W3IF7Qni3l
eo4zHCZoPg0qoRA7gNc0cSZS3IOhnKn74P6HQLrw+DCF/sMsJ9SiuNzPJQKVizgUQCPMuQ093L5v
taPYXjL9QamBpWUcCwsl31tamygrKECX7BayRuAR8TgFufP+sJgnI/uMzeA8ktj34qjGWRvEkNfl
77oO3LRKFPQ996JUjFzdhmjAzOzuUvRV+DJPtrC0TqcLi8KtdIvvaSIu1bbjqcRypT+tFUH3e8Vs
/rFIEPMZY7gj71iZyFW3p0whsQlqxURT+/PzBC57x5d5mDU7xjKxBN2AZio+2uX0uxVV+UHt1gI+
TRN1YFyswoz4ioKw/8YGnB5vsqWm5gUPpHk3sL7heJKbrjtvD08fFI+NacNTEU13Qwp7f365u1xH
QUjcPYHSr3+LTY/jidaYLYz/xBRMwCea4hb1ZTFwns+L98QI41ytBRhHrMxLyAxOAqTUUR0PjrrY
Dk35a/lCoWZk8Ku2HPcto/+em0KT98sA0u3kGeWBlofPEUzOD3V8rGCIGyoY+IrPKpcAmjQNCQiQ
kZkd7cPqcAd2a7j6n0O7kKOAvANJcubF94k/1BNsWMGN0cf1t74HpYqz75NEANfBezrlUWczvvVv
x0IYBXuJXLpr/GwwNkjD4p9zfoF0Naf7JH4YuleiWodU6K1i8NAW0TOwkppUT2c5E8s+KKFabyAO
HDczku0HIlz2QUfN5hWbQIyPCsjGljNH9yCGez0noXqlSz6ybVljnjrmykIWrcSzCV0lLaMfZsci
BumiNsvxV5SygXLpt409mLddDFtFuBjW0V7DaXH/nbls53PoLph+Z9m3Pt/Ddl8EyfNImD/A0TJr
2ID2zaoT+RWCLWrzPo0zHIgyv+jbBK/1turwx8nEy6yYs5u22H/6sR3OCSmj19GdpAypxaPcb711
Y+LIrIl/khT9wWT3ofJaRwXJEAcPhdXfZQA9Id5xFASgOWlNGTW4HOEPFRmHWHoMSWhzVgMYR0N9
hyjrKPxkmL4QibXmAyYAG4r4CAHSvAGEVSnAbEzwUPZlw8AY0LytjLUZMIOgFinsUk+wzhwLXSBj
asUPQPWXnDhO6b9btyO9/i0dfPmXUiaPUQkX11JRhLOHrm6sgIHoRWg/KRgtCjAxjQyMAbPSJRh7
wDnrYch7Nu0ktqHtFxgx9dKNa6MM9Q6LkMkCeWL2PW96cSmYBtFa82gLyWxxJevWKXd0biAolCYy
WnueMOGC9xdG7PMU6sdUdwespKCMSaEHJFTzPQlXnUF6gx0byokY/KTHvCZt/TD4hiOlPCtMxVvJ
QcWU/XeKIzdGFcft95UnvSjt2Q2Uw4rAuXV4WqEeTME8zN/RIDsGzQpPWST2Ei0HW7zPIj6hBr+g
1sIH27CRD4quNHWtYsget4x/Z6FccvZYcqoIP4eQwkUNCN8wfOEhLCLmXAjccWJ8/CagdWirP11T
GoWYiEPcQ9/SJ8qVeP+S0IrV+pqsk3IebKqYBtAnJqjwITLNvMQzTdY+qWtriUNgM7JeUzeM+1EU
b2FcTXmUDu3Szex/uVqyvVvfHs7UeJyEJ50f0ZxRN6MBmPuiP8aUKodlLtmeW5+ZVia2nuFvvmek
juC4OucUpOtA6EzT72VueD9Jdev8BCJHspdc4oWW9O41PO6zoxvol3/8Cs4DiuD/vCjtecopKQ4h
uFBVKrYoK8JRq+jx+6mMD+0RwZGqxsu4Js+q/hRrt9i6U7rV6anMga7Bs6WKlTtsTRGAWDcpYDtJ
qaHQM24bLnvdnQeGJH8OMNhrtviIWBmbZG1oyi2vWBzflcW8xV+sKLzz1Ut4Z22i0GIZY1VnojXI
MTsAHUHaLnegrgXWo4VX1Nrc4w7676Vc9biheGGb1gWrOegwDzlkWQCvoySJkzajQsqlLshYip4a
C6h1/HRmShuJlRMzZ6b0Yv8GYFMeo0lGnR/d3SYhAjywTa2a7wUUFqH/kUhBVP1jItraA0RCdXRr
Xgc8S3de/mhGc8oaM7dInSbo5x/IscqQaFzqlDmENrq7j7Hz5/r+C0IXlhA4HJBq68lXRNhPMV93
gJE3rXQQssgG9sebWyl0gqMPKT7dcjytb4SPsRxmuUcc5SgfCK/HScISaEUIJDR0fBUHYHHA3LZM
vA1ZQciERYZsEqg6pWALb78XsuZrJJPj3jNI8hj2TRvOJMsUHd8iOLVOAgcC3dCPDtyRFMFfbmjD
PmduimbymE/xFiT8ftirE8CDVAlIXYhsFTa+XAcIJNnPN1AenqGEohq7P4E1YKk+bKRmFPpa5wlm
XBe5S/ukTAQX4O/DEuiFEO4GnR7zs7J76T/IHQt0mtrTPQo8a2eI3nHUeQSBHx9W+wXx/8vxpQdg
aej/1WBfpolHwGHPAklXj8PIcgsKrxEI5r5E6tUugJco0BwCB6AAbWNep8i/6PEbGG65mwV+kmRo
iGmzs+cpJxFgvtq5EvtZH9C+na5kVFxpmw0ByTWOSnU5lUEwx/CuaVV3UgUVJ1RRH513dQp2a4Xg
6Bc/qLblC40U1G23eMLt6MBKiND/SbkQzbdvYzOd/9K7x/68eiq8yWel8gzrNxSFnmiJEHi1CRi+
fKrf4DqM/xHweyd/0HurAVhJvkpOnQATeJq55EMwmjv/EvQeZkvrQmZ4K+vOvKHhjIALmcLsUlc0
XReUWXwIZggncBbyAzj0RGpb0EiXNUK12fQeKw4w+Vrg/Vl17zu5FGexV+ni0xP+ZUBcSGhppSJj
2w1fyM9/Zg2adcqCyhUPbcbRZzJUB0OOn3bDCxFH2vrYU8ibdkVuhimrS5vu2VLntaToxVNnTQ7o
uUJG8lDJnyZguN9h7RByShrSuT2KpQsTbkaWezSriU0ksHOPsRf+i5gGk3xUS6jq2UE+sVOAij0f
dQY92R1Eqd0GqO2jkmNfwbhD7FcuCPmV8zje4HPITLA+7k5OeqRET+ZoahEHbSemM5KLha0xXjg9
5jDCHGH//lr/H1qN0AvIYW44nqXHXQjDf5DNjtCluqCuaR474ZFCmpheNTiGK/EIrC757K29JG8G
c7gx1kGBIGaHTXUaActxIAEGj/hIjTutt5BZP32qVstRrTZR0utC/oNckcWV0eFoII5EisVGSwoB
DbOeRlDo249njRDHK0sI3izK7uKCbcb1GYfeB/QMfma4m2MPyVaKVAWVFkvAXpvPVP3bgh5sN31j
rG5SeyzYvIWPEqSGKWkad4GyPBo512v/nYtBb62FnptNsxgXD2S43EAsUMJzFxGcKnU1joE1ACHB
wBX3No8EVfrExCBDDH51cOKNp/OCw/8e7DZOya2XWntSwikEVXJOW+qysxP2fA7YKkszsLv6XKox
dL5AT1u0XMew69bEFSHcgwFKXQoETImOjMNv59LFWxKlejlLKLZ4e1cvPgtRCSYMkmjTdpA1M/Rj
jvyON6kkeBwtuklhdnxPYFDjxaBQdVkCTZQuc3/s5fwVDrpa6D9nKPYgqJn4YFR4L0uOH+mTDX5m
4era5Zc8eCVLzw4zYguB2fbYN0qPHS0NCKOonN80ZP5cHtRbA/UrzoQXS1ACbjtFq15FvxXSagqr
viXo0hefbRHpt95GfJZ7Hnhcq6YLGdib5sCj2EbDLmK2W1VuTTT3ELZLjr89wLsF/aPaA+FCJowX
zeZ9TzoWJQAk2vEo51XT/LHBx+CapcW7OzrWUkt8se7EYv1CxC+JoqzvRNThLxSrlGqiH/oVdxve
7Ljbyk23cWUzmJKZ9Nhjqv6ZgD0vJ4uh0LSjOwLfIufox5rqFhkPa5zbtHwdpbxH5ciu9fnP0Mcc
OLB2kHbF/RUqwPPi01lmjWrwcSfA9jERFY1N+mhW87OweGsnX0FVwnlyFuH9gFwnwlo8luZNRqTf
QzfN98TwutdUWghubjfMPp7G2bf06LckCUQRZRbMQzNtStiD1u69z5nkuuiphW57cHsaX/EJbkEY
UzviOp/Q2HZflruMu2cYG+DeAfwjXrBd+0B9XNDBOzjYcyVnqSh2yHVG6KU2TBHO6nagk1lvP30i
HYu6IeOoOUPPgrZs4nNpgnwFZELHK6A35hxbJwzcSSRXtoZw8rJZ6fZn1+Ov5/gWAgmnd1PaqlHe
HkEmKo7hMPd7ePxBjODNhuQQes5yJx1xMzdLkpL7tgd/jZiqix9Z7ySLHOK/Wk3KlzT0QdspGtPv
umqGMW+ody/h2rq3Mg1jq94Di3oiIipjNm5D70APmT4K2SgFfGVabolru/3V5rrhnLM8GvTYyL20
0FjapcEOBdOiKyFJBmwzZR7LRbVTpns6SWlN6izimLcdbRMVIyw9JQcGEj56S4luAWSTPCjMSbBM
bVOT6epol3x9DW6UY84Q+7vKzRH6/Xv2z7N2Iwz+Y7H5mLScf+2wT6odJx8j/KW4AQm+9gOo30gi
FrZFE9DBnSDMvF7lcxW/PSSA+XXrHZl0EQEYrPvv7JFtGVGbhxylagw1MIXmu6ocoevyqHuF7hmf
Fv9+DD49u9I1D/3J0ra8E359ThANaVaj92pnWqH4rXsgfVR7HbPSURuDHtdb+atd+eGaYs8n4PqG
zTJFxN2Yux58ao7S8kCEm0/HammPT43opq6GAtjIOfLAU39mkokBRT8EFH0rYyw5IlVMrFmvTS3F
Vrody2sK6bGQKg+011EVCAXhGVdCtcY19RhWQvkznlDblzeifDTprjkyL/tc/u3RizfosbxWzOWL
HwTXRTyFPKJjvN+NX3hh0SP0iKJnOKqW4e6cGshEIHR0GRb0RcfUOzkMizyeq2A6Pwt7T7hYdz5n
xUej3Zwg6Tg75+MAqoQRXQf3SPsANMXMSYyIp20ZLHWeNFwXNCP4yYkgsC/eN8Nlxn3flPJixzC9
1M0d+Ur7K2q8n69Nwmr3zwL/2Tl8IPoa/a6tib8koJb1JogwtH00o61Tte/8JhLdVYQz9ndmZyd5
+oyXF707mA6YZMAhYRgDSF/19DauZiuHtzyTnO4IObeWQDYbpRvYNAW3yFb3V7U8x/OvaySg6+vF
K9A2PLLeZpT2eQQeWd3J+c2+D49APEmi6MAWkYpxMNMnfbyfUYwJXtLvqkrNqPtj0hgUkzoVfqQ0
a89Ozve5P2jHpm3kWCLDcpp5ZKl+bD804UKhzBSMcE/MmUXz6rO+r3wFHSXKAz90hHdIPC4MaieT
3JN/G4DS1faR8NbXXXXbs2aKJ0n21infGJrr6y9Gm8e6YRXy8alEM4nXFlnztcTcY/t2HWv9omiR
6iYn2xh0WH+ISy+Uv/ExsPzy4xREwBFmbRVdtpLzUvnxs/pfz2ghjFhucG0Y5ambnG46+bMliCVh
H08fYbQ/sO1QXmqojKUzJ0JhcYKsO69fqW45qJyu78BmLBf/IgRkKTpfvBN+PFPs11rHo1wyiZnd
RDEGoVTRWc4dLBNtA2FftMFYFO5FdKmbsO3EvnMWB4/ZS7y1BrBN+b6gUkDjgQTr4EayV81DVqG2
6bRyPeKUIdeq/hRYNJBCU67Lhej14xOChYzvvBP6nMdaIWOogaFUDmVX13VaN+YJiD2xdqWkhLjq
4OiSupUZiIkK+BEqeBzclMO7KFKaAkqMFcG2b8ahRBnwv9z+45v/Tylp17gUChSDl4h5RIQR14Eq
AvFmznfHeobJAw1qO6/4dMYTh9QoCdiQLUkIfNungw7R4VdYTQSDUGTswduingy58Mgtk0csL+9d
fNxTe4dVMDTjhAKGhelZ91T6/afll/F4W7hqQTdwTAka/WaoBk2l3gnpfluM4lp3NuAQKlWW9JIR
+QmdY0BWAK0/8B7N3/H5u47DwP2MPcV3V/clN3OPayPaScvCD1VWyGQhMlGxoMWISkMfWSDWjWqk
vbmkiMo33WVSEEF8vlueX8R0KExX5p0aE2nWBhDnqtZ6FC6UEgS4n2z2IwpEFkJYyYJLtN1CC+vY
1b37GM0IIEeSNhISxthGUXDlcHJ1KsgyBQuW8aS35GecJgxBjmfc2x/jn+ly8QkM7quDDP5DRUKn
C8tlVTgpEmrDgbuh/qYA/nDt72xGHQXhwEXksl7Wpu5vpb2Gj2YhRqa0gLY8xJjPXFwGUtfVshpY
mvyzt3kaptdaTvhKJMcBKiraJ7ej7cGsdWc58Yn5Fu8V3wUmOzBw24mbPJsC4+yks8HRLE5lu//E
XishCTgQD6KBFUOJcR4/2jssW4xEcGGW7IHDf1e06yeo4Xcs4t81KiIOFn3aeTpRkChcdaOaHFZY
iYNl1+5fCB0RvpcY64cnlXN//Ppw3WpSfDMAcXWuei9x3SijISQNZ43HfaAZ50EFUl1jU7vzRo48
8loWeovq/P12r+wYb23tT4Ip1TpLV6tn5UegiGamha/EYyd373lqnupADfxeprRmxuY6tAK/ShEg
ARccYG8mbUpjSXOVUIljZNm351nbU3hYdTZy9nqepD51xDJOUhqozd/vnAj5Bj5K6WcDUeFTgQoF
cDAIPRKKLzlnbobnJPI+uRASeLQJqIS8cY5MwyNkZ4/VfGHtVbmZmlflnWZGoyd1TCzTkwEwsqEH
n1tFdaYVnU+f4YATsrTW3oi7ZqP0QFlps82Tf8CrxjZgqu1CS5rVPOX9PKDzgp51TU+jTSkVL9nV
yNc4teLAtgymE62gmNSQGwt43vhZQfZhUoNIYyMfAI5C8Lk1kt/kxYWtHyb0dh1bNoid4CzKgD4O
fE1dv1TbLIOUg+419E8NKVeBh4jj5Q726S5U7Pd8TmzjobqjejKukTgd47ngPC7c96VuexxyLx5d
cztF4N2yDZEOZ2RRndGqhVtlkYrfTjad0Meqh79hIO/wucEJMDvH+XHayonJixcxiKCeUddAfhwT
EePKgtfF6dUQ+oIVa7JA/e5eeNjv/3Oo5cxHfT9oz9yuQhRAZlTrgNmN424e9Ri4qMbXqdOJJePd
G7U+X/dsA/Go5Fx0AhYuTAT/sYXPm82YXf/EZWaRRmT7eM1wZNYmEyA7rrTfSGXuANeFqqfboN5z
QhojxmNVyD5bt3yqZHTksmvCU1n1Eyj5B90De9N2FQL6E066OAiPab25MTI4DNEDDWf0K0FdQt4s
/FCQ6oH5Poe1mrC8mnOr7xSKmByWRYcMzWVmqB40Mz6T7N6TkFzHV2Mzg8cX3mC05NBGCuVvyE6R
WYG6GF5uf7IKi0QCN7Ki417iMRJjRm1bPo3gSXynjG3wxYFslprQx5yFXM7uNYKF5g+9pJvU7juH
ees8WqFlqcSfuNcd/CSq6pL2CtxJZfwoSZR6nVqLHUfXj5zttRMyZYYWPhb3qTsv1M9/I4H3vzca
ufM7NKxhhCq6FJHTFxq7CWeGfm0Qq2FvVin0S1Y6FA2Qsx8YVUFUTMgjG9/UqxIq0b7ICXDXFQjJ
CQPVyn2EVp78BPTZhqLi6CI7J036gI2XkJohE+6AjwKV2A9jMH0aOZdCVCbqWviUe3CR0EitB/0D
lyjl/9dbIhleWkhZSBlZh0U5ygXMW9/ipLo+SvQ5HRhdr2Qs5JFXRuCXr9nvfKzstpPOjrk+Pti4
a/1tppZNKWenrYlOHTDxpFv+6v6fdFhd3VhACKohYoawM2UxEUmaLGrGw6DmHtckzvkKxeuqyYXC
zp7WNg+UWouKRfj3ZrDs5uAnrzHCrl8bzS5MsFj047genvgbJoVCzjwaOOwYhQCX3u97RO/4oFx+
qf1oJGZEFM213k9V8tVKm/44r+EPruj92ykmCoKe/xmxUeDe/9P1DD9mCO+Znftuvy9gCyhidyKQ
zZXh68pgerEjuh/wq588ku6aIqe7wvFFc76LtUSRz2AhsezyDEBjPfEklnTK6kCrPWF+bQsuGeKl
wwD7fbaj2kUIDMEQRooIpJUqWu6lbV1P5N4Dzwc+BtK33iKW+t1ux+4YLjYQYeyF0ZmF7CitfAgu
oyI8aJTHPYoM24LeXbQfBcjaFmx52gzf54oryCveWQ9V70UHVz9oIssIWoxecyA/++XVu5T2vRgl
hfqXLlXYsPQdDARdomqcBJR7QMnDCY/3owoaeYge8ajZ1kHrFHhnbEWh48IKxH9pnrTz4GrDqt38
JyLnc3cwgFsJQujbhaPoQxXHsEAxYojee7EYzfkwvtSE96r+/1ZCDa7rXy/tfRjn7Cz8qm7f/WTN
T+lwOPd2eGTjR44TqK1Fg0bmWBy7pq0pTGuSxhdn/nSUdwd0vUf3sNHuHVH7m5gWfnfN0FQKHpmz
+kIgzNbkxOh3/ghoUS20qlQ3rK2KvvOPNrzCb8uWXrmaq2PlZSyzqK0Fe8rMj5T52zl1W4qAo8l+
dNkbPm5MOaKJd1beNaaGwNd8OxeIJpbPoCqMlM19feDfoIISBDNf9d+sJqtZuDpf3PlQ5nmt+/ro
wAiWp0yaQ/JwVmt3tn7myVvpax3JkugjHYREOu6PZDu9ifVcn+HIXuNQQSbOlhfk1KXDD1QMw/BZ
XADhdneU4z7JISAP6jyq6T/YSxqNtyjk3qWrZfo/JdhAxKlPMpyX8/uP2qNb7F6AaNoI9icBcB5P
HuL0dtooT8Fl4KXNbFW49dkgsdOliANwumdbGTLn5ZvEWe3cJR2tuxTeRZDLlbYLBklXoTH5ADT9
Lro+Dc5zD2FwrDObXCwCz3MV/4y74oZBKgWQTX/zBBk1PI0rJpdQB416A6WMMqTfNiIebwHSwbE8
eEcTjHYB6SBnbx9bu4fKT8vBokVX+JGIuP8QzW7KcoNvUoGAol/hj4aRgvI9J1JrPLsNt2sS9ffg
FoYrrbVdGVZX0r4HGuR+IJgJfi5zkEJhn2cqPvsRSX1atxq3ZAD7S+g8SUDjC+qNO1jzc25NaVG3
3otTmhUp+svriqS/MQrdTu/hLOJdS8bCGjZKR/GmPkgGhC0Uzra0V8n2Dwfwfemgyu/CKSDTFoZR
2AATyZCQ6sM9R6aOINz+n/LbjCKofjEJXkhEixItL8I6j2mfW4TgxAV1tLhwL6HAe5btYp9vqQWS
tNj/U1IA9BDpCuwZTqhC5DtJisTftD4t//0spfX50NKHsZMTktlizcglZApM1Cv58+eq0V/O4zhh
eJrAIfFAAh/apMAZkjEpysW5AZKFCS/pReUPc6NDoLRmsBaBd5tnQb/ieNfYDuwcH0gknYMhSy+i
FnhPYrsNvPfjYUnz0agcLa8xICsLCUx8nDiahf+MnEXa03Zpj0ib5gjzBUc1oNdami3mHH7/eoru
GHPCqKGkcKqfAUIzrp87POGGJojd8kUuxUWlXz9P0JTqETPyXOfqvrcdtwPPR58/PlN5N/d7b+ch
uhEhiaoxc0ic9XY8eGZCgIA+bmFqEDUpgIPne3PzGQvib1qghzkhkmrtpOwmwnF41xTq9Uvq7akz
/Ez6/vm4yjQpOB22FJR2rTmbE259Bw8SM5jzndx481A7Dgq9Lg7HAX8F0MkVeFP7XkrXhLS8Yqha
cn1ggj/v0f3e58oSymLoF9b1kFXVeaz8v53ENjjw/MjMPmDsl+4b90XbaEXroe8fO3qirVkO5hEe
m7Sz5GFt64pOL9YOLBauVkhSezi97J3vJqWyam8R87yh6z8Lz3BCPPA860InI/KnDUHISOeSBh48
Cx3FWxeMNzc6F/BM+Df17mbBhBP7q9/Yiw3Q5UPkXZM4SToTY392PadWXuP1aHZDHRvC2uzsqjyE
VBtSYTWW5tEHhT5tF4pVH76DeBv6AEEMEBra4HoU5yTyhyQ6YPG6X4klDeU8rhpS/ad1x4wG5Vg3
gzzst+9/n/BKkckXhgNNHtC+z31tSIOcOXTKd/PmSYOdk9GgQ18JfEoZUKWKu/XwvEOXEWdfjszX
AfdmwjvpY79Zc23lODulsFTPx3ps+KWyEXfq3LYC62ftgA5nKhJUeyylNiknAv1DswQViznWD1qd
CZmjbklluA5cWdEX40IBZkYrQj8/TrpiNHYwugqLRdCbSr0v+GYnXVlBGHSL21DZetND8YASpms/
BuqWYbxqnn6BTYgaRa8V21/Vp4Ul5EnXhPV/ssA2dVmk+NaoXF+sXbIJ7r52VDe1D+F4erD9GJHw
QH6lveCXXkR+82DoFXX8z+EpJbkeKiTrOMUMUwljiEiBRZMJMJ4TkjVTn2o3sQPx4viqKSBoukRq
O+m5s8bsEOlZeKKQUgAvWf8WEjaHJJav67Rqx2Au/Veprsm6w6HuokBg44dA9uMMTOLhtHnB2yg0
f2p2S1AA/ktupCfO6M7Upf8o11tZz3nlTEJtpzipE9jIQPucJssAqdLY3ozU2WzIBaQuywXHtbKu
/fqmCAVhv3kgIjJw5q2gR5CxhS5L1+xPnaQQmkd0UEyf3DO9koXLIfpesTM3KjN0sc/2D3XJpQkj
BhcIYPU0gHaKMqpEWPJjwm4ASJR1iTJdy+R84x+w7cdxiGTU1mwH7b9gf2MIjhHMKvSgQ/4dQx1l
XNh4SdG8XrpspkaOmiUOpVzyer9dxNQ6/zounSwMOrw3t1Ol/JIoLHVa/nZkC6br24N1D3x1D9Q3
RexYSFZ3q4BuyqCg/M8zKYVPbUlFAVKSi3JZyBHZcjZHY70dX6Efl7FrybN5x2O9l3KGjos1ITeL
PpXugKdl+WP5j1AUDVEHWAgDBmN/C/nHPceg/6ii9l+m7evxmplmN4CTabuxI3N/ck7dW2rKO836
1TAExKDDgijv0gcNr2Brhlh4JzVyNP+NeUQBN4Z1aBeo+meD/zwGHFAOnk3cnXYMdUO0oggKig/P
Sa5zoyRs+7eZ6EsNe8kguWiQrFRKtgQ8RKRoHawaPi3BqH3552C5gCJ7+RpgQMibV5BE1noAmVdI
mm7/N2QNQZUEIeblVJhqd+RZ6szZ2fbva6GVDcgbKjQcHSb3lWNFauQsX5QaU81qhlpzv3G+8W90
W5KI4MGH94yrPMts5LsHANx1cS8eLI3eWIQtjwZ1INPB3uRsTBHx3WH3JmlYAgZeFqUJZZhtIWy2
6Vqlem3pxSrYsELGmc95Xlql8Sd9zRRUTa8/1u4kuw26mNS6F5uUWcVinBqikIWYhINzfHEHmzhE
mvRvF2hrDCsYIhyy9dJNjOI054aSXRXFb1E98EoH3BcNAnwtawuTk2J+meEcSlEEQobG8H9o4VZI
Kry36uMRmDILWYzDR1e1IhaFi/4YcMJ5EjSI1Ygk5YCKudLqMUy8hd1TtsHpk2C3ZgZDJYcHPmks
kwDQyUFAjWxSwG7nSDG5nExqF63qtt84OfGO5efsr92HjKohslMOHyVzcqqbpTqgvTTbhX9yxShH
yL96LSoVw9A2fZXErs+Kr1PU7n58tZFZn7elJWbZI6evSSrIrVTQue4pizEXh7/T+wamQtn27pKI
krLRlu/f92tKvPBRxy0aAkX8zFgnIRTVaAQtn3ksaabHohrCwhRwtym2WkdJ+wRPw5CJqFX9yrUw
HAAt4baZpBMeqkatGu8E5THgrXrTTIS01MnhRtJcXIgmzVUTl/Tf5n64K0Nl5M8nKhyGABd0Fiy7
83IoME6sVKeL43f//DG0yXBuevn5DlkXF/eiCxICPd5R9icnJKgcy5bA2cf1q2nr++/6+Qu20fEI
JihACni8EyNFuT53bRj0xh4+KWZLZJK4xSfjiLCKiZ+UepAf6oRZ/byEj/ehClRs4VUZTreuvc4N
7beBys+rHE81w0MmH4+WRExeCXXAFu6nD5kREJWoaZCFuFBHhrnsSKyq5L2ijEYShJ5wcquUb8Ta
wdhNBMxrevuUiNGYmgVpjr16Q1bFi0V+k7s7gGR4oKQTC2SGcfp20nWdTQ/7EVS7I03Lndxh3C0D
yKF6Hi5chjHStcopcLJCV3FaRs64RIvjmtAmwecFSjo4n9KYAmljO2Qlro11XEg5qk/v2J2iy1m1
igBv5tl2aanzjZ44+4ksCrkcUgaV1tzFJKEhSdbmhe90YhzZH6q0FQpS34WA9LIXHAy7ncvZ09eC
OGRBpByrJ7V5RDnClH2jAkdCa7IbsjAwcbuMAWU4lF74Tu+5aNeDPHpRWkI+yRl9Hudi3DUyJc6u
/QL76b3C3XumNua8O1TWL9ps728QwI7FJ0fMKiob0NYO7LWyHLg2mr80xwbpludrWyqCAlI5NiTy
BWvoAHJp0HFoSybNV8PRGjFIHHHPqDgv8MFyOZX/b22VWE9G7jIBOvkqMSe0fm+mK2+vV6SZhJFK
n3HBrC2nEIt3Jc9VGO6nofxaWT2OhThKw90t5v7hhMdjsmSKpkkDjyThGz4kE1Q8eJhW/onPPHk2
bWlB1B/XuU+Jz0Xxv//9o4acdz2U/z83VAETrzxrLLVBeK46Hpi+evfEm3ncE6puj5l+pYv2Q47k
tayA3UlYGtZN4PeUvOxfbyagBNQFbHPZLR9CV11PplrxSRVSRbbCnCJ4GMTIDdwwDFyqmDPoGwuH
HQ51R3ulFfNGBYi4i+K8Vv9/BhpsL25znSNIGrbWb2dvRsCBFajlecMV5QBotGz3xgND2LfLaFX1
IgGPAemrbmI3Fyeos6tjxrwHAWFS9/1e/RD6uJmk+8QinUH6EmuFovtLecPxx55CYXtyJCbaaM29
ep0RbBhWcgpdn9E+qHfHu7KJj/u5J3amW2NVz2xPfLDvTiXYEjcXrISKPblcwfKtUW3x1c/t/4EG
S5bR1HLIV6tFmAjkTL9myfGdMxP5Dwz0PwAIww3nIFUQ+vc1ApzR2K+6GqKEWRPzhp3U3Bk87K8x
8tBUU9JtfGz+08Y0YoE8rombLMrj0mih+v73i9N/Tbiko6EdXWaWt7iRL5gsv9wnv1KcZm3otKD0
G9BxxuZdG2cj8x7alNU3PGG4q1zC076aUVeT6s0U37Z2NqGuN6FxwcG91Jp2lFXm3JUHfM5PTda/
hDVnIwdlPFwGqKUfoRikuN9OlI/QDrWpDQgwCuXhp/juuQzVnM5jrPhe4p9la9m94gvHBLyHcgZI
Yni2zBVdUMgL3q6Z+/sqxNSDX79F5xH5eiXP6FnwLp/LzLPFSeAuZccPMRWWgUBsR7x2Vcwajb+2
7c+o9vvA99kk7EG861BZ/b328N5uI5iWmYr48oKOlK01NH7VS8qfv+hXYzaD2lifd2wqYJ4jrAqp
FmO/12D9DEWM4Nwquk94PDAVR5hpV3KxCFuRK0Y41yjiVmLjkhoZXKA6u7tzBe2FDQ61lpizQUhN
ZBuZdXWcIW8uigZIOIHSKakyZTa8qEQoXh01btlvQD73EhHRjfe5MFMWIaktfZxOkgnmC03WYX4l
cR+DUleThpLnHb9xpj/SXrV5OqConxq15hHWPPty3z+41pKTiXyKMFQAGUlJFmoHeu5RnljuQV0W
hox6EbA4WZtZz4oGriQgcbiuz2HzH2JEIyKqTUPrsStTn4cxcgFI00OKoGxeoIUqdhPGI95GPJyS
piHWjeEbLyMF+N8I2V/BPNtHLfXxdlZItaVCDxl2jS3JDoADqyyQrIl5HiUs+wySOBRh0DdeV5GS
4apzc7Qiyx8jfWhjYbTAUAhWhy0eLwrpmakHdOgnXRoEl7GkYUpht3bL64t92d0S4SZMMhQOxtT9
Vve78RCbouMdEvGeGrS4tNHiw0ABezO2a9J47WPIIsdKGldc0sYfplQ2ofY1R3r0saWLRFLgLc2K
0+CAOCUcfgzGh26lrEL/xMM9PX+xkS8/gYHLgWr+H6TQepp6qofwrOn1F5FviwmR/pMt6slmNx+r
l404AdEpVCF8E+6qzYOmjZC9B10g3EKmY5yY9eqORbZey8j4yU7cNN6meAlkJTLcp1xp675VDgO0
OrH/bAELgv5DvIIWzQSYr1Z96aggqYOT0ZHtshk4fjqnYASF2gtFWXK2rdkQiU75n0EvvyktQZpi
7QxuQofNdvhGD07MDw/afZbky9hZ84xBgH4X4itBybdmDNah7dPWtkZPN5saT2SUmEgTIvzP6ac5
5+rWrYMGUEWvB0Yz0bIh111Yh/rrdIlB0gENjms5m08ZCvzI+vQi3Dl866i/0p+J1pht16Y7mq2C
nCJSUoQk9OaHFOvXF6EROWR3tUYYR+Dv+echNie+671J+0/+V0eNyx3IdqJFp7+ZltezLunhvG3L
lu55UZeS4UZSE69tgZeuRZjUyVXEiZOhPUUXEyfl6vDy3VKCj+GxGeds/SIn28POZAqbhQ+vEv51
YLG2+KTbof7aON85ODXgsOVPJPuG7y/3TeLitLNgZoHkIWtFs7S++o/qILdvunD6k9kEU+h3c3/J
P2VjFrZoGq/DZ1V30MVSLv5pHp0W25Xe17Xh5X2fFICxE9WUAIdUJBFB/G8QYvGHtLWNwaXomqsC
gTqmcC5yPiw2V8GrLZObDMHgtlT/NlG9lLNV/kYlbhLqzt+iX9m7ilHstr80Efq3e5sLlpjBNhJO
tjbAfzkATWsoM/0y3HX0+d/+gxXgYydSs18qaxAV1Nt6K6+vCqDaG3K22NpN4Zk3M9kpcFgf1bTX
r+mrKu1cqRH4ZYcP3jwp3QudvGjiJiaprRjAMRcVhM3OPYcT7zrbCM8eyiglXjNV8odjJY4ZPn7g
mvRd3ECnIbp9qFqFeCsUXVbE/uJplTjLyJWcppQuzraqaXydgkbwuKJVad4XzbTpnhPeFYCPWaSG
/gXjUr15ZaTHTlBYB422KYNH0qXohisepHMFiCS2UxwYclLGmuIoLAi+9P8bw/KHSSAQFimCk9dO
0mfqaLMTxbNyMtE4iDlON2dGKcGUbkP/sYeQn/NlmxXlddxX+dz6Vc2mL/1CDWGuaiIweYOdouKP
wSDXHgYt/iXvuCJb3/tgPRWpNbzzSCCXllO9UB3MzDBqiIXQ0em+0bPHun4mOVAvOAUxX/mwkrxn
i2OUvYa1mlQGZOs6wkiBcAU5hjJMQAkKmLLdoc7HOxzSE84D+EMDvxJyDYmVwbCeAb6vSetqowe5
RvdYcOo2/VeLVJO1xxAKlVKkBLTVxS2mjzYtVI2+1kyesHxgUOZuoJv05hSrSBGNZ6IN9LmJ08Og
6OnNMcWqn8BbBD2wShpEyfa+JO1x3BSJRakVsffAz9J/RPrnhQX/gpnG9W9EFDXz3yDE2BL+jPTV
/zit5Y4HKxXeJkTrmlzNeCWgjpDwIUAMo2pgrQ2myCNXfqNqDtKbf4cP68GV/3GU2cJjTSnar0Pg
WZ7l30F2QFIGH7BS+v9c6lGp8fNjuoQna2h2F4b1SZMuOgmJUIBj62YBDWPmG4rPMz08IxbL0OyN
MCLtUabEk1jgCNB1t43Tqp/ROnNOzesRrJ7ZDCInLBW5sknAaBBXz/GMga8eG44fz4Xa49+uoY57
a+fZOqrf0wCYUeSkSR644F/etH/f/LWho3qB9efIsdTQscOUw68UJXH6Rhq2/OTxRRDUwjW5omW6
dZiyfzaeaNGnnWa9zDYdqRE056XjPJuIeLG84C2BK90z02FbaGRWPNcxYwPqae/v8Sxnvcx9Je++
fqCNqtV9ZSfdi/WTXtGQXDHqppCt2SqwfLiXOi35MaE9uSdkiINv/yVzBwvf8W8HfEKHUEJW3MzG
4/7kYlrDqxMfXYjn1KGATCzb4v4RmJgbRLJubZseBuQ/4W4zHsaCQr40okLxmeGrt4I9kpit0mL6
T+4ldFqJki7tGmLlRlwxNSkg74kv0+ttlB502rT6QCaBhQKdQerf4erPJGyjlAq4ehj0QulvajL5
pXp+K0dRN3Mj8oSI6mHq9mm2PIGNSK4pxWMKWzE1QIVwuBzkC1gUaCqJIebPVL2wfPankomOCXnu
yiAi8m9ox06wmSUKIwQlvNYXEsnabXPHD8U/nkLp0h4ZATkRnSfgpyQY+EK3WpBtktqX4zlmuJu9
mFYMZiOO/OMV3UM5QhO4PXIiy7PpHCpBoPmbcFqPNr46XtDKV/YAjtddNXe2m+q8Dwx9bsplZjEa
qEj/T2/nu7cFQs1VzGRiiADy3PytW1fBWeid+wVj+nAL+OkyFKV0SQqcIPi78yEzTJsIZ82Y114+
RtGmAUhY8+yD1K9msvfrBqqJPZtbePXInE+FfP9GS2M7nK+E8gGOuGSzHFwUHqVQs8PMiyO008Pz
XAb/kSH5Oa33mwcvIMn8XuFn3vYgUz00ElGM2U9Scsxrp9xlIPWpZzBmOJ7kFlJccaroohg00znC
WwtepYrpg3yDklXXPXL8EuGT6+hrxAH/k3QGFaSRTwX/Ysg8W6aDhgrwPxZvG7f11A7D8mNq48nN
1g9ekoR0bBSw0QPwaIGO+IrCFNsG+Tewz527lMeF5REGLFYVrGyUbNOLs5j4V5by9JAOUuCGLZeG
R6hNc8U4T89xQYdJfzuwaK0e+dBzz32hAMLanRtNx2RPevJMb2Xm6voiyq/UjXScN+/8N2wEMiVt
ex9aMHDHr+C8SyAss/iF04fpNup5TDPxzy5ghkfy5dXhLWSz/c4zvHDZXLro6wchdK292cLtmIEC
GRTRNernzGUEK3x9hShm7cVyh46vZfaaAoWeYHZGhgZYLA+pMWY+QyCbnCWtMayVBrUblLB4JiG0
w3krckVbs4+iOH0a1WsODDYEk8MXAqqg/0XRgFyiEJI4PbLFxxN47auGKu4BT7M1O2Lmtc4m/WNK
TnQftVOLxEj+kOWepMiwugIvK+ePc2gIwPLNt/115y7JgNuJytIEiUkkY6DHS77mf8MvLIT0NVZT
7ijsNACCUhQKFv8h+4z37rpKlgTL9byqePAjZPHIhcvSwaQmHFyyg5dkexi2RBlhxED2KoIvH8xq
XUMqnGI0mZWH41sZRfx9ItpxpI4WYXX3KPJEMgUks4GjerAdamuLMwrgiD5vLmBvvmgQ3G87mS0i
jNw+LLIa/p9E8CKhYTjJg7ihIy1DyX7+r7UQWhqFzE1H4JDEyUdyy2L9mqDBs/eZKWgRFg2BdakO
s6Yus+8DqhpMFFU12bbQjxd9nCz8R/9Acx5lOdSGk827GVtdjsBfJWS2yM74dk31MC76fJW8gX89
x0Ei7/zpxXNRb4qgUb76XF8cM4G8ObQy7UKYUUh9V99Fn/ZevROtqGJxoH09yU3pMyL5rQlDHiC8
ErIV1PuOR4tn54Gp0j+46SivvQKdmbb/Q1TjoIRwq3EdAoNByrTM0PiZEXgN2U8OvpPCDcNxHp3d
0aL61uFKK83gdaAdbS4hD62t/LQlxhaM+Hb4NKQM/FwTYWNgG+ssvO7rdhCyMbuyz2fV3POY1LB+
AeCRLbr6PXrNs9kHCAz7bRMNGl21U0UaxmD/V6t9Qvevur1olKC0g6zOGkxI+5U63ooMc8r/N73m
BDaRBVnFjmbS8GvqNTVcBmub93UbApAd2vi2WqCGEQSLVUK19xc9c8D1mrcWG96UN1iBA42eoVHe
pYBlsxa+nLrb/ICPyEfDjmb9MaWCvLdVFoQfzTidkGYJeqMg4AlDULpCyOLotMldCvcnBygmJQgV
Iq+z4im8n8pmnj4PpDTSlZw3OgScB7BKVeUtnQPosAe+ciGR6eSnZsX4kDyDEP4e613jlSsHOSC3
+YVGrqIbPQnZ/21PfYo6fvM9C4mGKXdyGkBxtmoBifQ5kwOvuzr1VcJfwrB/9RjwZfECYSiXsItb
I+bq93Xl85FUCiTZnise85IGSgYa8vAbhjo85xhu/OECGsutC0Tiy7oj1JRJY4ceUQzsQH9d8/pz
Vvx7p1UHC74B3yFZMof8v22gwhnMUbXWNeALdk+XqxPQ1STctH8tMRYhuQF6OQ7shu2tBYILjKJz
xwLpv05twxdtOGwm8RTd+nQN8HaQYJwpV6xHA/0akg/sCtIhn2N4VxK5efwEgqp7Rslpajhby8Hh
0A65HcyR7yZ2yRk49Q8ymIUYODv0mKlDePpQftInxjw1VqFNTbxWK9RSrp5gfp0GpDGcI3s9128/
G8UgxoJekQZ0HU7Ad0NlIm9g4nb7holiRVkCLkmQ3n6kbBMgcZPp+ChdBHgYj2Z/IMmhNnYEHWAA
lmcxYeVMvWq7DsBgRkphjTMVxCm3U/M6KYWKewGX9kAvoYXHC+P/EltKYV3X1tdMYR01F3PXubxT
4bhKI271yVq26Cqiuq6/xxix2JTrdbpaO41e9sJxS0mOCcbZYvYJOxhyyvFMU16OUfn+vwKWV4Sl
37q0ah7mE1jOkHCvlhHxHhPVLIezqotaPy+KW5jQBgacOsOn2r8plc71ETQBAwPAunpdieVlONWf
3mZywWbApu2D+WBOLxlF5FndkF5rLoIZI4nExfWxRNpt6eWazK2sFwrHqnOHlI582fHTDMqvJN/H
7iIBW8ROfBdkaneuD934KOXaHgQWOwHQ6HEwVqUi2uck06Q7p2PvqzEL7PfqBvT1wFW7NWH8b+4C
TfPIFZqft59kqW3dPx+Hra1A2hEJkvfFv1oJm58l9E4DaimSflQsxpr+/7uSChHGLIA6PsmFGwOc
tASHS4GV2Pfz0iMz65PPP+iq5uAzYsFg/9p05j+Ubr96EotPtYiCuObedmXeIe1nHS7aN+fd9cZW
TBNBL9K7+Qlj81S04YMmLGnhY6i640nx/FE6l7hLi96mHYXt8R82ojIxKa2HPLZ4/WB4FoGKULMq
sluF/TX3uWx5fyd8lfYsocDyuikaI9kJmEQ3hmwf3DMaUs2n3PcfLjOurZKjhxLYhiUH3Td2torF
IjC5Kd/2yUhdEpmymap2IyznWyaKFwaKQC/gYR1lhNqrvlFaWJZOqVlioRtJPYabayRtQwISMNP0
pvHKB8t48lv85oYgU3WggVZgiFgYgfuiqZKZgAHyeuxiKWY50OC7ZiSRHv7D+tEUWeHPA9CVQQOV
QRkHb0XP3LHYJ1gTH8vkhdxA2Lcs0MQCJxWJ/5KaEw5g4uRrgg9jH2jknnhPKrXNLCdKYaV34Zo2
QLwrY+oR0doMtEk0j05nV7r1C3D4RheIe0hmQOLGe1pmbuInbLfc4BiJA9SXoPlJxi3I5GA6z07V
WEWQHX8/YjCxo6f3H2q9Rq2eXc8uFtLsMOaoxB/f4i2MCauqr6vO/h1BkSH4AEn3WWzcsjIcQUiU
cFfciSG4WHlX9lkCbdc6BUV4pwwcFYekjXABjlgTOeiUgwqCaKnV298HZ57/xyCLz9ll85nueci8
kzFYUkQexGYuDqIKBMLCCokKcysywXqQBeiRSNiTeEl0b8QVvIuNCHVZ0w0EwRHG0tGmhu/MnaVp
GPNzvEWi1GSEkaKg2epRdlLB2MS/e4I4APyIlb9Jo9eszhOBeYJIenYzq1YL2cI8Nqil6+H0YJKf
68xGzaTQ9Ocx4MJ49EgaD1b1aWxABi05VBb/zIKb5K+EgCyvz+yMEd/lslkw325cfgi0ya/8dvAD
0bySe25ZxpdIOu/szdL4f/qwelG3PWbUcioN3iEtah22fCtOdruVKKQdZiTY6XOHWLhNnr1dEh/N
O9mZH9oxtKqXoQwOUgOVdt+wIUmJbDHORNhk4MIXEkbd3NOoU3dyI4JVXXx273DXRFM2IDPDXSYa
XyLqBKCA3XV+mJXedlQOaBEtOLupkLvmRVTQhhgJosOkhUkPfv+3GupQ7C4KzVQ93SR6uHSoglWV
9+hi4VHuGrY1d2FGs3gTASl+v2CWtcWTumhBy2crH95qmejDlNxlLySY8o9BN+Pnr5/PBLBoji3v
pB16nu02JWqFM086XB6FaT5Aza5xxUggt7VSlfgbsbJoE/mV72N3jjwKZsDn1al9rF3Wug728hyQ
FEGFpSkUnghaAnkux/n8KI7bO6HXgMw08LMWls4xFFQl3Pu37Px9jBLFKdjJjKGc7r3aiBDSPyhY
8ygrkt+byKypJFeDecVN73WJzQzNBgYtTS62i9/0pbj+JtCDU7oybblJoZr8UoQEjEuByXCdy1F7
rC+eeza5M8R5c2MtwoJ8pwv55ac2btp48JhtyKcPWDQWIRX1yApM2i4zf+XWAwi+v3D7ucIz1bcd
vtiEUbXprgDeizMS7Q1wFriWHhWXDR5n4FlGgkHqW0Jc8O705Wlz+Zi3+yIDZIXlGviHGvAa6OHN
cWrg8RhAGuP+Nxpc2M1A8xWzBZbTsPjFolN1pabiMap9uuo+ZwxvnGpuYDvB2a8enuP6K3YOTk+f
z9XWhtnrSTuayu+xZpJSQVRl7dxgvksX5NRAy+n+6usXt1H3C0i6SIxMrZiygi2ciM98LHJ3f/Ai
CvU8Cje5GQIWQY0QH+DMUhMeIWtFaY34Ec05dcn2OuA13zsqQDqx5Lnuz+JCsW0iX79oV5Oy7XO0
AEFBzFmGZlyt37qNjwuvRsame9ngXpFwzFNHaUZLYCGlkUiFjs649u82OXGOZTxFqDe4L2jR4zBF
P0stD6yngz4ff5lAefZLCbF9QfWFo4Mr8iGBj0KP/aO2LvZyyIaF1mBGsMs4ALTUDhKiUXoS+Gba
I2TuVCnG9V4u3Sdpbbmlkoz9sDcpgg9kDWD8YDA9aNisuSzrcikvG0z3SaeH2NVaw2NL98+IOmDw
cByHli4SbUNOdwgUV7PA8ZOz4JIXTqWjzrUR4lPiVDYKfaDloVQDcylQLR8XKJ1Vr2PGvyTpPX9X
NukOPAkIpUdzuZGIstcCJx4RYT5/G1uyWIbwRz5uFNIxaB1H/euL27tuEWK7+2f8M3P1PCdZNUg3
apQgZRb0PjIOyfnAm6zVjeSiKm39HiKh4OF/wRkmI+pMtdtSAAbUAEzFbW73bSIfjVi4iCTp+7WY
RlgbU9DkQRGXFSYTkVFtQAgK1Yk33aI8Qz/FhGspkbVfj+sDFPkAEUG70jnw3WuyJqc58qQaEzgF
NU1cWRAAr1FuPaG3y5V0LvxnSqdv0Lm9sKJyLU3xsBLYWTRhuSEZLLyJdItH7MMNw/4wRL/ZDmJJ
FYYLSmRQfTE6BO3Qs3nJSI2oZf0yyj5ETPRrBSy5KPC5/GaHKLBafzfR+exuv9jkGelF3V9Oczjw
TlerjJsOsSpO/FLGSemZE+L+l6Cwggg0gXPp4ugrbg8uipT8UBBJFY1XDU59eBMYJb3UAGdyoVd1
Hr8nx6l88rI9gGyHURmA5lv/DIZJ4VsowUOhOl4dzmAkAQvMbiVVKQvS53ULBxNnKCJlgHjqhb02
XdHmO/2ZAJ4wPUd1k52p1PCQK3ThwIaKXvgmqXXHJUrqDGRjkaDhcJYXIGKc9RtJE0r3Km8ie9CB
Ke9y+cd4ryRmvdPSXF3x6TpAGVLDcQqjn8/oNZs0sWH+YfVfKvTHKao6EEoYK+9XkNJatnZl03Iu
S1iVQAssLvSiYPmkxnKRN9mgcDHVpMHvqO34G8Fqk0c53PixnQ5s6ZGzpbqgZVCoInFouECy7IeT
hEMe5uvKQccm3DJ3Mi2doVct/AZUug0ZnRBZSXwucNfMu9KvME+9xmlTx5A1FM+Fb2dp+Ft+uQmb
UADiN6jyfvrSjEge6RbJS+VdG4Z+NDi/YDRMSNEYL+FQSyQ97b/uMmhUZPo2yqZweir1vWgYKCGd
QBq6Sriytc7S7N5Nfwn8LdmIbfh4ED7Q7WFl9H7TQqrxXW8YXGaMCL6gjhdEymM0pc/4/bePvgMz
mHgmonmONN1Vch5t0BJz85f6m3ftUWNXlHmGRNhGXXClH8MuncQ6r8pKKoe9c2oVrVfY34UYocKf
Lr2vuscGQNMkudI9Bwqmzr/d4ZDrPP0HQM40Sy4cmkOt4O/Hg5ByPE8DJEAXhBYkqQQqgyuFVh5g
AeecKQHZUBkXpCRhPxgjrVy9DFkkSSvArxPo0a7AHIlcwRu3oAxgRQ64om1Tnby8U1l+yTXslVnw
o+8fZE+ZNTaAGsdjOEfLd4VPXWMgjj41PtMuKVvaFlrLAM2b7yhVICrsbqWOt/hC4mqx7jeaYKnJ
avy/izjfOuvtAk1aviOQX2VH+9CJ3LV6Nu5mMVAw8pNoZg10CsUji1VcKIlE+QmL79bLDUEzrd4b
L/GdW5NEYv2tVqGatijDOO3NJlKocAFeIDojrTONk8EMU5393R59wfbRPdbRm13FaYNtyzSwF3bI
7Bh7CZN/7ctHhc/rNxGshyeensbmVtivuat+U62+HnX7WHycKfJu8CaSUNIJ+FJ6xifid9FkNSD+
u/a65OYUWgkmTFYudcXpDMvhSRXcRk7bPzBB2KIzK9F7oVk7H6x2xCUsrX6rvhC7vCvd2TqRcpFa
AhxMiYggopZxPP9IUQdpjQbR4bjalUc0ahpj+GkiFZgdcEK4e1tmIdLnFC/0/A+Z5cTkQhw/wmEp
+PrREIkATy09za4Fzb+Fu3t/LBAR8SYEBe3GlT+6I31bj/RteXs1LZAsI/+uIxKrSks+8eLRDxuM
QtgMeLDwvQLhS0iXONSlLBZyhcKuIGHlp1jv8A3hXpAv2pu5Yo4dlirEYrf2f2aOnViCetBzpQ4O
9XlbjnO5pPdNbnRLY7lDK9PcbTCMJy+8b2vUSFbVFy/Ok2qf+RrlbsbfWS4/GehDpQ81Gxh7add4
dEH09/257GNL+WpKp7ITdYyclkMcxImWzrgUILzcGc4preQOiLR7dQVQe3kM4CiLEuFagQk4xW3+
LoT/UD4QBIxXfYK6dAdbApJ+/tJzesU89/qhRG7YCP3+pkRBPJw8oVs+vUFBROvfH4HM/9otdLsu
mzcN+GwcBNu67eXZZ+FzBbYuaPfCJ4gZSNPlhpfJYkb3R9Vu/OEEUgKUR2XHiDhxZnyHczO5F5WN
o2KQnR+HyvaZlktxAZkBILN8ZqREpFDtqhzhIgZD2MkFjuF09nLMSLIC60b6Fuqm//c7aHka99mF
8miz1g8ErZyRuZpdXLHoqxE9YxqPDe13doWhLFqzJAxUCtPdjdy2SYARK376ry9g+YZRWBsv1rZN
vIjBi5jS0xJYiiQ31jyjOAlJHd5jFZe4mSnhDg2Zc5M5Li5lDX6FIXbDRjD4e26c1HRq1svbdTVe
f5jeGDyfWJ6hBInZtN9CkRAk9PhwIe7hcnhpVtweESweLBAovhNmHVOUO4luY8LZofn9H4AKADRD
zQHt8XJwkcd+R8W+UXXuFFQgwXzxse18xncAR9M60z5e7CeC0MgTk31rHbmVGHs0zPQbMYzhnBEc
tlY2O0LMCxn6OkBJzD0srPhXKp71V6EsJqyLpUBKbflTQKUUON3CMxNSf748qMSpzmF5Y+daV+lG
voyrQNiun/klwEsBN4EEhRqxVpl6iUAzmxl444a3vlMvJwxLTwWx5mTc9DE51dgWncBPuRXsN9Ee
XtHW6St9wdyH/dSpCe8S+gtixE3EAIPdRTsJl83pUVwrrR/d9jIP7x5Ss8RT2AoUO8S65Ixsx5tj
J9hjEw22K4b806MXDT8wK8neDrooiVqwSOJs35APSxEAGho3pWpgxt2hcQVRSJJkMef/+HHRtyHO
lRywqsX25sVJGJj1iOyQ9NCNimgD3jBqT0Rgn1DSP+DgrkF8vI7a0mn7H+QCJS2m9UfphWpcVXZU
pyeFPc9G6QSo/T7C39HBS3/7/lEZia9hgjSwldsZ7oClADNdA1qMvJ/jjtGR9dwAfwTwwIVqXtk5
vJFSssJov27WUUE02OqeAl60A5jfwGTpXdkVvtqQckJyF5ebf2M9XsIqHcZIfqpoerYKE+ak5iwl
rpEYEJ6EUI9690otUV5ckotlB3vvJWdbiCZeOVzxkbQDGL3DFiPqQE3JNwwqjU/4FE4dKxmJ8gPf
W8mZtZMIpavgWGaLq/t/g+jM671CrmIfX0dcaczosJ6wCwOhBEw1aA11drTpy/GwdZmFz5k2YU6/
TC8HohibFQFnmUPUXcg+KHqU1ZfVC34+Ef8EAUQjx/t2nEohHNloa6cLjxdLCSHCAvab4M9Vb5U0
ZzOwz2rk6bdE6SeBPvOZzee5Llqxv5qvQ2YEPErnKLc02HDI3F5WtodKqM+7hzO5SKSrfhKon0p/
Q826UvVGbppFQU+W/1eI/LGuqt9Gg/TT5cQlJGAePc2bzVRP4luuj7klLqGcUlwi3sdFjxi/8TtH
lnYcQbpXyWw3atEZsXp7qwaKlpbLiIkA1J6fXCxmplwMWEb6o9HhKR913clYDgTbEmZ+B6UtQqkG
WNimkO9x7nz30UBoCxpd0lJpuhQNhF0Y/d77E4ecOo9ht57YM1vJxKJuYQ1RimXh5ZOBQtMwoVfs
/J30+7r2/QD8c9+OY1gA4VRh6LFQx4FS0JWCqlKSMWHkFSeq1NinItF2hXLphP/vHaRLwilb4tQu
jjzZDwz0lwbfMBm4Xrarg74EeSn454/T48c4J9072lNONwScbm/ja9wV73391CvvxpUhd6ggULtT
wJj2ZhpKTQQxAIlYZvJgFhAZybi9J/MPafVD+tSCh1NBLM7mJVLazbVdRUr/TgJRwHJSYXCh4fxQ
IL3sj+XW/U3eTbxec1LZnX9cCshUy283V0dnaLEB8Y/HmVOueE7Dq/s3O2qWkgbai6JOS0Bhzm50
ucsQ+OC7LhMIMqNlAC9KdFVbHhJK0b1Z4Ex9df0xncu5Vj4xurQ3ohQ/KbekZq3P7wng3QlMWh5m
fmd6IE4BFyG3nu5FhNXSKQ2h+e2dYa/oQU4Q9UMs7EZksmW8prP68DJ3M7pFmuLxzJl0x0pbG7e2
p7DthAqEn+79PVv60UsbT3cbeA2h6JB+s6odUKdsdi4YO3sP/F0/9VKWZczv8YfelA+ocVljad9B
hju0WYJ/igYwCn7vzdDrQpveb8PcMO0O0pZKeg6SKPUkw1O9z+avi/qevS5A7t1cB7Jt5JtY+mB4
iwaI4iQoNtx3dHCtUipaI5qA4TawqiH4hNS7agNcgc4WrNsJwks8T7aiOsGHKKsLI282xLmjg1ng
OLB7Mi4bTX3ru383iB6xjs0gSE5/8QiEG2X2MkKd+rtarGFRHO5rLUks2wHXF9gFjTy3NL5qWmP3
6jjr8bKhb3oBFSRsYnxVQLMEKnAFHz+vk6B1iNcYeSg94Q5e/dqSmP4Q9hwJXC49Hgu14r14Pcns
wzVWRke7OAs6z6fwla11uZvCJl7ISscumRVnBA4KDyEfAfeHPl9OhRu2leM1qzO/NmlS9oDpOwIN
S8u8J8Tbv7K6S4QgS0wsrqex1g4jAD+H/r/hnDj5KPdRAgzn9gHor03DPbvD117w2APE8Ns/EqFo
9CcNaF3ORgrwlUZnYYtOmy2YcUB1UjS5MehjQWlYhH8Jn8m4YB6WxTJmND3qUEWIfKmIF0oQkqsl
d/WUbE/Q+JEGyUzTIATVer3MEL4NK1fqnnN+pSOOF/tXkyFQ++9XUoz5zQTZrLAAEYdByFP0lw+U
Ktx2z/O36Lk/S+3YrJ5sd28VF21iDAiqPZWmFKKwwD3w1yEWyR+FMF/dcGB88YDWUQeAKWD6YgPl
YOHvsgUk8OKwaOPJ94YZi1skf9vhkcvrYLk+uViXFwYyF/5/cXsBfErf0A3iFfdDndw29WQkcm9d
S5z2izt2+93lHGTqZG+oMovP76s8f1LA4inijCo7iVIFT6yWIqhFX01BLxzinFYWYJXeSkBHUF1a
UK2MY93n8MiemBlI2Cz1qg6YGOVN56b3ElCOIz8FjhMz3MBzL9tdUbp2MU5oJOWcJtHAQQh0W1vj
wFrh9SmQaTOy2wSSD12+2YYJRanzYHHfhg5yHOTc7zO9nLgv40U9nXCfboqScrayWQKZkaOhpFcC
ysTuOdfgGeM9/n4J0gsZWmCPN3Eqm+qWeJKjVpzIun3IP2FCJWjFkBK6IWH0pUcmS1D9b7qETj6F
Uu4/b3XZfOo+ARpJjr4+brh1yvZXg//yCw6yeXyB0ulvzH9OA/t5EIw0GE1zbTs+VANh3n2bqq0y
7X87O3xUmOBr61ot38wR4diR6/2gXD/XaJIureAATkGAff1auMWgIpFBQ9DvejEy74CIYicfZvVR
K1MZL581npCPW8IhL2YYI0t5+RC2B5ZQDwaODfqbUebA0zDpy3IN8KjQjQSeyMqcIoluj50so255
kwrhT3ju4/z6kBgIvqQgNYC2Q1AXLWL0aqQVrP+vx7OoXQtsjiLX/d/h9028F3uW7Ny3AZK5RjX4
+SpHQZPzs4yZhd1ebTgRrQjxt9tVFS/vHM1sBpPZjqbKGP2iFQADUUi/3GAhQqUuDpjJ8hyepp0e
lJkQDiQiKfO71aXrBA4JPCP80Jih1ik/vGoUWylOmkOboLrCc3BaEhV7RL5Shyqe8+SNHWUU8ObF
pQY5N6EKDcuW6AD2qYWnbUyyETl4nDHxROHRqAO1JAiWy9q61Pm0QPD1reweTjdNA2htHir7dtAv
gIImNoO+fpDQIeOy9yNNLsG4fGmIE0xlYl1+FppWstYYJccMlvxug8rFDpr47mH/cIx8uvG0i2b+
1qMS6kkoAiEaG/czZ/TUz53IJpAPK5PQgGPKEEIzt0DHtPgYoLccH4bWr/Hym/IFZ/458GpRYz4d
4JAI723J4xRK/dma7wRqWCoBO34FS6vRtgU9LAeIlQRDnwTvtPPQNov7WyQqUbk2jxPqYcQ/bHy/
4JWL+foEGAZXdGsbL9nFWiFirYUZfizxNfgxE3eJKZi6qmoV6gENolLgwoV5BZ7wWFdArX5Cy5YV
mIfXAON7S8ADrv2KdHSwRR5OegxJcrh65BA3Ha9xGAiaqiVNLfxhdJczeg14M2lgr5lXJNIPpnFA
GhNbIRzda2mRZATOm9LkmQRCDlcQYxBnhshy1JHdtFBJjI57lT+gRh/9IdGE81Hh/RXvbuTN0GAP
utkGDQAwTREjr1lYsHOfCRbW9kNIleM39i7v9UPKqU/XAbsRck0b+NdLn0JAWvNvpvJk5EKRcRT1
pPSXM9WBuCP7BG3jRfBQFBUKShRXabij8xasONVhfW8woPMC8Ixw8Pb7w7ADf6kldWjc2Kb+eFc1
+zIPfN/YNymlOBZCrai+S+yYdmH9qyw1gWkCjc6URTNqsaVv7YfKaZMsnU5MziOWx8C1hj29j0rR
Xx5XItQUMsTkpYmbnBNmRxSPwY8lasaAeQYoBI+YZ9fDXIjLGyWe4UqKD+Fb0lGtnQ0RVLayZp0t
+Ev5yVpEB7zpm6uIu09CpLU63Ni5d2+3KbHfhqw9eR7GC8RwIwGjEZdkyoqCDWHoqxBL4W1ZntKM
fbehNOv2YW90gWWXXn67w2PVueVedL7hdxx79NayZvJ4+WmMM+Ce7FZz722rdHLmaKVJidgeuwWF
Sv6oUXUnuLt6EniGGoHo4jzcSKT+olQ+S6eNSTwJsGGwkMOrrR5Fr0Z9eEuf8OyuAPyvxuy/nbGE
MnW3i3ccb0pnuXyuSnTPR04+SnTPNMdxVCKaQdNTPExdam8OqbrY2sdNiOAPqg+QQ5zyjbNTIrip
GT6kkfDB4FE4qSBbSr9Q5w==
`protect end_protected
