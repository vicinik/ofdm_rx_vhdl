-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nR2HPib2VdYN2q+0jzGpR5zNOYFSqPISKIGnmXc5rVjV9dEJegWIXz50MeMYNuMAGH5fzjE8bZUW
PQl1sbOr2IPZaAEULgB/Ratkied0JOf/Y608oeZVWFbr0dYeDckuqYJqzhuVqgyDSi2Zf+kTqiWf
4j5aXYBe4zq1UEslhPScbyDBM8pNWdrY9qnFRHPO/8bH0MO4SugEktRkifzkfrV/BUV53L4tx9J8
TyaCUiTfCFmv+wLn9LPPAuxX5BVc8bQ0vfXq3ExlP2iA3wbeKqb90DljRLg+s/X/0aSHMiIA9BnL
I9eoC5l9z/hYZj8lBPePo8rdvDiIpGzLTv4X8A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 71328)
`protect data_block
3mInpbsnSBRdUS3aGpLC/QDwhH4zj8TdFrH/8hC3A/zrE0CzUL9HXtbdSHzoznT1YV23SPuYVwzv
uDIkyb15r3ywrJvqYpyrgYocY8KRG2M4KnWQQsdAatNXoP8q9bOd5q1phPFX0ZY46Q3ZfkXcg0is
aAomJQ5xm5nxPzpuZW9Ot/SaZB/GWtpv9EG2i79PxTw8Ud6d8EXNZnh1zGQdNx0zf66mp80piN82
Ir89wKXr5bgdgVwwylbS1Iz5KqYqvJD/NxDcKgI9H/i8ymruuMULJmNMb3wEJWwcjPhxiRRbHR7H
Qv8GvLg8aNCAzBJz3InZgKWqxpmmA8pbEOjbWUH/+froNQp4ut3SensOBqdhr+zrYYp7CEHum542
/Z0jMJYmKFVfMcTjfmzIGg6RtTqW7+97HVoCFfT4RA8pk37kcWsg2abrEPMdWe9VaIV7hqBUNJ0j
/bKTtAw6OBJRzHidBGHxV2s6k1ScSfbE3Fbl3XAJiuHyifNhM0rbquczniADugQypNs4wp3Jllx2
8zrX220cDBUfxYB/aCOYfg6d0cQHubZ0Tg9HcLr0GMX5P4KB1rPrvgxwKNBzoGjWDtULNhJGTK5Z
6aXt6Jwavdkqj8d3U75k1l76AjMnWni4SDwyHK3PAYIYWAqKKVsgWQ7MSJ78V5ZqkXupd83/VZqQ
Zdwq/B31mbHlc7R0JDswaulNXHgWYVWZwQbYTc3t00AESvkE2p6j++sfQQVvTe6SNfavBHLnIdBZ
rfA+Q7giR/NPmz+qcsqTSih0lPKd4aELOyzx7A3aaglvQ4fzwqAZxKanFGnwesVdRdAysc8lgP7v
XOKWiF28nf/jeMt2IEqcNC9SlZz4u7vlEeig7upUA072MTfdYEUGDy4338W3AreL8sFGtnRxZFzv
cMK0jSpsg67jCMU1YTQUIjygJ+qw2VsJniMy5c3ez+tlAaMuDhgtCm+VziYImmdwpMW8Fl5XNZoE
5WkV8jGqr3jFqdDNbEyDNdSdgEUffVfRxH2TLzkVTkEXzpWePhKE0vQenO6FchoB1P8Eb04eEzh5
9Ztd8dznlDhKaxyhBkmvgw/nyF+8kR3/vA4JLaZV73SgFvuQVA+ooUZj+Ck5jS15K501CqkGEvG5
RdYwX4Xsn/Q5D2GGXi65C1VIDHmu3bEiYF3WG7+SbHzrpklopVC9hreRBIk1T2HYuviOKjvh/4Pe
6HCE7N1jkRveQ4K2yJx3r6TYbjSHVjHJt+6T5uUEWdak1+Zj1k8OuVfXK/94iu+cFMurcArWaUgT
nSFGQnbpBwjzwsLrcFyb/zU8BZZEvTXIf/2NJI3eIEEMsqJeSDWniTK2yY46niTwLA3IX1C6sjYS
o++T9dCRLtZV8ZjOlPPI0RO/I/RNA/8ww19vexALkYh/NiOYZt+LbypfT7ZkrevmPLFhnbTdogyK
OvajNQPUa/6IZRA0wc7G6uqpP1d6n/SnZTLnlKZUuA+efQSpCuq4wpIHTYkZviSM7814gjGIr+Qw
QurSEfvMLQbdEarpjHZxA+Yajd3jUBuVOe27jbvgRHii2zGHZi+HkSSL78xiBXjCn7h0g3zI0DJq
mZIQWLbjVQGW5JGrLVxU3UMFzdDIXt7fNbaRlpoXrxBKAC878djUz5gDb1ICqD7XlH2uo/5SIZcA
/hpF8tadQ3LqccUXNUc1W+1Ni1Im0LUmKUZG5ve+kEtGWH2b5g20DWqBkelEiUxiALYlXvhQRxps
0j1HZN99LWK36VYMhd4ZH9e39I5XW1DboO7kC3eeWzRzASQj8HYWBhKCTR8kgGNmoZ4ambYyiFc/
6XH2XVQImfyX8gwDijTU6JUJwa3ORZ9t8hO6mJ3c7aJbnU3O2tG2IybsOcJQprJ0d3qfN73O40GC
vkxRwLfu5hlOfZpj6ikUPqqRHrxQC+uJxSCNSK63UId2kGqyJq5gthVQuz6zexg0RI02SUeE1tUZ
ZH6b0nyiiKsNl/Ly1F10kTMz/t0DdtuT4JD8Qd4oIF9XVhaZKeZzHEC2UfEW2Mr1gpNyTIQJtBjP
FM4histCEpT8vvePKFGmdkseJL7EnIihyxfLIL3uNg0qcTvxvnZtER4ZtMY7+hkMiLDLlnhM26KI
53xgeELB+fnjirGQtIlV9475AT/FTaDubR3NeR97UwWsS4wzS+MJo/ixC/5w0GDsmXKDw4/RAKov
qSbYoy0fcZEmx1fWMX2We84J0PHiuTHVufHoOBEzoUaai5HTgRqxvip8I35PZyrRi3IibFb3guOv
hXTm12PFQorSLepY7e5v4j3FZkjSaJEX0W1bUD1CBYDXtyY3im73qjFlf+tSnYkAYxRIpL0ikBqX
MEKrTweztFTqOshrhzM+ewq2u3I+8T6C46yWWSsb1auzb+xLrOcgPICVq2oBnFMc88Gy9t6uhGB6
4wRwXabaYH96fw4mraSxz/UQcCuz2v6Uk01R7v/UQCiT1IRPms7cBgzUQsWS4OEXesm0vYXMA7Gy
6qTrdWGiI/F2//1netKO5y0SHZygqGa4DQD2oDOa3RShowLOXIu1dLIKnxHOHQueftkNQqYPnapb
xzn95TqN49vJQfd79KWF3Yg+eL5CbskPNJdUpOCCgGoB3T3l/yN/edYfoAv4gWhwiVhig9LkbaHy
EKg6AsLR0n3kpvOZy2VI4Hs0DADU6X40dB+5eNVsjYiv+Z+DD70YbY9DrK8VDH67FcSeN7Hz1Le+
JH2ArL5aLo8S+oMex9cTEiLIfYlt3MIW/xVRIU9xdD3oGus0wEtbnEAtWuSrdwPcZSg/fktEcS9+
+sh6K+79WJsdCD+eqz6pcV2wXAtVT1dA1pXyOeLeQ1MS+rNzznJhvbyfe6jravkhPzjUFKtwBih5
9blQw2+Lm9R2gXtJYLtb9quyQWdgR9C7+BPt8u3OfFcpSq1zt0acFM2rFTPQF8UNV0QGr70/94t6
hSgK91GTISKxIyjU0w+phwG1DBOpivaUocnpJLmBWquAsJF+z4AFMgc5540bDf1qZCnQiKpOh5mx
EVndAfhQcHARHFbPzVG3Z2uNHpbI2R7klKY9u3snBJXi4kEyHCId/1U6+gMZTSw1MrJ47ti1QvHM
PS49/PI/yxOSfIX9Ol26XmTBHaW1u0gLLGRPwhihBXECJb8YbS9Po/qNV4rU4jfPYrjs+QQBsy37
6kMjGihJ2MhvhyxQCAQ3O06WUP79io/UbpILsLhs8MJ3O0wonExa2CDU+orOv2yHc/88foKef3hr
ufuX1SV92PfY9hWZIiyiLum4ydmYlNR707f0xPFzfSMJf1OEPLoVdIMKapPBAJef1vnNKx3GYJoS
669Xr5U3GHNyDPFCK3NuCzvVIe9u8Cjuukv7enaF4UZ9N8jOdFmQ+7mXsQyH1z3AwzXd7rirNHCv
LPjF5bx/4EWnBob3rBDvGjEci3LqNHn4kl6lfjVvrvYiJWGpihmXzVQ5IBJsOLSUfCq1UxyKIE+i
bxarvSdz3ACVecf/H0WCS42JRotXrlP9cRSKFgEIp4dNnP/RohHFxfMI5aBawBFx/4YE2uBMrx84
KZIHVsVLndMsxI4u0/fSMUZuTUpijPuxc0k41xklSkNYyqYP8ZzMhBVGQPAA6kmZ7D2O5FKGJBAt
wnaW4XGqlAFG0EPz1hgEdJEiJTOQtxFpMbBqA8WHP4kufam3s5ZsWpwdQqbasPEj6zxnKEzpKvKn
3NAniSuvhMQI6xN0FvyNxnnrv1n+JXtjDb/7uAcCbVtuZoUuetveonGpPIQHX8YG/EVn6uHPHuhn
1HnJyyqlDWiwFkoTOHhh1JJf9xNfGJoitlxltA3KUWCIBeS4muzQICgAMv6HhjfWv90GMtFTIbT+
TijD2Op6qQAvqvQW32PTbR/7unUF+D9gKDZABZqD1FfdAnp2tnee7xqh/H7MIefsZL6T2nC7quv7
aodRG5bjUF8q8s/9mABffpHAqMR0JBxAyRoEyF361NHGdACgmpK/mWnPlsMfvJs+aYqkhx8AQul8
fnspy3YOLuHRO1/fV8/5nwy1egmmTX6YVphlXLpwnFFLlq9YGba1uZl7qFbAVoQWrvLhlT1xelmD
71fpnYu+oYKMlzJ5wBp1qv20IEo2VZ4R2McIc/tQsabiek8wh76H36BZ7kZHsvsg94KcuD8EH6Tj
ZeemLqJ4JRa1opdW6fmLdEbs1BCjzvDtTU70xU2WbFePV5qY3Ulntte7TPJ897zAp/A12qs2hOPh
xmlhMW5PBGd63mJgAvgrPFZHcAo5I2X9E9r3EUME3QkINLc/TOBz35ArT0XbJTv52PF6JunmTpX2
NkV7q4Fat7e+YSTgSd7cMSPHIEKKXYxkhv9Ka/18jBtvIXpnsEXjMOfvTVGltQg89g5PbP5uBWEz
8IiF3gHlYsmXz8pAIhuZrndGjssrkobrm6/8qLcyA/Z5TcwpEGdWsOV3HwfcWBwcyF9gQWSZ6DU3
xNmyY8AIIl/ADSSZ2Jkk6GEUjx/P1/PehhG78tGXhBSrWB6WbL1M9ZDGIMAa4tewsAjNo7WwMDI+
7edCSSIOm2GosgXDeiaYX1gWx+XCXWTIyOSnwDJdLRll8FUCupiBy1rKvZq2YXpou5AXGH4UE76f
6JlBJiNeOHefBRWoSfd7uCRmpPlyaA5XGDKasnMdebfODQ2T6lDo1kTyPYpju93Jji1YPrWY7Jy/
PjFCeWTw1I5OwxNxgTIstZCBP8mf0BHb7UBUIkVdeJ+rTNqsOormVRVzh/wffnBvCNCkdawHVm2o
DUAfbirdviE8vwQUJwNJ+4rhJh5ii9iPuoWtYZ8bvAo5XS5vZ0dliYLZ1ZQP1MNiY6PHX8UtloHa
L/WcYs6+sz/WZX9jWepgVhl8bNdPGIWhB/pLVJMFYilj9hRp1IZoY/Hvy+Z5MdZejnn5xwmKMNNp
tPZnwcl5aLy1pHLotXIvtQgllJP88LbE8JAsPiwNoQcgFauu99ccHSBslFUscFwRKEiOypjBUnvV
fxxCXy2OvpGXHgBcPHg6tH3OdcKQKs0woAbcOiMLvJtpiUT7wRnTt6K9ZGuTD5PzI6jWYsXawL1t
VH8h3l20NtIVOLhygqoBZcAJA5evCsxRyQtMRmz9eShrtAo7VRvk7Z7O/VZrMP1fjcC/y+R/Jcjd
kN2CMEs589PbaXbA5fqucn06sY1VjoFUE79rilagrqXNy9kquAAgt8bD6QzadGgT9eY0DMWWOcuC
IuvDpCpjgvjn/iM2hSacokyrWyq+rP1EBSiEG9TosZIiRJm5SrHOKqMpX9Fcy72Bf8j5Jys5KWSA
mBqziK6uqi61ExnKD1k6bjt3UjHqeQTCGHdAEVvCBweRjugVcuYYJ48cl9C/x5DPcLjLCopuH4+a
5vRkN2BSyMnU08nyWONeMg+eynVkZON9uyFSBFxCWdQ8kDYwMLtkspufnUNLulaNJ0YnhjlNtGE6
TMBYyexhfrDeX1bzVwW7CRqBA/oY822ExsNGpie6hcYw6JG2tIRR80Tq47zRvnnUo+XmnZbi8sYO
dDVYORVPm/cPX0ZsygntbmPW+KY4nkoWq+4AkTYrdLFMmxcGnsoRjyKSeBvXCwx80S27YsGngiAq
4smzsVqf6DnGZ0STN7+vzo11ZvZdaP9rAbvPOFop3ZgMEe7RVMQ+sUTB8HUkGE/Llo5zAsZSzy6u
RhmELUe1vJrmSVuymRxQMLyqEnY/IHKA50gsxJb2vhWL4D84BYZMjd2+k0l+oJ5svY6qYDwHheQB
HOWGEYuTbsqHgWZuun7iYT9V656pxeAxfzOO5TfkCtFIQcETy7+HXbz3gDmTe94XyHJnT5c4WuKe
0rhjS1tSy1dTXgjbKUvDv+3s1jfKl6VY66+fphjn2PijOqGirkZepo3gg0DBKksRhl5oYR4PUPzw
ciRnLLN6Uoa7Kx5tLUSO5TXYdSJPVrrd8f++Rk+Bg2CYYCqqcPHi0eBzbOcCEjdl0hhfwA6wUA2W
NZeTOS5BthpDmaRnuekHlQDL2FHms895nphukfz2fGanww50Ua67uo/ZLt0ib5jvAigjKB58Vv4X
b/6ntk2PA9lfNASKSDXFUtZldXpIxGlSEPEweMwRAxq+DMYbSu/4bwQMHgwoBhs6toQ5su5KA40s
gRPEPOAwAXbFgRqu3K7llG4sHBu/m7kG4p4KE1S1YY97hREFWUj5gtOxTxbdQp5SPuj84CGjjKbF
daCi24N12wDyUMHDp5Yimgixk7/scwNBP/QYoYFleme7V28vMUTXa/Nb/mDTVQy0OgpEbWREK8oG
CNvjeCpUT3c0XmOzatJUdyDL3LDXJnvI8xlQhvL2R4kDEFtPBAElfp2ggDjhbslc5GnMVAVHdYpO
v+r34aWw1AU3Y0h9BZM8J0GzX/45XfTtqAEyjiuHVlTx4qYqx7jvQXhkVp4lkVbvxwPg2z1ud5Pn
yO33jVPXRwmv/ajI4b4uDOXV4U8lSMCQM0eMFSPHlerKvuMgwOFnr3F4S4Gpxo+5Oyx3lyLU8o0k
tm6TPYYxHccVq+N8rZQxDPSIatdFfXB1KIaVNMNj3wXWGiHm3uoFSYjzHRnKleVWjBn6DYKm1fON
6O0lU3AOeOrZaFqcMdccRlnaQbS/6nXu7TqV5s4tQ9QWtHxd9isyK+6hFK+YVo5KJmBfDUkIPih/
/Vc16sdEvShCN1y68p7bws34QRAaLEEj13lvVntylyWCrZBgRKo5wRVt2asMRoaAd4JFNH1ESDnd
lPspIcng0VjsaKvjfxwr49bVBENBhsOAJmh5UvqNgF3yJkhuGw8CEE3UPB1+qWUWmghQQrQyqZke
hVIRu7Sk636GoNoTayTZt5DXpgrYeZhIZY85oLc6wUG9v7ifn/YwHi5EedHlq8KWbvNp7QskZ5ZP
05dA4BMppX3c3CEmiOysx3G/YxPjlQBRXBBTKbvPSQGEJpVrPUjYN54HoNn4Wf4B4uFZiA+LXZUC
CtUN+zFKk98AQTmAY+0N2rXA4pwAvw+yTvFi8wgDBaid2R8UqQDKD1OjaZgPOe3B45e8GvRz2MAO
rr5S3S9KTG/7+Qkg1sIDLzJ7O2n8LN4dKimxi2TOdLHZGoWbjeRUoYUwIGPGrYziQMsRgM2Ppaxk
Z44P0WQAvHL180QLcB0SSk6rSWM9eXDEO89VweCJsHX1SmyS3cF89EbzIF+Dgi7p3n7IyMPuMm2n
FJ1+PJ7ExjJXZCCo4/A/+5HXMyKaIu+xVzR+Slre+EI++NcuWlw4yYIfyL4fvoU4tU6dLDg2PHQL
v1F8vc0CAc/dYBVLO3BX8MLj5TTphFrmYXLcY9TK6RSVcbrOye4xiKCOpqrzqGyAxPI73MIvY1Yj
nMogQzMjHLNWXRVmQhlBL9P6ZQDcNLzpMmU2ceIgejHsGY7weNDX7/bcpGUgfyzjzjGKEu/zjYbn
iMUZDnUkm304koEXcnW1PyKAoKSwB/wykba+7EQDVYbbFQ1pbJ+arjdWlYOuvsPS+P/NdTsUjgXx
BIDqciMXnLjvbKvgoFTohI1DHfW3P32ejeAQedRb9lKUDOZsTAiVId3dRkqdbJTxt/9b/QA1Ympv
B/Tahjdar+/oetk3PA9J47ylZUZF4ir3TrFsxCtyIrjnHHZ12ZZN1yBvnLY22PHkhufU5LVGuaPz
BLUjxUgEusBFTJF7y8m8SvPQUZVstMT96j00ilJGHIDJOWCVZsoFHJhYXR/x/LVMWOPyvn3JpMKp
A8ITqmXpPtCi9Yte1zhRSYGVUcns1uA3O/Mf7InBJ6hYqz1YAq6eNLAlbiIidSzsRfBdN4cPMprz
0qxyP+Px+yjOohOtbaj0Kri4qt21ckd5R24fY49yuD/OQPjcc5DyhS0LCUOBWUy8wvkf31pXMm+M
0DGzR5y8lxdGC/N4dj/tXUfgxz5L6Fqu5jZyoDmH+BoC0hn9796NR17oTTlf4OhWSU71wF82RztA
eUGC5wVBjsLfvYSQ67uAJ7GI/AEjWTIApTnjEFWvER2VK0dmcreGkJHGswUoLiMObvActM7Seji3
ESOLExvVp0kBCSR+zny53ZdMHxkwdVTmYx7M4hfUnykTw7HjmjuVhSBqdDShzGp+UPe/CdvIPyrV
bQnITe5I0JrzbWIrf0PJRY+oel6ifVN8doF+szAeUw2HBPoxcNJhgbIAeL9+tgyxMZ3knzD4gba4
pXjSWpD7u3NMA06LXiWTQoAFVjWqPuDzHxkXRqOsD4pjCEUO0B1BRasbPTK/0NXfGskQEahSLtde
mfJXOlkIkEb2RxcCWLHOXf9IlMEy+yN5syjmspsA+ffYdksyXBOCck7w0q4yYONAzets40J6jNMa
b1YWx/XPFDLse/IfN9XZssfhech6X8ZVRJoIuW0aa3qfx6UKVhjBOqsyd15fplKeJigO1tgs1jaQ
EgvBpa39/3skcXFBn58/adzpeiuyaPgq6dJBkeJ5vOYdM3RSfKw7MyGF/zC7aPPXJN9/s4rDLbQS
KEoCB7pAzFLb608TBjtMUOw8/lKl1g5QCixxddTFcxDLzzNsXQzEPD6w5oVyHMsBU+Pq/bHqjuzG
2nL3J0T2vWAztGYWg8gcr+EraUk53hkHNjw9oqjyx76HYxiwBaZEJWvOSlXovW5+xZZeh1HHnAjy
1ucxUxLPfDmw4n0A3NntOJUcPv6IkkUkD5n4++llW3G0uUDDvowuVHJeJ1mEVjuwwnch80SOwr5r
h5mTDtqrPfOwjw2W5YPyufufOq7UzQHsaDL1uBIThpMcZxBtL/vroifM2rYMhDnM4IetqF0mJ0fL
uQNvZYnybQ610L2V3Y1uzIjF63ZrVP3sQldmHbbzMjsNm29HLFif1apQn/in1hkDwXdVyS7R6/OA
0k28LHxHvOFYqFmkr29GE2keXwQDhSOChtUP0If/97XOvvdFgarLgSDWWPgS2A7dqT8V8aHu1HG8
B76epcrTxp87b64KFuxakYKuh9+HNjb8kp0u7Y7Og4PgSiOSumuKuaygTKZ1OdKkdh0pzani7e0F
kw+StF6R5DlzrwjtTQY8VjU5XJ9wd34mp1N93ppey0SWt7tQfWBm7Hs5srKxn9c+fcHR9qGPsts4
0w+H68ezg0YOG9um3CypxvPF2LBwNWH2xk8mf+xE750OQcQjpMf1lYm2H3CWF/Q8shM1kmZ2Exca
3GgiIWVGs44JDBTOioW8ySt6mV8GTSW/EDevnroSndEpzL82wBJPSx42dlOH6xc/F+8EXcJDktuK
DtRLZKwBT1vGTzS7agqjETXZ8oYo/2n6qCEUOz6WWDudxp7BVcwoPDkdgtZfd8VD8OBgUXqDQNkp
L9gJpC8dgT8h1UpyDYcOgZZJSZAWFtY3y8nzZ+z0GV7kqtamm+A4s0cEKHMBf0VsTwk/NmpN27AV
teDGjKuojt2b4A6fkDJLOww+Wluz40YvPvP7gXIRz9Fmu+3/9FhAtUxkTsJZiYQcyYuG9UYUvt4u
AZxJsZqb4srE8eMo+YKht4yE6dR9hvx9/9DvBt+oCilW4De1v/EdVil4PmazWz9aCLyOpG/ec/zk
WG5016FiLbR1ksHEjEReBjNPx/tChFBZmdZ54dGXrMumsG1iz51L6GhQmfnttK6dRLAHC4WOx0XZ
hUSEQjS9qOKsfuUQB62ZgCXIwpOyCiMBy/AfsNUI4xd7xmg/s3aSgYgeRbl8QDFug417OPLc5lCC
47GbVXvJSMxaRWcwNdNmn4Y7QjN+YtarUPZjlc6f9Wu5+A1GAoFuntxM5y3RWGh3r0TaApHuFqoN
14L3fQL7BlHX6SVSV9mlmi3Bh9YYBQoMT8n8q9dkcJlGvWB/uRcmTYs6Eh06hPyaBF/se9gs3qAu
7BOKeky182+6FxMlKvSvKSf1U5/OcOqcgJY2lxNNV9Tv1dMAli7nuw8egbPECjVn2BjbaumMPLoe
Y8hDr5EutSbgqui7ZwI9/TuhUihNkoabdoX8rT8JMSl96g2oolZ5mwYdKb3cTkYvkDalnGbft/5M
XFH58xMOra08tGIgh2tU0jmS4crq68q+vL3AQ7hyrKwJmKl+xl+K7fd8Lge1uhqoUP/ighE824xX
Nv6GSyCCF/I7olxqwcz1Cje/ODeQGsxlrS7i50IGdFnjtFDnOkrmMiOm4TDmmRH6+J0bv5ETUUGm
zUgWd8Y5YuOsKA1RVxIVFbh7N5pjrpbnDz8PNVdRkTn1jGew+JiLqVvTarsWGgkRWC3iKxg5r/a9
tXZauzmhifWToWVH1v/c1Szfgtdy5gwdD6z+zWcJ/AihRM8usrgtmJ2smE3ndCPXNNUUyP5K7I5N
DvWzcotAjUVU5vN9LPJ2wdPYPrndLx8sWWDqUWLHAfn/YHY5q90qng/o/7M6wQNKQz8Dj7Gu5s2x
Ki0QhuJwk+cnX9g3yEJAdE6J5Q8VGaTDuYXrIxEgUhIPDK1a0uuPVIrAVirUsrFo7um4lMnLzMvk
SylSejdR9mD3RLtqtnYhfNDeUXsW1FhlO3hWbU37ihCClma8pABPBbRGFr1OwI8PiPxn4ZRUhUea
OBE6Ma/MRpLhoK0PSQWrLkBgjWd84+6ywK0+0VIsXmEAXmDStmXr9f+wbPhRXL+/0PCz0kphhSGT
ku/pnNKBUMlefHbzOtJoGWbrAaCU8nuZFLsdam0RowVg3Gm7yw07KHDwDBGA1L8l4StmeDIjs/SJ
1t5kbD6K07BrF1Gg++RHP+TacpXRn1MeQKA+UwT8i8MkUQwUl8AUEXcS8exvwxExJLs9sHAh6TaG
l3DR6O4bgEkyJ8Qae0FD+jwjHH86RoktM6k5nlS3stT3yzLUnapnXhikUK+NxLLH1mXeE+NuSG75
ENnrKeud/yD1G/a9UH6/uvoaA3C7nU6cUPFA1QPEMl4uTGse8LxViMaDhcQfdkvd70cQnkk5aLjg
VbuEsw8eEhBzfGZpKPRK1QUHx2FxMmW7RPStsmK3U7FSE2unAykAxI2KgdfO2oxEF5Qrkx+Fkiqb
zaIYUQoVC2weRaCyG4ylxV/7eMzzmrqzDy4OPw98L7de8NWfj8uhvAN5DY1LxX0hiIbnDMUTb3x2
dHACp1/9y5W3WlbQJdtq0TktPnozrowrGH/39cVfE7Ofni+1vOj2UYs8qKBXjeCY8SNWfAg8fCJ+
e0TdY3JO2ZRYT3o6nt3yz4RBMEKgs2Ead4BIIxRxHbSauPJZ6C2COxDXi9HpebzFo5dta3F7TJ6z
UQObOM+su0Ob7ThS+8ztD7OkOwxtbsbswL+2SD9ZkTyncVUq/i3/BFsJtzM52x5GI3zz6WXR7iY7
NX1BF6xmmuyhET07aXChGaWT8olPrLoZx0CNqZsC29DpPx/fmS/+OmZOxJZynCK515J+dfMULCcR
NN/8oeWLX/hSVHAPyN0faH1oua1S4uuLUKitDklIgnHoFVu0Ju3a8Chikxz0ht/NXYYA9BhLIWGA
RlZZLilyno88oHQAER+rzKkjc/IaS52qfSM0kvheP10CZe0Bbipe3Z3RNdMJ1GP7MbtEC6Nvos/J
Uqsd0fAAnMtQ/UsJWWG0KdKzQQu27JSHgNVVGLHjwMYNT7ZORSj0Md5ixp2BHuhQLhpDiaVpHgM1
AhOEECxUaLB/iit8MID18bZnkDkekumQ+acgV+i728xOaNfnIUq0tdWOHGM3IXSb6tINX5A8WnaW
7yGmKtapCQwvOCHzroZx9t09yhW6p+bx7a0T9+85i+1vBEfdEIZdoql2OzLJmpL3JWcGFWRquc3W
tYysok5kbG2FV/Q3Z1JKkrVPSbCAiYw/A+7GDu5gUOhfnl7aNzumZBjFQ75krv18pZoz1tAJYqQO
Zbom7qdWQB2NaIG9vW9DCHIWmC10A9QQuL+vkprA7QSVZroWgmLnArlZ1pXeG21viNLizTK5Zvxa
0Sce32eAKe7gUO/wp9B9SJMNYb98DuTREs1BY1m5yIoimRQfcaEwlUNSVWVOfXZAVD5oo5KsNQTD
pIKqEBdhAcEWM9HfoH1gYK/C5yV4mMymWH3XCP29Tonn5fWly5pAC4hDJaadnqmHcn9+U6CvM6lZ
cBWmtn3u4D0AcQ/nk+4SM4i/+bU4fA9j8V0Pxn7CVb3uyorxEgyvwj18C26uqyxtTYvneIRgwjqJ
rHQ7fMDOEXtvxkNwyUC5WIBvnM6C0inLgOLAKSU6PNIUf/tGtWt3/GoCj0+T869/lpKdbz0PEYgM
Ybsd9HGI7HbwCjpZQAxWupr2ubBjU8TuOAC4BWS6ZB0DAiOgYFgbdUHvv9vq8ketajC5hkaicgxP
/eH4GY5BhpcCYcNhfsGuWmrQ0HD/UUzVmmsjU8BxJljLuwx5KPyP1LshWw55SJNd1oPHUHkXOjij
wq2rOuolXDUVMn8QnBZ6Q2cxVdPVrJZWz9y7wagaKjBJO4ilma/Cee1U5lw9FhG57rSJ79ll1FWl
7rnoUtngxS4d5VGKAQEWtwacGfs2j1myOGuBbsMEuTv17S6ViRl1Pz7Y0WywqkT/4FECWkx00wGc
5x/LN3SpQX4IaWdZkONmBLT4OPNF5QeMhroB/II8yq73QOBSZr/yCH0pBbGIv1ZG0v+lgRdI+YGu
L4+4SsftStP47sbewIF0srttnMevhLa7FcvU6mdnP+ynzuYH8ERp0vpBWXMS4KQYE3wXarAvn83H
cCd/gYHCLDGPE+Uh7U1x1A8GCJVjlvirbBy0FHrGFEAhYiOVDqIN9nMp9NRknLX2z79zkBPZLJLR
mserrr3YveGKVyf+5rTAsYFMVfei374tqv5orGR8GPpjhF4gb6wTwoQKZA9vChZWzMNtk3MSMmeo
upupN7XOKW53MKOmAaJsYnh6Bkvllkvv+WsXei0A2ibPu1oEmjzs9fvTP6a0pVnmg9MsxHATfysy
l/aEXkf4fmStWaeH87zPXDEVXlG36lcbRESV3PZrC+YJ9u699JoWdgQsaeWoPiHBei/RTgQ8FJCk
W1LsGdlffe6HjZ3DFiee8NJpPJ/zGUniiUA4Zix6wkvb5ZkgEsaJLm5P14ou0vZ4Ek/hGNCcq/XJ
y3bIW/zVBQ/aTYDePj85kNnxdyt6E68UiVPJd/k9JjS6FRRdXRxf2IiEJ+uLAG902CIhBRy2qCc6
iMxxuuqXlBvijO2HbSxAqiPbb/HaWiXXopWdZX6phzzj599WHTYOQMteogxjeRHxbWLMgvmqzf8H
NbzF63vfFmUBSTj7UaXi0V3Q8I6T7DlBnG8bs8RUhRsEvRKVTxs1ueq981x5UjMBfyvImASAAy0w
4/t9yFzduqeoODVuTHlR7g9zkvYwtZwxVSdPbzHM7k/YNdIPp2ZvcNT+7F8gUxXjc/i8jRoOCdmM
1+lrVMERhS9zyribJN6MqEjoo4+7pRNk+iY/5F0KbaQx2je28Jj2PxIcwaTs/xISnpyzbDmyN6LM
DFRYPYI5R9UkJLYjmMWpJEYXthCG19qT/lDS2eH1+XM6YgrklvcgMS+3qknT77ckTilrWz8MDl0p
vhip0q3DyYs5J0K9BtqZvMNmgKBZwOo6byyACwSiavtsx0Tlj2xTmvq62TbNm7XH9oaKDuN3gnJn
JC7V7n4xVC+iFzsRA0kVSclYDtGOjrnUn7CBUAkMtrUjjtgJdeVolUImvBJlSgoBbHr3zX3i30Yx
8oGrzcf6yRiuH7icKzEMmGZ2YyTvcPPzQpEtSyqraqsZMa2lZchA4cTN6Fmw2knUVaoyTndef8AD
QkLD/SbAucxQbt+2YyJMDKhMH4NCiPxJGjaNgph8/JomK0cUIv96imDD8HVwehH5BFrOjwt2PKFg
CP3tdsM47mNAztEbBLId5TqwCbCBzmZuAetI0V6kD2XJEUK4blfTszdYbZpr1dgw02BHFzNuUccO
iK3nrQYsMmWAmTmg8vmOINpT0ql7H4TS4lFAIpNwby2ruW1khc5bAYNaUiIpv9mbnJDgT+LL3OvU
LVDu+q2GGunbo2yRWQIm6lz+tSffHmTw8iZz/eGq4j9MTG62kxiiAux/N9vPzoInvOMLYfYjk/4B
BBCbNdZz3jdtYlKyEUqLM1TySR+o03LIy8ZUemO2QynC6dUCr19ykXQcMHWXM9f1mtptOElPGAPX
3gFyaZQThVM8aEhBYvb8HYOOs7cHxqLnS/1lSCAW8rvacrkTFVBISMPQiX7w5Qfrr4mn8OBjUKvL
8C0HqSeQYCyyRwuzoHjCjuiFD/uHXSS2rliuEF0jbjQbCx6SgGmsFf09hKaqNBGMkGpNfbjYUP9J
8zz6PdUNagBeheK5oLArunOx9/+RwM5p91xS6sAbXmNCrrClaw21HRvzSaqMdZMNydGSKymYdXAj
LcgMHhrYT4/iRZVsaWFfsV8lkBF3pwHs/lXC8ibomGM2S3WEPnHi9h3Yps0SkWRNDzIYub5xgXUD
vHoCo1XcNiI6betLiZvvgMqKLfkklsgq/CcE9pcyC/m964NrbusSqSheoBrWbbbZvIORPOvok8+b
gk+K3dyvlNBCT7Z/bg+xzMGOZa1egm0/ds7WZ6so9xtIXajMmKgpNcVWE04KEZ0hmopQ/Od6lhgZ
DFoU+D72bj3GHDcAKHKG14f0FyPc2NT7mDUATmEcf9hD1zjVotH+SNyGuC+EzVv1L6WQszv6WG2w
MrzFIirmMldsHl2NNJ7p8Nna3rYyGuo2KNyyTCwIgnmlT21AEb1tRSEdvXY8CeteopH1DAPuAgmA
iGKLx94+sAumXtZbzYdJcx4fz0KqHR530GjeNN1XRKmkM8RWEa3hX3VlgkBiHEZPJNrsg31WGra3
z0j1Nf4jeXcDk0+fhzr0SRbwNhyL1KrJfLs3z1igEJSqgJGyk8ISNDQhSXi0X/RbjNQk7PHAWu1y
pNEGR3+2xzFoW51PE2j0K1Q1qYOTVrDn2URHlNb8r//cbJuFX3iOP+zA2cd0H3h7m6JXCIqG2PsJ
/q0lt1Y3X37E2cEKFMhcGuHhRKApREjQikwutGM3cbsib3MV1dfr7Nhno1ofFdrkSZIuQIjzHgdZ
wnOOR2h52H8M4BVNkUu+kiMjbQWozfGOEkBQxt0azlj//myfngus6vKwg9a9oBgPDzcFhwgP81T4
xNbk6uTgT7qNj7SrGkwnjro0ZDhdl44iAnTNJz7UMQBqN4NCtuXaf2uhsi9RNULQa0qF4I4ghrba
ofLNG75BUm63j4qMwdr4qSDSVb3LBrs7d7nSK6XkbKikSE9rV0iWoD0/8W005TkHy3KLtCedmsqE
Foc/gJSrkloV8DNEbgogx+gcJ0Ind4MSpV+dSIeAxiwM2XTRx8gQq+Bb18uBEylU5DyJq7c7qy0G
cRf+tNh4MgwBWdFftNdmAVkrrRvN0xw9mob74zoXOdgRt469L0D1nsuA8EkL1l1nzpqpXCi5pzkj
HZjIsEx3yoAdgShbnhVGI/0ssa8teqZBUJQH/kLoGFcg3sumkGcOJ3OM6rkc1ZfU6B8USdRjWpWL
XwWoaKnw/yIS5J48jdYtYAMWydwlvz7Lx9zcBzPPjhV7bxZ0SoybYnjXh8sIIRu9zgybYEkZMTRV
H3kmGR7OivKzAecArL+p1sisye01Fxt7nppybIYsioue0JO99PQZB7v2JIIgqjzMHb9pdzG0u5G7
kmx3DmVS6X3xqbB/aAUU4kNMBnXG13a+uklx1pj3Rnzj5YMsjjxh4JMz/sEKgXFCSvRtiFx+WzVN
31M/HP+OYnBBAFes+Im1OVcDV3wXFuHTG1HkhwbXW1K/Tcq0j4W7ixIvXMTfKPKN4EcwiBmh9Cal
dF9FnbZO1Acz+DB61jyax7siwJpRRFhTH4B4RWdnmoZmgRXinVcN5zo6jUwz6xuIIAsSjwEsYtE9
l2GG940mZ+GnIR1gNknWwgRh2llixXcs6IQG61WwDLiTvoDhRinoPHcedt7Rno+xhtsCk/HdQ4s1
Rj8TWt+OPaPfCN+sjfk4VLnn5jpykvIFdQht3pN7vOJfZ2uwJ15xTLVIM8RioNY/ogrlch+IS/8S
+hu2d+cn9Lcs93xU+IuHVgXio5yC2b7AOi6F5uwa2ap+BXDBMKHl8I6imtVTgtaxMUh27TlmEBiq
ukuQD2ewZQInv/L7vmGSE7vh//AWtJOlVpY99OZOiNwrpAYSx9ENXcaGw0TcmPHtM64fn+kBXBep
+60xq3Oe6hyrN41xfEtbp/aRtp1Y5TByhEq/vO0a7jYvwTiMwIYbq+vsgEe36KQxrQhFbI7ZhZUz
V6Ne8sTnPKMMmWSPXsI9jpHz0cZbK/IcDMMH0puZvlfH6TGk0Ia3OWIfP/A+1IYWxrIcZY02R5Dp
5y2m5evnszpkg6aRSga1H3BgQahCOUlkm8vle6UdbuYc9G0UoyEpbGsOoJ65EKCEenTuwmv8R2ks
pFeuDKdbWuub4LK00MSx8zBjDxgrP0c3B1dxaY3JcJ/qRe7Q4hiy45+7JisOk1uKCS2hJNPH4O/H
5r75U75TgIsNC91OLlx7zBUB/MVoqphDmvvKZCfObvt1SdhCuTiaUlN6YzuLw5V9tDC2SSZuOHrp
VFdWKEi5eexEHuZ8DFU8JaL999XNwzmrBCykBBNsj79/eM9jwTIRltPIdHvgYJjG/TDSqu6w4Gko
WNqlzl+jy2O2YYnbSgB0k90VRZQC3B0r/fEBxaYLjSnUMVw29h1MMWx6BvoF9OwkmFEMm9/2Vy57
5ySftCkj2XG343/4qf4dd1Kc12NkDbxfPdgUrgWDoDtvEqMD6XF+jYTPg1c0B6mN7xzlvv+F5a7M
cQLfLKOdAOEshIaK1wV/4YpoL+Np6+1tTExgbBjoV/18d0HNo6L6u3LpVx8sNwGNENhwPX5d8t6f
GqntpX2RTRyjMFr0B1tKsJ6zHK5tRMsBR10e6PDJWrlH1US+pJdIC1gveVLNvo+Hch59alC9kfrg
tiTfQ/gjDz+m+krI25JtFPBqwRll9ZHNwqDHVtIm2ld2BQC1ZYEo09Y7Wy0cnN1RqVYlZA8iP3Fe
fGDWamYwsoy6G9UCgQ+F+ZQOcKtNlGiMsXzE1V82aYNiXtgAeqzvOYuwipdh4/ogu1qZvhXSCgkX
xzjG0g3VnHFQTWTLPb9vn9eO9Rv3E4KPMwF1cDGgBQ0QLvgxEiDbXo/pM/+2Prg48Sju6GwbYCNI
vqFPHsyqdypZyO2yaC6yGAndRb50SrsqltMqBt5eudc5HHv8R4nmVigQDMsI5kTOD6vTwTSll6rI
gdiRohbIyGZRDnkbJ7sJv04lY+1QO9fbl6si2ToFjnfaJaYG8azlOh6xo1DvY2RNr218QY/BmzBr
fKoEbAQSBHGdGuqB4vDxqOBwqOIM8pNW2q0z2srw2oA3Jb7SKkWwD5A3C2fVWBrz9nXj505csojK
pHBP89HhAZMtsadRrNfZK7UFExWJBaXDOoY0qDAHK+Ugp53Fko58B9Xpn6j2Py+a3Qmv+hxz5rdI
6Pr/RBlLGD452SxygCZP5SpzDaXkj9H4EVJ4Et316ZnJ/Kt7729jq2BeBY83u2AeCFbjlLvCIcFv
uKnTyMwkQZXs+BVMuaiIKNBZDK55frIbJgiaNYDBf+fa1NktImlxfFih4I2NECVh+c++AzU/5VVb
yvq6x6AksfldeS9jlm2dZaplQ8s7QmxY8l9B2GN9LAc3jSe8wgyD8fFn+K2qUD4KPprIU7jgzM8I
xpj3hOVPSfvVDUnZ1x7M7O46/nqS3iGQB/JLzZL5NkJO4g7wdv7UPsZXfppr79l09zqW/VfqL1a5
U2v+ouncAffZIBOI2PRMjUmgshluZBhmRFbm1n2bbxXgJlgGxLP1ectRz03ZmUsIgfdkcWTisrLX
1WqELkZyePDw0g7arIYTRaQ4v2ZJzYAHEC4HztXprR+foA6UqD0MRfF5gu17iAaY1uB31REhZeti
R1V/8a10QAxmfs92S9D0kBVcoOqJSQVBZjR8YXdufc87vlVtkwXNqGW7MC252VqlHxxpO6s2VRy1
DkV2sFu0hVsBeugs+Y5UsIv73MpVveh0LW0yYFFvuN5moFJNM1IZ/dodP/BofjtI2pth+tRGbkd7
GgLgzCvQyZkAcbY/25SlQiKJrWfXRtU0HeV3gi/wZzRy9bzPxH92R1LTHB3oeunM6TavVg2UO8Zv
sGQuP1SReYkh2HF3fkf4cUaYXMfEP3UyUBkT1JcMF9qdu1hk4l6TuKiF6Gz4l7KqRpS662va3Osf
3dyjQOOc3cu9kGvzszQktsiB2xpELyDIKonE21fruNobE9uYxZyaWTR7lOcJfPqWt7k+7X8+/Pr9
9JUUipwITWvMUuAEI9oLhjWB75AJSMf2mKLaHJsYUffm2oOauMXvuvKp4baYc5GQXHs6wVSHfx1v
tzni2kITv0nHl+0uXbHQj2M8kEzwu+MwOFV1Xg1Hiu8+mOmRIqEOmJ13hvV8+ewJiMvD5xZwCC8M
nwjbbT9tyJSRpOfCxEpAUq8jzTmA9jGtB/iTLdKIXLzUOcx2eDlmd1qngdmZYMOlz07AgNNGnwX1
fEkbRV+Lc3JZuuLEdR0fU2+V3SmrEzV+yzyaN0lpUAe7M53rT6I3wbsCdm3zLE12cDBpgjkOXy32
rzHIsNZfFb5Ic4+s7dJ7qozlcTaJgjtJf0qOdo6EEm1cRcG26wNc3MSkwiHIZs6teBV185DmEdXj
b8hURbKXxaaog2jcUFQ4oZnJF448dm56oRbYBEQwRngx18yXucFp9EE8fnAfepHGZyLBdHYSuoIW
/zaI1I12JVRQOzVzgRRMJYnScvoerf2EF+dkzo0br/wkbW0fKiXtGk1td5nOtSjcxXxrjKJhAR6T
A4F8NCQNvLdvzrA/EQLmlZTj6EJfKikjcWT6sLWz5P3RT+owydI+vge8R/cP/u2K0zGU616nQmIp
SrdaewkqbLSbzTYM3kIAAPXG3i43aBfhKQNMnwR1xbOTTDuzXwtdv965DjWdux7f7oGZ+3tkfCBu
X5BTlutXkB2M0w8tfYx52IyeE9S+uwCIe9eIRzO/spN0o2S7cBfZIJs9pvjEJz2VR+PpYvUMuOhn
h27Mz2qAaJYvfR1XtHKbgKh65FUdjwXWv6/y0ZEtW6N1umaAqAdOX+D1rFH5RfzT2LT337hBJl+Q
fCX760X7gUjdeiRkg0Y3OogETnZ3RTd3gzqog8veGYdiaIL3M0FCbvRszakMwKKjNSGm8PoH+zu7
wxATgo/8bOt3U0T38venvIXtVuYxQ5xAzZxDVuSIbrRriAJkmP2zK8TJ52ay93OhjEU4FZZItRAB
WDYNPbyPsWKgbWey+ZlFySq2o6rp5dsqlRfKrh8YTer3vpgM/zlhmnSKGODzNNigwOpUl8L/XQIU
VODBWMLc8RmuMSzuOE+oajfuJc5aKNrK9HpzK4Qajh0+J3pKL2C7JjU0Iy/HR1/Q8A1aABNQE8Bm
V142uajDGnAUiXalpihcbXdCoo3GI/4Bl/az5FSIJsV1pceoaPiChw4eKBPcygaMRXHFKrnK/9Ad
eGjSm+keUc+6Q+j+HZo00ZhRwoS44FIBV0kMddRCJrby/k4xD2MeHrmi7phcIIBd5IY8VGRMeAvh
qrTJKBrrJUhs93iOyivI+15jbM3TvLT0VcP2P7lhvTKwf2bJ/MafiEt14CbinmbWvaSQEDXQRDl8
qn1P7aOzAIVdsWZezVrryKRQoGZ3EwCF2waqR3tofn8GgPnFpxYjSC5eVlo55hvFLqRhtdp4HQBY
i28ndpXJ8PA/VknQXbefyj9rh2hBvLd3rA3XTLRf4aYYhNxISk5236jjBQfGLQubV8E0A54f4WDT
qGx/+g9zR7zCCxJCEEKgrCVuIjEci4W2+JiP84DV5hVQ9GUFph7HTLt+Ut6smTvOZaYFolSLHmqn
4IW2FGf5UmUcobwoztw+oAGLQeLkKJScfP4xTdpbJ3R3Kpxn1KGAuueEQMLpakhQiGwZQzsW+cRa
lluP4UBANPQD94kBEXHlwat99OeIMFuaRXn86yT1vF1+6fycFqe+G5DHgMiBMOc4HukcUwIwS9j0
WZ+y3y5592Pk6htVCc7eVcNU+McE12y4hlZSMDdk3H4vJ96c7OC7cvsXbq6dSRFM4ySLhju/hPCV
XGADFC9GDb3mMZqnijPHmonNMgBro6UrAgTSuvoXP+ALk+eq4XGK24xTLUBebuKAi6ZdDUxGvHTd
xasryvcVi+1TrN8z79tvEtZMLtAECM/ohcGsA156didKD4hutIde4ENsV0+XCzUC6cq9Tg+rA4ti
Tg+8HBhfUFG5uCC1NL2FfLAylm8Z4KFg9BnX1Ng4U5oFz/J96pK764QV+by4QF+uO3AuJfvkW67F
mo1c+mJ8WfyF6e4coDzOxrCHFC3CATDgfum6FLB2uCN+V+KXcJiiD/brteSk6geIkkmJiJNTyhhy
dAevBpjYlDslT6LNG1eqCVEt8byZGrDCt9aPJGCxGT3DcZzQMfqAcRpFzpWptfSaEJVI/tLqWmEq
hkD1xbaJva8r4jmr/gKtWBqeZgySnkkFOkm1JkjvEp5zsIlFvf7f/k7Vpp1y74LMU1MXBqtOpp5Q
s0DHiAZL76OcKD57xtzySqoeeTuHsogfNCh4Vieu1nZgYV0MBUq1amTx6ffymqPNoQFsQfGVykdH
48lmEXH/jiJV6a2enLdrtwTHd+E6rCjTM2CIWIQlHOCaGhEkTw920PppZ//F2oAi4VxKOELJKwPO
ibz6Tp7DUkleRN5+duozPwETUwTIar9aFpnUS3EGW0Qr0VpaMdVc/xyA6zMu2obf6NP4ym9k/oh4
FaUv3qKTy4eZaY4uflpEL+zakteLIq7Sivof2nlfqfh3G6vmvS5WcYdxCg17XXfokuCB5ZNGGIEp
3qwzSKBfAxCWON55eeKeh6NpWZnYp3L1G9AcJ5YHaVovWcqXo5KTKNnAH5XoJnNdkzsd/xIdmjg5
bzs9A4IkWn4iGv1yQcaggZ+GG8G8yXDafacSU25h+JSlUT+poK8ajlkfoGETazAr0qn5hENYeX36
QqaKnbScjOdIdCnmRmrL4IKxGqBeBDAtb0ETvyWiiX973ymffn02erwUPqbPBLLHmpuo++Vo4wxc
G24uiDVEOQGji44TAWmaXArWeHrRb/6+zh+kMRAQzNWDJI5tKehF9y33kQBowynPT9FAZ9TV5wYH
fmQphPydy+5virCCTGjdtQiRLadcmUDGb/Fwr1RgpWjN72+E1nJxvAFazbYD69fBk/FNTzp6XwbH
7TY1B7u/yKiXOY8VzGU10zybacd7FCBiqeR3SeR4wzwHeE3e8yEyIpPJCuMH4QDo+qo1bPj5AchJ
4T6ONMHjKJzX4yLzOA+kgxM4cbek9p1DviN7Jiu+SY6nW6fPggJ9iNNAGWN09X0ifX7xS06Cp5st
wt2FUaUtFCiReastcLSq1Ha2xNO+oUyTUK0emhhwGaTqLQMMM8MebDE4Xc95z5moe270RiUjR7ig
QWe9JimURl75VjewTIMOOTcDD3RbFe+J3rW+BB8YNF/5zz+IIEOoV6AYVfvoTkhaTzK9u4egA8CL
0fiktNhjJDo7DwdpO/o95zIFpkz5H4NrT5rocedVyCXb95XbH6ZzTbk3Gxmj4w252Dv+8kSk/AwM
1X3F5oysfY2s4sCmzgs9oHcNX8taFszdNX80gyVRX6rRUJJSNhlwdKm+cwXtElHVf+aV0yY+nZvG
77ZX27MMmh5fVSysgx4nj/kOO9IWNFc0dl8L+gDR0JiXSGVpMWI1KCv5D8rFmv+rjmqXuCWjfDXR
BbuEHk6A14RAx3Gb9jZ8HhXp6SZ6+pp78ftY/y92+xAOy+rBgW4RgJqUto2yztmX9A8qU3pR/RCJ
hXR6i8lkLKyRaWlHDoV4IxxG87mdGkrYJqEIrvPCVk80/Y51w09ANkYIoZ/3dzRXz7I/e0EVcvdA
It/uS1UCgWGc9syDjDYTYCC17HIxUx/EpSyWgFV9qjfpFRvgyof70id/+SAOodnP2slUqOcjZsGG
gF0p5eKGHdpM09ErA9I/cqhapHYxm4oZa4XbcNgVYt+4CF1bBvaYKwh0sN4KfmJwjsX/rqwUChtz
kYdazCLG40D0L+Y8FhE5RMr0suuAa9WDWY8jpf1uKGSBEtB5g4OKGKVXyjrWo4DV7wQr9nP2m5aC
+Qfr0nqq5wltzeFEWrL/o4igPdqoiqkB99Uy1q/x3Sw5ziP36GfjMlJDp2DrWC2c1KoYKYiElsbK
edO1xxT8lUBsXo0RH/YtyAT+uXuwhBFqu+J5Wtb9pVlTFtdnspKVD0oCcgCktisO1BNFqdd1TQ6C
Q69d3xopYl7ulQaJzmEd9GglaIvgSKk8lIAJvW8uS806xapjhcIkTBH7Z44iL9fF6+lof8BGykIv
YI0mqFrDeHs8pk6Cmu+JmaTXtJPDo5qVpid+c/azntWfXVNtf6r143L0+bgB8YTYv8iw3Wp2xltt
bF5RCJBX/uHTGzCPN0VMRI50oks8QjUgGAICdAv+dlVYiIc11ngt/Ogil8cO0lAxNhkimeafOhMZ
/SyOSkJk4Lz5sZi8C7xKT7sIAJiNWkFmNMho9bdsrtux+3f310Ipunu31cAzFSFuFkMZxXosWLX5
HE/Tj/5LuW8AlemUGetaPK32ACKD5wmpQlmKLkNDlNwlXPm7L8yyoSjmynncXFp1YtsvU72jIOy9
IZ3bY0DZ2g8tXD7ZD3kWaem55454OeNAoo71RaN7Ncsb+XUMqAC0oERWnKZxId6aklMJaUP4UCO6
FsMSXYpqnGf3t8r5QPbw7UPWXoM354a2F479+BNbgr0tuD2h2uggok5F5to3eT5cD2QE0X7yiuA1
R5cLIjcjOBw4yM/tLXSbyHL0Ind8BMr+Ktixn00OSDHvOQhIt3fTHuUUsbmU0i2SRRy/pbja1wFM
SAghEf79Gr332QWtyPABSUQblRMpWb68a5vMHmpqvYoEjHrEGy4PjKoTGX4HlAUfAdrMBGPvGFfC
jQPy3bLXSqlz8Y0sBQt+hDnCm9tNv0L0LDbMyE03jI89fMHKmu8SUXU1qnKWxDcRfWMoQ+5ykfkn
y0GVdKas2Qz9GCRYAQsKLA6J3bfW3qxb5fHK8x27q3D2G22tM86AxIXeUVyZPljuEJoyWS1RdDm4
JfjjzeluUl5o21stR1U53rWev2+qiKVImo5XrhdaBzn5VxtkFUgBkyPpFDkvXchqhVQ61NzVDnMd
gXkkFfESRVGdlSbl5iCzmlunzyy+o9t5d/a9A9pKXkz9zgC2B7E9Xx6jSxenH6Ab2XD3gLEHtJpW
7VFczKpnLoyt3/zhPMVYd2fbcLCYbqiHEIuBB8ZbfpRoAmifo2gMlvQUxcjUdg++9po8IoAD28Yh
cQOF64FDUfKFOQTAO4rquEBaB11F82vNIq84SzKsS8H85pm1k6gHtkVZn+Ct8lbcWJomD1YGrlEt
n8pOvMHqY9AYfmzLSvLsVt6Rqoh9eaWAXRL3VWXqiTzCKffHgJWZ9ysxdiE2uXLVg160HKITyusG
z8vTBaSBFfj63Y/Kb3ouvvVkoGIq8hGrKSxITzt9CCH4VdGa0YUTjlnwyryw/+AHvYJ44v5YJE8G
qZ3qc0WR/5xca8QDAY6Og0njEqptUGzOLbW1TcNuLt8EtqKBZDo485n+eVAjaF0/Re0QxxQ7+Mwy
CNyevvGyhgKXIcUJlT9R1A3CbRjvxA/AUsVvxMNhz2mTHI3M6dAhBuL3ffpEVl8OBSnK3WnDkwcA
Au3viod/yzwRfT9IWqeSUH4CmlEh5e4QzyITSMlMEDyFnz6b8soYsK8ovq7Ha4tIdIIcTfp38NVh
h9uNnxAzvIgkNxhZsuOt2pxzfZ++h1wnGjsqJJ4vP4spLADO41/MYq3KfFmPQZ3ve16E4P8f8Ozz
B2IgO+oWoWgE48KcRGtXYKqG3uMopjOvitHCOO5p2HQUCEOSj8w5wHrlBY8fQoOWAr4ntCaJHjS6
cq1T8obo60qmhWW1yaDeD/qsQ2VvgJAU2heXdZzPea5cbF0Ivd9AQyL5zK2BzFh6bqJx6kBN0pY7
60O5OEZS26vU0RalrQWquLB0XxQAGsyWCDVIFJo+xMEb45DPaoVxuVxEJjatLYAJH9f2kevdZHID
XDZjdoUqqgVJgitntbTqONeLDXqUqyasjasz+GA77pGygdLwtkhimsuHdzv6+59yJ/OfjMM55yQ8
E2qMMW0CvMvV97zHP7ZKPzO+R/RTPud09aZSEHtLyspQVfgjLhf94Ou7EUHzSw2TgMAO2hk9OYJd
m/EOS0z8ra3Iy6s/Tg73RkJooOevWs80kTl8KRBtV5SI1uqbfeB1hR63AXzgF75bYvHBE3+1MjmL
8qxWOEAuW5zdTZwWkMT2BZLQq/dj9GOqOz8h7kE4uydfD2AB6UMYeiEzFnsv2orjErRf7MVZOngX
tBAOoj1G1aYTDsspKgIEZkh4XaON1wFIp3Cgb8uS1NyRO53cij0zeNTCRXJeDuzl7tec/jC4IseO
DMLGCsSNwR0RDVcZkaywmiLOqsVpDSFnq8jLWmA2NWiFQ2N+76v5dw7S1MUhlXwtM8u09p+fq9ti
Q4LG98oYFFgKjzx65PrJ4rOITUCV1ZXXWEiexPm564zc5rg3txZI5gz5xhS6p6kAY6qDK/L26ASn
TbWvKlM32hwsbimoq85gtvVcgdXJBZfK8KIxzmQrzK/vPKZfaQjcO50rvuywdzXrlf+9K1Hu07vt
A8QXyjRDD2kOesCKU/H+2pLdIbeex3ZnMrXUSTiqKQtCbV6CNH0mHMh3GSxMbN8FQdC3qpwuZ+nR
DwEMwmPd6j8eyv8GlBAwZBG0gzeZIPTa/xsbVG0rspUWL5xRkVTTx1jtwC8NiUE56iFUqDC6AjaU
EkVHkw8ke+My9uj48be10aK59BbgCHE1ISIOW58ochjYe85ZAiJ+mc/nGMXkB36QJ1AkazVhON59
DV+k3dm0UvOSmj6OpQmEupYbUc2UxaWgq/Mc0TM1DX4o+u9gMYHoNC42h1uiaT8TOW4UEOhCjuKm
D4XGKrVDV6qUxoLWvHyWAZp0TFMTi4/cvxRsiZQZHkRic09421dMhwGA1g0JjPCmbhG6Uyxw+G2e
SoC0gfwDTwLGtaJGggjpO9cmuHU2R1WNY7Cr5t2G6+6NdFAurhDF5XlKifQVVthAhWAAY+/9Tbt5
8Upgnb1+cq/m1Muddhrl1OnJOFY2lLkniMVvv27c2jb2trVmH4AeZsXA0wlGZ57S8JemTEZa9M8h
iZSYAHJLjS1K1SxJzWKcrdMQ/huEtJwTmPG7gBi6Pt4bcelgnPweqpNI0QMp88KJP8hviUCQDjSR
w4YcPJ4iRUuIP+CMs0YPCo+99JwsorptcGGBqOI+OTMChkrIhyLRIkgNU8KxmegotUMjAp+C1FC+
IuIqLkLhjOjbM7Cuf4dyHtMzaKpKsUsGoOf00nB2Axw/BW1duTETjl46KBrD/YaEkJFYhR+ljKfI
7qGpJ3W9XmTKBXlOd/RfbMeFirdXmmrzQ73ZD//NkM9ZEX8nlX2XX+4SbDydTwS/zXO8gf+v1XRq
zSFDS5zjXZa7k/8BkgdDQ0ZYjlPNKVU/1tZsa5ab1wjLKbiOkNWFReP7bBwV+krpXBaXv3y3SnEX
BRuupJjqFikelpJie8+RZY5WrnugNUB4GsekIVd5CtSG03LbLfvg823Voxs0nxEBd+8FrfcGRN5o
bdCMsLZu8qoqkZDYPPL6lCqx84nWcYhDxM8xa6tH9vY62Syori3beDJwQLXJOpAVCLLr2b8ES/ap
0+eR2t6a3di0iRY4O33LwXsL7/8ILDts7jXv9LTfpH5UE+0leFZYOIUx9fvgu7kq4miZcEBybVQA
VXdJZPvbPfn2eAkq0a87w9LmqhO3xpWnYfQS6+LHmIGXysvjXjlX/ps9iSHHAQK8oiaqM6y9tKaC
v1RhcPt86GdHglvi+UUTLYsoH9p4wFTDvh7HTQsBEtFfsW9IT/e6cLYpDpgeD4Y6XVhUrlzZWZMj
gE1r2qDm0HHo7/A5tvshZLIMqT7BtgXEGm3dTcU6onDAK3foxbQbV3JpM12jLvqiIBeBU0C0Wx71
0Da255JFd126n/C2cBq4jybDT5rWf/G7hsMFSiPrHgI4IliDJ/R0dkSZKxhh07wMzK5SNpmRdL76
SaKeZ5K2osmzptbuxdMKELHZUxNpmIUTCPT9WvpfUtuxCMmO3YY4nrLlwJyH0ZFyUEHwAu2A5na5
g2zMegL6nDbbDm8LU+D8jHMK5JoiOJ36e9KlcFuP4w2uM5FQWdSOdzq0D8f/3mZqx0AqZR8vu/Qm
l+hE+q5DYcYQyclV25FyBJ7R4uDtx7og52LmItAgpcIrgKhrwt/gpuQaKFuA1G6inu9ZLChCIQV/
O+bHU1l5q3kL4keNLd+KWY3SnnEhQgBDRJPE51HU8YLbGyQD1HnDUsptNXPrOWg8gk/gU6rcKhpk
yFiwz5rkqaE74+phM6OmpBzbdqukxFdoxEj9aOX6IX7tyRAbxX6XAwBoVG7mrd1mg+efeCp3QS8V
7rmSledcRUMMWdepJjTWOV7I/Bk4peGyvTWJCaigfPNUKrqNvy9qd78Gb2aUtQpuF7byD6Rl2ZnK
ShxUlaCjqC5OoMi7ODaS0lfGUd3dcqepB5lUXKwAYJoPo/pyU2NPMg9NrNr15j4eVbvTbCcHNS6+
9HIF+oYVmDoqI/j+pNnVGcY2VPyK2htHeEHbJn23tF21Dm/YaMq2CSWUS8/XbftUSnFS5J+7D+qY
OqlfmQz6MFdQBjMsJ80CUi6E3/wHwdKdgJtQ8kS3pcMdzguSehqzx9tU0X2vOOBh4fCb6coXwNSc
zs7ceMktKk+vwO0LtFnYmYEdLy5x8JS1mS46/NerJbG45ARNMA1E0x3zlqDgbtBnLALlFO1UA/0k
W7B8CBPrc7JiSC6AFIWdymplo1uPNAzMyoxEkE9l4dw/lcp3ciZNaC4PqwBHon5MeL1YB9KL3KXF
2jDm1QkYWk6hh3LDDuEMSujVK8X7v4f9VDlN7LYUOFvls7r+m1qAtme65kG7HSaafcoOoVy1I5Fd
mncjrZJ+tojQiWkVN269OZ2mXFAnl2pm9NdTgX0I84sChqZFDeBS4zZHuxvP/CQqkDg0nW17Tgrs
UeB9ug53sqj45jkeBRManeNnCrW3VuKV74zSUN/v11cRaAXlaAfOfxFlpyD1KQ/uabDMW/MWWHGe
zXMdXdnoM85Z2TvVtA+HW2xYsJNZhMkx3QSv6BZrAgLHNknvFC90vGcsUcMLW3f1Z31BeFMI98Bq
AqG54PE+TL7ngv9EumshkMOAJXRjkRZg/cEoChowkKfh359KqvZGPEx1AEKmfLIP29DUWyEBHcrJ
V+HrDpMqgKiVjGJM74TkqSS1gRVRKb7UaJCO7jhwjeE7swOhomA0AtBvUp77dfJYz1EgQQ/X+85S
SfYDUOD2roIMHSMifNlaZHg+LRmGB5N6a5YIF6LvxQlEFUBCz8WBAgsx0Xk0N2n09IMdhLYGuSv5
hJhdp/fHX+CcqIeyfFGOLoQcrhJa8j+hF+g10xlOALlmvLt5D5EQeLss0d1JOgO41GKjaomR9ruW
iPRSrZ9i++fgltTlWsspRcsP+aKszzSkEU3DzVKry0Zu46JLMcddFM4BL4uz58mt1Bp9SoRIzCcI
sc3SMWshfqp9IgTR4hAPb7L7uX6Xg4ejgKlffN+JwgGsafoVYQ5VwplTxsevyb1oORjpc+vMq9zL
YZLPPP9RdkNFkn6oPFLjviU8CBr79dZ0UnwF6Ar+AUinAOfG3MZEjtLhPybodvjwfFfgxgcHz9lP
B9790iS4LAqW+eL/ryhBirk4x+JA7xY6dU31jYDYSaob/WMso7sdsPPjLQ1+R1IN76KoxyalGdC+
QtSW+qW/PwPf6DcfbK1u6fdyI3hzXVg94v9lCYcNRw/PeCyC5+SFb6v3kRuI58ZWSLAe0a9n/En2
jLCAurD8y/VzQC+UuSTwEaRlEPFjauXfQgRCUJnVMCkk5aTl8qptsYYMZSHXg9hpdiDyfc1NlU0h
auEAxD4jEgy/9r/jDhLPYKfrF/COtDmILTWXbU0kezwjLCiYPtkf3TR9BCiKxIbcEOVYcdjqdAs+
rTds7DNqz6xyRe1HCQHLqG8oq7YAAwUkkRTTo4RDSbeiVa7XEpIMYtUwNWM0RMpQuJvvjPrZooa6
i9AwitRL84D6eqSeiBH4qfTlosTNHYaf4fhDiJDnCeANai8A6KVInZVSljqcYwFlTkB069/fm+nD
XA80CCsGWBZun4McIIBm0HfE7fIPAJrGHy2SgP7JHlgsImOZtwqFIVn4g29lQiGw0lSMU6rkvqn4
dWRGE5eER9bd81xE13fW2VpiklaI7wR0eCeOqTEOKzV2QHJQ3BkmCx3HYxK/6ERmsWIAZ4myKemL
weZRfREM/1e+ApmlGlGGY0/K0Tj0aXitr2rZynd/eW9djEOQp8vhDooateXd6XUCpDngPdpPNAdX
caesrs1NSKWa0nsP2c9IOPNXxyaD+lOzicHQ4TRWOVQFDvgAcAjtsNVXFGH0+mDsRCm1Gzpqnqj5
pms6DqrlXTW+FBb2moET15FC4bPA3HpqbQ5wRrf33zPHOOKUmlP+h8SuybRqmg3eHIJ+78ugwzB7
OVGC/7Sv5QXoxnaWaB+naLV7fOSDblMqC9YZ4gkL/Jf3TEA6q+bsa5ifHe9q5QcoqBna/HiA+b3D
ncxpaIfX0J7p1geqzypAJlNme8RTloLqxD4CQ4xl4JQJ8HqugYTGNYctdOZFWmRzWGzdJI5cLDp8
C97N8Nx076uB8GlQHE6pgtEBjz8gFlf8OG0g9ilmx4Ftx6CfK9stdTR0KHpUyUX7fIROJzSItHoK
bjqogoE9+mEuTkZdHPqXyvJzAm0kK6hhK+lKRFqfRGTL9k+ZJwzJkvEZFl5ON4QvS6lVg9frd7gs
/aSV7wijmamj/fyzHOnMYNaRWBH/EjYVPXDddL7p7eqsuHvGoxw9P6b1QGAlw5wF9H9kPSqa6AAV
IKF+LAXuCQGtW1NUDixh571jue43EsCG2ai96P7dnnIxKChPZ1B8TVGZUn3rOcrGwnn/kFkZiN6v
VTDUrUCPbS0weVkWL8FfQAG/cHgbAAq0y7CG6jSTWisZAKU7ZFt3h9x8dL5GSO8Orcb9+ueSu7r3
2ml8vil9e8ApV+m16Wk5KiB9Bd5DhOUX87Sx4SJSuCd66p2dZ7nx9PVciC40+FlIlhrvVKvQZ1kR
DiQK3JV7CEWxd2vkjra2Y/248984JYsKYcWKJrOtD8rHvuTB5M45ppmk3x6NRGwQEwYce0OcxG/I
FVDWveGf8P6lz0UV8P2ap4Zk/Z3EiH83ji2SDTvQyVqqMuP/vmaQmLmFgV8h7hGhlID9CWBTqV5A
5QTMzexS7scEGDFuqTH8iK4KBZUH7rrzrZ4QNzCfMOw5IlMcxsdHb5FmC5k01CqNxssdysNy0VWz
XMoYilnF3r3yAHtnTBj5Gnip1JCvmBhfkSrLk+TwHRHu7iB+tbBKvVgzc4hghRVrwE0YQqdj8UHC
Vmdlao6gp+jTjv0vK31lH3Fs8ZSO6lXwPEXaK9eKQkTZjaQzPhKf5SUsH9AnXv68lTIi8KaMLqU5
Tm5yijEfQU9aCCKxSJi+FRkzJZV7JEB+KTHfrbjWml4FF2aXlsU7iLlH44FyatHmjnhBEYm/RlnE
7G3G6VcmQZiujk8VZyBiMqQ0mTEcvL3aV+qYWgqWONMbgYCWEaSSgAfsuZS9XjV8KLtNX/7qpAf0
SZ9hmX9s4FwXVXEB9x6VrRvi180QOUMHJ7D9I6zRVN7PYymcfaZr0XBXIYNcGBrVhwbU265U8M+S
tVeOOBeajLclnD48WplMzPw3514w7PG3GcnsfdPtRKF9ntFVHjC3NFr/zraqvf3vNzLQnB4VZd+e
i1MeOLyKMcjD9Nc0Mc3TbbkKTa4h40Nrzou+Hd5Own4Fes+R9NNP2nMsG5gkFo4BpeQVE/NJ1gBh
galg8mpWjjeLSoamJ8e0R6p0MhwEOulUAUcZVqKVH5pC/3sBNc2OwxyOLYyz5nXroWQ/Dl9omL2q
bpQ6FUS44M2RPoeIlFXu/8/MXO+VRiWUJItGJaWrbefDNETeVPlETD+CiepJeaQ2Nkch7PDTs4ht
UycFiL+M5G4JGUN2trImU5qMEWqNyMB5prZDdVhgRIGf92h+R7OZQgyDS8GBggNx22XgdKrFXlV+
8rg7SOChPCslgVdBZkkifXcx+cGBofCJrFrT937AxGTEiu3wUj9lhGHxwyD5PnNR3UcIEE6vgydV
sjHfeiOeK4y7PTGAniqIGLIq+9cyu7o30RYPENAAKURGb4ygpVnxB1Ux/9MzKncOncrfxP872XNr
2d2j8QnIIgLH+ifEqDPLqxLezcta6ShSbhuOrIyEqMEKD0u2eyKHBOdg+YlszSdjKhlzogP1HEV7
6gh1HIYt7ku2Jz+rJQSID3AweCijNKw0f+s91lc9G4DS4cRSJ8ZejDHk9T504S19U3IB3zX6aETS
RxwTjZE0QRcXOv9NCTI1PLbngwR6E+mTknd4+SUQDub/fhxAlS80jMWKo28Ju/yMk+x3nk8natvo
sDBVQQ4ow9LtZhkDbaYlk2d7xZEcbrBrVS856u2oPN+mLOH7JdYkw+1/QvHQO5rpYl4DmDJS9Dmq
Dg86BQv5X5dXI4BcF+tap05sswyVgZDYgzAwoz0IsNMY6iKfNoeqNcTXNs+aDKTP5/R2YwD3+RIL
MMkJE7OREoiOx8jorbv2IPYXuT8NU5vZCI2Jfqds0C+e6ICH9cNRRuH3q/VE2NeAVDn51+xNGBB/
vr9D6jMOZIAiufOq3MFCzsDPQFM6/YrM6+0aLXZObjVRkIf2VN1Uean6C3YluyX2lbTfEerR2H2L
FBELXwEcHPX8t9UjcEo3ocjBhfI+Jf6jf3GS/8lA1IekJna4+R7WPVB3oVP0787JmlztZ18pfjjy
8UobixFLzHZv9abNm/GmN+AsAgVW3CYq667JhREsMj5LwA1jxMSAIlrbCOLOAPCPSEEyMqNP24pG
QPmA4wpIFnFEQdg+qAb61IIGzxLQ6WG89LXUxyNCxHlBiQ9lUt9IXpawTaoxvfXxVHjinlSWyXjX
OuKIvUfHohTPQ4N1spbEvsuyS69n6CHzTz/U7fWaO1FTwKg8AAllNn/jaUdqkOuFqJy9pW0WKdQb
4vhleiJw1PRWEzo7zDC8pflrFuynqhxyG5sjeoGh/+ZdPqL9hqoJsaVlHj23rOQXS+sJfDU78+3T
EM71tQGrl4Ubi7CdIAZ6hXWH1eci5gaYe0HwLpxbioquEV7ZAm2n323l59aLKu0oqawqApeGCcC7
tLYsTs/mE74OKzfdHfY5OvjxADDt1beKSu04SHqCoTs+fz9R0BrqA5QTPR4zGfzRzZ1HDAjUsX8a
6/U+lzMay+xSRRRYcnitDclsxl9zez5KqS2LXFnIhv9pAkdrPvfQq+eLJjAojVrTpl6UH3D2Hin1
0mdaCda/9uuTBQxNIO3cZ54bC8mnv97DXJTk4CoDNCn1QSsCYUVCD+Z3eB2Y29mPpOri5Wqx1PHf
rgB0fmTL/xG2ivRXKuX22z1P2zh4e9h3G6jk3o5MLnxqg00Qz2TsobkK5Zr+Pn/IVvfNSO6CEeJw
MmgoWPcUSAMA8G5zy6VTKQh9z01tM8gAb67/gfWj2scCHD7NdfdK4QKqLTmfoficC/sFqWNyK5Hz
sdgfksNZcf/DUCHggN1WrWXKdrmtdgC7r0xYLHJ7hMBKzbGtLBHVXsLVWz0NEOVnHmxYt/sQSSj3
dIGrXlmdVXwWRSCM2oKjQMBmm1Yj2wNcsQwITiaNzdy0rIKJ92YBJpAOtnnoogga9dTJEuAvXMFR
9P5h2M2VBS9wnPbDux0o+KhLvqDFGRyLqryrt/cQZyR0CAiD/dD01y/lIqaLaYEbojW0wRlKrGIN
a09mp4RJJ3fXpit83clGRu5E9RKJq8wXM8ttMxeLDhN1nh6CEjwcB1ViaNcdLN/UpG7TmdQ4Dcz8
0GumaTnvhMGW/Lwts7x783ILUFE7FF1LOkernn+Rl+0fyeyBu/dMXvz1XrNGY39bKC+zcJvNZBA9
NcgVQJ83TpLbP3B7n5wUwf9pDZmR3Xu8wjoHE5CB66RRIolxfZHLCHWsYUdCp4rXE/YrcxJU3nFh
cZUIyRnqe/lz27ilwtNw8k9kFY7zHI74h5uetuqMW+eOeDkuUxHd8ULArGgjov+bYNwT6duVkEX+
R15SmYWSWvpf+ARJyOrJG4H3jmgfUmZuTCtzSb4riPE3qfwuYvkNY32ICObjqp5DNJxOxAmkak5M
yuAO+JI0BBQwlMlVPcMpiobpYQPU6mlkht/1ktKdNv44MLsC7YIjMF+zluU7NwEKONlaoLP1/xw8
apjlvPb1eAz0ljtqqKIX6YfgQLJzHXBccu94zM/kZ+oaNpPmo9EOOAMb4cw5sYzTniyeKVzcJjOI
1v2sAY1wxUTjP5YtpnKW9rSramGwiuuCPH+n24MiSZ0MP/WyaPWZWFSwqowlPEgDtWShcIGRQaxn
4ZJ3Ag98sS2NbdD0yO+0kdsWYx/dhTs/3V1JI+Jzf5NJMfxnQOLldwpFcOfTKMYw4ncFix7h13Ag
1pVuatEzWAYrb8wq9NJq+sHOjvZ1l11t24vkGAkyj76RQrNqCnAIq7rMJmxTgiGwEJDCJlBta+GP
wvNENBrMwMY0iVXv87syaqbDt7MgkHDxkWL0qPXB/Y59KkvJPTclzmIMad5aRcYUWip/LyLlTuck
pACW7YsPrb9Bi33Ulw8V7qdoRaGrDlRj1Uzb4A+p4hMjYeAFeFwVKxhCMRsFqRQC0+QPe7iAqbL3
Gq02u8pocFCnZ266cjgogXGMClm5tR44X5x0RDlAP/5P2TwCgI+S+16gYh/LbodMbyYlP/fPGhdP
1s6C7HD9MjlKg0+zclPGRiSlL078Q4fUNIc0Sz3hEacPi7IoG8Bn7bcAzCq+dBZnaGNck0utRB15
aFyTaUkjfv19ofwndm5RdQm+OxuUTpMaGhffRBSckmWcIvUGOBNHN/EK+7n8wlleuHN7ZmseShE0
VKlv6E2S+4Z7NHRcW+qExQBvF4q0LTxavcHvXq8Vih2VnTgchte6lpslIOOa9M5YM7g51MYZ2nBj
pAGlibx5I/5kzMnwDQVWsH6OhVfp6DRaagAOXtTOxb2+trzxdM63QdlQAf0dnmXRE3QAr4PIiwxj
tUBPdEjrHIo2f+fAFZb3ntanUWm6ZJtmUJz/T3KB1KavFkDwSg4MFm/KywF8Vi9aup9GE49fHuWH
8DEln2LXsMt+JWvmCOpdhw6x878JzFbU1gBojpjyVGAkD/s7Kfbk42usoirsUSsfRC9a9umcqS4H
vqU/behBM+do2PqDZ3TIFXYJik40MKbPbqy/+wbD0Ajjw5+n6JTDrRDkmKgFp7QUaI3YEF+xxcaM
R7gXAtzgB9I/ZjI0VhXlsBxF3heKWUWrr/26iCkT1urptsWOh+FO2ooh+muwvMUnferaPXzGroLq
/poxWoNmqjLg+krr2Rikfa4n2JakEEQbAv3pa0s1qxH+aLT9nPT8qjMP5vIpN4khke8vbEgAsn3i
NYxGCD2Zyj7dnKJDYZ5L6B3pdc9tibJEm8i12+FDX9XuGtr0q3wzeW94+QVOcNa4W0TbTAlkTLuo
TLdELbN9XGazkQ2SWec4GcPu5AUSnXZbJ4RTNGjEuSwYVTHmvhwrEMW8DBIvImeyQaNsu1aVxrvX
1sIF7fCrD5cFqOSIobkZRodwuCw4j6kxYa71cAATIF6xH/NJkBj8VUxjFB+w74XiKgMhIdhDWLkD
sIXudItH9yMqU+TWRj5MaepWbBRexioqk68iiVApn9pJZ+L1IlWD/bka5dz6vad21YQVXHdC/9uN
O4fQ7gmRdSa1Gsp7squ5aDAUj0/5R45iqmUntjwD06PjjQbwM24iH8MsbmfkEaaff5v8hXQhP65e
86yEGEpAl3yoEfmUCHywQoINCtcedrmMnb9Vb1TSgDlq9emj20xxheC+B6ru9OMz+rOBFHBdV1aU
DJYQbRgiSenm/PD76UWUk+ixNjORntUz8wvPITAZNpiasy3Cd1XuHk7CS/Tb/t+9kaq+XnItgSeN
wKVFe/tRg3/5ztyW5C+Q4BAwO5MzVacDjz7taBmZ8nO0OtvLeAFjIdYODLBJI+mo/DVDPy/esZSt
fA6cslkpkMStjauDNbD6s5ya8PpzsfCn831/AqhLfg/WLfVURE6C90kR+mr9ni3xVsztJvOeA0x4
sLMaWaYG10+7oB3Gy7fTGsNymvTAPZheuTEmKhwNcrlYtuWFJK5Q88KPkZfd5MyInN0nEk/B54/I
ile9ZiPwp/z3f4emk7WkhLZnz2F+/jCkQlGJSUpPVb5544mknr4WujIfFNk64x7C5T7eZ1Xy8XW7
sgcIGuPEQ8LNM+usIdoWw2a8yz2gSGvrbPeBjPpuhE3M7NSl/bWZJfblRtqv4AvPCJu2akytoIZF
KOAUt8ebsR5BSR5t3j5dCzhTV5U7aBWrTKSlxZgQ0AwSyQM8o3FwzVDlYQ67eAjpxPHXwVFCBCyp
2RKlJQl7pmOncyZ3lB676JHHmbnUfXoRbZCRmbiSx+MbQqFqDe8/QwdxwRQ/qGua46tnNrbKXrBC
gOA7vFZZpbsSpPOMJn3X6bxwCCCaQGycD9TzjyOPrislC7MCglq0XEXYrZGMNiUAsR/7+huyrNEk
gYYOmlnaSqgH25zmaXkLdP7ieVtAxjtUhBzMQ8OomfyI2qujVwxKpaufpfjRdC4lIlbUvbltYjQE
xmJSLyt4QwZmPaNwNDPVW0rQ9vQUe7B4NwIr2ThUDcwQdB2Fe3cpxhtos3ASN0nYQoeJl9euZG2V
lvbaFO3K8mRvFQIWY6r+lCcSZ7xbIzw3+gKMWdOXlqUt7F8aKW8R4seXlXllMHYgklzvQvs5iHdE
JGZ/4kPJNYIRRv01xrpfvJWLhUZmXElrOjbK6Li2CpUaBiIf6KhwM/nFMQ0qzxUoR4LyD33sLcEt
uSqO+/8QS7HHCtM40sRYEVsu94Ui8bz0nDi2VGtISi3LS4uAnv/uOTa5alu23PGZDgw7n3S5q1Ro
Fvy08J3YXUBMNNLzSak62LhEfFatnfrg32Uks1AF+fMRvZMg9FKNYqZzY1xICuSvYGIpGOz3faVU
PlnacpdDQFJniKGgcdnHavowcpjUBOsUeAJ1AlMR1aVTRH5AFRdXaJvT+oVPlC7A0nizy/aCH0yA
OFXGvAauJmNHt3NLxMEfADEpALE5mjI5YcRdNIhvA1UUpKufxMCb5bTedVN9z7el0ew5/WROK2mP
lX/wYeUMr8JhyVRj2NO/XaORXJwUYy8fvoMj2b9AJcEOCxRb9AM0qj/25st3i5R8aFzuGjtBvoHy
TTDOlTu/AlfhWTj1FuvB/nrV14Mtll8Z7gjxj5T296wFJL65J8wZEPTcEsdK8yx/1vdU9Dw72Ko5
UnlYVX8xyWty3BcZk1peTq/ajFPxt9bmouFMR+fzAKuBPyByWgpe2052yvWJ5Ag1UoqhGZbT2oi6
kl2cmUHTxxWDNYbfdpsJ1y0z9ACQkxCS/MIkK87lYjvY5agENQv4vI2FPWbiOKYgVaG+VFTiWzGB
ZFAfFXpf4bt6aJR0AZMaPZu8Y83Vl4ChrLq1LVY8FvCHRRbbuF8GO2ZHWwjwZvlDnmMadbt1+tUj
v09EyDBSLe8FCKsRIu891G8hG/kPjLfYoZMS/fDW7xPmhqtEHQoPdLPDvpdk4e3Ur7vlsJZeVBcs
xiz7k2ylGF8+uwkqxRh9AfjF2+AW9Wh/goZtoUNJfZd5du1Nind2INtGfsC82UpA0kHukpzDq3OK
xkEgAo+JrNfsLFv/vo2vsK4ppxut8nNCOL+iM+0UocniHJ+ibj64y8G/DzPwlBFBIbfoCe1PBYfS
5UNY5QN30OHR5sy9OnjUgNu+VZA5yU6jQMI7Pg/HAeBrPYQjLvnN7k94vdIGDFeIBxOjkWZLkHZR
f9/AdeK6Bo+4cn323Yv4eCvTmvcyHoQogb8QWog5j2oOEvhf201G6wtjZoc3gvNYnt713U36OOQc
PqJFKUIR7m2Un/cz98PLwDTj8PYK8oqzRwEMvCXfi8DRQHdjSIwmnXvyVRgOB4iykj8UicdOe8+t
YQvSC+NahYWTDUf3i3atgj/FBq8ldGoeehV3bi6QFVkcFncLAMMS4eozXyaae0TvHysrcNrkc/yI
KKbVqnSMOoPDcq5ARkRwEkadniYJKNcKJrAG35rhvfnRhQgSmPIIn69LvwaR5Riog7kP3J+gos1/
+NIpS1XgpjT2o3N3ZbQr64xgQs7Qh/p3d/wfSx4UKax8XeEAdatmyEpPI+MO36mM/z0CLUtod+Ha
PTfctCN0xvGbQ9cb2cdrRCQV2JAaV5Rri4f03VKtJDuGS5oV2K3lOsujBST7qLAneCDkCvnvFutc
ZZn4qfG7lY5ujXLqBCtKftRha+an0CFCuUBeTirX6+bPcKcdLhVxHmCIXfrOeBXxsbyMeGw2p5K2
f0w/h3evYwXZeo8E9Xq706m5DkXsE1tg2uHR0lmM9YVKnsFbUlC0Tz/fTL702iSvUOZpFlSnt6bM
6jyOSEGvnXd+DQb1bVyc5+4mw5zXEEA2FwiK6mHkbKcclAfeSVITjLPin/+4tnTBw5E5M7Anq6G4
ABK0ZdoGhki3fUSU8wbXpCusZE6w5Bdjq8QqJqs/Lh234ktICqkKwSdAuG1wEcLakxH975CFnFGJ
gjE6ocHXs1CE052CdjuinxN4Ez92UXDiprJH685y/b/ggAqhq0OG3LuOAS66ht17f/m2bfA/AhtE
xWRNVHwMbX+cnuZRmgII/wlB/4t5KA7BkMA1vcAGCkqMUqyUKiq5bIo7cdV6uUltccqJiYR/ZE5I
XJSOcK6Bfohb2ojGtjIE3fnGBrnOUiNDo7i+ryH2DzAd/Lq+mN0D4M47v39sNijYzpHvUUT0nQCs
R+N1vUw0iXSGd0Yn4GMvIehTeXf87Lj0F/p+tqZy5iikeyVGRWkrCy8eyVxgrFqfzmuAFMUtft0+
bvL1bqbVh1X+zkITRRMV0oDnLrLQikxB+U2ROKpHm/Rr7qC83L8S2AIAUmb3WlXOTqS3Jx70ooef
5G1LKQK7nYL6p01Yh38tUXFwZoEXDCuDxdqC5Or3X3AWarfBqAHR15Yt65DymhFFZfFbnTN/Jg5q
Ci04Y9nn9ji5JP8QMpv/oHPi4xyF7IBfBr7XJjhEGyX1xwX/vsFNc2BQPJ6R3/Ew0EtJcFiUZ0wL
VyE6e/kSHN0sceFn+sYsGTHxl2PgJUAMtFxb5m27wpwXGPeIAXYD0MucOH3TBfLjpqqMlCha122D
xHOFMq9alW1vfFlInurtvzbXpFcXeCF/Hs82eo8nfBNoEMyR+PLpXvZJfYzHqC7sIDCyx2SI7uX7
X/QMCuM6rBgbvo/6ZtIzSwl9z/qw4zW6Vt02ikWA9cuGrsrjG68k7P2IVOIIc0GsRs5EhjQYY4Zv
a5tJBCs4ZuHzuD9J13u/uX3AfyHI57joj7sNj/WtmsAx4niv97cU/SfbK6rO4afMOMvRTab4GZUd
cuPIIU+bTFqlxTW0X4aciO7ddwpVLw1SDjMOvsTkbuiCJ7nGyFWZ/VKip4eaB/ibffFbHalbDxsp
M+OPZj4az+Jx9LOjmBdG6apONuRpVqcNYQD72EiOTGLpG2tnzzGu7PvPGE6jf/mdnJJLqWTFHQGI
tnD1XYvotkgdAiFnO8nkDjWpBOP6GrpCjziws0+SAxHSYbg1bhwYg8K3EjMkUNvV0LRXXIbETFIW
42j5MhIuQImXK2cYxhD6zEnJLPmV537OuCc2+D7AQl5JBv1A3iLNijGiijOCiitYPZ2HfpbHH3KC
jDqJEmMOn74rsXwXihHZQJWfGFuYraIATrVBCcDZ65ndgvIZ/7WgYDTU69HMLjpWnsRYBfVXf/G4
/Njmvz45YGqbnbsWOproRLMPhxOQRFb7haDp5li2bYnHasLwqrbgm5mvLJpNXpp623sJLMUDZ8eO
uAzOgzM6C4/iSGTqDKO9Ot1cNzql/n1qBHnp3qoSZESJtHzJvWO9cwTz3nmFadRQ/hRuJkT4Q1M5
tJpL9xorAxEFVtIN7koonuY389hMoFxse4UAt70bFzVVy1oPQ+Rvvl9gq5c5iONO6DELet+A71SE
1uabSsDOAmrSwNYHsbE2d4nHfR/IhVDKNrseNDbsj3auIC5MvHVrhM2nVui3T+kFJNDHM04YzKGh
WH95iOVrbGN0wgQI//w2AeBmNjX1SrL6VvOy9u6T8dsEe7PJkLtf26nJglmoHI45GulMfNxdN1rP
Q2Fm2rf5qA1KQYV4YQzOOP26C992M2k5DjGkBGosSJTWIjUdqzdn9ITEIPuyTZOljGzZ9GcMHjBh
RLj+cjOm0U6hohUaR30rN3Y+auPVS+ctUyLr2pwWAYcBvU0i1e6w+tJIjdXhlmfrNsUio6snPyJU
CQQZ7ctAkklbb4wr4K8paP9sLCZ77ld7nsWf1FkCkKjWOm7dOYprxMpAD55iKd17FbWQysqHV7b1
bM9zAngg7xztLq6JBcV/jlpBiicjyefL5lXAQeuR5KX0CsbovLwqXcv79JlRtzoLPgodUCxR++aq
NMeRrjTXZIX2g8GO/UzzwOBEoHwrQcV7rpTaeCMrirB6DJhS4p11hfS96FFijZUop823w8AeK4wc
nGuDwIM3aLOROAvzXo0MTNVdJ8Vxi8wMPBKp8mO/msJhhuBua5FWHpqX0POPtN1GTHPJn38Ym+40
i4hAeC56HvjpooBz4ngCltIESJCWQfni+ayFWzKB6GyitRBsIBOZxgEW6J9jiU5/1u4D2AwMGR1Z
UJtHM6nuN3bVFbBiwFONnWYTRcIj2XEsGSNVTAJC6OajFTZfOQ3qRDZv7LeyjTKflgQZ7JjNECDG
UQy2IpI97iY/7Q/TgfIx3YVJaUZ/pIfJ2zim4PazDsHJapp2HYCGWAe+wIDIVG0eOIqWgHtcwNaA
V+glr0hSdqq47kHLqTG4kRjLn3WpVRcRnicZhRY2SM7cQ2qDyV/E4MKCj1wnSZm2yYOm2ghQE46b
RTolIaW0NiEETU//mUoet8YSwc1mAUW2zPpsj7aRTTK3BzGVkQL+7/kCLfsCOiq/XhrgiGAQ7YqK
wAYjKyKtsu2Xex/wR3aMb3yqxzHKZUS0eNRVSxf65WNpu6/17wZMI6loo14tjOLvEBR6SgeckbiB
usTsupdvopgYtajR3hRpIpKB5Lw4vTbWmUHqSrd2fMchiS7aVm1kcNBx8sp2VmIdayHHq0Wi7m4S
CLN3wGLx1i7ZL5SH5T1w3OkCy1S8ZiwpLF+TzBXjIjwIAR73DcEDiIE6aeMbemTIhgG4PpJHJeow
LeXORRdZ05XD/mmRjBTeobKOcfwgUZ9JimhfFyMAMmZFZULMd1U7KfoX3gaApKZCdFKZpamy0BO+
hDEcdq+55diQjV2u6JOps/DH0ABK1vAaW0HNR/IHTPELlTa2PtxvaMNBefv1aTi8VY0P30DrL3Us
JBKEYHpuBLETWgaB1Zt1gJVy4pGbbnMx/jdo/uqTEBsbpZyMuK14UFkxCZj/MPzOS3629fKrYvym
E7mkQZ9S4iDKLvg6giiMV/9kuvwEpu5KwIqcqlkHOTVd3iCKgFi0t/IG+3kKWhEP7z3TiqTdkKIi
zYTCFltitivUgJgwQEwAjS+xllCYRBmKOz/YuoRwEfvZL/v/GTHVE564hGEEAXuJUoMKntamtRll
s22ePXx66SFZbiUnz4sNWcDSKmtl//rMCzd/oif8r3MGDvP/wLUi8ZpaDxYwRZl+XPE+Gg8fiRxb
T3oRIG5+6Ax7SG+6FioQi93Db1Vks9Z3ms6O2duKh/wJi1Syfl8YYAaGko/YEHvlMzXm3BPaWU5R
qiaR6rn+CpC1/eLgxnWHfoRQhwkl62+haj5PdPmuVEZGAOgYPV6NwgMnyTEr3I8/rViimf/pn+oG
1P0TkzutZOIowpcJDJ+8zH59jX92wz0DFBc9oe44J5rNOG/ZWBfUkrW/FaadwDAX8RY8CC7rGxCP
zynxCYVQb5hp8MpNdSgWRIWVXKFr+mqUTFfPkRfngiAAIqNoTF6tXnPeMzhRHft2WdJumf4H8XkI
P2UXn0Zp3BiP/mZyX48+8HNAfLO+WLxgBZYoi5999OBfiOZfBVTx4LAVfT+66ymjacmvwf6p8gHw
Cz237UOtmMga4TzmkJsNd2107tS/MCb18HwrGF+nXc8Wb8vtea3gnKsPbAwXo09QdT8ceheDXP2L
f/LGMPsybO8RFtfk1s7DkZLvukPp3pRGewUn/qPjkOA23Iwo03Imb//4KjlzUyX4PYIc8TOivz5F
dLYQ/1Ulr+Xx5m0wxR87oD4SQ+snqmfr10xVMpIzE9ZugjWirMGAyJazteCh0qULuNw9JYp+8alV
uCifM69E6oAQyR3rqTZYjUDNIHLmvTnSCm13hobXk7UGiyEEGAto9AkOs/jsZkoaYlUVqRmuQbPw
Ow6rPgR2EPuwuythR3758Wj94lPcUFsZly58NDugf6UNJAd9loTH+pR3lTVbwHvI8AFyGe33NfwI
59E7u3p5obNfbBX3zKKjvCyFo7MjgxpSV9w1DhfJ5Osh8H4VhaVzM4ql950oTNI4GNYwHAy/cxzP
bhy1eFa50igFzQy8TwfqhtaAdQNYHdDVVvsqjqoJGA92eAsrLOOkYAtHgbO5PQQtZHOfjKmbb+wH
DNY1ZCS7fSvMKS+yzcZFv4mLxvD7mDsL5DbYCiCtXApJwAoiPIWEZRR5UQmCLKvVhTWQnc+Tcfnq
E47rV+PzjBoAfnAKjJm6gvUeNhSI0+QBWwDC/fByMlVJVrrGrTTQ/gfHenTeJDEVnXg/Vh4+9yu/
eBchxHaRRHyTkkhA71WWPhZHjx7RQLd1QZptt8vxhFfDR0r5XrwEG0692vhDFmtV5q0BOKH20OuT
YjhOuQxhOn/oc0IUcZi+9JfwQcm1Qnq3RcQmFCX3j/I8Zmgwh2PU7gi34RAGTjE/OekC/T5z+ZqP
hal/+YG+OrneCkObOJOnS6gQhjg42uJNwo1p5lopWVA5GGy8/kM6QWDQA6UjgMNFAKlQftSCAP7v
pKLI7ityf4Cc1L+hdHlh9n3A1Za8HujLKYIxegiTAFZCA0w7ENgb7hgdyysSX/UG02E3V1E0iv2J
nQVEJ/gg2RRi6NeiR/PomseOwDFn0KcG7M+tSwh5KoqqSxL2LD+VY5UNAjs8Tj1a0X8hdBS3PWq2
JToI10A95xFfC99wYYi/numOjWBwmZ9x+IovpPPZ6qKXCgXiq06zMSxg+faDcJqzjmM+2gUr/n00
6Bh08HCnp2Bp4v+jfBlfPJMgAVBwhh5ACMKpjoaP3tuId8Fa/7fgNT8eRrmu1tEu/Uht2lMqR7HT
J8bz4W0miIhqJ/qJHotjs5HNTUUgODcBBufJK0QDc12EV+P6gx3o1Verx5dAhggEClxd120JORuE
qxwaz7ZkdT7WncqjHuW9v+MSKjNb9JQTuPt3P7Wm3/Ko4ic+dModP7IbAnO02R7U3ZhQ2O0dCF38
UpBDSBO+rAH4Uxz9Dl2g5+ZU8Sk43m0+8EtLWadOtFlQyBQYIwNZCs3CvZCfxSgc2uHj8I8xZzSn
09yuxygxtPM7o0hNoZUdbuQcGJVA+znHK/TfYdkZ4vnmBnGFYAzu2JoVGPak+OE0tr2G5aGfWFwE
50Jbxruc1ELLOHxVQhZ5XrxwcQ26boqGtTOFlmUff/lIqPs4FHFSvrwIV8ie5RZJDEdCVdreJI/O
E1WlIPGFbThFcurE/WoXaPPCWHtvMP8yX4DA+mQp0vOvENHctwKYJRdCp+FLwrc3l/5JRF6Fzb3c
2itaug8cWbA5kTn5q6x9CNXieQ2lOFg7A4NhAIPS0RYv7r8f0rU/Yc5mZY8EYh2yvL2Xjs6Z8N33
/HD0yG6AC1odvWp+yA0pMt2ELJmRVq5XHd6/YTkN+5oVPivNPioAopkLm7xwXLo5KrwXFQ5+PXaz
E/odfP+XiJodDkENJS3EgAHan0Ek14GE4YFXuv5L44+oKESucx8HKJc4VNThIf87VXyV8r7gzWYd
NXIyg4TVZH6AoXoVf64UJlfe8FV6+WumP/xb4NM8zgb1ob1dsoWNaZkOoLlARLHcd/9yiilxKJCd
NT6v3vhWh4R4U4FCctlyN6PT926AIC7LwlWBP1l/mulK/ko3Pua9YcZM+Njvmm1IunTtZwgLxvoV
2OBJsq+E3BRNK3HiEsH7b8vhivwO/EAAmtquUpziVsk5/155Ica4gdRElHMHA93v9U66p5OSjJpf
cK1v3/lABXvpEIYXLZ9w8zEJZTjq3bvsh/L93psXMVF/BLxu/1x191eS8MVeRZxPWIDunoGnvvEs
y03qG9pLkKO+9h9UPSv1y60GMTo+h0AUndPAh79nunpCksf/gQmLt5DUSxNR2pZfrpCy37fB+X5d
bJYd4tNh7mmcQXNxbsLk/RI6zvTIJY5XC8SQQeJw9FfAQzTYsyhpHF07HyIKpvgmJtE/4TC6nvrD
9CfnBokUhOViMxH5kXg2qRHj7fRYH8Y264lHbrvrZkdINB12a+TIldjo0x0vHECXFofDa1Q7jMJD
Qp/D7xIymDrovrOvBzAf0L3DQsRRPecYGQB+IernZH7/V8dZkYCwB+g1PCBzI7mAhy3P8P6YIQA9
WYycbmVRhUPht+4tbM8o4bMggr+Z4KgqnaFZRhULP964rqYrNooK584gEvqBXPGTmjTst3zF+1HO
5waRxez0JIpJXC74Cxlsg3QT2hBFkhw/oYQdTUXfnaPgmemQDq7r1SXlkKZ80QICTTBYhJ+5MKWg
GlN5DGosXfPq3gki4xJyAdvbqb78Di9asUetJhiKVuNCY9qZNoBRUNCf7L+ZDeqrd+05k83uo0Np
ytxsO3h+t8fnMtlqUb7/FWwVswCKRNbheHMHDreBXUn2JB+ZziFTR0Qf2lLzzp96xkmYU8cw9V9d
HfNgBIW/VitcLQzUOLGVoYr4GFB8dWjGyCCEGxqoK+RUVTxv75zSykCUaF1nL3n48d2kwUr2k7bI
KAEid4Qp4io2aob41z0y+Jd/ZMwSY3vIKLquc62wa1KR18L3mdjRanePX1jqYtLvuCYRhwgkE4Iq
Z6vVdilxtZfon9Kg0MLtsg4z8yTRvgRpSkfc1+4rTqPaYEGN+pi2tZC0SumaGOTYseMgMYiUezXe
miqpyoaeFFEMZUuBUcTBURESg3KPddn3nVaxv2CiE4mg2h/IIw4lFyJD7ggk4TH8d/wfnjL1V3wx
JZY0IfR7yF5fvVJPckaPLZzXTRQvIEAMbcH7TDpcuIv259t0FZw1kjBG0wGiY4XMHO5SEjkDaXHl
fOnwTP977LG2di9fJMZb3e5HlSw0qccnMtSm/11CFBdq/Qv6x5Sk1RuwQ+y12597eFIyiPNqgVii
NYkk2Htl2hAtXLeRiFjO7E7x4PwzC9TOy36yEX27t0vMDcayXqs+BClCzZpdHcKB8KqMlQ/uZVa/
n6lOVxUyed8CxnqIzUMYy2bzvQ+McfqW76yWf92UiuALZGQM8iU5ykFOsfSD0u7mId4sHldSpVCJ
RLH9Y8kUV87Jm5qF+1b1NyRnzSxkQs4/ElCEtfbs+ilBLorZqlVbd52QilHEOY4rvcii8SI7cLFZ
YC6wf1pkDcIv1Es6qLjzJvCbcwDShGvoymnpN+3LYs3hy9h+RL/EXr37jg+C3s2gSkrBeVXehtle
O9yuWxsQtJu4TA7iaXJ2eC6vgMWaxix4WzZlD/+B++VYqjioGSQyBnVhyKnIwvc4lJ/BLHNdM/RO
duWGV4WTIY4uUFzxjgPpK0ds1xiTUGLQLSEcgXAvQo594o9aYFxNz8mbCEqXjTyUCzmdqib/WNQ/
05l7f8axrTFkrRQXoahnp8eokl7bUsnMiuvXkgefc0o6mI7DZeWPsGwZ1pJfnErtl347h1xNM3+s
4lyIFOb2L2iEfLhZbTYUbqAOqa+ozoHBmnFLMlBuicJlc9lHKzHDzookm2Z0OmPcpoXaaKUZ7t5U
/imd7WAyKW6jo3f1pSqtVqSp5ItqiHvYfbVgKGftzVzK2qIMDl+mRBgyUaJq5VaEU0JB2AVG56Bc
l71CwQB9DalmM3xJ1oZ/M1hRktsUYu4MgdyxwTMs7U4i/Jg66TCiWoGfgb0nrhTI/V1lexbD5rVh
7MDO9PJddqFN8TsOCmQkHuBDZSpW2IXgJ+2sVPMJp2uEZyttTnyOgTkyfECKui0WdkgIS7lCmvt4
ELEzNTFfZ73TKROuC+CAcv981Gh1YnXTr4Yq7Hl6dqz5P8wHCXC91IzfBAja74I6i5F5CL05VVyG
2FzPrups4HS7nyL/yt/T/zXtzCaIG4KUR8DbKTzClsdf8jUwfXaiOI3ySWyaT0AJf9tF9m6AuyVv
gxWV0l2zDDdrKj00j5a5shM4ZScG4xJcLcJax0mZ1NYemDSyrv2VZmAH96wkH1eDWqFyrLgbJzZ8
BC24jxc1rFL8XmoUfLa826a45SADDcEAGSEOhrM7kXKuq1Ln0LFDNPXejPn3KAsVVxqFCX08tyXv
u2R/sqo4ID9HfYnZVuylJKEsMtFAhyMhdWOhg91R+SIGk0N0mVq9zVsRGIaj2l/GHosJD16BM8CV
6SojJZ8Chohp6HqWfB53ixD3ZbAnDPQSnWMaMW3uPiXew+I4nPxYD6GzTZHvvYMVO2GL0PphUeBR
pnKTMiNFbjJv+ut3cKFpdDXKYoaTGIfK3OiMODEbX2OWebjLaheJxP/Z+/CKuWun2NfTAQOtZpWu
VITBmAxTdoVlfLpZsE6zCpCEEIuOVCcbOihLfAHN8uQpy0DueB7lyrEexzpA588GYIBX228VzrDA
zeUx5uyC1vcKCJvgYky3bblodFGRGTZnreYojE6hCrEPZlsne3Cx9Qy429Q3Jai9jm42jY32MoPw
/6r6OSnDyTw2C1Zv4or+xWxIVKPd6vAX+IqwLlOuGge+K1ZMnqXclDQFE3isoTDz4T3Yf+v9gv2z
TdpthgeaNSqxYuGEqSeSii9Ni5ab89RGEhGFwHBcnBImvEIVvbnrlKv+SIUTYa+zMV6tzXjXbtJd
frYOApEDtUhnZjkR6sWf4iWhBjqCUaArzR10ouwwa/AzvZGOzaG9r1BWIrhJh3Q9D0tUAvJlGDFV
DG/J3hXsMQ/C3espBx48PqIMBjAIESRJMbedKd6j40IeQmCL4jinCuy8HzWRIrdN4ezf7wIaLdhr
H5I895Jj68Z+Cv6nz8aXTbFLAw/WcVfigK4gy/7asSX14hcZPChOqFtCyW9SOYHcC8XzQoM24NxQ
uO6DrHfhyVo5YjBxXeu8W67HS8Zms4ubSIVQ20zQglDJz44O/MnB/890300A2EgC3n6q1RCiniQG
pHMN50gRaCgs/jyuAXuzbUQ0eSlHetv67A/LwuLFTObnLByat8yjdbUKIGTFBpfwqsX8KoeeHc2K
TME5FawsGDQiqAYKRoXFTy1yn35kKEyKF4VEdFux8fEn4WpLDv1v7Y0uyIQM/Xxn78I+rd3qxHMN
U/GikPmSjiIr97y4jo7j4wLdUptVzONQs5WDHV3uTXYHsuflx9w8z0++1CmygvXxFZM4kWudkrcc
drlYqdazS29bFNs1EODJ8xe3XN5ZiQeMcsg+JAv8kcJZE0MVo0daHdC+5BzK7D3dZon8ud18KBL/
q/wd1QZev/tY92wpasTZLdj71BPHmDrbBAZYrfmeZyenNuAyD0mHa7z/y4fGPtDEWPoHrztnzt38
qIxaLFMkSI6LF1Ec0rqAQ34R39gZBDySbcZUdaKLn0tCArH0zZnEvmqhD1k8KizkCyGS3sL49Yix
HSV5wFjZs/YGtZXqUqwYMKKKH0SkWSbDq2f9toyy9iTW9IVl8iAfO4QrBE+ds74WaExMrxUZktUj
JVOinoxaihvZURkdYiJ5+ouZA2HlbkrdWUpOGwGwXhmkiNgYMNCwEp/dISo6fUjbrXI6Rg9bSuJ0
4MbcS/2AG9IS6ZVvfBGDBcUjFpCiJhUzCwSxnS8l0PPZuNP3khHjZoTJZoF00Kj7O2KbE+FJ2vHB
EM/4kNfy/yWeACosHepCJaFDfBUlFCK3mkTvgYZ5Tk3w6M7kB3DjQ44pZZ3boQjEkqj06UgLHrAj
ecZVhl+nkvRSr0iZcs9tgut/JZw7UdBaRnr1dUrYtdZp2BqxIknfI/l+8pcTEFGHiD28lAQSWcoi
jj7uzZzyWjq117YWDRaJHKMnSA2d7MoYsfTc925bxqBj39u/+Erpx4QZCrd+u3o37CT8E6pgEZSM
CtV4AbWWsrDO7SXRFpmuJrzYMrTq2ia0SZGxrc2Rd4kw3sW2fCWyvUuSr+Uu+/wnRpQTKmtRcbBn
rSBSJwVxO40d/Czo567DPqR7x4Irbf2w0oTTHarIyMJAlYrQfq9sI4/aM7Mq0GPKEwvfz/lTdIK/
x55rwd4t4deO+0D9O96RutW2VTuESG2pf5P6w8pf8LcW+a38DCKbntmV0fcq2xiran/sCMuvjgz6
MBgGJSLbvjpKEzAZaGEyEhEs1krmMQ2y/WP1inR2Z9edwgz/hChU1IiHRgkgfrViEt2o0upGT5cE
IRqVZUKblMbFlDP5LAGL9LsqudsAJ1l+ObnwIbT1Ik8hhlItrQf6Mhus1ZkO54bJt32qiDw77iG2
LEcYlW27crHS1HodPHN41dAZ9A1XMgOIZzsCeXr8OQ3YJgj6vqJ/7nePHsqbujGLoUZoyP6yU90E
RASZnMFLQbM1PFAq2iQYdXZmX7XlrQjFI41LbytogmQKsTMWiRwF7nhZ9Jy997egWUOwqjNtv/K/
iKz/T9wTzBJ7CLk850tTVWbp1YSVv8cAdcY5uPEHufzh3WD86NDC6YrZVK4/rFTJCiTKhfVxDIUM
Y36rklgsxXU2I/MAqw/71b4TwRcAp8sZXaY3oVUyYUjYnytQ7FB4LfQzhIkZR38sMAcuvO8KVNjR
bETPr3JNvei4fSGQxXzxJwkOd9SFtDKt/YjlOneyixp3+srQfeenAzf74czFt7VTzZ4gACEFjAQW
8lJ6JMKVckmiXG72VnN41KJwFBDuOeBdT81eAL9nh4c4T2iiDvRLIobBsXbrSR+rP4uA4IxMN5tp
u2lH4xBIaf3jc/kQQlmNoT3o4tm2Hkp2w1pOZZ6lg7NmHNMZ5CM7sDd+X/YMV3r0keZ9qzAn6S/B
uSXlPAC31V3VFFujeKQuScwBooOwJcGoLhsIWgRqg6cvBDL5MXqrjh2zRg9/RO+f5x+mQ+VOu+WN
0BBJF2SB823sArS/K2m8UJpYqKSfAb45QoCnX6NUkFX7MaUzd1r7DBJ30E9pBs8G23CeJDGAoAcd
qQFzwIc2EvsFDpESFx3QXf41vuMA/8u/LrHzFpTu3WFC697Pwm7ti87LnNyyi+R4a3jyuWbFCQ2t
ccHNNpDuKyD2dAuy5CjVXZE+WJrJ2y7etWkd3GPUkoCckykJJ7/0AZfiMSvEMOvA7y3zSPCMoST2
4mQW6UnJmZf6W2tL7R1R1Xbz8sW3aKE4HHKVQp56/WFHF0K2MdFw5Ah+rPhay6Gg3W0Wy5F7lMB5
YsOzT7SfzKVaOVVIA89D/iYMqElwKlC/KDVzpY7lh5OkuiHNQEhIQlrgSaX4Hgj6KlPLCz7nOQXK
uI4OpopeOelhR+ShzaRvbAKdUZ2Xc7aekY4U9cNIdVll/5fHsIVvx64nbQwuMagdgJeCvC9+v37J
hQhGxrNASEEY3h1X+BSTwHvO1+sOw4xIUoJWspNaZttBHq4a0yX0G+SBNbgcHXepXY1yvFiDRXOn
1BDI+dJAWxUGagpuqqXwB6h2K7CDY3ibwZDG9zZZ8dzFn/Y0V770O+yk5wpXKBDeFq2rFzoAJa9m
ZB7c3stci4qTRVisEMSGh2OZ064ssuQ+/9QudUlgjSEkuZBO8SpbtAEPgL9H5J5BTsGGm5kVZK9S
e/cdxNLRUZh1E/cFqVu08+Mi0joSo9O5cNgGGRMFmt9fDfcR5neNNsBjaB244F/01eCh54LpQJY1
DFdfJU05iuhdbPD8E7M8/u2bcfjbfPclrRHplbhvRqroLZfoQnTy9l5QCb/h2GF5q5fhzGUZOe78
VfUcLmQ8qT1qRcnE7S8zFUgs7bxyQa2LiNT3fVxvxABR5L09mpzU9tLEe0+SL9+VGWy2uCDlK9ts
knLfGH+OKUOaUjkxBrQTlLPWy79ya/sjhQvR1h4HcFWkM+XzPeAJoLNHcNfi1NjbWwva8at1WSca
kLX7uMt/Rmy35iVqFRkS4GXxJ5OSSqekzwPqYkncYjXAlUPJxVmlUmWgoit87K4JxCJ7+PldAH8o
bj+mVvfmEhWabjlEsrxNtrQuFuzi3pDO5lW4N9EDaSiMqriP7mgmT2bXnakeZaJQ7O5RJgsUiv0F
LVBQTb6DneFRto8yjAaUmKOfXS5UXVjVZ2Dn2SIn2K++EcrecsLqybnbW7S6mwaZxz0l/VcffIjB
SQ7CIZje68o6fyLz+8FIJEtZF3VbiQ6DynjxnHzHiztVaEf8TLwyDfu31fcBjzKyL9ZUVGao2lnv
xlaAIIjbHHYtftBYWTo0MsA4z3AMe8evWf40dq2ztfeQmKF+3OBsYtwkl++UVQjqMdIG7gwKuFOJ
FDd8v+3oNq68yOAXEVsb+OjEZJKASSTz3kfS6SWRRfeqea5rzwkZgI+HfSKWs3V/tp7ernfn2hSR
Jk3ztnZG2B10QuwvMLmOm8w5X9TtiqJuO4qA4smkKba9nahDYyEYWMpbKj0YwTV8V08ZggIkoJzY
CMpSAPunABgSI6l6cDrjGUvgleL4E9kdXkgI/cVU6fZ4i4+h2ZCCy5kA1gJEtNC915vmNQIOA33E
b203CoD4Ww3MoUF1mrTXhNECmxf2F9tmdvBaWeLekY59o9AoNcEzM7dxdDlnmW4WFq+2ZzjjYMXz
W2PZWEdWd1gexuWV0fzzBgXpEVeR3Net7s1vUTV3tW9rZzNTg603o0/YGs/aGUvwvysDYBzsavF0
Cm0Gp6WsvjK6AVox5nvAtwuHyQDiRTVgGLKwp5Ttn3pLYGdeCLFmhEWsmw3LJSmnlN607FLQ8VJv
OQxZh6w28RdpyEc92MP/UrobbK2PbdgoSS6nZNthLAkd9AflSinGpEUiE1d9kHayCoTXVdHXSrDo
s83RShUjJNvYs3OfvzQMqg01CAbByiUf0ptmtTu7Wp+bMnBlVBbu3FvyTXf3Um8Wa7OunqXoSVYc
Kagt1v89pVUh7sdPUY+fsC1PyVqW/XvNbqTgBxiO3dSVHFLpXhezN5aaFA64XdJFl+ojpXc2vJKg
cSLkuB0aKnWsH9gFJW9EHItRL3IFG+WMGxJwZ+7G3KXzsBvEZuCS0c3znK9Tykxvtw5Du5LLuycp
k+nQBnkoysVOJuAtheo+kX3lPq3g7x2H1MStBSTiDxCWgrD9Op3WEr/TEDZTlNWh+trQArG9wxnr
MWT11lTqONU4vhmGsI/dEmoNSopwLdBrDnSWpPPVpF9dxwe1FgRIIIFsXALcrIHqLGfYA/q7Pqi0
m1IK38NCd/Qc+NBxzNr4jIySbxDImzZNtWcvtKrKuzoyhRJGnvF+zGAUDJcfiapBmwZjQLAuFG94
hflhiRkwryeuO7EHswQtXPCOMCY6wMARazwJovaD5jHSppOiadGgBMbm38ermt11X/2xGQyUUQjq
nFfXTPE2iTpBZLJQwmOzSpPpP+UNaZL66f8U1mlw2oZgZOClh9unTDJzpcI3+WGOwJ1hMHSCdukT
PXYyq/8uouomB478WCdyk8puMXrpaP9YfGvYB5RaZ5nd9C6+NIl7TgcgpyPHDzxN5ctXaAxMMsVZ
0C6pRD8ct4Xwu705lMweT80dKNjK9d/5Mj3SQ/Fo6RRxhl7YQ97cR2nwLQvEObD+Ne2tUAA3tof/
RXScDzAqdgsIKIfZxFYT3QQ1b5afZ9K9J96Gbpo6GvUJ80exKFahx5xmrKNxwY5VC/BNyG6R5ZmB
VJpyGPyCUYQeT92rd3E+AgDcX0kZsdm6cM9fzZ83nH9YEbBli7e/DcRkafHC0arQ8RnLHRn4xMjI
+U9eYDj2XX85bKvvN4vfwMevL8igW2N+e+oU6iHH43O0OfcGCEwqRNRplBl2mbtoU4sRjO9xqz5j
vCFxyJx+emajuDjQznfEkkJswbmxOzfTnPbmujHUqj0TYWv45hOnkMbwlGdebgyS+QkbWiZS7pJf
jg7BRBoaPZ7kNTLuGOx03jEb6hClCtlv340jNxBsCKKhKTAAojVcpmNsWPBw4UsbPpD0DYmfuHh/
p+pOwAd05ppsNuO3n3Q+gRecRm6mbGRFnpsHc6VbDLC6faxZpvuToIuBvPX/BLKoZw8b8AFKukmz
q5eFjamG+evFgQUwOQXarIpK6cZoTAqgUcvkZ28v0kX13hiXV9iCGt6dLv/5NLGmpcbrMMmD79ac
eTj6eLKyCwogz4SOLeqFF/Ij5piVEpejEq1vV27Dv9AUCxOfh8DF9G9tWRkK95GRFw0f/2PJgihe
ULZygsD2hDdrrZwiFs19hzqFL4cJSXqrPaU+/VlWU2kNlBHKmQBYZ+OEqCRRhYZsw7rIfxztXcY/
v2V2lFC51pBDYBLxBjYzTc6tX7ItE+2oDb420wctRlyNTVc6fdNixzEzJkIILr+jlOfRkk/JPs5B
qB4/V9BkKZknaEbaml/vC3Fx7pcMW0Bp+jhTPUebTJAIxUS80AhiMIIwzc35cjTxvx6R3rMxhjdC
4YolWrjhnMqT8ESSedYQquLArZ3yY2NMfWOA8CZYZSDT0nJ6fmHl/1PFs2zLSCuxG0ZAuFrSZrk5
4+kGoxlSSHgGCH2i2+7hk2WFNdAdnaQ71AkFRGIJZTTJWrnJxlHg8LkCLgtIQ+hl9ho3P9mFT/3V
IQBlQkIcWSd2BmrWeYdnSYeqcDUgWtxt4H6KKUdCFGTCbLCZWU2wUV3H2CRrGPQo4JvfpTOw8Rjv
ajgBoUE+UOJlgWm8uLplwFsjVtKDShKgW01kTGAMkdnGPPirmbdT+4fD56jXZh1QymiRKnFcxKY9
bEGapYnMGodPMativHM76XTx7EcaBgAdDrsV+n2yeqNcE56Hj4iZiWqZzXfd4EfVFm7+MVPhNHym
/an9qnCIQg/eZXqIlH7Hk7fAwZThtw+R1dblGtJvPc43WyOfHcyreng1S0c38D3BGRswDmSP7Fkz
CDDbt3smzD0+jgliOMTci9M0MsjPD9I1Y3hA/JC4GFZKUZiFlwoI8J8KyD+JMyfaj9Qwnot0W+Uy
b3PHkPjstJweUb6bMN4cAlrb2k+PJoSm4anqEyUZvpkTMTNpwhTAj1sw99F22+NIaUNmjCZynoNd
f7yNV9OgKZeS8tAZsoBGI+Vla4dNqws7ZS0un+Kd7Xg5Vfttabm4L030qwbAqU7lx3gPjDrVuLDS
b6J3Rzra+OYC9APNJ0aSwrfEGGryIhVUAZNGB3v47+S9Hm8o5Mezpc6L4GLq8VJlRZ6jLFfxC1oN
yMfu4K43Hd79QQe2Gh603s2fJzrpsc5kDqZAmw70LToeE2YnE0KmlGLG93cGLlIMkQmApzDPpUYH
4Jp8yhrKDX9xYcLVF4mBY4vaK5s4dO9UY7pTlxq5gdgbJH+S7xEwah588ioe+JPtfCClSEvERmg0
eoJ09njh2iRShV5zcJ7x2Jpg1sY+pFXzAQ8ysiTA98NqomEsUkZXOVsKdKP2ccL6vUfnCXXbgEBC
rGSoxOhzBVOPjcIURx1lRZYmgMgfKq+qG05zQfCo71DySTmqDJI023weUFnGFfzWWSQ2SGAGi0Hi
pTDelAtDKMfP97XYNsrIhJwGWQlyKU5NGM2RNH+x3oftZr+G8nUyz6QZLfKLhRBT299BtMA+Vdse
IETs70hmCKi+OGmqZ3TtM7H3IRcEwY4R4sQfztOdV7whsFj3b7jg3tHd56g+lHw467D87pU8zKw1
B8/E+WFzaAXtYRWbIqwfpEAopB8mSNUAe2T0nWn8VY9MHYBREro+kFxrfkXUelXQR6qzYzHIXyZm
pnZPqtILyiitukniFaiuflNBtbI6NNHs6KoC+mB49b18Io711k4FYEdu44+dZg3g3WxuWAkZSyD0
LiyxNurh1KnYQ2fJ0c9Tde6DBhWpJeZPprBdJgoKJexDAYItpthWbwcK8snXa34QfS1IDkYmBuMM
Cm7wt6a7N1e4kkvu2ezgS0PmgIa3QH9Jxcc0SK8y3RD+tmSohN+jQyiwjFaWvs2R59GifgeF21Vl
y0FmdIEpP3Sg5MVi2d7gi3bApDZcu2g9l9NceXTB2tKajGlir6LPpKenALwwaajSHeHcPRB2Np+/
U+xsKyenD8G0RSdVuB4r7XowpBLURfHcMsiLpvjjK3DZ28bC1BhXXD9EXBq8WPK9swd1ZcUK7JKp
4HGlBz5P0S07Dk7lomOLpiV8h/sUbCKTXfjmXPD2h1qFQJK2fPMnyMsULCQYEcJc7JeGjA2VAH3A
3J8G7wYCXtu+oq4fEHCavuCA6Do8uU4UvMgHgdg2k01RfgcKxdybv/7zeFYMjXZsr0kwEGApw98B
NCKmjOPtJoKuj8L838Hz3/3mAHgQ26bxEX/4eQ2lgsYDiIj6OGQc1I6Y1gBGyojYW1g9aVUvWl2/
uQoYgi2QCBIzWN1HkxSwQ1w/AK610WagJZYXdwFXZoR9r/l2ecjZI6EBT7qnwOp6LNjsZV0xr3IW
jTFoE5NcyeyNSaovV5+6caHB8bCHCO0w2VRSd2w9iErvbURUB4UDlm5j+IsHezVpY+9THlq3LDtc
0z5Cvo9xiP6KKity0j4v6WCnrkwH6gNC20Fr/6morcRtdRjnMPoZUZdM2Oe6/i5FOUKnHkRr/L+K
OGU/nwwnb2wkKEDJ0nlw4HWNdQ2Qlvis31OKw6XrIT4WuRD/CaCVG9k7/cXIF27sF1jS5ZPAeNv0
n3Bmfr70PIoXbswIFmufNBHbRSst9XjeuM4DWQR28kj40mqW1kIOWWBKDNc5lQxeyGbbzNh0K5J8
XlVhS1c34ia36rikt+cDiirhD9a9XWuuik2TPGxw1yhDYwe4VWXBlTdVGhXHMxwJWzkjxlqrrrPh
BclUj1gXcUUwVOWpihunFBUuVuMG0c4KqsOMXQ9JOWpqXs7aAQ5uLV7uHAyYWEsUMCnEQZe03O3r
qvwU6+mTI0Z6l/eiNzdOnJZ/xTm7HfTU5WOueNWXRUtrrOMxJlbZtKTff1ljMJb5zHFPyt3XqqI9
o4kR6fDUlDz3vukIYCDC8HtRg9Un7nXBP+MjJEx6C21PBSVIPtrSEH2qcj8aba3YMw8iuyAwUqnO
zPoeYupr60Z0EuC4+0JNX3pb53QoKyKmqHt3jdTGy45rb9N06P2eICcSztH4kZFdiBro91BsZqNX
QgO6uiMUWncc03rYWyg9hJIBHdNJvgAy1ap8GFtlDNnWpNxBMxgJyjl3jOeFZkhd/Hlr5C8HGyxV
sHgyP9vBHjnYzI6/pFH1ig+eUFnhGWp8P72tPL7sGstDfPlUJfBP2QSo08GSnlW2ivx26oWSkJsE
Xr/EbgmfQZ1P80V+SixzHY8e4wAqwD+Ba9bZuR9GFYrasBLM23XQzVN3nPMhjjRfag2fnBNSSdwT
0qnWYV+w4MawwL8Aa754umJXOEmjWsxgn8cHikq/lV4X691eCb4Sh0UoBCuiehDbh93fG9rYwQDx
wys5/2NVd3s7OQbS29gJi9LOrBMzW8TD/c/94NxjcMqOZ50PN/5WwP2lqDoMZp8BaYr6U/5Z3Pho
MONPxCTcTX4vigWhvffL/KR7rTuAATqAQ8dp4pJf6Ymu5wN8cyi2nHE4YQKOGb4HiuLrmsd/hsAh
5pNaXKex455yHurRprkCYS1v/pq2w7mnPSgJDu4gPAZhWZvSQtJDBDqg7QINKZ5rpHjHEaLZwauv
eLjOT6tbSnj7ZHGtuzRYn6p19jpjMG7634Lkp5dG2gOGsxlqyqZ6naeup4mmJG1liWzuYu9QZOcy
K8dNXgbIJFqRk/Oz6674BGT8FowNrDV+s6ajj3zxaKB8q4FzMxkjwDWOKM+4/mnZh50dofcIwHMt
mHBEHCsdM4GfMJEhK0wDMWpm+3ka6FO+uHhaEWwCC1Xz+wGpTEa3FviF8m22bsySSUqb5Fi+VjCW
k80j/JP0C6lQwN1UYsoC3sczF3Oiisxva22HsPs5GG0RkwhwQY1NT3WUuWUNuxyFIeTIQXG807ZY
lJd5o2hZrNfnTmoblQAW85GxRP0+jZun0LqjNk/FU4G0x9Lzqs+Ic4bMTlMQsjAdfYEJFC83bbup
J7WbIWjqNppPFKETKhCGbZSCrS+bEKdTO/lmDPhq1jc7GM3tJOvTa5n/5jo0SRnVbfOkvZhV17ol
1zAuPBvCQXl2VUSJaB6xx2GmITQnA9BVByH4yjnXwgsO2LrbfXatFHYFUsQbZoJBBbiqW/vOuN6U
SEGfrAHvJUlRKUMCKwFzp9g4jtaWwQ1uNhiaD7EirsTL/3Diusg6ctL7IqHG+ixI2Ovbks4RmCxx
1yv7cX+uiXx+yhWgyc3J9oCrt4rtHfAIkhT9aeNFXPustohj0Rwdo7CqM14+hCHH4kVIdLDC1FIo
4ue/cqrTiTCY3DGm1mQGpxgoDzKQtZWNSmWGn3wnDqVaPjcq8e1q021rq81YRmv1KP/gPf+K77w3
7AGveQP9PrZEa8Y+PkTTbdMqATeYD8SpXzTKIRgF3FMUA7jJZpAIVoPHSWOSbC6bcJx7Ot9aDwcn
WgVeu3EASOwBKaP74+0bousKuhHXe5pDVUejqIsBjvgyXOcWSLrlVzvEM2lQJcXkTlEaPI74txc7
tuS2coTbSLAHvE2SQ58pxGU/KHtlmiqaEDPozQx3rPivxjtRcqdJN2IoJeXuuMI6ZmROYgG58Ohx
1Kd0vMjDHRlz4qNviLB8SOffKrZs6u5BFFPmVDBXsRQNRhq2nge7/N2HzJkm9bKNN5DhRRqweJVz
yQ0Cqg6creGCK98TmK6QrLVagy80tcdiphF6vN+/vnJUf98bbbkAlOwcm0rdYValpqD0geFRBl57
l6ldMWKSDcHg9ZRQic2QG+MMcexpY30nttUTBBgm5eOHhL1jd53uYGNBqOJgMAiI9Ylc2++UG/oS
1q4CHovxVXWcKoubvP/0RNBRn650Ilz8Aa374leAaNb9c7TqARq+RGC08IE8ncSjAIi1IBKczNl8
8u6VrYjl2Up7yxVW8Pop0F7aiv5r56K6vZuZvz6xakN0CWbso1ddK2waIXh5xXGXVuM1Q5iuf/ci
MUPIO8lkQYurtdrHtVd+d8v1b+WyLB3UgUQuhu3RDYMYP6M32eqFf1c0IZjpdGrsbIJlwqH4LvlG
/hZicc9n9fuOO1vjXJJ0+pRTHly+ysgrJauBlcu5o3M9dXYv1XFcdaj5MtuwFPedb4WZKY1Gf4XQ
Xut1EqP6KNGktXItsz6wJ/QmgMzT937x2Rk0+IlmB13wS2HKtUBZ+hpuVI8WEzBjfVRjO3LMIx7f
cOPFUaUmOaHcVGBRdR/4GjihQ6fr1DMi5DJbp34M4HPpTLZJ8csKshGVDmZmgut2moHOgAp4Jkfo
OYlV3I/6v5Vy4UtBHMb9r89U2/BG+o8YzFTISZljKsq4Lgg5OUjK+cLXAc6Hjm4QD9O3KtKZp/iE
DHiklZOvwCkaDU04Y7gw0ugj8Y9gCReF76iRPKwok4oXDO/+3dM1dk83bdr3JE32ubmcnu/6w3xg
mKbvfOVnbKEsieozNekTlBOf/IY5czt8E0GoY7XdFvLUtcVyNKx/fq7hk8b20hbHUeHjFjDS9zZL
89X/psQtqsBsK0pNVa3qTm5VEvVk4MscG7CNgyg37qYBy2cI3/UPRtLohTjwDp7IZsfZiJfW7n91
c02pO4nLH+K/9gJTQs9WLdVU8rZwUWRPi01lOJqq3oTsTyY4cg0hEs9qqQ/Nxkn7VZ3sZ8i8iGmD
XozKDz07I2nEK5tMeI4kUJWGm5jd7hEhsBOsB7PXNdZdE2LwTgMctKvrksDbQAPyj+g1bEVaA8Y6
jCXg8TLmFTeTfhz7MOsWaFlipSECl+4Ek+rrtL1mdd5eZ9vlLWNVk9Hk7EvzC7esI6JO2dTy/p+1
0sZoJrL6G6KnMkPlN6MT0xBsis7qPLRin3e2NBgXJsyHQZelAkK3DD8sRy/cZV1vH4q0Kc8qmJe6
0lvP8udiZwARP7crkeVWVQD8Jq2xD0iUepv2ghb3uBr0rYMO9M81lH1pW4aK40rRNIAmiAbggwfW
G/JsMPHBYnSt0Fs3lEah1nilaIFvQUA0q26rncjRe17f5jY2w1ebqVqwLZkhYZta4/Vtv1qG3cUm
3JI+szzMFYOByexHARp5kth7XMkHLvpZGKfo0HI6mYHCtJMHdEIbb/o9R9kCLVeTCNXdZxSdc6xF
nYpAT7EWkT4qW2wZk5H9wattqdjcz7qqcURLigbH5yWXyAxDiS626I0XWuysduWQYQU3VRdTGEwD
M50lI9XA2E90/Da7PfhkTgXriYuFUsdci9Q4mgRLa+NR8j4AW9bgkx2zuyVlvYBch5GpdeaQTGdh
yj7Mroa9JV6/nK3wCf1s9sXd8YLPfd3nBuRWGsTS6nTb8gKRMl0wC477InOwu1wdywpWCUb9yV3h
279BULI7jOGMtaYQazQrmmfjN5I+8JgWqVz83KBBK36U2hI22855XbEODGO8x/sNtZPYK23N89kI
bB8Qu1Nv9UyLnilaZyYtrSjfCSsC+E0VxhY4yPfgWRQYhyZlOKmB4Y/gGe3tfqt/itc1gY47jJo8
KMpL9wsrfVGDXtjsNP66QaC+ejfQ4rqpbUjFlo1Gl3nmvca8DpYsVhcbk8df4e2t1VKBZKzYBnpL
tMb+nE4DGmc1VoNpqZNQma8an1JxaIjwkvw+lTeGYeSlMDoY118nBJllezFkmqznvIrCwoH7Ov/i
gmZhu3HfS5FGHg2xxHZwLUAEnnvL8brhE9crO+U2O9w10Q1Fb45hj9QzMUW3QCBQSwpAROw8kLEk
nbMSuGyLhzybWRwumwgl3IUmDRjlEj6mT7hfBmr4FRjP65cuZvDgkHJDSt1x4gSLr/fLCqE2vRhx
ReE29tLltfF7UkLIaoPA2hK4HgaoDnc9tBAKQxv3nHPjUVSJqEC8BfT/ofQxUZ+iVGSeksZDwQgG
bhGiuhHch24a4e3ZqeDtCByM2/61i8x4rZEr3FHOdImhaM8odmGc3FdJBsYZYyk2UoMHwHeMRKHl
PR6CDRUTv5gr7Z2hWHWFtT8vPLO06PcIDURUSg8VoPOHlGrSCh2kgSZpT6tW4aXLtzShwlKjRJWi
fKrFZGN8ZsQC/kmlfYHIhgHVx+p5fG9AVpw9Xqlw3pK6v1mCv5u5fFcDvVrxC/56YRpE8ExZt/NV
6qgBNfaxOq9RJy0VHejvXTqHnFNyQL/FpbDMS7vBQEx15Qe41yR+cFQbaLn8XRy6yy9jNZisn8Or
lfN+s6Srk1snJbLOQJwqowhfVDR7vII5hMHE0JF84Wbraz36yVKm9BR5VJySuYOZWcJeYw51paPZ
OSoVhvNU2HZArRxkmMx9BsR0vPLtAdhmWiwRsap+bW98c+S3VamRIA5ruQf45dYLnpWHBKAd+TcD
4u4GmriZVEeeKexqSIBrIxKvnaDwX7VGONUANUvNsXcfiT3LWCkCDKYWhUCwC9ChrC5XPrhMnz73
GjBr6Z7DC8eifxqYexBF52OKqaDspXH56/XNOC1+CeI9QV1SAX+1HgTkdCBAc2mk9fZNn1oFMG0c
/xrgov3DOPWenG2A0uqxyJ5lfRMC79TGSXMdpryr6BW3mQszPWGAH65M8QG0CCy2zFztUHG+0uHX
hwDe+VAPfR/HJ5TzuQnZGbS/wLek9pqr+fAEH6cFPcFklOx19JlSHIgOSMI9PN/K0OizvmNqCvd7
F+p8Vtbz2wLSQJcXGBUPVHN5FouM2QlXDbjC9e++veIIHj7ajf6WMvZKRjRjOdzxSiqHXVz260r4
+TXT7Sp915eNdlYS1PfguAMXPKSrNPkPSzs+MQAeWxbd3T/WvQPUruMJIR/elbEAAMjzD2S0IEw8
LsdTu5IO1nwsY2Wy2kfAhUnOWIDqGq2e9TEGneKN8pAoFWzS3sfIC+R/H9HRPCWxVD6NkjO1RHXD
d0KiIwKj835rkh8OE0FYfzIbY1nzpLep0grhEDQZFzw4yXqMtvw7SA9WlF/QSk56voCukOC7hy7z
qf1cEpN7yvwPcuNiSkL6mmHrijWpSixvNggBqVxomUA/ZKBpVnQv43JY3a7jxKaw0ffdILXvSyhv
lk2oyF7pxwKOix3oZDc53oODMdzrvWu5rq5GdH0u+yBYEgT9941kIt30PueKMxcpPjp3/GAFJ+Cz
P4wUIQObfblt7whQZ6O7PRe74nENtAgQrqUVStDAbtNEmXkaMEard+LQ9N76xMa53gWetbRU56ov
5CjHrHMNNftJQZuQVAAjGN5ONzSdnSZz6ousrCP8Cg0/+M0WTv216EHlpe1obBKFIpXdQdqz1y2f
1pC2qYhbFAWkdmom++KY+r9hK7nBYg43do5BvQW0cAEC2ryqno8FUrxO7UeTNukavf2dwZIChf9Y
F9LEXp5dIP8DcW4UrbE8RmNZxtMxilABbG2fULtbwqhaR16YAD/ar8RCptdUlVKGSTFMd4L1bqmZ
NnT3YfLqEjIzjMrt0xgfAD15XGpaR0hRPKeoHj9pNyZOOVb1CLKoyjVOhB6yfiqnRGBrN4PW1IX2
S0QvCUFufqi3S24o4lg41LLEXhrB4OO6LvD7GI4oYulC/XeXnKZh5FAfeM0V8KXlky/kbIV9RXNJ
4R6rE0VIN6OZd/k93CMpFXHhcpGHaiXC+i15O4fzMZKanECEbSwQ8XT8v00aAIr+CPCsNJ+Hdta8
xi5h0WogvBkXAUy8S6yJNQt0AOz1K7QdnFCn7CMKxi2Cvoqs3Yjn7gvFtn8xidlkRRQhlOTFuZfR
cv763n9VqDOrZSnC8F9R2S0vStORH89HItVfYdRWicghAWwpJXw7M7nR8rC8fAVbXdGlCT2j09OR
MMrB/EUng7odZnxEjzEh7SEhot+BgNF7XaqgwB6S63+U6dWT3t17G0a31Wx1uCh/xwyhrpYIllbF
IfBFx6WiJwWDZV1qEN6CCR4dXoqFVKsxT3ka0HiXGONSle+INzkjjFpZQ4NeyG1YfCo+jmmLDyEi
rlROa0kx/ctYtx269yr8HjBL4jmbWMFdRrRrhqlGNmW9zLAShKCkaFy4JWog+OFXAou8vRj0nim4
YEFcU+y8gR3KPDoENK5If350wxhBi3RUzMwM0Gn1KJEgokLRJK3krBIA1addfJQTVO9PSNwVdefj
SRw8aPmSMqWeI1LJBuSL0dAQlRVSBpMPerbYPXVOgXakdrY82YJIWAw6sHerwjm3ZvgxHCqmt2Uj
Wi/8bh8KyzrDPISXC9tNulUYeDb+SDDLCMAliMfVzDH44zRPRepWgaW0TmL8aUNhGsqreAwNePQt
4JbrClZ4iIExQatHT9ZM0iIoVtjMizd2FVZS/E7ZzKNYkewKQD5mulCk+QizOXNShBXkagvB2uT9
u1QtFgcf1DVzyvAhWWW1r56OTvpUhBgdCTXSSSOIweHcglYvJ+WvArOlQrMxd959hlnVKONQ7V0L
1uXZ/orbB3H8ZLbfS8IXzdNRhFn+DcMdjd2w/gGua433ZghHD0ZLhHN+gwaaEC613djnRwIheMY1
4+EGxN4miKlJJwZms+LQ8m4n6US9lf7Pn9K1myU3YFNgVoaCiXEL9s7ppmXJEtbAJHU4j8G2XSXf
UTF5X6qRkIKgbLk0bmfri/CrCtujS7dVYTd8x/4TJzsa/m4c23z/lYjIc9ZgkUNpB4Mp1CrgpZOZ
lIjaQBIMAtouT8eRboPJbDW7/5BHKaxbS4P8s+d+aLKOywf6cggrqH+MA80OeR65IC2RX5clj0np
uRHtvIZgSVwvZvfsp+x5DtAs6axWRhlQ2LYtO0civwKVjG3KprAVcngcgBNu4hWa0e4k64ssVYSk
tOkQ1h6YF6Ocn50MbZATwmA/XgqSPJ851GUEOP2DmEJ20TlAMs288m/4MNax654M7PFQ1Sx127QL
hzaOpaPa0VB/NuWh2Sg763z4/VOIorw5vLsfgEjGhYv7Qfmb8rv7h4ZNMtcw87DSWA7rLQSWsif+
57KMzniv6wh16iwvEIC0kWkizgeEHxhMa7hEERtBYMvW3s/7ab0tcRK+IrAQBhwgdErvP5+TGn1D
kewdftfBh2HjMEXMmLLoPm3C7x2bMiR+W4heILiXNyLI086AEKIMoeJtt/hSCVWtnyBwif7hEe9m
e2A3K/MrVe4X0j6uczRTPt3zNCcqRIjZPtkJc/Kl0758xmFbO6lXhBG8NpEv2I6Gdlht+YZ+/qYZ
oYGLUF0IBK/crdz8ezoKNtBio58vusBMX6b/uIkgzp380XRrLU9nslWVtLtcNXxFqClHuEhiVyRJ
tTzGBkxb3CktwbFUqJKGex+il4yfNcgdBc//NnoHFM1UkW8HTF+B/bUDkZVL+EkuWIFScYofB6Nc
5IpJDaQgGo59Tws/BtU6RuoSEBDyEUTtVWStNNQD7Y8vX2PCgeLP8nOZGoZE6Bhotgq/VQp4L1IQ
dpC/X5rRZ2G3VEpGi6AtAOUXFtiEIG0C8F+3J/MjleQdTsb5UTkOdSdQwBanBNBiBhgcfd5Oug04
bfuL08RwNDCxiWvThIhJ2AuNH6MHOZlPiCadpQAun4q2XEvL/xdMgNP8eN2sm9XZoa4cQI1bCAmn
KGJtpXDdESNhIhsbgAGXq6JOLODrrRZ4ToyyVZ2ShcatylqlxwrXTapP87WDXlVzjNat+7YREZs9
QWeF/7Y7hF8ENjaHnXW0OsTbIYvn5fz5GY4fWay3nZv5T0BUc2MwuoK/cKcPI3HnOIThxxT6g+aD
rIbFF95YLMO4TsiheGO+6vY1rg1ykv9TyGGDMKPG3pbJu1CXV3mC1lMPr+4zBEMCUU255B6RqiES
o9GmynB++Xpe/ecRAuDA8EbkuPFRvxJ/Wo2o5bgCXPYBOISdxewVTh4sSv00yZHPu+4UO5ipafMb
mLFVAyZPr5+zjICu5wdMrhBdSrYiHiU1S0P701iP1olITFy+DZWvTAQj7jjtiD40B5/gM5zH/tQH
oVLDDcH0fgWqAEG35aksWhpZL3w4h7mHjMLz3ElVdRtmHZqMMRZZ4g5X8thnK4REoGf1e/1knB2j
An16cNNQS/dGU8UI1/26Achpg/WY1Cmm4uWExpcmC7ikb5yLvQdNwXPxhhaaeIq6J5e4ODk8gZ20
2aM6Gfef5gtg2M09SLZPU55Fu117pU65oprfnPkz2L6qhsZ+zWiAgxnamtKEVPdJ+yFVxmWCcnCR
IOuBk1fPMz02EWwI+bqLKBPPy5t9jvF0NBqNoeEh6pGxGN+IEd5ik7QWEYdCPyk5JWE9KYhIBTFp
BRANYZD2EZ1en6NxFHfqpi52Civ1X/0Lo+delQTjSIqSIKPhrYcH/2cytzfEcWJbYpArFAVv27Ch
EOcUYfWeZ8tln+c5fVEQ1J/TfKyRj5dGJCJrN4Kb6vQ2OA9OvVzQe0SwCyNXQg6KPXck960tEB7Y
sRuWNgOwJWWpT6MISsUqDyWAS0Wpf0a+yW5q4q4ASDGokYx6Y68df+WETLeoY7QVYyCuluZeXj0a
V9I0BtD1t7lyg0yy1eUBMojz/eBp69M1heoY9YOXr4kdRyDgq5pUcNAjmB9slHm6pjYQ3BwTMyJa
kuQ+1JeOPj7rvTqEl/Rtc3ML9vhd6DB+LYILr2+hHDlHhk1KRkFrCLIQwO4UPYj5xSIan3OFZt5/
FYXuk3/5cA5XIlyjqpmHL/iUmyg2Rc0wMRPVDgaR99uV3IAipTeDKj61g75lXIrWSf2juk6aY4s+
4fHD8nRX6efAviW2TdLaNnTi9Tt9eJtzASUzRfMg6gJKjtvU/atnppKwwOQYSUyyfxCK6RD8T8sS
UUl7//JjIJDTXGQoVDN1Z3MwjzFvz3UmWaEVB/0XHIxWsHhhLnkP8aPyIyMYXTm1+BWizJOGz61n
tUFmdMJ7nHRLXgdzLPjigruNn5WcLmTTVaE5fx9QhaGxz19DS8akmxo1YQXXsTAYT8VGPSVfsZYb
+bxqdk0hXYQw/oAg7vWe3QUV4wg7k++/k51FMX2RXIHwhfI82UAUGcKhHYv+uVOH37nJeGchqAPp
gb92yB1IxQ1+ben+cZQrFySuoay1DqSrVh1aQAg04vz2NVyyJO1RtFdZQbL9Lu3moRbk/cqjHgWB
/fNAMUq9xpDQo6FqRTbTpzu+rmtVYr5ipgPt9+mtzZWbSSWL9WRzD++sARSnuLjWqD2qHJU1LMGk
I5SlZIh6iSgbMo9WVOS+XWx+2XBmDGd2gNEMChfEocDGoRixwCsoB9nWrAAnpysIGOkY5vG+U39a
xY6+bl0FWtM6ikR7SbZFa6Ia6thT5eGzYvAA4nfbh5J1Eq6f02rEa7XlSAp5Hjk/3yzsZ3KEXIda
dcdPuqjxYYSYQsXXn1t+P2rCGev37JnGWLUOJ0F4SqlCzc1Ot1E69YIOM+QfyBmeZrAZEYdSNEy0
dqiFmeOBYD/0Opg4BDDuI9O/zTG+u2xmzLUpaQlUEJhUIkFIJFuNzt0tSvZQNkp0Di47LOqTVaJ3
+Dq6lQpxfmU3Y0XZvumI4Y3eazyK0PJ7ed4EgiWAstbl05D11If5zMvK+TeOupFuTaMql0L2P/55
IJMQQfjgeJNcb3q9rxg9wzeXFjTIapQJ7ZRl1iXQaxlyuT6boHYpivRDw4ZmiuVldbHq8AmFiIlL
ChniBS45q1Et4HoIQPc42UzLAcebKKRA85PgNlo1QOspIw9pbmUsEFF8dOAz09erMWa6/Drm9Sp1
Oka491d4vC2UcAXI+IXgIc5wKwcSClk5ISynVTNYBjgC/6kni+cII8aXROWzpAWsL5ypnQCV3JC4
Gi00mpkzny2J+8Tu2qtXkR499Ka5RcDQ/KzEUgUVU/INWvjsAbCbFYYraId8S4Fy3vuIigw02KYg
bD3hW1O4Qz4b7A3BUa26YKm+I1wzDdqObJsJZyWCvyEC9GhnA8YcdkvHYOrqxakQfRVnuTmLO6WG
8fzuHJ/MH8WOAWvoUtZa1naS5cKyhy5nx8ztKwSDElU+q40fCLbs8A2gh26hhPCU/9biLfUrNYSq
1YIjOfa4okF2veQbaZVD/s3iT91T2AGyGMnWN0xIjVfdEIJdDT8wTM3lIXCfG+zmXzq7lZOWBQdS
kge8Qn0IGd3AZX3o1ltNXV7y2sLuGeeG8JrT5+8/v70GchsDaMRN/Sow2x9RKKc/jS38CB/9HYox
ATnz539dhdB/K2AdnLaxYAgmN/zppFQl2VJUqjG36jUU5Ph1Y4w80oYai+0qh7+nhOSK4Q6JfKk0
QXKgMxakhOBatR0kLFOFOYq9z/HWoKkL20WI2jiwX13cQw8ChKX8Zo28UqNzgjxkHTgbpeYKdYsY
6T5YCtJLAzOzepNjqXk7lEQ1OsT4+NEx0lNaPjfgYOahcX0LhxwYF6JXbDFtR42MAMtLrRqp+iYG
sB5AkN/wLp5xsx7IMXbITayGXOHSVEciOwX9xmj2xCa34LYdFzbVNB03RRFveivSw6mbGQ12wW6X
b2NQiS4C08Mi9nEp39S0jqWO9NwyuuNKPmq6l4mUifxR6uLFcW2/vt1+fQ+1W6GCAj2tlbr9+6gM
l0OfgMNbbpNi4SS5ZTywXGHn6d1Q7993RbVSM9JiSUTvfqy4A6K9WzKHkqKsQbMmDUJxUK/uaWSo
Fk3ODLnugVs4M0Rrl7iWCz8RRdGbCO+fH5JcUrnKHuGVoLsZ2gVujcn0EZufSPhj1c2CGXs3ooYi
uGdpfF79vzcVDNRj5osolys7DK4Efx1Vwmqg9OAL4ouHHTHNLJtMCM/Epd7h8sv9l7u95YCVHdLr
z6q69RjRIG1e0G839nLMiKTVy2Xf8HZaHNsF/6PlmsLyKWUP62ZkaluNEu4t5igpHzCIBt3FOU0x
2CED2AdHZyiri+ZR48EFsiMWlU9HoxWB3TFd8bVoD3Mbc/xn36WuwzyuUg1bO7TI4KD03uvT7n6o
2RmdFw0HtR63qxeEW4NB7jGyOzu6D7n9elr3ueZEtgNM1RzlXO9BOjpcApmlrwKrKoNMwfnZUscj
0omJXirqaVxIoynNy4hdexGXkrGXD100Ks5TpbEMk+jDQQRMYl6zyqO57x1emx3QkwX4gslzB+/f
uT3WSlqLzHA/CGNQll9F1+/eyGzyP+GqUNtFwJOlSvPDn3LWgUBHN0ofqrDOVtcXJ+i+89tOrex7
Yb6Jzb4mrvtjzAr2kueM/aM+s9W9SQXHo/iKpIsQoO9vIVhI8VU3Iy1SGXMnyMdUZqL00SIT/I2E
litwMZWZj71MH1xVQlwwrgo/oryFTtOdBXgQlmOMllEI9dgRNtRAgHX9eYMAUfytJ4TR1ckpI8j1
r1dYMwInf4i1k3N6aXrzKA+rgj1VPAHxbo5/J5fUAVPnp0dd8tZt3Vq69AcH3uOhEDekjIS0PFH1
GaebrgGMplyN7xZMcRw8uWy0C7bd7jtM4bNl3Np6F4bWFQ7FMed694IfBEWGD/teRfnHFx2YyyqE
aTXstXGlEJDmKcmq4cB0yjjgOWsrL/hOkKM7Phj/ykzXQ5pzCsH49+dPgX6BxbL6VPQ9+HBG1m2o
QJA2hvdUmKabCLsAirjaFIrGuNMeNpuqqdZp+IiNkLHI3OOX4aELAGX9wyJ5TulmC40hBpU07Bn0
0l3P7KkzfOBIOZrfImteQkt/aoBnlA5cdT/ASfzGIQYCTW9xxFv7BFduyae+oyimyuBecpqGdFy1
wVqp28QOezsw6i36aCA42+87mwwtxGkuDbKB3xX8LF2D16jGHgVWQ5KWZMhRmEQPnGjxFuucmlLC
IDPMzT7kJUsoVhhIMX06VmvUoqB/c0sBGWFUJ+srBA9UVuGm/xbM9Yjy3EgKaNvE1SySTjm+h1L0
GEd03SL7vLaPcWYUWEHQ6LImvsSsK2IxPjhbAXk8/0XNTaWXNd1OOGLEoyASE4xvGxB46VRAC7Qe
4CCGs+jCluOMGA30xdAlWo7XHJQudzT6zHyMK2274MJ0r34PzvHskvf5Q4xes0nrVb324KDzj6s1
V83eSUKTnZVNmtUdEGhayBcPGnhK/malXCAET0ONdjt1yV7BxbH7xF0FpzYY9gNoYhWgRRRO+hPM
BkBnURizvG/Z+HTza32AM83j+foTM3nQFF6Gp5InFlfBvU+k7Ad/F08z5ehOTKLf88c5vrMwg8xd
4eeAUBFM9e9SKEeIv37TxMgHn5EgkokmHZD+Qq52m8Ks1505eIVyRwW/VYoNWAX50vorF6WFrpUj
2bcXloSlFrmQJeKvzkQiIUIOLOCPMk1qwFVAwnLXAOyTsejvatIJil7+8ZG3xqgpj0GZhcO/R82O
n1w8c/yTfzyq94sv/tuhe3i+CvHEYzPjK+klg6B6uKgIqBiNkCwdCjG6cP49I3ooRTDw5x9tzZ7H
sPVWO3OQNqP6Lm8jXzoGS4DN4Ns4Mnv83X0qaX8ybzrVFPMK4psZwNgmDxUSxJvkT5BnkVYOLqey
60sf4oFvxY5bi3NiIVw8ec6FkH3fwkuzG+UmpdhcBHmJB/uuZrksvbzb7vXsghB9Ml9KqXdfgSXw
cS9t0dkHx0O/Q3fj2NMc+W99vMIykdxRVG576kEzwhdhhG4f1EVNH+eOEAFjdxEm2DhsdusCCUGq
BNm4lJpii/mrv4MIXHKXpe+Kql44vy6l6ea4zGtqD/UtRtVHxF1vsTA+Gc+r+1MWquEKVfr6sWh0
HlUpseSPb4E0IzaYJ6Z7jeQXW+QP/i6XpARrQsQjSlLxR0ET9aTcTTOu78W1Yo4GPSWvdiILbpXX
P3doSANHenaPEQQbPQnG946IFC6aXyxAIH0aKMXSG9CVXiszshbe56rnPtX/380NvNMQQHpSKqs0
OozN8HwaVHit6V2xlXEcuGxqMTPGUOtfI670LViikRrPoo2ZpSuPYOXxhfMY5SYP6QSeJ7WBvMhw
i8TVjb4Awr3PlT8Gg/SjQNYmwScFoLFDwQGk8bdEA/VKpsU8IHDmxMEqvaYtAL9WR7LKdVUVr7kg
bbFQj7onHwQh87PhE7mP9EJhCle9G6mNWGLZmbnjKOIWvKaSe+jMFZ3MFONPB91CgS7gYZwAUarB
aRFDq2Bb6jIclO20Bi3SBJVw/dytzYORdEVTOfGQhuSxdcBROQ/HVPw+62qBphFX4ASAQJE8p1CZ
MS6lWzu2X8DFxOCK8ot6wDvT9mlvhxHprdrcP8FLBt6z/jTtIgZgCkB82NmxtUsaioOpjWp9na4s
SsSbe1kBp2jjyp5uYosFkope+FZq4n+zoSdFJ4izLRFM72svkYDRsCE1QAYaxwyTGXfOSce746OB
O/EFuipJBfp5egQoERZanWu08VMWsdubjcBRbywqJYPy22deWxhvMUCKk56+Qz9hTNRIEJRrc8W8
4w+q81NVaDb/NSyf30UQUUjOG3sbHeMYDI+krcccLJPfhIEIJRNGLIoDeHgsctezXuneKCrc/DSA
3ohLDJRyn7L1xc5Y/vjBe8yxxpYoCDSEO+LxwJd8iTVVJUTejgYuoTyTIH/PdJ6Aclu896FnhtYn
rQ/CAlAwBLeIL/uHC8JJXRwrGrZ70glrp8NfajTJC7mI2bah0TuU9LwMHmY75gdgC2YjUpyB9KNF
QGDDSS6FQatCBeE/pUouA0Tqo6t+zOnqGBcuw0ncG9WMDmaZR/3r3dvUByQKPC3lJDcd5KLliFJK
UThZG7TirjJQBV9GgDVEAiIS6z/3xe1KjLqx3WZlw6ES2e4SEAlMWyPxzMMeMMnfYems74HS65tU
hroeX1YjmsIVAkoefvvLs8qZias0tQBUYFY50ZyeNqwj8ACMEaLB9qJAxz1S4hva/16enF0ctAoI
EbNVlzsVVrpBKaER/Jj7IqnRugtYBzkCTMBhzjJeiKm76C5JVoOKB9bxndsdOd7lPgbCcTzhhPUm
BPWAYKrldeBOn6HOhlycvnFdD4Y555r30V6R55rD3jw7uO9kIyny9lvOKmNuEIQjOJJVmTuWRQ32
WvMfEGcwMVyCqU0ynykaMYCsabqGJwgmivIcx6SHS1bj0Os3WzKkpaWze5FjdeQhv1dK9n0yjPMi
b08zDNGRWVA3hLvVDRXVnP9SIYZYxHB4H7hEmHOqwt1JQxrUGxPVubGYGRi2VxJ/sJyKhH195EyA
X2CPo8WpXB90Jt4PfZyWsoETaawgo5/vdfNtxLwyUGmSVseEL2JVxmo2hWLmvHk+5zFCjXyFKj+9
kDPUFT9MYuEGojuZZSM+qEnjhDnMPeYDmJcgeBY8MvwymickFIg1uybCjjSYfVyCAM5BxBTJNh58
RwY89HDU/yXzYm9TvCsdpGwWC7Jr5zMxXPsumA+SCQutxMHkP+9WchYOvj5X+z7PTXw4zcqS8iAr
cmWkH35a3G9amoanvudKQQLSSzzSPwShIliTwq6S3pJW5DykH7Cyc9/IALEyZ+NPUp/6Qs8kpMZ6
2LLprfJLzPVI2BAJON4tTUJK5zmi0N7FqJ2qjkf9b9oT3ocmfMQI3onOCHGyxe0FfQMRsEcs8Y/P
2YxJJfmx5yx3kj3UdT/SRTJ0oCani3f4hAXlcd6rky3NyFRxNKVcDXUHsnag0rKeJPBUIM1SDgGO
W84FBOfXpZF1Vf5d2o7TZ1l5Bldku+aZsTUi2reSU+75Z7h92Wa4dHg6Mn5QG0fzsKDuZxy0aeE9
Kbx+Ol3aFtkRkBlkgdMfG12Yk2wuCtq4pm8fzcKaBWLak/wZzsgrkX6BdZD+PBe1e56EZNVb8hhn
OynYpoRegV2A3q/Nd0h2eu8/ToGalM+3G1v90JHFK0USst7gaBVcvGXbHINOncRzhVVQaZPjvOo6
5w1SeM0ZQ6pZRfXyxVfAaCui7TapiHAug564UyCX13NxRGoIfSH6LNuDmAr7nXp9GJJ8R+iZZW8o
eXnanCeccUbKe9HXh8A8wbBQYxnOJV10NsDtsika/csKVBnr+MLb8n17Xl0+QV1st+BU68bgDtpe
pErp2vmMC/z9p7mupRHQtFB2f2ZsUebrF3p6SsCJCwjZq+ohOfBnt4Uoi/wDz1lrbBCb+8P7955B
Gi1Vje/WoFl03XbteNXyNDcEOe39K/qunaLy0wozuiiUIfcFwL3rAfYX7pnbAj4cNR4NEYleILuh
WVLt3dQZtX3uSTqZ0BiEovksz2c5XXJ3930x5xN+Anfylcu5BbE9L1mYsPQ3AhPcdhlGWRXPzJvB
Q6qcU1iymuPzLkpamkGEf7tey0cINGO30IgyzBvdUAmu9LJdRq/ad6AzjqJ5JrQuset7pjcjHk1N
33aesH4dgKZzNzm8rd3eCshLLKOkpRGhUu0vW3FPAVUEvj7ZYimKF58uYpVY6V37jTlSa/IDGYEJ
LbaLs+Swp6JXE8HmvoK9pHOOkYyjNBDt9Ke9D3cBQYoM+KV/UjYGW5FUiiRShnvDt1aiF2xzMQO7
9YiwSMiBt2XxJdEQ9BELD8kwfiH7nO1VveEeNUsuaRWfEakqZ43hFP/2Zngf3hpQMeaXAbRtFxo6
5OuNidFGK5E9YtaUcPrTnYTUVE8T7BzfG80dCVhKu3L6T4X+f+OO5b7O/vbdKxxaPk4LGCI0iC5e
Uikec6e4QAYFdd0e9tScATmmOZGkm1eqbu+iREQQWXYfyd1QvKhITyv2kj3t7aDLhRteJ9hTC9i1
Eho1DpJGxdr4Qra09Kd/fQfFBnaO1ZG8HAr9SAjzkLF8DmMezPoezkNIXU/vWtIWO6kCtF8QYGIs
OkO0iZLlX3MhVUKb8VEILa7EP3jJ6ZPV+JzK2x2diF7bZgXla5LpEI/0oucj9PMfsCb0H+jxh85j
3qWj2277XPi+vdga7bW3f2v71q+pqZVNdGLZoMtVoOUg4bn3bruw3wseeOSwEyRQL/5+wUiFaPOP
1oVJyS54QjOw5sS36W4DDLbEii8RAkTdKUjX2VN+/On51Qw8oGrf+FsAA7CNN224lW2n9RZx0Vs+
2HHFqIcHC+TMXjk/uoaNrSBqxwpN8swaAMrd5k9WgNG0T930uNF1Uybj2xq4Q+WTZmyHFbdlS8fT
tZBeTKKtj55fzZQCnfYPsQDemnS13ZYh/M1tV7sZZrG/LVGNbF4EiBJ3U5UqOg7ZE8kid4HjcabU
N/Z9WpZ0PuFoUX6vWBDBnykfGEQbt583U+4pHsVVbMcKUxevmHSYWNUUYqgFwaB5hkNd7cWk5QSs
BHBuFvrF3nnNTcFI7HYYisxCqbuiEfOduUh+95yEIQxKhhgPbnvw6yFTMqUvOYMuQJOdxZp7czje
z8G8S2yY/Bcr6O/pNndhVGw3KkCP2BwcGDHzOII6HY0Xo0DIO4POph5CR5m2XZveR4iYyY3Z2BuC
O0hGjUjDYVrNDMIfzVg23k0E/7V5NAtotZsYvwWzZAecTW0z10AcHvKDSbZSApAIEvbfbFNS6eXU
Hpj43YYjEw2pTMMiv/Zumag5B3khVqqILFu3z2P/oDT1pUjcUKInYDq0f5fzBhKA/rPTi1YF50Xm
v5WGw71AtZoZj4GltLdSlYe1ZqBlAFqGsqaWNFD9ENCNfGzm9SGQvQwvIvxY35/zln5jJ3L0b2dT
KgD+aYZiQXn+nP1Z9StPAmiaQ9fJbmrEcKsDfazoSiEcEdKEOTsToF2NifX3fFX/HORUW9KJgq6c
d6+DLvG81RBeBrxNXn3WFZy9pS+kTVSKx9m79Z9IotQvUfMbBWjmjSjKNeBs0Sv5GBnRo7mPBBv5
jEM3PumwML6AAZX6mdyXENBpLinQOLWUH+wuH0FyvAnpFlAGMSqO9pJtnnXsXdq5BfSWu4DFl/VR
Z2g1o194eAFA+qMbMZ+kc7bqBlMrM1F0JdQeYBRB5fXtHd+rMfm6GHc/0bISbpuBpiXi1eFxLrDK
W+ePsVZ3yuN7Mg0jeztcMH15eFzRFnz+r4ajkQgKM7sRQQ7Y7oLe8OC2Kcen0HqhgOBZIS/8yQli
f3ADokTmLkjKTizMJ4w3y+vYqkq5W8+vY+h2X1cwr12XIxZh5s+cq62xRnW5zHbG3/HHu4Zn1Dvx
cjleVDrfOi7lSkwklvWq7AY9U25BucoMC7POrodV9m2YIY/a5N7RQz802yftjYeNjTpls6laR3Z8
eLxyHXEnDrZDsimcYRZJKG96WCeMj1Udy65uvYo66Ai8BIRadfbTLVHbnWJGSM4ZlvLzl1SsC/bl
UgBTXmeW6ziDAUwiIvh2FOE5kZdHoYCWPk1Z3QuAHEIy121vbKmSrctFzmh7k4YX8Xm73qur1qCE
9ZA37aIPzB5lLHEJa/bWjP93T0gRV1mhq3bDfDkv4InMQkkP1CMQ+XPmRcP+2i+nH80XfcxI3mzO
WU42wtvzVnx4ATF6Qiu6MyQSdZZ6GgbkG0j2cGuDzrhKIhxRQ/YxsJwk0jqk13kVW0vk5wBUTpOf
yZluXEsY2+t7e5ihHOPD8jLa1lPEKBrDd2kgn+hVJo4bvsq2R8z5RDkVUSLn30k+zEf/T+F4oebw
25HtrodogDu8sRNtdyE8TX9MQEF8iEZTSq7w+jGTgwdiDTVTLYgFCiKjJcwYS8C7nvtJl1ib4Li9
mRHvtd/easuxA7y0jn99pL5uYgk9Bbb1oILNEw67bAJoF95/dOh4d3epA7N8uh4H/Nf0Oe95+zvx
71cq/z4Ww0dlDKbjC6gjhgqQM+GnHDmsv4aGQ0boXZ5hE0ANN2p+4+HtslhjJKaX/7iOf/YywKk8
EglBEzxtoVkljVs9yb9yIptLZabQK3Gz05bnM3+dlQ7oJGagLzd0KyZogxSrsu1Pcf6bzEzDPBmQ
ZceMAha0g43eu+24cRoHehU3w6F+xU03lRr+0Vzd5xIspFQx1e944SFm+OPggbXtoWyBjpgG2w9+
LdIFg//foq2CIW7YfbV6q/B1iKXGhv7NGsIZ/Oc4g40mMFn9kA5sBFmSTjaypg3jggkSld84Y7U7
z/0sClBcd94BbbgbAP6imzueItWgZehfwbcdXO39qazP3H3w6Uk7rLxv3y3eshUd9fCZRC0WFIpc
wDj4csoUmEZNyszsH/nU1uj4WpliL2N6jxY8SbKbOFkfXvBIvL9xSRqMh7QuNClpjOpoSbdAMGm6
3kyzCTx9wPLjtovrhJMXFw8FH3AcAvhdhZO5fYqXkhPEGkc/rYMCLFt8QmFCKy8uRit0YhN5DeKR
tUXRd5SMCta5v5QoJM30XS0CwWZIkFoMLHvDJniOONnvWWdd0C81VLGzm/ar3LbAHz2tl/wPYVM7
EMaSfiZitUfklBLSuBZRxBYBlIqOJLHDH938HboIyOcFk12r6ptN8OMTpjJ3Y07kLXi4egvPAWKx
O2M1h9PVFoY9LtB32Vt3WGOJJ0GF/TTX+dmmABRQh0sn5B3BZFXyNROlO1+pFPbNvRvx2str9qcW
uP3TcJJLE8pZpJqlUW5We+HG2kMiQFcpCJ4nbEbcZQ2sSHCs01jAZ0//qf5rz+eH1oXlhpya5uA+
Llpff4GjPHgxmuXi9SjB2Ap/O61NWCgGwe1DCcGxrFxAT/xGewQPl7eZHnItrn4Col+gWltLviI5
soiKlLjbAbaLIPtuIEiQg1dAsWLUlwjLbqZb6CvelOMkDV5I8BZ2bgvghtYfNm0GydT3zCVHG/1C
zqRMnv5zAP5JaBUrVnuk+kEWILxv8gmS+WbG3voQMoINjFsdxqgkl5EJLQAI4b1kS1SUg3wjvH/B
0AigYLbkMxF+BpyVgduTY5xzYlgNDOORX66a0GSDUSldK7EZHzITxkfkelQOZmHtaUBI8rQLISfy
KTg8o0mEbnvu0FlHrDev50l9oA3ybTUnK0Johlv0mvJRbBGlf87wFTl87//zxLOeJsRQS7QX6eDJ
Bw32d2L+k+rMGBrcPUfRFnKcB0L7HZ1jXu9yEisr4ZH/Miy8QqwR/dBfdcsqVbumwL7wBV/KAbeN
ydxTgz8AqzC6MbXenBj7L3Ewg37qUlfQUWNhmxQJyjy5Kbv3aXfdKHibM1Dq5QQtW9Wx9xUJZgP2
Vh+oxNnyP8Uw9e2DgFrmtllttWCBbQcxQkbFSet4T1POeopDNBcVPth4T1n3G4zFJuXLB6+Bu+MP
YM9viforasc5vLZC5tJRQLGcEzLOLqc//X2xQgXiPzf5Ea2R8yAYZP2wCAAz2pu0K0Dy6qseyslA
928Ho7iS3RkGKy0ZK2xcaWsLN+aSOehfSnxJnK7ZaCNybHmxYVF7mc6gEBJj4PzyRaX2LbnPPXj9
HFBG+aIoaGrMxoYL9jmMdRwWckcDO89b6s8JoFndWan+Af2Z9HZLjqE0H3cHXGSqDRV/QJ5U2Wcn
Kpd+TAY5HSZ50Bh0UkPQ6wbXV/0WerRlENjUgvMWmfPKy9qdLbh8R8PhoR061w3GSlbBSWJn/IfW
sd7YN7YjxDVFMHPX6QfKL2aDT26+oDAryrs6zYm8XVldkAUtxotjG7TWl5qlFhFWODvjXSE+fAlC
ggvCUqpJfvv159kFUczHmDH/clACJJ6ElNvKqD2duatRB6Lrf+ZS8Y9Q5ZpVXPdJKw/k37+qneyw
Gxm8Y3TPn+K4jJwwf/iz/sebauVM9J0zDqqW50giDHGom9Q0EqhNMLNRceVuaOyOrsOFja3dyIr6
DqJJymDqCfVLY9CkClprRt343KzPFkRd6e/JJREFP8bKN6fJWsHZ5y6UK/TDhCVkjfmn27ZNHgOJ
/rjklX1ibKvHLHenPNSc1m+VTOTmhByxLqE6Z3B4kJfwKpnkUaD3k/ihb+JYfjuetNF883dhSZEg
JojC+71sGV+UqnlhioiCYwsU3vmDJqNMe2WPAnueUeFkrmSHqS2XMUQUMcs5CGHHXub17R5kmurE
glNos6LDpfyrfJVp2vfn5jy8lfVwPF7t99MfXYB6exOyFzTpKV+Z8DfsbJk1L6H6YKiQNfRvOmIB
aZBssiAndvh77cW2Uk1jxz0nqBuizcpNrhngEpiFcB8lypUJOjzyEfG/rgpWeQuzvFHDtl8f9Wj6
gU4SxH9Vu0VnxlcOmyVl3mWY/vI7EExY69vB2HT9a5jg5vMSHH0PUluJbuzGSvnExkgsVBnY+8HI
iuaVtDOLhSa8MH2GAJQ8bHFMfdlgn1ci/qFe1hkFfUCQfiSjBGbKCnq47sAwLVU2N4nGk7YENmPK
RnpqE8aKO1xYQ/QcpXMghUMcv99BBR8mtFJRWSJDq7LXFHfC4NdhRrIIAOqYN9oyGzzaKfcNSlVe
3TpqsZex6rU5Y8+/AXDHSB0Yof05vXvpbs/H5h4+FfdU/RA1iwyWjaoa7zTz3+PJYM1df5d4XOTs
t3joZH1bBSHWfUYFPOVzRyy5V2NS5POgOXaz8lKQtGjVe2QBWEzN+jKtAu3s7B58SHKgevoFSW+t
liwLw6B+mVw53UcBFN8oX6fLkOx734pQiCqie9ykshKOmmng3dBElnGgkoKgkxtTNeQ1dEPPJI5H
qHvhAAGplMDW6F7TgC4QWVzDXaUggHB3pw9U/G/8Ah8qx+dvCvHOFiXSc7XlQYINDE1Ypg5HrY9c
DhYm5fe4reaulDqyLSk4W668S6MSbLhT/W2Wazg6KknKqjXqK06c1wXDGq6q9Mwy3HSlbSZKkKKY
x18r/TQ3ELTPoBaHbwulhAM9F36ZOqhAhy49xJnJvBRKsUPBdzLVn4r96aAxLGqHro4GxIcIfMjV
9OHgVyw2dTRGVqUJtw4SCEoj1e6xqr5XrOxtUaV9s3CyvEtCezmOP+xQchYnG2JgkkhVZPlRadAi
nFxU39JpnNTWjKSl9O3OUQLIjSagS7Irg8nR2YBrM7J5A2jVKRd+2kykksfzPZ442eJgy7e5HsPu
CZEz/50XfFd1qMTotTD6VsXhRZk6HHNSmGbOmidZdKiyKjo7Rwi6R8u3rEAO8dSudmgtzVHIWRzs
V1hcpJwG0T7zU3rCctX1l6DWODGf/Ud98+B1kVQvLzm1nht6GYyyt3BMFzCgEVZrsExeWYEPJwWh
88Yr6g/9S3tw4US7J0PQIPBmexgQ650ftE61pSuxaQDE2zDNo+AynK4B/mYPXGafeSem2FnlwSNm
GnQYaVnMiQLwZXS5aODX3pAAw26bIL2T4AKgZCUwJfbrMvqT2HSOaWFm3uaddZclqpBW3p6rt9am
OxS+F+Xvy186HjJShLWSv49LVwQvleS99YPc3NBuaKL5YStYvjMXDC2ZGWIj65QTng1zFB++Bow+
feiYWpSEZJfWqmxtsG0SNGQbE4eJfg6Ho0znoNyBR7TT6gPEQ7xmQe7KcrtT6+diZnhM+kVHtNJo
DRQYStN9hkAIARMg8xxrFYLXOcsVZrWpDBkx1tqNmvxMNeDugax5MbFwZyN6HRcGdDF9HGFo8m+R
kSqPJUSGRWRiRQpX1Te5QXOXAXyPH6D2CTnIQrVxqxJ78FOBUqXWQiM/HfWHff/FY0DL5m3B4GKW
0JvUnRrm5a2HIIxj0NmlO4UhTUzBvkfYqa0NMUBAEaolaASex3iIBbX3Tcor+/2Nxt5lwz8jVOd+
uBAFL1ZpbScDWIyYiIz3ym3c3nEZtYjt0kZwGr++G8ee1p4M87swp4upLFU0M9eB+lsBnFemFfjk
wkCVYNdcGXXwXmKO9lkwvJnbFpyiUopdKQkWEVrrDLG3IMqlDLfIv9ow33sIbiMF+NcSCDZ85Z4y
SUVtGtBlIfobn3nM2QVo/FJ6Zbii39oAGnFtATGilHQKCv+MbHwoghF5XcGfp7NM+1VwsXsCiA7W
Lr37x2wLTKGHn0fEqBCNmGkpWpQRTP1vEvnsOISHPOLNVh7YzoA6g62uz83YP3gbZ1erdRb5ppub
IsIu7h1ZRNG1/tQaqE1hLwPxOuBoKsJohxwWoAH/7WvQ32DqK2liuNxCLR5uqYB3dslY2a8po5Dq
GUTS3zF5EcUNPzP6r9sdah9kh5gWAylAj30QQPIg7wGz4NA5+RnV1LF0ID6lPz/OaUtHn/E0GGwv
v6laYejA/BxI3v2HshOLrjULVbuU+C2chGgmzAjlnLPYBroCmvpZ4bxEGfJ1+1coB8QrmayZqpZT
I5amp8rnXPMcji55NyL/C2fFQCMHfljMShx9yoaVwHNaFYoiyik3mApy8CR0NztVkAnSdP9KJ86H
Gb0EfBNTfv5IXtFIYPVitSJZmg+080LQJnbF4mhyGsHAy/+Pq+RXRC4ayOu4XZExgzh4RckeCQU3
ah6Aq//FiYQTTeaDOwaeDhxq+agOkXtwHAxZwTi8/qIDSOAWabVZ97yeszWdTeSLT7E5FlAB3DPP
koji9n5oEN/px5SglATjfRa3uFjzaxLbKdo0mG1FLmWnRPW5gpLiTCiVdfCv/D+HLg65Mim3g7mN
80eAPIYVW281wT85iJOmRhfQeGQWFP3hxEG9TbPExyrmMTYfHqmtF7JD7WYLU4Xyf9bKVxCXsKNv
x4BMyqt+A0oRd2qbWzdmuo6/cMznxZdP1nfHdvCOOs1ZC4tjsTrgcVOHT3zUpm9Mm4VrRPLDPnXk
xk+wlZ2dndOOrPrrReemI+8NpsTkFKsNpWRAZ539V/nAXOh152GwKwu29+JoaSiY/qbmS0w4bgUN
kk7d0/HvWqs6mcxA1DFqIZXo91pprQ3s9FrhU0Y56zCg0SikXR+d04alIga2N+xdDiuLSL1rTFro
oWARvum73UJQpLwyy/QAppht2CS+Na8YRz3TWQ2v4uq3VyaKjZ2JmD45NbwrIjUMOzw7bfQJVjqw
hEp5CxQobG9TJfbaGJmhFYJTelcTHJLW3v9XWSuuoipOFunIUKbAMuDHIXTVDkTmJXxsNEASU/KK
BpcbSV4B3GyhgWnLTiX/r0oLaQimSqhIaojyJuSoPiwUfFPuxuvv/WxkzmZVkGMxgQhxz46dcUrZ
XSW35ARggPwbi1hmEq/4lWP2pyKrVObdj71G6Zr+3Ly2mZps/dkD6Ze8CW+Tf3MoJv3tmaQ+UlHJ
mLbQ8KVpvmz7m4UJmRdMH8TFKnUgu6eM0VC2Nh/oTAG960q+W9I/XwI5llG9X9ZX5+ClIN3s4qD4
hqweFFUvl3xLwcT0+U7z0r0CfbssSdQwOIlKxJ3tBws7uskl1grHzybqLyv5m8GsGE6iKALlM6wc
QbdEZzbMdytqcLemebRv0ueAFZn+vlfMRkiT8YrkfUNxljy+NiFmH7bd/42bCFxPa3lNVJqfNLsw
1gelncHHf5ykp6eosBX2Tgy4H0GSJJWSgsX1pJxR6JG/12d0P6yP3iJBk1zZmfPIKX2BKq2wEA0Y
65msVUNScRDOx7/J9mUNFdM4s2Xz+b3RxviNQL5d/mAT3b2s1bWxlhAQUM/RE7E9fjweCVxsO3nD
KrdhlN5s6qa4OIDccBgFCGTrh6ynnfpy0lAIOhpuUYhgTctnX61IbFChlbG0me6LjxCpubOKibTX
ycjMEvTVR748GyEQZ6HA1et+GjslBZ4iduOMPT15bmOfq+vD37zi7ILXHVthg42YCmYdKgRCy9vJ
KbMqoaqu9e9/LjziOu6LAuSvvJ5A6xvV08HaHtxoV2RAJQ3uLtya9BQmRZpaiyieEk6NkdKU03rC
c2Ywh/TY3Hfjbgduz6CWBTEkQegzHDJGoYjlf+xtpaW2LPYjuxzi3chgG67SGhcOuKUFQ+e4pHAR
AXrT5vlFedzIWgKRp0h8dO+OWbe2kqlJJVq1AvzXgYKeTJuF5z97dWDTExxrFYCJoyjvqjW1Mr5r
pH4XXGKENR/R03cdwMyCTxEi/nZeZVnNqxV2Ia4FWViJ+HWWV9MRf4zxX3vUJfcvsykizZ76r12/
KSbpEXP3Ywy8M/9BbYKPcEdYW5P7IPXrkslOAXPVuxH7ZCUgA/u/wQSBVNucSyBtxyIiMiCjrZWA
oszW8HqtXh9DieNoaol1VIWVcpWLOL9mWGNYwndEBj6i8tlXl76on6m+0MZOQPTx1AcnmyFKSH93
ulyQL9RL/Z6w6kUBwQu8Jqk+9Kt2NZ29vp0olY4YkoxKnJbM8cDlF4hdw4Q8iVJvYMFPYhWl32VK
Qi9FcougktPPEcrdnI0JzmX7tfMFLolM5wEkq2i6xPDHUlC5dSTICulqC7zXXvIHKnbAqFnkRZjw
pvyJZPBP2LzHEEHm+kBWrkkauLSiilsWfcmu1Ump2uIdp5c2g0WLnKWKhk5XifbFPocTeGr1axQw
s1u5aT7xfxBpFk3eteRKTi0IGC5kINzwDkGVSyTsdCfFF2LIfRhv3i7Nko57TEyQcvWYj6hEXYDP
8zqNZqk9/u9NdAxhW4uj4Hi508p/DbMt4Xcv7H+DjGKbNrMOP/a4UQRG21TsZzsq9hnletuULrdv
6VJbfpsqw3faCvki8OlcohKc3gl9pE9NcthZ5ohiKXQz9Z3CFrmazinDL/OhsEyjgezUWpQpI+7Z
X/3ZRZCgA6/L0GdA+bTOuzS1060WS2oqvUzDfmkj1YHpqZwazueBstDLkM5XmVS6f6KT917nHLsz
bDWu5of/iVz0A2hEa7Wmk0Q/obFBYFryiEj2h5LunNQk4MCFGAO/OEy6aTT3GtfngF9ERYWQ37J6
vDdlXCAIEn++mVbEw6PrJPiLLH9/YHlmN9oW3uIy8SIRyAOm45Ut1GxbOD0tRSn5kjo4r/cPGWJr
08k76K3eggQH330h8oZn8hfkXkXyEW8J52DtIje2WyzPmCt6V1wy+EyJVKATR0SGZK+3iGuXPSic
uQ427BJ97RaehECXZEEXa9RFvi+5qMmLaF+PtUOd3G8HcBsHjVzEV5pZD78533QEKtLmhoNbp0Iq
X3pwyK7xH8xka9EgsSZfbZaQ3yoTqMPbGAZj3Fm1B7+IFwd+HU8lCvhXo6+jOl6IdpATQcgpWgpV
SBVygybBVRkEei2olqj7YvXWIsW9JVZNmYOZEhghfcjn3/sysdkAI9jRdW/9iRVQo9boFB/hGqNJ
HkcdjppnWsXHg7ii+ufx87M08P1eQZyfHSGdqZ5YshM6dECb7vfawnyyFJRHR3rEek0rOZ3lAoVR
qr8LRnwu5TlXmIao8Wh332pUgK+LHurIsmdVAtmvV+P7oWwJ4tgO4uteAVByFqfM08iux8V3SH/j
Tp1OnEE3KNGtGazbamMIt9WHapLgpQBSNGFyFP9QmXAdZF+RzNKuMzpNiFPELI2E6Yf9vlmO02Tr
bhODcgcG67thwue95YYOni0UA2wQ7OpVVb8L6ywLpOGE66e06jz7vTEr0gzVRFJt66enWgcKOoId
K1bK2prs8h1YB2nk1PbsKP3EIGv8fR+nINCDAeY6bfpmn227GAIRcQ4otqDjmSgSHdgIKPF/uVwu
vedg6XKb5QzUx2jzHx9bESMveDtMYkHZwG7oDjUglTX96kE/pp1rScwJgmXuJ2wQlFAMc25uKq7P
iIZNPnuYj9HxcEC/yGIlcDlL84ErYfwq5Ys7J6WcGQ/ReyS/9CpulcXjb+kr8nLdqB+8E2Lg3wGB
35HCDzvqglVhJf6DhKHinVGKJPX9QAOwIsvbhnfxdjBteLWjGNSvhCoH/PwL1YSOCcrz1xMkOiuK
UhiwCfqLilxYpxI68+i0D4qrbDiLXhvv0Ql5ASiQAPgg6UWcgxCM+xJmqklT3NEgfxNw86FWuErO
0D1oHqjqEw8zNUw5SDzsE8LDZbw2xYsxFoNuNdybcJ7Mr5tfoFKZ2u07BG4KMgDxD4Zuk2exlRsY
Wl4IUkL/mdzu84w8ZYpwv6Iw8RLcJrIXa8FOmCyo4MXJKvmxO5mTf3SUMXcK8BplyPyAY9oSYWPO
ctu4FQFZnHM4vlMbXtDdMvbDthm/CAjTEhys/piTaZ3oJ2ls5F0MYZ7Y4+FDxnQKRG6t7wS6PsDB
mVjdDKAAlZGfNbOWebF+RTRo/YLPkwn9THBZJ/pSOrO56slQCA4UDxlcDnknomy844c6vABNgc20
5bSe8S7HrLHMWSTygriCcQVX3SZZ0Z7VTBNbHpzDowBSyfU4XC7KlQ9nOha6fK/qU3hZGfw6rBbl
jBcbOermyZpUcPpuF+Am2DVRBesFLYKkVX1mvRzKFP5JUX3lRf8Blyb2Q3mHFleJEwLpbSjG/Wow
9By8y/7K0Sq2mKSMlunwo4CZpfDwZR0xa7jXTzFQyy00r9btQNj4U1XxxnUFyaV6t+ajRxTR/MaS
EY49i34VXBI167ar1BCDRtrNEwnmTKDLio7ksqL4c51ynASR1BbDc4BRWkb0ed6K3p0T/qyD8OfN
cqDCMApQ3602ss9hNBsYqTMBINRttJixzhd61MoWGgRfXF5w8WyyBgoB2H6C0bx6k1RfsNB9Osk8
XyMGeWqtq3Z3NcBb6HIvyN1pQCg6VyArzGFJQfGuyGOZD6xByVYEDkKNp4xwXnH+HeBopzsQHK1T
m3m8eaTBtd1X7RaYwzY/+zqVRLhrhY7QQEtKTZynOHzkZNFShc6Pu5RjHLoPS+qhJdYxNQEHy7T3
0qjZZiGHWxfNZRdQel1R57Daaif8cgwomS8byxdtYDO0imcXBfXOAmKJD0B/b3uOd6Xe+Kf6HbMQ
IBpOtwYmyPI5fdjyDdjIMCoxGNBlFX2Ht5GnUGObFbwCSz7QXC0mB1ypScKor0WregMvo9Lhu8P1
Wy6tBdf/DSnEK/0BuUKuyMgXFnH19dTq6BBcEb6nSd5GhKRnNOQZCFqlL1xUgah0S0vOPv5tvGTS
+/4XCdvG2fwoRcEBLKD6LfupEl633Br6O3l7d3h1aeTafOziTw85Jj0vFzTLWp0pssGQ3y6/n69m
hbphGtXQqRGU33a8IliT8Uro/lT2oChqnkUXJ1GFVfZRUhyVB7uAI3SzgfZ37BRXhwwLIYR4FqtR
hY3RRfXJT+wXvM8tLMBwNsRQtYQHszOKNWnBrbZFwLlAk4HNzMqdQEy4KxEqA+Z5dC0+aEkg87L0
EaFbUoRqydmxJu2HAi0NSO9v5wrbppTvL/v/n000FfCMd6obbwc2y9q8QrZVLhiI8tbIOSsvN0iE
T1kXMS2/4vqrM3t7+EpaNd1KeElhYgHK1WLVU40hs6HhLoa5XIuoTX2VoJ9mNtT5KmqLvY57t629
EXRUvB+gDGmWCF+3+vuMMsu1fjS7J3AuqMS5AnfEuGc8GZBTRSAy6hBL7IXSjHfwUsUXUolNi/id
m7Le7h0xnD21tUdSPxg+ucIyqw01s7oC3LOZWQZpmVS/cgJtKLkq0f7PbRcbvbCHJHDIajQQlhDS
3vxO3/wvMBnmO4r68Sghd4V+bSPPRh2ml2+0afVjM8LsyVgrb42hsg2zoK5la4HkW6IBtedxEGnj
CCyfOo9w//7C5eXYsrEnKzdyPODg9hJZ6zKoZoPdNy/yCLfpAnEQU4GXiIxW0rOWfyPD+3U/d+el
QoIW2zuxLO4qcrx+GtDXislSxeB2U/7SrmbHezol1KfPOUshAJyX/mt5GJQjcVVlPPwmzTPzrpBT
tizWal3LAymKvz5R/iWXR+b8Zaid3efo2q52YA4K/YcW+UOyEzCpZNeqH5ugaCWwc2QuzB0cwGRH
Ycl6Hk4mVCCmScgXk2w9UFveqykD1dZCbsYh6Sf/TtHtitTQly+CGtEN2tLJ1vBd8qiVZ2Sr2IOj
qiDpDKcE3EjLrwuUiAV9WSLMv+mz9dPTMX6t8jrskMg1dwc0rIJY6zXyfN00s9htraB1CQtv3104
pJXG0zTj6Zt49EBo7X2HFljNnkiMK/KaiAXyCN17Nlh0J+hWXHalKmI9sFy0Eiibj6+cNEbWVDcB
UT4Jf5nwMaADWfb1dES9u1hLIY0few6MQ5fCraPP/xJbK5DSE6k28ltHGtq5ZvcGh4u9n6Kd6JYc
rXzzcNn6fdHvTY+ndidAIMJ+z7KmMsu2Lysckav+j4w3WUo15BsN/m8oLGSzWpok5vr4N9BCylob
dp938PpLZB9+pxRwQPGK8W1JRNfcvuacXMr/wSuig3iMFGByM1mgk8pOV6teB1Ta5hotYrf9IUpB
N/YnI4IihcpmVMGhhhuIQ2UiQNThSBG6tq3YbrXsCzOAHqEzvfjdnKNsiooF9TjeG3qfEllRkIOK
HfGWvocewPeC9wRFEIHFDiB7Vmvy3maBKkNF0X30aEQlrcFNzp4qKQ5QfV64FJLJOlEYLxcLB9yF
c0cQn+Emt9R0Oyqnsh3a3hENFoiLxHYKwB1ToU2r+eidHy3WSEdlAq4Pfh91ExIPFCG8IOj5msRc
eyV+T3z5sIZZ0taT5NtSTOXFl9YhJDloqV0V80ubtCmYVD28PHQHiXtgCmKCTMdHzVctTc3OLJzM
X+MKyeV5dD7gLWEVyDyp147/Ck7+V6yWrn1iIzkDOI9AGZOSNGDOLcnyT6hhXu3I1YCZg6Shaljz
vOSvWd51jFbJ+sx4mVNQ1ww4fVbJM1bTfXY1dvqGBKmp8DeSgcm5RJltNxyKzBNgnp9ZGG+Du3NA
Z+xCV3SC4LV5ceR86De0LqbfosZLVTncY8ClqQgcSnQyTukbWwI7peh86DZHy8DlnzcR55rMOLwR
czllefnqCjDrdQ69/ZWhwjSnwuUUj+ocf36gWSae0msdF/Psqaa03VrBZQ8W2jDgBeTkbrzBvk67
j25k+kjJYzlKHqOTOFLA1eZPwHoTxaI9hzWRFTxrTFf1yGCAVmbNH6+lb057OYMVO+Iy1Sy6dAiq
/j9IPMsDZpsFQdNPyvdztsjaJdJT99jLPlbBOW+0iIbjDWSG8HEvdCQaZsmmCwziJIqzLmN0Buo6
skbJPBABLC3swQVRvpG+n7rx80TwLOEoqgq6SQlvrSKp1SrTfXBtJKWYNRfQZkPCzc/bDy2aOvUs
aAazcdKc7S0K0xZSPXsIdQNJ+pSuXBwu8IlA87+mkCyu1zg4O/NKJNCy8s64lhhFGWF9eVg8+hIl
J1jXmp1voa0LVbCe9V8rYzH2HQBpg85aVhFqwyvmk3VQujHS3ImR7sSXo1VWdfmMBnqk9nsM0kms
Q38L4q4NFrFCu5Wng4jKxbtLtk2e+kHt8xDtIAXI4mjBJuRMU+WZTxciQBEtKXYCZ+FSPMAayXz5
RUKwFr5aIJCK0mugJ3sbndM7ZcL719a7i7SmgH2hiGF7GYbuSnOpZr8Z7y70E+tIPZByLqXxYFzp
L6geyLsylpsjdc8WEskgEJaH00HONmG81jvAr+vt5Gt3LBIZdf/g0vs2PJ6RGVo6ppC6KJ3z1Z/P
bKnNVEAtcjTCYBGE6vLPU03XHaWkBKe0dSKQmldhqrExk05GqGperh2gPs4f17kQlUDTvZwg33sP
ZptqmqAF1q37xBvCj7FXRHa6Badhp6RAdVf7FKq92cEZXx2RsZlfFw9X5C808yjbZuyYvXzhlwIf
73kux5HwjGRP+X0pN8QF4baNBVpi3TcwvS+G54TuIjDQv/8Qmy+0Akusu0x/qwAhPucIt7cXug4O
5iGaipq71YpB2uhOG9vZO/vC9N+xSb0zv/y1o1TgkWrU6UypwNJCOlDtA+z0+QmZYs8OHnifdp4u
W1RcuqB8Ocdu136s66lbVMo7U955266Dv1DWccZfKV8Al/RKpNz6Gm5+2qNKJZgW//IepK6EZ5Bn
i5st9TxS7F/IYnEVbUvfrerxQP40DDCsNgUf/6a1NowTGbmNJBEl8NJqZlUWpvaBz+12NY3AV3lL
R1yyynQY1TL9vcesyPdS/e8jc9G8Y1+B3/Itx6DcNfSryejymDKXJZs/CQxpOVyblJHcRnMY/lkz
+MRUMcqtcvylDoIQM5a00WkLXcPEVF+jHiJLbLnWBCpOXK+ILskCwHgR8GOmU/B8VZIf3Xeg3oIF
Og2ASs6fdoNQwaac53H8D7mE90J2tVoNfqJF7ALTsZ7trc6YdfhoKZoBhJLhMyQAW2XEEScLRgv+
K1QLf6fMvj6r5K3X206f0xUZS9avlh8Wkk5vy1H+VGpQI7b5TSl57gLHfQYUQiIGeSB8T5crmkGL
m7z8B04HoN6znrQz+gZFHs7+6DnmpXweAsp/OCMCW8bMkXArzkolU/T5aWBPXNC+fgXF683eYBBK
G4uFWh0TrzgQUwIOvKsyP5qDqpGJsFI/R89tpoEV1l4EcIMbu9gKtgIYvBmtV8Rg6GH4j6zVpf6p
W3oNhrJEae20bEqUU6vjH6N+ddOsq1uAIlKHDM7X1fg4H+LNgQcsUegaa3tx2BEAyEvBRcHJoVLg
j4edRtaXZwXP8RZnAgjyjErLHS4OWBK2wXAPJ/OpNet8tmy6FTQXQslfL+R+aR1wA67HMU5/Bx50
U2liVEWXEODtdEy/qJH4rFc4CJhfpDFLi3fSWFF2cPw01caqTmSWFX3wfsGREQsYQ2XfSjZGtA7u
7BBbbPST2rAs3nXoIGde2Q7Au31TE5re3GYFEqgDqH/A8KZQTmVlR9cGkIIVJTCKwzYEK0H61HZX
fkERrkI3O+3nCAgvk9w7Nsx2jkknHqVcOAmTxEIXk5fcCJmzYalVVDlprsqqV6xbmkCi8jvwNjTK
xnMUMKttRaxUk/pwGk0tilUJqINwAOLnr18gB7KpDo7R8i3Ytc/9kwkeiBLIXL/Df6Vlhcsy1gp1
+Z1lfCpOwwI/SM3kWmV2U5Fe2kZsZogUUdeOzSZbBqELMIsfMrhQiNiz6H0XI/dcly96gJhYksI9
JAGHBw3G5zc281aH3ZZ6dJrPuaBJhZ7tqkBrCqpWZsvqkm5XJH9bkn0dCf+a35+2WMp29loaLCzX
wGoz0plCr5d3BRjPQQkeYlvrfKMFdS26xpeE2GgW306aNsaPVod5HKlPL3S0Mgdg6oiioz6IHaVw
wZ7Tdzsk6sclx7OW+gQLcsKg4XjW5VjLYPGRu3Vk7SDZoQ/Ns3lgctzrXk7enTu7Oa3k/jY41gJ+
f2XidKpoSau4NU92j+L7CYnOKzB9PIhvwNqrBEtrDx9qO3eCY3CR1sxMOymDHS7mwVEgXt10v41c
lWxGp8kXac7+GRS96hL+XQIzxY6Ubg9hjJ79x+N66acG7vZmenzbE+VN4oh7yrX7xwpny1MbLjey
S9mxPWuzgjAFsAb9zMlGgJrR4Fyzgv1BXTr+gqJBMqFeiIlRdTPkQozvTLJFbZYf+HwFzFEKkBOg
IXcmBhr9V0VX/x2swmF8fkbrnKN2zGWproDOKZmJ3AZv29/bJW/nHKXZ2GIM6yJDtbefbI2ed4F9
qnI1Kzqob+ExSBNhNx1nuJNw3E5iBxER/6+70D2q42S7Ia+6i8cnmVXm03FbDnkRcZVwdRu91eGH
UgS9TIVParMXt5lyCwkiHJ6RWmUQof+ZKE2WMKqaQ0Sf17x4OviHCVnMbFJWK2gOkxdjQzvdhc/0
XI+fB3fW7ApTI3YxRAl/V2jaSBfBnZSfmVWt1l0RiAj8gdpNR10gY8Xm/i/O/wXndi6KNvbdSR7p
wP9WE2gy8o0LB9Dcx66PztOsskzOA2dkTV+R9MDB/+9ANf8eHi5NPpTBKVRgwEagqjBUrFC/Ccn4
cCw9ZL9azDi+sXntyWIpt3iY6F+QE9hQP4siwieSHp44VHJWrBmcPYBLOpRoS+T442eKHdP3eIEV
13siSIem45ix3hTS+5CuRXbuRv2LBagH8bwSqGKq/0bZQjo/tdHIkj1qo3GtUhBRCdS4GYwvkQNK
9qS/R/ImitBf2lzJEuUnizMdRlcO2FV1wfNh9y9aEqAXXOfKyHbsgYZHUITYwBIXaJTlXH4M3QRL
2BRDC8eJGI0mEq50U8lG8+XzRuq1DyuGa3jL4KXrD1JxY6+f6I8AW0KIzhVuAXFz9zpVvn8QUwY5
Cx9ZaOQcbX/iEuFYVElCWKzxAyIjHHRClEOsQf3JptRz+Uv5mNayZ9O6TN4FOe60tfsrYCq8u9PO
LG1cEY7CBoRvLWneI019G3s7PkchiLs1iOV1tW1+FjVc7AQA6LOnAy22TkNxBdZeixUvyaKJZLdq
3LcztQWZhV1yNJ3mvfkJGuTXtvpH+nKtXpPnFxYRTjqmEX2j+fcJmv993zKMmnbLxWUIAj5NPlgb
PNeW+mjidzJg111CTYi0e8/jBdx5InL2+t4hEMbC+RGXecNW50Dzk7H0aHqJxRdU2JxKIji1x+wm
Q63eHEJ15D92TDT7DmaaL/TNFoKX7XaBBzLHXlWPBadgyZc+FL20yQCNDMBnFSWIxFDD11UXMV2C
Z58g+IjRZbCs19pqzwv89VDoGidnccM9oNb20EJbmhqtS3GZoMepABXYMhmP6lSHvU9xlQC/C8F8
n20MxUkmzq6gJ58vtR9qtcNCVRxORL1iZd6ETICqgShYutS36FbaAPZ8RB4qRRTKGVS2dL5seqIV
PK/dV62ubdHe8D3V+kw+HxJ216AnjEInVtwqlOR8gGQ/1mFIbgfQ0e1JEDaospbHpDO5Y7K21oac
w3m7SJLSGgMrNI5zx2wbeKUmw9Vy74niqQN5GPBj1iEwKrqxd4xPnSHIg8c/6Pl8Io0dkprHX6BQ
8SYHdW717Xs4YjSbJR+AwFUf0icMCs6epRnD9wIXLpgciVtvrRm2VJw8TA9ClwDUjA/0GU0QTXPa
3zi+0+/k/skPBqxqA1bxU1PETScQaPOtbc/Je7i9GgVTPKt110fgHzbL7Ppwt9v9sAG32GCQytMw
Ve9oav+PnMikW+SWtsO9Y+VMZw8e39ttZ5zlpZm8NKPb4MpfHbsZA3070pgKUxIPJHQYXUEh43ea
Xb4cWkuh6Ktk2lfpvULiY3eNvk6PPnoe8Hyujdt0KAk5G4/AmINVRUzzmtzgyFUU+5E+BanxMp3m
H8CZNehDh+GxWAtoHlbiGOHZZ/cRDHrGp/lXEq2SL9pNO3VmR7B4cqda0I+e4JXTkJZq+3acDFLH
26GKvBitemeepC/3A1SpohoRJVPbL99xFSAuTYJcuIqCwy3gzzGTYePoX+UusBcivUMoAgv9uhxQ
LKTCgkrTJlzdHtnEZ5XUniLBntuwkc8KmrMIaiVKFkDrEO5RHJgGtDkW6OgoHzaMsgg652jil2lx
DrU3ISS38BruPuZuZw6vD+dLJJ4xye8BSuEAEcvIPa05t0SYK7QvA3E2T8VSTbGzRoMY0EpxHAqm
90ON5+1LoT4nR8vIkDdof6pD1QNvSXucpeZeITQ242Kj4+Opi0XaG3C8TFCxpkifWKQ1CIBOPAJM
3PfsY4sVeQkUd3GcdfkEHRM1/j+N79N4GHrJ6qhxkIGxqVWVpZ3Ja939qOy/qUVKF9fEznVgrYIt
C5UI8VkG7M+vn1SxkZirj2Hqt+kPT5xK+UzDnxDioejWGSbP/iyZLsLG+2d5ZjHwOza21l/mLCZL
kduT1CW40nuznIlApWMpfL6QBa4OQf4iK2la9ITZbh2n7cy0eV+GkFdyFkQgCXO+SEWNjx4Zy46R
yzYmb9x8S79eyxE2EZq2gI2QUGBqaAYOyaLRoFcxe7cExllzRwzR9XR6FNRsj4wympQnXF2wkEeB
/9YRv1eSQJ1QTQiU77XtHZbjW5H+aH531XPDQKOGdJW/NRJPfuxcW4OZIGbb4+OQUH1lZD1snM7B
5pspid4lutdCTUG2YNBof5pKink0O1dI/4Y/mLgO3LILedUmZ/7h14+YCrRG3GpsgO0SzQxz6rQy
s2+e8+uY17fv5Qsa74bTgLP77bfeLEQ3s9OdVsfC9p77H2XV3GlCYdAKc/QZEttndOQXFGexFyvg
p+AiR8l3YC6QCDDXMSpx5rQs+w1aEy7u3Kool0LKO/840HNvYBkgHZybxBcErutuYZhE3pbSsJBK
DnZA5DLjeMXtYKGKMNYF6+3TjtHQIK6kDqhjrn6QorLuIuHvheF2vLPlYLax8TZETtTr9YnznQD4
u3roxlH5L6Q/F0V16+HoBomJc2enyRjBP7uZx8UxS8jFc1w15b0Y3LYcHHsKg2zWLD+84zjIrYi4
z0HcQTSfXEA7ZiUBlgs3IzdVcffMN9nXdHCtYnuIJHAqdf3ZywhvqeTChFAqri5oPF+rob3reZ9S
tH7ZcNtGzjwWo3MpAONvA97o7wF/B3LV21JKmXCcyAzJ68FiGCs3h5wzLiFNHzgc3B0Gh1L3LNaW
UHwJi983sUSAd509mnFt3OoeeXOiblkgysuhynMLCi4UHYd0bhYo0XE16Ps/mdLChfG6kqwA/6fa
ebvp/MaLaGR8Se/UY3DsOob8Md1Rd1qm+RC+gxMahi6jz+o3e7hSg8nLFH/CCaMZDYuJ0XN8+jcW
x8JEBaBMFi4+DeuWMHbaM5z2FbWkqkPBhj3ZOnzxlxGynzgHT7G41acMHQTEFXRk5wqKJ0odSVWm
GyfK7gOXwpOgq2xN4s+0QFLB2iCvAuPrzvSvwsjTjKF1w9+Llz8BCpXVtV0ilkigqRvljYHDRriM
1L7N8jAAnN/nWznRJrYUboyJSxPyIpjwenH3eJ8ka/NbXIwBoEAPjfrrntxjq+KYGlhoGzWc5hZ2
xaAX2uJ82uNYz1MDF0TG002WHq6q8YFTANXzSxvuSz/LXajGPQmdDtiDCwfV4FbhEXIXxeWjvwLu
NZDE8tPdOSEjF8Y6SEEBmyb5lv2UqmNngYyYF+b1YBLrfUZk/8VPUInVSoytCRBz2+fxKJtKAYtU
phouHRb0ROYdWvOrzEO5mwdax3h23Vjs5i1ligYxa1IrhBGXY/zAPs73s4q7kWT8DHmelAVEjDIm
2NICmM1ABvot+0ZtD/uxceQtrgcy6gYxEM7K0rtaIPg7erGbR6YT8L5GesdOiH34rHdGKxyK5enD
/bkTQFnxZIOqKSdclqLkSTk37kvwHx+GHgdRd+2377w+JmoIyxCGuCRCaLhf/OqogwlNPuTsxIdu
C4VV8lHySZ5JWKg2k9mQO1gFnhnWMDbCdH815D6oyHybzFNFCbuDv42wy8Pw/upICIBxSf5PY742
2O+GSR9EriG5mKzouB58/Ebo/FekfzS+c2mM0P7Wb1ufDDguKNzedjxBwy3UwM5pAg8k7x4jLr5H
laJC0hWTbYt5vqECfuShp2TajoCnBEda8xG+Luv66YNUgojDRrNBKDob6hyXftGuHcs4uAIHgkU3
IjaPkDcpNNHcuSKPSN38YbaWgzFRcXnuig7uUsyptvPOyq5wkbZblVW2ZYAksaY1PxcL1NbWLLn1
mS5rsSLs9qoHRhtGpTA+/H8DaGTJRLqSQaDpiPDUY2T9NpuTyehg6Nnugd7HxxLxF0OqHPlCzj7v
HUYr4gHxQM6+wfHQ6gFvRDDotwqHb5AWG/K1nl81MPRV+pHG2gMBQK7GbmaRT5B2pPXrs/aNJ6nP
Dr3eqM65mwaYf0NEk/IWzMY3vdTlRXJE1A+7KFA2wejJtFTC1Ne8ZrWR6KNvZAqOzrdavyS5o3W8
Kwmcl2T4edV3HY1BvTQz0Dvx87aXkEsPC9orWrg8YQKqODa5MxgFYUz7S7j6T9OO85HkXnkewiJ5
0FNRF+z8hM4Z1eg3tia4rpE/ZvuXbdX87u9qD+3mCF3L97AGHveeVuph5apJUHfhiBadiKmfO1Jn
S3MkUtOVNOnz9ZS31bfOfhaFbP/xeCtUDYlOkyn8+UZB+db0fdaYtzwLG1zOez3s8pvd9D0e2KkQ
kXWcusZe/KRjvAajfRcz5QiQohp/jGy1Nx2QmZPHfvzakad831j9cn5ULicoIHIqYXgTIsAu5wcF
fWZn6/0TVNCZ+6QelRj5/iRQtQRRZkHpii4z/pLiAWD4uYOkEcC78l1D4q4XOduufRujM+OPGOO6
lp4sLHGsggZvPAYyYeK/44l1G3Is1TuItZj/V8ltx6LhrcTwjBgONr7U2UCXQiSGj20o5aD09dFV
IJPgfzZU3HU3UXHsvrNqt2EZ7BkqnHM6zqMOl+wYJsBBAWplP6CqQINfRmOXDcqdJkSJHcweQ+KX
QlPUmDl7abztny8OxCpQvmGguYQM0xf6X6fcEpEGdPXh+J0hLr/jG9nt4+19Gy2+Mn4SHarN7Jxl
hj/B7H2Q8dMwCa793lknFOMXYOnbcTXLA7eF0Ba/yn9G2JLQrGGPjInlWmfW+cf9vX5jMcQwqq8I
CEJ0MtmIQ31eNaLHf6HQuOmu5OcSBdFeb7hcUQO7IXggCF3QB6yOcLwqBGxmakgMik91Ul+wb7TJ
LmT8O3W6DV5tIf/Q2T5pVBAP/7/6hGHBul83aC62q/E7Qlove7HhOSdqZ/kqHudpSlhauff7YPpe
aMyRhvrFF5V5Wiixj1sE/J/IAsxcubkyLe8GHzwCsMkVJGFTO5KkYn3FS+J+D8dwP0ViXfzZHCSA
W7Re+hsH2hQeHTMOooblt/aFR2vS9xWFK8c5R02CcNcqSOdI/XnJEGNTMHjijxArJLROp1gSngSy
KJ5QPhdoQmFnOJb/7TCoZFdkrf17/SlV9uUFZAOeLZG29vTd3b739jWBBRRi4JQb0B4T+MZ2vWkX
B3wxDSU0my5IxEmD1qJNS03Ak27BhAioW8Mac014AzUiXRC3Y+bZ6BSZIZJf+c+TJjAYFXSv32TB
MnCftkyrICdF0QfeJGwcmGP69WRs4a8X/W/RgiDHsdFzXCKMaftXDrRADGwGB+YWgUYaWk1scen+
bUY0P2IVlnEFXWdhmsc32o0adXch8B+QbvGJu2UKXQ589cNEQ1mCgGWBGFH0D6W3+kW+PSIraelM
OA8HEtBGo/9CWl8MJ57J4eBHjhwbvFuhcRiqXRSscvXhSnJXJE2Tzx6kFssaa5zyJnFchiTSB/6d
al1xioKqNyKUg8ZbfeUj2w8xq3XCkfPXSfQ8uJQ001z+y7pBbw0g6+FM2dIVI8tRTIcK25bp09lC
QTdaud17bru6/nLGSCgH6N26pqtOj8Cz3N8Zjcs/C+GvrOvFTwya3zTLsBjmMl1vSZia5j75+sQC
RtroXq/p1GF72NVoLPRu97UADh3bud6n3lRe+sipZ9Nj8UvhD/uptMuvEz5y1oFXBZSegYL6Gncl
sfoUfxUDqQZA0mxzrl7soGRHsdu5eDV7gO/D3zsh8L+5jzQgsLB0B+i4gKUdQ44QLBfmr+EUGEUl
RmhEpRS8ICIrllkQ6OTiq0aXyj4NXJeXD5MfRKNAit9ASLVFIDkxc8pJkMTSRFpSSeEimScwqT7U
TcU9S0L9eTHrueW9PIg4lqdCUo823svY2/YYRH/PcxdGU11Tbekujcu7NIrxGPuUykpOtJQkRo+Q
dSHckCalrYJalf4M38XWWjYjHMBmjDHJWGuAUZJ5bmMVORozyjqGcZtdvUkhSx3kttSrFPn3t/7q
viFpb3IPz0z7+1n3aQT87tj7IcPuZ7gu2D5IMJmKtV/23fGz6eU0SUUiL/7EwMu6AF8UkvrvaASv
VLlfh/6yraXqZO7Lx861hLewhS3qGWuLyaWPnM59pGQa208+6pdC/u7hq8D3SJ8kuCbC23xzJYRU
KV9yydXI3mO6qpyRwQMakKoqKfSez30WZ4I/Wf7FAy6G1uyrLsgHMgCJXIl48OThRAPp4Txtpmxf
dWec1+Z2sk1MW6cMacFBNRKJF07sVzcXz+Bk2cmfz9a5vbgLvTFfSKEDE7VXxbAYsd66DdHSBcB3
/VpJ4AgDQzs2OVpPsy10ffQFijeSL1/rLpk+rkvW1ISFevwHjY8yj2mkem3QujSoXnbnpPSTsxk5
lk6zvJ6zbItDO8poQUap6NyLZ393Tr5SY6JEn70TKFnMcbf6DQBHCGWuYef6XKA63L0oO/06JDez
2eLf+ExcpcX0CnVprxvGaDezJIYOMQMebPewvS4gXjAveZqTAaeeSdTOEDx0n9XBv1JNwb5A90KZ
oAw5gq+UembGcYU1dfXeszswzklVgWI17OsTcCwROJYqsjvzEnDicHAj7a0p7ahp5mr16AundaMQ
yhjQj50+FmIIyCf6r6/K2T69pgAFGO6jc/9jVWerw5P4VclfRTL58iw50Aq9fe++77sY8mjSIYBx
avLk5qYau6xM/0exwB7z3CIi1xtF11ZK2FPxaStTmRHwHKhYz1iiBhK79foqCAcEQVSN5v0ENDoh
w7/IXMsncnkeUYUEGlBcnuyCYPEQqFKA4j/YFqEHcsKO4+5I6GakfXSffbjx4J+/hrEEg2lBtne/
5eElTxtpIwcxpjhtyIkVDhIlQ6XPVJYhUHEUTzlrOeTywgwqZf3rHgt5a/3ucxnSFIUPxa8vW8qh
O+eBcTpDggDhjoufs0hmJY1XRuGpjAyk/tdmqRsfXulZCow74fbMQpUOfoX2WwPxTb8tIyUEq4Tw
dLcsB2i0mUX88CJqAKCtGf3/mZOKBtuz0zvf1G2rKAIMG8vuetOMD+ljLCeact3NCAylnRvUs7nc
7qAWd6gCeHDB1ozHsXKMVAtpvTqkdDu158kxR8Xr1fionQt8cfDVwe/ZEVIh84yX/JHTEmoJXskY
qHcLiTfPdHZTIHr4ZiOnor1TnZBPfqRrIm40ineMZe9AGJnJNfVNQur5cqb0FE7MMlKO/kmQ/gkL
d8FYFS+AxW7WmhwgdZ0O4gQcE6WJL4XHjRxWn6yExx2fyZCrr52aTOIGQQSDX9eiKgIo7NMwKKYz
Yv35GG7gsgrbbj9WVLxCUOIFj0WFK0J1nwuwgb5PNglot0DcVzlb7WuR/6Y6dUvB7rUHFzcQ9S3j
h+7Rjva9CNUiw57++CFKFVa8cPUGL5uttWqDmVqG1qyxZe/Am2PA1euTCxiwoad1n0R+reiyG7Se
IX4MxMADRj6I6ZhQ0metRselNGiIqdyEwbynAVhFXy7ulP77u17BXdEaYbZWhhMLKwL+P+u0DeQx
7tnH38vgjNWSfzrRDeOCJQPTO7fG5NUK5QzY8AZozw/vrTUqK0nTmBNyl0C2fDZAx5rHVhrqwL2c
64CWhfgHh3wFAASm9PN0BzktKVtiRRs7RHT12usNkLPo5usnNQhx80RCUy37pULCOh69899a/+Jl
sq0yrLErgQYK0vrvDhgTk66jAt8Gaoiy6qbMHnxLoRKC/FFRQIsFf6XOiR56CqyFH0YIfTq0X+hP
7NFQC44CYTNaYAdHtuZmnVEVRk7qJGGtJwl0NB23czWx6gZldpSqctolSbfOZRu/n7M6DzWu4j17
eBMMsfKGefao9Rp9IZkkQM0Fd0lSO5k4eDWkS2nhomu3Go105jod96XGKb9xAqEM5jjyZnjy3soT
crDPInIENEnBQgTIKB+mcidIt9yRcY5H5WL/sEaWq37HeZmo0SObLj8weZOPmZXwd9y4+0xVzIsA
fEq7K6li0s8jTX0M3syW+fsZeZeq7abtyCb2Q0FPHRC/n1b68Tw+vIu5U+T626Ebl+twWpidj+md
PiqSVrEnd2rsxM/TBJO4uoJRiUdSWZZ3/GkfhiTA9HB9wKz2ZJGUllCi0iYAhuOPePsOYluJwaF7
2glbCBMwgx7sjtW7HL5Rnp5cXxfErR8Ktd1ea7dTj9+NY1bsmDKA3jkyE+d5so5UNpbm/UhfuWlw
N4BMLNdNRDmY6ll4DzOotA53X8rNEUVYJq8fz021HrZAhRopZZwaiMNBIWZh+5NrFn+sPuo/bDMY
l8SjsCE93uYZFL3KbbK9LV3RKX3084naCuWTa6cOWjHEDXc1RHTsxXtpHUBeyPFOKf/pnb1BLdZZ
Vw9AVbjEtRDuivlY2tMXlJT5kusf1mgy/PYmSofpfaRson80A0DhRAYU4E098DoeslSFmv4alUQ4
NfyokEmzsT6MI7CrjaX5rtn/U7X9xaN1P5u6dTxNVwcjOORvTb554p8cQ9MNKJUD9O5+QOsW8BDg
Y/rR9xtaLwDX+eQbJ+5YejE7H11GjKb4oEq41ktEmmHgBUiO73vNceIQJmKX3dQ6aMUQ8ny41kQD
0z27yMvRlceo15iE69GDNi1lBy8TAT4AxgXonBw1mi9mkFIYNNHWeNuDvqIJl2iNFwc2aKG+idTb
xXxtp3qHowYV2pikxWwovIWR6J3r7nDim+mJ96q7iq4HtXgIVg151XeOfJrdscqwDTeTeta3V0Qe
9XrthDQHxevploYAFeM//CWFLLgRKoh+SvvXPKOANuIxCRexeQKiRFzQvUcpWusLtWAX1znU6K+y
d8jIO55UKER425AsoZHMm4Z6pyu9y1teYHwcerrBXa9a9I71pL50LJFepFudh+/wMEcjFVp+Tadw
rHwT0EkJtPN5xHFwDVagIb9wMciT9PLsQyBqc5XU9hEGx9GmlKpjCPNUWkR8yxo1/P38hEhnx9tl
xIVWETmrlP48KmSYOP42qtafir+LQk4G0qbbZUWno6pBLvBHeGl4Knmcqs0pYzi96HdOQd06RBwz
vFHcVSSYzTyExYpPxvReTJI3dwWkxjUnQvfXRGMCK3+jAoAUI5VQlbhJ7Isg7aESmtIPO0FLWsic
vuoLBSX4GEsmo1pnUvMg90nns97D+uACiv9Au1dk0CB8KFJi/fS+ry+XR7qTlsSjrDPrXnbLgn07
5r8UIPCN4MIZrrn3rqG4jFYx8knGpSsrHQHZkuVDCdQlHlx07Lfda5drpQmukTFNIzBhZoDCY4tW
3jUBCDWxJmcGmkOnfrc8i8SyGHB78iel82tyfHoXi81I3hlu8QgvRFrZB8yda4dkDdBYqWm8Q4Hj
ij8//9FdrXSGGu4rK6r4WxVjTAygCZCIJpvQvsM8AFwaxVdCt0RL+Yu6OOLljRGRq6TzQRRw2cGT
k7HvKttFBbRPMjALAncb16nkJ3HRnU9DZ5zdePhlBQjEr9Em1KSYdUl4ZdLiSKjB2bwm2xCBXcvF
EVPYSaQtyOUFZxhFa2Wt9aIrI2DwujSpnpoPWMIOTr1ejOV/60UlICC1E0VIlitiNjh8eoQpkj2N
zPHLYxCHHNGKsv3Lxc2wVpHJxax1UkcYoBV8MbpnTb8jKsSVdF7bV43MYkGrzYAMmXC3dXCSrN7z
qRcWOM+57ZUfLDi1/bKYd5rMn4dHjbVvcstRemMKJ5dYP+UalnC6jRY9QdJwSeRlUFVV38q5eUMH
i1YN5MiVINH5jx3e4GzMs75LIKvL+IEdHhFvT2c2dBzy1DQffUPxpuk720lEyJC18tMxz4M8DIlU
X/61Wq6QJrOIYucq6nFMasX3TVi2AGzvdMOP7zU7k4b47EsYA5FlxaidXICjK/vCRcC4gW+krtq7
Z9KgVPYVGbdheUQkRKVrE39uM6mT95H2xVmQP1YEHqmOxUocNyacE3MX00225TEVr363nG0zSDUv
WTzGSuZUnWIwUPlYbKJnynklZhjR52fxV3bgLT4DBwLirV0rNAY9ts1mDuXfMvuzHmVJ08hhOedp
h+jiId70gkQLaPuHbGzQSRHzdpWln36xS4yR/7dRtCqk1PpT09IMbL1SZBq10t8j/dDdnJZU3Zjr
R2wHQR1JCIk/4hd463cl/6Bt11iul8oU8UpcRe+AnLuwxcOR9xk/txXJIn9YrWjEx+hz9Z/sokha
EIrKSvU6Pd0pGpFh39BaHjOplTE7cC7w2TZxQcR4cRvdtZcRY84gxEEnEXTOc1/KOkCw3/FbmbZu
vct2ImYIP4OFKC7JMqE5wcxych6f
`protect end_protected
