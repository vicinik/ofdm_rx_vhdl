architecture Rtl of FftWrapper is
begin

end architecture;