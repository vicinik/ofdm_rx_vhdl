-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dqqPUt2mUC0FhBOCa5Df/aUdX6ej7ggpQwqTIjR/AreO8l5pTWUwVobMq8BVdVRle33wnYMj0bqy
gScAfySa79JBOnUUswyeAogqyLg5Wjrf7O1BG4hJe8XgyPIXEgiBKSt0pnY0lLs4naxmcvmNwHQl
nxxF/xRDh9yNaU/dqQCj5ljW/WrjBnDimQo5/54nSlbELw/3EcmwCXf74lk8KKRRKl33mRf5U7Ib
lz6zKBpOEMnssN5ZNST/6ZmgSWP3yw7SjhscqgJdXZfNosjT4NDnEYLgtqUU8PB9XfIL/HZcnnXe
Sj5p6jUw/SFsrJvM1uN2w8hkzhMegI13ckqwww==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
OcBm5J9RRL4dhuP4I5d1r0rf4Rh5FJyGljBaW2+VxdlgmZex7WIkSbZvMeHsjgy+zANNEvZ2lh29
F8Lb8S7xIXXA0J1XPXdATqqCk6JbjhIAfUt2C/PR6ARwGNlUXIzic1BClK/IRfAFJF6pw3edXyVv
vsCPYyozVVqNMJJVJj55y/bIXFjSDr7ZPP/cjOW/URutwznczTIdoJv8RT9TtYw5xjOpN7NTF+UT
phnXXTNUF5R1JDUgI1hpI312RHnh0p4LHy4louIUWwbplAaNdjdD9UiQt8f2w515XI6P2lbCfshZ
JDZkmp8MGQKmB1+xfqMZyDFanapZnDHq3puI5XecOE1iY9Xzhxl5+xFCw7LnIQ2pbPQgLEkBYLuN
ij6k1GIfCniLHax0Vdti7tGelQRobpQj58XKlu2x3fxDODZPhqJqYx1NE4afIKhfUzPcA0mPBr77
Fb4+5d6yUK132ZhnSn67je7oZ3SibSxqz5K+fTqneVk9fe9WfzYW/QN8pMQaBOUVb3i/0eOGZyDQ
5WnulRlWZzzURh6JvJ9xVKCherPGCj30j6KY/1YHgGAOIp8K634zRJBzZB6L6AfbkWYe9VHY5WVh
U1av2bltGY6NiKQ7jjnGzdrUWsi2prStWJvK+NcyIV6+y0zQLHDjgAEcgAx2GsOwjfbQmKKBnXp0
shXn6HvF8R1jTMD3dQnzg2JQqb3rAmznG04b6nU3l/hYJrxXAajw5vRuf0P1zH5u/JLjE5zjP6lE
l/Y3OU0dVpFMaMc4C2XFEBy/PFr3tAYSPWOG0Ozjp5YEf4dzic2LbZKgS1t5b7lSm7F2i/0il4iE
TsWn3AS5YbxeuNcuKxM2C9a9WiCq/vfHb6W/1ru6uthr6S8+pahAc34evSiNwrN1TeE9/xddyxfb
ANkWGb5n8+VZ6MEKqoDmQErdHLaklNCJMc1aRl8OI74L1frLzFXE7vqIVujktXSpj6thMjReMTcZ
yZaifefpOt3gwzulkOlF7uveb70ywVfYMAVIP+42EzsxqldYvDHJO/2hffMIC/chC0YMraNA2+Fd
GuF3mof8Hj4Tf/vxl272bIm1lWdwgrHjUluS7fGiGVlmxjCYA1OPBZPaX1tDrRBjdMMCuMGaQWcz
YuvOhbNaaJZk2Ug8Pe4i4R8MyaRcwBdsqu3skiiYvvyjnPLP93IQxlJNxRXaTt03KF5WSedYsn2l
nhPOMm1cabIyD89G71/sH8kCadTc2n7/UtJvK1VZpDKFCgMIReG2VCF0i9RsYai7RnUXAJ7H3BSU
EaNsa5myVMMuD+WDU0cpPnVJlZ6pW+42bMviLk+YVEMkQ8DUIZgQpnOw3fLDzlN/Oj0jVwmmX892
a9/8tzmm2aOPeds5DITaMFQJwSLRLzxmiQvKqoJbWEgMhxrhDrcwy6Pr9/ae21lcnfkNlRMO8Kla
wn72/w7IL/EG3zhKGqJfFlq3ndWSgrcyKSb3/jkFJPjiFQarem4q9N+qYi0eUICqCTGxhosbM0SQ
GmNr6t0PbaGU0dmrdETTp0ITZIZ7a+wMTKf+upQCWUdZYnlGuErvxi/ayovhE1gjLiPvl84Fsw1W
/soigNSh9XwuJjNo8DQh+ROLy8xTTBnAzgHjY2H/jxR9gbyRaAevJNAMbQ5K+LwjAEhUJV7ZtPtm
I6tEdDo0wxA9AVZNBrfzS/tA4tD8q5jdp/P93XX/RVRWJEhl0l9QIMb/zYnh6WUDB3TpSg7ZsPNp
0t5K7XyquZJZv2oGC23tb3IL5BLM2/tRH9Msbkh5LFMCiusOKqOY9g/yGnPUC8FGQjfsvaqqVF7t
YFbtmzo8MPIFbgR1bJAOF5M7/M5Emr4YW7BCNDar5Gml41rBlOja5U4wfanAR15E9ldW7i2UGZU3
3rNs3nXoPyRq7dIXuxvMsFHmJdZKl0+MM3Uya70QzUhn2N6iAtHYsU+rbb8TneRRTf+N48u3t4w5
v1lO7nR3q/0Sfu5im7HQdTRuV7k7P+tFFxBNenxsUyP5xTc6bHMTHRzXUzDZakECtWF4Onz1H+CU
qZjav5GRDTynogD4MD95qTe2d8Z0Z60fnMI/SyXu/Xq80y4HFJVegGbhybb6YrGCE6LLnLLObgrQ
jMURWVislOkSkP1+rwrRosm2nd9K9khzTSD21leAAj795NgA32AN5XO3Q4mktFKIqvgC7GrRcqqO
yHOYawOW2jYgda+mev10mmk4XMSojED/Ox8Wq87tNLe3eymQqRUcH6NpvDv67t+wraZoDlAXwDoh
dIE/hBNGm7+cxIqmbs8ntCCQz18hLZFfFIBpbt430w0JLQWI6NnJLPETIG07sp7ehXe6SAMTOuy3
WzblH39bHoMDjzT+rNDdzblT+xAKpj/dMia8O0ntzISZ5P4PJa7tOCHXr/LINE+wRKLkHn8n5Pdt
V5YyIwYN6X0D7kOYkSduLcM123Z0Toved2KeFfSpHpnZCzLhUTuWhmKPG1NFQiNYxNam1U5OxONy
Rrw6rLElLt/sfMr67RhhU+F3CdLArAHtFU83Ni8QANZhSqTXTNkgk1DAVS8RaqLDIwsZh8sg3kLO
+SIoyzQ1yNBueMO9tmubEZFYf3w41UfQc6cFsI1nGFGc/pgVD8er3nDUAROVus+kshqLYXyvTEyg
fjaxQLHwFgfRcd36rfNbHZNXSjLNJKZrUJvnMgPO257tw3rc4UOOR/D9Yszg1ue1X1LcvdCk0KVL
Lx4WrPrVdJG2KrvJQRVfA1gKu87LLwflC2q6+UzvFdtUcgMnOX8bsFeIeAc+pvKD0TLIX9spmCP/
FpZEiGOKEmDEmt1uo6psCNdrTIPAmJMEv7zfMUmF61o6yVTiMdhLlS3xRqbF1oZfwDvJhXrCHG4J
VlaUuDIUXNFghjLC6kJFjcRHnVS8vHnS++2g79oh7y81GqpAorU2+nlDlGCAZdFThTWX5L8lBDEz
kHAQ0dsDSHqSLg8cR+s2DFasdtnGErGHxtni8iqKEIYmnlRRsa3l7o1u9MA+JOXc6wBiY3+nFioo
Sumn0cqwyQLU9c2QNTCtRmnsj26jLUCUCynd8sruV46gRCCDh86w4vUPbUeLLh//3mbWv2pkxfye
QFsW5Ycwn38qUQIXwy4NgHTs6hRJJ8aKSFnrN7aCFrfZHWRNYJETLAqSot0dv51fAH/TX4C7K7jE
OpWfJwfzQvOXMJi1nuwlHtDNpXUtm7cVoHbWkhIL4R29E4PeaRgI4byDVdOCdnF8wa7jLJBn6cgv
YSm/U56XRVgClpOEaIV051VVO+jYATukzIFTELfeaXBsrzpgh/Pt1x+6qjO7JEfrCzKDmS2Ek+mf
27XHkysLRCcUoPCRkRi7vUqyzF6zqyCjKUf7yxQ0mrqrZ2poLp9OSlQN3Yggaw7gbauPscDFsnMC
SPyl+cNfd+I0CRrap4aB1JMCjZcAPbyssiHN9sIh6kuLN6LyljaiCEbNaWE3Z3hNJVj1445GQeJD
kt6wPqSy/ru/FGJyZWOIbDdUKxCmQ8iWSXPU2RXbRyOYZlMeXG/rSKbQiXktob1S64yds93Uhovm
zs1MpjtSkV0QZ0X/HWoevAUMtqhVVmnUKSGUyCK1xpdMx10L319/hhjHys/pFp9sDEGfRGRWiZZn
hReqH8gQxR1Q+BL7leoliN05WdSqEsH9/Yoj591UPZEtCC5ZQDxvtVGtBAFJ78pRLbR2JBKtH//6
Uva4UTRNFAd4epAG4v+upK8Fki0a6L73oDprZu6kTA/Nz4CJbau/+SP1UP+dkQg8NB/mMpt8imZW
6ojygM1W6ShjlAOuDFgs0Gb1fbzls+LGExPZf1HWp/dGNYHHZi84HNHT1AhwNYOhMlhbETa/xnse
YAMzkMq43zNaW082sPgJw+PhHMzKww1TvrTRWZV0xnvkd3J79Sjzqh4P7DUDdvjVr2+m0t3l+OkF
hzedz25LoNJ7rcQ3QvpZm+bWObOUjQaSILxnSwhe6QyZ5lJhn1vCQIqxUbPXTVpm5S2vZyvTcaGo
LwVBG/8MCI4B8iF45X1n1exdiloYEbdVaGJHZR6oGwjDCtcUj6i7eUVP7wzW+jXuF+jkcrvk469K
plAStgRSpd2bO+cgLIGvjD7bStE+ZZQLyyTuKGJVoakwoQPqXzADsfskhz4C5l2KmE9eyDVSzWSG
Xf1t6mp8lhiVjuvKLUtUZW391gdwQRiEe4G4PRGL1VRFZ0VnAMSmuVeS1TvjTpe4Vs7UYhblA3nY
px+KtnnIl6uRy5PyKlCdIgIwB8k+g5LXMJ1VMW8Q90h0GNYvogBhqfGeS4JiW4MaSnJHxZhBClBd
h69WP8/r9uwlzn2T+ngxK58C2zk1qzOHrbksW33uOE1CkRDzbfTwcTfXRxYNT/3tH+cJ9gRRv7cB
eStoxpcL8p8mFuXj8yXiyzvpS7p3JC3o4iuME/5nNESQCthkDZahjObI4SD76mhyBn+BCjt8XTzr
sMKJvel7SM0ZtNdjG5zdH5D9e21gLbIJOOW66CjYpkoKA+r313utP4uisRwSPgLdaCrYs8mRkaK1
gb01vdZa6w2EyvDJ4GhWrQ8kjivsNfBc6wqPO73DkwpgljbsiBToaUcQ4/DkBRldyGpgyZIXoWP5
Ovd+8jjjKjND81hSwIxZAwgV/U+AYr5uLWWdq13gxkmU5s1nxNF00oTvrc/VoNGxyOvbC1EkQHgM
wGMVZwJCQusX9UiynSTs41gY7LPmc9Uld/9yFceAfPD2pNuP1tuWZmxhv55acGPnzF+XLnP3VYw7
/2qZ2ABEfHiyRgrUk92oHsjJhhYQ/h8AzLXZEYPgppzBjun3HMiBulRb8GKdYwsfN/nowhSbaP08
A3gnrzQc/pPaVs4zRUGAFXVMZGXij7P825nLZYMd6Ppf1iI1Eobie8uiZzEiO8oVb+50s0qOCIgA
BWFT+YWpTysHm7IzbqdTmlv8bb1Ih0pUCax888eqCodzFGeCmdg3NHlNZex51tfc8clEKLt/jtyq
XYJK9wO3MnhVrK+mLzr/ZJLz0tNRwnGOCNk+TE1Avf2XdrHdiaxZqhHOob8iIy52PU69B8Umhlbo
Gb44ep61N2yHBPLhtqKuU09gjdJVo/yRIgRJOvO/KOKXOMUAn2d8KxJFanv0vY+agsMf1eXiN6jh
VznJ2teSt80eGk4O/ZnxYAnA2uGHHsTEAtnTS9vfQe3PF86sxjn3Dtsbu3hOjWDUClPJ+9COBXXJ
wKD8xLUEvArmhpzLd41/iH55xm5qNWR/MtX+Qanaote4v2YSzxyMehJZpCe9Vp78zxaG6wFwiLIU
EQ2igYeoTNTgzZ4Dc292yv0LXG1qQpyLzUIRR0GTXuP78b91NT0fkHhfMqAAo//0iBZuNgYJ+nQ5
bv8F/omaY7uoF5WBtSmbJ6Jpe4tZJuw+qez4rACfV473058meNL7M6a7VFPL//xyypG03aXq2xHb
MILEsA2Mx4SwneUkdjIMMb5K7ntb/AKVTKNrD1UTdWU1DB75ijQjYb0TwDHV5gB+y5ApNxqd1uK0
1J1z96KQR7N7938SMBrsQRH+pUZ1Wfon9q6VpA0zW0929/OVndLY9Crxsc1yaekoM6paf7rKv1fF
hFY85wB3Q5dgbgfcEOxge3oQjQFLnXbJirQo/S1YaRbSRA847zaDMBkv/7Dra5rLf1k5blV5P5nn
6Y2/mkNk4gO/P8Uiw+ANzEilas4aQtkTcaQ6d+ujGMJrgwERKh7ChQ6TBPXXj3/pRUvijIVFCnQM
YiBICGkSRDpD8tPjFvDaIBY/xqyDng5N4XF+MzbwXawEKNZZXaqOiUVdQBqCvRHzs9sFb0Fd1pVi
QgPMc3TNogAwyd5TcTjyK39UT6sJi7yWlV1DeggSc3q1OfujHx9GScC1uWKVBiiBtDhbqX6HJ5OE
pTIb8PXog5F2abmvA5t9sBznBwgjxoHyFNO/Hx3V7en9tUL6ZA00CoqrGO8/u9NxgH8h4ZLkTWyB
pz3UAu7gH1iNAFoCIck7YIrRgtvXTbJkmD1XYWBJV8Y61rD1439wtZ7DiaEXlDwS/GKZr0DhSsnw
rprVAgzR9eXCUrVWvHhFKQivItRTK8h1sStV7bwweCdovFlQJqMFpKjs8E+b95Y8Irsdy8UeefOu
jak/phW2FHKJG2sbzElj9BlFBjjwbQ4HPTqvlTg7yXU/nbnxok7eNXAaUQayLQDCZmGP/YfNhORy
7lpTpRyztVqqa2U3DsqrjbAgm5h+cjXlveW3hQhb1iEdZ3xCPGxEGsDdC43+DbnbincT25cDU00w
6LJAnkYaurxcdzlJaPB/mYM0MoGXYPb/ce7MWZbjNU9SufC5ZgjbXuBqOfAR6TGRmupWqmyeNeY3
l2ln9+ZkDE9QE4mGuAsDPC4VxtdzSco219hlcCdDSiwLKiinPN/1h65n3ptM4UQvwQP/lNwULBqG
FkkQsNJbsgZiOslLlVyw1sT9XrG9YNhSqoQ2LzxYY4zUpFr4msCm/pOWMKbtcUxcKjrLytAS9AwI
r3KKN7xIfFl6jEoRhuW1a9mfrAQQIMS8wpn/W5yBk9E2ttaZdIx9Qa5k/umbqN1kwS3+5NwuS47f
EUuEOTQRECzLJ6F/kILaGXYSCFOxbj8mcgBwk7Kmcn+MN40aR9pxqr68uP5Kw9r2Y3WGggcmwhFP
zwF3N4KJwb0lwJOVKmEb3saoMkxe3WftfZmjHhgDwEMcbkCNOWdbqkGamb+uf/RlyCACLPl1bual
Cg9nf0jiIl6BC2R7IqcALklM/S9ck8Wm0dQ5qg8yEHFk0cK9TS9gxd3g003/CmWB8loh1gTHE7J7
76YR8rcPyNmWeptVZuZ6xfyT5cE0HpRCVTCiXN1by0GznCwomqp6qgzZvWvBLL7uQE0eupHGp9yA
2sy5T6qUKAKB2UmG0XAGTkCm4qZkTKQTNqipxNalRU1rreAEqAYpR6WIxPe9gPc6oQgFZuP5CClO
AxG+ZXiTO8CfkMJLHv329vjweZiLrIpftiP8Pg/nCVCWIeySU6RCmZ/KQzNF7rNd7cIkDHMbOFuv
q45nxpi1V7DOilNMmMh69UbGCKuh3nxQmokPkOeUkQwhyaypgKp2gwX3+oZKRrL74c9KwObUSQOy
iK4C5PzHloSK4vuHKKTKXi0ehlNntFaURGMnuKThS2Rr0CXHBz53qrxzDPj1ltk8WPTRbN9bBznw
REULjEB1HgbTFgKRDo7XlzXp5l/5JKTfIAMsjrcfwo2XDwFxR0pTsprfn3FGFY1ph2RBfUn4GVGw
psE8IsxfirSuitYpVhUT+DpiLMeCELCfW4OzPzeKFEnyNM4iBYQ6VQpbdS9npQfkd2Hejyfi7I6a
JSTg9Le4rusnxh1LnddQLeY2SUMgqgh/JUeJx2SrSBm/qSU0OeP7O49E5TgUmhjIl3Yx4J5UH8b5
gQRQsScdFZ/10fyA8jWYiiw+5NoE4VckhDT/Ra2P6JRjH/aFRj3jjyKl1ux2dQyAUhDKSVn9+FiW
LNhGpVp0BW8blYUKT3eju205s9P9czHgLHK2keVmfWeG91ew6pm/LOiLtCb1PDzuhNnhRc3rwKZ2
yJcZVf10W/bbCZS1BsiF4UG180V3vHI2WnC9ec9AiIGffTKmPXwVRWzJqQnYHNrFFMPNYDU0r/QS
H3KcrLr3EIKxqmJFAKN0E6Tp9V2fg9WotY3JWBYzmEnePoGWoRE5Cduplr5XhDaeMVpgAy2Xika9
g8eAfxL6dS1o+LEj+3erWQzvLPokDR8bnOGAt8EOubvX3ldRUwisYrXaca/ygadbQEgbU8wXjEdz
axvyQ4qU/SH/4XHqlqiUncKnTy9g9FHk+IRJUYVqr4Lu0sRTUzmoTscm/oY40gx1TZze129eOnED
xqJyW/g/a8uolDDk2YyX3yRZ1YeHy2N+7I9MzlW1mBO1G+deMIrwDCwDR9GVQXVyErkdAhWc8xga
L9vIckpBeacjG3/tHb6VNbtA3MWi92PBo5bmtF8PFlS1LIrKKDMlf4J1Y91ehoZ0o3baBPsPAdgS
0hHW20idpCndmdbWaUgAc0MMM3LxjIzRfW7nyujUDuNwbqTxal7sYBdIdkOOncf3Ss3qFSAzAdHr
Kcbe+ORFK/hsgM9Basa+SAMpAA6gSQbYLcosoOuTRaIEsVZjZemkek0iPlK0f6VVZnBiNn9h86nE
O2CFJXscrpIxEhm8tMxh1LtwwCiHvVZdlLrGrx4UoswpPmaWC7Y6LjxmUFhEWiW/e0KkyzyJZo2M
8hQVSakHrGXiyErRjoJxW6RW/KdLAebv39M4oshKvlK4swRtWzMjjVtMFjz4aZgHQDCmg/RWboHy
NSn0Gh65bOYNt2/ButNp9WrB1djWlsroNrHcYB8h/nolgvOG0vbq07O2yUWCiXjMuD3NpnVYtW/G
KtQImxhOY3YxgLt66PKR3eZjbxUpiF13OrQ9pkMdkrg3n4sm0Mut99udHyHjGlWOKWiZfmhnjmgj
LGAshdu6LNss7cF9TnP+ojJWVFeVbQ//QwaH/qtBco87kYpWgPNWis4ubmRBIZ6JtH3Fw2DRpdBQ
6dPRe0pj9PFaiTI6RPLvxABZOHNLIFNBFaylKafkkp6wgYlukUc+PEFvX6YymHw6IPShziG6Fnin
DV6IjrkHcsuDFCFH2LTDYh26T/EQUeVy+MgyPCRjxIvITR/fJRWuOXRmA3zuTdrTtahcEXILq7z2
GxB5GZLPol7ATeUPNVMYYembebLZCrOCu8q0gRKaFfHd/pYdrPFsjZFefcTcxQ7U5GnwKr0h2vuQ
uHlsFPtHCx5bDOgTPYeFkfcATx91F1sbcYPDPn6zWYheJj5e8DNDVrNzQdkiNUPA8PluLrQctkOL
v6vn8flAH37qklIHMvFRQd0BL7AJgk7DdjT8dMH0hjAOYHPi/tlRLm78tc28yhJyHdcwdP+xI+Aw
Empbo4oqHKKmxzqaNhiAWLvqVg5bfwBbpGejgZwn8O+k2gRP7Xewu8vu2W+tq+MM+u2oXcjod9Dy
HZSbOCOS/8or2H9IS08Jhv/0356VvEaVAf43tB3pav0S3b3ctCp/+KQgFNfwlpaIdgAwOOi/M4P2
3P7JX+gzEucxbb46Aa17zGmN3QUYXpb/1q5yd8tCgTP1xYf0RaeHu8gA6fhYQcXLWcSa0Srbajhr
WiUoSJ+Z8g44QwnWpRfkWkxLpE4+AyCm/7/bigmgICbg+uBY57UvSQQtybi/E4aZNAXrzgbYI2Il
iPMv1IwG3FX1u2UPWIS0KY9fr+GVmfVpDuT7DTZjUNZmwyIFLRVlrG0TRctWpGjCjTRPT0RDle8y
XJLNdBLYNFL7ESq/zwEjhxPwctmCqK68o8+LWwPRstkTuXeXK4lC/KHdc7bhsiGtCcQiJQFDxnGZ
3ONRK1O9xOdZZxVxSGKneFuq4PqJd7W7a4HwiJ0vm4DYmM7/uXsPkG7mlEzrlX3dItH7N6RyiRj+
/PFf0zDJ01th1K213t16dyrgeRnZxi3CW5FduZykKRk7P/UZAocbOFw+fpiZNW6xxIUuqNu60VtU
qaHk/hQqe5VzzAHiHPTRFZlfw5JOw98cYZnb5MGvMEhpp5QX11Cmy0qhNvHrBjJAxlrh2fgkmL+c
TlGb24cWonq+tOtAkAzU05irXizS5d/FaJ5OvZuEuUkphDGeTW3CsghfOVnGNcOWUnaoRETRKzNg
ht/XlSpN6jMiLjg3uH3x93wRbO8xLc8E+1Ugj+t02TbXrCjGbJH3cZmyLaBV1v3hXg5cYzk1lhrp
lwkEYRuFDJrQr9j86Svc5hfW22u9r014i+xalnUaksyieSZ79vbO78qksyHl2ycAYMrgGa+jy6Ag
eQg2ZxCy+q5HkCNhPZqe+BrXuoKF2CD1GAZwEfAjGqNNhfKrn2DGzzYM5pzMNjgbauruj4UeJbUb
0FGTenKGFoqyP/DHxPK8Gsx00ZAWnQ69IvWrU9F0a7eyupzFqKCfJwDQoY4cVoNc/KK5sGvAh7I3
SK97K11nAKzBKIoCM+bIR6KfaJA8WvnUNn8VjExqyGqE024JNbY7C3TtrxbIhwZCcTlAwqDZlLpl
8TG9ITuOldVF0qv4aCAb9sYaliAqL442+khrgXT6xaJLhodgwq47khhBXarww6uEw86bVqqdhSnH
qVhmw5TmmarTsTwzJEjTYNyliX4uaBywS2zoIb9bwquxyARLj9J6dR9j1gDkTnumRhCdEzEZhp9m
Mz0iX8He/TEmkw+6OLv6D2m163c6wpXcmPnGAidA7RkNFHJCbXX3DcXgl7h4bhXlKRrMn/rs1YaC
dGImlcYl6MxxlmqgkrKAXOPZEoxuHwZblJUdlYrcPhb7K8irgMVusdgurYc2HaAJWULcp3Dk9lSQ
VghiYcnH1V98PD0N9fT4haHWl6kC2gqOr9DEjWTNQFhWSlAnkZ83c+a6tEdrnMz0UXbQNuRU/IkI
IqQ8MUJScBlmNGJVCAOh7AsY5b8om7SYu2pW2AFVUd4tL33ygfIeWL4T0xN27oZMvwpGHqWf3ONl
m6CBJUWonS8nwf/hc9M8t5+CoMgRYCoCjaifXDf/jfFIc2neRPLNbUfQtD7RlEIie7C7dUB01l0q
AqbPyfw+sN9O9IrzIfKhIsLoJguMbuxAU4YCN+o7Z6f+zvlZa44sqFbfpZ9gG/JNhJjFdItJLLyE
3no3sSFt9hhUEro4Jh64XCRNqfa3khuPfnnY6caCF09H1jG9EFmu0HSRZJjMcxQ5YN7BbHBNpkON
f1usYR0WRLL+SztTD8WhUrucqI2ZUeSciQVhPgZVwpNAfE5mRqru7nufdiDuwy12r/VyCa9drhKx
8s/jOH1/X0SCZGMozCCkkaIMkFK46W+iZmnTvWuyqg8FmYJGb9nokvf65wGHUUTzqfKOCrzvkF15
W2bMNGh0XonrYARoRRFSdpNX/Z6hIWLUJm8ph+OMVF5h7T5hXSESB4CVjcKrGOJ3nlF3pXST5Vyt
b2yTgJyB4AvxUVV9n1Mb/LuVGzr7yb3z2vzFtCfU3Y1Olq0oy5Qwi2F/5ZsDxTTcIJ0XxfSR1051
757EfxWm+crEnSHNggoeizahPpL1SDWBhgLq0qNL26KxmR526ShWw+1oa9yDT+HOUiJm0n+YctkP
cQeotpDf1+whbu2C+912rFmHn77mumi7gCpXo9Tlwnun1j9CLc5u2ZmfvLjA9JRb2IMich3GPr0d
73NpWh4PsPgWEhqWyTdAto2bsJA7GESIXRLVa54TWkOWwZ0UqPktRNQH1Yi6+b1HZ06k4Da46AMv
hYQ1MRsr1FMmqr1Flo5WRFr2yvp7ASEXmJznyLObNmEz40RdYfyPikvWx30wjMbqcyF5gIFUza7t
xZjj6/UQuBOqo3jEpl4R/+XHdkJIT5Xntzfy4s/yrWny1L2wHUE8JeLmhHm5kcWBEl00DGoDXbin
tDcpCnb8iV/OX2bSa+rFu9+KIv6qXJXiHz3HqopFpNIy2RMRbpREZ+Gr/KyFIdAWjpZ8EStqSEbh
4AdZYTylZpm+I6gb4F5mQWoFAOKvuN0rI6MQfQPxMbO8spE4ZvIh7IIci9Zo6KLMqKb/Xk6RIFYw
ks2EpJocXdibuk2vfjivcj5EZDJJ8PHOZxlAB3xjgHTcdZYGITjCLLFigznS67YnuGaMJMUSl47j
PfIb/aK9Uk4jmJ/BCWTX4acTf17p36pexylkjuowWTMZsxHA5lYJpOdiIoF/zzkwDn8clQjgVZuG
Djo/9xNpymc5EWu35Ni3q2+GwGpy4leJjdkuiw/fbMHZwGoEP9Ag+3IMIIgK+8a7Y4iUp9AVC8Ag
pZd5B8Vma/XpcMcmqeVbdc1IzySF6Uu7J39WeIrBro5saruwX/8k3uiG6KozpAvoRJx1IHsq1cR7
CmNa2kmi930Pyv4SsaoedIaZ7CGM0ELIS+LEYYNmR0N5YSkpPm39QIPrifypZA+5qKv7h05i/Ch9
k/Q1i/mJMk7erdlTFrsBY3aZ+IlDvzRrJVeeU2rTBah8sfQQVmJxUke4ZMIzXN6ZKrau+axgzoyO
P+Y80aKWSdaLVJikYmSy90yBpZwa1Fii9JdTGNAF7oBrQ7w04sDdvLEdV9PgU7KHqel30+E+34wM
RT1pXugOmtQZW8m7qeVTk7c33Z7lMCsQOGgBrQ4YbPuJCf4Y/MvWjWy7NmLDqG7wx6BZEkqz1kAv
o2wH7HTHfIJnjEkKBxi4MgxzEoaSjS/a/bh2qwHL7Ia7gn1tryQPej5hbInYevduJg3sFejOqo1C
D1Kypb88CFdJjOUXjis+Aj2diBu5VRG6Qgg4k7RWpa9l3+s23De0IkHRhZ07WXjN0MYwbtBDVtxJ
HW6T95/6dj7TKIYK6i5gxDyDVboWGtEYQAtbS7mwcllOi+E27USkYN9MuXg2N3/hBZMfsJ/3tTF4
Ubf+2PEETQTtrkXBwtWAeAvjTlOcfubCz1AbtQ8Z2RdHlW+4b3BvV80/Wqy9ZvQLxbzqfDjJlxQG
u/LeJJw0OkjPnAh4yalra2CK0aVPLJfaq2tUkgPjtXeErq9HIPFQDoNEHdPJBGCWd9WIXzzNZFkW
+hyHtw3rwGSjdLLE1Ng8g/JF3OT4MKXNwfk4nmmYYpH/0IioCY4NU78fd+r+WZslkG4vSZM6g9hC
+jY4j/ajIZnAJK18uSY7r/Qrr8fMxBqN+KSTh9zepfTdWMrTlWmYppK6I0KziFu4dtKCP6rA72l1
nw2wMTFEoszgG5J86WvUaX45b9er7iQ355FiJOt9JVvF2PpQvN7EozF/m0M/IKytQ8BwIAxjVn28
mom/gbc10s8ApQ5HUk/KMgTCwI6mgUN8Lt6gKZVorwsXQH65aVoFzBU8WWm+H0uJoART3xQmlN91
unXT4wPkFoHkwfA4ZAgzsUQpntc0RoOY/9LVUcWILBKYcPGoTi2pZ3pNi38opleqz2VRdbkmy0Gp
A2WVYqYPvOKMqstI9bObjfIoJed1IkA7AZMWC3NZqZ0EZwAovvUpuXALumHLvQaAwdgPWCxAC6D0
jDP4y/u5O9lyG6BP0sqffhLLEVfkpYLnjrghWuujebTBp/FHFTW1A3UtXpvcekmIoZIPtoGssJ+Y
XjERV6WlVitbw4AhW2hK91Jes/NT2VfrF7ab76ZeOhs+BX2/ULsJyGvFfhlDqjd9w6y9XH9o+lBv
rMVSy5WJvO9tUKmvgN2MkGJSIVavDIMIhiB+gjRi85EelFC5HdWOT1wzEzkezfTdVX5FNUB/lh0I
57B/h+g52N0UN1O0sMOlykQnnD5dVgiTHYCKWHNLAY3Oa0ddwR/rfRzUg7Yap8Xw/zarozHnerF0
Bq/7nH4dv8UoWkxAq3BxSiKzblL1u/9SSMJhhXiXjwwaGBJyUSz6JyKUwrFQhydQCG8pLHDM1vF1
kr4mDH8jv1aGF6/sL1HdMIsDqn9MUCZhoMGgp0ZagaeX/8I7ePlK83XTAwz6w52S6Vom6dBdgZ/C
WUSJOZDYxKE+33nz5SihLw2RO/uBeqa8rrPD+mjUXjILQpqRZas+ryTWKTHNRTK4fctlSi7EgG4O
4hNfWJkInd8V+LfpAquhS3Pl000cZ58/6zuDD1H2inHoTB+dseS3n3YcfFZ3Eg79UNTM7/CztpDC
FnbeDfcX6pIvOOlgoHExTBVrAImH0N19v1MIFXQzowvECdNmrRFVNWN9xoNDlurqSPWdEESqVA2n
2CfB2l2U+u+q5T6RtKGURDDxOqvlMi4f9ujUZjs5fijX/4EmtX1w2aWj9htfbdjt/DTHB6oSXpx1
k6Vl8l/jRp7WDW9aoaYSqvgPlw7FB/PzWFlqPe/N+Lm5cf1gNj3am9tDlisW+xGhAe2LwA2AIJGE
VJGpp8GqSDR71jCTVInWe8undBh/61/au+DwjvxT+zPxM8UbiCqpv/CxiXqK8zG8oYmcTPVyTuto
hW+dlfLOWnDb682qm9r3MHNvLrr0qYkHh307B6u19/Y4aos2ci3vpdm4oIk86os+GcEgPFxq4HDe
SIcR/ZvW3GLPqQrC22oSYA0aemwk8uPFOx6c8og9QbOGiTVFx/MDiiMdj/KQiss=
`protect end_protected
