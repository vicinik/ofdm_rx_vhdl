��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P���S����b��G�=i7_	�/Vb�f�AT�`K\��rߙl�*���Fc���3�x��ۤ��#��:]����߀��X��
�S�G��P�UU���^�ɧ"v�CT7xo-=���	j�C��k��Α��Xn�Z{��Ó���d��G묟����A<��b�)S)@�~��nXqZ�Y���E8�� 8�)Vr��n���O&]�4)d��l`�mmX�E��e-��[�l
���kg�ə�}��Vto���kZ��2��کRؕ7�x5���5��1C[�u���������x~�E��J"D����^��;�:��ǵ�]/P,Pf]z�F�.�x2p3��JjUi��EH�LOK�`1�3�vXތe�G(3�M%�0QE!��Ԩ#�M8�uV$-4et����4�h,:浯��3�a�z���^@ �*�0G�Z5��!�?ڠ(�Wn���א�[�>?Se�8%|Fj��j��5F�U�70/M�T�F'���q� t�0���-�2]#}p�0�le�;�
��,��
U��9t=�q��9�i	��?�]!8�iM����J� 1�R0��AJ ��#E���!y6%>y��Lo�=�t4	�]��(�[P,9x=�ҎV�X<=��\�$�#���SFFU]d�u(��m���8�~����u���{w1��ʿ��l��y�)Wv�3�e9��8���:M\#���f�6� �����/���y����mG�.w��}�X'��l�ۖq����!u�v#��s_������
�dX�^r	9a-CU��������}��f�u��|~��yyָB��mߟ�Gl[?��9���K�a&�\*\�I���N0��A������Y5��i[\8�H`�NS���@�(��1RD��S"����^�0'b-����� �M�<�A`��R^�֋0tŷ�
��e�WZ9*��~��[�/C��`Q=��1��y�Å!��A��#����߸�y���''#u�P��}���|~��ۤ�/,d���G*���W�R0�̽E�9I��C�v��o�8�)@&0�?�V�^L�:����9(�^����ʍB£H��I�ŕ~����x�lx���4[]�Ǧ��:.�.z$���dG$No�����ҩ���V��:�W��r��=��}6)��	zI�Q����+lH\ym���(�p]�%��#��q�"qO�{��ogyʿ�v��j�#���>�Ԇ�Wވ/