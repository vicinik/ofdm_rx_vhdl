-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HpdlIWTODPk7UM8VWvOQI436nPOjCBlpwCxG46Z9n1AmmFOdbeYD+tY0jSTq+Ak6+RVLWEWFYAmS
ZLHvMpnD8nn81OfwY/cBMJ3UgIHxS1r+9J1h9hqktNBNsYS37lMLshh9CC5nawU3X9CGXj+WTH/A
ZzDP7SsPl3lNpXaSpmx+6VwxB6pBEaIWLdScU4b8FdMmOe/jNIe4RijJ5Rmi43CT75ymJRNfq7kk
I4VygQOUCggqw9AlbAm0AOOIVDnhwLAYYQuvPllnLaaLRj1ibcBdy7pDsnEKAaPGlAXDlIP6HRcI
I3VsmWmx8dHPXLdA4LXodMLPnMx/CHY3xfg3Nw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 72832)
`protect data_block
Ozvn4kWOu3xpiF/RY+YheC+CnBX4Dj5btSX5ubZKgb6sUjv2stYF6NEnsSZLDw6syDf+YKZ5JcAT
uzxiChIqozCz3LfQxn9ckBm9f5BSGvsq+kKs+JLKcGftHx72KmspIu2lQhTVEmbiGpaM/WZvar94
UZUidwbKkdiSJJhnnlOYGOGDh6EbzCrPlEth4PTz5vaeiNR+MfCkTayitquNgX1a5TEDFMh59RCL
Zu3x4L1Ft1/DVrkgoF+VtCC0+loOpYPVofSwWnA2KbJLgmlGbwgACYnH8xuO2QQRrE25FgcMWstD
72Or/mD98Ok16rTJI/E9z3GSA7g/aa45jXREUTHu4JBvHq3Ltoej/FPVXaD4nkYj2xWJJGlhEfKE
G1EsRWjD783/Np6OCcLVxnm1qi4bGfpTGK0/S/qvl4Cb0hF+T0Nj5oPGBlfy0MO5aQqOWn5LXGpV
J2TpNT+JxiOHRhfD7LofFnwRzJ9yEwF5krjK5tbY23A7ZoKqcGqOjsSVxSX23L49HYF61ITW5mi5
weXfEM+QSEyAGgFyokSrsKiikbvPv2LAswXc6kAhQ2K7a9FT1AGekIEkFEY4LPgXVtSlhXbi0LLd
R/Ng9UK/44hW91HmtktcqT2xJRYeATwO/0RbT5fic5F7gjuZsHhMCZv/E0xmKnEiLoL8vbpqO46L
8+qvcAfiUALREMErM1mElN2XM6f8XsZELrI1drux4dkkpri3piOL96nZ9TRW7T691QYzV4mwZW6v
OAezMa8Wi1ec4fw1w573TBjtN4En3lJBkQ7tIStlFeF9RLMQMjeZyT/JlwaaXYC3gDd5znLqhNcg
ZRKrg5T7geo8FQNIgd6ZcOBBeZ4qK/hGTKdYSUREcAUyv6HsfsWPB57JNHtGjkV5Jv2JTLYUKxvx
YRfJmXI/EGHOFgAfJ1PyahyQ8/JoTyFTKYCbD/sVPVWh5c+YL9kwTFbCmHQiL9q0RgqulF262gj7
U7jr8GRQMufgoIw0iDBrna/jhPwRINOZQtPpHc8AvQLwHUU4xAi+7CIvimxaz1bSHv1A8+T/Df2/
CQ0xUUhDmFWlKiwcUtDoUueNR094pCyeHXx5tDMlxLSM2OwsaHYNyVW+pq/zK7+DyeZ1RUI7Hy/c
TATP/1o4ryv8tkQOLtNWv2uXzXkcgXFkmrdfwi6UBuYvfAwhx4lASirkm6lbzxakwP9lMczEe7zL
yzbAIbfAghLp/bifDaFG7+wqQd10NBNp3qwZUoZ8saofhO1107Q1IR7kPbv9Rt0Lh7FWxtEF7fth
QlON7YwfgbCa8RlQ6aVDX3Do/1XzpDTIIN8tmhKdYyiQ9rL+nF/MmUWrt4Fx1HsPJeQmTYWm8pMX
JggUw5gNmMm6CwguBECRyvgNqPz15TztVY1A3sQ5zoypYsS7HEARo8nKhD+VqFOL/coRIClDoYJP
W32Riofb82YG/RcDntb03+Ar8WKn4UuCrXDCtQCqJhNCBh/nbbYf3IeP8wkExdf5H7/juDPYdvba
3STDXdR/wExB6dWBoPa8ftMKf9CYwYEhlUKVzjiXuevbLijt4ZQWR5Ev6AfdRZiHtQQwNW5CPRqO
0/NPcOisbGmea/6BUaHU6NrKzaeOWtZK40d5HN31ORD566RFNloI6PQuy3ZUrzuXvCVhIQ5Ozp4X
IvCbIbp/Eloy7c80CHyz25uItFHLPiiDpRMbrhJzrZeQ1JCqUNMZCUQ/0qwIXhtwzWTaHT7ssx3U
ISMNakgEDwvx7wJk2pNH+VwtJn25+syVPWogU8PnE/t8jWXcmiItvfIsj/XYVBC+ZNNR01sU/60g
Glqw0LLBwKmBKiU68hYdwEGxNmQYSQAJiUDPTpOqdIWbxKbX9TeQMdZoE1aVoOcKQxReXbXFaTo4
dRrKVvULmqa6uXetMfv9NoVBpLvFHTUW+eBxKCaATncv0ZTWXDtSRjjpwTxtgRa8yBSDpIKoyx+n
KUyTIsYuMUc+3uVc35RaC0UFhqX5WaK8eEDcd7M9zUHoecdnwhc6NKgQugYvrWc4wM//YkTDwEmp
3+0UP6TmK4fF1wOUaYFR5dyooskF7VAYaBuhnzR0Hnptpv7cyn4G/rCY3njnELphhyqpYHJKSFcj
9Vcwzk3aLIpFN2lT6Hzt/AhrAklIDkqUSf1NohfT73OaeoZDBPfB6zpx2n41DV8FnRERuwHnrg+I
57Cs4IhKXfbd4pdXsqIuhoVDXMnfWssCFRlljkKEcjRLlaXFiBdrv7pPTHmH5ifMJxwZpY6gig10
ImC667LTXk7/B52IZrwJHo7dUZ7l22PRc0QRlbU2VJHz44a2yFB+Oy9HkOeoJKGZqpJsze6C2Hti
QwHuMEJwvPLMWkvKt2rx+D2fp0O+KIUTmgVdtGeiKZEcmAiDH9be+79A3lzbklm6rac6j8iek9tF
YyNnwtY32RSI6aqGrMehC07dUJ5kCSuas9eYjUzdrj5RHBDdHBkgfFNPOiAbynqbSfRD298Xi41N
cm12DLSRHdi4bkePjVZmsQH/YziPhtt1VxTxns6aKQvAMch3/2gSh38jMKqEaCc89Fg4zWQoTwcE
fggtjy1xD1IDaA8XHmbQyqZjtLUoLZIJSwFg3oSZTfy7B9ldMqd8qjVsVBol/U2BqSWiu/2GFVKW
BuCIMpnbhBrG16OJYguPE2tAlLTfN4AAuLZA0FPJTD1iHGLxnBISGAuBaBgS7M/mwrCZujLo1Rr4
xRFmCqOJfF/WRctLgWPbccxk4l1gfLgo/JZypb40cHY6c1PAOyYPgb0abtPPpPjecWnY3zkAJaG4
b+JbcMZZPrHY69lOJGNmOY4YcrYjV9yv75Wbx/vjehmcS8hlsMVVvkvhqQKCCb5W+scjMd05QM+S
KaEoplTXs55iSH+bQg8mh2Me4C7R1taIiArIipydtSNZMJ1ZPfbKli4EFYN+Hpe83FO2aZ9lyxOp
uLqMYPqJvu+E+FEqmPkIHpwKr+d1M/V14aslmfhIMQdsaV2PRIiL+boC8Pwp17e/UFeo7M9fE+t4
7jXb3UrotcO8FJs12r6FBV75bTR4x2j4i3RJjNdZCfC3Z2FXrfwSRY01j2TrgQnndrjQfzuPeJNP
7w8+9HdWlaBuIpkHfagnbzLUA7MqkH/r3eYrvphPl9Lqj78ujy0xZN30viKvEu0v0J1hwXs8GzYm
IwX1HrRrEGBdopEjZrvlQnVRnOQaCI9yYXUs4AWm2N6W1hjKhfalXi2RGQ6/fHkoAWExgiqhWZ9W
yOt6H+RHpt8LlJJa2IfSCSMiylbjKDkRSTl9MkateWkogX/OeS4FFNNv4cmDfE93pNjsm3DUGrYd
FRy7dYXbDOBh5A//T80fJ5ffaZuMcz8hOQ3F0+QlQ0KRB+uY5oXWVg7b2gWKfgV5IwknpTDwZQSS
wIG9sfsCnQJ7Xbhqatp0fu015U/Dj9JoEs5gKlJ3j6TSGxEpGsZdvlwIUo063bZtavPhVk7FCSzP
qyb4unT2nAoA198791+dTPZ3DH5CrYOWa6eIahHCSA81gwTDVyHSHNCbi4DTIeFJ/3FPl1QRtqRh
u9e6bwCwBmbZhVoQ6jTSkYBwLQwlsI3QPeIcWAH4CUiL4ALxA28LhGedbQsFAQstZlUnv1/mIizx
xMTPGz9dU2Z4G+Syq1LCy/v5YDjUkVuzlXpeqxqLGl8js9qQAZiNHNoED+KC8ZabwSPfh5zBgOE+
gL3HxTNewwhZCL21vpMoxhA9OavPO2D1R+Hg6nt1hCF4EIg7JANUiB+YgmTlqk5eHdO7x4nJB4Fd
J8w36uWibg3ZiVGZ2ga9TqEoEIAHpBgPPueBGsp6joBEF2IQQr/LoWXK2krHVVND1WGkiKO7coDD
k7Jkf3gXJKv7KoYA8EO7Vla37gtnPWe0Vgf+1VESV6tFZCD9MSz2qT/1kbkzN/BVzD2EnUqsZGpz
f7JuWzwqrxPDRlsuOxs+VJtoJA21Fbmk4zOBpMTxOU7qlg86LKQEXix59/KzCZ/SGY+TQc1NLqub
0INm/i/rOz57ZCrj0KtsaiX47yX0LhuZYT5KFnFtA530M1sKjyVB5JbMyHA5JV8gzzPwvIDahocm
3XqNkFcKvkZvNw4e7C7y1WSGVwvR2mNmpWzDZdiw2oatOh4U/QwV+h2sPIybmU3s/oUYuk7R1Q8/
1NAqMd8y6mx23b3RIFI51M6M6siP/mV7eGTohkbeNejGudeiaH4DkeiEicZRi7lOKXycTHPOqaMT
lekt6OD5Dt0t4Fe8j9gyTJuAXUmKPAQbzUE4CTYCmo5iVU4qRzgiQGUvATPaQi2cccGSNTOqSUeb
75rjrk72YRzALblAtN1NeO7pxBkXLwUKF9Tqzed75xe4CkxC3D1cOkCU0og9JXFmprAgIPHLDQ7c
yQsjXOZ83teGUMhpeW5a+65yBMS/ocKWGia5irg/2PwRDClvASIHBoUUj9kojaoeKJy96LjnMKUx
tzDrSJzf49RgRSmYwo58g3DSDV2PE6xtjRlXXHvmeEqhR80z8qFf2gaWl2DwPTLKLM9JsMGXFUSv
FZwlwBHYO9FyAINYfYMtg9XMQXbqOPqNTBqF4jyKyEwUIqyZDs+boIxtIH2xvCdW3WOq2p9BagBn
8LPLpwQMEaKra0CT1PJnRyDwZbY+WapRne9N/nnp5dsHgPp6PISfgbzGAsL89cxmkm71IfY3Unol
x3gJVSGyvelOgFVrUpcDgIzNEHiysuiY4x0iUtYI0sBm5rCY3oUzoXv0GuevEEL5CjZpY8Axipo7
N1YZmVUfjf1FaMJggiv5FKpidlnGRZSkByHhA2GAPRBtwPBtw7CLhElHh9VCWzX18pY/rUVvn1Sz
CPor8iXNeNnkiIT4nP4AzlMjSZK+OXtUZ70cGdoyjHlOsDVIRPl9K34OJOTbx2UuPnlt+A7mQdZW
6Y1xxc9QojHONzcGvIfWefpFUVzQT7knf89xBjMd5VUeuxYo4R1igFDbpMaslLrpRjwzLR1dzoVx
28krdXMGorkWy1FxOQoitlQbc/+FFY+D76tyzwU7AOsKcBz3bjudWD6mhQBFcKXvHqVJnGOLl4eJ
qiIMONxVVeIYUpa8R+p9QH089rE5KEtV52EFmDirLBGUc8fYdO5ub/o3l8b6gMEUWe3CmgEWi8UF
9y4Qez/UZ8AnnyltEMdVtk5Mfg5IyBeiz3KXHuX7FVP1sbPpGvEPPY9aix38c/Yhd4myKaat3WAh
UPAQBZV78A4pUyHKnCiTXSf7SovnqEs6SQ8XhFpWU/cuTW4wHkOJZkBBtudoBDnOHdGMb/Ahy81f
UMYVmiWsVARJnVeBHDCvalTu+qYhjUyPBcIb0lkvCx9bt5f8ZlwVyJ155pKHdG7V43F0n2hX4D/7
Zms+wo9iYR4lns3bOb7k5fzrcRVEiSZhAwNG4aUnJdPswVwSjt4oh0v2XxUZXtEJn9jnuMfM6T7S
qPznESQhgkZ6b1Ai90tPSAjdpJVsXuz/RGDmTD14yKIAwO7SZihIcfSHNjx55nhzUBvBk9Hpl7bU
+9lWp6gtTnLUo81qRd2tWxkPa0oWMX17TWrGn5ufpmyfAOwP5IQSNg1HPD7N2bXYHnhbm1wb5FMi
+DN4cokuZdD0wVqlLDiEVHB0R99L9GxyjxuU9KwvMKl1oAjmCbyqgjzDvvj6IfF5r8cpJaMn2ShQ
PQcow1C0BAwfaj3mesomhypV1tQZijIIUNbrzZc6UVHzTt2lzkuh1zNHLOwlNvlw7akA5Onnuckz
fziA+OSug6criCJIenO0dk59ec2TvMsm7PotB3smmQlcw6YOxf9DKtABHNtc5bPyLfBAr3w0/WYZ
nJTdXxX8AiBW8zdNPP5XnuPKdw2nJaxUHPek7MjI8xChPjRryTLhZJuUI62wUQbHoRYu5Ex28OEj
i5mbZaAEtsnTWmDxks9e1CGtd21wBhKa1EknrSiJJ6heayfmN4wVi0XJe1jlwziL0kK2WJhAc0/p
IlX7vIWVsVbQ+yOQhgG//gMgyp2BDs0uMtaXYsoHS6pq1jNS8JJOVjsiA6WM/I0u4q8XB+hJdi2f
1r1yAv/VI/EHWGY05D8OsQ88tlmsyjlTXCtPJrpRef/xoDD0Ifl3y3kljoNlC17oXvI/OsPGNfTZ
qxU528+Tw/nYNdUH+l+GIkXQVN+tS3SLRAirNNVGf1kk/Ovbrt0OsXwvf6K8XiM4+np4DW4Feccu
SIuCvmGhEW4CUx0eLW2aOLWVe0U8FKGM+C+sr6aQ1xmJOFbA3KvMMLuRwrVzT3sOxNDXK7jDGXIh
BmONuk1M2z+WpG4xSfo+YkaaBitDjHGqzkJXBWZVpC8Ne2/wJeANkhIG6RIPIZnH5PVmii/8mgtU
OWz/1N0OceFUXMSF4zb7XZZJJkgQ5mzqTpY4goVU6Jp1G/7FgxeKZ4SJtR/K8qskkszMKHodGzrw
VFNfXCTUWKtjIDZILArJuT2bh3Zm4hJrUHOr5E+iKCbAp5cGUZ2TUunT62ZeQtgtZ6W48Umcq+xm
aeEnUpAfjGPxZ9NfHPQICXUaTUbDgWfuBRHe2joX3uH0FLO7F0TbQEqUxsB5XibDGcPkgVzeFVvm
yilQME2LoUGpdN1yfdCQJNbLFnyc6bRpsHNhz4gxgcixl2Ks27LFCn9D9ArqFOPW5e4i1cuBmpAW
M8IVj0z98aSeQPaB1MtDv7fgdPsmQ+1nhGl0BauLF21H0UtsRvMvvUdIvYT0B52435PVdXFgtSdz
9hGdJ0Dp9oltr8Vd1Ns7NYXdn93gAh15YxAiac1qy8FLzGnu+wjVIHjmlvcIEQouqn375+1upyDS
u/Bbh9ifFrGsON+z+XoJs7E0StWhkMR3v32y96ppZ+H4kgalAvnSSr7gzDJBTpNWh0t4zW3xxs9B
Eop4nBLk0vQSNelGgm/78Jui88kU7DYHexSKjoLewb4fjRJbEMF7wManpARQCgghv7OUOr8Bdc7e
/ZprTCQeUeARNPqxUlxB5WagVUVX/8vF0wg6/XerH1saYZ5c0psMwnfRZlHjvpEctXSrf8YVfFcj
EeP0atTgrzNbf/EDb2CSYwuzh4W02j4IPmv/6mMcuZRii+4eztvHPnZTq0DXR7HZF29DUoMr+hsl
ui2SNFq03fhNHOYNicYp61pBEd3Q3H69GdokJuiR2OzbUZUOs6J75M8MkLeYGRZ0LLNLR0JluTJB
Ki9cZrLCk5ym8SAPDBqKf63iaRyX1V5FQa+65PjtCZxc/R89jld3NT4xjhMsdOdp/t//9vGOVpfz
cGTuNG7GVQfaR6FShsAGC533PdEDjzQRh2pL9WuJLAh/uZ9GFk3kw7kcfApUeRa53EqdFs7LF0lk
Ena6zw5qcr7Hqyw9yxO+rHgHFp/bqGCXRbJ8hwlUit0HOyQkd22d2bnGh4t6wNKoODDY3PVTxnPf
m2IVk7smeGIxz1yqSPuqyYxCT2IYblhf3+neJdoQRcdjLVhcnivOV934JFR3QzxzRIwiy+cMINxf
cD2efsBCRccsH22fZdKt5/QZgh/NgwS7qieeNnC0mJH1HJSz8NyrpaIj+E0xjuE1/hxAN1aDP8wA
oJrs5IJ0beiUaNxLyjgUvI2384rHPXcl051ZYUePdGOM/qrYh4l9Z2zn2PocytC0H8BtwgsxunQ6
/dTviBfFvU6+J8upwuqu8rfF6t+ApDT5yfC2e38xrn9ENdk1FNkH98FlxXTb9n9q3UJrIWmPTOHk
taJam8IjvE4lY7Ri1nrqpTN64IAqWTKP9wh7FY8+E1QqdsteHHCJGL4l1hQB9/qBqDha/gU7wXdN
/uPqB4CfGpfxpy4HhKI1ZVkZTR2TQw7UHvYUamyRPVOwe7JCD/dgia9hUDclT1QF6m9wuYjlt7Gx
gh9FAkdmgIPUseBhf7mUp7DbH6hqrnC8VFvGYElorCKdF+XRDJJRkGzf6x3nqFSd/wcWReb50LJf
sKcq2QYibomjc+YHOwRtSIFkA2gLt5CcVSE+tcZ87zIAtqFV2cecrpY+y3ZCB4x47ur4EFMOxOhW
4coYhYJ3DgTXpTHfDH8FLNDlofHYhMtukMy3YptB7ZUEKwrwobUxQL6glp1U4tVqWerLSw1T/mVZ
EDJHhqURIZf4XvKspWejoEDjMruNoc0ztO7q3+u5ibJqY+C8vyr0a3PmiLe0QHKZfnmsh+Lu6oE9
x7yXPggk7VF58ImGPIZeC6+Qgh6W4Bwwo2nF43M19vSHts2iHjnFb08SiADKPLqWCz829ag7XUg3
yl68Z+vatefH/fItBeZJWWEzJHKLmJxnvaa1a4BlqcYe4hXdrdNhxPDaPqZ7GF3Ts+OzyPRwncPA
OCvEROdb3rcPRt7d/Aimg+a87oAzx2lNN/sU4veUqH/uChH9dIxOGOolQ2zP+vlWtkX+MDRQlScw
wq57OyyKniFAOAT2M3BIhW4t9NfnIwQKZtNVlLU/43CizY8asLKtyM7xABeOt++GcaemAzPHbmVH
CI7+gOlKYqXrzsm+dUInNAImCpd108i0qwnc+u4SR3xkL8MPcLSYijodM5y0bUN4SYZZDU0fsA2q
NhAh2zRh2XHPYXMfHYQQbTrh8zN6gvrYrPawNExeM/0/20FIKtJDwPGzlVDO5L+k9Zji048EIs+7
Ji/X5hebwx8aqSqMw9+PeDOK033sm5L1Kd3mkjbhLwAfX6UJEFAyoSi+NQdQkSfGPNQ47zL4vko9
eOU4Aj9qd87P8rd2+u0OxIaPbHNUuOloqz1kbX4py6n0gTNDlX7d4bITxZsSfKUywyhZ7EP28Vy0
7x2rZBzmAu+mnAfsHXwKWul7Ba5vJNLi+pc60/F1Q1SCwsHDOPa8jQHP7+8gAYgVHvKEpBUOjIbe
kdo3CLwfV8VmUvf3Uc0FQSmueTzKo8Vb5cNxnOfDrx3Sr3bIghE8nBXPFeCPKWrM4CeXUPNc3Fgv
lKY2GcNz3srpRvDf212KZMnqo1tHOZeH3FGJ7RLhOPKrDthDcCVwFiN5gS907a2kivXKIR2HcVym
o/FQVkjmATwEtNnvoVJzG1Vv8LEM1xtDcKF5q7AbmZequxF0RckijtCGIk0dSknb3nYbjFDFTPw+
o4F8G5YQ+KZAdeXBtjkH/EZzMcWqfwfhJzxx7e8/liKhrTYf/w/RJ0hAvm950/zTpTPj8osZVqpU
N8yOp1HWo9ZPRBsSxS9bJwNCa184WseDccXI+loY2JvyRdj4KYb9vgn7aZxg/K6cHx27+vRAv0u6
KK2SPCsNbg2jQ8/Aze8B28yk2CrflcPk6WXmDhdeQkB1EB3useAfg1+3nANJ3VeTyFlrR96H9pab
BNPuWPFOxT3uXRHLAOocNKujAQFZQ7ES2YYEUlqiNxpGjUtlm/Tk0HQt+15hR53VfIqwkOzjPOeo
WUX2Ql18mvZon2DCtkz9D6vZMXtPOsxlRBNQmpBNA/3F6yC8e8t1F83HGV8xxQnWCeQFbPwS83iG
cf86dswF8VuLKPg3xuPXgfOLwO5+LBEG6B2caExd8cb0NcpVLi4ZgEVDw3Qy7Jhu/ttWSqlK0fiP
WRNFkfxXU5+ahyRqn0GM/xYsyoi22dVEJscU3DCKfzRex+5mSq/fvydiZjJ5mNpM433PJAo52a43
by7p9QOlGI0YYOGUaelCyUDyHam0JkZDCLX7fENy7iczvuF9TdJKN6sQCEQn8CWkFjKI5IQerqzE
ltFQWUCPXteXh1Jb72jcBTpuqOgRLRI6yhDhmWaiMFoODhhb/mH2CiDYitXHmF2F3P3FjTATUf9m
QFEt/sZrpRB080Wkk1i1h5F8HS49siWeup/mODKqc+Rs1DIosKdNn3IhUhXMhKixzn2BEk4v5Jzz
H0xvVpYWJW6IBVXa/IRCfcH7EQ+5AWZK//8gW42Q+saXA4zzyurHrsIjRLyAYCdQl42k+aeN3IDN
szDuwdK+R4aC5eEsMTLVmimyIV5Cvmw7+h/gtEykF4jqlWEVPvt8MIrTLGlIGT1tVTWNOdTYFfbW
OlGSEUmgd1ucOajScGenWn2o0CDqfEOBwUNsjpejr/8jpbe4S9g5LCmOISZ2la4YtQLuQnQEzEUJ
0lyOoVcNMC5e3gyNzlsUtxWh5Jm89y9hHCGqjRjBg2t3PF8xzmonB7QWe64q6XtrQHfxbGGB+GnA
kvramClDNPD82ypl6p3SN4sF2ugfWE9D0kPUfwU626AS1EoCLI281ga/zFgXl7mF+qLKey7cQMtD
Y1ZmOLj74K8zguE+BuFMn/xTL7AAGEkSIsHQMlPhCXaF4qX77xjBTZ17U+J6zWxyCE3iZ5r5JZkL
4vj0uJhVD+RWI9J0IwitfvwD/oLCDMMhLY0b8dVh3PKWnWvbpkZ1bPB14VO2Hd/HzQW2zC8rZsAY
y/YKONfwKjKKZgsx4tlWXa1H75QmaBYCoTRt6cKKG71cm0yexXUKz6ZlGEh2yFP4Wcmat6TUhvMn
HNQfJ6dhpv4Dp6fyFdOSuG+czzki4V5OxX6XHbOQ7eN59L5V1F+nXRt4UWpRz9xQwQiggQ2G/3AC
OprbpcQS7OL6RNCznOcZ1HBvt+1VpFn8ldHxzsWj958jXlIXtwHY5idHuUycbRRDw3/b3542NgWB
jBE1P3/fdxSxL6THPJbj1hnysmu00vnkq9GhpmvtqbTN8UwnC9X3bel86Pv0LjDCCnXkPU+XIxPx
YJF4RRe0NXSbpmoYkfK4k1+RHhqKIJ1sQt4bg3mE30+edsF4wjS4nmkR/csCnlFiaqVO5BiSOTNk
C+NGiUlYfpZqSQOwewjKAZ4EOYYkjtBZ6sP4gstj9p03EHjaHGsYj9/qOjtlQ+G8REI1c7TqRhfp
9sSVryRgh5WX8Rr74uvmpC2eDqRPQhJTNfda7Uy59nkyRJHhQum6ClUsTqb4qFJPH+TI2Ssi3D8H
FZCTMXlq7eNsnZYSo1lYEFd975Ac9jwv8AbMg0nVVb60RzmhhaHrXJGkVLNXKIveEOn+yxnlSxMN
x0oR2oDx26FFeTZd3aK6lQWqkD2WI3Mpf6HWi6fPb/hwhnI5skpqYOsR+OWhCkOuXFHi3LME7oPO
kj26DQ7fL/pfSfblzNBDxn9pF79hOAa9BPEM/cYW2AIYLrkYEzrQlalzs5Tu3uX8SZthCCCBWHY6
ggIL5m5QNNsitCTChCkjDAnC5dh5+ui4I02CCpCZW5X2/nRzL1zY+2u/WkL5KehNWmJBTWbmPsTZ
8QLN4roeA9BTe7T/Don5Tkmac8STQCXeScwbITFBv5eiSzipc9rKGGl3HJC22JhUhpB+PHQ1mY7J
UGLUmRMHUWNucHWXFJecB6Y5EDu8CBs2T6rD26U8ylVOcSkSb2cn5Cm7/WMfrdiWOZZMTJNIcRDR
Mid1wAkYIn/CjpC3uVydZBJApKyvRGe0ohKb4joKyVacIe48dhuSzNrQZCpJKGMX5+1A7hQwY7pD
WdHdpMTFOQ5crTG39SIa3/ofmDFkrXFTzrhby8C8ywSYINNg5K1xB+gFr2mLWAWmjA2Hv2iwGgjS
pNEsXMzFcnlyY4G9Z386foQZYLCnDl6aCicsRwxs/izX0SHvQOfMNEdXCNl/NksoHY71IcXdKmRG
MTz567IWbJ/f8FkFyAt7HwxA8PLSdZCRo4A4MO/aoITYp5YdOBb5NXgJcVRcoq6Y9R5FoRKjP+Aq
LmOtjKorIZWlL18rA4QnSupjLeUnIjPBo5qpszvQRwxcorlm0WJWH8dnt35i9TjIsauFB/2NtPHo
UC46ofJ+T2r1yW5RNcgSag+vXUbqmienIMM54RL1AiG5hdIMNwwxxDdMHchLQfjMaDn1bwJaYKNs
X7xWqEk6bqiUtMEBGoYv7qmZmKRW72mwCGRDU/2LjCfL/2rQTf3bZVXIEcbAksvsPeE4Wn02Y1YS
isl1iMyeMNXPvgVCuUR6p3tjq2NdH2nS6OGFjkbdmKlhiLvsl4KGALGd+j/gaxwdKO6eqHmEPMMJ
TB+Nu+4mIKebcT918CFgwxh/H+XVYxfKlF0cgsDI0heiud+uUc0RIdic17ecGWLsPdhWJTvokfEi
khGcdsawld8cqrDgQkJfb6LvFQoU3Wro6HL5xJZVpLk40BBLp19wz+ED7DQytV5nxNG6N4JPh24U
CZBOoEShdqkrP2cQLZlA0wfwyWb4L/cG4yNByOEcPgpPpWhn4PmFCHEe24ap3+XA/TQ8g33+2uUV
JuQwueezXheSNioc8xBt4E7CMDNWro3oRQ1bX97sQgGAb7Vji6QOvfiqm4ydm/blUMnhXotqt+X9
dSYnI5e8w2pUJZ+/lo6sA0fCqF7oHkU7dePxPNDjbpffyPl4OQ4XMAf2Eu598x2EW14YYwKUlR4H
+Qbspalaitil+ADQAm1OsBqsUy2aPbw56cgVsxy92nuNtTc6msPhBlHGexrtnLYdgn2zOgg0vvA4
TZt1dHlJcqhvrFrc7pv7oHNk2cEERqEriJkBE0pdQsfRH7TZIMv5VyvOz4xDyV7sD+mhBcc4If6M
whFDwWlNCxyVlmWVQPrXRD0Wc+pg0KzCEwqU64Z6VGENuZ2b2sx0XssCZknxijueAQGGnoQN08KS
EulAHUFD6xsvplH34DjidSG1ke5Uu9dYHxPaQ+LubxNJrr6VGSFpo6xtFjri+CwFZ83jU22yGazR
qJF9WHpT08oXueghS8e4/VRNjLxVEfVTsfk/1kahsxfSUZ5XwRonOp3OitCyNmpyfNdnRXue11sl
HbKO6AE6tiTL7z0/uHjLI1PrzTWpFGDHvX7MvX8dp22LS9cIof/h5kTuDFh8erfSITZNtET4jwB5
Z6eEcK140tsczYG4mCp5ysaijEusH5buEico6QjjGlPIarnK5EiAKpyy2PfprXt/nBbeS8fTkNz4
k12SilwyrogGyJG23udKWEUU/NPATzDOrsGGwJKBUrTPltKx3nk7Y0LGd+iyd1NICjGPA3OgWPpO
gD48rCwm3mCOjuV13q/qe+7cZjnVUnvL6H+6GIBwPcOcQa0voQ2q7L/UDx2ZKR24ZInDYYo6l2tN
88xDRFP2VQyCWpJZQjb25+4E0+UAINAyTF+NrQhTFX8/voF517nbvySZ4qSTqQWy0OfLRxsBu96R
VjXiBYw7yASz+pUjyW7yDw20+w/5zbOTftMg6tZJ6la+IIGSCS4pJsR/rOdiL51VaXisZysLx4zt
H2WuDxmcT/66R7xZj7/F11V1dK2SXkIUGxOFxJXVisQRL1GW/F253WmS6Zf9CKH+eN4Etnak+YUa
3TH+I30PWU66lpxcycLjdPPmyONtPrlNxuPwdUqd1LHElsVZBImek3I1r9bdhUuBrADT3TRDdt/h
BizUtv++stBuIreR8svQv/2MEVjHRdrvu7WcE3YenNt3LQ4adR2GzBcHrohviStA9RrumYYFM0QR
I/9LN9e+pTJn0kbvbmARvsP7fVjlIOHy8F35O2/fT/uEoNaQCiYECZDvO7rAtTxq0aIQs3SMyjpd
e96nsSi/NCoa+MIRWt/vYqBxxI/d1WZ7YrxOqDGs1CDEKiA7GkldwVJHC/pzT3HKvHHnxIhOFwxd
vSocQKLixeTuz4hbRRkcGRbe8eqS34AJJFydI2YzNmu2bRxsbuhhtfPcpSRipqeuDWWVFXVM8UYO
6A/91IOPr027+MZYV+BdlLQarS+txN667/oRj0HWE0z+PeTCScEDH/wKt+9eEehzZKV4qGeym+KE
JsS45ipQLr9XJ/aG8oQosFA0ueyVkTLgUj/M9BwrE5rVhFw0shO8T4owx3Ot5p8avf9x3QXtW5l6
hOKeb2Fddt34Ja1oWAz74NMudIcFeLxCnCq3Z3NbYNEL5xWWcSAJ4xg9wb0HLZTykb2fZXVJwOCA
MdxSKbylk9hv9UbHe9txPLFs1hAfoINOqIgxCJ5G+miOe39cROCgHo2sIb8HKYWNWpHJ9+g4i2Qo
jHhL/AdPuf8W3yhZZtxDJiDkihZIkfvcFKd4APiSKtWEA/srw1k1PrVv91mJiasAYlwfm2CFatmr
OwEdo2Y1fWdoO/kGe5pVH4do/cebMpDDjDSePlMt9R3B7ckBqvTfVsENelZjYP+T5flO07mwRtJn
sLr6Pab17XoWzAdxIce/vizKwhIPrc9r+jybVR5NWI6o6deKKPNsdLx/LonneH7zoel2CPv/pVqn
v6eIieMu5l59lNlmjCXxo8yf1tpUW+6B/rArtX37uKD5aG+rKhffI7AHUTezaJ6x0cB7GGHGosKO
f1kN7qsR/nbiInznkOz0bIaSr0zR+gWoShKK196SCD2N73yCXluQPUJy+3CnpxEpDX6Ha7/OEPvv
lbqGqR9BwF11DDgNJTPe1GpQK5JwYLH0nIxAnbOYhE8qZkq6crdJ4IDYfCzBu2Uv0U7mwafTaaSs
VPpyg4H2qC3CxumqhDQ0qb1G7BOo09RX8qGjSy8E+7jtyxW79QRyIZmiW6KRmNTQogR5aMzeVVVH
R0G4Z1sVQW1ugq9ddeqDjUMTgvsvK+SMYn8BTuGbLXKqFrd7VKKjc1q32vq6+BukzLOzn7+hQdo7
WTDz4JV2WjkzEZocx6ZD72Th/K/8qx7NjruRviiCGIyGQgBI3+MUt8n1vJqd2DXkK0JCEaFDPogJ
9IPElLmehRBak2+VZfrV0Yetxpkit/VvKUkWHCIrFtRq05XqW2nHe2E4YAVamBnxPQpI6c4V6whR
2shA5k6/ClysNcyvkh1fSrFO+47DGAQ6fkIGuY1Wy63zcTPyogl/RbbVHUyd+2pSR3aEYrKcmBh6
gQdFX6qSsob0z59GThmqNqFcMeSa7L+T9bAoDSAH8vO7C0LHWMc7itQPBuAA9ut2mL2M8tG7TgQm
Fo7okYX5D1x/R/8o7owfnWPDsaR1U4EitKRmsTbaUyCXTIkzOWo6bf6Za3dEcy3EM3wk+AjrnQSl
bjLhTjThM/9WrFkH9x3YKFSILGeADX03EydMTxQveKIm4Riam6ncNJmdOKeiYJVrcCFayUgmdwGq
ez6dEx7UL+UT+RFeUjvZmWFGIs4Ippy/IGNKc1ZtOm416vhBUwbQRRcv9XEmOI9rrwB++ZSQlxrQ
GGj3KxUptbpuZgdQrZPNlJj3oPLTsgTioXr101ldUpcKJlXU7cNqLQ1wlPRaLZfNiYZkAaotmWZ6
UyWHkxmQLl5yACAKoZZnXuVUzziVYaOTZkMjFnJQsjpgdcP4QFcN3Zolm/wqnFQcmruJoG1txd27
SK5U9G8UWGKiY6lh54LJ6t4hsP7z/1rd3yhVdkBDkZ7pmlqAmIE1HQQMWwII80zntgXs8XDI7I5X
1JDV8y9qGghs6VI5xt6tuIsXRPLDLdEK2fl1EwwExioACF/uv9/h4PS4LNip0acvfd6lnVswpHGU
KGG9yYWpxEP99eKn6REUFjVZw7EK3xeoLBx38qob3I8iKafEtfiZI7ZUse7TH1adRqey1q9ViGPr
U3/EmTifU+jqt1+zHS2vWLFOX6lv42WY6ltprIWrbEVnsLVFQpyCT58XHUnjeg5j+QRvT6OQOI6U
wJgFkFfc3x7aPt1JBaNocEk+cLDWJJUNF3NVlOmwquRPwGEcHD1WsAa13mGLQm0pjzXDoM/BnXtx
WW/K04I/PYvDGHSVPAFybmUr0kDlm+nRHNz+S+d+P+CZ+qkz2oV2TYngpDPxa6XaeMUiwa7+GZxL
CSRLw7J5qhSx7eDlItKhTKdUU7pOMeJMFG1eJV8JHn2upbGPGAaUyAf0U4DymbcXLV9Yqr7wYQ4f
TuVFYxIyl2JnSJzqqQ8Azs0xJyjhraYVkTC+556O9PCLlG1xo/DLkCx6px7xCxHEqtezJ7B6t+ob
X2JZGZLF6Gr7vbWF2AyF8+HMON8LehhTl6Olmb0VtsNINMcenzxVRVAVG/UD02IQ5AzjdK8X5NLt
xD2v4dB00lhYhJRwok26MpOvWF4p4kZOHGf+X8yS/r48fOShXEPzY1KU6fNjJAT4vRVeIamLNbwU
5e2Fz3Aq3O8i/RhN7w95HmL3PrxSLeCrfDSiwmbgm4IdvhL/QPMzZIeWY8EZ3J31NAkgf5Ukx9Kv
Z/3IULo/KOFSQrzUkoCs1nYPuhRO0BPmsTbGhWGPCAETMp+eTvg38J8e4L+ICnBadjeDpYzIhpiI
FCPivqoT1bbe2CBa9rcmtfhdIb+CPw91KVfjNIJlWQiLeLLUjqUaSL//cSY/yCdHBw9P7ifj7diT
J4WdL+6+lsPjMkD+gIDTq9QHE/e/hFmsrksq61yqz1LPTzYtecO2SFVrh8OKPmz+6vpczcNxlx0A
8Z7ab/BCD+8SOJCGPYnw9DrkOBsjtXLI24HEptZSf6PjqryR91yJYcIlbzbsDLRDpviKyJaV3M6o
MtStpWwoV9uxtHHfUA0QMw/Ykgmile/jFBjonnNPtArEB+Hz5Uyzvj57bO5EV6vf7P6onuh8bCdX
09emhfUvA1DD09Yo8WVLJg4h+DAUGqaPCqvPrJ9F3Y1HJDT0CK3twDh6hjCQV/aEssymua4DAd6H
aD+Y74mKJGI+JdzQg6St8pbCYC+R5wFynjv97yTSWF/z9+oe0ZRpAgVYotLsjTZ4YCjTy+iDILwH
AXpkz/qHDrljl7bIPzwyav5rBY1V2H4+SRQ5O95IFZqmyS07DAc8oPFK/rC1cU0ZYOijlhejemAI
lgG5YjVe2ZcM5jkLuA9suCh8yPxusajw/3+VJyRsD7NhfiW/5sW4HC3SzTqD+69NgkpXuVTdDoPa
GAKLtsA/W1RaJlmM4E9Nm+xJDkmok3+FeN20aptq+w7zCuo+T+zntmyFJ+bzdZuPou6eF3CrG1L+
+ShKAj9pCccGpNP7pSPtQVnRCLzM35aEdeM1q6UooDqi5VlpeL98YBN5erRtSzEI30+vIph1DB+D
aVP00dql19x6T2bsDeokydmTKqeCcLqqRYKXQNeH29QAt8pUHRIV91NRnEv3qObK/JM3sKnll9O5
Q0ptLchd4gkvE2dOKkKhGLh0SIgKkSGS/1XmGpv5z9oFbxGTSRIklQLKnA+CByDAVDioA5e/mq/m
dxgxhZC4yTEMaSYDGdVY7hQurMYcNuwrSIytFBRBLdOJ85+HWOyCpoAJUeGyZR11dZK0exivIJLd
eM+kUYHCTP/x5Alf8baXDO8CcyKPc4KbUarDhcpYejFF5azjuNVULta0FPfb/2kaBEs8EQikc2p6
6Rfixpiaa6pfF53Q6nkSUWKFqUh9xV4ztI7Udv2uy6+YVRjorUwsujVo2QpZoRBFT2kH7lMsvlb1
an3uUuTtcUqOE8BW1BFLERAi4t3NormdinGPj15+GjrRPQN5aS+6CoWdCtMQV9ecfCbA85C8UxvM
OBgH9GrDRC3HZ2zmCYZW6x7icME6Xet4kzC6W/mdwMhqLd+0p3JVyoQIxN1QL17YLav9Q3wl9Qf+
43EQ1w7J0zbrWeVvTd6p8RlZTIMD/wlZ/GVImemvOMuvLrnt2pkxdXIBFSC0j3h1bDxtQ0ewMwET
GNeNtRC+1S5UFTKC907LU961OpJvuQrUvokKSisDsxz90OdGUNhnCiFCF9GwGsH2jw+Zk71Syeav
bqPhakxYR29pakTHlKphQZ4jdYD3jKU801il2EI1PySgnnqTGRTi0IPNh2+1q3pYb7qkO2wyaGzt
hJ3yjJFDZMLwUcOHHI9PUs2731EuF6YeKxt04elU8Pef7M/2vWbTL5cZL36OwkEhrEIPusdvKuVX
yHBqabFU8EDvPxRWTTFvDFR3La/Aa2iz+wcqRjExhOBrApZYE0yOhC3xq6+PkgrAwmQpuXgKU6nz
CthHsttZPgc3ipw7+Qwl4wnPjTUga2DwoxIClvdZFHpgZodq6UUlj/vcEfNVpfJcnW/f0ai06b2E
HRvK6sQqzcYVAnpfOa1HrZN1OSsw92kKl3b9xxGKjdCRBYHaZUWisL6wDofDB/EpbH6Y1zOb3jx5
qAo0nlTipFAUBmodiLPSJSs1V4fx9t8rt2J7TbvfujgbPGb3kyKwIyyrvMTOQ2Ku+uPz8rfDwKab
3R4RfBVtpw0rQwvCryE8gGkl8TFI6IiMhujkTrlaD56zzyi3nfw3fIsla/2pOZxn5Btn++SCKRBP
IsUpNtYMo+5NlQiUPgeKvTfcvTIR8LFaSaHpu1a7cUqGcND7ocWWF9NR+6roit7gvirZuL0Hwf9j
pJUS3eGs7niJlHOSybQPM2Nxry9cqiU684GV9F1CJWn875QGqHxLUAfeXPoCsF+EGy77EcLWHhST
xV0+9ZxHXZKH9LqhnWiUxcGwmo+MkratGhybXFnjEeoSNSxUKhxcJbJ9dxXfMpg7AZsf0zTrCvI5
3J5Xb1lj4SWHEvgWMRwZ56QxAVmQB4W7zsePQnnFviFBno9cKVbDS/bmpimzIfJLguZBggPPfZsn
l7tylL/FfXCVSiwIuWlFfmATQI2ov2G0ToMyCi8JMGP1vH114wgZZipO7QZU6Rw5qiEE8uTgr+kC
2VVz3VS0fJQGeYtSjHGcmkpMNg3wuPHlXm6Tww7sJA2FwCWkqZCcv/mEBSwjAhwbdU1oHXDIvho6
5anQ9ivAd8xF3ulbyNecsOjevUy0jc0JafcG4rfaXNx55yDlpIzSf09roFjhy0TDrGg2GK45f3TG
7oRj+8Y49t9pRjpM9kvCa8dMiGsiiDmCp0a00dWsOS4rmRckYprVsDDJINFZo+lWBfLNUAcTb/p2
7wRPVi+Cd7gKRk+qVdebRvr94d1Y0fbGzU/xQjABT3rEKsh/UIBZKl0G6xaCpL1srtno9hozUlW8
meHbHpusESfHbTC7tu6B1CIzYDHsGDwywpaxXZ6T17oO9Q+YTAHF91ijIpdWzwSL+NpL0zrC3jlq
PvY7q+3xLzn8JpMkttM/pyky2TlTUoi7IWu4SJZYguWZW8PMc2Ag6K7VAfVNjq2xWLT0nvcqE9+V
lLxPo/hgFUXuwvF8vvx0OHjPGIqe6+6hS9RlP9bbDfACxxWK8uaLv2DWaxky/Lk1/Skg0JbpPK4H
n7r/7eJMa3ys8p8FyqdRGhPe2D7VFQRwrjvD6fVETO5qA4C1yiZsScsmmQHShsGUEGRtZTEouKYf
M4YR8L1qnCKB9VLBXaITkZqvysSHoEMUdNY2neqdHe9K7Sz2VS+K4gaLUcZBkQ2Z7T+TmUfsC0L/
Oayi14LzSSkMc7RDADxtY9ff55UIkRGb+UiPB6z4tS7sv+lmv6amkuPt3WgNI5PIrk3D9MDro6Xb
bOk2gDF/x7uyS0txp2uRw8Hxem5pWXQEGjqk5u9Umuw5Ly8E5CWpeiLa/o8NmaSTY+yeb+Qb3ubG
7KSkEzVhwIbJzaArZvZ1ObozV0Flo5RqnuK/2tDSYLpBqi0qb3JTrJyNfS6vQwqAf/y8bOLFDspy
4sqdrEo6Rew4VtRs+xfKv37V0a5Ncg2QoZY+O3fqJKCSizFW7LLHkyd4dHu0Vuz1lZhbhg8v8n3U
PP//xlziZCHCktthOerigV7rfGoTH8cTQzDEvBq7PYaFLthy6LAOt0HVowh6VKqHDIShglWrpzur
3YHGDadUH6ItFt9YaIZ27I9IvT6k/5vFd9fo6j/hjeK0b17g9n4XhvWmZAmg2cMwlKjLU2rUGGyn
6b0a5mfZ0imxM43RifuWtmmm0tMVOEyytsQoCPKeUozwJ0Cer3HO7zow/JjbGEgY1rKdQNbZY5vu
LssmCCrc8ByZjvY/GnriMG79ahLZ7EqJnexJmWXzJhBK99Qpeluq3AUskOCJZNPusfkHB5cXziqR
uF8M9FENmztPu8pXwi94f/fTJV2H+NeBXY6Zf2JI6F+uSXQ/YWcCP7arDHItvbfFTh72MLboSznO
6eJ41R0twvP+aDFA+I0d8aJnG+OX1YX4g93wKokzNjeuPObG4b7Sr8rdD0OMySmzYkBuP7+6z0mz
ZawxDaA4vU26oWhYuMZLUbkZZ7DoHJaFE/j//KL6+zwQZAly95mBD/Hqdp2Hd37diHRmVvjCUC0I
uri2sIubT/IyKcHora/6q01KtgzncgZn5oES+50xiW6+Kelw/946NdEsDxOSCaFRUHaPlT2IkZF7
54neJufdE9l5nG0CgCiqRhminWj15++l5NzV0roIYqDhq3luJo2X8lmfBhmzOXjqqE+5ohgKqS7c
orkDhmz+rJl1i34ux/dj1UN+6q91JVb6+mw19ZeILQ0aNGq6Y1tuSXv1gFB1TxIPiJuJP4qadfWx
ZxW+1FuC91Ru8KGPaFPJ8gCNL/f3WwA3X+S88Y3+BDFmvsQtZAF3qssAZhyIenSW70UHK9Gok4MX
ci0w+IEVfmq9VwSmogiTSGpHYPRGiT74sChngBCW7hjBRxYn/0Xb5Pt6sXjPWLfl0IPnilNlg10K
yOiDGR/4WU8OGya3wW6M0FRJ/AZySFRV/H46PdyXsyV9o6QsCQl2bSh3K2OCG3DRelF7ZLJrAtSN
G1xyLIZW/Ny8RuLgK8hm+ebVmA4u+qiB76gaCNSovAC49U7lr0ramRmuzgJX96jLDgUZRU0f3erU
8p+wAjXJNbNgTKvJE6WNYyZd4LZ/EZn7Gd0+NyWiQbvscPiPHd9WPZembGmSpYfN8Od5UNbIUjBJ
B37G0QwhdfU46Fu4tlvVi4jvkrJVuUkEB7wvuByNwj3vAYdjPAMUG+KnNJvrCu2C/3lBZJDvWoMV
Be/QKyoAG9+HXDTFFPNo2ZieLGQKdzwm/kvSTkIf20QfkQ3b17pM0lYSG/poh7AdK19kQQ7+US28
5tjshnP/j15XFxtAddPgBaAN2zy53S4r8ze9XGCMFuQLzFCJ0bfr8+6MUL8P3O+IB7nVGeU2Y9FI
rm3f6L5zINU1iMFg6mrCo8FQ9py7mJmEFLoyS7m7RemUBPFEfeQ8oIPez/2+Ibnfokxm+GbBUAEd
QCrXC1+QnJc13ow7IcKVtFkHy2cpoGWZSBQ1JNTZg/UKVNmOJxRexDimdz3nGQ6mylT0o8mGeSUk
5MepGTPIEvow9JtZ00yQNiAAoflJroie/VNT7H8/17UkReXXREfp1vmvLHFjJqufrZgccxRTLxp1
xDYWG1tHbkz/MQIr17UZXQroGLDgeMVltF5kA6dgn/MG91d9CfLbBrkHm/FEEMSi7z0jkEi/+2tk
d2AlVvNJ8D50E1EIStuXLzP3d3kWV3J6NxTegMXXR9kdzmMOk4yQe6YiasgK17pmFeAxGRSjn2+C
BZXTmLQl8Bh21pYCf2u3YhNZa4Pn1bF70X3eg36cr+cWyiOdFDGCH2h+DvHaU0KE+te3VmsPqqCq
0pkFtrBALeEj+PuYpwvDmFtTPT9/tpiVqJSOOMs4FiXZsP0UERG6doaxZlaoJDfeDC6/LQk2Jltn
8LWNWlEB/kee9pGheKkyCT9j4qsiDi/XdxpUheLyA8gdywFDC5XWcBOXJLWm2DX5IJpa6zvKotLj
H89jAWmD28C8MJgqGvy4ZvKtAqo362LewFgzReXxKvTCnGTdMMgAh5W6h/LXu9/a8F43JxpxM3jZ
acnrKd1FZtGr8BwrTM2VXfemp9pP8r67bXgaRsKEgesvRoLoVgaOWWo3MogoK4NktoIw7CKoLzzY
AawwsA8fdunRWvl6GI9e1BHMS1PoTlzBgGIRdKKSxBhhKMvjuxR7BOP8SorKLJO6CXeIa1jlDw8W
k9UKaJR1HqITqTeWMC67c9qVpW9l2NUI9h0hEOJJ4Z4NX5uQVllM6MfjQZj+Y0vVBc6WRndDgRID
tWqfKDGnyuk4cK8csLWLM8gq2G8vbklaPMDsUzIrxpCKZ+DXrmdUfrSASXadjCX0aqb9oPw5+7Gf
8g1WuzuDPMOVRdFLryLkl5/9+jW0qjUA/3jixWY2HfS3NGeNsFTlDIUKo5MsoU3BXYPVqlcJJT0N
RYsD+bj2EbvAc5pYeTnCzTAm0FANu/N7J1Un+dpX+arZy0FAYZWfKGxHSSOvxvfPU0bRgQ9PzANt
6uBRQTjRXx4V0YC1S+/3um8lk1OP2Y8baEDezXU1c444Re+xeefJGsxPRnTGQv/c1ACZls67o89L
1j/tQZCBOC3P4JeWtVYU/mStRk/0jO0OZJa+SQkQWZimSxcJDrLk+Edakyoq5ybxSFtcsHyaxlW1
0z/qd2XzSeX7fK/MKFsUhjmLfDvROdr6HTGjsaBHwSbzd/slUf/fEjYqNc/6lOqNJsTfYH4c+5nQ
ZKMKjH6xC7Vp7NKHB2A6D4IC8WsRCbiz/VbUEiuqRuF2gtSSwlcEqBHmawXsqtPQj9+uvP5UMgtW
dXvbvLdKhHaV3a4nnxzAO+bFSE+J7+UX6VEbRyRPOEnFqHJ7H4R7ol4MHMNpo7eSOrtHvAMADncn
l00IgNDqnOMgWfsUbrjSYZB82+WsaEG/N2eJlvSGJQT6W+GLE6vySKrc94u+VoeS9fp5hmVy+7LG
qZpU5vU+D8wYoeKiMNg/ofVH4jZkrcMCqhQ99fcqaXwcxrvfle/b7jj68PaK9oawTTexN7VtTUa9
4wguM4KYsQZRripCubUX42s4frqxf/tnMMT06AlK0Yb6xNUIrLni65eGTlpW9K23kfKHq9Egl5oV
kSo8xCLueiyFW5FP4lHjYfXSSlf67J5jPQrhknHYRiyQwnMIOZ5oCW5INLh63bruCiiKbbjTTUBJ
4Funow8iPdJGI47Evt1VTq7DxodfL71DuhQGi3VOs4UOl6wNjraHATh+2tnVVCpwdMHvJ1gLwAST
r16Z8Yh1O/QRUs1AGLuKoIlg+9ic91Q3WXQaOkyUql2q/cO1dNfDGaRwB9wBzKF4HxRuNfFanKe3
FqHxLr+dgTfvT1tUR1tfE6HXqZ/H71TG9T0qfd1HiDlGgIsQ7Er7xU8732LCRFfgsu8yqb2y1WMu
JF3CUOWzbSARq9RTrtEGZCjAESft/SDv0e/AuUQFesa1QxHdmAktW4oDYEo99iyfDA5ObBWT651Y
EKFghuzf2Y5TnSjuG90hrh25P6pFO4GrXpSvKFeBYWyuCuaupJvXZ28JU+FFltvkmkGHGldtRYK0
qVsbwHXLGP1hIZvdg2x1A3YBaqOC62qB4/ieCyc5zaaRCirkl+pYwzHVDgJC8TLmxmGdrmXuNKIq
Kv60bNjp1U84JJD3eFNKRLyFLrDoU4LJ2C3HOexhDdQOviJvv1c4IY3ZiTaYD+BLallet6i/E1tz
sGKaSfg48z8PZWWNcx/om/qglHxU532ITaS/rMLlosElCBzLUPeeDxsNgv0YREnBaYdJ3YWzHe3r
1gV6YPriqQinWxtnssD9EUkUgsEOezFW5XfC3lYOco1uIf2Q/TR3UJYMDD3k86AjCmpg3ZW7Q2rQ
Gv0C4DJPr3kyWOU7zbIduYcRvmeIFvG9sYN6XGFwup5H+Efo2Bc4rtPfil3wkmcYoRgtXuDdDDDs
LBZggT8zTpAmh6SinKxXXwLahtk3Skyp5qZ4eNoSSkuE8IrUIsqjZcWGnqoB8Von8kunZ3Exn0EX
w/riCUN812cGvAxdq98TWeuCcOGSssDyaF44z21hhrrrcvc78c0eAEHo/OLfsJNt45hzqRywJ56W
53NxMpQG7+hgMDDTSf+m3FbXfdxH7/ie2sw5VVKkAmElejG+6KS9AvATg9QxsnoVMS/z7cMqubth
8p9aoyIMVnMiZ6LfYJVwnLeu1pWKT0FX6/0YVtgfWnKipTel/+h86ssBt57L+LFfGIzspdsxp0wz
mv9ytDPdQnpr0DEtYG75piRAN1daO2fbIHBN2whwMz6jXyXefUIcpBmfpwVXW8kbUz7HHUqUN70f
Mn+Vur4wsl3pANyyLTDXuDkZa3pJHo+DmbTHP8990tlPmRLVCOrGBHeNpXnFDrE8BJazLA5t24nB
Z4Tn9n+CZtYuiTt3m3f7kZ/Nxb3jdQ9kkDXFq5jfF1a/bsz2WzjR6RAY2ttXkuTn8K1GHOq8yAua
kMpxS4NgcGIeznx++huxIv5LTw61/O5tkaN1BTI+/YWuBoAahAsD7/TnUPNbWanCKfJfR7I00Ocl
vg9X1cRQGXonbZV+1EJ4huzpubP3XxkmmOUMmM5LwOqJywyQmMy70mvdWkpnwO8J42uupHtGKrva
Yk/s6WIPiAiO+WDVmMtGfWJ9u7J3pkt6LuyfrLdanzAPdUcX6jwyBDL1ondJ08DHuMR/qV6P+yYA
ZuWlbEcRu/w4f9DtxfXYaj7J0BTdF2atzV1rFkJo8U6AEnpy3NIdgEbQxbDqUG9sjvY4EGm5fUCr
5Q6C7sIqukFWTJHHsnD54bFxxRYRZo/OTom7fLJMyVIb0LJCQpR8SsS2UIUxTYuvfk4+Gg2k4UKe
zV0K/TIhVHL6x1u12n/OQLmzam7cd54+DW+RP7B9R7wqryNWVBuhJO4cX8l9uHvRqR6gYaua2h/h
8UUM7yUMu50wcmpN3Pkvsgc0P06Su0Uok1c2cw1pSZ0+p4996NNMLAzr5IwAP32SoeOyMjXszKGS
Rv+rXxv0kVLHTh7izB+BP1MNR2XoxpcPoK6c++iu+2BRvwuqu5Vq7+ifknPwf4mKtAvU4ZJBYhJF
mc+sZptrbnhCpe38LIxDbm9dKBDaZiJfQgAM1S9IGmkwcHHsHeJSDDOc1Q5GndLgW9oZRqdCUSlQ
LAvJ9/qmlG1G1+U2n2CqMQP5FEWKmdf2MoDtuKqRuxfT25uZASzfHm4q7cSZQvLE8Xz+nvDewLdb
YTAJvmpvqsFKnYi+4/rpJdyxc7iq4wycaDrJCdKjQOx4QxXbkzL8TOtqDL5T7y/raAD3+klho1wx
f2+zcnlkgYRydP0xkazcJnuY8quLFzasWUpNeB4+kVQTO4dOp9cUcRxlJ/NigNOlih0pOcDcZe/8
LlCaQRC00xPSd9eDUteKFU2QOu8F9fGor8r5lTOI5w3NNJfwah/bQUxpbnYz1FZlmCwNsTJ9V7xX
JEBtjEJrDkuvBHkuYH/0a56Gag+WeF6JxfJBgWz2h7lHsz4AV1ffqQ+ZL9OZuABCIdB8Eq0PSXeX
F85wZutj8oM17dXBF7ac7h+29v0PtvAFLAwvMWkV//VTKwleXAmkzL3yLqKWXyG9OcJYxpuvJjoi
tX2SrqMorqakxyiWlAFATE9/a07pggSEdxL0vagOnpquPuL67haPbVKW5fkwBR7NjowHZkz1ukPL
PW4v0OzuWdQz0XXv1s2dAmNCROEHJp6ipm+UUGZf8n1VlIIINHWtvA/uetQJeW5jdOMT/jKMgbYc
Y9z8xI8/fUSDNW9ra3db5gxFGK2f8MaP4YupbYW0m28x9UC9+Xhy/S4oOcGqTICUGBKUDMtoLLv+
Oousn8UsXm4ZIGDyg697xlF0gFvf1lRR0kpvUxBw8bj7LR7aoyHbT89C9/MLqIEi/cUBy3ng6X2F
f/1G8HusMfAx7G7tKI90FhYavUYDVtgatE1tZEsrG4Q6S/75/3f+PJ5GLLFn5V+A9RoeP1QLp98q
IOt8JJaqM0tgS0jCSj5v6Bc9tiWFG8hAG+97oU4EKmmY6Urgb2LKo5dzp28yebU9XEu0rGX3GKPL
YVDhOu3r4+9hVyMVi5L9iJeyOBvPVoyf4CjP1mOjmChxAHstDqKuXaE8H9JgWz787LGzLTLohU/B
LO2WkQsT1fVXsXl4nALga09sglAI49E7jIn6n3Jiw7yx+60Bmu8cCzGbgbX0FUkLmhAunFr15G/U
aPjEQVg4UjwAUwPvHiMfG4prrhvUCxflvwtwCBWxriPkkOkFLzdRv+nBJuVYrKshQb9QwikP+Igd
q8pllvXmu9O8awUvnfOiO9JYKKUIVVHqdaE9ABUuSwEUygxBv/WXLVjIvc6xe+84Hn8MAXD819JJ
6BSK72b4I5QqXAz6D4v3kUXKkryE0Xp+3v/o9FlZ4sM9X5FUWSAc0s1+HCE14GX8KMN1sVwMqnQu
ccrrfTQYPcyk5IOxt54f+gWxpHFAB2VxRkUAQiHboAUnNa3PoMVE/7W1iMl4YgNz+J++C5YcBZxN
+yCwZl74xoCF98upHNyuPE9gotUyLZx88S/DHixZCucR6m2Vt+a1DJelq+q4f2PtlzcbESK0gSv3
Ir8zJVHsu6qIStUS6BRsN9f4MeslGhmOkJo3sx7a3tkY3/mZhUlAq6X1kjhbcm9NwNj40bG5TFJs
AcOjkLHA86fhcJcf4e84xxpS4EeWQ6t33Jw1Wy/Ua6w0GzIV0yijOHXx2nd+seqiIZUZ5HCyNepG
3brRgTC4cdfTDvGKlOGJgAVjssxRUWbFpUV+PRzjlilhpdpKi2VL4Zx9UasJZRnWkrv64UMuQHTf
MsKSzyD2gd59cpwNGKa05Z2BIFySeP9dq/v79QiWEA8RT5oT6nUDtHncxVGWYlawQqWkEV7d051c
2z8oP2VFqndzE2V/WTg+MzbBSDR/Y+Vh3r5I045AYFmXPc+YDixL+lDPPgFYtEeCM5c7rL552V26
l0lQ9BWGdbzbV4MHRfKtHkCwlqf726R2wST7lNauSxzdYvAJTyTwk47sMxlPIhrllnC/i6V6FBmW
hvMRA8k5AobosnwISfpp8lyEUhI+TyUo63VykxkRoVKN7+Pfz225dZjYFoXegPXTSu6ihqMXsbIg
1O0JSw9IuJuCjlA51ebxyJ8TwVMI1vHoGUD3iW/ByQsJg+2uGWJmPyT23lI1vFFd/WiVqlv1CvcG
z5TeJVTS1H4yN5FujEqjJK/aT1LkpWK685mPC2/+Y9yPDc1vOrXqr7okL5jJCNynfZJVmkX0ZlCW
/wwDcXaclVD1f9wvSdsB2k/ZQ9Y7aZ0SswTymWGycW/989sV5arZd4fZba5A7fjLAUYIUIPAhzKH
H+WIj74ngWWg+xCS/cxYoquQXiq8uGvSfEzSvTSB1tJQiNtUlY7KYeE017q7l3NXefxG8bVjtW7b
dw7wMiUC71Mp3SBaDKm/da9BbNruuQNOnyHKih/CA25bm4JrU+UNDGqoiemXPQD7GcEJFCpKIEXY
YTp5dyU16AboaaU2PocF0kl3X5+AxgcMoPrivkxapsjRQt/CuR8Uf3xtIk6kIiFfnuEbS6impqWO
FJ6/bFxMbF8BhvJXghJysfw93wi7JTCDCo8tOQx7Hp6emH3rkzqABQ7wOA7oN4e42YU/+sd2N7CC
VCxgAD2ui98Q/+Swn63esiAm88eqTvqWfXV7FvY5WCGc7pI9h9RW6NSgzDg33l/DJvwsXzfN3m1L
EV/a7R5yah+qykQTgGke4Aps4qrCuiqdIfSmyLTJK0rHR/BPDMUmzos92EfzdCVb2UTM3gFUvdv+
GXO4+/d0CmjmjC9WJtaPLjAkA8hbxl1Vld/x1Rlvi7ap/htxEtniZHZWLxcDRaittZnveoqRbrWb
U0g0AYwqDcOLAhSpKOE07jxk6RpOanLx23A88SIcHIAlitFhK9ddvvm21Nn91HcjDO21xI6gUh7K
YivFIZEPLP12L+HPxz+kfUnu5le7nCbozJG+j1HqW1WiMDexyNTyzeEDLOmqpG8lD9nfKVLHe1oS
65G703pqbaeA74zAW/xAIpTJUordCYSfW48+/rwIqgUbLChQiz3zuCOxKZ7Y1XW+AtV+GwQQmWWy
jgRd1pEhZkwnC6cHozvY15VCMjEHTpu+ws0UVnZ7v7REQ3EXmPWRbKwBiWEUmaiUzoiFWt0zaXV+
OBDQoXHLhgUhEh7v0jSX01nrOVT2f2fkMWCnKQj8OFGn95NlFO2dUFv01mgzG02e+jdhRjkgcmEe
Q0t295cIixZXR+RR//963lmQ8L/wiCM2oQ3+6NUrK+iXfTDqlOWxQpoyx05tx66zwZPbmvv015kL
j7O852zcSbQf3doBu0Jw6LtQnMmVQpnL32QvqwyyzHM+pLHxTCCf/brR+T0qA7RlN4/ygr7g4OIf
qLfD9u1MHbTciNUfimyxFNS28RV8wze1Zu+g7IeZI8mIy726rynrjGVyVkMCE54s9ooIbTei8uf1
oFTrZjPZ3TTlTl+eA6c8aZziCJ/6/WoaQZ2wSqxG/yY2NIEPm6naMwzGEr0NZ1dR0oK2IuSiO7Ry
t4P1TKKIWVrsRBc/ZW37eQSYKvuMtrngPrEl1JesgCwtydoPTSiACqF4SwDk9dgqjDAD6LXYw7NE
YTLBg5BHj1vfrPv/0byFVO6+xmznngL9OGSshflxClQT/G7xD9blOuePOH0GJTvQy3c9sfNM3aRp
TLaR7YgyaNnrrhL+s90+W2qLMpwUlOOzlwJ+BH63jB6DU7GdRzjWdXgbYk86n5Xvcr51/p3OfkZo
tx9+GBAtl/gFzn2cea64mpfDW1TtDpogubYPydf0SsDW97AojBru7r9sXm/xeY0TmBoLHQ4i3xj4
D1W9Rnddp6kHwEIvj9+BPLnW9+aonQJYZzgVyajsIlJ7LP5KUnHz5qKyOWX4V75mDujUdcNXlQiN
Jj9n3QJi2aougnjo3o6dalD8ZSsZv6qomx+2dbCoiSgOBSGkbUC/21ota/MaAL1NXkcqUllhFdKJ
8uHSY8HrwG/VjApTK7f9tgfb/6CJLOS+0+ES10bx9t1bMyGJ51QMNpzmipcgig/BkTZtGr9yyqiW
iLEYcEpC0MfGhcZUnPIn4t9rUer/3aZ60zqV9W3WawKRKOkKn4lIOVTKdv7RQU3CB6MDTL9uyXci
Ql+om5c5RDPNadR+kmsMuI+/IngZ4WGV79xY2Ul5hd3zFKm8+h14/GcxmbhQQmF+fZJOAzp37e2w
+Q1AbrwgVc6ugTXWbOIF1zIxhVw13E4MCuL38848bKdGlYUls2VyHQjjS6+vaCmfLreKyiMlmzE9
E8ZSl+6nHamiEwXNdLLK23Du3katvkjVDdpOwgB43mPJ3utNyX/k8GCG4+2IK5drwKRR8LkjySlS
+MkrxmWjoc4P4HLCVZ3Ih2PEXgD0QpRvChmTyoM1Xuldi4DC9CfjRMBFRiTPNImXjUbsV6w2iexO
VsFnrQBtXg06eQIZfoXNotmcKCbNh99I3MH0oMKyl9UcnMvOAf9SOspvdaytl3GgOOxlhqiXnkFl
inNHvGSgY8ran1RByL/ILTNLXOkrK7eJdsYv8s2TMJ9XaYR3g3qQkPhD2lbY5WP7rAjRoY3wtig5
vd9O6HhBBpWrd+7MVPddqEFvyd2epzFBf53QgEBUrBiD7Qlq76WduG4VqkN1gAxUBi64S14vDLP7
KPTh11BxVPHGMsuWDIyqzX+MQG1aM9mIpHyAwwq1dHiQ2Lyomw2JT/1T6IBqSy+CB++SFWpm1VGn
7rvzBN0D7tct2XjzMHe/LO7hUvnLKo5mMkMgzutByeHu+GqyU6lT6g4r7zIUtqvMcw9swk5HlWX2
du7WwMa2s9YYaBjCFMgGQL5/lM0TaqxNCy0eB7XbHEiCTCkjN7MEmA/G0iQNBbufRo5pmdv3o5KH
SCE4MdESOf/D8cMhc4MC8bjnhHRip4ZXFeRbVQciBrwRU34RRzzJMkPUhHflx8dl3hbjQY8DQkmP
NUysldhn+FJ9S+5kAyPDJRSR5BPjjC+pAdODr5F48BdjrmF0j6yBPWTqkzsZnurmgSO0nmObbTy3
OZqK5+2hQ7jvA80ixZAr7Q0VZEAaKJrN3ZvytTX6NzrYRj6kR7UpkHpzM4XcdtCR1i91+W7gqoFg
DH/a2AmPu61Brfg9NvMtkYDhdMcliPj864iAMzSI7ZnNW7uVlTqlErbr4dLzONUPcR8OB+1jE9o3
LpF8N9Xw27UtGpVL4pTnwc6s1X120pO7MBnlxc+UfA1Skf0ISCSgMFoLXqzApTpZq4sXSai2gX0c
aEbY/VQvxndeKjxkZ2ctDo38uVZnLKRnfNon5VLQwj9fyEX/yYZ1iUmfKLUm/sSPUUKqhndbiN3u
3u7ZJNj3AcfP+pVgettjHZ9Y31LT6sAgoDSTXKQtX5VuSonPXBDvzTZ45QTTk+gdkzfN3qFdIiU4
h+BQfr1Z9Par356r9J2qVyalxDHki71MB/RL2FnpoaIT35t6XclAJKsEiJPNE6wAXSnBfOo77aQt
bTADptmDwLOFlN1Qxl647OxNs8v/mF/h3kF+UdwY/SSBZa3k6PdeOnIhA15BpP3whJ0aoK/CdUEj
o6Ihk96RIJqQSxl3yQxnlq280Wtq0ddQtNoojOXOjP3Wt9xIjVMcKDOnVb/3RcdkYkx9XvCkkjn9
KzM5dTRUSMNwqZvPqictQpKSDrAkymEhzD1T3wJKzYqPyL3CbGagkl/x9RZjGQdhvwOOfRKcA2J0
xMJiGgZddBu4Wr6XhKO7v61xqoCLCXSRk9UPxQDt4Z0BfrFIKDKYMjj8PPXqSNlx67nwGs1W6P6+
RUE72oPGVPuQ+fkwGhIsnrVFr/6cwgzK7RxmOTkrcgxWlNMqsreO4/PqNUrHuYpxTbWUCG5VWs/p
M/JV9J5vZUiYxmDWbDi3iurZcYeEv3Wd/QG+KfTMcCb49QawvyUqG83vedhP44EBEsx61VDX8C34
6gCrniePRlKOOsO7ITAIBPoCojoXdoWlpMRe1ikGuHkGHxMrk8sByUyUDoArogCAPOWkl1utN12q
4Upez2TlCbVt2mMTVmJFxmHHwtv2miraR8B6gVBjHrDvkIu/NfbA4oii1KXj+2nXdRUxuuWcv5Wy
9qZxEjkzaeNu4Affis7j8yEnqfEO1L0FTYHe7MMq/BdwAQypJdFlhHJMZQErtUPXvGkwYKMtIZSP
XqaASL1DvBPnqeFdQEpMacOP5wU3cMObNBAB2seHwF9iXqsarIe7pS3naL8ZMCfYO+X/HA5QBhi0
sKVAvo7BQf0kB0UzwrTWkSSHtWpXVer7a1b/O5MZpCWOJQl4ZB/hmzx1kDA5729J0PUhVbRDosZH
EsCXmwm3V6vF+D/lkUNvjucpLJL0wxDFfb+vp3tYsyhIcTEIm+NYXGcDrNltiiwUWtIA5GK3MMXi
oiqICp2yWP9/Co8PDLEKaF0gjFnMMV9a+4pBVM80uKNNqYgni0wqeA32fT3ER9KeJ4B1oSrsnK/p
trlAYTbYuGTNspK739DXBCCaEyugg1omb0sojSa2aZhd+DXI2sI4r3cRbkUKvs9aeLZlE0b7/8jF
oHdrt/F9Vpqi7eLl6EVwZnanJnMLNaHnwweprrTlp+XlkUG06bNsapW7qc9iW8wXELr1/M0/QvY6
08c5TjfHAZCOLVvP1ZBIwyuDbd7mFxb8z9/MAaZufbuH5yakRDtopu7uZjXp03Fw1ydfI39rhsr6
yky8ymo++JikiYe/2hIIa0YGtN+i/K6bfgbv2PPK/u7cUjih0pL3AG0Mi91rmHXXN1UKdazDboCD
KWboEHMEE3ZgmtqQ90Kbo6Rmpl8rWsgdRvibJSbRdOEQnSBF52x53vTGj7HV5gWBfSCWA3I9xFD6
rAnlSupw3fjtL2wAog1XZj8mQtw6XX9G+frQ9Ety47vCHEpfELZNaWnGANPs2F0gO0RwzaDCd7g7
YENdVUWEuE4bfYORPgYl4TICEZPCm3LH7EpsD1YBinRaAHhrEL8jnMhlN0Vx4cINWjft6he90hZ1
Qy2QWmydWw0gdpUY4SUv+zhCWQGdy7FnBSLGYaHZlf4Hegx/sqlfMbLLMnibI8/cBGQgZRPSFkoZ
maguS/Va5QqdXSnUQYgqW4DyM8NnETYVMWWugdVnP8ROoBhsyk6eVzynwCUGjvf6NkiK5f6CN2oM
32d0k0VhoZpVnx89PmXEZinCeuPorkHvoipv67gSv8UyhfuCch7XlwkZ9jMb2JC67zv/heOoGVjb
DXgqXsARLgxQ6MALk9KKUWm8eY7ObMcZkaBeUY2U1FsvvUl8NRBHWY3kSKtsKJ3BO/BRREvzkeMr
SQbwMGub+7sE5nXPQGQsz402RxSez/xsc3aZyQGLV3qYkdgOlBjnvxuwHZTeKsveoDDAl9R4qFpS
JfBwHIu9um2FvJYiUc7Fum0zO4xUJawlssY/FcBMa88VuPo+Y9QGD+L11grbHdrirKptQAOFlG33
89BrQsekCw1UQlW33oADjTTkgAxRHTJlOErMoNr9tzKGvf1EnH1V4AQk+/v6qnzvyOwm9g6hQuc1
28VC0idguHOhDXxU5msKJL/I/x9fvAtzx6ZvgkeOA/iY78nG/OzLVYLTi8zDfkATvmowsiQbhM1j
r+Hz790PujlP6BTbDqPIqADm35Jmy1CvYEqoniC18PQ9JunI/0kHAqd1aKVssr6626G5sB7oWE7T
7FGfiFJFuthW3hT9JWRJq5KMIEaFa0ue0c5HPYYfLT7+zQ16TrZGAqatRd9n7h4ACBXw44h1EUGC
K5x64SeaG7tztvSsAq8HEZry5sPZqblnDVDivO0MEvA5n0gc0S0tSe9Dqox26Rm9j5H0lBoGbdTJ
2a5Ue3sDiWhYZGBebdR3EQSgLJDMukdGOEQj5D+rTdMiB74IHBH5E8xg+R1gGeZYeu9TaVwrC+nI
JxxRzmo3rRfxEW56e1U+1pXQvbhJkK1nSEjOpiZNEgRRgXOtmL8cB0e2H0wyFqNbaTWpMmkYvpxP
PF8X3LTUDD/zC/kwiPUu1fUCCx4POTZ3TfWBmtFTyNyQN93fHuftopA5iT3j/DEMpvD95o9CCkMT
K6b4cr+paNlG9iHiaDAG0eHc9my7U8Ii52jcRI8hojCbg1giESlpJis0nmPintJqNesIHClN49x/
37F29DTn06GYEJcR4CNyduk3ZpBYO7Z50bLoVKq4wrfMX2XsSod22sfxiDT96Rak6HyJge0PzQ+i
sFKmuGoKyD+I4ozJkGbjc+zcoClhIU+xmmGIZ5XzohkZE5aeCc6cUhcSNWaUCjdcyMqS+gJLMw+l
47TlpRN0HqpFRbsZXen822VjP7yKaNTLDnR5qnnAPHMqFkC0+bBlKHOBhNIXYt7vAH/vLQU0in/o
H1it7bI1eYn1yFpdYzMqKB6lXsAEiS9ws4mdbPdw2zLn1+fwQSv9/vP+gK9usOmXX8tSn00th1Ke
Vy0dpm2OtHkAQ3Q6lh0daKbNvdxrnBzCvpkos23+9mZIeNKGGFArtl+1bizuX29xQQtR7ZiL3E0Q
7mSfYl8YCwha5HsGvHcE7UH4V4X9a+6nJUhTFuOoo8JqgzUX/PSZ/IUALmnN0oWgtk+k6r63AnEX
uRO3qegBywQS/PVv2s3WqthK2LtjkEr7Lb7QJp6FvETpWnqhD5pd8t+rcO565Q/kfICZDeB7xs6H
ebJ1oUx/X1JcYuBw2QvUSQoAH/uJfYqSs9advmoGZx0bxQR5TJdETHFypzG9h+ZKXeSwkzV9u9kA
CeVB2/CCEyXiW6p6lCaMLHGIJG96HFNMcBPJUK9RTi0Dpb/6fwYxba99xOH6ooQNCJz9ph8Hy5Cl
nYdzbq9FD7MWZTDz2YlyiM9Kq/hZ2cwmtpJKFdvYFwEzrLc4/Wl6B7gogqzuG3DIxsfh/8+q4IpU
5dAKIZgQ1Y7eG6bf236sy+Nuz/QUhpJYtr10OEC2mfwbIaec57aEsSEgEz3cuqaQQrqbRpNuMuwU
hmyrPTkYHW4ldCdocEK9YH4RYFXQ9RSlB7uW9gLry3zUcnUp8D0WTifGvgv3fMqhxpA1SKGZhCXr
IqAawbPJlmCP7J+uJpt9CST4BKgTZ1DMA+/7iCFCl89w1R6PC8V1ZkeSE0QhXG4n5f8invM5IF7p
ilwtqxWtOFpf2VfSFyRI4vLOn57Khf7oSGTH/Hk43Glp2PfB6PHQMIMpMeiG8m2mUO5x6lPvorPZ
aE0ogoFJB0V+NRg9VhRcgPnpDYKirBS/4yXq4hOYmxyvS5XImt+l6VPxnYHKQUtcxyKn6t2sbb0T
zfNQYh7fJRKn9zNFAQuhyd7b5dj567cZDXPOYaCsyzEhUKrmrEjVdDBeJzGIJsUzuf3nwA+kE6ql
1cLFcY/FJSxXFa5lCm4ZwiLXAo/IRteOt35+glF4KiZkjT9rDnYH1LNKl4fMlJ4opsQ68MoQomQq
/FJcYr9tsEDogzBaINph7yd5TmWDYmt8a3EQU7r7PQpQ2IZoPYLINhg7ZfhLJJ+NYZBh6Cqc/f8i
XGGiW9/P1oDq+SEFf4xbpPTFrSZ8DkhAqA8Hos8lCPGzGGNlDk1CPDAeV6wTOZ7bsJwHxQ9MOQ2W
cJNGY43rX3Fa2PhXkkijoNhj9qbJxYwnOD7+HEiap0IyNFJvEND73+RQLTT7QDKAq/2QoMeMAI/+
CdCWiKK/1qeJgqDhl5JGI0juKFQE754wiH3zforQVdK6G1xBLaegaMwwv9xFYdBNpBxgCQvdizjo
pzotSORJ1CXGIrL8CjnGicbP6acKJCjy4oxc9CuqCGkEJyOOB3Oa0d9cbjgJWVsRUD9HxeX1PzED
cZyzi2AJpf5lvbt29pmNfsoKRXC1GAtLH5D3kSjDRiUTzvvmBuMMvTg0cD3ImlBGcdFhhfdvSjRU
dSdy0u2Q0twn3eizoHFvokAaPqs2axQBnevTZG/kmMU0g0KHVXNEJWOhdoW/Tche6juxFuLoKofw
pkhTq8myPQIis9uAWyeD3hrDZVcS/4qvrVySZZ4ZKPKWMvhhCh9Ws/UHSPQu99rfU7BcVpKWUlB/
wo7qyFisC+sXRQsnyMkqX9mQmISVESmwbkr2Vx5BWiWcZhhviATOfWqT5Q/6Jp23UsV/UG6n5p/d
20ZZ9f3KHE2I879Q+q+oYgxVuWMv9n7Ji1GiXi2o/fk93mtdTsha3lO0aBT1PSGenvxRZ29jY6ST
4c8rAL7CR3N3IHVEW9KJatH6Ot4ktdD5pBez5uYPvmQH6jOolyg0rkpjl21tAHcO8aCCa2aeIGun
QzOZ3kj43kAos1n3bidddk//cAmUDhfEIVpDc1IDCD0Nn8JhQ9nS6qVIzP1ky/vrnDHB09dKojdr
LVmVH5CPkYHvXGdvFUXTJ9l+t6LOXl2OAG4Rz3VituVPuYSnWF3nqlT37kgeB3rCMMyXnnUPBou+
7IKXQUhSdKZr/KuZZJ2amQFtB87pnLpx/279lif9Kub9zRyik7Bh3h27zNq4jA6x6DWi0WBGKqNt
qlcZecSzL/ZUgRTGOlHiFbfJt3jVX0KCmajuMDueh+hJ5t1l/m4sOjZLSGLb8NCGfYkqPHrkvsyV
D7FNosTlX2+2ZiB5FGYix42hd/JLoRyM5jf3wICr+MnLaLSmeG5SznXqNAyJPBhyr6Z7C2qYro/O
Drv1cPzlMYJbJwg6A+/h+JL9+kFsluIjrAGs7mmO/QqH//BDYD521VVZXiRdWMVQgyVq8rJ2sEg4
BNPBfoQggdZaboacYpXu/d+mbS8WjXil1u3gVbselv8ILriEkmwhwvFZghM6TX6ApAnWPk7tUZDu
21cPGsx33fs820nei9JPcEUtUlJ6jM1hyk5RPsazCmOc/RseSUsGW0t9emllZBklBbUrbxerrtUx
GsQRQc1bG8MIFhNnUqbU4JEIZ3GzrHHGTtrDrowDObTkrVhp42OCcv654UDwA/qr+i9pVVDFL8iF
yWtN/kO7EnBTtp4NKkwcQzDN1j7JFKFoJRGhLZRJflOeay5t82jaLgp1CJtY8/BcmNh+r7skwxsE
GyvxyC3Fh4Qh1UFut1MzUobQyDp/nbWKZQ/BjNTH4viFn063kYMAGTWTt2LeKY9Z2idMuqaKHY22
kzgeIxEpT4TI+G94RhiG2+nOSpwrxKIBrL94NLCQlGWJOUfApEjMkA4pBv0DkxyXBb5SvvLmNC8k
O0pvL7u3oWCbCyJ4P9SaeyqOK1P4DTc8y2/cQx2AH69hgsulW26NwyxRFxwNw+t6uB4Mc0Jcashw
47k0fGZO5WQID39iEfpz/o1Lii9l6EnW6W1XJ78KtEOTKmyf/HM+/XfQl31wuhps/C7OeaG5p3s2
39082a8jHb60gkhklLKaVsvVJZFIiMyHpQJHkUseoldCL2+GZlA7aC/ZH5b6ZuLC3U82O++3AFc4
v+LZn2LgF2FnrrA7Zqq5Hlw/dH8ewdtP0pzbEvkJSpewTx19Xz+sRPq8ImLcBACwjzGr2mf/dEub
/tnEiBU+bfR4q3uV4NKXd2QwwMIEtZnJ9jWfp/LBsTUvfDwtBbutqDJVTruEzgY4OpGlRU5+lgiq
1OMZgiUdWGKvuRHOX5utFinHdSIRIzKSf0tPySPNnN8fOYVWzOfFR3LekBtD2KNRFoRmb3TO/qtq
1dblYcnE8sHPmxfBccEcXQmK5Gb8wRATtP/oSpY8VtB+c3Mj2zSDQi3FmzgdFBBanGpNUIn5BM8r
8xtklD5fqaeLphCefjK/0RQyoihG1IR2Rwvraa8t1xlTR+Y5xNzw9pG4FOA6vH1NFp1g2OjwxNU2
t9qu/JSks06cIAWcZWiyh0t3fnlpZst2HeHRm3IlZKVO9cdY8Gr/cULODrfz7hrMroD6vmt8beO8
9HGWrlN7xNeqPd3nhlMdOeQN9TNKwN5fWMa/1bAoFC8BMm3ZAQDkhb7JV7qQ/JbPyW5ao7h+dqhL
fAfxfejq2r+vOP2qmWcb9CyC73l2tN1sst9Qsurv8Vn9hD15lc2kWQZdM4Hd3Mrr8uojSkVV70ti
+ocZLcBpMOqgw/XvoxXc87vSWZm1iMfLlBlbKDWi+f1uEa/Rl7cuSqzyplCmjfbjFXhJx8Yg7c6y
+mNUBHzNavqgLolMeC4khs6Y8i78iaRbex4y+YkugSB+oQbLoITLJG9aYfR23T1lXOdsgSD/tZ/1
JgcOlAEnnMdqzQMXAbF+KKGPDVDBw4X3ZLcXIryeFb0Ui5I1BGVTnvN3AZUt6l0+NPIHQtElHVH4
0MM9x+gOCraU9zwY3fmxTK02tAgH9FxGFwy2H/6A9gWiG+T06A4/LWK8AD4AUsrGwzeaMO8Ezugk
chhi1/2x/Wg026vChjBvCCvA/X3nEUB1tSkXr+d2fnlmJv6jI9bmaga98LzF1w3s9xjaQ/90YvBL
sK0iH/9Y+HhSTBXOlYr82IspRnr7EBkXA8BxBHDEqhSqytjh7rWaGIuONeZZcLTN+Ytt5ZSWTXcv
icdoO+k5HcRqGhAHBhu33Q96Os+2YH4HyXM44Ecn57FqhFyFLWX0daSZaQhv8CGkKNvAgaVRSu38
j/it2E3Q1wRYb9fpFy0V7f+zzsEJbcpy65R+RSelxnxzHkDWV9L3F12QsPnP8wNyr7fdWJeu/WO6
vpmIPASsTzw0SmpuWYaX5OTI5IQCXB9DN1RXW5DpA8DuhbAHnRrB5puK+yDZjGdgcByLV9Tnifrv
rMHiosOQhY/9SlJvR8Lcu5N5s5xBRZbqrUcBIvRRcc9No02BCy3/LlS8GA7vw0RTV8zFf0xYFbXP
fZPXZPbS2DHQYQq66F6Eja8fOyu8BpOnm7zzuixFGU+ewRDll8feefIkDUdVmozLBKQxqqzMSRFp
BaAGitDuTWQtAUXW+VrjD3WvI1lvTz/iLnfD3d3apZl8q0tb9gh1WXgBv630kx//WkNDz2XR775w
hmGCIHSn2AMvV5VSdjpuutIK+GhPSejwrBu6GErXGhG9cvps4CIz1aPLHdvd1wEppoASZT0fKw+j
Ig0KWwVN+5uRR9azeHHcFubs5MewBBvSkzh8cLB7DZ2loOAGof1W9vaBLMuKWNomdhZSiWQ8pxRB
MVGxvci+lZ00wdaww444Q+muNhHNMjf2UN1afnRrgYv69LOqo8sKZ84N7RzFtS43BM+mV7HMhUJo
YxlCvNgkZbdPguWW/cq7kCTJTLi+FJqPEMVTSGjvJezOWMXr7x9YOdp9gd7Xi0kbLC1ze4LRiC9q
zb4FjTKaFS2w21MT0JiRyMIc8LArEpUwhxo0u70bsxpgm3sAIqW8p5y04sfjRBk9QPw1+zQAX6FE
FuThBA7K6INcFsXs51QVTz7ZuOUeU9sgqKgte9F+lGOhw8fnELPSc/Ff7+CxY+BbwnJVzQYu/LOl
hKoHelIFl597k4GhvwoBUanFUfHDzYEpt8zCLQytFEXOpI/CLNMuCRx2Lj/myK0WMnkPlV6uCnHl
lpOm5GiIzAyfZHcorm6n6nBEarzVpvZCylClEvt2ktw8i0dqa5JvMdOElQzoaqF9wo/dUbRfGfAi
3Lh29SCzL2dxy+QxBnJgmfCy9+TpkylDJ8DXoZlWEA46PgkvPabAiGoC+mzXXYBAmGFkNnA9JICd
AabpBcrCAIGGEsaGqP2IONkCaWzxWBADMSVwJV7+TJNaWXR4wixZxwU84fYWsaNI90XGmyf7y12Q
AmVx7kJptDCtIxFfWVt8ZghBUdJqK6RCOLQXkwR2J0TZ1eIoP6f1+IfETla6zDwDqqG3/mQt16+Q
zZRu4zv14aKeOsNaNKC0Dg/71WdscOSwOFy3ADgoQM5vHJkxh++0/p6iGVLobDicalmZ+TQM87vH
t7N7lFVIokyNx+emrJlRBkSULZtnxRjB2MsMFF/bW8i7apFvUQ8kn222XxRPxcCO6GcoAKLMJjJx
cbOQ6ajtatV12RxaGQBPRmPnx0DNcDrVUkWOBd62eHJegeuqGN0eFgC2V+UYd27yNzMwPTBIz9f1
zpMUIAnrVPRKLAhB97lBNsIlNmpVvA0l66ovIz7CYj8/RdCHGMnaw1ih/7rT5KxvczlIRCLcnmDC
JIYQjmNIpVknD9c1sN52hdUNvmU40ewAjqGuvxC+2GILqLSzdMOtk7tHELPBasgPAeZovv+gFKhq
vmpR/eNgPgTHHm11Y94GPq5Kcc8tnrksReK1DxmPWpeDgHHApagWXjN/BwesZwdtjkfNJiemC3dz
k5+qJZ4XXVCpDSSms5q3e9uKBfDKmf7WhkhjH4fD+4BgpSJY6r505uzqeOKDmIJpsj7GX1zsTDOA
cmwrH3zlupdGcEPIS+8WKoTZj0NksfmiUDjV3FBCbdaz7GaWgJNitgEc6OI94/DOmqiimL5oRys7
LNKW6+gb3bqAFxQQF6gnLR4mhlczV3LqoMXTgXYMS+/FNbpx9o1JjfPM/J5iK3oALW7B+QpMLxjm
KHscfoomIzUevT6nHcNM0bFmV0R4lRi8klUkecTxMj6LgsSvEGu1whXbDwEkCocow1rKjvlcLYt2
ukN8lEgI3nFdMSueKYb5qPZzPNRY/xPZli6bXExLY/bYOwdtPG8giB6g4AB1d5ZfLJet+1td5cfW
dkSiOIYuC1tr78FLX1/IpWsQM6YNwTnJq8ZjViPxAjx6OoiKOrZYFL+tP7WAPOqtYfjv7NspJWiI
oBwSeUV6dqQhPdlXPuVTQPs9QpgwUe8gGrnesbe9ax/Sdi2nnHfJlj+b0Nt+b3ObNpKyPMMRVu2c
cXUZDnIpK5asI+nuA/fDtIRY4CX/jvR23nNMXSm9X7sRnEsjue5E+sbq1dM54SMpg5v6PRZHMVi7
Y1A71K9Use3kPHXTTeA5zTqAUNnK7aWgFEn/2wgW7p+ZUjnoYzTR23FBpGasXptmvePiFsEQgQBb
XWUlo+o1wKlNbWfrv4f9wLJ6jkZ+9du4R9/DT8oLYKgpzgubH/RTRNxi4rq6QpzBpco3tP3kPqSn
xBN0e8+rQ8vlKPfG1JNlScrQsRvgJQ9EfzvRQ/ovxu9VOT067nJxzakJzjV2V8nhmIiBhNzOFOsv
DVS1CdNxclenn/mFW+jn9sWLz9o/smazH9um9C+DGcDOWqEEqeDhi7o/8ZSKCZ7Vqk8qG/dRYrXN
or1par5qtzIMn6liqOlxJcyRDufBeNM3yLur8Vrk66UTewDwaDcZOPfGzoPjth17uMzLW/48PxF9
rFKxXevgIbEWqFMwb2ofrUTiAkSvGVXb+J7/JbdooN3A59IO++nuco9hKpLwtJNiuK4X49IzhDrd
wpNtL5e/WjAsLbpC3hdecyH2khL3MT7gCbcAeAs0OhAnY3Rqy/p7vjG7lVQ07eURcDj5luCByq2a
+ezeFr7vUoaKGxxbMRAcIv5IJvNFlfTbUnblWXw05p1f8OdmMtwfvgZOcPJ8C2guR2SWgKhjeLVW
u1CpZqZGP8geplxMfipPBhUQn1wpAGvunF8QQaEzdMtSNHxuAioW0fm3T/oSZ13fV9lQhKqhj3cq
+4nFmEIok4ae1izJckIgyH39qh0yts0wqJQ3hNOC/bKA7Wjx7zuJTk4IuVFfYOoIV4Pqda4PV4Pd
DaZTookFZ6wSSAM6tOiHpRaE43QeDNU6piBkrpznG3TYnpoqxyTJUCeMxTV1Y3T+WMIwy/t8zB2x
EslRC35xNqcxtxaTB3HpRBCJXPccqkVVw18Pdm1AL8FP0+92RZZn1IVxhiJ9Czk0ouPvniWjiBA0
k2aCvQWsLMnma42hlwU6rnSph8MHQhUVktX0ujmd686cs3HRPtIjiTRUJlz6NLGaAbwLWhZgJxmu
Yq6g0ESc2TAhke1RNmkJpjRru4tnoqHkm5a4ek/dMYHlHV3CBLgxbuCSWp1Y48ywJ4W0K3053sib
IXQXa2Qlu4iJ8Bl9uhR7k98XkXWVDsDJzPDr78+v86Ii43jhT5wBGGyOq6T5hBnhhpfqLaoZ3CNc
PNtVdjYi3H5OvAeSdrrhFCqC8qJtweKpya2DE+jClYg+FDnhzwsY2NhI7ZtKmKTXMShlaYXcbwCC
3qinvfhKSas6DmAyowDlajEs2C8+uKx2nV6JDJyIX630NIJJmbH8ayhKFCx/sChm6pQAjJBxZ7UI
s9WSUHqwuT32oG1r7tkpJqc9cMSc+U8whi587sXfsYGOta5BuTe1XNScxuGB8SZMKn+h+asqqYOj
/xsm+VTqaX+yL0pWBwCZt4GQ8SC3efv+ldyP+jo+F52WzypcjOmv6dcP+z5W5qnJ9QAgiK4thGx7
bhfOqKIk1Njn/4dN+glmZFGQi61HlK6QZ2zRhqWU167GS1ZaycLIoRQKd+Gq7DIuTMhqW815wX3P
0M66tzrm5T9EV4vnW/LVT1Xs27s0FZI/ITWUbcbmz+wpdXOpUgB+D2JOX2fYwVZ1baZkgaZxCJ7u
TJKfZP5Pwr1tzj9bx7uYHz1GpKB3dwA1/01tDov8ccC+y2+LuGyovOSCRfnij5CpR3Fj+r4B33Lc
09SIeRms70RApdp1Mj8VJgt3GX7GJfftKl4mVnKg/X+iBO8ZwMu5aMfDNtrjNrM3PfBmv3PmKCvS
pEFBl3GiQI34PtCurDLf/hXOjnqNsc7LfGYMvs8mJvFifcY53rSRNUKukZ1IQQWvOmIiOt0oN5U9
stzJlLHmVTQ0be0wmfiCLHcMQlN5ePzCWR/ZG4IixnuzW7R6Ijx3YqJ0wU0Wcx1grPHqZtBMjUlT
Yhm6yTRo8b/85fr+ZpfCTKTA28c8soVaPXOskpajPXMXEBW66LDHARAKakOFLXpb3nac+Wm8MBTv
Pw2BHEm5xf/YYv5wes8FvXuetbKcY1eDvCsJVVCfX4YuIjL3g4waiGoGloEa/0j9G2cb+4Rz4rD/
NTdiR/qQV+xEo3JRAMP+YCIhiFgbGYT6L2ATgN1qm5jeXCBPRPM7mnsET8fJER3H5LtRKfJA5kL1
l8gynjVEk4Rr29GdZAB8rCANzLO6ISrs8FHr9Ja1LdCbFV6Z9OLn2i3jmhSiEwtAgAlGribs1WUe
YBqqoxtcnlwGcRHelcdb05JoMUjhko9PpV4voV7QtWnLt1NHgjaiS4uAs5EqqrjXpyNnSfwsVtFv
XWG8pp5YRAW0X7qrCiZr7+c/tDUJKJF4hTczhdx5yNFocKWJ+xfzsNo2kn4NhSsHRqL2c2n/iu2q
Zj56bfnolHhqVG/PEEHg+QjoTwqkvJaj/dy7jafAt5Gqh7xRzn/OezxlpaiDXfaJ47GGXNyorX8N
DxFg/bU0Hn8Yx9ftfJ8EvA/3sZjJEF5KRqgFeK+LSCB+jn/b24hY2/ZFmfPgV+rWj1RnwlEE0eKz
XFyQKA0cQ8O/eZ9YOebfq1WsH9GcPk7izOTsza0XfN2838cJkPbjaMU3j2ZfIjDHz1jSgisParhc
nl3BUrzZeh27GkKxs5H5rev1rfZ0hD4CAXYS3Op8gEzE4W30lgPscqrlQK/YGgLCToheft/HJCPj
6C0fQy2W2DE3qXZ7VX2VfF8SZI5RSSvVpg8/WZXtTN7RZlPMX9cwqp34lFPYndxPrn4ufcATDaEK
SrUgGgHP6a10NrsVcjBuPCnxpzq4TJAxAwIZxWfp1Xk3JpX3K7z264873jWQ0d+Lk4e4NdbEfyUz
9GIhS7TqJcGATZK0FHndqMco10odz3Nll1G+W4tPzPXvcr+W0ZD0mhbQBYVNmnyjvufJHEDfbAKc
ncipD8XxHy9FPsmMWCEUnBfOKNZ01Kw/69W/Xq6iyxOBRxN0ALGK8ZIFca6aaA+3VOmRkW9b7ZpV
0bvuPdKU8qoTBLUT8pFfw4N3IKfH8yfKs+CinkL9MspmrIdNzKerr5aX4dQ1VIPbwgV3IRTsZyYz
iqdnXcg8k5fjySTpdDxLLtqh86jssYN8Z0OIEacLIUSGo8JPkz6AbOjsXwqFdByNrHNfk521Ry0p
JsR3W/slJQmOOHt4lROHeF+wy1SZJQ0zWcrjYAI3wD/l345LSlDuppwNQCjqhfERvxk3hzC52lUe
Iu6WBepJaUn6feN61KSFtRKdVgQtckVEmkL/HctCh+CKuiesyrdWj6Cs5Dq7BLMsEcXBMIj6C+c5
NZTubLncJurpaG/mydJqRKaZKQhZNFVrKSAphRo+YI4rToYml9V4ywDxSXm1kMtXJIX70W2qqg8l
uvWrtVK4B9IeA2aBZXODHaLbb/hyRFLCPWa4j6EDEQFFvMJaWOTTzUQUQL40061ITvqxMt0V0ANP
ZRvJy/AdeQJUbRnYWBz7tjnOxb2xHymJ2IVQ7Df2wFV1w0aiPKL8ytUEwEuvJ4dFG00x7wQ0kmJz
S6SlrmiwyVdpa5MoDmb+ZsOlrBMZIokcbpsz6GDooXOkqm0ULtsdV8dwN8GNHRuHuTR7S/jmPSMK
2qChqIDfHX2xutT3PauBdfoFvdJeysddgTdLmDRa8/0Ef6bLRIs6EmUOSOfsy/8m3FM7QcvdgSm8
86FOKmTW425z6M7m8dOU0M50AcS1RRelTfVf0qnL3Yvmyyl9uhd0Xyuj3PsHI3pYLFH1GzAQ52sl
sB9IlEqhZwITKwtM7xuypE668eWi/ua4lxCbGGq7OTKpGLYMeOJ4UETeVbXtjHwvjkeIHwYmH80l
t1uHUcwZePak2JwLvFkiFTWS0U5jlxwaXsYZ4ehYoqeYvBOoMBj8jdqIol8vZ7uZS/OCPJpvuyNc
/lBRMwivw0fNB9XVNZRYUYo0D2I7QO7McN66JcQCTg9OqBl+x9R/oAKELJ3rmUipvPH0bbgx8NOj
mJsDvBVplBLmTT0rwcNqIQRd0hUuRBF4ooOsw8P2j+rGlLVCsWKiGhyOoG2kSGnefoIZB2GQRHXi
WeKm4Ytd3RUs57iENv+TBGdlgKDvuC5Ky3VC+3A2asv/DtIY426lNncYc/emPtuHq4VNdmFH09jK
rsUeH7cP9U95WthPg7Nmo5yNfi/Jy11dp15q5Qjcifqgkbi3Sd4vqxV5dEfbwhNrDjmMcyoAjxw+
Ysjoj8fA84RDq5kr3XU7AxVNIfKKfyjEk5eXh0mMV+YA/PHKMhOtqNJoTXZJwQWvp1i4QIuENkUt
l36FbnizonkI1r/+lm2En9II0mIUYJB5iJbTGkGluXVaxPJoG2SZVwRqjMi2AukKosHMwiwDbTMo
F3qTFpwJ73Ztb1PF+SPcHYvjczSnz2HgesAtbRDz/ruHBAnQ3S0NIvM0vCXlaonB2EzfL5XOI85T
2GN0rRoK3VVN2NGHa1XO90gpsGZpSVuhA5eDnO1EgY1SXL8r8EpdoHJ4fx0PYxFUU73LoMaaqa6Z
4yhkPoRibUskY7pGD+yr7A7FPb2q/PM1ZvneM9FIO2wTgLxRCGPUV3n6Beg77l7/qsWbL9UgxPsc
YzFCpS5J6J+f3Jr3r5Pm0FN99fC1bR+gtb3z/fa8K1Riv6RTw+ThDs8K3qKhZU32iap3r0S6o9H7
4l02intS6SXn4JlrDWdoIyQIXeKrczOrQbGt8KfTaUYa1zh8mwvqQjq5laNWotW071hFygMsRO59
mmgF1fY47GMkKOvLo//GqakHP6/vye0lRIuVF2YUzdMn/Y+RFJtUm4iaT6F1k6nG60lHzDei+vTN
BGgKW7ckfnPs7x0Sa5so/TmRB8h6wqc6jyHGEUsGaMxbDztrECFB3tQndXYJeW0l5eTt5eNHMbMG
kFp4/7IA6c0CckJdnWzod4He7LBjb/gntStJEhzDWb+gPSozsDZuQdxgphkGhBdfmm7//2O6+B94
36p+P7y5UHtF+BeoXgJ1glcXA2O8UjhMErR35IFJbo1znW6sOPT/P7m0nKBvMpLznOP5kpP2/iYP
7ht6FI3UcfKy+wxm75vojKr/xahJOKonIRQEjU9oBEXXg0FO5DUuKAQixEhaMkWuIFR1KZcIAbio
dEwySfVeKXOg9rdq2YEeRot37jDqtmFVzFsoYyUNDJmK+939kOVHO4vnqdyrLBBHFYjQh4sq8Q3f
L6l/ds2FVprxKLBAjE8lUl0ayroWBIghg3CQ90f5PiEOw9qg+K9mmtTdjlgL9SxJ0x5FT+ZWp/aL
Tfs3zqJIlyJRoenY31mEb8v/7+YmyxyA8PTeTBhUleRV2ehixhkgJGisUyT2BkClEsRtuXEemptU
vJydKYfRIKXvcm1dnz+SdKoBzcibIhqnNKVLKOKOxPkjya1Sse+WhoquJrg1y+txFRu6hPjPMD8S
n407mwajbzVCHqNZqKX948GNDKQHpZgyBO2FfjihtYOP7LS/ts2oYPACMn27/I55q/ITue23WJsO
G5/jnxGbpcn3BfCAHQJmydXxDxLi5cPZDrnmJc0ap84IXsEYWwdMKdClJ8BMb+IQYFGvW24kiM+W
+WfBIPcXsIfE/qmjwGZIiTcjB//vpWtun3XRiLUUoUwpSYp5RnUXDGcYr4S/HcLdmq/PYzDV7yAj
xgESTKWTsqhTYrowJS6Zshf2OoOhZe5K2H7ws6wFqeqbDSqK2vAMVtRp9vaS0njstRwyLQtXb/A3
+FVpExORJVQ0XS4Q0ezLcMhwbNY1YMWFV0bhLvAXko2Io2HmYaPkR7Nzai/8yShqzGXXehhJS6S1
82E9nvwh39Ywmm6ubC1C7Yyoz+mFi8onVLvshwPlD45yNV+DvanCCWiKwuOULmoFJWErnmReyNV5
kfa9J/E68qyl7J7pFhRO+lics+m+Oshv9CnIBN9wjExsy3mx4QHdU8d9kQN9Zzpqc9ixhVWDAiXw
UjU/GqqIQRamLgCe/Y3MwXMDUYEdd68xyFOHAMYUgbQY8svnNbY4yLvc6mU9cWbbYEtQNo2TXJFv
n77BmZOqXodN8lwqtKzT7d69yzLpAsWN8pZVqRxbl+m62KBf6/XwKrTC2+yXYmizR5SVpb9hdH+g
QjBUdGDROTnC1d5jmTIAwA+Lrzh4EHwnO8iqpTqSePJMFtZnpoEz8Dx09BDm0T/DWSKPhCWPupx9
TUiKVdWF6ankH+Qe8yk2V66BfqP6lRdL2VPa0yra2SmD91VU0tJ8pZaqs+hXgk1dI+sbthFix3Hv
acyqx/DZ2gEw/7MljnxHPjlDJ1mS6P0tlocvl5TGVlC40M/N2S/MZ0tGi4v0ZpUdV2edlZO7F+Gb
OrZ88DoekqUctCcU3Cy0lEUtvdcpQ4lrJCc0lgaD3HGaJ/cP4u4mV9KEl+xs5dnwfkJD0h7T+98o
IN4fl5+GOJfZjFuMEnFs3WPJDMiJrCGzxenMWZXs4Iyr4J6f9nngHXDMyWaFprKEkxGf6qG3itx+
QQiVJEK4wsrkqPRLWc7qPNq7X7ZFN6LGfDeuFtEYY9sCJds5Hl31nXAf9uzN0/D+tdE2B3HikIcC
C6xlSVm6SaneIt0RRi6IEt7dro9EbFNgt07erYvqcD+TlL3drjhc0iHYdg5GJ1U1z4fjy+yD+RGK
6WSOeduWVpAmqeiCXmrQgU2/ZaC86gr9svYvwsZlH/tRCXQhbuDQoyIHEqM46ksScuVvEUeUUqy1
4Q2RIbUO73sgq1DXQagg0jNe3k8DqCwAWPCL37ph6yW9OyF1ZjLOgYpF8oH16Ci+yo43tsybT2f1
RD1X+zcGDh59B4TZH8uUXL8WIxcetUYTDrvWaBytozyjrXzLGTL/ewYckfntAvOl59f1fgJsZRSZ
iDPV1i1Vr1bVqFAkVk+RoH0XhYOiUp9uP2G4xNIC0zYRG++drceLKzk1y/1b1LJBGwb9c/GTo3TG
pA0l50jNCDfWny+KJy7d1/FrT58S8oJtWNYfMWG5E+RmCMeRTnIE+HdKkt/PT/aTEqMqCA+/AZzt
p3NydXlD3ghfTfwmzCwcXsybje8kouJOp4AlKv2xkVTDAA574vYRX6zXs1GjMwq+ROQjfSrShQ6j
me5sXbZhI6KmMEJKl6VULpz2o5NfjUPjLtayYM/jX9IjQUNPGKlnvkSahnQfonfcLPtyT/7uaGp3
CfErze4mr5jEhIvDhf7b4v95yBwmRqun1Tcmm/72QMXQoZaHCLYg39GJ7KFIgvebtFtS+H6UNMY8
Y9iND5tsY2HZVdOK/9rWPeoflbtlHEdMpQggWCWqYeeGyzzI4axJYe+/7GkA0q0xFReZxTwtQrIM
PKzNIb7yCA4UsVjfgvMauOzaGGAViSaM/G1D/7e6SO1XSCKXA8W5/sfkcr5tKGZajZhnZbKKwieG
m8/qTIzzdnszSGQKel8nktuQfYonqw6Nw9WStRCXs77MplYCX8DucdEGg9PxSl/iNQfZCfzLV/OP
sANHBwfbXrqfgoVL4aBQ4qIBwY0Yr1SmdbGcNUcWtVz/aDpo2QvQnKd4BwbJCNYswe//v9Bpvci9
Ur0MxcS18Wyu9ergmvSoTn9/QF0PtyJsbp1I/Q2BEZ6pMfRMR4pfNRm5z5P6IlgGvABt/KZRF8QM
jGjFbog52/dJzTi7g8NcO15KtDR6HTq3St+mit4c+kqQ0ljP+l2okmYy5vzpSlzhPCzkJMK4jZkI
xmX1Wf9+z5pCD/aVfMOih0IILR0gtJt5KeWB8AcBQgoq0E/FkBEWa7uGYo8kaQeYZZjtY4Z3fJ0+
werS7LsAkbTEnQfFCVhY5epAqZGfR28RVsUgOrtj5ySPqHpAo4o1/Ao1gFrfQDF9R7a1B5sq4PVk
X2C1opWBvhj3JEQfG5yJwm0CKQ8kEbVPCrv2njC7BZZrXspmIiPt2yXnGNSPIQjjs2BwxPnbD6R6
FoG+CrxOgqPTNMGBJmDHln1/tYTaE7eu3NP1I10wFlAR5ZkbZja/czVuhfwS84smkJr3Wqq5gSUd
dE8Be8uzT/gR23RRgSF0DeusoFUz1s0s8RpsWeNjz7EZaV1gMLghAiSvu2ZD/BMy98tvt1do4LjZ
j9lIwOgKwEMPB34VV6bZXIivBSIxaBFQU7kbAbw0c8CGbT5lMPCKr66P6rYioZRlnFidZoF6jhOI
AgNY1TQrv5VUkFc0TV1IVJRlIR0ZuS9buLfgzLpFYyJQXuADArqnsb2hVF6ImhHtSIhPu67cUt5R
WO8FYB34VwiKXSl1DjrNfZDEZSg7QX6fIBrv/ec+9rCTUKB3MmeCmm6QttJGmxb5wpPWTG7HLe0s
Glb+KL+a92Pv4svVsspvVuv92ceB4ZOc0CxI5YwaSylEKh6olWjgYNOq5hJUhBleNkGlqoeACXrk
4CvAmgRQxVjYX8Eg5T0FI6CV1Y+gWgbcB0TC7biiskYYO0AZO4yNq9f+UgbiFyZHAREjk/tuzy3M
tufZ56v3TuogAUhR6n+7qUXC3U4ssXzLsxgcuiilQlilUoQr9qP45tRjbnD4w/gw+5pW7ci1wb2P
rNwqVBoQeW9+/lR59mDpm0CDcLMFUA0YZ9+c4hLuDUabyzRJBVTS1Kd3KdZy3+uFiF2MN/teVFb2
R4iUfE4YLcN1J93UsXQWhWdPU2eIJ4PXyQmzCzaK9IsGQO9W9+8TNKZNZSm/j0Cnj0ANtKX3jovq
fvKwqaQ3hxseX5LAVvxJUKEWouoFWtM6Lu7UP3X8k4Ix9wL0ieoOwKdh4x+DNtUQWrtVeqwTamny
L7ztzXBFrBOveqoZeEAo6Vik5HYVlbHGdB/8TrvU9NLwLhvAjteHAlMgCBejh7dmeTv6p0RhakIw
TSlSl0VajALnQ6tYw+e8BzsY4Kkl31widKWN27HdQxIeO/1pSy5xbiCDlcyOar0zmgsnp684arrO
HkxtHh0UhZ/pwKIV0Q6uwCsgAe6OaABKTIbWCY1b8tA42nkHV+1jUsU0o6nhkbrBxxY6foI4duGK
GwPbSPlAe3n78JF3Ebcrg5IxXrg1pFvNI8ntVwXWzENcpZRB9NIkEJBSitv+cbEDvpPSWbJbkw3I
/gLJnoGPTr0HXEkVrm3FS8cohIpDwh1zhBbDPCbnU2G2g0aWaCNneGClIl3zDTVI4Lty7sz/N/00
/+RvqdPNLOZK0KMxdTSC12FG7TYQp4BSaGGvHcVAt9+ak84m1M2vsOEf8UtFJr9Hzf0+mICis6YO
aRIsDHhkmje4c0hPeCZt0o64UZVUDCX1w0Q0HCu7Vq2BfPC4/A1uGRgPYwKH5mxP2rocR9pPpnyL
KAMkyLrHiHp5vX9RSR7Gj+CSW0xTTOKT1DePmhImnAwk0EspP2VaIGLTcof+DZONwBYkhxMjgVqN
DVNc1s81wrinruQni9A7GlSiGsJE1Wqq/JR2J6x+jF0CQPMvHFpwhxu45tPAgaGMt09mGvAPBW5+
GQWibcMguaPVNVEUwl6SwLKVOylIMx1LEKOTwenT9K12Ul/aqjoSxtOn0mdo5zk6qHgw7pyGkliU
49AvCFF6PxN44IZkSLbJNdrN2rftBk4pRoFsHIPb8yMPowiK1c9XXQD55gl6+f+tZlCJxZCVRGl4
8rk2AMc0SVfrPfXBr9wdpFcfKGMeNpqVYIE1gYrG45Z13+HnDtcrDYPwDIC9VAFITqtxui8qoMXp
bQWmVAnMtKZ/c4i0ys+VD2LJdsOLpizeq4WTTxSKdc0+j08ZxczIUMVjQYjDDGyj13KSB1TPYrCj
YWIJF0m9+e5tVeQdIEReNuV/botQQzY9jucogOQbJFimSmWby3SWOy6DSxGQzJSI9bEEXW7kh9Gi
n7XLBc9r39fkmy+I89sobsS4jB5YO3tXXYunE0HfuAiNjclQWNplXBnUXjW3zqMSMwI7k+esllss
IrUAycf5nnM7ICfE/bFhIC0nPoGcNmGdqOUk0SquvGqRR8DgDhqql7RybEkDuuPWBiFRYivyVOne
EIGJrxQS3HjBBiLJIVBQeP1W1pHxIhlMdRc7n2r3Qdhf6IEt71K14tjEUIKkKhyQXJcTdcy6T1yt
kGJW+d5tknAFZQ2oXN9po/oMo8h8HYqDUsduS64tm0VymCvRZPGjICpAEIL0RGIJ4HdUBCohvkGL
GyVKqG1QNpoHioCs5gM4KJAoQQp+U78/FUGCJqWDgX/ZXLTfzG/094/vAAgYspX7gORd9J2g85Rn
iOuMJ7dfRT2Dkuo5gLjHNXwhLocm7zK+M59VrnVktWAIt3Q5WBap9YwJPHvqhxPsCn0F8Lb6hELQ
vG5oY02uWRrbkFcmYexlKQ91xXoo/Q4A9D+3HFU1D68ntbcmQYl33dl6oSimWxOLDbPeOXsADs3A
fgtweo2qyw3kK6n/Y6VE4HtmmwVNRWGI3sPz7AhmBcoFxuAWIEn1O4zuRYBFqhgXsFoPGOV9hv0i
OFdROqeuDFH8/ypyUSjN2Q8yefGY9AvewrcI59cYMYFoEkEq0R28CS4JBHrNk3LlZKsfol8Rk9HR
sNEmRE1iLolz+a2A/NnFedmGg44Y/LXVnoU0mnAEGuM7NJ9wtyPAfgi2Yd02bohKK5M3R2g9nz9l
OAv0HW/VUp/9mWrNOsF2e5tV3vS9kd5WBcJiGE6HvVbHsEGcmFzFh7ZTgoB1x7ssx++eaNT3nSiB
zzUmZAUoN6kR2auBWCgCJS18Xvqyc8RGliEz2VA+0488TJ4i5YWweH/OdNaLq0KAvMgt147KUq8A
xwcK65QGqbqM2ic7EysBHysW8eAayJ0//eiGSeML+XrSOdon7EUTK3ve7M6vh/JgcfLzBHRWFUwH
rNU+pjOZstRHPR9bVuKa/7ZTF6w7XXeLJrTl7IOwYH3T8Gzckwf8MZHWqrRRUhk30EnjCubNVUIu
nNxDkjNCQ2EHKxkAcSOxKGzX9c6z2ZbU3B9P/9AeU2ZyjZ+gZzfDkMYqjUpXHqsKjYMN3CNCJn7T
2yq6Hp4yEpsGOLBgP3fO1Nf7Tyo3kG5Rn3O0rwghFV3U5GBX6ynQfQ+Yb1Gb94blsE4vHKtSrmEc
+JFwkAuDcaLuoXj5Lz11nHOTaeQsM490eFmbJ7KZuNZR+fFSmHeTL7eoEQnY0ot8kBarHRfFJM8x
IbKp/5mVi9Q6T95H0YCbgZGTugaWL8PmmGi13dPxQbUuKgIavXQqA96XMfDUFzwGcObPAIoskTPI
8s1ydLwJdSzV2ZWjcF1gcrOxBqfjS/f/6CL2MNkEQ0CwSoKYa0eE1Spb312sOkevEew20yOebzDd
w2gf11xaxRI61ZdvAfPB0ZJDOJqbAgzNj6U6KpxOpTC/w5Delyocr5Lm6HHaGaVvxIA6bP7GHHjj
XB4PambuzUTfSIO8iPJWGJRKfwnO4mZ37pweGhZas/VofnY6UkrCeBx09tf/IoniDrnKxXEgu8gr
loYiEVvM3F80mD4wC9fGyVSLB2TV42X0UTmcRoo8QqXNb/4Z5yWOTctFbeU+6ts3lRK0gkUbkzOq
nNwIeSwQmdOHDAuXhyJSHhUM/QdMq/I+3mWm4JTx6X+KH83UmQxValZsli/0cwNu8Yj4y6H10QVk
jL3DDWWm0cRFDCRRqGE9b7FYrJOvIQ1F/JVEOZwVP49M4mbdxfT3GC3wnZVMQnjeC+6qlTF9N0Ms
7SAB7CfjkCWojuxYFUllfvFLiw6EDrzy742LPlFxNOlA3gqSzXy09bLizSZZucHZocpGy5IBszw6
6o1bJDxot7+uAC/hC0c1bpqB1NCQ8zbog7Sp+hB78byA1nAllGGW9AmjosNhNd+9SBxO16Gz94fU
kMwAByd4BQVBUBGmcbJBh7h+Y37bhLBwrZSnhSioSU7lc5BKKzAZNr9TAfvJX9c6uFk4ZT4gI44C
dWmrFXhLBz8dHSimcGC5YlxMgak8NAAsbSwS0h9kRJj7n/bTobknMdjfgsRxfz6riSlh+XAoANv0
deyiesPj4C11Z3y2g93chVucdzn5ZNYboStsJ9/y7CZTsl2UeM9nU6ZN9owS3wDmpimPS9rBeDWk
WX3IjJqiW8aX90sE9P8pIg0WEHVPgpWoBtniPaVlSWQnCy+HBHpxFNGffiiOf1OhNYSkcwvDQ8Qe
otvxWS12G474dHSF8vKPQPiXEWq9h9F9bBlwgqZeU3rZ2wELmjwzXPAozaYmJ8steOAhnw1unsN/
lQGiE/FG6kh6/8JVQaNiKZrRLwbgc59xrpzhAgpNakyFn7D+IxYLhIraDtvrqMgUA9RC74jpip2R
Mt3ofNrVgmMZTikAfyXz6FD1gJtOylbaddo7WWhbz8L/G07/sZ4lIepu1+mMpgjQls+CcEE38jp/
18JmjZ6jduT/eQMNr70/ohbNbRnB/BAQtXFe0xwUdhHz+wVO44BSsPyybmIidg5panfOmqU1FyqL
RN53vY1hZ4btoPqrn2/0EegscTAmmU4nPBnyyoPmEX5nF9bZeqBBMQ3fIHKP7cxcmUB0bPR3NqP3
JRQ5P/5rJhxPO1sKhEAlxm//Lmagtodrtybr8E2BjBmCQyywucDFe6gebsicz7CVEKGpTVKb0SmM
dQ8SB07X/HQS1pb1MG6GV5an0LZlopra5A6aLHarn2+CbQvCxYGY2TZnlSBzvR95EA+mVZLOEukm
DepodEtWUiha1N2e8cAFs4HM/ikG0/e6uT5s1svBO8ZVn9TKDcNM21/KmM+66CDPRqTv1UkpVRoN
eGX8L4pFzhsEZC0wJ8R3aIOenhdgL6AHNDvvY9F74X3TguGT/BlvEX/gnnxjP983c1XcjR/Tq6MY
zRIwJYvLllxgrk9IAj4Nw3ZgffuDWzOIr75sywepfuAS8Kn96o4JVkggKzpjOt/5DeEQ3qr/xEaS
cRei4aFp5Opf37JmT/7JLpkslUAC4ZN3KJxEgI4f0npcD/yLGK2BxPnzkMfj+km+LsPZSFyhZCpO
YYFFkuaxPXC4uxqG7cGPHmJ8hcUS78EUMOBgNkIOK1YermkGv93apZgy5LMGe32ToXhLLODIWczE
J+qTKZ/V2K2qRrEnjdrIwvfW+xkikMFx3SZqqclYjWK+BK2YYG0haaJ9E0wi4b9/8AoUU2PrPmK7
dWYXI6dby/FRzZjqhaYkzOcuMPjbfzXnQ3mlLODhF8LdVeO3jg/HDGt8crMmZnIqgSiKNwnf43np
Q31b9p2kT0AH1irPi1PdqksTtK8gpVxp9L/HydvNH6TWyVXZwI6V2Yz+Zjh7jvSBQH3dpIKGKyxE
cpR/Qj3VTJLVG5S7q2lirr9UNo+w4rGJP79EUsZz1sz3ALDX0zA20NwPg5sUIPO8YQgvRzIQIY/h
QfeIC8/DqU9Xb9o2A16jKcyXqqMn5ILP6IiNFkE0+sFgHJL2+PZExoc/XiBfpEcE7iFPZpZ53qb9
YWEwdz4O0nS+SMO+kWl8pXXnmnxQNqBc5kbTbIQKpTgHb2EdgTel/PAlSuG0GihjXBN61Y61wlDf
WB/lnDJ674PHmvr/6FqBF7x9ul9ICKt91AD3rmTg/9rQ1EzJFUO1KExifCZzi/vgYTHRaZGXLVm4
YzyLLZD/QkSu8v9zvL2S8Ea5XP6vkTKPMzm9lLNYSAIiLGS+BkiApXRlrN/XnD6pwvKMiYpDEoTP
gkUMhYZAepkysVDvYr8OgxbxiqQSHF2Jw0hxavU8nTVmxTOdAuok8bCYs7wD2zJSs7iuWUKpheBW
Q70SpMHBrLbdS6hKeo9uFtWYuxxvW9/yZeHMoTLjPCRfM3mJcSYobYrb+NxWTSHLmJaqYOarm+RP
JJEO/GwmYsN+IW7YB9zWS9nzgx4EHT6j7YSMRBP4rD5qA2QovfKQ5trg3xS8UjmIsH/YqVcIaVDX
vtGVU1lC6npU+UkOAIAB5srDMqLmQyC5qBIj9mhG7n0AQ60BG7pKC1LhJfXyRLUcsdozqzCvKZrZ
Ned+rvPSRJJjIsJmJg5RvSDxwPvkDfsraPUsdjolW+3rceVwcm4lYMKi1CQyu1p89PfI3kHmP89N
Xa7xuRvUwFvhN8ii5KiImAigwz9I3pISW6+HQaonn7meeWpCyt4QYGhG2or7mbrh+J3Tviw1zoEw
PHLY3bmNc+I/M3Cxdw9KW5tq39z5WQre6xGj3HTIBHsZ/f21I4+kgNVCW5tz+UH/KBpGsnrIDEHO
9Z1TJoZQ6Se09amkMs5kPZz43hPEkzs8gmjUvWtm9cGo5bcaJsqTweMBV/xoobn4RWchEO/+msTL
/EKHeEyRO5OR+qMuC1LMNkx/Ju+wTcuT7fe4XSEbDHyFH2OfgNcWLvxMguGYS8oc0lYjEgPBYYnb
MBFBEStLoZJ19LD6AWltOUljcJO0CkepmxXo6XO4vIYKsoDN/bnRtdYAa1gUxKwEnyevqPexNhxT
kcMAJ8aFbN9lsQfDaNq5IgeuHgczgNM+r++Wp2seFPE7hlOJUdfN+sXTalH4gdQc90eJ15jguKt8
P1Qycm/pHuvV5fdy990ZPQtQ0V2hSACuIcfj0EpGy8912MjnWfmhVwB+qrAZhOqsJy6G5gQ8kIeK
8As6oaXs4lIeg7t1XpscSrEH8LRHrDI5QjhAfEOBwBHAWDKB/ZX8cldBuIpS2anEIiRue2iXybaa
LIC+BAXlei7meniwTSKUAtE7zfvTwccdC56S2bYSIvaxF/sVZJVjW4/SXPkUbeODdRA11bARLNxj
n8a/AMSU9rpZBcT1O4oprSkEX/qbVv/GI2uQsywvQUr6A87g52efvY8kGIAWHHFN9/kwwPH4EY26
brzhzdHL5QYPGZ5fSk9+d9dJKdxuh3c1WRhGNfSBNR8/8bemh2P8hZK69lvVwlsc4ayDfIzwlFWp
0ef1Hz1azY0rslc2DGKCTi7f7OeRfqpgxxbrumkH4j1rNadzMQ/3H/BJ3yhkM+ESyL2asrJOj+50
Nn4WohS1RhpcmIT3C5oSKOArNycip+gsOpjnNKvuUm2fTGuht4Xrd9R8/l11DzeMP0Zxzov6QeNE
pM9bDKtNfCYRB3afE7RHrWrKZJKz0e9JxlPnZMNzhAskEn0mRh6ltoMxpbi4dMgEDKmu5UiI+Hw6
bG0DKXtsqquA+5kb039JNF64Ie31Z+2Ne65jOEW3hT11xTZnlFZkURTrQQCq9b+QXQ6ANNSK/K87
dL51NRTFS77/Q/6v2sQFBhhCLOXpgZDnP93A2HHGMLBIo1RDLttS+4typ1uCufBt9nx+p3JJBZTk
sqIgfqySafc24kOlT+H/B+3VjYNwzQ6L0K9NNY/edcfi8PBOyX13xx3kaI+/qYj9wEmEB9I9x1jn
FygoSden+OQam6aKEGsv9wJVvWGo18vSsWbYUoi8/k/qRRU8hv+XF7QmEkqBxmbxDapABrcrZVcg
FUCorgy+wbfJMCnQDWLwObZxiM8m/Kj3aTuMIX/unZlxjetKV3k1Ccnue+dOZ1cIg0GoysN4A8fH
YuETS02KoyX1SVUvoGaeJOn1buwzZS5SWwItmtbfXxQgsD5nf73wZboxZqONJ7a3XlHeMLLsaCAR
keKBbeGLOA/J5TyXHl4ktqxyQPQh3FSvExkJ6croa8aVd3RTbfMomqjy/IhmapA3aLqgJfylqL9H
UaySsONhWphEusPK/up2kWSqHfVQsAVgadvYqWwdX3aZd7rBtIdtYizjgFrE2fY4a9mtialA8DE1
r8MQIXHbXiS41BWiiyPZRdobRhqFKl3xtmue5Bo7H/11IzUxYkmOVLvxojx9+xJT7mXhzxkDcoHw
zytDko55Vqy5PGsTQmAuRy10jw1EAl4Fm6nwe5/7r//bsxBKxCgb08IYDDAE+ASk5vRzSRW12mY4
Y3H2sNVMcn5dC5mjlB+oCAJd8v8iKqzjxfjMxklUDDlvOfzOiJTOXjYSbSZB57KX5g52Da3eilFi
ICBnyBLq3JdUlKpdauM1SxDGufWQ/jghxaqVIBxze4wwoJBxQv3VecNVDV3PGIsfmK1nkBJNvoAO
vQK/jJQ57tKIpw/WPCsYQ25bPVe4g9kKzvMqBsiHdgbrD7dizHIteZTvzlwj1Bxm5PGgxcopjelJ
qHIagDWM9P+QXGh7CXY/E5zS+vaS8PQYanzgtj7e6mtPet0io8wkQHLcGn7/sgijQ2RRLc0EWBqn
kjEhTmo3Kc5FZ9ASR2XNVhAyTOq8cwFzaAaAPeLNi8+YMQOvG7YS7ABcHjzD8M+4iemxZWBhiTbc
mYDHnto+6wa497bJL78Z2lFCNmN9g2V7Xz4TsOYE6IRJ94h5AY0tllT82xEg/wYn+AJb9adWNVZt
N+gh/K9zaH0XYcOJs2D3OhUj3Q9cbAzkTs568NBcmDJJcl+icYAVHo1kEb2lZhTmegAu3J0RfP+x
6rVPpIEDincUL9aLFnu+SfHwwDykkSMQOUYNlmiVR0OTF4JEeXJN7p2lYGd7on/s+arF3W5HffOq
fI3JuybMrlIw3O0QP2k6QyzV8aCmLr+fosXlkuoFxgaWeyC69UY8ch6od5Jn2muFGcC69X1khIhO
Gbc2cvXLe28RgcBQACyWnec5ViIWRIabnAPYcXyAiqx9MfDpv3NasNnyrS1jvoc2m4Ehzq58Kq8J
g6frDkM5GzJCN3yxyBcadUhYD1E3+BG5i295A6TXq25H2KLSdNDY6aXtIZAeITw8RzUfGgvAY7MO
sDJQWjcow81D7d10fOr/ETXK+6ZSj3HhuD5tgy2NaHRqSsZDgRgsrZ5zC5TsYyOEXYb7DcAOHZ9r
nP1FA5jE6WZHM39SZPlH5IWl8LKvfYbEosXdrNTXXGeBOlGc6AYDdH67uo2h0ToqDBH4ybusl+eb
+XFswtZZd8FDVK0PVMxfCyIgj77YA2dei/qWPVezlqW1bMELVRGlnt50oTSGeF7AV2gMlm9hamJt
wIpY0q5hU+nKR4OyCCSD4nf4FNrCKsnCVoKyBLNJ6BtvKn+GQGpsGqDujqFam0HaiWPIIDYdWbiF
dBgQSi7OMjWkDyUklXO3137Iau0BQeW1+6F3pHYC1+v1MXwss9NG2ZtkRGzC2EexwtWL4ul6l4Vx
cEMaC5c/yEgHCFR6FpheaQRws4EfoLnoV89uaV8+alZzDBmFCqlcI8sfrudjt67z8VEVkGin1YIR
oxJw2kZDwfqr2WRD+o5iUEk9K5eUTY4PZCsUZgl56PswqJQRFCrqYQqlKQ5ymkR3ftCfd+VL9Jxk
G+9CavQ1LKVRLxPqH3TelHG31olF9hWA+qzle3M6D+kEUxFo9q9w8aep+iL6dItmdnm2bZYQA56N
i9WFbgZcvHLEAhp0lZn/KFsM0/h559HAG6GudX9xRrI7QYRq4ibVNXJNDxYZImnn/uQUKOaLsXlB
Nrlb/WeYreGPGx2FH65R5IF45vLnKxeRYFsrIYAugiDGtLrap40SDtEZhRjJAXCAbr747qEvB0Yj
0ACJ+K4gf3Z6UU+/CBKjg6FAlhEEF6Nx32SGjJA8pUSwD/7AUnyQlIrD0EX+N/gtNl/CLxzcOAUH
AdkzwJPM00DpqnAOlm9+0lgr+qEvzelTbAJQu6KvCWtxjxO6EbLWOb2AYeCb2y+JxuSp9NS/G4oK
YxxGkd6GLh3kwADl8+w+lD/Rqt3Nujn5cPrYDOuCe+Y6RNvuMZeT8yd7pmpLu1fRgAwkHKdxQ0ut
dY+iuixvGAXQkdXM3feDCwd7zTiztXBrue9jHm04Rv9iB1SDR002llVV2X11tZpjdhoC0Zq/+17O
+MkG1f/P/Uxov62yhLl+HrYeqnBiyvyYRXZSVkpRzWg/IFGp6u8GgDGl1G8rC7f859BAolWvHlvI
hqhzcUBBxNVru9Pysb361OGDCoAnnm/jiRZiZTRGZpoL6S78/K5PQeqN3HTyl/y27Mx2TY646LN5
VeMdtS5bEveCcnxsJR30pZsarfpdllX3CgqglgELpgIvKYq9KlyRU851geF6R+ajBxS74luB7u/Z
x27AyrzFRKA4ylUo+sx3GwV5DkbdqvqaZIYvRNQsMdBLuLjFKy+2ZAkdEqNCMQ0UHZkIl2s5Wbns
VjrYwniFrui5lAuZxa0DeDiUd3ytxon32ReZjEVymoM5qzDFqlUCqm5D6K3YJRxGIa6eO+zTCs6h
HKq3rdDf6V8ohIwI3mlQqgUiDs8Yg7178PxIUZOlPwSf7YVu7H2tBhdQT8MW9Y0Cg7BCxeknqgZo
PhXtYE2F0ul94cYWmYsTPSX9HHzY2riiMtEYqoUMVlIkB1fLPfUeF4+wQqIdTWGvpp081elVlDYq
YCbEt4IGJq9Hw/Hmnd73X5fdlQMrKQL9DT053xILCycUZJ1aDjsjFJdhddyuQYEcQMz3AuQhoauE
9MK789eaD3hv5tpI5V/JxrCsu+3nOSSEPjUmCVSxOFDjMAKzbIDCUB81Pb2mDZjHXYagXEfTDG9C
w43IA0LNN9dwD8OpwBjpXQoXuKRHw0NM75t8nI6lpvW5rHG+FLREXjmbkDTfKNS6W6unPhYmTUQX
6pwvrHvS04P/3nbY2JczJgXaYjPEl9MJIHuzgkSmxAV2ycB8Js8AwXW55zPTCeVV8fYR4el7vn1I
Aqbf0krydxSR654hS0ATGt7TklQuqiBBQNVdfxYGG52gsMICFf64SIgAUGSS2NKZKaf9vWfns+xl
3E2vHafEuLqbxPWZcg3F8TLxvz0nKyVm+A9dCUewGjuwLoU+UYPxZ1Wn3ULQEZWfFLWm3OFPAVmq
KcMItqFfQeNETH4Cx5KemmR2gsm3PEyNqpQoNQLeuaOoo1T/+4xKL0GwGvGxUyotCnOP8VyyLKz4
uSJNsVKctR6rcLwuVRDLKeM4hcrh67hjXe48GRs/vgeOdXBNwMhUrhzQWqei49zhU/fd87C3D87y
FC8a4xu3d+ZaDfwRSC9D1v772oFEzYTN7roHoZz5u1NZV6cZCOHrkKMSI9MN76EhJJs3hcKoZj15
XiF3C+ZlXuhFuCmOHAsy9Hq7pgRSojJQnhpJBK70PBtrln5yUMDxCmVizuQmsdNIPiTREqSRgvlX
budyc2OB/UIc1gOXUbzhskyncgqBo/wlbhK+iFWHX2xchM6tGAz6GXGq3f20mIjmA4pjaGuo7spF
TbcvRwv1iUMa9K6Zpd8yHEdzhP9Eh65SipKmc/s+GJpsr17PxD+vMpSmSQ7UqQ/i7rYqBgiNAkIF
GFtAl5BOGk0Ft/bEgmy3BjQCdi0GwbWtr0CnAcZRYtelhgK7nVi0h5XCM9U7uUxbONjSwgsHoUmh
QBwNW/LxFhCABesF03MZ9WQbhI6uXFW9eQGRLMVIW5ymOGfqnDgxAKeNzcG6X6mxdDy3Ur6VouBn
BzDpefVpMf40wBJgcyKaMbOTuN/3i70NrVI6yUZ3cwrSQAR5rt0ILNQcMmEdXS0pSAKH0cqy0DXz
snYZ2kJA+Csg8csUB0eRaRHRfRr/XqjuGDZFIlEH9W0ZWxiG4Y9ImB12wWkfG5kgD4jOJua02E3+
jsXLvIdsetHc2hauKuvcRh0RzYGrRpPP1/peqfIrMl3mzcRCdmpYpKjPU2DrbHmHnvUo6KaogXAw
N38HDYVbEjC2U4HLQ0+9wpcXPRXuJk+q0whiqke3nwtDcJ7WdRMp7qsuYzTh4AGmUEiHGMszknZF
BknQBKxJ6kfEhANt3kfkUMl9qDTKu4bFwe11f3cckx25eCZLCQQx1GAP4H7K64MGj0kO2UVBGzkR
pLfO2ncwl0XaCxsHjcqGWv0lZaD0n4RBE6hweQ6oqdmUEk045dy0vOMiZeIa7ORRRLl/1lytmXIk
AQEzoeMRvYp59sAB1u1VvUeQ2DT88Tkk1b5zRf0FQmjpI58j5qMkvrWN7gon0v27P9B3+GgSPPsT
BkDI7RL9G0g5E6q4vBe5PWjJOJw711WQxUAnJT/7T+/H2xx6vrydh7W0kA7QD9j/qtGFDtWCBZ3C
XaWcNFArNWXdklwfthun7YerxQ0MQocbB4mLBDWS6YqFyuyfJLWqOJjMBsHZl8QlS/pY4UxHI50E
PHcbbZmv6OEp6+awlAr0My7WW8GwcfC6zeHn097275jtUfa57tKuZdJx2DLkzyym23dvqlWPaGsl
rxC6tvxXiGu5i8GbBGbVBYEt1XvX5I0O5C16FTiEEElIpKQIeZtTgkjac4pTn1B4Fs6uEXTLxB8i
7G2+Qd1kw/BoyDXtxiJSkhLZGaHSsMS6SWjUvenc8AAYa/R/UzDLtkAtiaDb/LdYV6myHS8l9kQN
ROwaOVr/VvMskU/r6Hy3sRTFqMD6HiW7xw3/sWp1RQo0Iz8H9a9sjFAuROyfkz7cVSoykDn1ByCF
eUQl6xYDgKLDiaIbqCyISAvFOcbnwJ1y6jSKcTf8e5YFEZUj/c7nF/hijw06cbRXeko7qWNCBcrg
qoaz80KPtaRRfdmJfw+HkdZH5/YrZVqdmpjk8XnDjhinAgvkUVdGnLu1V2fAuKeijyBb1Fsk99Uu
EUhJi83j+NGpuQZ1VIVzyVVLCWBfRgYqGlz68g9vlAfuCopmmaaud6+Yq2uBji6t4q/V4gIEvBfP
r52TkknFu1xYonhuD92FZQL1g8nLN56SkUN9yrtH0VuDcmWAMeFbJ8Wp/zky6i5M9N6btwhjuifk
DZS3BoPLU4yMm0HxATWBy13gwigEC9TukV/7qIVWNL54bHms7cExXh7uh1Wwa/mIlXlcO7/6HNKK
S6JM4Ahj7gxmfWa1H4v0q70ACJG1xyrDPMnvaxTRdYO2b1JPQLe8IjEgqFFpB5el6WNTAe0hWwR/
sdaDgTa+3WYGWxjRcXesBSpnp24Mk+61IuE0T/iGldCk93O2MWjsu0q5dREs7RX5GJ2vBSXhBWf8
INPVNh4h9Vz5FMcPtzitiFPaIyP1aTI1SZBx/fqAFhOiiRiy5q/QpDCCfbjTLEizvikfihbg3kap
5uvPfpcVQMmkF0jeiGszwAcsYsX0mzgYRLGaUblBi1yiLQJFSxgldR8zMQE0hBmgSIpqLJiTtKG5
2dosYIxWe748uOE5PWaKEfPslSIgF+dSis0+O8YWCt0b4bIF3NtnblZ4RQW1cSz4SARFwA9EWiDC
WUcIx8FzK5qPO8dLJy06z7/ahNJbcUmZ9k+/7NlxAotqxRdCtHgroj+/ZVZ//vOj26zNfs0r9Aql
HtDmfyfjqicPWnFzIgzDFWLa4R3ahjTBUVGQ0OVw/LWUjZN8KMP7G37lPVPUhbCsQE3DAMTbZlF7
Tru0x4qmHpwOfXDTNV9Fb0oYdNpUikWqZJWtGJCPjQJ1bH2fgwKcbCheaaneQYwGLN9shT+r8DRR
1YT5fgQ1g+lPGVnhGigo6swgahVn9zGT1tS65YfblQ5f95SxWgzLgS/Lc3IXa8xFTBcri9Y/6JiE
5r1hJ8lcuLHF32k5Mn6W0zFyUehRCy8xJQz/iB4xMMk540QtDYy/NbSp+UHSMcs6+s53eA3IPXLG
OcAWCp7I6kgxodRmim03ydGeGvnrH773NNulg1YmUFE/6c6zFzBl02VsIaL3B8/qxXBB6SO6ofdA
kNtZYOSRowg/QnKRAbitlJgPuoj4yPIGUtFwJVWa2EqIicAh1lEzIy6mBdJ/digiWAznncp0jDXT
MBr4nDsfVA0TCYHo8vrn7lmBRy1KxoR8GIH9e+M5oSzZ1/5geZtLR9KcmIPx/RBIHgQNBWAr5rMJ
C8zhMSt7wv7+LJWqsdMqC0KULyLFFR5+1n+qmtZd+5Ouox/XaCE7RSOHIGi2AGMsEFQF+TnWM3L7
ynkCFe5raxTJMY0sHEp5VgC9CVbTyNIPQBw483QlZcojxLoNWE+5qu8FvWpRAx0N0myiRaPKWltc
lYXNuN9T4sGxNwCmPsYMX1SYxdI2kcFfmznqzbIg3orvJJPrNg/LkVl1rZvgImE0dKk7vDMeazGg
JFFflQtvrhlUnttiJuU2OEpvVMtNY7La8YucX7ObYFP0RDNaeeNC6/wpNMEovdW0dOattyiPYbcx
LIHYjF+aEUae4fSwBgf/EM20L8H2PYEkNq46Afm+B2yPoXbOnzcUnwG8fgkr74nGV7WljhbZOTSQ
YSU0wMExxsp/6VHIvITlGUfW0BTdwu6JfELP4jKhJFs7XIezlZNhQ3MLUBETDng6QjHzSS6C5El6
LKIHOBB2ydOWHqz2UWM/WzriXlJxGD9U0eldkEgR+37eD+x3WDR3DnfMqCVExAIhhVkqW9tcrmTG
2V9fVB9OfS6AUBKTVDpoNCKog7BDeVQ1qEMSGViiMI9Vfeo2NbJ8GQL4+4t3X72y/XLoUyA7obGF
gjGx3feYbDebfdvBv5e4A3sSClc9DxIVC3X/LAMfFMYMzrMVjMUiqfiCbCAHciSZ04UN9O1xxcjg
coGHtXQWNIRC2OLoVvVm+f6Ug8Wml+x16zFwaXXLOYmfYL2ATsUobp+SbZQFgJrwwyJuByt05EEX
WPAY+XZU98b+tZWSEz/SHEv93r1CMUr2x4eOTQpuKSDIZNrjwbb6KVaC8j78yngfTLiLgTD2sjgN
Rvmq4GF+qnefAydnWBsAryOhmMqeLqjNKE8h0ZU1yMsCK9X8rXqbtyERnQST+8gvOHXrXnaH8OJn
RxHb6EabOX5DGj696+zEBk1rwgzplPc+USI/qLyu+3Y3Mlph8fJu3TmRSES/2FMjbStXD+OabMm8
KMziU1WgZxi6DXQs35HplZ318x52s/I8/Zw11b0eoipo4dZoLPUjh97Ic90gDGSGU+xaPqbXWTif
a+Vjdtv+YnWx2Jr26tfqut5QRd+Q2Jscs34bQizznYRRrBKbY/IqxwYoPmUEDwDJRFYCMO/1gc82
fBAh7Ept2fC0jysT7Fzqh9poz7bwH7spn5NYQ2Y3rkvUXmuBQS9jnoTymoDgWAnazQPW/TYtzbBB
9/B5CReSTVItgta6Scc15q2xcMmkoOir6x9thI5NLgr3AONrqmLqGsHL5f5mi9t/7/gCaMfos35/
SgArPOz7gPJXn2kqDfIBzDEHgVgYsqEqW0NZNifQc/ne6iZeH1u6+I+VlGGXeZ8thxD/+AQnGbyD
X8np1Jm+CqX+3JlIfUMlLr77LnmeI/rQC1Zas63PoERFoDiXXBDjnM4A+Lppj0AMmKm4qmZy7yMr
hFQ1Bwcx7tfN4S4CoDXb0U2cK4mGXO772kKT3WKhip4Z1cy6aS6y74NjHL7R5o1bRDFCAFOH1PJU
qZuAulk7I0NYoB3QYpdPVtKnV6LudS9reQz0zx/uZq8g4DWGPNfOZyUFN7ENUjbVIhN4hJZdbylL
ey6NyP612j5hNWZa1vvrtsbdfSLDxkw98/LPtuMUdQR5O5tgYOme2Q2doadqLXQU84g7UeAXfGab
rkfqBetFvADhRVB3TxNPMKiVGw5AQERBadQ0eUBKDvMcNe9XNKcYfr/gSK/UoOos5isbXL2upqCh
/U5gp/hbI2h3SOgUXIxwTXv3ZKVreLpDh+a2aM8BUOrMhZSGvr8QpAh9FnvGG3QMS4be+ccTsjA3
FrhyN2fkEL1b/nBLd8z3EVe8rQY78U1zbJD8/SOhrxMt8QmrsfJsMOWPPSe1S4GYjeTVnefcANdc
ohHJHBDU57j4F//vtaJn9WlIuIdZdzcCyQlvB3R7JotGgP99NBzA/MmmfrbVRPnApyzpmV7kkqTG
QiBukOxKRgG4Wk2DeR+SfvM0eSURdTpk6QmaJ0a8EckBJaFdeO/6s7chENyK9ncJ6FcA/jooE1GN
6xry7Q5HC/mSOnwWJqXUgTsyuHm+8EaIHAQKglFa9kzwvOhq3piziUa9MVb4tdAAFB5nvLB/OemD
lqdKnSh79VUGhPRYAnNcplvA+lDQT+s2q6y5Mp4rqUiz8J6nlA9bPuWMJypp42NuVjCdM+56CdRO
qi/O0O0DfYVWVZdJe8Ba8y3PJQK0rA3oChvnxk8EVU7lEY2Oaj3sWq5AdfHiMKCEv09zeUZuC6Gw
otd8l67OSUifE5u9cPHeAV2803dgNBuo47Gok6iZEE9J/bgWBxAHRpSGEn1rHHmbHEqWo/QX0F7T
0DERm1i26odxDxr/xUN4UdunNWVxeD4jzrJhPW3vjGXMyDph8mg6F+TIuP++f+7p6kmCqHP6NBzG
0wtBohgozLtiz1FEpqTynNxLlxeOHS/4DKavEYIZkozupLjGtW9fnjyK1UaXqn4j0jNjJrU3K6mE
ZE2o4kB7AQqtzmxXj1S7rdiZkhOsiakF+Z46y/EOtYGnRNz/g0x6mg61tRvSKQD6eEiCsuHtuees
cKGB8vw/2qRFZJihZ/SsXBP6T4s03Sz3Sfq4AQlkgT2Vpgx8SLV/gcpaioTS0MvT6WRKkeQwdLBf
Z2UJziEfyVq6S594Z2cZPXXiSCIp9ysvExqevKLPX1cus7V50bAdwP8u0qfKocvK8MpMe9bvPE89
Mnyc+uE/KmMbla6jIXQUOSkUB/kbCmX1Ye37KcpOs2ZRtp9u2s8eYfClU8eEVqvnrgoG3BgKEIzP
XiCThWx+lIxmzQwYFFCDc6ShOLOHD8m8Mm/BlhLi0yKGee3wmQPiyBzhzUuGZwrUzQWuV6Ir5D/2
UjNTv0ZQJT8BsNHo1WiIkUMWMmAM6P9xgxVMNFb/7vu6JatPQxc6F8KyRgyxoQinF6PjgDoHaDE7
ejlcYtojlc4yZsJK0oqWAHQWce5fkZyuN9HF9LhBDuJDfpxeJad+KkrW4um1rRv8f5FoOXdsb87S
E+eTMarTwAYo8S8GgVhOTh08NLCwCIqE6y7OKTblmdloDtfYm9KOq1T9SR56Wz2wj+sX8TFO3VeP
YaohiP6sCZ8tceXGUBAJFx0nmFAc+U/SzZaGpj2fCOy0l5eNxR4wqYouyiPJ5r8tvw88g5bF2axx
BLH50XW4EN+q8On/tAeQw/IoE7Mo1pyrkN/6pcsrWrTxAcOZL2JIbVzbhR+3yZKddZ/f+OazQWbV
W9xYBT4sOcRXv2QPxpF0SXyEi4K5W7dTUc2hoynbTh+3LAEqFeQy8pWOj3cE9Tg9FHUqYO6RzxPc
ZLN60C94+1t/+K8mPtV2NAUhzlzgVRxXLPawxVjim+wgbmp7eAU99evrO6GZo4f+PjZVfKFwH1Pz
8Nfq9aWAc53zhIwvdjDzTrKOrlvCVn7TQBae5VK0WHYjZbt1za6JSmvrDMyezklaMEJKDvaQ72iZ
WyMF1w5GQ5JNaXcux69Bo+5SyYZwIfRWUPe0qR3Hd9aGzxudj11j5IyT1okfTwRu3qgUHarLxViL
S5eIpytbQTKVajYq7OapfBR8JHsi6FMgHq+pEAfohbK30KGAkW2+lTyrDw9InWkGmaDvrvFoie+d
FFYZbw11cXT2yNHj3HVTrr0spDMpOM+JLX5I2hBMLqC5gdzR2UmKLiNO83DWiCOu6luIAbekrOIz
L7DMamNN9aZ7qmXjprYlLRCUpOhPpr2KKq2rBe6jdwMS+0J9ec0ulH1WfeK8WrZ0x9p7adR8WYRa
CY/4UZ8C45vC/K0aTsl+OM0IPeL6g3vmXtt6lFVFIRs78VjKBoFoNMgW9bJSHN7H/dQ9iz8JecQm
lFHgfLmnzSvkfqtCseis8dp/sMhdDlBTOovIdhoyILzPJI+2u8byTBJnXrAvQQhyPM06R39tHqMW
DNcHxJUHOz6iqaJBomr0aNblg3VavwSor5gAOLaR31OfAIZPikUQBlkQVNzce0nO+T+Uu244cGIR
O7YnSqmAtqWT64D9kGhWAwFVyLx6/BdV0DGGeX/KbeGJZ04x6w/yUfoZhTCj//crsiNzE+3aeWCy
gEcO2FRoaNVa/xujYl46r8gpM4mVceAxwJbvjXsi+utdeDgL1KDtpyEgyvIgp9aLZYgNc87VG+Ue
o6BJS26xWT+qDnrVPklrrTXqODtgYldj/9wcy/hPMWmaMwrw/ZoNm5R3OORDtsqLZUu7DaMLc4Zt
Ld6vi4KpnYmzbYNJlBgPa2ZVBr18YMiChWsLlxiMRRVOpBov0eKgNK0eIqxMOJzBv3hfxkRseAdf
72bbGV3vTA+mc4aXiEIqjJ0BQy1HNrygrLhuy0pkBv7Ar+5S7UN3246JWHpTwl/uNKOjQ5UWKZZb
IkKk2zKSbtF/PhLueGzkJDZDFiBeVB2ux/389dKTupwkvJujdR5ubw2vQEQBegEofpXm8cv7yix+
LTnmEAruhukUVzG6uMi+XateorRaL07mfCrCitIJkmLf24tqVQq6LC9KpJ62nEfRL0NcXFsyzPVV
DgsIPRuWhcLM7M6X2L0T6TFFiNsugaBpdqCix+dsXZVR2CruAtCOuo3ZiSiPAUxF0Pfw4rgc1VK7
gVG9qrvBMwNwRtIFSLoo+uIJjEQ0uieOWoCv4IwDUxbf8Kr3GW0jt3uC8GYsVHX1C1Eqr0LBlhV3
pfvuNz2bEOlw3ITiuE0TWFafcBcGd2ooCwmY+uoDXJ2BGXQVILnjL8kWvHIXJiaXleSlaLB6BZtB
JkNA78n23JCOkimSiC5Oamcm9GnUpfEZ00LoZ6UEkdVPiG3cPxSf8kAGZO8ixVtLKnAaqIK+y8kr
cd7VG7lDwjiqSCQhGNpr6tNeLCVjmum0qogTSMryjhSxmrdCflkopXPp9lkksjgjZuGuSYgomToi
gZGE07D20WxtAz7dLQ554ftXmHX5dhn1hVwPLHw2S8SKGMVUBq4/Gm6Vpn0XrNU3oA5/ymUnMbCq
PEmJ2/ffbOLNErZ66b1ABUCqNW46n8Nuzr9PH0uzZp1FHbjeFrb8BNR8J2EUI0KaUKz3d2vz59jj
KTV7fOZPJw0rm2fTN60LtXB354lQGPxBRREob5zTEl8A5/Wv1mlWK2TAqPOqF1A8D4TbisC/f6iq
NJYYtGGPhS183ZybNDDueekUC41G8/evRgYk+qW8hZ7MCNF5d+EEbOvFOjWSAuFUxyYqsiU9aL8E
XCAWrOwqch0mUdDcSSxv09zVnOUheflOLLWUYj5zR+JsR75kZJBd7jqoIgSmu7K+SHG206GmR1iG
gcpJgDbMt2+BLs/DxT9IXzctL786RqMKVZkNKKFCkx79pCwyyhaPT+ZewlNyJ3p9TJo+HKU4tUTC
k9b5IzOzhNyiwrd1wank7tobs1LYomBGBTOyFD0B76Noifg75p/1bDgQwEAly/Ad/4abtmk6nbAM
DFsjsfkB1dIqhDx5YX2n/ELmIi/nX8cLSVp0xj1Vcf+brqHOX/dQKTEYzjB986VwvMHgDMGijBvm
fa8jBU/IOMNKoGtsjF82cuAMaEygQkPg7TtgHIv+TFzncywQ0cC0jMt+GDYiZE6UDNbA6IXyD97Q
gnPgNYJXnvxQ8KJDAly4Pihz4nhQy2JmreesJzCY8yJhOvT1vVF+36W/tZWeuSDi77t6dGrhD469
G0kawsYtm96zZ3UafkYhRly0O7d3geBQhN1g4fH1DlxlixyTdOI1awSZodTtemrQYIrihQSVFi/e
8XHOwGKHwD0ud+jlNcGvJATMAUQFjsb8HY3mAs9YBAGxm9DPrbUqcucf+nokZaagFjNb7MvQ6Eep
rMX30ntw9uBriXsKCM0akpdhKmWxfMBZajIUWVoqE9HsnG7RNAFh0oz25jsR2xxci1hxjtovyhT8
lsy4IHcekunXP8oQWAtbavvsx+x1LptvWjoshqXjtqL1UlMYVsAQJoifsJJOizBbL8agXO2506Zc
3673i4wycMq1gaeWpsFmtW218wDdvx+2Rxzxbc/JP2e68mow2/puGw3Jf8chwhk0UBFXkdmUzFJa
WI0KoHQ3kNAFn4DZRxrBzGfFq6qGOlVV6pxExNXZNQYNQC7Pcwie8qQJGEEUiHO7DqGLMOiNDypx
njzdVIZ8l5gpwt4ddeNjH0Tz4sQ3Qv+YJgfrooy0KlRQq1EhmT4YFtj71+Q+e+F40LCRy8y8CUrj
ELh/Vwd1jyo5JRR7nrH0Fvlc1fInWddAAOYdxyknId/UpHQ1Zd1fCNlyAry/5TRMlLlxXtr/SJ9u
g1dKyr6osIkYyaHzeYack9giSUjYR+2MfDeEYmnB2foa84lMe00ixlPAqghxGANckSgRL+xHEDZa
Hp+8vkRTLkc+KGUzQho0KuRHbm/QR/SC5X+l5YwZsA2mrKZflv78TG3reGhHJjbSRSheAUmKSzx4
XDsEp6i0hlM6Cj9dD4jyFSp69v/d5Mu3dth3utjlYo5k5hs1pi8KcB1q3hFHq9Wbi/rNuWMuhDc2
GBtEs2PpWQsHW3rhjgAQMGQlGSFoMn3URFwdXwzE06REmSkQXLRUIECnLSBoOdgL2tW2tPg5/5g5
ORD0bKA4bgvTAp9GkKXd8BqDBmdWy9PK+xiFNWzXe9b6ZK4ljJP1hJI+DQ9S8KiyCi+NS7UtdwhT
I1edntShLfafJDSDyaCNYP3LvsPZlbORbkcR3xIFJ6qSY6pcjBR2q0Yokk6fTebKxH7hh/VdaFRf
GFnpk6F7OUtnJGHQ+i9KRxw3TjGIxL8JCLK6VkUaoC+pjHPDum2ZhJftJjWQJhk6vhpM8MdlId0c
QGs5ve6I2+EwnL94o86u7g3jzT5LF/dARmfLcmGr4vl3e241Vr5t87fBwPo9FM1giESHIGXtt/AU
Rq/5xWSoRTw/LCkjf5mn0sEesC1cmjhGCBQky2bCP6nAEn7OcA042zxJc5ufqvyzSOKg0PzXab+d
CDPeXu+uO4pOtjJarJSNKXjoZ5wWXURcaHrjHx5NGdbVcKUXCzL+NVz+d/7DcnkswAAuw4oqvXDB
o9GFL/+yevksQHv+Cue781PGiM9LA0c19lJGuVFz0GRLDQfmnmMrlXqdx8nL10mCjkfFTfLj4X8r
u6v9gXSn/pLYzOn2rEhg2IVKO9Qal3oAklMJO1+Awoqhv1PiMRWUkhvVMqFtrDbutUlcCaHiMqkz
ToL6rf7ksTZKHg183zlSNvDAftMfAHwUHC/2I7enAD/M9Q1psBf7YrL2lfilym7J5SfFWi//IJfv
1+7zaHX9KZVBpyYa+h/C4WKY0MIE7m9YJjwTgr/vPkNd+qoTB2W0tLuitl8Pva6v37MvSsYzfJ7a
8PKVUgh7cm57RS6Eii7Y9KHJYUReaWN+rqhkXEJUDbcC3SRWWdKTXW+7fxgYVZHiabQ8zlbGC352
D9Mk0kCI8FEblzi5mbudKuWfTjehHP5lj7NZlKlQJw2OSm20GDsRJxrZpaBtMewUY5NvLKlIIinQ
WuN8iM4l9jAlEj3bChpGXdqTtUHw4/qkqJFMg0rdbWBe1AiyCAFOXogMxe/igWyTMsoElO9c0+iA
T7NmCqXSS6XAScVVP4CC3jULDNDtepBr1lT9VvoZIA2ruHJUHl0Vy2tNZ/sOh75zWQPu8gsbkBDc
+Bgky2JU2Hh4JEhVyExceoDB/koPZ2hu0Gwl7vZuQ8xnbfdvvm1EvmNJJ61D+f41jhwa6/x6KG1w
DNMXdo+bB1V0HyDD9Roq6J5jjLLVAbL39A46cOYzBQ4iisB2yiu1/3eyXC22OgHSvyIG7tp2x0Pv
6TKLpm202wd0PiMh8z/ARl5yQ+dIaVDRUh8JbzMpNyonILnMKdDhnIGfmXB0e4RmWcOoyCmtJb4B
OZ4DbnE4RQjLBg1uiEdXVqx8bSa+/m984AYhM+DI3lzWDz0/h4tT7dVn0xuUXUM0FF3p4DzspXdL
7xbrjZI/cedV56gQhY3gdhCuVYmdutb7mYtASXREXFYWrAADkVYOhEaVrAPPA9Ip+zLBfRWnwfxW
KFv+xtvoLpxdLCRmlUZOsoL4DLPtp7si/nqo5TLEWTgvZwmF1cJvO53KrbDoVFS37fJTpNtJHrh1
9ZDVoQfuUcrhykZBmhEoR/yLGB5iKrOAY4Vq86kQHNNUjKvjbX1/okOkNQZxfzRSKcBFt+mnGX0B
yJ7i0BfqfLXwxvyFwH6aohJNAqdEV63d90XTeDaZ/it1sb4KjYpwEpolMjBE7kd0WAsWswYTVdOL
PwWZCWBWw6ymcKmmllMn7jF0mBdpx7F80tDX6KwX3CAAcDvvbtdvA8xhy3Kt6RNNStrW+Qz1wpJI
lYZEoN1pE6x9WtdeT7pPy9vqKEJ+Sms5XLyzGkq2CEsmHG9alC8ZdYg2mhP+SeEPs5lgImAMwOqN
SmxJqbzqYu6N3uVXMH3ezIQ5a5z7auiMR2gy3Pse2n0FGQLZYekVRWg6v5vtULyo7yu4klo32wQ1
aB/j43Wv7XrOMgVbLdcW2JDhqb54V2Hifd8++gjApjwJt7svY9ohcWwCwnL0XMXyr6iSu6MGu1NS
POASsjTGTtYdxloLRwwzWKH6RE3wo5gO6f1ZW1TjggmfsJJoQg+Qze4oPfLvss1SrqkX7ga2LUzX
KCzR1vYNLmakD6iJFfy2wN2o0XzNgS7ZoRuRE0qGMQno0fca8mAfUdQRkrC6bYLf5n51sCelAQM0
FbpalGdxW8O7skSTOVrp/6u942qkrb6dLjUlwitkS15fqr1iaj47785wJwkPyDwvmAvqi0GdIbvm
cePQIMnRaV3jnCt6FxPvOyeUVvn1WNdRUscnqEGk0nHFZ3Cmapcv7J0SWWBNlMrkV/IMGNkZzIfJ
gcbE0Yv7Q/SfyQ8gNgQe2Rd2Zqgl5qgvl4bi+9MXGtxPmvC7QKKANyHZO3Xt//WnJkcVBs4aB/ty
YNmcjRZIHV/xAVIa0HIfumBNvblHBRoBD/XgCyOp6QI7sHJ+Bb6RRZ5RVF2KLp4mQohyQcZ5zeZ5
xBhpI0pVQ0HTa7O70VYc5zbQZblWiCzKfA+OzRb1J6FoQD19ux89asGB/ABvuOoK80QuDcOcnsjf
6Qvfd7i6kJi27CtPEyHSsefscLeSZRTsrCTcx2iN93whDVFL48PWgvWGrtX6dxH0fJKJIFtdrRuH
8KiOa9tSav38u+yWy0YnmzVKBF3y0xkImUUGz6HwLSDBr0HYPj7u6P7cQMTUhVZInYwl/9laE9ez
WI9FarJjiU353slWE1KG9m1w+iMvmwJFxCVLl+SQ6dY2xmIRTwf6tMOze8vId2U5iD7kJpFvss+2
5sw/16MbqQkEcR5aKR1AQ9EB9YYHFgPy7ANfphRhFJEEBzGcsfcP9ke/GaLKZ5dezQIgEj7qqzdT
+rBHnagzXFOm7CJQD6k/L9rHysemkgSC7/gWnkHy+naawY8i9XzywwEDxABXNmUbtCaahKFodlYs
w8J6dgdZsSvtzS+H/MrO/7fo7t1LQeIAliixeReIYV0rY+wFu5rvYbHwCYFPj5MZG7GrcSoPrWHe
TfCPOt4+efjKRBpqxsUbLBl+IHUFFewgz+QjIzAehHcdCSGI7H8m/svJjYMIexNLUUR1E2KN0GTb
JPdfaXtCcqtrxVCiAnG8Ish7yCnAErC969Obhx/jEFxafIf65WpZ9fr5Q/blpdDDqzyOOMmlPwwP
ZGTpm1SqSOC4XNCRqnS9qOqAaWW3pD4sdX/UjDMsLnAod8tUvL6JAjUEuzWlZQPlZ+Vv1y6Lhqmd
xJ8/5tdDGM80JDn1U11wdQRhsH481joXmiV7z1PX1LvqfxodiljJOBUCgYTjM88sEwfgovz/8uz/
O2FAvOHoDrQrbi2yZuQQIkLHrhqtrM0L+iF/eN5+UD5mMTauYYBdXl+tqwh3oqokfhJNFS9Rsp8b
dNZHIJ/NegPBGgFBZHIHCpA1SSvkbbdA66reATW4xeGT66rM1lkSbmtFXbMtQjRDyEkSTVLFU4zu
iqEBppyxPsI5rOJpspbgsj03cOSqtU0NmnudqNBXbJpo855RjMBBdBdjLb/orgGXcFjdG9tybU4F
Uu5bDZuaN9/PIf6QX0kI9aUALoNLdsvqdAchL2DgsL2fPIZ1w/PaVkMeLsCWhQ2jKjIzgvq16SkI
HYgyoZR/SsuZ5kT04GFGR7u8lu8k/pnOORdWMaOvoXaQiGKY1Y4jgLfYh5GobBNzLkYSCpZHMqXC
e5VBkqc2NTy64522LzQ1ZLnrmGUcUZk/45aup6w8e3n60mGFNdFkTYZo1IviPTwq0VC6SbOL+Kow
i8Vy58ZPkCfXfPOYxbymPFqf2KE+ZbenTUwr1qN4T5jEpV7QA+rqzIJQ6McM48NbHVuhWxCgy44B
jZnhVpM3/U7KvZOKVW/3uf13sgWioxB6M+qYSfrY//3oJccHDVw0dczvR5Lw+3dXb0yFCmaU698N
ZbnczRcn3Vv23tBOKolTCVrYg5EctdibTCvVElhcY1Pgxvh5/R5eNY3XPljq0/a8VJzx7PEnF2Yt
FvkLsWMaUZG5BeRc7auniSGFl+f7StQCcbd2yHLRAROdLLOaDspgrg4mUAZZUiCmblcsa5lQPC3I
3PcQVtXHyv9UlZk12jdIE8kXF9fLkZhfmjYbysKulmVRe27bn+yBh2mmJgzrrkFi05SDwEKWrXpt
wkNuhnIgaj8vY2AvgWWyDvTF1q68W7x88GmCCvIJUjRqS/D6F+srrG6inrT6UwQqe8l+YwQWe2Ho
P31dXAgeKGLhzvK6N4icPU+vwNiS/Gmkg2GsQP1yhrFvw7pd+eQgWoeFMryxRGNoNcSW5KSCv8XJ
skrJPyjYMl/ywrl2C2MzFPEvyukY7W1LnOx5i6QG6m7Rxvf64Iuh3UKQXMT8ot1Nv2Bn0GhVJtw9
MyqhyW9FNM2937sXrXVY4PgL2e3lzfdTKAfwVtd1JZzO0CWM0MOaJ6w88uWvDuy0zqjJFueolcsl
PKk1aFJs5Xe5xsp/KvU1XSRuT7PMjV2XcM+l2e1Z9l8Y+0fdwIWEpWen3n1MpGYtxn5cRTU4KbJD
GMYC/BrdDihMYawQQC74InLZNXQbzDmpjawwYVvcm1ZsDbghNW9rETjmhg3FEzElc9fbMKb9aQQx
UJyBf6DgBr3Y5OfjzsNI5FOOpkrEtl8p1VA+YRbKeI0oLNMkGZ2/cYssJOeY7UduV5/2J3ttXoRb
Y+OFUd0FRHEfEpYCKc+fRrwEWTiJM1SeoFeUQFvgIH5glGyLcPUbcw052pptVE2dIHVW0tH/nW3O
GzGAyiJYLGyIxySBKa2Fq5xz/oeehrNJlGiulqvtd4DSk0ONWtYHk5uAKkyUyxEFDrr2UiRsF4GI
OlFub//BxsOEkwqpSFm0Tl78/RVIP/hLZQbI8TAgVlHz5zkHrFvb0EfvrLvxiitXfc0w9XAFBiWe
FQbdWy6WKYkArHz6ThGBtp822I8Muwx9/fggXXg2GUZonY0lbH6b2+hkuteZa0Kpj9XaMZWbP0vG
DOEt7SwUSLXV8XLbCvjbE8Y/Ul4gAAeddVje+CUWrchteujnmbEwZjfpiyasp6sPbdPvfHJUQSNl
QW1Abajwc/KPVNoNKq0HPB4ZfKZds8ADG6xxNp51wA+4J2+ooQ59JXS7SjIdhs7Czp1RHYt+nBJ3
5g7PcaBAbKBh5d4qt2gx3iUSkDw5Q04QPRaZ4dFZF8jxzdvHLa1xU/KNYPvzERUkKTkFTrd5jrwn
iH55CECzXtsM8NhDRn8JVWEJ3756dHEMIx88hnk0vIufx1NWdF1ajBacuXbd6L4yIhZKOgxlTbvH
KljdkoJIIpaM8W8takT4OSiG0Zon9Y8KymBOhsewnwcIr/AAvwT+qf4bpKqZJ2xwgxPOfb6nX/jx
6rL98Cn0vC5SkusWWYIYgUZ6kwart3xCGcCqEGO1Rxc6zPOEYvjoG6ReWF6E57HyvsFOvj4YFqL7
2VJ6o1H0C5XsI0VwBtoN4I2K4yf7Fj5XvRsJBo/oxBQgOTBbnJu5FWHfqJDs2NOQu1hmIRuUHMtJ
8QOa843/ECJpgvbqKO375Ub9AvsaQw6AtbFRk4NRoyYjkWhN82ljgAGTESiwT4mmw8me5oduzuP1
CIdRAeFxlc9btZkucJOoyxHOItAGsLZr+ieny63lcggOb73uRh+gw5ftCXwTN8mkgTTsoAHbsWAO
/peld6tqr61zuE44+sr6s8k3NsSeD82EB6gq+gMjqM/WrKahHlCDnAGnCVJnDsI0mk8el/NLJHFw
F+124Y/rcLQdam7HM/FVJ6Yu0DGO8ojFp+1dZ2weoHXAh5cdUg4vYtURb4AhSLJcc2oq6nk13WIE
duHyaD5AZ5ULU4xM8eQEkznkg1jG/KuArnFqDIaQX7w15m+djSrXByusYM+p2nROnABk/tNF5PgW
c1krh6sT+Ysvw/ZGrC7cuRnUJwilOHlvIvWTwu8FyS7gZJ5ei7x967+BRFIbkosKbLWULkc7PfMK
DZVZaZvzOMrk1N/TCy9NO/1cZA/amAIEFlQCSPNDr4Pn0eKKZt3kera/ZTQVFMwC9FiyUQyFYL1y
vXsPsugKJo1frCkBLKZzGO+T6QM8Y7pU9E6lGgWQ8iW/lxSlziJjs8NnqvqaKIRREOJajxWFEY8M
BTYVZOtiL3fb6ojhuR3lL6G2h/c2+sHASJtiuYU0KXvEBy+7y1SwA6BoSl41PO1iZs28SkyWbsDx
CtlyBdJrcqbxmaCLSL5s7NlN4t0mPNr2QDiVi34E4+YsKEKHQxI9XMCtQgpcMg5iBdvcO2+BxCqN
WxcHFnFHVIWMc6W6nxYF+0Ycu+x5+kd2HeXgjuKnn1seJTFe/Frz1yuO61GDaRFb/NLH+k79wGwC
aYOdSXlzbv89aJ36ZO3h7dCAon61hvX9E1oe3l/5+g1PDp5yHQOFPWlGo1dFKt+iMOjMidJX9O2v
bxIx6x9GaTcTzUD8pl8DFA6Bm9eJjEUAfdWKvwEUPxOPOzgFoMvRYFjZwR3oRE/HbWTrZMbfrB3z
jKw5uc9iNNzE3yDbM+4luWMPmR6iWvJpstj/pqwNonag/c/nDK6vGpp9um5LoUv5/MXtHXEcvY00
zXEe5Vb4sGEl9rn62w6MIshaeJHwA7FTjyKwtx9NaEwH0n+g5GOJ7h0HWEuuLf6QENRJZ47ArwwP
4wtGn+qrgAFhX4u9adffciXBvmknP3SShxbm0M9mMpFi/0J3xrtIUKxwMM/Pk3QZlrEQ34HecSo2
LB818lUtmpRXKKL6yaylWybXy2bOUXI6c/yClg6A9Gn9czrstqT9PFgMavXHb091neJBWdvIIPp6
z8NZULtJ0piEie9z3khSViAUnob1frscveh7v+xNPfuYzvu1hivdqUGfLzGmK+vCHAL4rQmxdDUY
D9uvJf/SaBXtNfKq/hrhv0Dc1ZvT/cfo5bJgj71X51EnuCUaP2tQ/1yhUoEsdQXeo01MNDDj+Tmr
sq+pqmpGGh9y9jfuDTr0/tgRWFXOZJYiNdKDVwgK9W6rsEqPzXtedVOsYeA7Q5nXYrDHxSFqQ5eV
QzXKE3AU1aC1tcgQ5sSGvMRtKfGLgPxEXgbW9x3u+Y78LYDGiyuvb47yToI3xXnlt8F5pij1lzK4
Pj1PdUVJMuyLgs5xN9u5g+Va7AXRyeLOy/UremAnsEP6ZP0nvTrK/VWzO8Up7lm8NYO3jtezWo1c
sceMfgI0YwiDYTB5mRGKXOQR6hFGIjvJF4bD50d1ZzJiwI3S6yvxbHPZKBDR59R9x/Go0fSMa7pF
K0Wx1B9YNbbCay0MTmpD/x4efHxRN/Ihi6BNikXDjUwNd7UvTSn9TuWk/eDK8QzPsYK02cVEqJo1
kQpzaeuk7382LttkRRpoOFbkZb4khq92A8TTy5wozt2eyeVHHTT3U3F21iCLLeZ8iTZwuvN5Knva
5TutbF/qy7DlwXWKsFEGr2o5IiU/OiV2hB+hKR4S+XhXICx02mJKuDWqNr6RdW/l9RhOtr1rlNpK
5Mo8MohqUFfmaCsDVEbt4zpIvA4wj+D/GPdwcnRvU5mKW5F41wDm/SJJFVLHeFM7sOVsEMzkVnVJ
9bpm9Ku+B9FqlOzXUbWHB+mbC6UKcXur4xhLm0L8KjaAwcInojxn7RSbKE+RvFZdKgIAJr6kj7j4
ece7EK9D8K+3l+vKD3El0UsaaLALa7Wh3LACI89qths1NUo3GOL9alVlQil+3BWIzor3sbt9KKC2
zKQ744DVYJExW+9NjtZv5AbJXfV8M9404lcyJ8+zgJFEzn4Eum1zgqTm37FpD5SWcJBZxkZEpL4L
rs7yAYrcy0yKirJb7oR50tm6JLu3J9Ca0kWRBGbkB0Tki+MFA1pSkg4GDChVAZr9THBQp2hSJqJE
qS+dPEhc1Q8a+w1M1DTmU++5v8LyE6lVVSnxWUlOVgZB+IJf4dXKiJ7EQ47L1QFhUP4mXBL12fZ5
Z/KUDFalQsbnQ2CHgQyirUSbBpAEtFAT05UdkqxiS/olrsaczNA8Hua+1S8vl+1rxTGj9vGTeKvN
xyp1kaW8EARRAO29qTnTntCvA6V8uoj4/fgfB7F+3yY4Mq0y9d7UW8F9QsEyVTbZ+wQXar/HdECH
wRVdvDNLwezjNs47r1c1JUVDAVfsAeCqDnEjXPBF7v0CylL2QDHIbmxcFT4I0HEweB6FpqpZ3eC8
bIRkeaYhZcXhVJ3ZYDUcjVfqtihdCsUY9j/p2b9KRPs37dHmAgKZlVPNZBr48FWvxAfOlOcW2Cvw
MxzznTDW3AnwTtBZq23HGxVPUGygBdwWeQE7nAlTHYNiGPVTrUsOktedfyTz2mBUXeL0H8Bye1sL
dSsDLsA9pIZ8EDkhr2LgQl9JmfltjIwfnKdEeak9yk/2z0CHo+bW7GOSZvmxFOdDX9Q/FYPVsLWW
SUJXfOm+OLlePEYyNHm9T/pFiirMsvcV5ceMJRipJRRD148OC6E6z9RjoywGD9/2WTIQmOSkIBJX
9VJY63AfTDhjaDP53ZtM+2Y3TellVgHs8x1vv2KMlJ0AnllE47PeieLfeLS/N1Pb3Oa3070Szsw3
5Hx9zpc8ENf5mH5QN/qw+KlllpPb3+cLny1NnxR9DCyvuCj8vyA/PPG6e3xWGJxSziFK6MLA5hzG
Kc4b6czu8wEpXAlDLAq6oJ+GUI6aV272cFb3aaqu6LpIM4Ff11fqUACi2fdeR5d0YjJxgDdYKbB2
kjgSKFDJL/alJpVX3Yzq1/qSJCSIQAH+g3vnK28wD9AkUzuW2oxj8QGqtnAeO9JTp3Qy9BIEGymB
9Z/YZQEPEHkWYVjPsRooWsvUYteYpNeraRPojLP0gwQACnZQP2Hn2/KKcz+eY3jua32ueJkZSKU4
R2Ud5CA8dZ3mBacXEzivAs4hBT5uNdxZ43jucMn1domlLjiCobUmCoJ6Yfa9e1gGc86dBdiIr2tu
8l89Vojmlp5b6yWSwNo7xybNgMvDWymc0pXmv6/v5NQqxIGXdDmlyXOiVSwtdJrcgITLO8OkLBUN
chyrucGky8s3Hom5elVbaUUlD7tvqw7Amy3i8NlVtbhJd8SVagkz8NhC/E1Hh4yxgu0FZndLzMmn
3FAk+IrAafZ/V0mGkgIS8Jr+806cl6rf4heAfxEavMnLS/06Hcee4AHrOLNlyynqqWtTr/llfiVv
E/WfeDGWIjnbUUhcNuwG8NNClyOHeAq3nPw/AJnzJ3XptzvYPgx8vk5ocZaMkEN0FEb24w3ICmxU
2JF/hBIsLCVtN4O1aW+U8bCkfUnp63AbwOXI5toxOVpv7DGQAwFwM/4Q6DzZvGIPrvileOb5ZKv7
9oaGRvzEq6NJCevBfxLukBGJVh/0eyBr+o50WyTx1YN/dMutmLDcAmmLrCQDae5peuNvLpeNPji/
SbSRL/FGwMMSQKw+PnCQDEQfZDlH8RK5EOQtissGlWMLFuVVbGCdPDJh0+Tiv+LuJLZvl6AHTYl5
J2uCzW3NSnbsOR1o1sorD7x7uvOmtR6eQZp47TDDhssVLOx3kaL3Hd+0gVd98a37cp+/vt67zj5z
KvpTj4lpbCyxN4V/qHAf+5jEL079IT2PQG4bebmF0huu8OaCVurQEIcnZ0cHOG/Quetkqz0DtAZB
Ft/BFqv7qRyLOJvDnEvOE7PYgZ6thMSBxdHIi57E2LcTEWQpvLX9PP7s2F5Ngfbk6n+mxP1cpNnv
8GF5mICRDdktImX0OBXzWon5FMM+gufN9rufQBjsMjU4hsrMKFOdSPIH2103v5atsFLJAUUCeKGV
JyUGpiIiziRdX0J776mcCl62wa0mvQ+Rh571WuHDW6uhxaCZdz3vVg70N1IN/ZyeVtDSxL7OmGan
BjveJtfjPeXdPok2GF5ztbdB/yqel+KzTfV9XQyQgzCIUafttzck9boQ0vecAcHDMT9+YtuSxOrJ
PKskMG4hwvW/xmfjiHb3mHPUS4awtmPx8J5YOOGPyxA7QNXFQsMdtfIkrBexiBEniawdkHZgru07
1Rf92BHIktsZnd3ee7LICSbm+lfRh4ep+//sZ9vVW2F5lwpsyiFeG9keiH24/SqsSr8qq1UDX/QN
+CIDVzDybxk+exZLR1Q/WgtK7QE5JopfZ581uV04dNblTcxq65htZ8ZhqyMnb1JjJItHjs2/hViC
/TS4Ta/6Be87a1uOMmzRuPOLX87X9rhHyXkIL0b4fUW/p751X6YJe8WdCiM9Zirs3xS9vvoesUyC
2KU6oYQQzYOOcDqcLqVby+Pu9mx+e+Q95jetflMVxumOKrZ1piappGOlEjtXAsvzPg/4nj2qTcQj
gA+4hYWiWsm1mBza32wjR6FyA26VrxiPJuIRsdevAx0BsjWCqfUWEukqTqP9wlo1vxhTAd4yf4og
iOTt1VVDEmLhfP/LEnl7tiQHcN/tcWiLcd+XbE+0U35FeKFwFZ7AgKZ/NLyYArcWMRoyBddSc/IL
fNSyR6qTyzQHrfJTKQqFH39U1SA09BLkAgGZKE2pVnbLedCtuLCjVFw1VYLW5CLvzT19n1HNu4pX
tXajUFkPdcYu3Ap6RnBxA86w50U7CH6D0Fl4uuZB5NjjmdIUmTQhvIh/e6DgaApYYdezVS2hgEao
Bu3h4ozqy2SvgKQJdGjiJvCDzAwucsgcTRHPE8TkqG7Vi+RPzfZWWithuwlKbuOSyIMCtt3ouKik
SE78db9pCQ6OEaDgEHZPY+rUyRcZMlsmxTEaKB8kWxNwWV/6Cml652FTUDk+2k/b3lNYto0J6Iqg
MX2Q9ZxNDGxkBRthykHZPkJyhoOU0k9S9JYkZUdp87pHeu9GWiyis0XNHKgKwOtUmZKNVHjbPeE+
Paj7AFkvXFWZJAKdDigbgAI8MepZLFTOZR2f/lIo/w6BMskjzJmEhEQN53v9oCAbnZNteM36fTnX
d21UtdRN9thpmg0nc5LZ1a/HcxkdWJTzPsNMspt6DQTml8ehi1oPaqxbY/v6CKueAnoANmWPGyz0
Q2PL8Md2t7VZGbw8c+YW5Yz3QDXMIwAR5DCqfhsAk4qTfJxuBVVbH8MdjrpC7f8h7717nNqLVXXz
id2P/XxVFbGoEIbx3p5cOD/qnDBkoE7sfqQmdOyrcYLdpEbnXQWT6pDzeqGZZlmkhWvCGlECkOW7
O6IBhx4lqV9LJf6T1R4ZyGezZMt2orgDRpcV5vfB7RVZDUQ08vztAZ0UK8luIEROTtAsGh18fw8F
4mlNkzlPXtK9xe6emNG6Eriy92M1WjIx7+8j1JbQl7G6k++ebI+fbmbS8G4xyUCYJUPXYazUKRiD
MQ1PnQ4rZMQy4/vQ20BSukevVJ5b/y4DlsHThfII1n3XSWhNJEokJlOmrNyEhYHgCXf6f7l8Oc70
3YQO2pooiFIzaJVT6Cn0Ta8/VrGWLhZjqSPjw1LQVqZbqkVfuCWoGm4ZBU3Kp3ERusl/9tEGlVfj
MbgdUUaTaCj7c3A+/1VkBSmlly65wnMdc/4HW7oel24lBCEsa7mdtNdh9tLn70FGWreDzLC8WIlp
mRfsQr4qMKBv2KX6IxIjLnmTsdCez1amL9CTsB8BSWZoDjStN8ccu3CPG5KLN8XcgWMlJQIKGdaK
H2GM7/2MwlJqQr2FegO9lg+EMG1fitG8cFP72t1thvEo+Rrh1f9C9jKqR1nv1zluulTifBJVAWBr
hiHzASLlmfPdj+sg14UqOmcqxJk1FYVyOW1Ww0XuwZNLVGXrDweFqkZvGYR3Zi0KBkID78b0S+VP
7pIFZaYEjiGuEA/F/ZsBf6d5F6DdVTnoMUzRNCDUsyDk/IlPOYyFHxBBuy1HlKw8gcx11JWFwgW3
6pBOWaTECaIPW55XiWKdFzOLc8gpMq9QKPL4bR6K6FJj8UawU/bzHtYoxgXeEgacELJpxQWpChRl
LMO30R2E80uET1UxDjaSwk1u1BWrD+dxgvNboCcqpmnCpaO5rDOQ5ALrD6hTWhiPZ2EuL1B2YqmO
DLXKhFSrZu0Ij/P+PDGdpxc6zezV5iIOhLP8v6upNQQFZBifwZV+QaLzhT9+X88k4yZF4j1tJK7O
5lkdyZ6JhyfLPH2URzvAHt1aCrtVYDF4R1Xzu/lq1MYZ278qEwM5443Riy57UlQc5Yo0PUMBnM1A
izvhy1uvc7ilBec6kun0+ArkRIDHVN9jC8AG44LtfcHGBK6MLnFYK0F1gQUKgZuxQ1kK96Bi8svI
z//k7AQJX8giURtOGzdvUk30WTwLX5rKY81+uW4tW/aAYWNWl4MVGan3sq9NPFJH/7hbYncD8tv4
3cWCg34mS7266t2qye7lEfPn6yNxWm8bpSfGdGJUzAWdTMoVmjHg+Qcxujpiy1gY18QcU+UY7ltg
w4q6OFCEwFRirrAJz3CrmHfE0m+VMQUJ5Q9NfRpLDMGEsOjJdQMR74Xi9majj77XRPlWyL/ZRWK9
eksS90OYhQ+nTi+xBGq4rzvVY6/SceX/5re+Vs89AragvTM2WQkPf6LCzvNkUksu573aFIagi3lE
lymJuvJdjMPaekSvZkiKTe9artFKrw5DG8c+6RiVTkbh2jKBdrMu9UNIRc/5brRCtMZfjqRdBJ3M
U981qkiRu6ymp+5HcPe9l/e7GSsLsYuCXqFXLvAvw8xVhfUK30CPeZtO/lzAcU+2EMYifRMvfImh
vtATQq4loUyQ6TZs9jHUuy1zZYUWAHjCYZkE/BMpkfhgpbOkOrzgezMQZXNiGBNdVkoUrFZzSCdX
HRxbXbm7x1PQe9t1SU1AK2AGNOlGG4ZqhTvZPEJ9b3OLbUWi5/zJplUUBaYVQD81coQShCUqJSpC
VaJPJ3/ekBeFISvvC//gQGOoo8daGoe1NUkB5HpXrQjPhWBMoV/oxqL3vPjVz8BiU5iKWRMWwKsU
ZVwcoO6FaH1zC2ZGdiBJwne3v6npxv8Ir4sWzNunK6MsJuNt90pT2vjraeXntnuE3bj8Oj17rx5j
xbz46qNZW9VrGt7fa2qPBNKkinPkVfHvGyC73Mdlu4OTui5RLz/grIzN3qphd2f/u2nYe1AU8UVx
1FsP98hYnnh1cJYKkvvPdqN3KpVzvwF7Fmn1fEPP6mf1n8Wp+mfnLtUtvAWP3vCtLG2l6VRxT+eW
dgHEtYDFndrN+yNIrDCp3B4anTsTFZnb1iz0fvcjmok27geadqsGGggjMjDgtu4tVmFE4uj22gRU
r7Pc5oq+F2LhXZV83tgNEfJqQ4jzFSIefqfDjeUtlDMV8bk0OpHrO7GSxWuGUyL5eD6Ae8KnBxhf
s31cGz0538oj6d1/KxHrNfvwgagDg1IN23XRqkaTl2K7OzuEnsE5SuT9uZs1v5WJy6XObOrf+AzI
SYXeYdltc4XjQHIT7v92gVj8sSddVxZb9pwcuVVBg+rp67AjdyiiCu6xp/A8CYT2Xcghlnq0uux0
kd+jwqttfukKCP/p+1fuvTyko7jZxUEq6IFDZn87o2fRY1HXrr/LYPrk1l1Wo9Kz0DbfD0IGJ5pc
KsElDjQEUUNZsPi1joz5ipfP7eiaUSJ/29EeKEQWL3qoeoeiZlaZhg0NvOZK/+nWDOU874GjjRX/
xNkoWMyuJbdNeQM1vM+QDg4RkWt+KgyjDAjDqAvJmOIOSUJQ5FT1f+R6wIS62L12LRvfBITKZkqW
e0bPWne31T4DCBkQA1gtO2o/gB75omOoAk8vlHH2iLDHkmNWSJtGok0tuK3w5xmMAjPlqUUL9p2G
jCb73c1BFbOaeW+MUA3yhTAZcvgajmfxsl+BAzB/dhg+pzPb8wIrKTh3fGIq7hW2NO+QykBm68R4
2gYJDFjxqamFrTF2BCxb2WLicpMkqXHzHr7Zl94dr5FFhGq5DamUPdmCVx0TR06bBvWF4GUnkEYx
+vnfMHWhoeWlniQfLvkhdNviKw6D93EzYMyBkfdkCBuBovqX4MRlWcwjhXTRE9Dh7JSsZuS8TFJ3
9L7HcK/HPGPybjPAIijK75d7Le+4orpBRCY+nrxuqFj+RWHgQ275aApspIEJgRl0RBuXaQfiJ9j1
JMh7F1Q4BwG2rQBZvl2sR5mQdDQ7sHzftp1LC/EFSyus29trgKqMmaWjf/jaSLwRIjNQroF31G8w
GgmQJNlreduJB4P/ozTGOfQyzJ8KR+x8hBfVfcuLlqJ46Loq68/KpDAZhgwwJGER3vs+P4qYMLr4
csSvxWa0YNUdYG85ut+whmKK0FwJGJa9wBxlfKbMdTwkUWQyl7ITNUK2nRMy6Tmi229x1E7fUuB5
Emz6yo15Cxnaq8fF9+C7UwwmPV1BAa4p7zGA2SIm8bLN9JZlb2ybVdkq1HYe1sOx5zUt/Xovur1E
AFXoUcP7LA/AEakcOWfujemBvZRRizCo0x5NKtdrCVDkhnks/LxmC6oPfGzn6lzVytZ7MNWkZfPS
4GhVZLzlSuSk6QGg5I3qtVeBb7GMDLd8qv07yZvIqw/wC69fR08oR2VBbfNL2aJp9kuh7GZlZJd+
I7Pi4WrdE6NlkNJfDbyuT3gWvMu2V0zUSMWFm3bBHxLHKeMA3i8siLTyBiJQjPpK8J1n0I3b80jb
Z6dbmiIYPvOS9QAhnsoWvVsB8c9LbIPZrsZDta0MRZbhDNSdWdgqD8Lt1ehAxI5S81iz76U8XklT
VOpLuVwMSMcUkUBp9GKx71Z9CtDFOGQ3Ryo2ABbnD7AnnJoZeJfYq0IqWKwVWZe3K/IK5AHUBFcy
BJ0F8QAHznyaV6Zr/kP8CwnDJcKuKV3EpGVjG3x4b0JVvPcWSJUQzWdvCY6tbhd76JXLLJvLBtCU
hbfSZwPk3hNxf2hUeJ1udFuk3pbcddpqrXhyDFnYQCY5aoTGPPVOBywWVivZaGppmaPPmf7zcrJT
F1QSC4ZcDbbE1esC/rV9CyOS5ArxeR0PECZyPIrenh4HNvWUjvCYaha3OA/QEU3mjxfy+2ugDw1e
VdWGLLRPjNhd8Wd0fWojwWymKmteu/hryaejRkbFr2RXXczFSFW9qM3JcjAyFKYkxCnSKauM8VFm
OoUnm2Yj8inVWPje7X0xs/4DGyl8A2744jGAHyaFF9BR5EaDrIXMcAOPm4p+7qL2gaxgmrl4R90G
3WmJgTvSfpA76AJOBcPc8ezXcQWNl3rbE2kmET/lb5CzYHWiZfgmnVL0UHOVfKoh4HsWPCH5OqaU
aSgkIxVlxAXUuGjXeRHNOwOpVIiVZym3HTlp1sXrT3xqlmuOHVDfycnKA1C8p2yX88+ySh26iCPP
tGpKN0s8gHpmoWR6/DBerEM69X/1QA+ah8ht8Q5nG+TOEB6Qf9PHBcyQemsYkQKUyesYJJDKqhzE
PEXtOerxYiuTRmikwp6S3cJlYDhXNimcgSGxNHboxLgqb8D9zakBGec1hNXOELsJLVnIQ2RMSeGG
QguTL9jBwvlVDvHYUOHJj9wJXmuapYW1yZ9io4IfPT3sWHdcirpDH0RAeDp+TNl6sDcrYhFy2I16
TG2Yn+qAQopiouPTn/n8FxPuFQekFOJSpI7IyFLfxUC5ZfBLfa+C8/UQwP3pTkKhRe5g8q3okVuq
0hkvZSvjETd6Wa/ADdlXACu9ZSVmF+3MT7pGHDYitONSyxe78D7XHmoaEQFHWUviIjVWh7J8MjcC
UfnSeGsydAIQmXM1tgheCxifFDjusOGMK1W++BGBIsMieJlUiz4jFUgiXMDpCpXghan7KVE2lpCa
tPyi5+OGURssaA5d9dtxlDdyeIg5vqBlVgcwVmfTzFrNhBvOhgvyBPDsBWN0wHSr/TIe8HT5ktRT
l5FBv7F+OeZFvDZv+imuNgohkWlp7aVFtNvrWLNNvENTgrpyyivh7X+1am4DGwD3tg5uTe/c2K2E
Bgh4cqUMQzHVq75/4Xjssy7IzXLfTpvAAA9RSNHbX4Uk4zCtIRKVnpOANjwoIUW2VLw4gKAagpho
TBNnQ7nJH1HDp8JSXomyOcLET6phguYsk+RoBkgZtp3fmZjyzAXBeOV9b6qbz6d7jtiZJuUY6l+f
j1I4hA5KP1AOwtyhVGmBZ31M8xGou1a/qbMYJ5+dBp7sXoA8vB7bLfREZHFSwrP0L67c7VG80r3p
CnE1LJZ4AG/5qiPP1jvV4D7nZmwl6gawZQiAJUfyzvfwdt1B9wt+MwL52sUIo6G2vV62Kjy6CctC
KtSDJPiDjLJDHSPJL3IN8xixzDdnE2rCkau10q0rju+2N9rboJ/ncz28jIUx9fxhwfHuU3pEI5IA
uAjC9A35BgQAduVp9NES2SjiCK54uaHAmvBL6f78BdbDpbC3082G3ml06ERNIEkB4E9O6ReHNI1H
XpmytYbEYXSpUhfJk/hljM6aH00PGmusNq0ExeTRZ3FaMktmkWRsts8idLfppV4cHpVB0opY9vWk
Rb+u+Y9KEEFfpTzOtXkGuY3iHaeGHudAHRU1H4bRhIeUbO4yBHRNfGga61fbeDik2ES778+AjT6B
oCoQq09fn033bE6lf/KeEegSv3vL3jRf6G4muN7rSkxcvuk4iajjwj+q53xIKMZJSmDDzKh54NUw
4YekdoOfuZop//4IDInuCW3Yg727E4B1gL5/uzfktxFAPeSzoEe76vLqo6eDMMkqAKVJ3HLvnYBH
EnTxPHnkN7kr4b7ZgDY7Sny2OMexAkDoejeNNyH9X1nOSUp/L2Q7TFzQSKUi+dveK73r+Ji30PFP
ITlToQsO63zfeRmMDICi+Xj7Kl1DLsWvh6p3u5HeBV5AT4kA0e2QdiMzR2eX5DNQvgDzBOarlUyG
GRL+guCK2BtAeE5nVKBafpDEJhGzuYQ2CSZWwC6hZvcQPLvFr9Lw5GR1LMThB8IaX9u+gABVrFlT
cQ2QU+Y8SCl2f5RNjae4IG/CvpmKfNgw3HE+G4V0ueHvJRQlczpbmzXHBrvCMjZruTifFVaYB46d
6qjtETeAkD3fkwz+eslnO41l0BoqcE46OViMXq5kAAiSiedhvmSpsJZ5akmvzQ/LdC541g9jEz+w
HyJ81zkhuu/Dmz4shbbyvP6oRVCxqXWAWZ/s73eC03bvw6bMj7J42b627GRY8FaxuP/eBImywaMu
cqHMS3XDq1HAm0KH6ACd3CgmaROGXH4Ji8ErfquECBP84g3NXvzojAeFJbMv31QjMfoxRXDInPgB
vOMBKkedLv5aPeBZiHB19+uBPVc4+zB/eg2LZ1h6NYjsGEC9/zZeaoYrNWAJLk7ImZK8kvdnOcYu
2NET+CP/Ag44zsHxc/MSTEa/SWNrB+sf3GyV0pD3+1+vFbGMPItprGf5KbXi20+ZDhXJAjFVoGCU
Y279k9jc4TC+CoPC8WpfTPqhK2yXW52QINR4MZohyovYlpAunurKA6/Fjnhut5MGhEOWEVJR2V9e
g2KvmnIRGjDdCSjwpZaRR+gk1HjnNtJuTRwIupm0JvN0hjsazVdEQSEICbnolbPR6gYb+6OKO6WP
QVyws1RDf6qSao7a9rdbjT9gNdVB2wjrftWiUeXrwA3yLmwdD5k1PdOXTjLrEn/cEmSPKnb3nhtD
Av68XLhVFNtZA2Y8dMQ4mXtTehciv2LT6PNRPZOYsfCaHfRYGCjap0y49y3EIkXjSf09Agg7jBkE
Dn9zrROEAVv86Ki9pK04xZwwZZ1pnl83yH+phaz+IVLjtTmCTHAnGwYg/qvuAJjfs+A5DfBIphu6
RuiSX69Zj1lkliWyzAZz0KFaHsf1M1iuEIp0fwZZYO9lHLh6ocPE+iALUPx1YuOur3ZR8T9D5CQz
13tITb+rfmqvy0oYXWdKpQLCcefeNmgr81l6uIthElfHp8xL6Z6EuoGw3463YVzK3Oc0Am+H9lXQ
iOG/A9oZPS1shYYvUlBqdHWGRfuk4z517VdrHaDKe/zIXQo5vlCHd2qJOarZZBDQqvyCHI8mBX+z
xjnVS229wqg4l2TPC2/ojDmoHsEmMStTsX43RaHK7eBWxvjCTC3e+0BuPF1SxMYXUE2lRzlC/8wK
EY2n8KaZ9cMp23LpIrHBibPVDYEH/0i3LDR7gMlHgdWVJltCVIuiVPMXfXs6CsGPBbPGlJZ8YTSa
VG8SBZQW+IAAH9OCP9amAj8Tikd3PkULDRCLsnjC5ewlm7ossnK04YWpMcLiWRlvGaVFhtsen/M4
ynRGgFVd/GIcNJOJWYRvyKhj2pkHAQqekqQ6xKBONrLNGHv6gpPau9/I+8N0kKx1KrHbRjS0hEPd
mDLaPEDFa5By9dZb9gVsLjIe9WuwgSs9Dc1oTJDMTP41G0BfnXBmktJlfRZQPOYW1mJNUCFOjYVt
CBJRTVO9b4i6bptGvbN6nj3XHfdLK5WziqfnjX5TxAbcNq+/K9pEbDJghoEw5L4vHQTkgbYNFkdR
MqJj+B9dyBSA2GbYetgnX97AM6x1nnMgkBGn5RzUDSJ3TpD3Lwm8CTFTRg45A7XBhDkQnH03imdK
104flUI/u3FiMebO+4SbyUmtx3rBDisExBAjrN5N+n0D+iTKyv7d6zyMrOYLgMQYZkqrL1P8je3j
hpZ7n9DbqkAg7mfaoDQTeWOU8OSaybfrhKXzVnnqGv7x0kRCynQJV3JCojANOz9Yl2oor173eYEB
BFTDHs5Hsaeb1nvs1F3Nf2yoKRi9TzpD/4xQCTbMYKuHkMtbD/F6W5I6CvfG+nbtb/TVIdXevRFm
Y0xIwqQ93FHD/W8g/Hio4tLuZR5okdAwTBdvLovdlwgfS6WwHP0bOFuYVJGhGmP8Ejlpf3kdZbcx
TmvU+IaeJJxPe7XmU1Wk0TwEbtuNmimTbEY+ZuoVlvUemNAxFIHVt7ZtXSczYENWPlBGa2ckqA3g
rPMgv7/gSvhDKwC45AMMyn6v0VBosWjl/hr3D1QeFBRnXFKHhLR7P/kDLQmi1wjXyODvbnlhJlQz
oTiWxcWd2XJ3i8sNEDQz32hXqhlhI3p1Pux9M3EBhXbjcSLrfsm+57Fg4aMu3yJJFxAlmlH1AlNc
2t/t8BJX4rP26sW3o3d/ZZbKvuNTexoWQ6W+QFnGECDMW9NI+3lO5pucQE5pCiDFoztxv/rMwKMf
YYa2Loe+va20PGlMYCFAr+/5THjthn/aQU2aqPrs8SVVljdVTyXM/cRZRLfzzstF/8prRq2rbRTh
nTuXUDqjWup380T3GPCDJGGw760QlxoWNi8RQo8Fja2LKrTwyoV7LC6Yn+wScB3zuNOHTTcTRh+V
e9ZRL5k5hpM4Fj7IP5gM/CuKFTp+wRng2ct2Ez9Dr6srQM5bGKFaHYe9IeVo10hTpp7DzPqfI+3J
4mKJ7GQccnM9F2NJVQQSNBhN59HtYo/5sPywY2wM65cWFeEI/O3BkVbjMj72o/i/L8uobhjwKioO
BJ457LPIAkS7OSQ3GjO5jWQ0yyh1hhMN8KUJgfcXAifO2Yq2pdExI6qPvkUG2ubJCLJUd/KPN5Sh
QEIhrcW7ci16S1Z73Ae6uQu+OVGUxHKVM/DdiDao0VC1K3+WwtRXQg8w9scbZ/c+o6Zf68+98fVH
rFrmrhuQxoClyjDbdv0tcNvM7etylT6ygRYnMF7mquDrQzLeEO2Ko4e10v4HSyMEFYo4Oohj9yA6
5V49hwGK/W71zQGvjgRYeF4LPlkKalQRNR0le9epWeQFLQfTKtDSUm03ehCevGOtn6qL1bZkvWxR
ES+wXojlED6gAB0KGGrhuKnNifZccKXK6TjZ6CMhcSmv0cLDC4134nH0V6YSzcLdD3nyGZQ3xzxS
ZduoCBAkB5UVHNyXM4BjVK7Eu1qOyH+BznJBkK1NunIRp3tFRDiKm7uZwA3k2L1zoIEdRdOv4LVr
HE5Q8sMTH9icY4CjDUbxRiGAWwpjOzcwMaesQ2fObcZWvfeT4rJnvdmNLX7h/Ouet5BR8J/nSm2E
IufeMS3QZ+AolzfDStNIREo04+iKvrasjFdYcZmPid2TX8F83xUKUkQJ5vEHk5PKzBOSa0sF4Rsh
/bEB6uz/CNeNESV9qn8sc1FQNPyb7st4FGl6vCJY8Rju3MsGGPg8+TQIWsCPGzV0zJu76gayNRWR
HyHbRDE762srQejojoVzYWrr/WPJ1aXYAw8r/Kv/VOvrJ3tGBtYa8ByETSGd85yBqmoasymPDo9C
aKXB3Cv6cvJnhZRFsLncbZ7ue6nGcV9j1AbouzpCnQ8gYmQKL6/PHMtlTEsdj8/W/Hp2DeefW1LE
onU/gTqE4IzhttN7VA7OKYsPMHExHr587XjJCAQwnUtF9nsh107vZKTwV6/xCRDIu+D9CNrACIek
croO5Mc6jKt6pR42n9kDWndSHkjNa3zHMjwI6DED0RVENh03Ebh9bIWRZxvjBkoD+bVmeWzIOvWJ
NSYk/MiMrJtXQ0+XlqS+ghYnw3wnJ/tdUCJt6U4QCLQaCQAZPRIe7RgQYBCCTbIOXRWi0H6kavQY
B/rJkvPlJHxKEzh+TptjInDnaPDCAhvHBLtEU8qMJHbERi1BmtRn6NyHiiUxwTuMWxlPyuh83F61
qYlcnwn/ZdVpDaveMHAXK8Pye/e0X12RGH/nA9Gg4l/RK7iNP58l8esm4KhIZwfsliU6k7P3ozAl
ju5Dp1w8fg1Ha3zN7ROfiUv8DfkGI8XoB1b9Onxw/zC5uKhGzpvnEcFHRuif4qTYGmoRMXdYzweQ
TSWf4n7cpZ49aS7z/nekNHw/4fZKqy6R47sZCeY01rvW2XhwxiKzqA0dIuBR5SFuji+YD1v5ly6t
MqInmMJAKmm1+i4MasU7Xixy+tAhRoqHIasGuJvTq1TnJjjKv/TPGavXsrCXsbacRrT7vwf9AoO6
nQpY4w7TwaIB7vGH9z++3guGIXPYgsqeC7uJGVnuyCKzZ9hrfil2g5QGf3Zu9VY4iZC95Vc0/9/x
E6ORyXuynCZ5V8fy8XJa/zCpq4z3oHXtRPJNk7j+ifT6HCXQ6yhGVuZEE55DKB6tTFIObWgYYnqm
fwMcY62qedfYRzDn7vQDAZfj8Olls+wLrZSxF74O8bf7rmRiaLdZNymoRpWILAbtEdV5jXXwbc+8
futo880+Pbc35hBTyIMWbFg6VInW72UKytb2mL+C8qK2MyEpQOu1pl3Ffj6pj6026pC4eOEQYb2u
RBJOCqv2gGBmQvfiYC7yToZbNQRcXyS/koEJkKkUJUPox61ol+/sI90/GTMctKDHuHUAXsH8Y7xj
p2bSKZdX0uyllAvD6Oh3/WwYyVK6GzAwBva5q4VT5mASuaZsFzzaCAhShtoP8WVCiHZWiYNCGQ6y
TtPS6QtJVSebNAjDYCagDjhjjLkF9XyvLx/BwAg95tpsVjCwDeWrAZAtfK5OdCcO6Ms4BlwAIhcx
NNi4lWJC8HrjtHApws6CNErwZcYe87cgM/ymXvQGH55nypPGdQAuMIKC4a3TddUgyjpULsSItpNc
3EjkzzCGNLmHWcbb4TqPEUP85wlzk1jFhGN7jpwA0jyrobiok/ayVhb5lsbHYAAKtNsk367F8kUn
66wiaNaDrjH67ozC3/9NVYRXejYkbz8zBR2POwQALwrI8mVkfTlP5OO95lPFPGIRusX2KPwbzig8
ZXIcorKLfY3rYRa5AiaUYhXkkDwJoqgypnYUYCbP93nvWX5dsogHVE0qLQivBfT9q2Er2djH89YQ
PLSOP1wA9eUn3PJ+5ttSWcQE7Uwp0Akp2YQGUowpPnyuXGhDxTGJoq/AGgHXR9aYw9VNFzR5dI6v
hHv/c3yeWcCEbvT6UFygUnxYwqy/jegY/sey9EvzkdZfkqPyWw8Wwm+ZWkhWeEp2kJZng1k8o+ZA
MmbNWId/kDBtXzj1TqTXUwT+/mz11BkJitwfixOmIuYmYLtBGo05mp7JND7thb63BKWzoRajBBg8
UCOWaMdMq4GCg8JJpY/WCcrw+op8D3MP00FbuQeJtfNs+LWODfzbqGdA3jgM5k0PYr0cVfW3EF5o
XQGM//YdFUjadyG9lyrygmpOzqJ2Q07zdWXGNInvTW1UWjcNTovianVp6DK8Hux68els0XWX1WeZ
qavAjE4HiiQY/jZdLPSMeSQewXoCAAVoyd6pblkppDZg6iLzGG3fZReMdPsLAoegQnOmGpDNbUJ/
xHtjKzpPIoLPoTRCroIvq6Cujd6vPXCk0UDC73KpN6fEQ4CdRUtigd8fVVCIEv4M9Kyz2+VSRWNs
3r/ya2nLsjXsp7hNwjI7IkZO4LFMc91HvRagUT+hW30ObNydQwfqDdv0nV50DEtcKYdBheUyMpAz
Uq27fidRCq2JKYlfZfDMoodkZw2Y+HgYg8QaqCLwophZduDYhUqHvPt/8hwOU+p6/SnfHxs0cqe+
Y5oMUr6ziGF4ajjcv4wFXSv2ndcpsehEBnKrc9vFz4AfOjpM/3lPkiWOwDxonM0dPM80o58Wx0In
a0OyR1epNZn4mKKzV84sRjfmfwC+8MIa4vUx+mKyBafoClIu3iO11pgrv2fP8wmfRbAPfWEjiICu
bHcMR766d7mqP1qT+N9U23Arg+bIzUb8hfUpMySRAmcqpqQ3SRR/+Y51/vMsUDlrLOZRMYvjDCvB
/FuIseDV6uMOC64bUrnSNhmOFtOz+hOldvj6lWMymdtEoqnLsbSalfNEjS3F8g6WTCFRc5uVMy7Z
8r9D3OAMe2fVlb7pKrTNOYht+kddNMEuz5EcQ7NWgQqy0WSqMlpLhyR74gA6doesLz2JQ37yxHw5
8mQqWyHqfyLVbVYvXvMRmkCi6A2UyMe/bZFMi4b1IkZ+wDngdH5of+utlmK4crMPL3MEtA+MMiFn
8YvAHDx+A5UCN9ow8VLPzU409lIKDjEmfFMoliGzJ9pTZrzDgydgvi3b/RDyaxE7i3FNxTpmDNDL
KI/FKN4x/pZI/RkeQ725HqMMARdACLMh0wI0CYxA4/Pe0bo3s3T4pHe9juAda24VElkJIs3a0ywI
RNFwVoqWo4my7x+gpDGne9ZGSj33Ewy9ZQQeuQ7tTZV/PmRBw8bSxzegJxjRh/7eqaggSnbFdNIt
0S8acOiyE2U6gIZz84s4voeevxaNBTPM0qgJI1m7jfB2F2Ic1iJTbTGfJpHudtp6MWuWsQiDTMLS
Kanwt4NgUVwTHnWYHrzGqI0Be7Gu6kdBw1rUAdOaqrcEZp4Hs1NzaZ22djx3n/fvRXk10+KI+Fs6
g6TEADJHVGpi6tFhER1mDPTQ+CKSu8GOs9PqPijL6Ig2QNiT5WIKSuUMXPwqQqBe3gT4h7ZokDRl
tBjzWcsymdlhoUDnzoYK1ECsUcNwmgvqR7tcV5MhFJuskFtp19bEZfGUVADKO4E/C0Tikyj5aOos
h1+VTUjYZBI97dE3NO8rTjmznh/B9jHe1d4PfrDMD7z0EV0Y5Ua3TIbzteT/1eeQKbiypoF+7zlt
SMQxz9oBRsmhoRmt0A0j9yR67jWlUnvxzIuTjCcNz93peZYX3ScdBEdzZGJEUaz2A6eIb3ysUVrO
RANmyuNSxpUzk/ylz9mqjaPRWFtFFO8dHPgGjOzE47e6WWiYEWiwGyGo4m7McHxKu8NxdrbWKbFf
0/SePWvxQBz5089XoM3ztsEmjE/Kg6wfRDHkqPXoKNgNex/Hsm99UijPKiVRmE5bye32M1P1d5RK
NFeunJWtmbrSekmGUWXMtqQBSS6t7jkKRbfre0X/qXwu+ya2CPiAWAtATFyvbZE/LCd5xP/v1q+x
xLvm9ixQpuXSrbsEdo7XGLywSym2DgI7Rm1Lp6KxfuKmce3h14ruwQ0JCulQjMExGbsEjyIwClTQ
kFdJnhCKpQagI8+PryZ71Hdo2zUdy2H5zT3O7kjayE6Lp0AXsmD+6hE564KQdOLioVIn9x4Ejc71
9X2jEM8MwSftQFbrk/am/ccS5cjgddWgbg8kKoKJYm3TDGn1M3zum0tpU3pJbPG1CKOJeh1zVtz6
rloBluzMmfMeL3mW0l2inNi3oXzNfDIe1RL79inNZ1g8yHFysfLPTIIQvqXVkMo0VaAG+vGeZapH
JZTK/8J4co5bjkt9ffO4JzRbKKrHeglBP0iA2MpUEOGvenoFqNyfTUkDtAwZzscPNO7VrbTefJ2p
vFhoQFM8Z/hbOKYetqDfsRp40WU9mlaSdOlFZJIFOmYG8uI5rw4tozDHrYXIWDebyYF07szQxQ9c
lc3w0NO5pEnyYpgmlPTDacrQU2lfJpInb/BWGz/hauU5//wM7sOjiMaglJLR2Cv4CdfTJhp4+ByE
wg0lF+OgtAbxPdgSP3wwgHs51GaYB70DcOKIqKbQjrsQf0G63RITGK/ev5xiz6LK97+TY9AfDjZJ
4ykRM0SHQF9cUplULsGqySUDLsA66u9Cm/gGKUNIs1EoSS3YtZSA1lL85qFQDln8MdYvfdlm4znM
M2jOIOpBxJqCBSJSTXWAwV4y/4eF+E7vw58K9cfI6zb9IuwA9092JGAF7GIjvwnsZRENN1yEapv8
aycCbLIde0I4TvEUD4mZTQeQHDqIyzD/xRFfxXHyOQRCwRaBZXy1F34D/tN0rkSUhH2zF3E+G3M6
bt5pXZQzwVEsIyOZzNAKHZ5dw/aWsieT3ka0bwVdeVwmG793p9P1YPQ93BD3AbG6yWPp32jv254D
+HkjF9LE5UURn/maMv/GsaJ6ze3zTkRq88LO7wMMJeGkXRMdypVUIz/clVO1FtWxcLI6i/xEFn9l
wIEgHBi2WQxf9ennLiabLPAoAJATKl3yfbX7UkeyHFkhqlrGBgUBV21hDjaO8B0UKn9El3qIRS6a
H3/Sp5LmPVmQossRK3ViLu1sxtBIIyYtc/HFKMQHGKq/uy3X8obGpjXvRyCfD2hLSuuYlU+Z7xhV
nYvGbgBF9M3vLFECDVlZyj1h0yZRw3vF39NGLKIXcdm1x2C93vM/gHi+4I+4pGul2MSMJ7KiQUkh
RDgcVWIEtjYylTlHK2Hzm10mZb6gXlFUGMwuyIJeMr0S/jyG2GNEQI2Msfp21ZWTlLHgAt9GWC7x
X5oAbVt+NYuEXywCjmKVrkRXzPOBTQkZqOMntSkTHZZVb0lEc0Y7/SCGg7VDGurUXhf7i13k3ySR
C2/eZ1c8ry/bP9rw9fvcKsameONaMsvB7RdrgI7Vq5RV64D4kYCMSuCD+1xWDlWw6zznxKpWL4Sa
7SHBe79J1lNJHPXd3adYHFu+wPgN9jO64f3SOdJrfMcQLE80fa51vGWrzvupYguxmBL3c5xCiMQn
LNSsnyDaLcga6UIg0nwVuymQc40Bkjxj+BkB0EmxwB1i55UVdaJJUG8lMvdR5+Rw59HUVR9t6hFR
u3qxfJVoyMkZxIR1Eg30MEpgYdq4Az67NAN2M5I9ipZeTE1MWRhLzZ90JZkJcrYaYpGY0U8ZUYE/
3zx/UN9XvimxSpchEcjZbB9RFqi3LvRDdN7GAjfS818vb3D9sw0xa56cokNuv9tTOPjZmZDyigzT
4ubz+jEP6PnHRCDunk+x0Ku/FrrCkWsKKk/9EUVXdfimw/x9cH4jiQdRcjKvj2M6zqEwp4ujhMO3
vgZMG1q1ML/ndUb5yiFH1KkwEB+R+npDLipFywrh6BUhaim5cdlOfYGDMkWIJZpdXegY0iAJFjlY
cNYWQkpNbtSFrNDt2X7/qj+eUGP363Xww7UwZhQnyZ8C6cTPkYLqKPudbMZT8yEag6qIYl70Gs9/
tYYaTj2FMPxNoUL+4RxqDYBd8kJHZqVPNKvjNJPOeY2DI98EOZR3fTjHc5d4h2GYlL3NyZudbFPx
CdZ5ot3/5/QUf8XRfhv+RL04z5qRNcp4WoYuEzsPB3PapSv+eRN/hne9X9H4IlC1SdysHTlhu4dL
2ZBQnkRAHPMksUCiVtW1rC9Po88Id8uhQ1zoUq0A+wvqqqntJcAJxmWwqqekdLaRUvvTXNpzn3GQ
rz0TvbD1jV1JXrx29v08W9wu79ka7NH0up1i+1uekoH2UQkF7qrApjQgDf7kjC2UkmOf4mTvODET
gN8JjgT8hwdxMiOCXGj2ZcOSCupS0909a968tOJxLCL6DrW1ZMyRw50MpK6rl7neFezOC5RMfQvX
K9b7flDwGoqCtW+VTXCu3E30+hcpaAM3MKJaX3Lg8J9Qkf+bex1ExfraWXON4+nWzWn/1dyHaLU1
+tFAuYOZsgmcoyuEYJ/U6fsuI8Yrms+4DvZbTwfJfg+Uyll/VbUkNxiJjoAMWPUZ18dR6kTLcfz6
AfQVsVWTdKS/8LwcbCcunzC00q2VzHG2PlqyfUD7TrtL2lPJRLSO7DnqRMnjnStZ02Y+vAdc7pm1
KWBLQDxMWBAOyAZwWaoa4BY5YHPYwwAnA/NvsdOkKu9Z1zYF1U7hoLtNsY7K/88ZhspjcCRoYeY0
SYcysjWb08U6GWHlMb5u+ekNTMckGwE3kLIjcZGwIg7ubfYoM1O2ySVxR7SgY7wBVYfs8uX12eDe
NkBMnzQqhuWAImWezTkjaJUyJy4A/k2SgKpf2chJ7461AgebHCoycRDaLt6mTqYHqkA47cSC7Evj
xQ/w0I8V2mIrx7R4/mRRGAbHcYIj87gsoj65uz0b9bPQUdrvuwNwXT/vqbn2hzyIMfTCWYOqAayM
syPswuP+OWnJFEkPU6AbQHva029MxzAB+fnX62z8S2PFofEUlgmsuJefebgJqyz5OJgilvbr9AXj
QnkfWFphSn5p+YeywkSRuEswZGrDhQHztw6ARAta8aSrPo1NFEuMFIOmCS0ZMpw7p/dUUhlzHbgI
bsh5joPlrZ4qA4GDP/Jfyz9zw2TWxBO35UbPtab7wuAZhI4C02QY4V4F6InmG55rcQw8ovvxJCCl
9fAcXynsb/j2wTSBytaXBoZRI3SBONyx0fVi0IEF2akBqHu0WPCErwrpEEhSGViMjIvC3Lxo3qKM
k1WkOnCwSYyqMip/xS0h9SyenDlc3FpRd0waZ/Sjqzxr168TI/Smg0kMHPQpilGJsJczpKKUEaVD
f/GsKuT2jaQGx41+SRFji7F3s4pKZluBEDqqe5y7HfXhFlx2KW/h9UeRGPA6iKEUE9U7tH0Qhi0i
lPGgzLWHaedLIwN/7qr1bw30oXdIVwwkrdxSyaJETF0AeozZLpSLwz6brhTtnseo6y/Mt89L9/V4
P/nCo1Zv5UjRO23/pQTzEPKfZ6DVR5S8aSolqAdWgqhF/Uqo5ea9n/9HtmCiUnjMe0TTXMuGWKWv
TbWV9WRB/hoFnRRPetO747cXty1zy3OPd0tcdEc+hhxx25g6aCOMsS+0dkoipK0fpuDBRghFwgna
vu1U9U56Qh1IwfQNfjB6Civ9jh65utyptw52DP05LPiU6hwlGn07Mxo7KdyDbZJK3a6VLZ036JDE
SRicIF6IYynebewQcsplbrRCyCx0DXLFAsa+nCIjMqf0qhGywSu2LfUT/nFbhBPIqAYpbmiRFJGH
QqGn8r23OjCOpv1ilyGT9BZ4Iwu5egYXGZYxpBdccuRoI59orBIjWlPJ4DuFrgWKw7fvApv9kpIF
rWRowDNak4nx5JE5U1/V86PXgkvTZSAc/EJGt6wjRv6+D4h6I6C6IZAet2ZvAQAa1gK7awGKTAOK
BTfqqYsqI8uALNQwE94Hhd5vqjZmE3VIxedcfh4ykzC1jZgmuXb6IS2P7YR/2CgfnQEb198ls+zM
b1jKKozHH6xiMWMz8lZEMdZRXm7lZh3cLoQ6gGOj0RH+2yRLy7PczH1JdJDKzGYrNI3+719+Q5AF
k0zx6wsOVpQpGfSIBKy1q4d1eH8AHhOxjLTrK8N4K5ANoF23AK+0EDB7M6UvoDtn/3quSbZd43vR
1ZdfClRw2N2wR2q2h/YqS9rNrJp1dGlJZ3GPiLD9boo5hEGvXTpzU+6Rsxcn/O3ZqTRG9mfbMCFQ
UAnxoAX+gj8lY9VwlZHQ4IV1Ik1xINXfA3OxHBQlDoIWlIN+U0vndBH7mpB/G/ANpJWLa3Xk3UaQ
56kU4lgxw/r1ftpnGdJQpxnwA9t0DWc6QQ56vsoGQ0KX45ABrwbTG+R/c7fKMaCSgw90bRHodV/u
QgPINyv14NUENkj/RCfb9UX1jAwE4WLX7y3ZYGg26/7ltqWz5XJwX5Lnj/3KsSo7ml/nZcUDB3Qy
cLiOBv5H2HT6lnpOOKlG/h9FRdBntrFJ5F1ppxOJs28cRksPxJWAGoJg3d5MERTE/jDjqZYq5cfp
Pt/5tameDu951JcFLEko6fJs/k72PcgEesbIBKAkA+OHVw8TQ5LI+ME4tX8FFBx2WH0NUvbYXERS
tSot6fvUQpH6jP995NTk7OOuSg0+fHLJ1JS74ShQnrqU6boB7Sfk56T5E/a3MCf/wHMYJWeOxdgX
84mi+vFpoLIWBEytBpXQYkQJrFfkIrJ5f8Ys68YBDVQ6/2emhuNSdfm+WXbo9HEmFIpugRiN5tG9
bLvQZCF5H2iQbxtn4c8PGdmHvSwIvmXDssWL1iUJiqdy1FIkdUP18STEY2MZbI1dP02quzFEALfy
n7gE19TpYJgPLcOB6ImzWpI1n3XyOxChlACjzGZX2qCmjhMNjp0R/OX6utYoV+bduyRVYhA50AVp
qpnjX0WLPTNKmo5VDZ+2esIBTUKYlEUUnj/9Wqz8HaE6hCgS/NyrORVNJ8tiWfGc3yi6ifcdMn3P
1cJMPVWgFL888D/gQtL+tlDkXgR2KK5qmOFuUpiSRqoUZ9HQ2aMbFaWL/w4sWtG0rMhprrosUY6A
zNC8y7jU8dFsLt75SfkC5Ms3gL2bqeXMdv47dgcWTCKtNnPMpiqRzda7fQ6FM1tqrXIrCh+HfET9
KGXJiW6NntSSBx3P0jJGqqEhQnuwajNSmI4vNovJbGrW56lw7kqZQr080EDn5pny827EJF2Z/oFE
ahy5yjZKfL3vTzY77idcXdVMKI3BG4rDW/LCLSDh+2Fxm6sdOh3Pu2yJuo5rEKRmqzSVbQBTF5q5
CV7w8a4IDEDLDOYuXQMudOmYYWY01UKGT7o7/jOW9YzlCV0MUVKmKtRxFk/yjPIVSPfe4+9/BfrO
34lBqYxhryVZ9ZlWWEpPEedZlPo2uxB8R+ubQV5Yaz5TG/U4R++YdAqaPU+p35sRmkPnGYei4AAA
L8mrWTTCNLLvpgp/EDM/NHxBggZcr9OniJx4JWm4lQwAe+GVaKrvT2TWB+oyS/l3uARLABYehhvh
T4FEh7/4mpns/6Ju8Mao+6+cUdW9Kkic6HsjvB5imbHJfZF4DGDY80cTRVsmwSHeXkQ2ODpoCw4Y
zDCyVoImU7kITKrYUzt3pRJt7QdJ9ONvhRgJ0UPEYHLdlPwIs95VxBs8yyWwGG5MKiJLysSn2yeK
jw31ozUuRQFB86jvP0FP72cF2PL3eQoI6PkGA014BRpxY57WjNiNuf0sO8Ec0BYHtagVEH/hj5tb
0X0PivCFHdkqA435lihnRyA7bR4qgTOpSBZe/9/k8Uj/G9dD3zgcHHoFFw==
`protect end_protected
