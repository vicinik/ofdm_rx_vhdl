-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SZJkonfK6lW/gt5dvDTJJIGn/6um2xqEZBCs1QAdNSAV2NOl6Tbr+jKyIIG8Mu83LMiP809VGSb+
iW3WEGJzKEP99W4FYtsfYU8aSPLv7g5OS4d8kKO03WDhwY0Dw6Y36Oix3eaWFCtzBsz3mGq3mP9g
QvTNHD85t6AtqXdpBozqBlow846/UjR/O6SJOLK+8ojf7BPgKOphVtvsJsoG3TYDoHhOCjCke4ny
pCi1Zc+q0z5f5KSPp9G55tfkzzTYOHqq/RTl3vljCioGDEyNK91CllDLA4oK0ZqXLaLE4uhKFClb
no1zO30HSg7yJRXy0ehNF+Gp9/t+IkacHkhxJQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 194096)
`protect data_block
+kDfkvzAgT2WJNhtn9Qr8cM84GjJC4VPZ9+2PT946/0+Ob+q9b0HDMYSVWGAc7vJHpFVs1vqmIv7
bPOPZlgzWCT5wwxkNsEl/xvldcjT5b8a6Lhj/9KiVU4fW4DhgsZb0jL7TEo0QdY4b/D1foLwR00k
A+yXNkxnzYxGIZGzTm7a137PqhZ0CWhdmoOlZ6Myyy0CGy095m2jocUB/LvrzWY7HrK9NP4qz+pV
ATxm8HQfwUZDFYiOWNNPW2G6NQz3+FxlxG6YKeRHqdyS61+5MQ3gR8eqy3w4pgE5hkGG8eDRf/UZ
hNBo1kf78COewMSCAekU1sARlB3BeP0BAkwoa3XdnYln8PEJC1maoqB1iNiimPFktMWZj+/Mx4lZ
xegurbjR79QPJya0KPMf42e6PL8rEPDutfmUPPDeKZxypA+Z/FAfjTQzzds8u8kAzkdsg8mbtXNC
iQlSV0rufHRusmAkBt+dLmNozG4/OoTbF3mPKZQw8eOWCEQlx30o+RDGNPpJmZ0g+gtwfSukKzpx
WRXdVqKnjLUxezZZblVRrElAvO5SFrR/1Ofqe6N52AmOQ5NpeO7yALnIQXoRxsdPcIxALjlGa+rq
qQ51stZ5Xv0p2vgCO7Pna2Hx0JVGnLgrMcFsrz/+i4G8A0UlQ9z8a4hOBPLi8Yp805UCD63stcWp
yUX8LBUO4nUlxHmrbIpuNrMMrdguy/Fg3w3wAVsFXP6XpfhNqOfcntSlC7zLOvmXKOccS0UWClMr
ufs5Jdi6hIUXcZAV9WeELfuOZQXQDeeMjR8THbLRYFUcwfEHYEAiY1LF2eO7rm1cWh+OuXm328Tq
V9Pt+XEF9bpihER4dNlB+x4qEjKgypYCtuT7eR9iX6k0behgy/jv8BeGFeav1gOLbNtJrW9PDHrO
8QCYC3ciiki3h/IZsH7BwJF+w8C4AR/fe08TmFz4G1nudABptXITgpBj+sh3rvwXdg7v0z1lMe6p
gYOXolX0LxuJDZ4lsHOB1YRGfhi36NqLDNNstV+XXW+Aum9Bv1t3ECG9UyteyqKmMvar43dgaduj
Juz3w+Lf4ww+d2O+uOs5FthMJ8l94fqaoHN+6WtYkZGgTQVZuT0Co6da89fdaboercRCasLeHAt/
hwBsG3L/NW9wJPO/UPT8Vc9KIjwBPl/VbwRe9dchaScd63zGZ2VK0K6KSR+LRoBp+qBP5cEN/cZj
jJWVnMC4yoycL3awa/6IIt0loQMqm1MQ3iJEEofi7C3mNAaEz8iue0dyZ40H7WEXGFWn5JCnUEfT
xAdBJnKc9///6Aecx09H82ZZPE0Pi2OQfJHWcnvtTygEKfeHK36s7CZoDQipMdfelEHw4InSMjML
SoNvqShmGoPCuCJvrrfB5f7B4PQWlAUkYIC+ZsjbxEnonv6eKTual81/PPcfOnAvvDT29o+MZpyZ
rfTHn7NYzjxPpOw5D1hZxQK/upMDKV5pxQEJDYRsRoITNXKVyjP/JZ/xy9wUHx+tnW1u2T1AeKZx
xc6u/EnTv9Kvglhc75INF/H/pmMi8wdgF7QlXYtq7s+szFP0QPUdpiii24vKdXI0kWDcmHg6U+4j
OvxSIWr1+CUbO0l5/thgqJnEVuQ3TzTNemxoU1SOJ0LOV3efaGcR20ofqqsnHaMzgZgeFkAeynfz
bAR1oo1sNVUzmqmH7VlzYCcRAFqSlVvVlBhljs6o7+l3Xnr38w71ZHs//E2Kt+dGtS7+Vk0R7rEu
Fxb4ut5oKCseSEox2hbv1Fc5aYrgmkJjXJ7dmrtwjXH+M1IO4KFf52LEclhZBZ+FtyMn+/EofZs6
scNI6CGTxKhuqidlMLQ/4QMWQNh1IJmRXAiZncgTeq4aY2ijbGIdzYgTOpvn4OKQootCwscfhgju
KuUGLQJiw7iUp8v/Id6gbp4CMUYOlxkxlA31/h1s51nHrIv5kDfjkZxj2baOmxVKJvMfn9q+I2ol
xQHM3JtmiixqtMbBVomx0f2X3Mr5agUltytxW98ayfj3i0UBoN+eWRyC36gId3CA5GBUi+bZE1kg
cklap4qt+yzbjHUjPTEtU90OkVmiIy8aHFq08EMbov1YT/rYUUDGgidF0OIfNxKSqGUAejehmPaJ
GRv6EHsKkQeSzXsZ/sAhgQXKYwcGOh+n+OMO5xEZAVD2kljBJKtcW1quOX8U0aJJ1esGxoFcSUJU
m9wcEGGZIFCMQHK59AtJ2Fm+JJps31xtxjhRii4ZswwVWlAFtN3vTTfOIf2oKZE/mzHWP25HQWBj
31lbjoymhE1nZoY+AI1RpaxLJU+3xNsitFoz+nJa9Bf0eEYHPYdGX9MSgcDHXdp6AUokmgalCom9
dG4Gyv4ZX7AbDKz0LJt57BOI39QkwHblHHKLiVt7deljJAdvaQYbXEtHRe/XYAkZrsuGbN2SNfTE
DaWMImTl4nmBkxXwDX5AtDWulzKzOxFlxe0eJakSHOPtjrL1vtdhZRfCRa14JP+vw4mMOql89enZ
LLVwx/EXnz023twaXQZ6NhmqXZEHP+OyFgogTIExTeEPxKZE/XpBS6/Oc31ujtpP5z0QzwMXh9w7
6yqQ4i46x4BHt8+FE40iLyxSqT3wPYCkaCPO2gZU0H0hFvu+t3US2GGfeRDZDebpobIcBM8r7FHK
MY7psm6HJeDT61YjR7b5ui5+j7hluvd+bD5E0YBHVPTNkGior899EHm8w8xhDXHevbFPuuUjCSl/
gPWHIF+GOJqswlAS762JbuVM+Rw/VNru8154L0XLh6lqH0NOJaNn7yhr12+2UC8w+3llODsCe1hI
6Bi/S7Zctp6JTrb/NsQAIFeUpLPhgVhDBDMxI0iTUuZp+XgH5K88uPQOF7W8f0rK1QtcPC91LzdI
1fx6rsBSYt2Sfo4eAgWrDqhuKSA92yb6vvXFXILa8wxrjC5mqZPmWXjevEUH0zXJuXgg3bqm2HJR
ZkBw6NRTAm5OdEs1OUJwQmIHJHEHcueBBwhz1aE8dpBloW62meJ2h676omjgl0xSoaea+b/Z2eGX
Yg8Mxun0cv8cy7+zWeryPpPidu2E7v9dC4XokK2dphKjSO2eyFd+oTKrM0n98b1+2t7aDaZV5i2t
+W4FL5nRmmwYsyDjbqctF/pL3iTb3JoSKVwgaHX4mnE8bReq8UeES81Z+kBjz8L68K/ASB12K7Jg
0h4+x2VITW7hNDMrjp6HbYyQB0/se+hw71co+ZyXQvGU2cz7weSZ/xuNRui4MLTRWLM49Wvo9dPh
yoJEcDcscejV1GrxllAy8bX9uF6ib40k5Dyr7tNryJ+8tYwrzd1DD06ZO+IH95C/bfvQhcaHY1RG
qaf9kwtRnAKgw7IEeGCCscCtCbLZE+4xdDjLibXiZs5629TuAV6stA23O8syAk+KSERK5ox3Zys8
eb3YAkpoZKZij8JGBoakUQt+cDbHnYtD2yf6pz1UOkw0tAFB25eOqpp2KZ3gUIvRJIV82gDasNic
LL+psGSlUIzSQhgnylPYnlFSecfIRc8trvaUbhoF82RiwHWX0EUA/F3UrFMU3r/FmVDMggUuIyRo
tTRMmT24Vn3q0KxQBCR5Wqhv6rGg3/zjoBlP7CNdCVUH7eRAHsp8uMwwIaR1IFts5RzdsUgGxHW2
FRLA95OHf5gEQbbcfdTFzUbysNuQYQqxn0rQu/xx93s9Hs6J0T/pX5YGs28bvfxxeVsfT3EPJVWh
lqH9iT8rk2WGBS+TLz5WQ2y/wywvjIQGqpO6spZpzJIYsYswnpdRB2NMolb2vAZFamag1YxGVkYj
neqZzbyYePOcj/JfWdZ4kaGS0tkAxKW58ooJUWUJ96kSjVnNiQnkSj3zrBlYGKrAtkezAt/eWBgF
5Hw4clJ2HjJ59+h0fmqeZBqlxBjgoq6p0VNxIGeumn6MzpegPbRapVL9OdQbldPi/NdEc2AGj/aD
uhqGuPeHiwcFktmudzy72eLu4Bp73/yHRgoLkRX0uE+stEWQh+tV2Ec3M1/X+bwUDwmjdofUA8zI
adgD6CbekRYosBSmwSXhJ/0WKhkuytz9QQCI6taeLWiTDjmiHTWrLWwGCFejn3CIXCS0eYBdYPAn
znCmRXjFBulJXoBOrd+NNNXx9oIgRDKzDhrcFmQJVgAQhAli/1sJiJ7cyqO0ocJuE9adzDysH+vQ
Prbb/I32QGljMaW05ZJVEdDS05VnawKEBmCGA7EM05m4wCDMcm/4JrrIdIuMavwi0r6ORBPaJOSB
imH3q+9y9xnKfICGtXkW0UhtkTv7CjOitG5TNoYHgYpfVJRidhMMYNQ8KtudhlluKDuddeg9pSuE
tI32XuQ2h7PIx0KrylWW43hJZ671MCP1SKKYmwqlU/mHvFi2bxJTsRlOhFnaVU52uuUHUVxgmwXz
7E1XcsW7lzajq51genU7F5P+/8dFn+9ISeEFeRf5Jse39hsXUdMMCEGXK0vQqUBZDO8H0yG04l/n
KdnjG20B7P5KtW+ZWG5yy2Ig4ifMbOtc9Rp4ODdsxc5ToCiT2fnzbozGRLftiPH/7LY507Nn5Fos
+nfUQuXRW3pAz3dWwIQ4hg8+awW8E+3cT4hLB+rq94XCDiCT9mEyT2cHeQvAYMDxBdZKFWeSNf/b
jE6cUIuuZFCCtn/I+pFDjAu/r2kwKExjwOj0R/5OJM+TkAwWSQ8Ku6vZ+9PQF+1CPM6a4wFQ80Vp
TuRxigxJdtGMZij/6dUwnz9jXTc3SiGtpT/T8P0GeZaKeBDytJSdkwFxup5yzcV/C1vDMUjRUvwi
zrpEKQ0Niofbqc7o+nUCE0sHYR4GKtmBI98vh3/wOG9VxZ6sequ/1BHxq8gNUnbnlRmcwB29gmwX
Rp8ZW9i0odh10sMVdizg9zUAiA7WmZP6HJrc9Emq8GkGawqdurs4ALp58A6sPW/f+xw4G+z5zFuJ
lzyrRaTRZZHHS+LvFT34qHxJ9zl1FCXnHe2+c5h15EJfIjs+ddMDb/43cJjWJ/ziRD+bvSPS0ivv
rkjBRPiv/6DAACurrBzX8PhZyir7c92hldS8XW9uNmDZa8xwdxtJTmwndngYJjp546ESYmXpC7+S
WmYiwbyq6EEq1vddCEct/RCkChighek7TaRkR7ElqcwAqKw55uYo6wuKcnmYiJezI8Vfnk1T5F5c
bQuqkmPnESt9FUqCd3SAR+hXSsLNT0KUBCD8oxXe0MzKsI9GlbpHMaSbcZbut+WHK8nnoblo+VkX
Ks6lpztGPEIw/fMEa4YAJ4t8IZ7FBl8rpJ7OIK8ISYnEA4puPYjY6xPsqIwL13owUF2T1ccRipTT
ZEgTnUyiNQ/rawYPetNxrdom8f1sHOqn/Zjj8Ej0dGlw6oS4mqewM+9saRRhJndz90ovVmmPkdwT
ECcOI8OjHk+rXjfGCgi9NpVVfw5JwuxLVG65zrRLjuZ1nJGKFkCmY5vybdyiITe5hChzq08LoJXL
oA0CYnO7co6R5zvVc3221kTaSXdUs2Otcehh4T4yajcvmibTxmAnM4p5pp2fDJcdA4lgnLtMsq9H
Ls5BKuhqts7AWv/R+LUjOqaqlRevRnUUtkj1ialm2PnFzlbc1Mg5vE5ERdmzPefoAC1ufnt2TT6R
Vyf6ftNYjvqNite5l3RGTsret7RKdpd1wo6ogN60XzC/pDesBUDbx1fQ18EfNRyx0DBdPvDSLu1K
lKQ2v3GBeveEkWzMCVm0xhaIw5fQLEs8IHfi38hwc8l5qeQwnwsThKBRD1vK4lCudBsG5Zig/3zV
tHJepA+dwchu4QfxZatiq3yGIRIJ3MFiU2y9AGZGjkkKKLturBRwzH4U2g41Y3OfIz2s/C3F8my+
9cIWgHUfDYr9Lw18Wj4tJ/MCx4vd4DlYJifkrYvtivNRRqMveh0wy51Jch8IW8PrHPumh+pyUNAy
vTvhd8u4XM+PDbKhUQlyQB7Gl8HkQgq7EevmwqLwUDZX4idholjWvPoRI8VZtQevhLkEU2pvg+fy
k/wgTEXayXAAkfphSe2XVSwin1P6zLpbdcKEBdA2wp/SfKUP3zAFJOrH8eRb0MtjZTJmXA/KaT9S
ccZ+98pKfBUkyQhlTWN6xRkjpUczhOLoRPA96Cr5ig7IFMlQw7fafdZVLpdMeWj2HtFhRmAz2WKj
Kv3sNhVAXyqfzQ5hT9rrt7yCuydK2yJmY+kkMuWKiLzaumuN4R9GrfhVnmz1wJvQKelFzYnEOzBS
hLvyKWMc6B1P0BcV0C1x0X4bIQ5JZHD3sjoZG1FczUYo3nRPyAm+UhsZxa0YUg0TuQL+f5o7gaGa
GFbX+dnvUYgj/Lr857B0YlODZXo2kWWbhPRkNnGWheSQ7t4Gj9P+K3O/NpYHF5JQJbHjQ5GXeQsB
pTglHz+/B/3wla3qcDMWGJzHnf8fzFh4nlRjl0XHnUKWiMkTe9FWYyg4cYLc1LxGEJhWCYsNsgRQ
M0qxyb9qZ2aCswdSfT9CJF6D+H3TxxCSW6ExF55rQ77bp4+IhXmTUPpyWNIuFpan3V0qt4Rc6L86
QGOBpuV5sXyaAMB3Q1TWnFN6xn6CYtDf2HRHtz/gTS35D/J2QXVEQE7biy//omIkPemJ1HjpjD1X
iJEYykCGhu7KKOIF0YhCTAfi5UKPf2C68SJ5yR4SmCjXs69WQsYgAkkr4CoPMn4OkdwPV+4Qw2gH
wBg6uu8I652K6m0gsU/sEz4vITGb8hW3/mIFY6gSLUpPsv/Lu8AinR3C3byL4mNcDLProDcrlKne
+yX8Q2nlxiwzZugLjtgXTmz9tAWcKJ5BhQlWwSBR3fTNTNXVfsKPOFcBgUePcWy1lXIMBGM4TaGA
U0lixzu9prcfTMjC3DzZwHnQauFPz+n2BIzFrSuXHv0RAr3os0tMO6QTbvGBg2lRXPmVT3vag/ga
SvpvbU+84G6ENgTUXLjWTN6K0JQtF/PF2K8983SXNvbLMj3t0xtSuNlhSIln8jCSgC7zP7Bc6In8
NC7tlQYtReZsO0xWLzu3kUQV76EKcDDFnt9qgYlag5GhmJK+o9kd5fKB9lJXhPWMwVqMswMH7Niu
yk30gQ4ENr9rszSmFh146uZ+WKiNsnusnbP8/Pz2HINJyTkCJyyfpAqdCI6r06G12+8jFH6nHK4p
Sfjcl1K8eNDVMB6HfXql6/dFdrQDE68Z1EnT3GN4bWptLnn5l5zj0u0gSXPqklmNQYTCQxsY/CLx
GC9Zuo2iySO7ECQgv/oyTARxA/AYFX+fsSg7D9dPhH8AGYd8UJHe7cFzwHi7QGieerth1Z2Z5vfb
t8VPNLJxlRKBCWKt/nYTW2V9L7c1Qd53Tp+mlJAL3v8uo8MTyRSRptbEWdXSL8FmAUWSiIbo+t4R
ssQTHnCh/XEcsMAlyQ8sD3MIIUjUXbnSTS/MRs70ysj8ck/XAbeNvvfZBYRHWcf2bm2qbK3i6wcm
wVuegYJkQOIPiFu9nnDXd5OIW9aIP+0bA+O4WqYjMLX6T9xvOh6Xfbw/a2zaTkkeHefSSVFJsTD7
n5tLCCAm/4VzcQ5ziitR//UQcfucyuf2v4j/H4zogHtv45FXc+PPxsY3Cvj+ruDByzQX0YbLw/io
dvBnWqcvCdsMebazMsm0tr3tiwg0lwE3MP414McroY/Bw/BGn1aJ/5bkab2RsnxOURRabvMWEamc
5AvHJdXeYUhTSKvm4+8exbtG+TJbFGabu5FUI3utRxI/aA8KD1kCgTnOGOCiwro1ETefoTBYC1G5
hLYW7Azm8pC5xoiKx34RNS2VoRLGe+gUZPcbB2YePEF9mHMUuMq/UV9J9v144v8Piw9vYQeNLxNc
vmgOgK0T7pIRCV0VwU6XbzGF+9znNxoEGWpGxCNcnzNSkVFZCnUQkt0b10hrEAVIySx0Jf3EY81G
XQiSdieuVVray10P6fXG/xs1tKmnSn1v2JrsiBcYOYxtpbROmcd8UHcv5iG7EAiRYRd2CZJP52M8
2BdBmrdhTkHRQMHKhTz9zqaREb3Ls3XC/aTEPSmIGnDMx9W7B8FN2xgMWRSx+N+ftd34qxaWyC99
9NYat5fHNSBUKIuo9moJMUFZFea2Fc323hOgkZBhqQ9nt6B61o+E+fOHa782ZTdag3PXzqAbARLO
9+KbSYyhNmJ3wpXALHRC21KHY9nyDhWT17e9lQQXOMOlDe2XUeXFcGFe4SpoXKh1kAMs2CwFJIGv
ZA30xgvMh1tI7fKr4BD6/X2eOaj5N/8Bxwj0xH4T8rm9+3VBlT1VfPwnpANFXUQ1RkC6ckA5lpIh
84ChMALc0E6Bvi8cvY9awkvwOViLGF/5NeZoDR8zV2ytTzvd5xrxeEdH+Pkvxku6r8O3+Uxsf4n+
g04dhFihC4Y25ffb0Udo94HaWaq5ZeVM24rGNYWjNjpjYLDlKFjOy962obHa06tkA7m+fcCVEC9w
zAe3Gk+oY4yzGPdHvHlIBFSChuA2OEcwtcNXVhiy+raOPtq4aFZrYWkpied0V5Uhlie+B/MuxiMt
DEQS0J3jniuSB+DVO1rCEeorDQcVldBZ1wnUYjnQvnUGUVxO0cidmyIkBZ79qqXRNLKgWnRYCKg4
7f1WIc5E5njHLMRMB/kGzp9tkzSg/4mEzI4bLnl1R4/SntLDOg36WsGGlXvUEx4yiMe7IbmTYtt4
iwhsMsHsLKU+nCVVtWycHo0ozZmsxw51kMwG1Kb9WJWF9lgN+jrTBhVrq2qr5cpDxPW+cmLWJLtI
bKLcxGCN1B1kKdM5IFHBqljjlimmwnrt4lesA/4KlC5hvDuwZAZqG00l9Tja3hpXtV7tGQA32pKq
DV8b0U7odqIQMfZuCV5ypP+NbvUFTEAEohCF68tMklIwVh3WWFKxGJNOAYoW7qBALu+LWULFrSai
j9jK8UKjoWLMlK4ftvD7cpnHO5Fi8eBiFjx/8SWk48mZq3h23GJl8CKOebyZ+6K3eIit68Nejpef
quZBiZwBoYuniv6fpgjeLKLQs/dvvvlYgSeLLxLZU0kIUf9Vr5EKVSWruWRctjOV4p3ipoK9IA/Y
vonJBO5UcMu/yaog8X+GUHKAEX6rbGm6xvQOuqFalwUgZwZlO3OeHmSl8u9MVHpUG0BewbU8kpwV
UDJY+U4IYpmkbB+g3cHrNn+lTTPB21vChENhPjf51bjHoolhNfepUaGq2XZEadSb4sGNojJ4Ha2S
rvSm/dHi0iMkmJY2uQ5D2fo7aMXBGEFKVtw3Eyg8AP0axwHTxZB/Bkri2GqfDzDZEeHPqJUK+SuC
VS0FIHKaIg33NK2fe7GfO0y6brDb3saaT62hFMW2+TT3IATxqoxSbjfkdZTIbCtZER8PTtMLzEYK
dy45fsMpzfsNKg6mdI4Sp3/LQfeDvPlCYxRqxlNuNawqzoxWp2fprQBKSDtsVBB1H5pkr0+ycmOn
WAvy9PQ469trLXwRDR9GRwm0SLSpJDG/Q43/z15hJHhZLbUqlx1vuMJ9d/xFCylxpZAhnVawHI4F
IfveYTq9UIc/nOTs9yEH7U5ru3Y4kmvMd1iI0yItBq9/hjDoINfhdow3cGOeIWYGBndcgNx4PiHY
N/3eh1C/KI6fRucscGoe8e8BkDjA6TPWJdS5QXID0+W/xwGzdf1LaDGtf58gBe1aSXrWXnStercu
jbdfodywkhCMJ2VMzSigVljF//CnqqY+cRMhyNxZffiqpdAdb8JRBsYNGbSYqUotjCFaFF4aTO7g
Y/u4WQvlx9BFWsMGww/YXQsJuhswT2rs+P1WDLpjAaPVJxvxkjQePZs+uyCTV91FOC83vFqLfWwo
9FVetG2A2WF4HlYW29CaQxCRaDvuYRvfgayE5+S/+UWehV4AqbBfHxzBf2GzhDAcekGyLu+aD1H1
Iz7bUVQeRjbKvi14DkTX+87U3WyzV8AzFOHNI7QlMuZUyh8niYNPY7IYuBYbLdCA5x/fPc4uAEjO
VT+D5lyu3RIpRZUw/ptqCQzYZhTxOjpEzOyGSWagtmZ8Z05uydj25wG3lo/ja5VqQJJ2+KClj1r8
/kpb8V7prIA1JJovgAG6seQMqAFMZKb7P7ANRAOKAcriDTLoZU89SBiZ90GUIjVpKDuqSrYUDFyk
pwYtmlghs8Fm+3dBE9WTBLHiPG3/1x0v9yvUdqRzNgdilCmnt1R1/EzrVlXKgdgEZgnLU1pAOtrM
5eOBdmSIOi3xfQCNwZ5o20akWxzZVq+dL1xJzrPKdBHmnL3kdPkvfbElG12P7xErA6oeixeHSJis
T2oZFp9LXrQty/rz1/gYLctVyFUF6YFuisXvnTGm7POCtJWQvaKv6PChYeV7AHMU6W3L2K6KtckX
fOSJQghig9qN0IwsHdP5jWS7NdTgSg1lgQCmvmibP+nbgPMacSr3hWWD4seOiOZBrJ7hoypR5Vmm
kg10U2B0gQzkEYLj/1uffy3XXC5zLB0PfuwMHBPuLFFhh/I/TIk6iLUyHiFdY4fY764gflMDPAJY
SxA0mwp2SYaWGZPkIv0iXqEmQ+BgA8CwL1PX9Am5U8JVIPCUBY37vd5oiUA69RqNuRQNuTUg54Tw
HlWD4r71MS/F7GOZV7kNItENwHI/zO3xxUjdgsgyuFCyd41K0NJJjx4UZ8kZiAWTrLSHe3do6Ed8
xedR3/4+G4rxKB6GBmJwTk6wcPjd5uhbE1ozqF8PEICmyayi0SXiiRd8rjqSHpOwF6DfICRjGzHp
biUICDuMrHah7ELUQhAVjgY59BMQhkXv0kMPdOHb31vRVU14vAgR0ViNRSLeMkEL2HKTBgAbLEbK
dF8mWIMRrsGU8c7ZB5UG7MllV5VfwSf/hrjHkT+xzfC/Iz92d5MZXM+DORjJwxjfvcsMaaaqst1Q
aQqMu8KMcTTIGeWz+Hic9kU1pWYc0I5v9+Xo7NQyY5/0uh0r+MslRaDb9+OvLLOJWG2vMa9F10ur
DU3+uwIzoHWjDXVZPpEhWZhaFy3cc5JiQX5F0+2VM+zi1C/RUXKHQrubz7jy347FOG+JGdQGcucu
7oKnnGiESMdrbaJn/273G090wgcSgpj744GdL8pgb81aPl1yQFluXf2/VotSVpHtsjOmB/EnvZJ3
1tVahIclsONLSrwDOdvF4xvcEEiyvXglgD8xCodkO6WfOIuTE4qvJSpL1SW+4ksvF+8prTBULEpj
CPdrzaNzXoNPYn5vAwRxS3Hr4AZ1tREW9AztvDpHYOy5VlM/mspzIc56NWrTNNu5CXRKyCkF3Ccv
kmGxF4R99qQLfuprLrEFdXTeT6ptnmtFBCRchCzoYQgZjIXdpinjc4WFrww+wKr8+8pfKVZcgrM/
xfE+BIxVk3A2LKLafCQPrRhQtONkd+8PwoveFqJWCCgHWAgNfQQViFb0K1AS7tk9nA77V6QJ2x2B
Aa0l2FBNHeQmNATB+hr7KTnYRyPkw2QIv+eB/6aAShnHhwJx8+rO6wNu/KAJGbE6lovupHrZzuRM
rYpXg0OxDOy16/RrGvjdDITI0wCrT475OGhUlkLLFwa9waGkzuHBX4F4P/1iaJ7pjuWgmZ8sxRfk
TmUROeUnlg2FMIrkxqMAq50StWuXNChhLYyP+AtOFv7crHeqUWF9R1jloYUpHAFX05VGBIw1d9G1
narMZp0I5EKbhZxEXsO4wtRxOALPZ/D+XpRf6HNMAamwId2i5FMtnBcVqnkdLx0PT/pjbljaBd7H
SkL67iLl5+4msecW3S53bMJQkpSKUflcI6vnnxgD14JN0uR3AYznQUT9sG/IVyRAoRjz2il2NN/B
hNX5g2gqPCFJhg1FqIr5Y1MFaJr3wegecX+QfJj4FlGqISqkvd0r8azPIPDJ9/0i8aeATz1q9A24
T9STZ/H9pGyq8cZPrPQebbKbEfkkMReHym6tW+dES0yx7XDwn+CFY2RZQKob4s/3Pd5xabXGmQ12
JMiIwpJayE3tZM33LTa2+A1zgp5pslmi6SEC6zmIftG0/Frrzg9Q88k/Us970yRxa8ZYnKP1Kx1n
Mz5OSfCGvoQ3YFQwWXMKvBsEF0PQRjZ/+gvVOzZMmhOVVzmDbsqePL9D+8oACmePMw3ra+YKWgs8
1rlBlgP0y++rFS3IvSvzXjLKL22Uux3qnCksU+y9PMBf7sTK7Vgk9/kKk99zeDy5HBQZhLS0JNv9
JriLo3JUvQNIng58J5eidLp9Fk4RWkiLzV6oYqBeCYSNn5xSDoIGyUPstD0t4SOzIQRhWUSa2Q7N
+ZiHvVLWw4/zwmGI7gwF+9/ud0YtKE63xPiaxmmjYQNwA2H89vhYqx8M6mum3vAosLPh8hA0DmCW
h1C4VRfMn6wxwCjb48kxl31PpUrRguQQwujJGLakVtParTDMyHOkspzMWrklOmnHlrrVYKADC/56
0bxi1xbVKKfOg+ItHf9Lxn3Lw2+q65BnyQnhZyadahV0EiiuJbRHZVD5e2vDcKK6jto1j8dCsLtr
3YZ4LLHy4U0F2bKYD4t9dFayPbHsuTt/A+20EQBePuAPSPpIgteYcXargo19cvsPxvNEe+oTV/j0
dsWXMO+PCKgf6XCeWPkD8QjajMf14CFMxjKCaYsIPMAoo3nSxxjDQBFih47w0SzsVZg77fyOiZss
4H9ZnnOAFFdGi6T+JGB5gOEsM48a5OIGhJ2RFPkXlHDq968T+4MZHJS/JghRAzNIBUDxS7NaxzST
RRPubJ/Gz4R7HZ+rttZDjBIH6Gcrkx/bX7dX+54iytYKnd1cjoq3wzOn4+ou9oQon5wAGx9FRVyj
UjvWyA3Nzitj0bh7/XvwtmtSJDmBXRQtxz7+Hk/3PZU912QA9V2WvLZwsAvLy8y9Rei5Rk89R9ZE
cfTf2WXEz+bZBMhKEblZo2X2l57j8Qlu4wEUkb2ou6h3N8u9FloWLEK8ocXcjzSjnZM+bXlGHDIj
20PlJTa6m63kHDBhCTKRZUSfW0X65ovdRbFWj9yVw4CTjVHvlxOZ7CAgoD85t8z6ms8cW5OPhO7c
1aSLtOkft2o/KzA54w3Cuvv/UhDYuHeEgFMbbwYUt64gPRbJEM+LBs9EUQ7Hj6W62RjOMMwGwoTI
0IUHvXBDrS79zkKwj3LZQCWW5Ue3HOlpw8CNj9JkVAGOdqvDqwamuioy8jyNyXSof/UChNSX0SGo
BhYw5QWzxrPNUhqq0mQ9kJzaaaGjC3l6eqO6cE8FCU5QPAp7VEptw+b4eFm3m0GMW8Cwh1Zu5p5O
NMgjC+liDD3vE5EVq9n02xZTeEwplHU3s3ctg66ZzkEpmhdlXaD9zXgNtqLFDyZgL31wCkLtiiKt
AF5qPlEEfEL6aG7ODiAYW6KsgJiccUH+LtJfjmbf/ogOCC2KQyXoy8nxKLPpvfNSsbYF+Gl0h92O
z2wUkpxT9hTtRxth4S7ZwNPnq0bZiNgiHsrXNL+YJuWP4OBjImQgmNepyfHgWcTbupT2fhE/k7tU
7XQNDjmBw5PfT4XN5K+YkUjcZLEKI2JCKemghv7KqRak7q4QvZ4SMcik19JY44+nQat1WjVFqBqr
LT/BX7N1Bs4XcyUTtvr8v9tJOcLcnrnSmMTEv1itsv8x8/KCk48so/8XHSEISdVeMBt1jZ6mhX1p
hBHxv3gXwLLUQDJzumuNZHdZUGHwvCx9pPBhhHho8JGL1Rd04lOGWX0mJ2/EriJ8h6J1qcGaG8CN
8+z2/hVGclhJuKWHtGVtEFgCnuvPoKVZ6GUyU2d3N+TDUg11QGEl6VxtG3iTVVI6cbo8IjvfKy+L
0eMLtV7dZgnGxx9XzDgazN4bbKmoMJuGj5lte1ybdgKIXZG25Hr14qIdoVJbYzGaf618pkzRT9kK
CO9EIBJGNQAcLKigyZ9RgyFDv3t9PVk09Stz6ET4Ksow7zAwQRAVvfo8NAm6eqaiIBsNeP4iM0IP
JdYzAHWHP4oKPDa1CWtmczGxJoAQdwaHyxpANQYvGOU24aTlAnvgrus6qquLWityjcuQAI5XxUkR
XViMOL6n9i8BgUjaWhAETYgvRAMMGkQ8IkH3zmFpr1V9JTcuaC/Fs2Vwcg/AEpT0P1ms81qiqwLz
5SeW50Ykl4DnueOGX3wwmGmqgne5X2QSK2iw70aABtM9/WVUXeGBvT/Yv4p3vo0EQ4zDACmuthlZ
HzuWiybb9gAV4g+SoN2DBXxOQ2bqMex/SWZ204kx7YbciZ8e4vIDAaYmgjyo0i6+TiYGwavQB5LO
UMSK0K/ucIgwky+9tU7IGcvmc1snq56qtAWW1X940lN/BF0Luh+hnfCq3E4mr5H6H65Rlj1UX0jF
765SwOo5lhBtqS54rAcKKtqiAXpJec9SAecSaOVxfTnm5z+M0CtvPt6s5YiMzwSaK0GYVLD6VLmM
GNMrAT8iX6Pwxojl/CpkmscvtM3o+28UfaEiOTthyS3zzeGHxr5knOnU6S1XoHZ2j//y/FaDmnyW
yOKre3JsQcsl5iLtTOHkTuimVicBPU+agYH50HTbzHfgSYTUGo5sBX7R0mjGSc3fOzOlziRKCPse
mfuCBwa7jpWoixvzIOvG3bYjhYVetNwwOhCzibMvZnRM+NdHWAHeGmnCxl4fHXiBWRoAt6M8BAvD
IJ3jewZKPw8GklWZEo/IqsF0chuiyIHNqXnCnUF/n3W36aUMGLBrjjbGjWaZtZFissuHdqCO2mM+
8l8HrWgwwlxE2yXH5+3DpLHsG1t/ahRPh4BQ+2iUL53PypGSiXNhgSRENs74MCMI5qxmhNzA4xh5
lBkcm3beNTfiB8AJaQcSHXovhguB2tZUBk1+MyqF7utZe4+RLSdfkEcrHQkv8TDjls7YMj1ZRez8
rkyrkJmbpquwWd/dunaFOCFrmfqQt5HWhkJvjoFGoMmi7g28SJYxlvvBAKQJYkwkxbhgRyhg7ZRU
DuQvP8iuYyDbxMRjCLn4ScjQdA7wKBRGfBV4KkP0PnVJtao8A/85ZnjvpKuqgBJRNQpTfPx7Gz0J
FgBqovYnIny0c8Pjm7loq0nTrCJdc0szGjAC/BA+l6lYNnOU0qikN8LfK4vjS+1RSq4ydKRRaC0k
26jiJRzqqaOvd/oft940loL05KprTDNan8jaAroB4bqyifLrVsUu2gOPLhIwXmfnbL4ElYglZMPr
sCy8XHYqpVEC7PTQFLXvcdFpgFeSoh+zyx37LBkNSaM65toXzmZ0EnpIlODIQpcNcluB1VCsZB5Z
26C8HAaQXyP5zfg5yGmDUvhE9ncbgMjUZmcdu1N+o0X/ZWJ5d+IJN612NuSfdrFDrXlZcraC8ghP
krb8PeqZTfIvkWz4hnR4VgAKdhMEZMzIl0DalwHzZaANSUkMbCKxFFX3GtEI+qmpTSN7AdYj8Abz
5i+Js86n/kOV6tWudhDSW00ceFFWIAw1zG89w2ZugpCfOVgSkh/uu7TlJV2YGVm1eGGPUO5ax05g
dDgOiVWpbu4tQOGnvydNBM5+hAnBj0sfTmmbo0QMUfb0rGXrjuxVL3HpJEZ0tOCui2/iou8B3t36
3HKvytUPVFvLGOQ7ZkDDQQDlvLIrDNs4/8PpctI8doEzYPnmxvYNfX8R+AkX+4KOieayFe3yIHlI
bef3OPb89Ydxx/2qqVOV8vEqzrsmThUYAJyG/eFdH94zUuN4UFC6DGOfKCLyz5REOylPY++u5SYF
KWrW2g/owgkJYbnER+CTo6DWz341zORNxHsdRVApq2hgmCXB49rxSe38snqXYb22an1zQuIHgFWL
eGp0s+ahMawydqIjlFJW+EVI4JUxC9UkxZehw/lTRyaixX/BRx4xjZFcZYpku/jjQzKnVgMj6fNK
FAorWiKNPb4smWAMr9Y9H2QwIAzy9jTYzvf0xiWUpJOp26j98GFi8bKzPBvVvqF1T5Av3bwt2uGS
A9vi91KEQ1H8agx1Ryo0M1gjEAeW+UafasO02pUc/qt6uEi72JPm+T1Qs2Nqpq9bSymfXJqk3/b2
J1TR+pxrSW1BMFmxMWV+/x3YrAyv573Z5JqRMOSYmLKRUbUPgeFhIhPYifGXeg8cp56Fu8gAdQiS
m40Hw2m+6Moavf8T9WQoM3fL9yFSMzYJkkRTX9FhlvZDB9Nl8pWe9s8xClhE2Wuz9MS0F6H8QzVg
H7vVmsi/uNo/PPoZJnSi63hcjdlVLze7ynX/N32vZVRJh64zrTXcGbWAPJEOswqyNClPbMY/0nSJ
GHZwbm6kkE+IsrR4KOT89OJmNsafBagdl5SjDPr1M+2PIDxVS0DsuYb+hVX7PlrIrzA2O9bltPJH
HW/FIWV6PETUD8Nm1AGbLGJTDXYRJ6UF2RNZsxgMiX8Y2JioE/jRE44BAZyoVwJMHXjLvX8z5h+2
33AEzfEK1lsytRf7mFdbVlDgkKvaCYvVwx8+3prFCxu2+TU+Wo3W2axhqifWmz7zmygFpDA1ATca
mrhE5Sj0tsB0OnT3J4iKQAJ36uaFGP2bCnIKpBCk615DU+t5KDhWDCp5NUbgSQ4PZ6zCZ9ZSCroZ
YwSLvewFU9oCVawkvw5//tX6HsVGgki2/6RIfbtXJDHDHdmZQPfD9B2dUvp7e3AbZKViJtSMGNfE
izZ/0mA5vXlRyi73M7HKsUCr+RnjG7rm4/AfxOqrAEHyOwqi88bCzRYr85oVjfvwcsV5VzrXwwnS
/rlf6ToEmDr0Q3l37i0PO1iH+My/uREk6JQKNHhrz5gUfZxc60Z4PaCy0UtQouc3RA4GqoEByCWp
H9AVifhNEINAStCsaCMDOJwU1ix0fbn1x3FSBKdoMJF0AvFdLIEt0LYQ2IBupIZNp3omulDdiK1i
SdgrvkAk4brUZ8Mq1oKo+R7Mc8TRg36oUVn+01ORqXzE9KGq1882yzQY4cqfR0/eb4MSRxpynNYG
dXuzJSdXOznOJ4GGl1Yhb0yGoBU8jroaXxQUb/rmwf8nwGGdLl8FkzfD/zO0ZMBoLSNn5Izr58o7
5andbdo1MV/hN0cfzAKuBfGHWiAE6wFXO7xwVtCuTUF9xMp0XoiAB/7YTBI6k4bGyMhq/MBmgws2
KLtAus+9f8Xq70TVUz7BZqZ8ss6uuwMQEPnwW1Sf/FSeoil9GnePstzQZzkwZRMREzaDNDbEIBys
JdLbt/aE8qGFY8n9PMnPdtfL7D97HJtJb9RdQGBFGr2RCTr0ifRxyf38n7Z1HHrpeRV4DxZul+WJ
D+aALSKBR3nRiLBDpgPe1GCbq2ZKKao2q8c5l/7Lcvi1VtQb0/ogykd3pR1HLDGcG5Aq6sWZ3Rm6
KjjNnk4N3OCf7RbSokUZ3d1r+F2L7QDuJlZ/iHfSg97EJA88ZSMfRDrJfJldnhjyV3FJHrC6YvuZ
1S11i/WmZ+jMp1oiULnSq7IB/CbPexFECWRawCjls0aDZzp+TodL3AUdngJQX5UXPRKapAMlXMg7
rLtjE29uWSnCqFHQphwR7dwYoam5Tf+YCnn5iqjEyHwrxciIUPEDwvgBh8h0EgOkHvytUTcffdpG
RM6fNcVkezcrkRS7O0sfkLx2DTZ2TqYvoDI97Tt5HE4Dhlo2S8Mh0I5n0gaxQp9SpJSax5gH3hCr
Hjb3mUqdaDdJdLUho5NddG7obbv2uJqx4iYhjTpFN28O+VeWsz4f2mrxhVjFtgTWRaCPeeIrp90F
LgumdfsN4GiCwwLSvW54oG+sEdE2x6DzOXKlYhQwdKCDYrH5nNw++LNpJPrFj9f7NiQjm6sIbZAQ
9GBrXRP/nVDmDb06P+VK6MZgh6r+Q6oqDuOklVoa3D7ugpyQr2VwZsQFBRPma7NYDyQrKLwDeopp
7QDg7ddocKPka3v9roKVtzoPehnfhRmnh1myocC40lMcFHlIrmWVa9AM/glJcHuMP/bs4ws6I92Y
JmTnmQYBwP+hdPmpYubw5SkU8VS/6FL9gJ8bGjYcq8z+oJPz57WopfWypS3/HgmPdnTJoq2Kw/wF
LDEw+nfGL0BFbyCxmxZ1iexunj3fz9UF2VxuXxj+tbFguSlLZO6C32UZpgtLP8k9/UB32arzFOrI
Jm4m+5CPjR5tT/m99GanZ2mMKV4rFbDpCwMrLVaxgOhpfQ67HZuIHj/8h3RqqKHe2Jyw1fDU1/ta
AjPrkvyd5gIzNZxkAlYIOQuXCjNC1pNa379LGiajP7QIwS/xQ5rdvOuvbldt06fOPBqREAuvE50A
xEIjXSpC/9qa8UpWys0O+W1i5mwcQwFE5bLjKrGnMnXjmTHhcDstM0GUlPb2+73f3YKHhp6rk7wc
eTkdDdWxw/yR7cOJ5KjscLNwGwst7kkDR6O89YY+bm0Sf1jsfRasPysBXJQyjv6uco64q4v6WdH9
Rnh61Hr/gmcklEHtUAR1AuGQSVdnSxzibmJjpUqUlUQDvoI7RCnZbFouoe7fOcC3swT7QZQyRUng
IvYGH+zv3JQQvdlk0M/a5skBzFT8HpG1k3D2OAiawSLEnqyYi/Ak75hT2CBolSz+MsUcOekdba1W
Kq/9O61NF+tdf3TH88lKCbxeby5fRna7GKi/ndMi1ciEfLIvmjcuWAwl62QQzLz/4+61mDoU6mLh
/9AX/leWPry9lRdKO5gP42qPCKI+26ej8n/B1jgILsnXP3zlbHP2znc79Pc6j1QOT+cuXPbdfkqs
WmJgECZ7kjc2/rdCWk6mNu58bbiuAOAKwvZfvd/F2b+UlbZK5p4ykwy8XR4Tyqsq58mx/FJBnf5p
vsprdaUs60rsbCsP3uvEextr+ncRpaA/hiURHDph7QLnYI+LfygbK8Ynwh4i19/YHIrYtN/Lz8Jo
JtmL1iTsTa4Edrzf/bJE3HD8jLH3t3vPT5qD6EG9lJW8aJjYm7mJdXd+xGC766YAvNJWbhI9Nq9q
bz+G7IhKdXUUI1q7icsQvZJzc6qtvJKM4JW0lM/yY4alkXt93/F59z9u2bawtd+V5sHEg9yUPWak
M9o+ru66fzxXm2EwEYQZgixHYcZcnYFxNmZnzkMGViYnFKi3eNtiLTIN4deS/ixuqlOR3s+DMbHI
89dR9hEy0GvGK1wUNoMYoNhZ6brt9gBZZwDD75456+X9g+4ZRS5ACkUnSGQ/nYod9NPy5o5zKivS
DicIX56O3lnE2rKOnaVVnx1qUujYq3vLPBHhKC/MeLGjULK6rqKOkK7Da/+6217jMRdG+orm1UpA
FN60OzQ1Vub62OSU+ML2jKcqVIzPGP8GjNcHNQq3CYfmceA/OIQuAG+N7DQa1zfawOrbTsFgxP4b
rE1oqI7jDyxXQMerWkZ6VH3Owy5DAdzhPsZExwoI1afmYdJzFUN2ctMzTAO/TiogZKHbpX8aRysz
u5JdO3DF9YylU+VX6UASyDYUIhEC0OcI8dN0xeLhZnNuSOEfe8JcqxNUiLFHvCznASX0cHlpj8Ru
kVrsZ5quGGK9WzEhJkyCy+YClHRkyRS/VZNOSJqoPsRD2X59XlIlAzh0heNrXyDy95R+hGhzCMza
ncYw+zCe3TYbMjvnUTHfhtN4uUSiQDbh7lmmj9i+q8Hf0LwTGIGkej9LxrbXx0oLUy1lojqtBwtw
BpN+reXbIjIkYEQfFDSCT2NhvhwOkQlAVkKd6L1T3KJUkHit5ZW6qAlRzy05qg2Do89mGLKoMbVL
aP8OA8GbvBp1WIBuALkX02hzAkcY54AOxsQL4l9GZ5VQiC5wAjONgHGXrWBzpSLHRxbVaanj1oHM
2FcASzSpM+7pnAcjlmlIpAkb/9wfPl6spDCGFPkMjBUr2W0age1E3g6YJB394jS5mmywcKC+qZw1
lP/dajG22F2um76LOYMqJ6rdiljOoYlZ/IcokW5jKi4tLdkhgj+GLGVQdRAcsz1t4qaZxbinI7yb
Q45UIFyPrubc6HIP03oFfvIhxQlTMueFAAJH7Gd+jzdMT8uxiDV81HGntWqOv964JDbT9LwpkKPv
JFnomqtqZDQ8ASvM/zPiILMcZ6Q8Hrf+MCqDtPX9Wrfhqnl/A9LW7g+vFbXXu5na8Qx6lomtK1pw
FvOODlvlVUiq0v2OygkVNBiW/cD7x209mP8kI3GGSMO6fRiusUXCO4ftTB4H9Yg7RpjvjHk6YPB4
tbrunqfkcUuX6juGdy8g1VT4/l/LxxtfKFlZp+KyPokOY/ZhwHtoqfUnEdEuYB7bRU+20U4ohp2w
hHyLzExUU2zFoh5dsOy9/p0CUpFwru219eUEd8Qi2yY8AIaIJ2f1djl0uElLRgYCzDSm0ece5lwV
fsAGqTET+n9qVSI2Mv7LsmZnxG1ZvNK5++s3BptAsUErxrwV317orXZgOpQqpF7n1C42BarF/0l3
9qpmLtsmvQJ1rW/Hro61KQpN+LSDOMHfdtqPOonKJgIAzidnNpyLs8HXSnA6I2dMTsObndU00/sC
xcUw1NPBRbdAxohxuXUh0TU44nBxZs48rxotg5OtNtQhHapG93UGnTnJbzfIa3L6G/q7Yqx+xh9V
pjhH4os9IlsbXdpWgQDM/tLePVFY5+i7VoOzSevHM9ykQA78Lsm4rD4VGC9zC9Sf9P8hSyiEcBTd
bBQClyFW1MSLp+ko6FaLvAi9d+5mmU8H+DZnqjziSGyUYsXnh3vRd7A+kkQ/H/tW+tNnVcnAiiU1
CiUuhQzv38PqFjIlM2irJlIAbDqLQcuSGQcC2Be6KUvtTSWldjGznb+Sxh4uJS5Fm1amp7Z3wsor
TaGEiOaEmI9zBSc1ZT3yB/lvXmH2K5cRbRu0avzwuOTMe2/y82FPSuSVQ1Mw8T7stUr6qQUJAWrs
MZk3zaABTBows+kOoZhwt6xUoiP21Bn5nF2BuwJTErrYWctz5+7NxUMNqQ/uZNosQcV6R4vkK5t+
1YjyHDu0cz9+aF+hklT8dQYj9pFmIo99CEOFiKwTiS4W3sh9RoPUTtYH+44Cf3BTSbCYslE//V2b
9Bk1I909B6OL+7/08ZNO6hTOm0dOxTrtFqaifRGx1wSCcFLfNE/CAgiHQ3NkWg2KO63PcMJ2uRxC
7/AkoAlQFhHKGJ574cNDdnqnUrhzDNi8JW3+AL+/Lc5VR3HrLMxPCM29spli/gXSmoD0KfUIQ/gG
juL/6XjTnXJjF/3k0EOQzjob9PW8F5sjzwxJxg+pyG9EZQUdDocT7Efq19MId2vtMhLm0BNcieMf
9CSlypkcMi+jywy56D8EfUuzGWFmtn0CIh1zKmbH2quibaR9u4+dVbSFH4XTlWOnGoJY9tBUVNzP
LkobY2H6alicYkGy6y9n4Me8+8Kps+ISfHZ7QfwZB8kuMh82CKYYxEkym9od2WkFjKDkpxStLZwK
tOcFznsUc+W4pdxmRZBqebkcOgddJJ7mgpEHLGeR7ETcd4Bby+suxPvrKIg/ZO6CDRwmZAyEGTht
9iXLNDmtD68B8bujF+jK1t0KFO4qOYqnM37Sn5/0HKsJzTtfB1+d7gZ5gR/lGLZtivGKTnGk6Tjn
IDqMhSiUE3ksvZZ0PKm7byX6+j/Mb3hLOzZfmBuOPGUVBeOXGAWvQDPcZsrAo4TOTnCKHkhOcIXB
fgsx3ZYZSnCkht3k4FeGfr3xYKcvuwkidNnNApipro0cCOJg/8DfH/vlIkOvpAteo8flOvd/iZel
mXv3Ufsa/10FackVVrr9bTIYZ5acjqewC0N6gPalNtdVeDZJL7iPyJExjbEJa+q5FqiNbzAQ8rgE
4BrfrQoYCaTC8ntK1v8ajsoIciSr978QSjLkphY7ceibJLlBU5Zwc+CCFqcRPeexHp5PqEttgiFF
SPKtsZz5zLn0JHPvAxqNupHLuOZl0BoJj8L/BXFYeUeuMBYEyJOzCydJlWODL4jIwpnKS2h+A8lM
JvV8CgMhhSV1RMZsiApqIM01Ycxmo6YXInpSVFUr9j4LjkC3uIK2SKidfcLvA3WwXrD+7+aSDFDl
DRWQMOi9FEzdEoic55b7SdHKCf6NohAw515MkdZWWeICqT3jDn1T41tKOQ+MDfkeLP6IDKd5GrC2
7FzOlF/HkCF6JWUlutlSIoIXwAhSeE61aeuJ1FO9fddHpgPShfpJzmmtep4LRtNjkJcF7tOe3nYS
+yJmv2nXqZQ0NMeYpr+jQdTJkk4E2UlqipBw0UDG8mwy45iD/9qbIHm9EYC/GVo/AzWN14Iv0htZ
aZa87bKqxMV8IdLnM4wMOHNs5dMETb2YxJTmaYZlMFPJFc/mSK4YHMu5sGDTPbi3/oljlIzElOU7
vUWIqO0DzXTIAzJRnSpkXaBxUo7SDhjZZW45IaydohzLJ20OBYbz7XROad7/TT8+byNO8UwjU7Ob
BaKDcJFwGof07vHtyY7iXEHnfcVltBxYBhPz1S/ssBj9ikSP6+CIpwm0FVPgR0GhGViQk4wUzV/h
EkRiJIuAQ3VjJSbz+KTXi+ux1rOK0Lt6LwRQR5mm4VnGOOJnbjiz/GlRlrr0DCBEsbYeAka340eB
Ri7rKl8tE1Tdhg5o+Bf7lIhvtEErhCqSJRIA8rLLb9nT4HUlvZRKR4v2i8vzNfB41thpgy0CQoRI
rn3SryvCFpp1ngHVe2pc75uedvGnVgyvSNAPHvVypOd8spm0jt5HJ94DE5LIlSzOVHxMbVuDBL3I
mbe7LCKGNo/qMY23UHlGXbbt1VF8DG2U53mJXTIOJl1JNtO9onacHkMWApzNSVDAyFnfCxIrgrN7
Gu6PBBy8re3/D+yzKDLJBVWUg1aF8xWfkW3PZI1sxuCrPXIAgkJuY2SRCQR825HUWhWRQOsWpGua
vhp7e2+WsT9Qc4VlE2jgliKz958cGaD1yNMXwkq6mjjx0lGNJ7+WC/l7yUbk2Co2LE4RLNtqChqH
rVpS4KWQlrMl0J67Q8Fjw6U28kss5y5tNGqo3Lq8bFszh8A7fNOP3YSpOByNUQt1eLdvHnjZ8+yA
+jEEVcN+KTHvQgp/dOGvvy74Xw1O9zBV8IpA1hp8yWHQoYQhyTQc9wQVrTohxR3gf0PeWeXqEmDm
jZHyX1Z8fiVJYdpf6FwaXF5+3MN2xZCzh/FpiIAZHMZskoa0lYg9rtyiyLf4pukbsBsKDJKkL/WK
/4L7J2JRCzyDwydZAvtsaYXTKj6W6+ewCjpo3CddB8jvKhXIgayCjFRUyQwj0JrXGzt/YEHHkofM
JbpTzWTk8B2LvVDL7gtEtaUTqyuE3p6BcRB6/Kt1n+oA1ylzKlUcWYNbcOoSV6d2/Ai/Ha6zNNn1
WDD0RNOeb8OGIrRp953oS2XO95gujgQqG7FC9PhivZqQ3a7IfsirM0yhVycrS6/CvUu0triSVJ2d
UCffw3WoeAGGz3X08UtzGR1wxnPmyrmd7w2U3ow/r5d4xJMSek+k9R6rdOcx56MlI9SmYdhSbiNm
xB0Tb7FvUmf1FWAWOX6Vb2aRqOy/CkpOnIweY86FPkbMmaK7bDLLkmXhN4fhz3rimGw+ZXzU9R0v
xPBqi52AutS0GumowYi3rrx62Y51aM9cWHIdq11MXmyJZl1wTH6I5qsKbZrH8LqIAENG+lwOLnGB
7Q+HrM4c7ACSVMtYjsM1mGu7tYvi3FJ6LqvDtzu1RtCC7uIvWocEmv4qveOcA74f8S4qxD95GmG0
9vqZfaTvAHL13qI+88Rt97Wz7OTXWfuJSaD2rLCDjkVEB9Yk0c5gBua/JIYk0dHfJ1xHwQiKJFPm
moc6VkrdZpFuo2b4tdCjy9aX+AYXctUCMoupgmSPmPSac9i4c4IXayjPR/SbSsLAMg9h8Yszfty7
x+U7raKM8OLXCrbRarEVeA9M5cpqK6hSREHq/0J5/1pHIoI9z3hzZCF+xSA/pLgQqqkqU3lz/nrv
MmQ8B6oS4QpLf5XuAZ+Ejzy/5KXAr8vIhnsVpxXUxIlxdEE9Vpl4geRszDK8dPRsQA5NSU1wh7Yi
Oppg1Bmpp53qHLM0Flgxf+HUi51usY1IiPER9mL2l/0xbkXsBBExOXbF5/nkcBlT3dICjByXejRA
nbPKGsqnDzLxGF1XfJQigQeUZCvpA9VaF9k1c9B5qcaSpcHBVzV/iSfKc+y11B2pjlORKnIpTpTy
u2oaY+LAAxl/PfrVJaVZbWkj/5PVed+onx1UeEpE4co+0u8oWJjG+0Si8UCx5X04BcG8qcGGmAkw
vpxi5eCrE7XghII5XL3t8zYlDhEUy53pjfDhMhAKZrx1cz0oFzEpN9qCmQWqVa18lgmdYcUzQsQe
ftqanRYdEkc+hdgFifSEkgyYd70enETn8aI+liFAtuCPhLTS7uFSo3G+SFqF6eY9ZKgaNYfMmUNl
sBGyil1bBYuScCQzI6UYCVjUVp3X/7tV8+tvDINKvkww7UNLI0MITYfz5P1j0HaCzgxjg4fP4VRK
nlPom+crhMIJpTwd8TbTDqmRMH5vlM4MJOFAss0+LTpaf1Q06RIHhBMffmGmI275wnm/A122XG1u
1qzSzsSHHbSzL4RHzjCmEJZrM0M1HXqZLTedgqNKVdJ0YTFxKhATd6PCFqlBAyBJ52S6bkq0Na/G
BweA4lXrrOnMLSXTh+cfKAD0KjNkX7lR8VoOEpJ1B1NlPGvM0lvxBs4SJp+stVqlKGWuhKFNNJOo
Bl3ovupxse0jiNnZz0JhT8IE0Ldt4T1lj4qEymlxQBMBwZgo29v7bhxK+/wbvZkX5RvNTkeXeTZZ
lzzNEBNpNsAqPnyrLjOGcpJEalFVhwC/T6u6yUrKqZVSqWVhhEOLpKGx41+Xgi/D8tPdLOcrEA3W
XDXR/ki+yoIc+yK6+KAHQ1HG3iZaMMJP5zPDvL0yE65Pq0j1vQy4gBk0deD08utyk0fxTtvMfz1B
s98uVH8TurPKCLkq9Lj25puAGeIFIIGg6M9CKwwo9K+gx0NMX8h9yC79+ZzG29wNYtAcRADq9BRD
ZdheAemoAWxSiJweBDHo+kvHyhBkfLkCw+rd0+BZH0oHxe8PtqjECT0ZsmZFI1EihRZTpIgIoI0X
YMM1QGMgVkBtF8yP3r5fsaVASZLCekCjAhimJgVYHX2CrnAcxQOw26Df+zwf3PZOjV/SrT4Uc41v
x2ECROsAPfjoKnDrDgg1wv9RrUIbODj61MBJcBUObXdwE1enH/Lov3vtdxgy8bn6gZqfsGX2RoRE
70JVw8QB4EQEnLb2VwgGg77AHONZyViqjxPEwL7WYQBmLUH0jAmvxuoiOT+evdkKWlzNuCXI8qze
R3fwETNg21+InCq8B733ueVmxql/1qyHXDqdR5YHC5oho2sxlzkg96/SvMj23oIVGI+0OIcpe6A1
K/K/7Sfmv7axhlEKXVQktBdhlb6GGRVw5HFjwOUV0fD+FByAkd/y6x9LtEPANfcijZM+8bTf0CFd
yqEkEM9b68d0m65ZHWiHuJ9MzA6CLLyzvbMb+9xaCxsMNY9dVBq1tuEcRnO3nTb/z2RIX9yOI2SF
1CoKXeYdu33iUYIhKSIOMa2b1vTiIHpY7iS9mdTkOC5CyGsZAVrJKN7m3T4aYVke4LM/JYbcKqLv
KVkd5AyuZCi7i4FQcPmoqnhE2Nv6zcaRAJPsVtrUoF+KnUVcCx8hFdDjC2g7BFKt5HtKb6KFiPp9
jx/EQGTXqaeqIzITjhK396hAAb+4Ar1yhhsDWPESHfjygstg6THzwEY0UEl72h7B1JXIOY8PfdNM
K+Bo/pS0b8B+o/dkzPVh6dBKNNCKApekzY2n+7rhYGgirgEvBaHU1/6YENcUzGkFJl7yhGYiGY2B
Df2/koMK5P+B0GvVGHOlPxpsFtc48B0CvUX22ueNAtba3QdW2hMeuneVPDihwvDW9UqZIjIw+i2J
3uI2CpDD3MKjHbFJsi1fVlwYRWOSYSfJKzT7cuuz9XQDDPq1JLjeXJ5MYGQ2h7NzfPWEcltYF/zO
6xvoQFglR9D8MLXnSYmmAdSAF+ETTiX+YQxGKPgUXWVrzmMvGB7AvBL59prze5m/xwGnZOe8khhh
jxbuV7p537Mkcz6Ich2rEn0R5cHNxgYqMHmcpp1+QilMmCEOmJVhLGOSRC/+Dwnul1ZTFkZe44PQ
jKw52JWr4v9K3pGdLfwO95usMowmxYTSnn6w0RjXCrIU2wHhb6qEnZg9CE9ucW5gKegwy4YENNmG
GUdjoUEnoA/SNgnY0xJsPX7P4hgC3U9QC7XSRNu5dpp4CgU31Jtw84x9+XSRJF8vfEhxbod/JN8M
u1xQCQx4g4z0wvWLEr/RIWDThI6gM4+evi6JnzeP2usRqZI/TwLk4BckADCtO4LdacLoyU6/6p9n
ahwZHpLLbsECXKf9PzAiBP4UbEPvSUZmylj2JmatSpIEdip/Xu+5llQveByeVaqK5FPnUa0Lziyb
azf+QmfSS+VMpGe7PcIFq5AlhHjY41yRJb2jnjK7oS6Xnoipr3jZMac9u+4GXyKscYGGpeYKOFnx
2FtmQHqZFJyoev+dflcMPQJ0TGNqvin6KsAAra6tav4aOuqXrMUwYACf2XR5zal7upAv0EiKJSBP
/3swsYfp/o0LACpNdKwYx1q+3UCbvILNOrWRd1cTw6O+ruRhDQJSizKmBBWOQYVj2paa1bVPm8HS
Kd3FvI2wTInVewBO89i9AIFMNVVMkG8L5nxWdIWK/TGF//rSOJbskxnJVpN+CcDXloE0+L52YijX
okglO8RCSY44Rsf67+9AJNKmhbn4sb5NBf6aGcBWnzDo2Lk6jPFCqkGwjTGXgtbEvVjo/TxryFiu
GmBNLUw9lD2pwfpaHMudE/C8yJCxs0YZy2m/xPnncduCSS5RBEIqy2UgMQc8O0O9RWOe+QKRsRUH
oEIGg8bzq7MtGi0x6+NEfXTyxnWVrbJmlzRbWRekIlBDnDZlgQ2R3nkOwEDYhtpWp5b0NDg3cY4x
ZeadEtI0hNA8cZ2273bjQEbpfKOWg5zye/Zd4ByeW+mmIJUbTj/1OP0twxWpkRCpDE/vs65pKKNy
+EqieEHvZZ0jWnzZf48uO4Zqqf5CG8jEYfx1j2PYgpyWm/Fq23SP1Y+nH2AsV9WfrDcsutdC0sS7
QVOcraS8k3X9LYr+DRBJg2ReyAGqgMaKULGUtSlxA1VRoih2VZgKaFrETTK5tosOG7cJPhe0YWHH
aHNHf7O6uIQxlgJPnoKDghcRNrSQGoZFjkJSq2Z+pTmt8lEr9iMPJTMPhOejVSAZnmloq0YyqRse
ZcgbJVCTBoNh7ItUdxfNu29jmfJVpNWE4TrfHBs9xHZ221BvbXJ8fiJLSS+4DmOst0ZQm9/0bjwQ
82SoV2tDGcIqh1Sn6RyBsomA6vN3EhZjr2w7giereIGB+Sguka2Jid9a35Vy0HBmwNRRhARj5uxI
EzdcEznCTFyBduyLpEpQhlpa+BCCiTfc5X+wmGyfK8RQFUFmrk99Dpz53guEUtZY0x1qHNm15KwN
Vvzdra68g4sZyoBPPkEcs5Fd9ZAadu9YjCd7nA58vdSFiatZKG+uryJfWIXcvsdQ8NFSCFZZcHQm
b7pff/W4vGngHN+ABDperyP1LtPLgV4R0q/L4Sh788JMCf1az2mqZPYjMkQifrqOkhtNtR1Xt+QE
1uD5NBd8JgmDcMRAEelY+pUuEFCgaduj+KKVdAYm5IoYuYrq5DG+lGnx/2b4q+n67xVcFNE6sE7y
hKn02h7gvWBxl+aMWuc+y6t2me3BAmjz6CaF4fAJSJjHsVc4yyHWFyQg2nQiTr9fMxxJkaCv4gWI
rfILLw5ESBUFIF4cXszzrT5ehrTMILOn0XL/P40FFVDMbZfeqwEmzczxrgeH54plt651XJ9zPWPo
a8P+HPwlTWLhmnRI6SnDFl4YMHF6bYZdwXLmj3rHs7CLtbY0RcuAc/mDNltR1tZ9EY/Vqs0ek0Na
GNV27+J1xHUt0RQsldrNVfA2ATpGngQofJRd39V1IgLfqvC+DpQydvQJrDPzMaxpnwZJM2pkGlWV
jpKg2H6QSCJyl7fpa06ym0WBuAXlyp5NMaOW6Ql+yP97pgVMsGq1vgJOZ9qBmm462h7WbW1w0sm+
g5sNYKoUwJnteonoq9paEp4q1SiLSTTiC69wm1EdJBnVBWSJczZpLbAcDr6uXHv8Nazu7h5Jsr6X
0ImdKO4aSvu4NcAPANZ2F69fwHNUaii4Golr6PlbUd+WiN6jBI5jb+HQkLTlQd8HbcfLZRPosu8T
EJNlhzKsUBjBHt2B49E3V3A7JguFz5rUKVFl15EVbxPxsDW39iBYXrDsAx0nt8gd/rnYFrI0eeSG
BXhTlrR4v0qBLYoqdtQbGcr2XDoyd96ztBsmlpigLhfqQgKB/OcRW+rgQgbe6yU3OQyW3SkOXVPV
VQVz0uCEofElHo59fpwheIIDoQ4yC5YTYMeszPOajrME3+nzlLauXfOXb9IxaGKM48SkgM7dlX81
69if2EYSEbP95DWsHOlESZhPFXprwz+5+twuTDRxIGfhomdTaHFYV6+lcCEy7FDQal3by/qzf8/7
7u8d8flkguQdJZhAlpKGo2GNysOnEnSZOWRutGuHhqlVUMMWx42pEArWmZAEcnCD3l0/2tNh4YOB
EjV6j5uPc2ccdYnD194aNqCfgVAOnkiLuzBC7QYx2xzwWSBtxuiKMXTF9pDsmCIX0/Rm+0DypKce
zKgn+KpSwic93N+Kd77NTY8lhAVDx2tuMJnJ8loEgXsI/gVkCb4EvYrsUhqrRsniAWnXvJaGJaWM
H7U59qr/wTE36sGenCuw1QQuPqtmzBWl23lc5p8jd+Ty7TWGaYNxbitXvNnp7D1ojFhhpfwCPweJ
Vcor7m4J32lUGKijyCFtI/qU+IRko02ksi4Y1rawUNBL5U8rYEXc2a1y8yGDCXkYY0CefNl3S8jl
PAtAXxkeIOVPPaMzcQZJeND8Fmfz2Q48Xsih7Jq7/R19FPLaB/pKODVbd4xc4Oq9j6C6nQHbr4k0
B2GpRdIX/sAnosoF234akIfZ7mYDdCepBeHIfpWHjUej0YOTNmiHJVi8XE+EPzqbNo3OA8yjPlcK
R0L9nJYKcv2Q2+eJFc6s0A8f8np75DMvDLf0lxSTy8Ub0hYFyDJWod5AqFNGMIiUcqdi0bOy9q3r
G5A0XWcynWn9vI6agZeXigsIQZPzRBW1+xYmNmxrT3F0yzpP3n6wefbJ91GsClgF3RKJIezOxCi7
5OcgWNea/VkOZo4LQmgN+hRs5GJzAuN7O4u36QLON0wITW0u3P97x69duPDpYRwiV8OHJ32ZqDNA
40exvcBS//YYf7nQSU+uuHOPCrEnqF3/BQIeY7up6Yn7QFd+A8+oyD2sJe9+PkG5FTN4pIetkAmk
gN2o2R8UCmdnCS5pCVv2ZGzVe5lPYZ/rWnuAiU5XzMboJ1J+njvg1iJQaXkY6bDE2lBwaQLsTW6r
DB6LbpnSQ/4cHxuSWKArmEc41XFi23OrsSkhUyWxGq+TYwhkL0EXNc/h8aHAJxSNofWXxUIQ6ZP9
pJ3J3DM4SmbA42QI6qnYHlUZP/++m5qX3sOv3g76O+NY8lRQbEvND9urZ/qY28mD1u1dKrHIC/OX
y/mW1FGQA78muZ3zG8KxBOQv/l2cL4kQDFBoqxV4HVAvP5xKM6Ngfe7omgJ+07SKTWBFw986AvG8
bliVz6V1MYiBiX235LbatJhKKXm3W8bsc/rJ8m4I8TPVk9aR4ZPWs/YPYmmSqmmTy9T015SJFWlt
z3dnJKgIqEacPj89NuA/WxVHzYHcNNPSYDEIEk4PKEarzvGZW0Yfj1oEYSwPL2gg8XYqvhxkrLIq
Ckz1r/sPS2BWqSoh3ah8NiIXGRwzAWDNgCUcazENXbykkX+/tbf7m+vHEwsnIJYq9Spc8a8SIvCx
+x9SN07nGTysFEPy3Y8XsDrR0IK7xW3FSOKOw94l/9lAzDfUfKvlELKZnpRsPHwEE+pOF+ewIkoK
BxOh8dk0lIlKc+kAdVgLPSeDUFWmRxpEX+wqQf0/B6Or7EFo/DA7h1UxFLTyeWzNPP7r4zBrzqKW
YXZLlD9yijiZgSC/fX2Oqua/IJh+CXYdM/7+3qq+JhaqVOkD5sG2s6KYTaoPnlrSB9V4HYJv4ue7
XIiDvfz8uvxqvKqPmZ8Bu1WwtYfNzfs3rLUVrp5gPo2PBMnfEwD8WZkOPdAl3Va9nbyAQWjG5ZEe
MpMfLstNK+wZ6AZlwZxtCul8tc3IXxsR0Fn01Fmil4P6bjL6gF2m5wHK7xMjcFo6Lx1m/z0gmxMB
HXjTMFs3bet0iQyT/51gn8iwQeZZeqU4MxX5r986FL/ezYyu5Dik60WB9LflZHtpJ1n8wdQ+E8ex
/LTHx9P0D9tdUG5DW8gbuol9NwVB9IrF6kXTwr08xKH7ZIYFXeU8X1WQ3KbTVXiASxWUkdZqUmp3
gv7Ks/+bLhbQCw1at2vaJX+schA/a6n36vmy90OA3+idzeeoQmKzXDipX/WMW7b+Sz1iMU6YV61L
k3jFtW4dczfTcx56e80n1Tpf7xejX5cmK6nbg5l1gEP28KyE712OKnmrcXG8lsSLhau0aYjR0aIG
A91H6IfNMFOq6JL2RHIRYjnY7EpOEVFqB14INH1tStTwKzzWbcVmE4hd25JM9zS7kQQKKpY34UAS
cEFf8/BrqlXraxkTc1bHsndBmc92Fi4nZa5t+4YPLBDrspAO8tFHLUEGrmddlPO+c/F9Ujkl8y2T
vodlAqkb/c04iT8RsnS2hL/5c8TyWLTAhJooGzzscWPK7R9DHo48yBveMkMayDlMC9XyBTuWOhJ8
FzA2RPe8oef09FoGOC/m/+/3Tl9dLrSepILb31rPTA9lpYBXR46ovouGSsL3g8OIEgtdAo9Fdnex
2DdarC+W+hwTg0zmP9FOH+iip/hkcCHxOOlsoW50rNYzApcJQJQyUTb3pjNzW6BdtzBTE6ODHBcH
KLZ1Hq2hX4FYmAcz+E3s12Mjv0+YzGKzMVppCZBM1jn08tV/sVZ96KuHYf0FjAm6XwZn+BVPbiI9
DVTTWPIDuW0ViUnxvW/bsyvJdYn64IERT0Jfpw5SGWdFRBiXaPRfV8djBg/thPw8uCtjO5A5tcb7
Do6jWmClgfNyKEcN7b5jv5sna0TDocudaI4ERCprwOxwtKjtNVTRfJDpro4IW9xS9cCAYxfQ0XPr
dtX/gG0lCa2e5B3gu3SO93HC6XfDdyaywFaU8w44sAh0koMLtt4+X8b1OcOZkhRLSQKlK8eT/OQ5
JEnqdnRxu4FqCdzOiKst4ZltNJ5IVJh1SLSmfJMQ8q5QvugLab0f/WMTk/CtkK2tztUgxE2XGhta
+n9YesDm/NmQ975XEcaMVHIUIFyn+mZzRf3qPaXjEfxgBwhjzQPsavs16oO+HZF4BKFkIRZi2dVM
wwohveOOCmcOVJ6DgcTYwW1e9/u2EIwDcSy/p1Y/MB3+CKvOKcullXTT6BZCtbSb+n6+faHwyYXh
S4C/CetP2nCyrHtBdrzGEggYG0oDsgN/4NzI3lBIdediOFVXrdBwz+zHp164OBbSOdL8d2T0g/M5
/6dc78Q7O1H3AqL/JWeJYEU8suUpVYTef6SPJvd9GYZyFxmGO6bQJDUOUBcnhrwCC9IOYGtnXmkx
siB21bZ03MKeZ9ljN/sKUqL9qGGslgeF/LcM3OWjjrB3mEiEnC2fhKy5jjHULQ4VzK9d8CGzWZAT
n3TPTQ4rxZGS7Wz950qAQsre0zDB2cMQ3cZF8bS2uJdMrEzYliWW7LLmuvPCZvFrr8FeIy8UQvTp
4tqCGtIAJz0FJoIW9QzsnO4NItrpYOksGklbbg5Wi69g8HRghEOPsEU7B46OLSSODrMsa9OPfvMz
DbVybBm7w85mEOfZ0P5StFe5i4aYqIrO3AA7MxO0xE3gZi3Il+C+OasweORRdK5HinH8XddvEHsP
Bk9i4RRM5Q6yUzwKqrgKsokvYF9VNKXMoFaLs8nXqQWzf0rmpyIkq6rQRA8F+J2LFdHuD3l7C1l5
sDL6SHnk1iAUwRwu4J1QDz0ec9enO1SMp492DFAFsvOUYpqOivjDaakiHJFVc442NZxqFu7Ajkra
Wy7ntnvAG4LD0I9CeegrGOi+p5yXDukP4M2IfdHd1SGKdC3ki27XLRSY3uqiOsDlXxkVKCeX/zrH
AWR4KexmrQwvf7uypiO+ALEG9ZQ5iaR+ds8kMwhP13z88SvNXOQU95mOPiRIQLBO2ienU7gFQi8G
RgkjAuz1QEpY2GHlttqbo5Gj45Ud8g3oFUmXDvlto3913YGM7cNRjUz+dh/VErXyXAcOiellVDxl
CEe+chmCxiW7yQOkY3Fw5TBd9dkRpHHB4Ld0M7wGm2kv52oDHOC5bUqh1fvz1ZAEFuckXXd0v5jD
4AJr+pMES3MLaq4BPF4j4US94mvhOYqg8BlspHhfP8fPPjW7kfwluKWLf3OOdcgL1COs1gK39B/g
HDLopl/KWD5QQ+VaCGIxB7IMzdvY0gI2P73zw2aD/1yzJaQ/UtFr1C8Gco5w11ZWDTSnQMSdzX/b
4O6scqfhzILIiDZ+wkKCqjBRCfR1im8ju6e3ppa+XpWHqUCqT/frRMhNuFITy+EtdvoAhkZ4wurp
wEvDR44zstM/pr3PGMST+RMMwJcNK0d0Op1VtTe2oPN600p44NtPI7dLHZJ81/COl1OaEHW3NN9u
He6Ta8D4+y2TJPD26FHEUFIJ0QW+p+hLQV1ErRXpsHiN+QjBg0VbdAfwL7nD7B08hspr4bjr9mOL
kM/1R/dlJILr3HSOleHoczq2boBzew/fVSgxMXyDlYd7cBgETmKHvOEbqkcP2QwmpEoWh69fisw4
Yn+5iahlTfRsJ47fE6NhjXrP4QSabZTjV5IskdGpPGlbM+pUgRxVuyaeW0O3m7NUyPkbh0/yz+ny
LTBmPq8qqCydmiLPC6ZeAubNe/UAs2BTwI57FSdm7q1phx/xxsqucEX3CvheTMhHqwbGgYz96t87
2VqRJ6WFSMXrIM0O3ZtHnSbB3D+ocFBa9j6iTVWV+Nd6QtAFh+4DZeHuC9oAO98UZPII3A6TdqYx
kFC+OqmtvDIPWqchrIY3GcE6fNw6zS8zkRdmvRfvJPsFopzKubGlKQrpo4XerJ3yoEFruiH7HUUc
mBxW3sTLL0kVIjIiHa6G4t4gMaa7Hr1CzqaFP1hY+XpYu2jXSO3JbRZDB6QiU2q2CG7Yv5mqxMen
lK8snn9spfUErXqaPXMUnIbx3IcDDIHxPSsimMjBOk+l0KWDyMHdbSDQXVSm7hSbza+8Az/YxnLw
+cI0gJTk0orHseHLZiJIrVjGQd/x7K8hZqVFW2XNmyDYvSpg4rE/Cyh6ANkdbD5NLp32XwZYYK8X
gjn8ooHwiZJGrVRCZFjrhc0aOicNhuv22YULw3jyvqp3hPRrME3yyjYqUanaO/iJ4kbR7ZbzOHjl
2NGgCCs1KyvXooXKUfe2vFJGlpfQBKZCEBCtCWM9S6ETNStx4ghrkp0pQEcbV28HaYWU0p+d0nqH
dmhGlR9L2pxxgZM0/SZ5+cDOv4u7SkpeiyhIRMlgGncyCHM93uBsp6mbnfEWR6OyYZDitsOH/gz6
ON4hFX7siMvWQ+DIt0JcUxcAAj57OrmbZreAenCw2EZpQit1s0741akirzKOjPcwq/k6FdrMbQ1j
XrEQh+TUmviNtwaVpnniBjw/ptWIPdhSdmGiiNPOTZPX9oghX4eZneWXB3m2vMi9TB7yhfKj68IE
uf4TJPXoqvYy1LRavuUqR7pwicuWWfMYygon/EKrf8H00R7AfAo3wZRAVw+C//8WrvYa9Zhh4Q6o
EmYgEZxSrLMmpMYYYqsHrsqZYVJLJ47nhWgqtex9q+MrezVofPyVBMPGj1kQpPLIFaHd46M8+C8B
zPWzlGrnf8o8kDDpRNg3D7IhQGfMYKMEz9TsroijY9C/7cEioQSHzxIxHZufk678PtbO+pQuQhfA
fhoYXMvyxiw/hi1p4ZZXFPP1ud3SnW9KCRzdDiI0CN2b+Y/2qJhPaQ33WxGZbKQLQXLAQypo1CoE
4AmCLyUByAcYIgCjTT+zXAQU12iwIZaxJaBlj3xc1IQa/YP77RlZjfP8jEF7Grl79mlmxhE84iMO
zHbCS1KE/P7UyXqyNMq2oarnO4VguxNRSSxe8cmuh7TWj8DPI0JF+1h3I+CAhn/t3X04XlhjIDtc
VZj2ihK7UXy66cQe4ctwhiX2eUWrCc56daVqJoNfxnvuD3jjC4y/8NIESJSYVVRzu+mpZH0xx2aW
x2++WV5imUt1IiZvTP+JN1452lgJApIFkVfk0MjeaScKeqIemQaszW+TwE5CBQ9R4cS/nRBV1x71
Kbh9UKEcSXQWEm3ZjZv0nqPWdeBRVhO1hD3nJO+XIuY6Ovrw9I6p7wfa0ZLp/DfsiFQfx9GtW+Df
9Ccn6uVUmG8TtKGYYLJ3pJqCf3ERNGhsVnnQyC83mz8zF1wWdHJhPNXv9i6xfLjA7WLnnBgnTGOA
OWEQPf7US9zW1jKXMziyjE2MIxdF1vBnw+3EBY0moVJtID3epR4aekgaK3BvJgpq9PCRgjLUYR7i
dg615QuZU+4LamrU2zKoHwi4Kimju9gZUXmNRyyFF7gzZvcR7xuaVCNxtAInjmECdq+2NrKriL8J
0V60QLNNcOBnxEP85bG/fcbPCPDpuARbgc7Wkm9DZmrL33f6CfFXbQPU2RA94ulyT7JvLkGYV880
td+ty+SI6PvX0UjB2xsXW2fuMrRTIeIsH35loW4X3mqQYzZD16rWpUEIVbcShJpga/djfVRAHXfB
lGrLJvXfeHR9i/1T6BTOvGiQCuVt6YDrTgDSe1kJLmf9+UWOlABb8L60NsV9GBzqe3zuqiujC1E8
vfl63VMYoYorBSXx7Lq+lDQs2MxY9TRnbXEAOLzBBtZe1nOgKCabrBo6R8dLgCNoPni7KrTUG2KB
+N5GbxAEQoHRlPoE5LK9ejALDJBttwetAlLk+/KygRBNgUzfC4B0IKNpNXZ9GjCWEbAVKlX3QaUu
3/i14sI75gMA/QA9KOTMGkZ1np7b9LoqoO7Oo5TDklH0z4BM45etq7eeVERynOjyMqkHEyfhFHpt
03F23MA5iL5PI7Xyil7lacKYKtX1aigNZv9rnzmUDfqojXaqhlNT8OXm+hHorCaUMd752rRGdmKG
dWP4s9pqjMgQpQL8OFhnFo5tFtXWzJr/kPZQzJDdI6vu7bKrCmL6csSze3zP+quz6pQfSBRMHCTi
KIno6OdHQm9QCI0qq+Bt4RlBA9XiS+73bTNq9oM9IJLKRohYdh94ctCvPz5ocoutCcQ2vNpsIRao
Kld3Ly0vKYFa/LlrYotZNM7C54uqoeCQqwE7HhpFvzrIKIzgvhDkgDEcFV4kjlG9rc7w6gk2rvCl
v6wh+OCHObF4udBBsdeNDc8qqXT4+e1R9GPdPJaoVf2/UnsAb0wdHVdXykWIsb20nFyGmBHWwGsK
A+MEcHaYVFh+Lh3WKLDR3Si7n7JVkYn3Z9zw4820mMaJW7crM50OJ+DA0+WaVKyz75gE1btTR+KQ
r8vENDzQBBiU5ScXaereuOxhd/zFCm1uxNjyqpAv222NySJ/FM5kZ7+LX+SIS88WXmQukcJCuNzr
Ydy0GDN+PEc1A7LQa3R/NU7VSUfecMnWdThIYXNOpORLI+uIQVOHRWLJknCnMBGB1ZBrC24TVrxh
SPk3KeU8GdWZknXi4IopEMoDWuO6eezItwWpSn0XqBSt8/uN6uDoSO9aYiQNgCfru6X1fP7N+NQh
VL9PiV+/jcYLX/uS1R5HzbSmUoOETqe6TzDGesFQ04ADNbyi9N0Kb8ep/9DGuRD89S5Tp6cwbxY9
6HNjgVKZB86dBX8FRNRcPvwXun60eIFKhhFpkErmRI4S6QZX6M/Bdd08uySkZOmCWEa0txVQHJss
BsWKj26appzVpVncZmL+2AHcvtaLXJFGNIVxGXEqZCmoNUNtR3pgPF+j4dGFCGgJNFl05afUritL
T8at674qPYk9RliuxYAVszWnXRLaptZt+Jv9yYGDqRp+EJaK6CdJ5/1G4+ty0oKMlvwT86w6WXdD
nK4Cwnk5XK0sXL1sPzCn6zoAiUUkmZjWbhGWvoo9hramRZkjJjU5nVTKIedZh+Czazvzf6oZNGni
vhRA+eemtiMzhjt8NzQJssCVPiPHt/QxsmRuTYD6bGtDYU7f2pM8tyJpU5B0Bd9O22Qq+b+nBhYp
qn0e0RdAlGWpWuPV0x+nDk2CO4Pe+9amVwbP8c/9y8+diBRPt3RbR2DouNUFjerdeKlETmul1PHH
Vqhz9Hk7KLP4sbUKuKGZljlW5ZssZtxhRjrBec0Uj73inYfF8ny2nmvWsxnJ6cojHeTnvS4gk78z
uCU+mtSoRzsl8RlnHyVwPqqWMjn3SrmFEERGEtbdo3gOZ7nxfhdiqfL0wckvtHg+BMZJG9emmUhF
5AvUkliGEbqHkFiTqbDbWuQ8EuwnzhpGhMabXq/yEK/bf4EU5jAssYs1AZ758mOTd4LcnEumtPbW
TrJzbx+nnnDbqfUOH2Jb8BUj1cR2gSwsHw0fyv94PkUjKTa/By22FW5Bu5vkBSIiSVlsvHRajZov
J3X+k4xk45eUvnUmB7EwKm99f5fkakDi4mZQnZ4/5VUPQcERLdP1pFkSo8hjAratDmO9ioie5fyo
4phLJ3kkA0fXM7OLppg1ApQXzez483AqqA4S4KWY0/wm+w37MdXgtD0irbWe5WwFjrmzPGrpm83S
LY++I+DWek0ri4S5BNB9ddfJwfpAsm5nREkLkRbiwQ5j7NP61Me59S3LRK9J8rMEY6/mkBkglyd2
lV8FwLNLns7k9bsNl4iRxAiBpYPGPCjaXBN0175RTPpvAXtNxauJOgjt5QgoLHrHMp7xuMAD6Zpa
v2IxaIkKeivtZiWtet56iTZCibfywwvykbAIOuDA/02mKJ9NVJd2ljZuPmmmTuOtVUReIMjeKEqr
YZdeDughHsz1vmO4KFRYExpyPgRWABaZqxSJsaMGokgK0x+YppQgODONU+NLKQEQ7u1PuQ6SaIDQ
3+x886FjTlV7b+4X9r8+HDdlNuqGYOJgP3+D3ewze0lwjNplJT+4HO5wVOs9ybJqdc++JsAeEeSt
pKCXv6VBAgFtynTAwS+bv06JqaQTkMe9Jww0L66ZYgl6SGopUYJ4uTXJ3B2wyTLdnXjuJMXGHw05
ZSVDnYuyHhn9liZwsisgAMcys4V62zKbIkAtbjSdzz50VGvPFVjf6b23lue1AsLaqgsE8GhTZqSQ
xCHAdZkQH4ANvdASm3vL69Gty6xh0E4sptrpcSUB+2AXDLQnCYsyPcl7qZlhPYTisz7tFJxgJcaT
iMs/9t21Eoweh5tAgmDy6iuyLaG5vCBJTnk65B/hyDnBJKWjCXpiF87Z0MRV3C71bDWFTfo+PJzC
Dw2+w6kaDH2BcCjAGDU8WLugUaKdabxZkvMcARokrp/zNjhoGA+gAxx3nhQJI0VH1ui/lXkWfLgV
zqFN0FEMyLcihufecdtE5Q5hueUC+2o+ox7Y+t6LF3ekVBipcXh/GGkLLMkEk+U8MMsmyi8hZHhJ
wAxEepF4OG41Z0KMxR7s3dxJCWHDFy1hzlZwsnPWbBnbDbu0vEKslTkReHOln0zc2KieIGmKJFXY
edNXK2o0xx0EPPGMir2WRs866pBxRIT01k08wiRu9kYTBA4Lt2miH/koPQF0PORSPzz8Dg6cbFt+
QbH++7DUfN3NTa9uIQrnSahqAELugYYwSFsho6RgEag5lojZpJTTvQA3nnMBsbQw2XZt9KwBbXFY
qFHZS853PKFG4nYqVkefD2dxvC0BienhkeKiJdnA1frBa0+QGSJjN925lZB4INZXBYTUQYDmdEIs
oW4EdG+88c53dCKEqT3KAqHaOc5MKT7eE7KAp0WY1MX/TWIknAYGp4VubYq85WPy9cjpeOmJh+Nv
pZm/2LG9/6WMT8Jyumla5dXoJGB8jeiI11LIubPDosfGrDC3pSGeUO7UgRnt9tOec5i6j6Sz/pNg
PTm6rPz4+2LmrGZTu5ksp8oXeAFW8M4Ov/0XRM5FVMGed5Z+5dWU8mgTDsAjT21dQsnOMMBqVb+a
ZCEeptL8VV65636TT9FKYvCgHxmUppGIEL441B1AueiCUcdqBvrNfJumh3GMJuInKR36n7i7WsMU
OewtMaCgW6ft2UWrnTQkTh33FzdIKGGkK+aIjHGRceOYgsy/xRGgCbTtyLvtTbdBfyTFjLZMNAGK
LXo0zCod6u/a71ts0tXrTLnbgPoflnLRfHjQdZS1J1FlldARa3PqX3E5xkbFtPTT7HgBnTdBdlZR
GvolzQjEjmt0tsT9hED3JDvJOaNYSGatIPa1wPgfVmOky9hlJYE7d9a/RYlQTGvyp5ZTDDAWvM4z
Dc1V+d5KDFylEcDs54iQa0p3BoFgNhY6Dd33DwnWADW9foz2jvZIiL9DNvrz6wjaEdwwe/iF0Id7
TfahfNwl20tBcPs+eesYEwCiuWH/OCcK43QwIqwhqiNMxV63NIhnp0eCCL52Se5bGXv5rV8fj67q
4pnq9a5oHx/YyZY/kf1dAabmDSnEbYRS5pkG+zA6O296jc8FkqFrisOMwEEKWVKnfhND8nWcnoBM
JGHWjd5jBD4hjRGL9n2eXAz40ygmnWjjVIpXUgKp5xbw2T9QhsfdpYo1bK2g6in7jVzfW3Rg0OQW
pTRSMuagl8n9an2+PzuPSGcRv7EZtbNZK1jdaGWK39pBwVnWHdTSKoefK9SOk499BAoZL12Mq1B+
WLRSyWXnI68ooENUsNxxlYOxPF+D137DqLAnZXbk4eczPi+jFRIxY2MiQ65bJAvbkuZe3pGJxpuL
9wfbtcJWfu/19y9RoJToV5fyOSsNtkMB/pfvk9P6UPCf5xApT+dLXg/hVXdxn/RzwuLcjCDg2TDm
LKYadukGWhivLCCvnktsk78TjG/oPZkHqEaLxRw7ege5x0y//LArZUskhjvLcokETmSJdAZafWnw
E6dOerSv20Z4k2f3HHVrmsrXKRe+DtUl9YquYGFuftbsEDkNTQlZRsf5Fdu+58vZuTGdLlbQvcw9
jKjpz6pCQIfiazQi1ojW1ueAW0hJNdNx/4ME6w8nn57jWf35PZj0RWoQPkMfcI1+orCxrkGs8sn4
rbhopBhBswAu2NgXzZAiKCdo8GivPWWqIecdrrHw6n4FQ5RGC4W0DGxuc/7VMS6s9vXW58K/MwQh
v2CON4RPx6yCsHpchRJHirJvCz9aITnL8CSaOhReyfFPrJHeiGgSLLfwgMQE3weeTZIADeZqXOts
DUZodJfKS5qeSHDHDbAvRHSKjqakXcu1gytjGD7WBqFtRGQlnybTAsrTy9KYDSfe4WY4bWemxg7s
BK3Q2RAfIWd7fRHL/U6c0SKs76kyJUqz1UP9y8AytalAYERWjRwbgt0ab/+t/2S0+pxvcQCH6nYC
iegk2ROYlyMgFflPo94flJ/VFuKd33isGNcE/5wO6TmVeOaH7ch9kgXsM+p8Si7jXR+guxeDFQ9F
PAq/M87JjW5CkHq0eOgRTd63yZKpwqz1k7pQTrkooBsSlIH+C4p29NldPcnvMdw8vruBC8PrCBAV
HpzpNCFQufBcaLsrT0rQelDzLzaFnzygRBatsiwe1zGIpovvC0jOrkcFLqOZXPswbWHOpGFUCl00
T+nqpHE8b3iUPYfkHUBMrZpnK/34+WPSSc/+WwF0tFKTgmJAIUHX51h9kKfyX3BhXHcJ0okulGlj
ed+tlqgW3lRP2xtjy0rLUoj2hEI7FOKo8Tk7uWdkJ9GVzpXYYBEQ/MZLbMVvCrm3zu4Qs4v2jvIm
qKJAz0iVvbDFJWEe2mkCS2a4EymwcfTa1Fc2se6KJMWhuQt7zhGSUFpsPIZZa9n2solieFql5z/P
eT8wLo+jYVKaedUpoH1/g7Bm+m2Vebr4zdn60msvXUGPbuf7mU2NVWOQepteeCERFRgOJHg5Xe7j
zzJJDlrAYtbL/fHcEzoetscI1IBwOpiR52/zxIkToTip5Pu/TG+uctuy2u2q33DjzsDHXAt68KQb
RBZTctTHPnEJ9RQ3/J2S+F7Xg7V9sJWvlcJTU6LnjD2/uENgmP6+BzyUYPTttndYKGIZaGIryJVO
BvUUndGLcfk3VkJw47dkDRD9aMdrePhi59phU+khLqHGq5ParUdHzSWvzyR1OlOi46jM/aucMhMk
nhq1Q4jmu5StICKD5hxiBjnNI2yQso/wsTZDYQcYWvZvlSoDaxcyYcMb+8YZXWZfFL62DSevUFtd
EapCX75/qkB80+YY2YHnLiVk39XRbLJDaTo0n1Uf1JglkATiPF0LW0AKsGRUa5syx9aySsmWyuZj
ch7iaP9RB2uuUfU0LsyQjQMWMm8INGYRH7W+uzw7sUcYj0njIbiTaG56Ja4CCX44UjGeL3Kk4pJa
12xNpCadM47XezFKuUHA5NQPmyHF6Pilie6JVRZsb2+hm1hKBW53TdxZgm5gJ9MVRx9aqvsL6rtf
etUnmyj+G8WnBa+sdXjS0G2gklnIatcr8G1BAe2satht9wHqSSL5ILOB7jIHDVeKevrUY0T/aGri
RtQTWp1manLc3o2tRfQsZS4BmdunT8ZHvx2uCIWKse08cYu2MDDnjbpdowggA01XmqDyPIO26SvO
gngxzZrZJOBLYUdM4I1ujegghXqf+kJLwqipaToQI7NCXzUsTdAdkGXeM8OPQu/t9OXsvuK3dTrx
KBy2EblP4cvc+8LOWokegUp4o/D2I8iIDez9GBxxocqigx43aP6ndMOk65WARPhoKSAOUnN+820K
f7o1tmpoXCgYIQKdGAOnNHvKgel8GD3lZo7bhjSY0WgCF4g4e2HmzBiyzLy4ZYSoKkBGBk2TpvbX
cHOV2yOzZas2ZL+92+8NBwTSGLcF2JTGTUox/E/EkY+PxgtMicbUTYQKcU+L9gbEaxvuWnn/lDUu
GvERoNnjBARWQo+1v8ixfJ/9M+xO5qINx+rwiZiTyTu7r36EVZlIgq4v2rrpQKjFxm3veWKkTHK1
+NB1+Fm2dWGzEKTvJXl1kGI3QEI+Jftc13e7hLlgOyHjVSU2xLzs1Ur+rBZVzqbhu1N1M3mzuTLH
RGbgF17QJEv9Q41Uap4I6eP8Wv9E2Z9ZQa0Apfbfnh/FMrTDzo1H1y+aYVU44dzvmZeZFbLGcmp4
+be1U6qiaFLBwoqbON+gj5EZXo/VY5GmmRAQum2SZcSO8HDvBdvjNcki3eB8ivDbMhPH6+EOvNON
w2jS6zjpRaBfofxRoydY7jexEafUCUmJFzc8LZMzJZT8GhjSDF2FtsSb/yjx8ni4PanLUC/vDkD9
HxX+8OiCnyFJ6rllhR3Prj/nVZ2yu6mkxnMMPBjCtTSFV861VKLecmyRpENQUzyQJjqF8nxX/hOz
PqNpYGSNzHvX1tWCvacHSnWkDoSliA94crWW9gn8aW1iusEFTGhwzK6hPirBmRj2YaJh4n/4Zg3t
7Fc2oz9ctofcbmKIlL/wl9BEw4yXSsum1ookIHRQ0kUMlmwy7ER7xENK7tSCEKA1Ml2yfHT25k9/
tXM6hTdkn954yKtYNOzGN18w42zieYud8dKluiH1zG/k0sAyDTer1nl273j475VtecmUeN7xkPjv
BBxc6rQaeXw17uVjzxcE1rsMvxj2/472BJ98eCEBvBa8uX2SrPgiUARyJUcFi098Mtm404cXBcT5
Io9Y/oMZID9svh5WK81oNqEMCT2VVUOKTjubcyYZmxZ1ZQvC2r47OqKwq8t8MIq5N+LKOWrKoqt4
9MF/tGeq+BOhlCIOmpZrwxi5bu2+Vpd3ADM39KzDoBgtLvMvop2VaImlc4dg1wmeigBNnhEbow7q
Y4sfhM7Zwa9Vxrqc3laHj2A38LwFx9fOY3JmVUS5QETskVcCeay/7e8Ttnldyx29dtRrVddvNteB
96NCaWo4ym3rEhsrrV1dHu+y0ajU0vjCsgzGxTUoSYVaQgEjoMMN0mtd2NoV+cA3y1JjpD0Jv3qV
Y8DZ45YQjZvZQfU2y0MY9VL/xyt8hDfq2Amyd6dGIM+XrUlOzocn+a7AAa+4l706GYS45UguCbFL
r8KF1QvEH5w5FiIYoWfM8N0Dx570lvFU1PEqAeuRNTfOFBuD4Y6D+Rg/lhpNKdKTxgPTEBcz8gMj
7Y6VYVECtW+JFHoR+JboukqRhVFpMeCfIy8LFCskwUPOsCFeLQ9hKdZsToaWhnqA6wbEzodbXIGB
Y5LQMPr5uFax7Od8s1v4cgSgQQ507cwZz13dPoE4L8zzMsPRNKAnPuE87upkyZ74iEN731TbXvgO
VvQVqkxd71OFcDzpGHVYPe2h1GWNCChMSYrK/aIFhIPYuG757F0gyCxQ8Q62ZyTXhRl09GI14GRd
3MYqBlhZNbXmlU5+YMEtXoAxQhmHzYUmM+izhNFGEyAzkynEpkiT8oyZIJ6+H50hxMR6ISM1aVfl
ojqGaVPc4mBQJT/5t4QZ8eWXp4JgOVPUBGs8WS923R022Y3f3WpYLuJBi5i/rkLj5URjnu/G7KKf
T5+s9utdpm3YgdSZNhIhxT5WqGwjvFTJs6zJXWCV7IXkXx8gAR2g/a4++0kwxzXknmITYS154OUh
omokdSwNiKVbKedGF2dOWFrXyf288+PYuR0f03AgijVF4rG6CunNTdSNvVAGERz5FBakQqW1x9Jh
TrWxsgdMrm1Qo0l0nj6ewryTGImL30Dexw4rzuCMTNHoPsbQobQQObI8aty1G/aXGE4IXV5HkVYM
/0dQep91bFO8BxA/rP5IZ6ywOgxuDA6Nu+FvhrZrA46go9thXos2ooiYwfhiajPZP322CaWhEQ+O
JfgeI5pFKbOHIcRXZYjH83pyukf7lRa3r14+TYnIY/MaQKtrLNBtYJOjQ/A/a+zYqwV3wHMkc7aR
kaRA1CiNzlkuo9iYiNsj7y6NKVe5Tq3hcbTGoReaatCeLXHKPcgqv+xYx46lZzaV6D2eoLQ/aRK/
3PN6JEiwAqTH8HMFDUvnSeTAlb1zgJWKLzCsxPI0ScnBPRGvoD/C0iJTybZLl3MMhZX7GSmMIAJ2
dJr8rXZ5X/BeHixxpzuMQBTQKcedTmThplQopkLwq5LRborD/X/1G0BO3u+APIkl9YSy7izNM8hr
zDeSx0qX3D3JC3eNjIO2uSkfoeEMni3wKUE3uzGd41IIrg4rl+dFr9H7YW1SnOOiXarJyB37f2qC
1WdHLe89Mnc/6nFWi8DOQKwGHoWwPRYmUiJxB7ey3voMR9/2qyaeWUejJWkRsdprTjOMYhILFNeI
FYBe9jvhHiofyi/4+rTHcXl9gxeo1ofpgyM/p2ErzOpWeRwvRmsPH3L2oz6FEaOPjyKgVJgUCSih
LcWHx3Y2Bum0gbDYNeicCVCytSwropD72qUfy6JArYKABzvr4TUu7k6TjvMQcS4OpxSxjssmt+MA
pZEEAFKWxC9elx65JGteAlllf1qzlk9WejhMw9EAmt25cqrWfYwHMexGkEl66c2+1O7MtSM8Sp8Y
nKJfauvoR+bJrPkG/XtKY3uDoq7AkrJZj7UmAp3pP6DO4HXI0bYizE19o5MjXDrjDtnuSn7BbBO7
xAZficvcxI4FtEvMfNPWv870wuvwBpT1elVx2mTmUWNZ7RgJ2ubYTgDC6F9K9CzrAVWXow/9U7y+
RICZHB57AKx3a+2IsjQcUJYlraGER6+0UBygXrWPZt16Y7+xh+WvbgcWazK5aM3Nu2SScmG1JCpR
KQ2nzWIkKbTJSzRGbzcFLo7Jq5rmgChL+VJJD1POmIoQ8ep1mpMTppX1doyDrNMWPnXZi6TDbHX8
xUSRNWR/kYDonL62kuvUbUv0MwJP/7wCVKXrRntlntRdItme/WxHnrRk8UVp+N8SQLvKLbFDstoc
TTjCbzmi4SqUVNFUFER8jlmf6Md3mlIPCmqMgA13KkgDu0eYV7xLH1a1bp1e8eW1ZHD1GwBSVOjq
A4RNvsMByg5ml5vF8tNdPdAiPD/YUjIOpP0uWznqSSdnJUpbE2HN82/8uBiQ50bxgRmsGOMj3ahy
yeEVDbCAJKJ9ntmAe3UkgYWAWHDD0ORwnpwL3biJohZSp8j85JmAHJbgAznpqxzCJrTX1okO+AvW
f9RKEv1bY4/GlDOFQ5+qPFDE0O9QbuqWoO8RpaYFikay3kI13V9OwWOprrLWOzzKC9+tVNm4w/WK
W1ljqHh0hXEHiTWf64z9LKkeTj7L9SgQqj3Bsd91jm5Q6+1pYmg12YtTq2rbRJb0suBbx9zjKyCE
AuwprYKYpOvMEfadtcRm1QV0+l86yL9P+hlyCVcL/XkQFq53LcXb2ib2GCxejZCmXxz0JnO+JcQ6
qMtJ/4O9h4HyIBeyImkRhKt6QdS1TiJtQ7bvocs28/VR+lsyjbczdIsq0u8IxiXmHE4h7HJVxrR5
h95dGRXF41AKXjOFM4D1cxBhQKQvuzcsl1IawbjqosePgi9WTvcEvqgZWLLZ3a9f6rDsspqwHm9P
o6sAUd7EinVamnAfU3lOC1rHHh3Id2yUphJcl3HDQrRgUzWsNcUmEIB9I8wAifhabEwPJnsBeDe0
tLC/Q1JoVIsF4aO30Q9Q95LRkUrZ/o7ETyY3CyEJcI1DsROBxDN45TavVsfF5IWrhnkEhlPD43DO
0PuO5gM8JBKlarCioL6fyFOUx19r9tDkA7It1kh5DviX4Dv5fBRGfWgsdTE1QMxlXI8KhxU/q8We
AHlZszwnyR8gQqLnb9a1rBAJWQarqGGdfGG8kr5Qbtgc3UJFxBXKtiihnxjyaArqN+GpCaeTsVbg
fFCXAceOasg7mHYaM2wsGJS6yRKbeNiNuRJcoEZl2Xiw1UTZV7oFss9k7qCBNcKUJcgDD3KwMdSl
4KBIKoCzlWPM1hcwKajcY3+7fuYJ9bBNNc2IoYft2F+zC1xOp4uPlHt9bCFV4XtfP1U2csPp2U4A
ncrK6cL65NTuRSvecU1V0k/IB+miX5fXVhl8YAiLfch1c6XtCvIb6DCR605qjD+1frw0lZ9VYs4+
pVEAbp8bGBtQM2pwNn9kChf4lgC9scbw812oIJUUlyn2kjIKnFd3D2AKr1RsjZNC7kIhatG4AGI8
zVMdi8vUOa5OG9830WqNCUgqElI96XSNXYX19SerIkDFIvnNydKXqs/9NV0lVIL3ID69S6ubiIDl
sfQXJD4NB60ByY41ghCFyvYPSeIOD4nyqxoeov3L+t7BuTp/NZnParbc0DDHZpesKQX0/upFH6Od
D4YizbxnKGg6prgrBv2ASHw+10h19A45YDp2X3SUOi0j8c8wag2FmWW9kbFOxVaWDZUmk+5t1Y18
cGV6xFYUwpdLvSXfg+h/G8HNIAwiAH05Y8wJUDKZaT2smRTq4fOJ7glSZnqPI+gMwb7624kFa08r
lA/FWapjbDXO+cHblfZYPXzcxa7ssbC6OiBrIUv0mJeoCi1tL04bn1WrHo0mKVWOkalYV2vMV7am
pFNrfn6BFx3LaYq4NHpWy4JK0REimSUWL0McU/1alyaXZAfK6iufvzcXIX7pDCL4rA43LehgBr26
uzQwB8ofEQC1uFjTlg1jp7DXIqFTbUjGpeB39MTcAEQPORNwdDepTr3pk+qZ3+vcWPgGIrUlcos4
2IkEVR70RMVmZPUPFClqy6N2e+w6CNOC+l0j5bV4En+OHSYtz4QmVlt2kutI1tgY5GpWna/KExYN
J30aAZAFd6m6Blhl12lC6eUJmeydg/lE0ITEP4Skv/sXM+DI+486OVM7g7X+VFEbLJXimHzledGD
37R6OT4gGB9wf1iK1M5b5JqP+a8ommv67B4+LMDhxBLQ7cyM35wSn5IwTvH1CVuH7FwfM62JgDHR
iuytpA7RShk997oPzCJITGBnvPzTJ85c5WBapE1NdrqgMem5EWDZgVmlZCR4C1bOAZQUU1SS4nzF
mTYEG0VvIwegbT1PIAmKWDEKFfMFyUlUPVbI9kwKmkE2Dj7WPOo4RLqcuIfz69X3erPBg6jURzhz
d5+P6udkyw4n1vRxh4rNYEUm1aG3Zfbs4hhJ6a3utzmKEaY7J8xdoKkat8Uzx5yF8NKvFBQm7uCh
JsZ/9k6SjNDmId4OFX5hxVeCYNpp7g8X50J2uJxRul1daIZc6NebpqbBmLoiOA50u7rNx1oNo5C6
Qp73HeU84E1f3VCyZtgfM5iMvF7rX+G4N/11lxmtX63OTosD+RspoRQcuBG/RihzFKVhUWG6LKMl
iFLe3irNuklkkrk1VxDoWXW/1WgrwOxY56lBFjukRJLMXOpDMwqbc8GqM9gangKJkcaHdsv1RWJa
sJAHwL8dGOfMy7bexUfdnUWl8JjFhJxK0IKnKrQgRUL433Kh2hdU3dEBecrP5x7A3qFqbfZx/i5D
WqnCkJRscXQSfwFPfNS9cGqw4eGJmPxVVw6XLTPy/O6IHo8rPGfBuDhWEWYUz67Mh06iNhEYIBCS
XVxVtt5kn4g+q1RzGEUgnB/w1+MRFOZ5IlltM9FzHOvFd7v8GJNzUHdlf/s5rlIJJBpm3mvoPhqz
Ovx8OZAsdWWkWdAm8d55V1AUkBK1ay/2aorLK5Wb+wHRX8q8lfkU91q5r3wu7mrbIkdqlXaluLYQ
0y2zD4ZuJTPXZgKP6Kjn2IeuiXK4SFr8S4VBnm1gZzknCTw8y8zX9gqhu6wZwDd1xqodKGdYbLtM
jRopK63NfJInMpT8DABDaWDOAbEcKoR7KtnvAe/8eyEVRqJ8zideXENbbKIKk6KeCgGXKpBHcuV5
CCBQH9GIml7pXdZyb/dNgtcwTw3HFLs4xRA+jH5nuS2wglr/T+XIGzIsSGvDyDQpcjf59tILa6Hb
Dd2TChDF15TddfJ0YU4oMfRIW2Pea5H5imupfEetI2fRaIUvXF9NE6Xjq3QW20pjvJa+tsuoW1Jm
s5F0g32EWtj2DQ94/mGcaK1s3ywgHDNNiO/Ewq4HPObTlFIDwrm7DTkYrh4A9q5n5jHSgw4mgrHW
FSdT3v9u4g/Ilz0kwY+JRcLpFSeAKkgMjiHDRUY+l/+o8NVcXs1f2zRZ3sD5iEwLvqERjhz1YJ3V
PtHFCxGMUj+EymZE3gydoBqFwMzywWsNmyVKDg2mgsIkHgoJDKUZNjoA4JroxB+xYKQVUlgYbZrD
VdiB2y2sV9oUwzNRrmSSDA9ENr1ssplEKcrY64UE3iRah26HoQWoUSehXrB9qH+jsEshblH1em89
QCZWTUleMzH1pJ9OigG1KDjJ1mEzFrqqhpi5/naNI3D5KlqEPh94dU3I9jngDfmb2ogSQLZUp0RK
mXpu4/oPs1D2dQlmV+ht/ZJfqu5cs2RolCrXEaDlKeybLo4tq9DLda1YIj+xPVMbSwbBNv23IZqI
Auw8KmXaO1fYbCz/wuJURQSzNq2zwQkvJbaZ6g9m+S77aL7xIX2SyzeBNmf+yb9Spf4vYoLocsUi
nFIE72jl0D70BO7vUMGTMcDtxNxQ156llEWHaMq2wcuzTIcCWpgLLvh+N7KlaW1IkffW1mxQP+hi
P0WVtiTulBjeCEsh+hjnxCAGY2Akvi6LvNyCH7QVAkopDF4Zuj3+44QZrdyBCzjQMeBVFQg1QhmJ
pheUdI/Rdth3OlYXtKMQla76jGfRutmYsNkvngb/qlLFMiNmF65BEQgHrbPr5k9VYhSxeBXodqwj
MGILey1S8N0gC59D/giSg5M9iYROG3SdV4LAbM+valoVlGpuTYWm/MQbUUjuY+z3bbxbyAsmdnti
FMUaglR/MadZW2bbR1lomRNotnbGPgqg46bKvs5ZDqGKO7JHM/IaxMFceRxwX9rcSXWDgWySEmDt
Iw2m6mZv+uNVauJqf4G6BGEBttv+DCEq8dufAB4RU9LDLG/mL1pcp574va9n9AgITCMRB10spq3z
nPvNqfhLNUtvZU5rBsoLqSzGCMUGrr2yCDzMylfZyp2m41Y+CXlgAcFuSTxPo+O8YukP7sZjRLd7
0cq66S4nGhjJlp0WIcsbOdb/MW2ZpIJxAx8yGVFDVl1A8BKqUwoNBaAsto5oni84OSmH/TlhreeY
r3zObkc+h3kFxGmejGs+cEWH+vQbALPCudp6NQ7jO+cVC2spKABc+eTvbnhimxUAbOeH00z8AFRt
bGYOZ7P0dRP4aB0CpV/ImJ9+L1ySckyPsVQeZBh/+yE4GUlg4qQlF6MsS1yGoBlESQyXVg9Liyj9
BqyBJsrua5pNV1n+uQtzw0wM1VVp6ISKRkOLnLy7HDxTbkMs7v9cpwZROM0cJjAg4NCKKhpY/gUt
KrCzuV4qQx1pwnYf3Pn82KdoJFyq247LarAUhIAo4jXz9LFQBz7TXedJq+PSiIUKSWyf5o3gEYMY
QuNv2BQCF5nyxl37cmQqigbZh6HbRpqnHqnHpcfCMQGGE6xzE8Bol0TY0K26KatoR0ULTu1QpqbZ
UidoUSeQDqf9nQXuHMgAMV59RfVBOAZOuBqGdpeKCGZNtTgBcRKdNg52sQAFIvCfr4yQwHbNZhRj
D5OfhnXI2rI/IItor/ApRhd8n/nydRQ0Jko0jqy4/KcvqJqI2kQYtkCYgudoMs85D00kXUPAqUDz
BhLRsBH7oCv5vMjXuYH4Lmrspy+lbdIsZsWu+YvfPR411N/W1yL1l0MExjyzlCSpXlIhXoNnJS54
sPuXDwqx/MLz6FQs5YneXDrUrv5s0SLuhRSfJGX2Z/6niq9nzvzqDF0U1/0/PGLV2E9aDQ7+WbjL
iw2F+I369BF7EMTpcECqmA5mQ35CWiv8oz1KRhZRqiEALmE5SXKZfOIjcwbtbTeX8FFjR6YueVg+
hhRt95N15I1OHso5eMKqxH8tf96VHKtqCZXsTV7Ta41ot6zSju50qFmFowJlynnfHYgxdoTMxnc0
AMvU1Iy1UenDM2XnBQEp2dZ9IJfDe07JRQct5XuQrbMz5n85QwnP9HHiphEpTTAiKhnpPSoLBOH6
sYq/P/p2NF+9fPmdKOidGrTkTqwhHYhtgwioPqwLUPhDG+xeIQ/GvkOTNC5h66FcG619QAaLhuxl
Yo7+ivKX+SL+v5wBdPXPVwhji2SxZQnZG4eQMtvchLyrrxeT86Ejn7y7OX2CdHmPfbJIPRoF6Hbl
7WxRf+5MObRxIm55Ovjdw9i6O7S74ZLmny1dMKae9AqZebCktbqI6HKdE0HUj/1mnj/Vvv3pFN8w
1OvZ+5h0XfHGZSE6jdylok/wTdvW04mc9592cSxV0oac0uBYPcZyRl3abyNS52k/svEypbqRHd1h
wLMt5FdhYO82jLQGSlvxeWutWS0i9OvBESh0CGJvXZAflNbgZi36AUd8uSSWuoD9j4RZSasuAJ1M
behQoopkTsJvhFlhnYxWr6UoVx6/nIjKeCFrZgCkWhkTch7vRCNu4cDqsIhLE5mgo9sUdVua4U4u
hg91WwRpr98FPQSKU5gX2dp/OIS189qGMvAB92e8gMBPXrweJT7IoGB6NY0H2TjTpftiRFa2/uPK
F7rdUURQo8/XMye7EX5sCsT31tuiev0U8tpF91Q6atGSwEKenaywCDyPzVttgZogvD1sWx+5G7kf
N0JC139yH36nZ9v4sdlfRv6NrEm9G9o7rUc9RSXKHKgfpC+Cg8C88wZtoX+Z5GwIF9eNYSL/K6fJ
dqG1ljf44se8P+UyaVyeYCu9g20bkt9q2cwksQkpVjD8Cv7xZVpD1rXJhKVwDE760V+1UIhZGNE8
HHxas1q9R7E7q7wJaYody2xoxFL4nSw2gjsvskYjvz9zEBYSvA6rJhVXUsrC4YvRUfDFH5HgAWPb
/3EhTm5WfKGMyovVY3B11QCiemIOf5fCd1c2LMIAcYFlP4ggSAyFEqbEHAlYKOcOHih4Aq6YQ0QH
YegBMRSUH9GHOgATRLWpCjdAtkweWLSeek5Wyc2lxZekXAMPty1n2b0dAU3PpxVsxw6hfhMHjFmB
pISwHQ0GLKXRtqrWInI22dQuPeAQ1fZYOms2tdm0Xi1wEvElYpoI43sMvDJltv3rNPFukSHCQlYn
Vj4lYYwwtCSVBULz6VJm7fWCyDl8dc6ChC7uHmkxrtAT0tr6lAVlP961yZ1Mc7awA/wWgz9ih/yC
SPV9rwQ+wNdbanYYa+gqGfsNw7IYxE5gbI+iqSwIsix79HtWcCtr7973+USPuJB5HCKm58YFFS20
xSAepqMu63/wsHd47daGqLuMkR4XNNgTiOjnTmI2dWGQzXFHlmmKOzkObzyIImQ9Cl7YPCkdIQ6L
BrZF3B1IgtWFvnIWbb59X3NIJRB7zWGqdyUG5D3SHpSpmOFVUluCHfN3ooOI6kIGI0bMO20tbjeM
yhSr04lw7FpA1Ej7fjF1wgTvSmNg9jxoYSo44fs1CIKN90lqePdxMbKjwE46yy27LmhJSyBzg2/W
04l+omHxpLsJIuzBNLIrF3myE4yeYX8x7dOM2YKr+4LqiUXtzqmM2hSuEle1TrNsghUqv0Peuyct
tUFqxdOqEwm3pE2foFaZSsEuCaFeZn/QvPiJM0WQ2FAqsmNPi7VXDu+LQwSegxaH5kDzMT4/3Fa5
qOTlvrbXLxzTzbYEjx7T+vsClGD/3VE4K4zIiAzqN8EmTBNi9Ph/wLnu2IWDP4rLCGlUCxp0uE4Q
Kyd6JapIj22ou4Krlm5KFAK7C5JTC/Ilomm9AH8LQfcLxqprY0zSmIcY5j/YJkLW93yVKcELtf64
bVF5DAkGA3vqfKVaQ4WFOTV0APecmMSv9YIIHFGZwmr1Lp3r6vPTDCyQxf3lBWTp49q4HHJHp2Om
MHAE89jV1HENBH8ygEWjFpaQroXpTcs73ASWK7PWIQYLaR8jIyf+NNx5NWoM1G6iCbPIudY++NZN
1oe5KvWKufE9KdnsDf37+wVeT9qOcpj3sJ0aqWjEsfrUQqAngk+ZDXqTbhHwdosGiLlvpFXBxvzU
ePaf0K7fiv71bBLHmq0woGsst0DoAqBoTCU8bzOjCkMiZ5FdcTOUNlkNiR0PKWXaAZK9171U1+jC
dtZLF9d+6F35PUy2poIA6MIMjliiiOXK7gYRt35U3g6AVeqAz/fKnz3+8vdrsqxWXIJ/B1Di8GOH
VbO1cAcOzOucyeTQ21BZCvhoCZ+Y+SNmJjl/aroytcUWi+LrE3spa2w6+HPY6y/E3Npp1sqkfoX1
VpFi+moZC8/WaRDhUUYJgJEwDC8jGkXuCJyuRNI/jL1mh9S2UCORv+v6jlT9UpVc/jpi5v9Rfa18
85TMOKf5/pup6NlsUEfANyXx1htll8UcvIJ788HTYJcNpm2Z6mVQdHvi4EGC+Y1aTN/Bw+DXx3pI
MZpCA/7HHV8EaVztbXFB4hSN7r3l5f58l778lXKrKj/KDn5Pc1DmKiQBMsA3xKpN8NvvZkZbBNGN
HCcii0up4DfBRJKfdcamJ9cBRO3LY2rJh/rKrn0b5bPOX/MDdvVBvGIUQvO8D575mNP7ipUm1CnN
jFOtRFF5vv6fQT8izIufuYwJPpu1hDFTmpwbp0ZwoiNj3O5E43pKeU0edD/IoTt/rVsFaYYjIMhg
AvYhd+5PpfEtHbf1z5W5cloWm5HbiTUCRhpoqAAJ4Qew3XV4mBkoYSSyc9l/EIwowm9VZ85ZUafm
eGFyTAHp4gy8yIqetyQIT1ew5AXrjI136A6aBzzk7hWVro3f7tUbV4HQlL5SulttBwg3/mMKwN8o
m2fIqWQlfRqwFa4OdrASaIXWWBAmJ5H4c73skcQjTw78TpQVkc9imLyVCBrz8xflufxxi9cC636M
SukKOPqvjRNBJ4Sczi4GwgHqZaVVIJkh4xo/MyQ0B2+h3nhZR7rhM8Qrp0gWKZJwEr2V56GfsEhN
Jpvho5xg+YeaU0Kf6+kluyYCn/1ARwK7ru+4AkYTkQWe1NQMHFTMRz76Qm6/7JA5sxeIf7bf+MIg
TxDP8bRQKUqfC6vaMZEU8dJCdNVMDQ/0bRQM3fjL/R+2MDx+M6PEbsNzL7GRWiwwIvome22AbjKD
WrvSwpxF1W6Z8n541IaLTDlb80W80i/sEzyS9s6y/wjARupSPhdmN0exXa+x7ymxxPtURtG540aE
eZAz8doPa2c6AhesvXN6M5lZt8Vlbqn+1a0EpperC/gALUKofLFvKRhYY7H8rhZFPgPHQ6wO1ZHK
50isNAXMzNjAQU4z5Jlscve11U83XRJ8TWdjY3YkuupebkFRb/zHO6tIIoeFPywisG6cY5Ge1BO3
i2ahOnTlPdri8gtxfDHyYbwPyIcZnPfkXv9B32gyOb5zgcOZ8b4YHecXNtZRPW7FQ97OxXtxAAe5
l0ltQ74g4ofW7/p2dYCwqV3u0XBcUxAPnm4+Ol3bAeru3zGBMugo8f0q7sYE9T0dmLz2fgd/OIkS
0NkNBbRj6PrAuYVGCA9Tjt8L0bZ3biBDzlTKaCXM7GWKNd4qh3IoEE6UCuKrCQ6ucpJRt+sInZk+
1JNRz47d0kAe3bqBq4nfFnIVCQqklhV5eLb04wT6WUrclz5SrvfSgxI6KEx0JsKUImkA6fiS6jeY
ktVLfDl/H6QY4hAla/P3YYO5il1o0R8ZQ0vnMGefdsF+3Vb/yFlwQvRoU8a52JQKnolsJKG0yYqn
Ct+Sqkzo90mJzWyGky6iBGxYgXur9Q+W1Yds/5iPoRHMpig1I3M8Kkn9yYqw08FPqN6ZqKwDE8tA
wDU1QHyLnA0vH/VSdG6gUi9xvtEPK2F96kUkoGQPIWuRbNOTezjbGeA25wNlJc1ydkIIUZHtdA91
BqVqeQAh8AZaHbolGtW3z3ZlKyhrOUkE/Tm6T15cjcyMrM8/DaRWJ+Lqm139mwxCTEAIjnfs2J4h
yEn47hd0883MRjbQIin1TOFvYrbf+AX0/N3AMFT0vdLgojPQxqSitfsKUGy/+SA6HAnN3ww5Bp4T
mPdyNDw6QtwS2m5qHHPz7XaZQIPygshlIHtihbT6DrCsHLHXlNqLjRLuJqb3LQ40tNJKHdmBA5RA
XvWna1v4r0yDsyGbiHr3GLoEf2TdBFWi8FEd2wSgI7AmZ4q+bTLb3X9lOIrnJgTRh05qCfaqTILU
SaIHk3ljEIMeG+s1F5aKVNrExdmEJEdHVDLo/NLRvY0omlWLnejwFnIRL9fWpoKv3cgGUMCWKsYi
0iuf8f5IdjSq5k2kUrHv+79Eoo4aAG04JcwBV9Hx/BKB122ZHnrepjN1rPtgR730on0XN5o6aiuf
Gpcr7JXd/ai0h1XhBvRhsRx2CEPzV6jPq3QbbhYm3BqyTzuFhHCE4wDQzqIWSwjTsbxqcTv/DiEO
X2CpLYfnBgT0dx2NmhZKqpp8JK8UceqKN//2RWdcFjssreWcx4S6ci9uAJ/uE8TcMaSrF7xI9Fve
KOSbEuMvf2H5AeUGGhp95F4b5bbUoxGGeFz0cMU1rhrP4kcKcxu86FpBxaz9l5DbYVyyl8kmWqgf
PYUJ9t6T3+NkkJX/LyNSVPYzktgUgVdzFqgZrgRDFTv+i3SgqrKwSnof6L9BW5xsLfhXPsxW5I/N
plHJ0h/SyOmP1AUyavW3LUlO5A14n2ZKLqzS89Hb+tVCJaD5oWlmw32eFU9NaFWyREVUCQBAupog
U5lUe2YVF1PojfkNGkiUak0dGnx/greEY1flz+2uo7AVle0EZkYf7raoBBau2BWL93etoROU5ZB5
ruJdQsgUClbOwaU58fezHXq8YpfzLg+24RGEHu1fxoNIyvpDLmA7E2nsQtOjF9xZtrDMYiaRqUys
+LEabPO4boqu9n/fBPSpLNwgIRqBUU8S6+/RkguY6Awr6v1mIwtwMjzQUG925xh2AqG9KiH1fogZ
ko5lSn5GBe4hhR4ioeDTQ9hmFKgEUiwyXkFWBPKl3sx0LZYJ2bnFV3UDQqTjW0kbE/e1QmRdRC0b
T6thSs4PZPmu9PCG488zQVdvYP3zdVqYyZ5yQ/AhbRP5EVMrEp6wFghx/boFU/36dCYGR7aM0Cvc
1IztlNWK+VUVMQ62o8ryANG37dT6VVZl4zMnX8lXb6RW/lEYHDDxBv+QdB5OOnbq5BxVtTinwqMc
qnniFIyYe8W60Upw0/9fg7AxmwkcExSDU9VSLL2K0HKpOBy61uNezx2dzD710D/fZ6Z86adLQJjY
OjOdeAB8F4TS9S44SsF/2+14D5WstaUlIHl6bOX+tcO5tigljq07mOM8TvuNKCQjyOEKj+7K9AC9
irN5xg3GS6ECoLU5m1YZar6dIUXNzcvvlYHWGB5YHEA+FuPFjDQ8GoxeI0VGK9hTq61Si5DH0e1i
VVXsQNfPOPNbEtJmOJUu3eqZGWF6sgJFbRLOeW+/S+l6lJTa8hMEKWgHOaYKIcAlNTjcYm/pC4Ly
ZapEC5pgnDKK7rxeMjdAUIaLnDSqwwsxRjbUlwaAHAbecS4XyoV3QUdqgXsvM56UJMnH9DUhFmMc
UIji9qJaWA1u1x1u7EZRCt5yQyL95p6Aludp5srB6wWpmNZalWWCv/s8Rm7olBovg2zL34tqh47C
ogNIq0xxoNVP34BkL0+0ZzCiax9sMLQnRwybLElD7Jf878w1DyBlb5yKpo5LkMMPf6IuD5iuOyVT
EdRuVEfYV0k0THrbBMDsLsrMC3rRhsZ0LIziBGr7ME2gpKeJ1/C4ZwblTXzTAA/MZS8RIapDhnXL
nNC46R//OCK9RNnKKUjy5kSMF4Knr8gyYiEY6nAdRMrVQShcKqTTnSf9W9tE/mSYh7rxg9Y9Tww1
xeTXmJ9uLvRuW80wVlwEPjaKoufBmOQBkYzitGcHPamYDztkoO8wZOlHACbUTXDoHHicoy1MyRje
q7aolrghDs03cD5X5QqlbA6K0pESpXkQn5JoEuxCH+cMNJLkUMppEqxRMw07PatxZ1Ag+4aOWcko
zPmqvlTp55vMSt2Tc0HW4aj+lwSPY92vtt58lnsYSaT52fhC983IFkVJOEjiJbOaNvd7e+APEbqj
blZdNy8QGcDVCVe/N41M2Dl4P+KSXWZXjAP0vW2TycYT5aqXSRuP4fvdJvwgTHyPfBE8uc2ZwwRD
tT+BvDtfRqKP1i5Y+WROOlEWku/NfqUzobWmoO+2mx9Y5PFJ3HHDDwGvI6Ch0j5jUBPPKjvXwal5
vorzYm/JHgQF0Y4yco3JOb13eCnQP6sU2q+d80Q+cCVqaSfTtt6grWv+czsuENzIVVoTCwfUQm8j
Fp/RtrNxSQZ0nt91Tkwi9zHE1fV44S+uw1R/bE9WEXw8sCfHkjiEkElWxmmjIideAVHO/vqPHP4H
gCROCRF0Cw3ecC/G0YPXHcsP+ujgc4++A+LDV6Wv7AlW0+hUmCswG/EDMhDYYFYpWDdpRLbXssGX
bYC57BoxPuYrRMQKQV867rDniuQUaQ04M0I89OSa+Ya1auTPJ6GDOim4sHmYiclTAeiZpgo1uyeT
jFmykTd2ka3S5kNa2lnEYQiuhJ5YRZ/aokSrTDKZRfMkZwYPZu+seAHZSi9qBkuwgQpx6pcG1kST
/0ucBut+B16nfd1XNwAYR8U1XFLZHNkZ7ugNXo1vM9hNy80rJJrjg5qeqg95BhJual1461YWEOFJ
Kmp1KbtgcGU1EUWh8PlS+Uq4FREa/DLkvtV+p+0z0rbNiwTdjdngAWEb5nZZVgPcm7e943I0Juwb
OfklVkwoWSVEIUG0j4wihSciTulcEccTX1TYeJPSyAyI6MKNvxba30Gk0I8WunSfkS4rdrVW75N5
3vSa+4bkqsVBLVUFeTR4UUTOfTtn5z8Pf0SsoCIT+f3DAg2C/nFSPjt04/BcZR9tSDiSrZrWsecA
LFMNDxM4OgN0BRX7dt6f8AnJDpAkit0Tr+tF+voET0fK6N3ndxsGTjWcTQaGv+X2k6NjTEy3Qgna
OUH416MslOkQgKnQk3cNuOWWM3AcPo9dep+SI913CgY7GyU/QqORyX4joUMw060blQsKmes02go5
J2uQmPSmpS6W4At4uCCj08aSlmEDziMVnS1xurAQMr+NEX22CjxPdVUV0DSdIkK56xJiORnjqe22
zF3VUCWJaKtGqnbHrICt0jUO7nPriIj8MtSoMm/OtBemI+ehx0QGZO4otSnxZR0gtVbnKDEOJkSZ
ZjyBAyCDBJ7OtENOEmgc60t7sBSzXosXpAw7LWaOIhlh8BrUhE542gR9C62wHsZO2xfGRH7bw5j2
K+D1WwMRYndOweQOi9qIwiu7Hfy3xieAtSmP3slUEuyIIZtMEH7AueysLykh61VblSy+psix+xk3
ySLwHWXwLqMAQTi46zxWVYJlIGgvInRx5EaQWNHAjGrTIMK5QzsI6CtwozRoozLjF+CzCXbsT8Wx
p5yKGQ/EAzGqsPDuYL6ktPwHoQbr7ErTVk1ylVSOyWn9UDwhv8ZBh5RHeqJoUDGNcrsJjH08GwCm
KJiRfIcfG3AvUq1JWnpqqUyMyePSDijqyS9xZYhGFc5H8HlGU83f3yMhlH3Qjvpm12hw3kyvj+5r
h9Imahw5HV8+SlzpIBDBWc1QT2CR6avbAPVPsLEJ4yOAGpIXGH6pMGpO7KcbUjekwTpmcFRddB7N
MMUsY4hAVsEjXaZQVMz7oslM/agLVSW76H+X66gz+tBrKkUa0F65VTdbQsvFTlIjl3pC6FnQzyKE
EmgdG29ypK1+Kc7mKE+Dypn41BZmK6FnW3PXQXL3rhkwbaUKtWtHqFIg18NRUI5dTNI/URwxGCfD
Kr6Ak140vADM5B/OjSoYCqSSJFdPbwa+cXV0nPafhE1S1WT1abuzG+R8jAbEx2a0mYerNL051lAf
qBy+eHbtlTIB2XyVPiULmVVIGs+DMDhj+04zAMK+Q2bzwh8J4SUwKyFVGyT647uagEDNYObGSd/4
d9vMPxGoQNoyj1lqNyPedI9aZG+7wCn7Frp48l5I4UQmWqNo8/jM+ZhEjnd0kcXMjvmjLGVgulEH
30E0/WQH6Lm+GjLycsX+V+eHbI2LIkPQ8ccr9OkrlQcQsmu0KK+TYV5yMr/VZhE/3qdrRS0rFnzu
U12FXCgksra57MsJ7htK2kMJz6bs/c7VHSz3/haf8lepkoq/QdDw3Aniy5+kgUwgKU4h9J48rxKz
ods+ny+dHt2nw44pO9EfUg3Oy41ZklJmc1eItI1AnVImPgzj2v01CfI2Lebq7ACMQw28NNzn2qCb
U2jS4i9t/RbYVjZ/ChbpReWO+k/Oi+jWWDa2dGya0E2zYn961iHnqUErOJ3pi4whKCJSE9V7OIv+
v3TleeomTqWzQF1D3ECkb2bNRvqyP2vq/q1qSTu+cRT/CBvlVALkmDWNJ5xrkpuZTFLgZ6mbydwA
OsWCyl5FfwjOMU72Eno5/JIF+ERlLoFT45KfXc31NcItj8Lwm0M3OX66AgOHkHBBZzvqbNo7fZSF
Xx66kZm1pzDOlCOlXvLv7heT0aWoUWiGUFfZHHNuQi9s1/q0EwGZ7nMJDm3XXpc9iZmJdVJ7VeAU
mr3vKgGG1N9/WQZnIYDFQn+/gqOBHmlHOn3qoXolC42zmjZM1XGh46zgYq5XV0qt942TglbQvwY6
hZQy4rVmHhMo9sKi7SDC3LRpD0A1SqWeXbmVrmkvTiyFNAnfzt2vMfHmT6w539lLti/Frz86opvc
9VwgYx/qn4wbo6RlRfwL/MMraokiL4WHy53+47u47JDDj3jWpH2Pm/qtzsIj+vNt0lhc+SotRwTJ
So003GaSFNT0jJkbxPKe9IjqMlPpGzPANWBlqf375SbyWdCjDJ/ACVj4doZ3EMR93HKAewr4+qZx
2CEHivSTXVtvqUxhWsHIJQju1QWnobYeDCuMQ03ppzMk5Edpsz2Qv2XDuL1Y0YIH3InyTDMEm7mm
lPQZJbd1ufhJM3Bi9eIpXM2bCvU1EFhxm9XyHACL+sX/daBhQJqbGJMpPicZNgI7pj4pxWLzQ7PJ
jdjfvbdNrSkpzrkGjJeR53oR43vJljdEEIiMiKv+nPtpnn6TORYI46e9EeSljaj5teYwkAz7HELm
oCdTovcJJH14mKoGWFCs3WSP+dOeQ1GtLc3EPCBaKtebTFEtP+gIg0m77TmOut9utXHYJ4yuGw94
4HKYzQtUcbuccN8RLgHjq6YvhX0K57oNQKT7FR9reQKTCdcUJ4PQO/8RtBsbAAibYgOC2r8uOK3C
7YEpHJvnIhcOGBDEq5VkZBNi5urOjkLfEZxh+NxUaO1Ac/rKsCbkpQNWI+Erz58Oh92WyRRV7SBy
1jpABO5FtFCb2zMgsRQkR56MKSkpsQYXBCM80SAjoa8/SFDcP/tCDGEqoVwFwR3K+IX8hEwBLOGt
6iJGEe33L5oQchpwX7tN/pGTlo7CzRetJKeX3JAGIYinr/MifcctT4DZ86xXB1xMWRynxVrwcrFj
KuduKZch3qWS7q733WCbocl6onqrownMlF67Nk7TWg63hzwlkOkrTU1NTRQqUN3/rXkqrQUotNtM
YgjMcllcN/SA4NfrEips4SfnUZZr5RY1nPrz2jCCoipFvfMK0JA6bqMiVOoFwHPmgoLUuCU2Fwyk
gzg19XrFtrWBQSXIJrxt/LAFhmGVTqF1b0m5pVH/KSQAl5EjFtdUTlAfjnmKaOd8oPzmysVv5p79
IVv3wQBrLje1E09Dy8WBVXAvPTyeQCfBuDF4TvdtezoBkGOztNYdvFCV9lDvWU1vsEok/aeMoRGf
orlo777WRgotGqu3GMdnb9Ny2uJIsxn/HINSGM1EYnMFu6le4ko1IaajkPDO3O7aYJWHJFspB2by
HlDV5n6SPTIhN0ouNuJbWYJg+WxObMhNDc7o+cz++jYPV04+jjslW9xJHgDix8oZuHq6yQ58ErRV
3DMN/1hMBNubxgn/7L4xa1Gk+rmJtlK5dP001i81wxN9PBnAjVu0gPKiqD2qpvOM95xeElpY/jgb
3v57y5zR7AYvEHl4AfLVs2QPL2kYSs07DBP2ieiSQb0w4JHDtywoRKmyM7pABM6SINtT8cF+DP5X
kFvpBXQ72oStbA2dTUXj1nEqw7fg1OcE28jZFGeXAgqcycxK+oc3naQ0N4rg4Dhnwa9AvhhhBxRR
MNa0V2DqluvzLaPK+6lY/HrpfLCRSaT9LB9oY67b043OUkuRdRhGpFeTAbNo2ujYxa6wqZ47A5ok
WrCHbvmx1WYbsjbFn+0D/2fzoEeMOcShXOtN33uoKLjQBunr929/3YN35H8AmE8Xb5zYeo/4NdUJ
lP0Dwoe+geNq8GkX0XAb0PFUg39+HMHKlEppv/9+/46lYrc73Hsda9PMx5UBDRUFgwTUllqC+YWN
dTahgqUUypKlPgTFsL3JWhvjVaoXHcw2IMxroXnFOuERDB5PnBmy7HVBKeJHsyxd6qWORt6j3bcD
Id52b7WYSPDh9MsAOtN6gOXbmy4dRfztZknMSpVYOyc7cmUL0zKzSgSsJCKuC5FB8MnQtPKhlkr6
XYya9bsyIPYlButhBfGih5ERPulgeYTJ0AXyvMoLIcetHqNH848DYVxoHyvGJlziFg4+Tfr2J97T
7VcNyL6PfymYPbmJbvlnbsHW4bhGev6HahtIwWwiy4sRK87G/my2HdG7e/u6x4mpgTkqrFjiYDmO
u4uI7lGQaUQRnD875ZmoguK36WdfBaNTi7/E82NbRlBx6/p9bRGHfdNkKphw//X8KXXwTVAIQ5ZW
gbDhWdJr0sdda/Qaq7V0jRKla2nIj2Qta/ZTT9hwyMEYyndtBeCVsesFn0ZvLOQ+434u6qX0cdGk
jXSx9Uiy5N0TtiTSSfzIJuPzIZ8XCMDaV6IoK/TR7vcwHnsTSyxCvkYgL3T/7hycIr18m1Z0CQBB
k9q9E1PAtyMAiHAKpNVhNGdqTad9f7xyNHj/cTtWxs4HaAjkt1tReTiHi3mgNjiPe0PaaA5J/+vu
ALKtqiYoMXCijk83rzsRCv/2meP5xIuZuRKK6rm+dJlMuk3725FCWyazdYQVVWYp5KBYIQPfaVLU
y9OdtX774ENFnjEnSzRcEccNZ2tPY6z9GM9eRMcps2/J3QzUg4oi0jEildvUbb7LTP1uoBwLexmc
7INoG/9kIc2ZtSixuiox+GOls4iDVDPGuEDfRmv5vG3iInhMr27jgtMr1SkyUdg5Q9AlQ+ar9UfW
5KRZmcfomXcq+5kwra3OIvp7vTrV93tfp4Ia3ycx0z1zO1cs7dyoyCco4dpREv0QurX7kEfdXpBp
w7E9ybOE4ESToDixMQbX8zEcNNXThPdALq7Oap+mxbYezOWuMKG1eCAcoaYhE9I0qKqEPx6R8IXc
KUuSaAhxcLvIYR3G46G5Y/hWNJs+byDWlQ1E0RyHWz0BeIO5mkBgW7cxJL3P/0qh0LNrV3FGtkaj
ZQIbWVw/+sXAYJXiCBYmv0RWCJlEU8TVHtwirVV84rwVbgIy6Kh25/5rTVRpWP3AuSFSAVYcLd8Q
yp17Wuvl6f5/gSbiGw8Ge/uDCL7jExLMu/kmmcwDSyeX+9OtY30bxjw7hzrY4pOSsdwQiE2eLDK3
iU0rIcDyO7ot56x08UWxyObBwf+g/lpcj+1cg420TnC/9LSDBGfETWJLYWY+W1jfI0oiNufccKzC
zTstR0lYiRAImiFxyvvI5mhnWY9TxdtcGeWeqTCrGMkbB5YaMIYdqC0RahlotayjLuauYGamQKS1
Ic0o2a/fk3Y+A4SW7Ldx1/U7Z8pbLVZqXwi2NjENCRHJPDANvsF0R5kYZaOATrppCBLBSWTSnd4B
t/gLabwEX+6xavzgociPEN2bK3wDvLEqixRHTtvqKMCHK/L08MrDck7HjxJ1B/gt0Fx6V/69v8Y+
w3qE4B+cGfrHvgv2LTlWY0AqfWEFLvMfb8JVRVF2GOElisTdk71vrj4yjqJXYnm3792XcD72ieXZ
ba+Q74vQKBDcFdj93X00aqm+/PBXzNlidWopC8piaKxQAf5lB6mep66cyJT25Qqsa8jXYXKl4hYI
ycm+FdidWNHby7c8PNK1PKEJZ4PjtXLLQuMpEFH2ssVI9rAYowF6nSnEU4b0ZewkFDu5QC259Q51
7JGlQlnWIqACL7HSvbELeAmG5QFlrTsIOFIccL8L0YtfKxU6n/bSnWdAPjlwl9CXkpAvPf9hKNbJ
S+54aG4WgoicKF7ElWW684iTgzEtKSz8xe7nnCk0b2Ze0otsPJwqLisd//gmZJ8CdUSXFQhcOzyF
v2JK20t4k3GbghRaMQZKjZNp7ACpyW793/3SmuoJBGYti2fQR3ELIZa52Wto36QW1wO2pD8SkwQy
/Pi/Na+AF8TPrRWXneDeh9TRYDfZXhXjoVxcN5moKXWbnOeq8xjDEigJD58Pikf0VIxvZIp2F/ne
01+iBcZgfdSZVppXCbA7LvQhLqbdgeWF+/G763SHDfVv++6NyFdB2waIoRmQD6hRR58SkZIjeISW
Nz2Jw6x7rNsRS33V7iJHtPo7m1B67ln0dgaFMDGrYQr7YZ1u/vBwHvzSbGtlnZAyU4lZAMXWg/ka
9jEX2sP2E3aADwPwIL8vE3e3sJntkKjijdbUFhonVuq5G+OUFJImJgIya2zee1OSqQuuPRJ8WA4G
f7FmtZs0co86bVDOQEAf3GOfFD+UXwrvA4rw1r2kpjaZsYSWvcQ3uVQ8szrmt4qD8aMyQO5uWyHF
x84aPKD9yolphPVHLF+iMzGeWh6DFBHRNZl0sY8X+dqxlVbYGYd0UM9AghN8o+kx4mrIOqvbnlgD
5EDYYEypl+6ZiPGGl35hRpegsHdsc/kX2ztKAFTUeE4dzMiVv3tq9pcljt95l9FGkcDUH0MoUWlA
JZCH04BwmvZlUXPss9j66LeAoktYoPMlS2bITx+USjSttyPUXjmYUww6Yl3fQxZ4iplWKaDeMMTZ
rEwHbyFDO9O89A+uOGtjDN1zgaLEXvc7v9u2vkmCO611tKlNmpHiDwL9bo2sJu6UJvsM7AyhSjCx
smDQyl9wqoPCEhyyK7A+q97Uycf4xC/7HjAXXc3oGSzxGcglir3ccFD0JJNkNsc03poqJ1+1RI1A
q9IVbVXz1sKEECGetpdNOjsFlNw8jVnInXxKq00yBQoVMqcc03+fEZmIcJieKU02pkUCbZkiM2Sr
F5EchKfX1WpjkkY106ozMHflV21WtP0o5D+bJv88x+ThMCbRYMlHIOyMuE0B6GFBwOSeBIyvh6lI
Vi0qWbGvhbQWvc7pUUgcea7I0FAcYpCOMtWC8vNO9WmStxgfRj5/SaLAxYSVgdDqeDRN8yvhzEfc
xhYITC2+OR1blIw6qJY//BH1DV3M+N/kLwVYEe4gxLGbjE9EAkTfcvpzB3547ZQNH54Vg63dj36/
hrBGoJVcyVRUg8azWcISG5nPyHoN8WrdvuLVTr/VrPTHc/PRkfGnBMqAyzE12YvSOqX/ViI+RmSh
ub3yKfNaSd1a/6VLn+JVd01CD/N7WZ8FG08Nxcffa+PnzEyDKkQMotpCTRd9eG+eUOq/ZolPnb9G
uNUrQwv8/l8+d6VLEfDpz8GzebV73sD+8dtq3xGhJVHdC5vC0ICmJiI0gBQYMZqx+zrJFdfEGZt1
ygiwMtwBicU4IoSnPA4YbsyM+6NWHN4q0xwUynosiprAgokuKI6KIdhRpX8/eOJVZvesVr4uKsmd
6F+c0k5rj57qrhZeyQh1vdGDBqBtnrDRlafKYsPnt5VUQwxZGePMR/PVkGSdWnFbSuHA2CNL/J5h
g/AMEl9cGMkIlyPBue7eoRxmHSUrXKWc4kUXZF9uc0IX4NSpJaxcydVBMo0RFSqrYP9G8ad9/Mnl
vLJHNY+qchuJzkahq6p0McWhohe4py1SKP//ZH/6eYflfgQFkEgGIPQTn7BkKiMyCopzgqsO0jCV
pSYxldp0GUGRkQS1S8Ca12zUA7FkIPuoLrCrrtx00pNvbmTtVZMPW8wM5ilwBEHEGssPoke6hZe9
1jgyRBpSXBARBcWE/B11KOaQNRfvO1MwcnboxV5gWL45S0lbvVh85h0QBg94Ht/ot/bOO/QrcpKt
Str9vzZq4Kbg/Mv59DRlwqZyM/69yVlBGcjruzLfhkuhCdrvZoI2uAXd2Fn/NfkTJckfBarPG7M4
2lDLg/5AHBbP48/9DQ7wx7IKLapGUNuw6K8B/3H+Qeu/X1WRTyvU+JuSGBqBftu0dKAATRkFBWKq
1MENs/IHgp0DYCWSrKu/hIfqqEPGcyjCT2qLYvRJzGht+2+6KmHHu7AzD4rmVQ4c9x3JH5HXUeUA
RCjzH8PFHUsTmViSBWtbFIsqiBcIpN05lc8EX6sS8lGLYJXcQT8VHxFuv2keRTr18fUt4fdp+0tv
vJ2h1OGpHMkGgNB9KM8w1T2FojI3acmz8zs5jE7gnbdAimtUI8001pSQ68MLvg1bPGik1DjQf8Jc
LgDZ8ZykhrqtySLBUVbMoomuoOPSRaB3uuwwMBkO5GGywrfKc4rc+s5VFCje7UvFjJM/h2w1PZQO
h9541Uz4bxoWa2MWDFyxRaoemamnZ+IH6u1Fiu3+Mnx52w847kuxA78smh0wEjOIg8EDav2D8P7j
NEr7T7082LHheW7UH3UN9Xowlds1UcNz3+VKq6pDFNmZE47EokxB26ztV/dGj0UTJmQPOBB6RGja
mr9QV/SsADR5WZlDcLUN3fB1oHmTxISGbN26Mqc9D940FKzYZjLlTtaWfcLAJSaMF3b/ASudtSKJ
gKbQjimpM5SWe2tgzY2yUXD05syJ69/ODRbA9qhEH+zTQuoxuTVBUwCe1lcp+Lc4X5R5DjV8DeOm
Pk52rQFHm6SmLddFn12mZvdnngifNygDWrzTNLlGgJZxkjzFhNOu0xY8xqkiOpn2jB5qIldSg40k
SByTdQHPoCyRDsAxZeCZlJn6mrTm4UkovWqsez6rGc79AgZP6dkSgLMW9YZ/8rBdZ0LcgF/xbPwO
s8tfZI8nygFozrTNiVdqUAdwBETFfwsPzeKn0SOqkx/HKXtyC/A9KviruP5keYwobrfiboYxZuke
L4tAs8vTvpgLsBzlnXs+6VHOiNALTMq3SqnCGK1fJCKQg3z6vxgCRyU9hKn7D7myUTeHSpxLrr9K
lbYYxjcj4SGTbGZ5ioAkPy/8htscd3NEdwztfkAcxqq3JtEJblggCqjB+QBUnRUKuZddI9dzausW
HqmcA/xOq37edYub7AD+21ZdeuSnoquc2pqwIOBsnF+G4itwgNQbkPopbuOt82fqKr+VwD10zN/1
1bJ9y2GrPFMAm3AUoqWp1HOOl/vX+Q7wRZVfXwKNcSc4RtID+xD2uTH9arnPa+uPoFvCUeanjLQ0
LusDKbVUjteKs4ShB7UIqcA2YiZDiaAtmHZ/CsPJS/BBQia/s7lSlYJ90Kuaf3c1CJZBohKDXW1V
utTtT5Ss2iV6hvwQqjGx58drpNDr9pFaQBp72RBYOhNNoqKZ4AgDDdEVnPKM/g9ziWFhKlEgn3pE
cqktyTtVaaHXI5WhGcrgI1Ga5sQfqpDTaOMDgG8/pHWhlUTIwoUohZzY9THcZcBYTk/RW1W2Yncy
RMmJk5j0cCentjRfV9vKQbr8rpwRgn2Syjd/z/a9/yBjzPJbSjGakKy6Q97+caMZsy99wvjAvPK2
rIfe6E0GZMeMVLPVnK5zC8Q7f0E5ThGezCqD+9PUqpUky9OQqE8gPNcWqrcXnnVI74T7XyPsGLzN
+LmhqSZQxyVDqWWM9+jlRQ0F9+X24ZuHxTM0jrMwVeF7CLc9H9m2uzSvRcEJ6Ek9jVI3OKS2wFdz
kcij4ct8auWjijVxS6N8zoAY879TuMut9Cr54DRfsvHbjoLlVdVTE5/Uaih49QghTYsKiuomsFs3
yBRXHPEdUr6vhmN004QjUbqUU1XJRL7krLy4it4bZ+AIWJn3FcWjWHwch8onnbYFlo+GxIcVipy3
SuoDKHmBvvk9PiN5ApZaCLaS03RxeG5blbqydbVNbw9PlHEGPr4nbVB6mvmYSnpxqmOSg1kYJKy+
lo1WLh7KFGBgwlZ8YNKSJyHq2fpCBQMzXc1sUUryCpMD1oOETNQrNtXg5jxMMpJ3lFKrO26tp0K6
g+gHS3Mj85rSVBuH4z1n0BaXd8+vWPp+/M+WhnLrVj4flS0jsN4WaFeveF/RaGbjdjKFGLX5NauI
cR2D0Mg3degPY7VuP3EbhCQT60qItSTqK57G7P3DfswW5zTO0D1LkaMmomTvn7/pqqfeGXpZQMAp
BR0SZMp31PBBTgMvbljJiiekBw7iKJOYUVgWuvaAgkbJs9uTyOlOVJaUpVbAuSqay9DA/mMaj6bg
0wLhj5oBken+KA6nQFRYTSLwjjc9Kf9I830cohzAqzISE8lTadFpwTQhb3t0DoAcuSas8KTRSEzQ
L5dqmNbcJN8ygiYcimqTfSDVMay1Va83S15xYzVkHtZqzWqMfuw92vlllI4iAcUBhr6XypU0toBb
+DdC4qa3jguurVkuBqpKeGZtk/lMGFkr9EZ5wHvBeMgw9oXeJFq+uM+5pbrkRr1xJbIkxYq41YFQ
TdBEo1Jq52qQzSNxZ5HYCPG7qdjXaYMefAz19/fLwXe848d5VYDT9JLOhh4mJOe0eaBkUiV29g9W
CQwrM1GBFdkOkXlyquhIcc/ZyNeftwGejEbvgOSPb54HkQYwqIS04G6nlYTaFU0F1M+yeQfwn8jp
Tc7jB0vz9l255Pwt6ncBSpMWgavKO+ALUiEYGFyDqTOTgOl7qs/Cr4fFjmsupPE+aCaPTTOVEI6l
I0tMXkIThMvylRYFYTXnRDBo1oaZNA7WV59D/eFiy+O5EwSPrOOXS6OWfKH94n9Xfn1vfWSng+Xv
CqXkNHFGgIq1TYaLxJTeyvxZ0zGrNoNbo20au/KpSptsbRr4lIR68vNYKiDxsNIxiceNrkrVBhaa
ldAv1SwHTc2RRr3rdUpVTfb8VHy20GFmEGwHzIPn0ZzLl8k8/TjUNmcAAUe6ZJnUXcdxNcC2VeMa
o+yipaZr0wLUvxzMa8wJn7AMmxRXg443GXFzjZGqwYXPXBpFLWOfoQ6Eltb8zsprXHPPP25f0YtT
uwIbAlJob2vDcM8iwWoB/bJEj+gNQhYttY0gvmUfYZrlpUCvbaXZkGItXU2OLx/LBqOINsv5hFCf
TQHJwH4R6X+YKvwDc9ppMl1PZNBC/5a5zj/dWkOvO7IHJ+YRxBJfyOGPpyolN6Bp8nP1mzGwyYRr
Q3+VCwtFmoNdbAqPvBmpWPHhee0+pQae3xcTyrIp6/eqFvKhAC1C64Y5rsbVy5nR+gurH0Tsq+5C
l3jTrAQ+ccyJXe69E2WcWJkoLZOG2+smqmoIpXaFbMCGgx2DHxpWUyWYehUhNwShvxnq3opSse2O
LuK3mDrfYUH3HUy33GvCgtDvspQqjesEK+etDHh5xqbqF3wS51w4OfV9m8WWgU3HrVgulnTtgV4U
ocUh26V8AXIawRLYX/FUyxlB1Q95974VzO+bqPtq1TdUSPSKx+tAbtUPYyTZaCZS5azvqdJ+aT+z
D95Ej9VfVukEynw26FRRf6D7JgE0WB7hib7zPtR3VsbzL3gH020+TqXSoAaJRSd7dUHcM8q61A5f
julr59Ci8mI8L2lJ4EV8IKsFSgL0yPlwhlHueFeZq1f626Ug9T6BaZpfuNyfaqA6NGXl28T38All
utaWy19WqR+8FRd+iRfwWEuMh2XqVvm6iyfSTFE8wPC910UNcT18QYo/u5v5Q9nEOSBCz1IUuSIx
bbR+Tj5dzdSjMoW1W5C0SmiZ6vCLHhxw74XwMQe/34s12ZutCDBycDo6DzMDIjeuUtWEFQyyBZJt
oDPLRlk73TRX2UhIuwSJkzvo6JHSHKsD+2znQrJz/AKexhTD/76iBaqZ7t2L3m8iFxStbvTKlF0i
R7Mot3W3mgesSetcvEK4RQyPLddrVuS3fRRl/VnhDXZ1+iQoPLcz7/UFTeYap+FBaT4gwCVZK+PS
gdrV69qwmZ9BZVmlVuJ0rqYZlf+D9L/5O8VCYFIwZPt4O0JiyLB3e//n+E+XhIRQdKvyO+g+CMPM
S0bTdmtNZLIf22xF5b2ws/Eiim3d0DXH0hQ08ZRjMkgU1mUEgrG+86w9s8+M4P0LTnIQ6W1yw91K
wrhRKI1XFEkkgpnEbR8s9ujaIXDng9diaHmz1Kg87Ln/kgk480KtHlxcpdTBWA/SdKqfaisZVpYF
d0sA85y0tV7qTH/g6xkWi0SbRmllGnEf8SDtoINkdm0R8P8jPIAr+mvVw+m0jNKYO1rgqCvfNqUy
Sh/tV7xew6yU9D/Br0Mc+fJxRYSonFRNKC1CLXW1CjxF9P9auKaHca1q8Ivc8LZevkJC5nuPs2+I
v6LQJEyc9ZvayvmF5SAblxQO2cPauLayAkh2+6dnlfcYUO0jGVVDRiJdFyLussfG4JOf0raHWvaZ
HbSH02l2u+Yn8Z5uDrjD6svagtpiqXhx4cHfHqtzG/WTHXx4jau9tYfXEQrpg1f4HeG+cBFqCAb5
hdKrWX6FSXyHh1UlL0+HPw2q3zpQRBd8O8MtJOJsrGxWMq8l1LzaGDqGtjUtnP8WuILLwVBvOV/w
Sq1DeFOJ1Q+SCbeazYUYOkKo3Z9LqEQ/VCAHwmBdE7KhPJfOuC3wLGqQui0ZCo9QQwAoK2X/bR7A
p90+mJuvyPYa45woaC0QHmwrKw8rZPfZZTudz8hst5r3e25LvX3jY0AU4cs45gbZYUldjrbuYXi4
qNP0EtCO2xZhAqcJqIdmZFYaRuJacfffWt/dJ8Kl0+u6zL+mv5GxAXoVoR5rO88jDCwxUXfhgz/z
1qUf5AOsF1L2hUKVGjob7kLjHsZDNQmngRVxPUiVeCSuIe699eIacvhPc2ghOvQl92UxrwInz8wS
/dNUa4L9yHynlwn6FF/7zG0ZQPZ+1xqu9wRmQ2njpJ5wd6pNW4imNasEzypn6OkoPLFoAHfdVvYY
qOeKTj8UIN1He5Jt1aKevZjHYBt/dOPXgJx+S8vS8mTf6YUaNAMUxNcwyJJ4RA2mdx3FkimnJn4d
q1oHwPiLog95NHrIDcLgfzjGa8Nh9oJPw68PmAS8TGU6MWZH69tcI74DcnWKU2Q/SdBVSkUFZgPo
Y6H7lWAqcUyX6yhRY9d2BsrsrzEYQf0vhCmWWFP+X7+ksOidMZ+XJcECP9DHGmwdjbyWCr4cpaEB
aXqQDbf+Df1H6zpsNdfBv5lUDsHSv29CA/Gf4ZT5MtbZDqx95z5AO91AAU6PfgF1Ce3VskoRHID5
Xg/J3QBnWGk9bAd7CjToip3mMntiNu3hJx0aWuY6rLRw9dF8b5fITO09iWpb7pYd1dioZ6CEEkju
LC2mU0AIlpOqGyYVXD4lDC7vjWJUyV80PP9OCQZonrFubNV6SI1KWkwcMiDYCSrz2fYAJjoNYMoR
bsxO6wSBGTEx3CNhQNa7Tklutbq0Ej1uFWQjjy7+qwSwxbpzTTHtmlN7OVpDU6U8J/8ZLHBYRPhd
gQKlEFTwQC8hoUO175DG9M7aNfDoHceA6nu4ufqld2gxqX70UxymIEcsLQMsn8F+cUa50t1iyby1
J1DczIenNkm+P/KmDUJ7qk1z+VCI7XQDfR7zccjm22DGChONDK+w+SjPfQvryhZq6yDQAVWo5Qhz
/XGqARMx43RNnwCkYjfjk2m3pCpeR9Jtf+1KfR+8GdAuJEZGmj3adlYvXPea28yYEk7sIGi9sHzl
ym7HW/fL7EPxzp/0V3e7fpJJ21WrMa5Ls/rNsOrwJJ1RSLZ4T0TjIz6ng/S9BOIsqhJBuPqG1t11
T8RLpMd47+0+OU4dt5PXw0zJCYoawjOQIShjmRRKJ4+Hh7Ux8mkRAri/mzasUo9IZycfLf4cB3lP
La+IVsQ+YMIzoY8wo/QGJkBhi5Zk+ayofU+hzuxdqkYO4F2OSBlb8YtPM+L+vBIzKHizOuBN7XTV
l3rCclHtg+161JYHhdiW49GNjclkGrbNeyIl2pwP2nsQLJK24jSQ15erBqadSsr2afyuu/0SHpHU
TSxrXuqz2IqJ5mm2Ag/9+6YO5TmxAbDe2b6qNnX47rrZ7mPcBpJBrvZgBv4nglYpfVW6QvkXwqno
a5pDV7z1wOULJ9nQAmvOjtW6tKbGDZQV0HlYJstxaZ091bDmtH4OcGcUqtXw+VWtUv1EXSv1VjRN
RbBvRSbx4RT9gyiO8um6aSGLdDPhcfpdWNGjHsWEpm8KAZhZIIJZ96HS2Stc9kJLjRyXok7YdGMH
ihBF4T/R71qzXoiS7UZ8CsDX6oOGXmP6IXGHRM0wGOIaNzbMyST2GRP3siG3hIA6az2ays76LgJ9
ddmnzuKvHP9zGJpxn7wwd3UimZ0sDJpzxiCl/sSAtzuHODy+vKiKT0pxvTUlra58HSaCnZEvJcSN
rDI9apJRLb2Asb7EK+ns0WkWHG01dQF3i9VEMOV/eCLN9v/i640IOHsa70o/8f/ljSkkmtmEFW68
B/O6Zh879xbj1wieyLG0pND1gzYBC1qBmdFc2Hajf2LbchJnFnIQMELRHK23V2CYvJEYbejE9J4V
E2GQdkOmH+GwGnB8hX6eZtSmRaBf0+CMKtdmojXQyB8qd6hCbAAWDo9nd47wy8MUnzjRawnOaiKi
u6iN97hC27sb6mns6GybhDvgf6ZQzGF3Q/ttQUKx+Rs/+OYyo/V5T5Rtj5kGiOacrOzL1GCcrJo9
+We/TPbrF9LzezLUgTniiJmOmyKS/Jb8WoIDz1r7uppb0jaUAw0kVF3lP12WvRqQjYGu9ouaUfKx
o7xHTQeqLnpAxTZcoUcJX+p7JZlG65Ke+Iimta5Iv1LyISuFIK3NhuL8xZZUuV5DPjlw2t58EOHR
Xzi/rng880QeLs1IqJkhUQTEnx5BxD5v8Xs07USPE+XMNhSbZvNkE5q8mdGWN9ca36KIMCv1d/DI
XhKAz44BKpNhwt2jQKq4db+vW0/mfF6Xu4kckET5ViOlDCsNKj/jvACaQ7C3exEV8epmYWdnYyYT
/ZwU/hZ3alu2cB7KmEHnHRW4eDF95iLfavOWJjdyvwTBvw2BZBqSZFjpFs0Kt4maqxS8l0WVcstw
eUea3fI75pxig3bjj/WD++5hKOD3pa44wNHHnbMp9ECCB+SXSMRjHq1M+OLnI8jWiC2/XZTWAin6
ZqgVbmo3o/y9nH0g/jq/iCJe/LOkehDl7E6r4rvkp/UtsgPq+xujvBlTdr2RJ/kJXhtHPzL0CXKt
Z/cKcxyy1IqdM/IlJJAZ5ZFKouz9KqY1TuaT7psnmX9wgXBC8F+R8kLoQtB9nDrkaHGtflaxWsYQ
uEVbp4a9LQuxEYgBcJ/1h9VP0SYP5p4sCO4ABSc59A0mpzoYv+K3mMa4nK7Ey+FjRtN7J9vtf5Bk
KOIToIDqDo6otgvyEScTDYpkPatP4wQRn6u4ue7OcX+QUM+tWNkXTb/r3KWCOGnODuIYjpKxt9Vw
l+hiZmViMj7j8qLa7PRTYjtxkaCdu3p1bCf1B7TZlWiG8hrYJiOPrdbrQJve3LKAOim7VrKoxVuD
xrdoG4WG+hjAFZYAuABfcJz6/X1XlGVaDonof6Q3PKMigMWyCe0mVTlT9E0DB6h5uhGJKCQA1/zi
VIQjuVogM0PAQ8ZhHIwzDQ8CPziwD7clJbMx9ASQwF6pXKZ0sF11uGfDUMH6i5LHDYDz0JFdqHC/
AUliIj+0x5ETI74VxoNMfcSY6NgUU5VOuqmZ1VkmiL2GMUuhcYFu8KmdpjAXfq7yrRll/xprl2Er
EpCsvB+HkxiPpOC9pOeMgOWYO1vCbvnKE4g+vY+RUYeFnXz4oAXZ+P6fCEIwZ3ISHs66Pa1ARPV1
KfkXfzuerdeKVNkS5CTB5OHQ9xnxK1wDzvkhLBMiD4KKL+KCNOHMwRUbXhOEcUmSXKCUx9LEDZ/M
E+poSeEzm1Kh0Z9TEmGM1yH3PBN6nXCOHDw+RIHGdgvX5QUXDDQt3Hem3YOXaE2jf4vWsJds9lND
4wMW0rNbQy5VR4ibqi4gaqy4v/+MH31cDrTusv6npNHzuoO3jykJWPIYTCFt+D7KGUjenMxwR8bU
qo/pjoD6cY4TifQtWZxkWfbceqm1SW4haL8BdOLm+7RwUqB5uuY+ewESUo19CUzvdz71//XhfnQ9
trZsCCOFsP5VcbotGVe3P/yCleFiBNzmkBS39mTi63tT8Fvn1dqIUffGJZ3H165xdcygHWC19HmY
My+ojzFFhOCOOaC4PLZjxqG6OtdMEVKr/LBzumiBBJzgJiE/JO/JSBi4+ywZN9SDwCGWn4zBaAng
clGEe9d+e/JBZfw/rVTKP0D6oaSs3yo2pYob+X/HHvo+R2WHnbTDirz/KubVrJqzYAPt++5H6gzc
TyKrmq1yiWCgujXSrdAtRj9gE/WLcnWYyCIC7AM97aU8tZH3vBf2Iz9Xy7VQDEEYz4LApsZsQC1y
eNtLOoe82JJRCqDmps8eSdr6mcBu4i5Hhaq03WdM2i4FMJ1bwmw8YyFnRZGFjyVF2aNjQQQWjwqO
CI9cDY5SlJiviFE3MfAgMPelhPhK/tlbikCXydIpydQiJhSla+VilDH4G0JQimj5zOpp3imTUOTZ
RjdzLCd8NtZKpa7oe2thGcJ1+V2cbM0PfiCvGpLChB/j5AlQbwovJAU4fY/ZER1CD/0r9jEp2Z4N
wL9cNXDb6kcBJH9jp54UwRKxqaoOS00yPG7UCeLqYTnbD65lfBOqCgKQduPDuURN0xYkglRzcRWQ
heiiauBGW6JH4nyu65Hpj8fSCQzjPLa1UFnmHLryhW86w7362+PHdykuOqTmp1KS/jwRzc4I2/cb
mOUkFMNmxWHMx74yrz9tNlc9ogYzZYce/bVEx8srvA8HG1/yrBeTcTzstK4ElUxq5Ex+xXPak46Q
/8PqpPF/4+gImi1Etp/0rzxhiycDanqyKomjwEMPIxPOTFBPgYvachW/PBBLCXe7Ux/6arZTsYP/
i2sFIxQ9H7T4lNVGPAVHwUwMyO2r4v7g2wHnZKKZMsyP+AJuA5HZ3qUD7T9x3MkmWfK4+TP0OoR0
5IGuh+W6Ndw5FO43lv0G0ON1ytzR9QdfWjkhEpm4je/40uT3YorWGqoyYehMcEA2st0dle/+HWz/
iKdLgKfR3ak7iNr+soDhtCijFFMIOobGscjVgIxjMAxF1gocFiBJqLmvcaOPGxefFfwQHcTOz1L0
V11XtbeiQk1RMDoxg+VdiWEkqWSBT5BvjG9RwUxv7SjfFXTQUFiK4xYrXtFDIH7Mk6650P7L5stX
Gv4+SSB945VqJfeN6OIRdm950oNOhLkuxFwzfBVE1I7lmAqqn7DEk/hTZE7ov4UYgR9lxIKaX65q
rbsMgBp9mvtlElqJLR0EZeuWGTgKyPTc06TUjBxRtLb1uxhef/CLlHPeByua14qjjy1MoNQOdCFh
23uAdbSnZLK2dRzkca/rbx5I5kIAW/xANH8OJ/Ph+pCALbJph4bxZyWvI5PIGF770GaH+yZ9NRL7
rN50nmrwUJSaZR2YZZoSGdBpd5SQqJraU0nyH45TpFiuAB9PzwbAqg++eWkVG8AabIb1RF446f/W
kABbLbf/KI6TPr17xtdJLaT/GCo9KOq62jZWyG91xmeQpV45kYycYZQ/aLbx2OiWgLrCvUlq236y
mJylTf8nt3X6k2WF00oWc8eXuDREPzLF4u/t/DZSRIUGqv9xc1hTJKecMYiZcKgsjb8KFZjIwARO
fkY4Swsniun4evVEM8wxW8o9OaTAF6dEkbpN+wiMcVt0RXTREM9xGn7lyk/lPdvJSzW+6VKB9chy
HStmEEnLAlgbo1rdWghvdrT1V1Zw/7u74Ea+bAtgL/0b+1sg35usbYSSfIRQU9fzjK5iPA8nC3OE
z7n/OOEmC3JfvPj8Mb9UXoxFo6V6pL2twXqI6Gd76EyjhJjHqJ7sCOO/uvKbZCkDTS2vXSC/uLgq
RfmzsSPqsreR6ilpjZu8xzdAjWNMFjWUdoB/v5zYBQisLwMHGUFzAhWiW6TiY0W8Zyxihf5Nl3Dn
xzjby3ZNDifBlf9ZtLkzlhiOsD7fspr0g/W7Gkpb7amqfrK9+t+61lN5F7NIbr55N1yp2/ZEz4IS
FAlWspJ5ozj3qF+KAvVI5t+Bl/R5+wCFZBqfEidA2RcalDDVoY+H+Jkhs8TAWkXU2PX5yckT35PW
ktSai9aJK69r+qtWWZuYXZuM8wUKKZnqObLJ1mYMshkJqC+NHY2h6WIu+DAlmJMveVgXKnOFdLhH
hL3fsoE324Ra8BOpenAqWmMh8/rr6/KE1YAOCLaFU0Jtv7x0TpnzJM5ZJspomE4XM5YArK3qxpee
Mauy8szvt3AgMF/m1l5u/MPBLM6AKfhA8w0bBa8qcfwASJ8QxvALRNGxNGwCRo3RW6VQSrAfeFWG
HFZTUv2Cdgm0NJ0nQuj8Sku9LNVZFUI+YoCbKQNjmz8b7Pb6J0wP7cN/PPIk9yW2tEKeuEMhKHiC
Mw6Z12K4/pGDsA7hZbukzwVGmN8o6eR7wgwtbFRM9MpFW67GAow5XOfQGgVn2bLatx4QVQVJRLGg
Eh9pYjnKkPundl7jIRufC+BDDBC6mEiSmJ0mtBYNcxYTtYLtESXhWIilN3baQ9VgqTjITsWHUyoB
k5amLlmnK29TTAyje9ZuGhIIFY+hUhsBxG9dLnaZj3jPxGr1bz1YvC+U9BkzIy+qdLaKc1iOViEk
QwTJtXzbuiP+lJCXPI4I1PbfmX9OJBccrmI3JFSFFYAxB7vYP6rSYfSTZDZRP0DV9xKuaqcgdwlW
d8G/0wPi62+z7p5+8vQNCns1IW7EiktF9Odo6iBQJqo5i7UiQYUad8XuSfiyEwklXBAyGlR/PaXi
ude19JhWujBBJS0o2ugKzZQk+kX3QGceGQUVLqJ8NWQz6zxij2jrW8TKRBmhfdIe587dtJlTKyPG
bJDN33LwR282W82u2pmrg/d2wUTF1y6K2RvaM8+oBprYzmkIkUG4Bh2TlNnt7AWgIMFrIWm+liTx
3xqAZFb+nr4LOYimYyIvbahqyy8GbR7zsRngobK9ViYIpXii2dYGGLa3AhzxAqt0iqo4Kb1x+aCr
bL75AhHCt6PnOxDIGDIy7g2vITg28FtUtw0nVqsGM45PN6xqV2QWawPzLQKNabm8PB6ZkC/r9rcU
cVlNghdLEORNDvHYCOkzWS8YmoLHMJi+3VzZxg6e4xXnQZvJaaP+O+GOcmzPyIltV1jPoa9auYgi
+7xVH9a0NndTqbteVcUwssFT9OyEZblSzFu3AxN82hrFyiTIY34sVkw4OT/g0wlIu53sUaAVCO/g
Je2R6K5dg0ga7XNT7VW7SLkAL7aqFHZIKOs9PoXojUTO52oTUc83QDWzSMc6eTOp2AcSQ6zkIGl1
G6P2rIc+zbwn+PxCqf5hostGFLxWOnf7MYYDL839vfMWeLjNXgaMrLHNkHQi7y+/Bz4+oNgSb3MI
wIq+fYs4gn8D2sK/YEvK2+bAemxieHVA/OccISTPiBTiWPdsxly7VyNoUfG5jGgJQ2BSJdVE/2QK
1O7CXlLhaWqlRoLR8/2G94K0vxBI+ZzGixDqF9DUlCKbiMqaNDuMIV/4buCMFp2EILwnESWIQe0F
/0+CV1c42UUHMQ05ngEqKkKFCc3ec3Cq3ee/QpDMeNlrlFXAXz0mYuucb/rxo3v3nEoT+5DZ0+fM
yqh0zlcK917O8WaCUvCj9vxqIsZABUscDg+eemknxndz8PNPR8AUsqFTOV9ZrmH9LfUkVoAGjYdb
CetePkPpwbXxU9q9KpKk54xx5n5159zJGda5UyF8DLWPcujIl59FajXH8kR89tcv7iRQ5b/awD3T
WJceTSPCoHNG9+g3U+M+jpiDy7z6IZykt5cIqow+E0hdenP7lDIkRFDpn3xcMzcRG86AXmBHGzLY
C9ahhAQHH61EY9pOWnXFqtM6Z3oujV26MDbM1hAWIaxpjKXOOXpqf3FM5pP1Ktwgf8K/BHJq8QNs
IlL2pPeiaW0cTiica1h83I25ey150PvSsHsFBMvxPt1wgGoqWNISnYew5rHlhGDAbL4+Ph77BZ8A
UTSyiqkgaaSyev2aQBQEqTNsJR716IYFLPuSPAcnz6nYtto5MIm+Nl9xTeEe5uW5nAK+ms0ywAyq
FRY2lI+Lf++xlf75wFBCW1cUuFlj0Li5OUNHYPld0JzUOonX8F/8Oc0WOs0eqyqFPX1KIWgjdmCK
kmlaNSP+c+V0XJnHaLNA8pEWFGtWaMsmj3x5uUxG3grFjpO6dUczFAdQPPEl1ap4dUvAKGT2sjqj
URbmeinKQW7TpyJ9+WpsYaNR66U56B7s51eQwBuYOkb7irvUSZdY2g9aNQbS+ZNXHsF/z8/jMYYQ
i58jOP9Mr/ORgr/SnsNZsyuQ4a22e5pqJDYc/9qOpx5rB3YWYtS085KtSV42wybMojOKealP51/S
3iRFRf4rjUmG4pd0hk3PBsbZtDlkDRqiN2Gv9eGycr5gLWZJyR0SEXdYp0ZRbZfnG7df8OO3sQFq
Wljbokv9NvGtQENzYGl+kXd3+CEjENgm6HFZ6lI2U1gG81Yd+0Ec9QZDj/VqTCTu9j/4B0FwCco3
xrWfXsGkXCT5Gq/vVg4DmeQtuAyE3+KKbNDUcVJQmYaJOAcq9/h+2qOpe8muaTuWNayuYFafYX7U
20uJbbTpG+klf6/z1Rrff4watAiMKkGTfSRSg0DnswEeA7gd3Z1ECeQCexnHHbcJEVhWDlZxeSax
8ixfV8ExWwyKd11i8C5u2o7VTJOqoRMW1fc3wPFuSj6NvG5OwoPqdbucmeG+Il4qoEb5DOW/rGvw
dItuloSR+/CxklUOleaoxEn2uX5JJ1K8uUHyJKKzTSxBN/W3cdHZbQdmsdHEKqtxQf/eB5XUmi6Q
KUuldb9ztAVjxcziaJBuC80H2XhLtWR0Wot4YeLUh1S8/mk0KgboARclWZn+RU+nkuq8mYTK37Fu
2bOn1EB+VAtXB84iTY9KvQGWaPy1JmqKW16mr3ASJou0LelwmnmxEWDDmY1w5MfbmtSOzA+p2j3U
+s6CP3TimnEVolhpSYUYkPFcNrr0+3+9BIAlx71H0CKF5cT92VNpRsv642rOfKHnlU3FtCp+u/dW
TdgPctj8PeFds/NeWv+ThkZI+lYBanlgJdGEHsq/VMyPfCW0DEmy9h/OKs06MIcP7hONwUgXOh3P
JVskMd0Wuy+Fu85+2kvuplHJMiJIQH7HQwrMGor0jRMLis7M/D2se0yTpGmW81TmBRbcpmoRBwZQ
tgOlueIqV7edfyGiV7j1Q9VHMoCM+q4w1IUbGjW47Mz1q1LRXVFAga/qcGktGa5oHZi3VcRxAr3h
dgHd2inq9dVyI9ZwPCJd/jS6tWNtN2GHQgnzz8eg2VK3014kELzg1MXOk1hYpduN8YF3i9tbs6li
QAFV4Mh1mZAhe1s9pwdTsqjxH3X0QzwPIqnM4xEeeLzl1bevI6hj3tgh98+UZDzRV0NojaIJDmoZ
WaML/MGzzgYYGwgFdHznM8tXAJX1xSIu0QJ3GWni1bFZjKR+fV/G0EA7nhwHVi6QjQIKcq+fGJTI
Px30LYAjo7wa5kyzK1d0OEjCPYeHUIvGj72XxuqOLtR+p1sPdlFnZszJSQn26Twh1ZPRDfSaG1KM
gbNQXmIKXvOpAqtPmYGzBd8SLqpsl/WqIC30d5OdCeRgJF1AebIB3YelrB8Y2JXCnLGBnReezC4A
PRn9jhXvc6thWDITS6ir2x3yIiN7I/D8/FBZ2DzDVqQvFJK202chA4UhaOSmL1QgJVP1L6bEdLTh
sZf5mfHZL/Z6L2q4zJ9N+hDuEtHqTToj6y1hZWuo5z2wyLm2uhMXWIetUbkRseD24DCAXrO9v2LR
62GUb/QTG7Eh6T55DfdzIvF2akcRjmzVsJdFU7lWbV8inkztoub0vaQwgu2eNET158Dz1Ym3Zhy5
y5du/XcoBWbw/MJTUXETx74Yj4WJ30CftVoItjqbN3d3LHPeVEsesZ507tMWwk1rpj0pGOGvIGHu
7gpWP0zSligfRxaCmy1G+M1uMb9pyP6OimN6pJ0ivcd0oONbj7OX0hmHxWjxQ+zjQtYYiTUM/lNL
THKpsDsYTC358Ri5TUknxYiZ0lKqTx5cWcFsIQFwf2fujlzz3Rw7siB/wVFJxo1YqPcKi6TsXV8s
SSgyz70EqaZXbqzHrnyPdRz5n6vDw2NKC4bpjokscGyuWvp3qdMS2JqltR4G64j0VjnANIlNMA8R
unzLuHsTXNJqE1/vH1OABo67Vb0VJSRIpSCfY+OqeczBHiny7lElwmNla0syZMP/OZ561iR7p+t4
Nn487LEv7C5YTQXwPsn0BOdsC6BPrW/coCJZCrTJ844EC1KSOKy0ItF6mfFZtfkRRt3lTkslfH8L
rDu9eINXE/6Z/6+wgcoITdOzvnru4WmqXYTF59/cMWuVM9Qr4+SeUQgWfovDYJAEP5nETv16XJE4
YWNVxvkhryYIqNAXZAemZNX3PQScq7xFpfxzG88TGM4NDFx7pFzoplwZ5Nc/SEqcvctChaZHFcDJ
WdVz6PsaEZZ7UFk17dXgEi9y9FRHFPEKE8rCD1hFQwOZ4zJPh/6bicz0ERF5RVq/LfDEKIelPYjP
a6GPwKgSGFQj3rNJFHN9kVn1aPHMx73pC9uhbXi/gcgLRYVUUihIp1as6ZE/jZiattrNvztYV1Sj
BSXNZh8kB0c9ci89cIW0OTFInXwbcQaniUUHTjGMVHOW1V3kvMEq3QMlR8mkWZMuEGW8OkjpakVo
waaEGed+PjoHxzAwVQCQbU9AOdxsEGGOsopzNGu37UaY+2pZd8mWVmzlJcKFOCYwm0p2vYX991/G
n++OY0SuB9WltBNA6msPHa9AgVYlHMP4lOxumcjea8n2lG2ny/C8PBXHc/lpCuqiIc3sFy2SNwh/
p267Y0XoCcNA04Ci75xv3Hqz3Vl9+D3hpNNIv8JSeTjm3MpqdxGjnbgeiC5VMaNi5k1a66IxalIR
YBqwBGMlCpqkuBKoJ/GI6TAipSR4GxGtzh44bqdmF+Ux0/S7BKJ76imobW6IdrrxGILmjbLhpc0d
jOWpNeMRN+3LFiB1ieAjq7XrFOj38vhZSb4FR874UAi3seF5/gCG5WZraJ9pamf8pLRf6OxoxlDI
GEjKJnKRiheR8D7SnlrB6ln/Ktx8wbl/thEDwrwaasTVdwdxILJhEDOJ28iEQxAP2eK0ZubtH1Co
RzFFukytBGtm8jj+pAKc8I/7a2O5q7WhDJ5v5Srsl4QdX08aaV7RTP/BtdZJ6cj4+EG+X5Z0LC64
P5gH5d4iXtIEwSMKBlHir/JupXW5wnM7bSjkWLYnqWIGM/NDGVFvQZlPmb8upO7qAHIRJiRD2Q6L
Gi66tXr455wmIKroR/1zg0BvzPLpXWL7z4IcSEcIc+yrl3OyNRl2A4twzyjTtuA6Z6FtujmPEazq
/GbrXgBGlcgkvTKSDq3RAKiwIkiUewqFzWPVeHBDFeu5ZedgH0EmQJI4bh7aelZqYEWGSAB+Bcpb
M94RXwY3XZGad6PX9itpVinKq8T3LBSVYNrpLximyFc3ixEfnyUMSZfO/KE9aic1hBiaHXVXx6s1
/uoUitNsR/ZV41KI6d+/Xh47VZH3umufurAeuN9/lrbSnf/IVvJx1bESy+scNAfNNPkRx6kwdwyc
3qnvlk9psp1JEkRPjLN8rhrCxl6wO4w3xNmpOorFX71/7TEO9/3Sb4pzcDS+cuYWvIUwszePF/Zk
+84CKIGqjYH9cpHcYU+1q4cwC1YSQzC6kB2PJU+Kko3giUXevezMFHPXgIdn5SjIorO02TKDcI88
XuCvbpcVjKvg03IKDbXtB+l0OlwP5Y4uyoidfKepXTxWJ6QwFPreK8VpP09qCEEiML3EtK2nbBt8
YAgd+D+ZEkEPi9liE6xLuJf0fofBFb/p4BXNGfJ34BTJf8pa9BL1sCmYrUgOBMT4J1auN+gF6DkD
0ciZhBz6IlzlCE0FgLmQbdd6BTC6204of3XOQ6ODhjD/OhhLTsAeMdWXwYE+Pzyx22u5tQQTPdhm
BcouL9qyVEnaYDV7LSXzoSwIqD5BDnYPRxu9SChqsbuLsevAY58q6ejKqU068GonWI5hf8QeAKqC
nhYix1AAXMnrXQ3saM0X3eQ2kMLfoFBt2yyCXdGn1vmBKAKNJvi+KAbxJk9PlU9XH8iOjc63cqJG
eZecxNHOoVdyMIjoY40HqDq1561toCaAnvryO4WO7GGUmiuLt5qtk9Pr9XItFXtlBPqSBue9oXiw
i5rcnObo8CeeOjRTTucPsSB0mRdkXjuhXm7BZqDOMxBdFPHFikdTVjfyylX+2xpnSfmVGB73+Pnu
yvtx/oU9xqklBcNzfRRsCH/uZmbvE1F7OxDsCSeopsTZk+tMZg9kiESNeA7ocW2woAqyt+qZy+Jx
Jkq/f53AcFqRCAqcC266eKGG11HBWXIbKyYxs7JBDycC5G2yj6/OqdXnC78Fef7enXh4cURyxNwh
XmhUJ7HE2mVKjrTZfZnZM+nyqem9K3HgaIuEsIH32Si0GN9uqe2tY9nr9WxLwv/9497d/KGdcfD9
zxN27fy+aDcbNkTQJRf8oTYFjBokCdt9eNKZ+uBk1OXWy9SmGzayWA9R0HEqAlSU0yLj811FvX/F
/WdKgD/YYZOWdBawHthdTA4El5f4NpqXMO9D/EcQc73Xlm/hwn79pxN/NCoEOsFgW0LGWIi99Jpa
6QbSBwg0vJm9rp9PCfJzf78Nz4fULmg8k3Y5MS1xMnf/Kb6DY2aL2rVJ0oi7qLTIyUPgOdnskj05
ZqfEsyDz/4nfXYfGknDl0kgcBKCMss5PsBMfG6VdGld+8nGjSAXBgiD/6liVn2JNWP+oWD+ShqQu
kVPyRdJdxGgr2ojntpfSvMPDeBi5WIiM8TMdpo6n0wtavOdaCK4cdHL3WtLh8ENw/1NL3Ui5NPYg
8pFXpZ9Yp9GAnUO/WbXnCwB47dce8B/ioMIYYOZvVCuDLhh1FgYMbhNwzsYD42l0JovoyQkBE4l9
xdEhqF+3aJJJ6i33kNIR/2Fa5tfkEJdmD4ew3sDMWE8+hQ7cSvOeM+cDV3wbThzaWuxgIOgkDdYy
UBHA8co2uwl/SCJHHWHRtXkv9aLBpX8ymvNPJJ0GLTNT1hnzzwa9DDQxDvbOXEx/cSTkTx1VUckd
arpDAyisg1SonEKeEtcUczv5vWO8ADf4iBpi4KQ4UdBvKkSiZE8YjZYxh04ntwUI4SvpPi0xrUnM
SMxGppyH6uGBzqdu4flct7Hwd/lvdTvyX2H/QT8zm44nuUhmneyihN+ARBNXRAdJY4z6bIrxGbPq
QJyVpkbVF2pY4wejGSH8/iWAAl0OaBxnmLeIGhZ0l6Pymczuwt98q/FvrCNmUrqLjT0ekHFooPzJ
xtVHsoNZeNk1YkAPMrPZMw6o4XsqZcZqz+lBADmNbHXA7CB5sgetTp3EqcCLoNeEPN07kJNj2hpV
gTT3550hl9QBXDcoLhlmBGHZOvEG+gzAMt8vEUY2btMRNPCiRuTMIj7MNCeljegudkW9vnuzGjK/
GkD7HTS73tXEUp1eq7ePr4Uz8aIy8rtL31HYjV1d/kj6vHJBePycPIYLTFyoUk5GGLrp0YIzJwhJ
5vxsiygxpQEkNgld9+4w1gjD/b+XLp7GPtP+iWaUdQnreirUeH9PTbZ8wLyl3XrOFFWR1N1JhLxb
PrHhCmS9xoBCEYipBX//o06rjHmkij97j3vKt9qoK1vHBjyvMAIdJU09Hs2zR49FB7Sm2hnA8Hc9
AC2Y2SZSEvo6DivDK1jLI+eocd/LQMYbHwB2SvsdPOcF6JIEhUrdKkAARw2r8vo6hwUo4Ow7+1+m
zBzqx6N0wHkGxEw31y9jgn8MR8+VLKNnI61ymgJg1d04cMbFj9qVuMd7WWnyVjhShvgkMeHvmJuS
geG+yWOZun5pjz/WEW8We5xUlE18KTIqBb8SRibdehYEfdJZgoqQRzPkaH1+MItt/T5pl5PwXXiW
Kga/5O1JvLBZkWR7S/f4Dm8G9ETT9JaNnINGwFrsv0Y0oiwUa9Ey0Dq9v8LwfjmBOgJ6fZ0r8UdG
t2bu4arPRQBicW4qLnCifBfwdKv6PbhSj67LVMU257/wcFieXLmb0FWznNUGVvU2QHTWJGnTlQ/d
cmqizPvpirdvVrf0XBj+h5tOyh+v7DC67gxmRpPeIQq6Nfz9T8Su77mkMCTk7c9CS7X5hKixN0Oh
Ih5GyYlMBCpfx0bOJKJ5KywArRHCgOvyTaO7JlvuLGpD1EB/8JFrDCujHmq4kAvCwijtdbhKpB0E
Dq5k7EnQcXdF+PprfCxowfe+bRkHap0c2LLkN/Y+h0Qdwc8FssVDhC4ivDZAFFq6ilkHwx7hq/vZ
AXVxvk6sqbU+ZDXypjfaYeZ1TLpEoe8QjsEjILIGo6FtKWDmheZMEnD0YE+4WvPaVaW2xtinejjw
nziSon5Lwjf0JMIOnxrKJXAv6Je1pFWWXbGg2V27L/5It8ag/87NWN1zIOg6X5B5RE34ai8/aqNJ
Sp+3IsnCwGjB/S8yecMFebkaYLT7H15CnQCmgTWN6lKGY51x7L8ruBzmi4T/HPf89W2km0Zd7bve
khyA8fiGg0tqRpSJiFvQiK0pZ16lSxMvF6BUxJqX+TOLomDeiLUSMfoM2MGjNROhnLh4XCEGHcNK
GKI8Pv06QYxa5a5aLM0vkpJF5a75+e6LpEB7f0ZK08P5FJ17J1ZvapHZxFcBZzy5iffyk2mxVh6J
EEL3qxhocOwjSUBwoHmYHka1ojsnwnaRRtyYBlFpSDCgS8SReBC1o/3aIjJbk/cfoXMatflzSaVa
Qmp3Gd3Fq6s04rbUctXthXYGW6FlqYP7kBUHaqPjEKxgCzmlidTQhTxhypszUhReiGSGveMrn7H5
PZOH4idKYrKqDk4gSJJB4vMONKCSskpzknoaAM8IT3rHYvqCEQTMWYb5nrfCY1azUMyA1G4prqc+
ZNr4KZ6no5iDVhy+03nOSYCMAdWyLi0hCgLCEFOSpARgARPPir18t76UHHLqJGPJnvDzWc8Y4AMW
AlpyXQ66kSIMPzJ8EzPtn/sbkZugD8lGGF3Arg8GfNkDtcH5gfV87DkSrFTmpMYStx3+SZH09x8r
WBP++WyyCACERNgDfYBWLXsGe62pR22j/38GsvTS5ZGx4HzzRP5qmtfxcEANHWofzxD7bLP9FYkB
CU4HnxH/mphx3UaRBKbQMU2Tp5sXaQ1odUJYteHruIIei5cexKE+42yPrcckhwy9fwFSjC4+abSv
aP3/K85KZWqgylG/aFGcy8IYyuc2eKqPMvSoCkArU0xmLTlTEv72b9RYlCCElnyDvOR38OAGlKU4
UkyWXAGta5BzwTPVfN3+PfN74aTWoilYi3M59cfUEZk+TCI4bCChIjhVhO5L5nz//O872tgj8k3c
08Mw5ARaHLYiPiUzquJGvq9OmPCv6pQtB0LfJG7CVA3ovCaCVkc3w3FBfJVjJsHX9O6mJDnB3BcM
kcsGWkRkzl9l3YOjcBcqO5gXLmurTDTh5MD6CrqExOS8Dzx//uXQakGAoZzqFC8YB5addRcXJOcg
o66CozgIcmi68YLoDiWrTI+TX9WqOWG07H3d6OpOpseqQ0kBQ4sNHwzu1Z61LV+p+gYDhAeD58VW
CPjBFR60ISXUeSdMiKwH9CJRa5NsQmqhAAV8IL/l0jJUhAcVtpRUVtgkydRY6vHWuRULWkfDR+tQ
EYMD+Vu6dulMSuEoRM5fDHoxx8fiGiSFC57rRbmqjZmeKIipHffqaR+mZAen4y04WK/fZ36XfSV8
7xYLIFzMkby8egSdjb4pmBY2iPYNO8HwqmU0b+x7hWwbK4vUol0whTqjHtFLoeqDVdo3YlXzz8xC
Rq9oxUz3Ph0pDbExZ75NjtzjDgWDyy7WKAHB2glQWXhreIDwCYKznfQACyK123Lz0ku1fnn2/gUR
KWGfvxOcI0cMOhIf1Bu8poKJbY9sqQUFTZN4newGceVA1EcEZoVO5ywgG9+Lr1bQMh4tOj6aWk+W
dk4AmaWrXMMlqBXh6fetykDqhYyQMx7jzByCPP0m6UfZW73nAN8OokYjuUXJbeYG0X6nLNjeoiDf
QPewnwWeO26j1T2+OG6+mF6Qzaee/c9ISBcxlIfg447/7nU+CfczOaXJB6u3iAaIMLJv/t5/30QE
bsfvM7J7uWaDDoqEOi89dlfyAN22QV2DqIDG/L0yP3+LnO75IrhOyo80BDDz+9ejLSiOo0h6AXrC
VmIvIkrt/y0wNng8clChetBu7yT456kzzX6mYeuj21Gsaa/LMmBbxFn1rQXnkJ0TbsAxGCcn/GqD
adpZJA+aZJLbxq9sFCckucZcqaETsHQ1huU85c1G4GxYeZ4vU0rMJ/ReNmphbZvpY9DOVduyueir
GlqP5XIqW+3K7isCzSSAuSOE7pijtOzjAch1/FAW0GuULXkGjvk1cpLqh2tG7swXXYM/U2fTlLIW
fQxI/WcwcVP6y90U1/TWYXWqKv47y3QyZFTQUZkjyQIS0iRr+WFzasYGxe1zo4RzcAoSPYQhB7o4
0JLNAQ7XOUD8Fq1SqQdtX69x8VhPEfVsad+UJFccpBNG2M/LqXqKkZRGRjg0xk97OjsOKgU+/pgo
XJjsB+Wu/YZ9Be8WCMSc5yJxKNk+fhdilBPTuvfFFwKykuB8DQVQcP5qSoPWPcuHnKwDk6axiYwO
wdTWLjU/rSdUqTtkljfsEMnJYYVsyhFkjQ42BEI4acMWJXF3Ee3EuE5JPgHP6mPcp/GcDHfPAA4C
zQ8ITKzgZe7bKf0r/XOKApq5MGia+bWYRoLo17PTOVJM/h5vGbBs0gRiZjc1UjZZ/AT29nvFZh94
Ej0Mh3y0h1pk7Y6cBPRLCuDtquM+qnU+uWjHz9jiaIrGliPKUcT61xNALwPHB/No3vEMJ3wfAQgb
ctiPnNyJXZJ5J6GHtbX+SOR/RGAlm/wCuwCfQIfB9LseTzZnKG4QpClnDEFCnO2x8g1g1rQPSqwG
wnGjQE1ja76PTr8N/8sezO7VIsh+M2DkM+ZEzQqty6UmHgKE9GqUiYA+SKlwUNQYQFsklfuQ7m0m
8TA20kl1Iqd5bXl3IFSYHYooHTI0Bf034ytfQWsw8RV6HB57IGyP+JOPw2kz6fO10NVwSDRhZMX3
00zknXk1biAqRGjNxZ/ACWqOIKeHAJzSxpmfryWXb3PJkk+VFmU8IqX4SofbacP/tSzGUi9Y1Hnj
KIFUjNPuReRkg9/WWtLpIW3qAgtYhigZuKHtpnyxaSi1FwsNnICTIHtRcnkANyawNXMh5599rSQq
jVb9gIUhrOSRD4Suom/qVviCGY1dGmI9U2QGAh0NUP+OhfhArFAwI7tApD7RyIsRb+Ych5r7gm0Y
dTXLp0QZAy1xRrUGLIjluJJJ1cmgnMtMbkkQUGJXNYjEsfKgBdk4b3dFPFHnieohuujDtVwk1Va0
zjPQmbLKGhNgZ6LvE10SgpnTOBIB/JMJajFA2ep1EYBsMMze5zxJlagZL/YA+Qz8DUsaeGOiO17u
hst6nTRl3SMd7Jh1VUkm6xsz0W2B9aGPzewIeNLUsZ35Ca65Wm1NGskjOEapDNlbHkNKOxgfa/4x
QT0/PeZH/52PIIUC8Spq1X6ImXB356+iyBkLatJFtGI8B0Kr2j/zi0/Bny7h6USkS/Nob8wfR8iG
jQADo8yQgrDNPqjrxxj1XvXPmaJN0P1J/l4ey6slqvIYvldE67cf4U+iBYDzb/kr4CcfcPJZ41LH
kLZ581dwM8EgItBVxiazeEJrrjpo9AMCiV4eTkodTEPyS/cZLXqDJCMnX+xYP2EtEGqy61jsYMbG
2QLzz/AMeYh0/Qh/oSa80b1FHcRRUVX/oYOu017ePTbhOobtM7xx+erHwDFxOsBzBg97t6N1cYxp
xFzicNQ8U/nNU1utd2NyiYTAwA5H28L2vhDDdYlu3geQq2CDJB+qb1wJTBwbNm02Hg7faAnGYaBr
CZf9XPIjpSmtI3Luj6nE4gkGdu5lcUwYC2LhzG4DV8Y5Tc4cGYuntL4SK8b+UAQbqCP9O1Fyb/hD
AMHFUiotq4NhHACHEWzjAwgD0aLYJpefqgDt/vhx2hPvAa5lREPZ3etoQf94XfGF5bTs9n9UUty8
TvaQn4tg/FhoSUh7v7ssQHB4saW5TeRJCsPGrrcSd7fjPyTE/3EZvAOYuyMOdDOieWwdEJ9lcPJY
QuPQoO24hW4UHDRjlAVOsJqf/FU10luR/q0vnjg8xgzCvPt9Kcqm3FGutmFcfutOebUIqqMe7jVv
Z2e7RGosTmpDAjBCV3WnTn2/dpyooq1QIvsq6EINWftxE2OB3tLPhennfsfATxHqK8pJw/s2HUJC
bQerboW2ekqmE/0uBRtUIdWgK8KJnO+4tuOCLYjCwK1ExRHIv0TNPvsEZJJXDM5/qdIoJBTbg0/l
QLPvjHXkcOX+5zpT09XwVEXGc5pb4IZiNDKmFFc5xPeW9BxoKH9kPtguoQYH05j2yOhMZlDaNxgz
554QzS7kc4Gj151wUwurHc4J4ELmuCP5eWGKrlrrJn2Jw5VE5yTvWHaFLz4nk9iNjKsjDd4NkOrC
/nG16xhqu/fg17Lhpf6IBrT8BMVVGYgSsPYIU97zn0LJiz47S3nsNPizJkKwL4c23thh7FhHWPzh
SeGwb6L5TPQSm81Se75kXwDPBWbVOajwGBbxZ36QUHlIG5Wgeg1nMEOpug6dF9JbYywn94FhObrz
5fI12faxgz9TeGm3zWURTXryj90XFzUZN0U1xiQP8XDVrPQg+JeV5v+r/EtzctffmlL3ywW70TS7
aW73BEfbSvkh6khOvLmTp6AmIBOQCRP9788UBuBcmbJUgrOFteH6iik6/a7PU20Er7ROkAmXPXgE
bRmPJPaIpPmBjNBi8l6XoteTMEQ7ZR/F4fPIOVXk/8BH+92xblrfNVTXu10KC77CKNa4NmX/Stw1
Ljzm3fCGywaMSxYlACpboxf8by52IYE9ka/TxbOQtB/JD4vZFqCgeaX+syxO6dJaci+759l7tWfa
qD3MV3tK9mto0A4IQanBorzHcqpMJB5iRpAHkg3hVdVB62yF+zdvjujd+fw23gLa0aRqDOSOr5pq
bxJLIk65UQK22cY4mGm0Y0CcsHNirQUF8QPGWE4i57W4b9ecsJko1UZVjvh+MetCmJh4Pir7i4bx
aNBAIZY/MS1CZFo+UiXySc4tAcCb0s/sQ/Ev2raDCyNGW+N+0CKSFfc5wOvmEWdQqtF8TMI3Ic2B
3aqYkStAaLFnLYH8cbiVplMLYdXLEWUlvmR+8VKY81Jsh4tY94POlcidgL62CWNAZ7vnUbGCPdFv
59Q/A+lWNp2th6oFi2uHEELOf/YEL5jRlcadNH5zMsa8NIKbd0TCdtY6FhfETgilLoEahGG3VJVH
qmDZ+Xj8XG/Q/LKTdKhE3CrZUaoAI+DaA/rQCFBgfyjTEXKLHWXbyk/FbWgS+HtwbxEhZM5hZJ8/
R7nUT2HA6fP3nULt3/EtxYfBNTx2HT5xesEOp+gmpC34T0mCzrzH2pi0h0qDyhj5xPzeINlLiMSW
y4Zq77Zzjw41Af5/MhKk/SfnKNjyPQNpxFNyFBsQXVAO/C6z3SRvW4zOJWFR0XPcoJW5PQMvnbty
MAbmKM3JoMivAeh7AfhBomUGXxYdYTGtyHLSXl/Epf5ESgDMyik77x6P14HH6bRWetCYnn3ayO2I
VO16t5c5B+wKJhhdqgjDVHcPFrDUM4quGxdNG0a0QkbKULZQMG3fIjqFJ/Mb1t5okObeAYVf4/Wi
dUy3y+LafLSkEsB0c/D+4FiXlPjZ/QdGnauKUxTXYdNSIgHF7nrCBO6PrJhq5B0WYoLpeiS2YIL1
3hnJDG/X/sps9pZ+lib3/kHwtcA5ePsGmU36hYXQ6Aw591VKn7rlL7dfmkpFzkFZxx0iPvP4Mf7a
Ij8LJx4J69obLOdbYyd7eZbw198Auj1ooD3c+U6GcmCle9QZ//QsDL9EkKu7sfghEAgOuLeE29lK
mpcpchJlg+2bbFbRu+X9hmZz/2Fz5mPLNSe37K2lmgcckCKCpPu/baRBfiYwMBujGpwHhYqC0V6x
Sm3aQYLB2LHkgKBgi3RO2NafCvpIP29oHLRf2XsNoyn6Is8TGo3+7aWGbV89Xr5jjL2btn6/wx+F
7/Ppu1+UUsSHOyiFp24uh9PSxmiFkGIiyXg2mBWzpYNZFXh9/zQ1znSo2E7mdNMKq2uTpGbTWVSO
XMO5Yv0t5RooZcY6bF5BKRX6hNjXlwp4eJyczEAcm7BDMxa2JBi7FIzSK4sUJ+Kk4o+GvY3Wv5EP
Zv7KL6j3NAIUhiNedqh8akphrAc+Z/x7Qj6IaXIV2YjjinQ+TkrS2Gy1QVToze4VsuopFLbBdj2Z
1l5AwzSFpZgnkQNh70kcrzWooAx8kGz/JP9kHAfFLbZUsMJco8LWYG3MkpwPveYgYaKvUWDdwl6+
6LhjEVul4Q+3P2wEB55zY0aDsjj85JII6qVVobIZftcOLv8lj0Vvsqf9giGWh+TAz8ZvQ9VkyiHG
dtgH1yFaTv9PTE96PGuDSHuH6y/j/rgW0K3g1nzZWNzUVSyT72NF2PkiBRkj1jHBjNRx1UrsDSVt
Xu+z62Pt9W4hyUcsSlcGtakBrG6MdtXhySUtH6w2xgxwEfgWE1thCjPIm2vXKknM7CjMQNg2Kt12
ZJd1Wnw+Xiw23K3TpSIuEGuHk4vFxIiWyi7TkPMByVdbhWkS7znSffpv/lgR0EPSGrssXmnhhIjG
651MzVtNv5jHygmSoyfOTwNSN1bSi+YXNveymCYlhtFSOXMEqOH7WKq7GVCL227sLHeH/ZNqgxpe
8o49AryJK5rx4654dHF0R1Mstt+7W3mp9biEyI+mTUnE2BVKyPSqIsd3ZGiaj+I9YBOy6UlBAfCf
2dh4/7RojtF3VUbWvdOI1T9kQG/zPrRZlQGTt+qiQYK0JgBLBA6azz/LA1f4ZFnhWDvsrG4wq2cU
HdxDxu/RLSvOZQnQR2HQi4VE6UNAtYXZ6R1MbGtY9syjElggbKN9AxKXMXDNmIRb8gFy1JSvoJx3
VkP7Ysv2cs5o0Dh+I04bB7Zs+o2RczXjp45wyV7Zlej7ymMLOm5UuX3UHupB9zDRO8DC8zENrN22
UJnCnga70O/DvaE5KGaFlpGYrW8RmV8UtXd3ogLaPAwIJktF6NGgxPq5hLRJTietwWULTUtce4di
nRCG3wxUk9vEtUmwDbmksKk2zw/OsYVnhC11gd51eWfNUI6q4SUkLQNuApqw/Ft+PXeUw/45cT4N
JBzmZOxEIvhCo7noXa/ehW86/OCaq1yNVecIL1LxG/GCrJbrrQSOLcdLq/Q/VtsXJENM0KZumFvv
WCaD9EwdPn0uxV5B5piAGGhwNbuC5D9BSTPTh5a8u747y5l8uAlh9mh1baLtmnmInoP2kF/ZyIgn
OzO7i6rkpD2zs/7Rw8zUS5Wr4v2f3X227JxP43R25pzqK6YDpV/vlWmq4w1jPE0CuD2oQngurdap
iOmyAQ7k4sbSob2N8BeY1TxpMBT0S8TCiiRGpLJTZJOZ9HQ80mfCJoPskplcc9spc89n6XSWh3Mw
QBhOVX8n+Zenq/VZZ2dvl9Hp0MDUHZXgbZaHp6VKV4/DvtblMNKr1zBHEjk88iW7VQiW6r2ML7zw
c2FdJGCAmBzwoxn5ljU+ji5aR83OzXRt/zS2/k5e+zqJNgKw1AHmdoi1nIHUZ5+UX01+cC4W5ggy
Ko9QXx6CmbJlv0awehiHNsDL4qLCl6F8rEHU/2C+cGy32shueKfaq4LQeaOpiChQe7b4kRYjj6kU
gfv1RA7cKxubdm5VMlfUO0IgcvLKiFYa1fWG6xNZx66YCeiHv3skGC2XntPoWD7VOxPkwIuywKeO
/M3d7lUm49Czkjmv3MV1vfqTdTfZuk4kfJKK2dlauGlVcRgL0JwKu9ZHgu7Rp845nGa8NNxwnqVQ
WjhCqcDUeEbCcZY6pX7nxgH1EBEoGeoi5T9p+NKC2k2Gd3fzZLT/OxPMtiHIPYL1hil19RWSXbii
y/JFQNFrmEXiIoR0dZKW3/aYlEGkgtxj2WQzUs4GeXNmJI4Cfwzx9rDxTPc7DzsQOvDUSPlM+DE9
C9vt0NvivZbKQpFu9EZdDwF3iVJ0AL+EMEJmfUVOapRjCvNk+mzW/I7CfxvRhvnBl1Q/WKUfFcmS
AA7oYEm0K+npg7ADpPeAA5vBEfJf59aq6554qEJawICmlHVUlifF4FyGe+K+ndI5avSa0jewn7SG
vF2WeMFM61ebKPk6cTyZUUvX4h+ND94GCmZNE+5Gtmw3Yh0mwbn6StqWxeID8Ovh0luhH0UTfTDF
0IstYrMKIBUiZakVq87vTBjX621OC9HG8fcQbNgoXyneqFt54gyvemkZTLlGwWFu9j9gzt45kh8R
D164KjKL+AO6f20lMi0JiuzDC99aABXAMucS0Wob2pzv09Q3QUyF1CbLHD4WTRlxmcgN9OAd+1v8
u4rjbkrenE5kNn2oPz6+ydZcSq2jWHPbY5sOwlxPBc+K3Z/Dtnq8hk45peJjnfzPXXlWFiCqMfCy
Ca+ag9jX08+LKsfpOFnO/K1plCP4lCZWSmJvy4c3MAi6A3F86SE5ACHAvtbVO7xUQVhE3Akvalf/
CJjnfOj5Qq77g/Nes58parHr9iS11M1zctHbBg5El5htt1HQCWL3zvG22Du2LuF5O8c6Rj0IVdZk
SausphxHY4nE+S/AJvaXP2LT2+M93KbYEfen2kRsorP872aGEUqSyLf6hdzq8cMk+SKA6Lan1I/7
SyDRfrihnoWr9XhuWzHSVBBYXxxLow423UaGGKBYW/lvviYVmrKxN6uaj5ByrfJ5Mch/6cDF5erI
UZ/vAcm0j3w0Q+He4KgsZSOawDcSjAKVegUY5wyeidM6vubJmMEIRy1SJyAPjrbTGY691TSHITfD
D5mA/HHaZm5FSXcVtIpuaS+kEL5QlfsSu3U17vPcJkfAmI8U6fZRFcUI6Ir9S6JTMpojMLsat6xX
EOo5xXVpeJy3/CpsXGLbTpkOJGBXd7RfNba9AQNN5gVqpKaa2m5N+dhrlaDrsc31tqBYelvrMzRJ
jhF0Xg5lbfpnSWAZOaRZkT3TEkUFsOZrxgJmZ3t1eoEB4OUOCjWqOEatgwpwMq30viBw7bxKN+B0
InDZUjVGHDyk+7gRfswQyv3hKkOt8yjYp08mjtr7e1ia7WzupIbk/KPvV1LjNwE3rJ0DF/shyyMd
5IDY+3eH4wqIlUe6A0DDV5Fy4a+UIhkL/qhCM45n2LuUjXe45NBnsd+03khxisAUWRzBX23+Bcs5
EM8Ywzl58cB99roAq3iOa1p/E85aQ5n2WUPuY4bkv5WWCxEmQMMrLxGSiSRy1OhRP18pYO8vOXb3
1q4iE7BNKv3kSpbcaVEkdlQyBMTGPcM0g3KLWYKsEdrJzHRHqdt233LT2fFqqzZd+0iIBAu7Sq8N
wL0exiVEkhK4d+KZUvyjaojwpNZOKpdEUZSsp/MOHrNBU0OAhJGuKOX3KOpg0Cr0JkLDGwoVInL5
deS8QTaFXiWHqxKVy8MBlbKUhpqKaTJAA3pINmkYSaRfqZ73ShPESpqSEItAEOVFA69MzfIL2g9E
3uRBLmPog129IgwOk3CMIZ1xyAp+MW2H4UMH32aVGkxHxTFWStYxselQZCC7VvMXONMp/BAa2MlQ
MQoTzp8ue57Sn11UJFgOZIp/ebgJRIfb9XMn3Da5rSkzsHj+14aNidRmAB5IbqoEWXrCcEPLwwFR
8tntDzlS0jn84q+Tfao71IHybUSl443Na6BSuLg1PtUglxyuGwW+Tzk8x616a05U2iXvOBKP2SJy
gZyB0AiNSBL9xt1iro0Os287Yuuy6T9Y4MQbQ77PjUBQIQnAtWHtmntXkCzAnvHV5GYu9+A9y3N1
DxKeDhi57yOuRFAQkZi/QFZpHsJc13NbCqXQ8IPbx5q+9IAonBXqkGsl7XMZ7QH7QIBfC7c1tfUB
g1KJPiQ2vQBG52w7ULCj7YcwWeiO60T9oka4V9OUTfRjPeGh+JWOhm7sFQ5dbZI84C7dUldJc2we
NIinMRy2lFmXYb3nJyZtybgnmPq3F1KPtjajkQlCjIiBv5kE2986ZnznMZ1OeLvyp8FbonhKoFkk
yvJUAAz5i2MvTQ5FGyd3IO24th1iQUMAMzbrZKj+mue9xobRMEEI+sbfIAghyYRQdYSxd8gMdCi3
W/4lzTX35TvNyw7UBk5XxwpiU1zPSCLZFE5dCPK5ZWw+qc8qc6RYSkitKnlPhg2scwWY1OfrMUxz
M5PbDj0D1jO8ku1i60jGRl2kRIIc1yKhsN6sqt1f4BtL7PgWyv/8O6vFmMWNYCz3yPRI2bjL4ED9
Q8hWf3lE8xzobrdqBxQp3L8bUwhTJGE8maY2wR+DJaD2xl8NLSx5zp+s9bQKMRn8FcEGQXXGFq4p
lFU3ICq+3LrG7TWf6yZWARBCJrO5uvNQ3ZlelQEEolOSpZpDuROJ+yr0q4OWnH6Op75pOz94KZHu
oEd8kwltlqKSLej6Hs4VWhNQi6PaeoOmM8wzS2UTHc2//zUQVfSCu7PcKRlnZHcdyfRMRYf9clsl
k+JEQWvA1z+1w0aRIT9mXBk12abjnixSg/O0GCemBN1BNlODeKeF7SXygpbfs5wHja2hGRIN9W01
JQWYy6AmhvU8YqfD2MveYbHy4X7lw8Zdm0uI+VlXUm6Zwh+h+KToYlsyzjqWGnFr70hQWkYH93Bs
J4bcoogrNYRCdymYCT4z2CIlVJ2JeImCKbmI8Rs3t63XahPOo7P+/+Qmo7R48BvI9Y+AI1e9iW3a
Tc0a42eG9eLF+EEzn2pnuaMveN/JgT9jKvvisgYPst5aQvy/NjtnIRYaWf3iJUWKb1e1+OCTEnpZ
XIOQfPTxN85z+GBZV8s+EGmPaM7KcPDIaTzRoIowaPcrPVOVxhmtcVz260t88Q1Z8bBL+v63LIon
e0zKgABoCCxVSG80d1IVi5x6r9/DGyS8FJs5gm6grnOUCRfDElSDkrNbwpvXFlkXBlNl/vYnXtrH
u1kn20hExIV7jK5gsN/9K54Q2y8PjyjDVhvo69fAQ+sJgYUlWN/zv3w0XNDzRlhquuW8Afdpslez
eX9MdIoaK2ETSpi0nu7EmBCvgtJSjziuTcQtcnr5CjYyXmp3guoRu7ncxz6acQn7T9OnpLBeUcqX
buiOe94hs6fSxFgAC2U3a6f+MPWQPG+7ztoUJ2T1aS3n5wimCbl6HgjA/B1rUqjZ0fJ53oV5OHg4
wMo4tW8e7MpoNwMTSmqo73A/7wPEo3BWnAihQUwxni/FBDzAjbNrJ+8pt2yURgYfMPhWyrS2PNAM
c8iDJUWi1PNuCH+DRxHQCPnVHZabRt9RtPkJbDh+Cg5aL7+klAmTqFzQsqHJx6kvncM/0BEX/fX4
GPV/HeycfsnkxyhbQmcIrL1xLPV49HxxZ7zt1OMMWxO7gBjCOOjNXPlWXeyuc0lPeJ5ZvRpoim2i
NBmaRGnyc/41kWpIZilcPVEOb7vBhEMG5++5mKCRCLUfaBaBprWrLEZAmzy7h+cP0AxWa2iGN2jq
L3ESAJbA2jz7aFfChWiHaaq4j6ZKaTiOPSvPI17PuT9Grk+TaLuPesFojqD5fi5UqW1ufXuOcrEt
utRgZnn/ao3k85GNm98XusTm1SRL/BxRpLgZIBiayfHys1d21V9RVgL7RnN6XGo0j1Xzxj+5hMXp
9gIslkSdoDV5ws+UW9ulYMawx8OBjUPKAdbejX6e6Hmr//wRm3fUi/kKhGX+PS+G8T11/6aGk50k
7msDJx112/NG4ZzeT8WM+PM0L1VmUX+cpuOhfttLQOnI+/WNXLzPHXiSai5RIMHU5/XgDQQM/iCi
7QlIO4oV69W1MBOotdcozuhRtOM8WOCBQEgS4ww/Fiqctgh1TTHSu9JWgGiPgJ30dGRzbThnLgSI
oYLhARsKVM+DKdsa5ziBkEhwqptoinq3PdaZD2Bh8gcVBpNhUvF/b3Fe34DBi2ravtGwvrbFYo0n
XWccsFUk6buezfuX9pAeVSaYjEDMCACJzVASZ66DxgAo3iBYKidlN1Zla2QEgH0E9LTs8mz+67tC
7VlLOGvQfrgp+ucg51JVmTt5yrcgZcSr4A1juayWxkAigRhnubcre+AOs5OT+420sGI8i455hwsX
ilNZesafmTvCz3QQI4rbF4FkUpyD84dvg7D/FBrSGoBC9hSX4HKOtZLbXpEB/uKVF/pD5vz4Gtyq
m5oHJ5ljO6OhEOCpKvnxGGikPwt2+G4/ic84qOhC4dYoYF405cmgEeefa/Oai9r4Z//e/+FuQkbM
3sEd0/XDzZ5WteuGqGICy2IEVigCl6KPdMHIUI31XRjJX+S4fyfpX9eL7K9UCpROuXssGHYLU9w/
gN2RHys+60hsIXDLzbKVGLZbStiLjYYc79msph/yJRdF7VKNqJjaQlFITNyk+gt68rhPoSLoIms2
lXZdgH2hfvSkewvwlrdQK4QwuA1aZnhuWtBR1R+BRXL2GT6hYmnQMvMjVHtJModJxz4/IS+pq39E
R6K42a+mfDV7qd+R4GqfP0jj/yfeMmSQxqxJnd01IGPksAY6IfXTB+n67Lk/sf07QvNw8KZk5EMS
sJWCpFPaZ87GMA2YwkMcl3mzVjqgabbrWdQAc+z5UeHmUC24ynf8X0W4HOmmcPRNV00qvKA3aQUp
UE99B19WhnHl/r3RfBM6xCc56kiad2e09sV70Ynzxwi4Nq50fVUu118P1rlNHzpZzpAeCnMltPjp
sFmF8WFL+iajCR+90ytThcO6y/GLuAWLRJ/XviXCktGe7JYjlHnaf1puqAs0rdnJ4cbuGIKUw8xr
LwWkeaM1Jp1hsNtrD8nxQinZR1KFafZlqBqpU1UYJdpdBhmU4TT3scAJqrKNcqMt0AB7zxZM/6Yj
OAN5aZUl40HNHvKX15ElCXvcXZlApVVja1c+w2y6gsOtxWMZnixO3DGAmfG6LvhxAo3KhF1E0bQq
WNdHB7+dUnMwNPUjjmpTZOkSMBL+zQxBvls4MPxrjodCzu7SiRmREEEIBP6ThB9F8Z9PponpM5Qq
04DNE01WOHnnU7JkZD3zaXYc+UB0jgbQQ7VDqINogJGCb70Wx5gdH5R8IUeCrqfW4zcDgwofvico
vUF8jCOjiTfgADwu1avIA9BXIPWyncPFKttTxOge591T7JukRsj5zuDdsORoYfY6owrpcbc1GNqC
F5jL96Zoa/cz1xBT/oKIi/vyDltkScFwgiDjUR/80HjCuN0ZsgYYiA7iNVdrRlywbvJ8NR/+E4V/
F/5iydylBt5wQuklN0A1FnZlPTdn0E4MB5+xcLK3RmDdjwmW/3VqqpwqJYa7rGDcAqAINtOtWvyt
5yjQN79lkgNtv2EkvVf9AWrAYwdv8bcWT2a9XhoCR+0wXrwUgmwCXaawFmGZg5cznLmdvRTztN3D
1E7cbzcGHfeDl0lHYAUhlXWgBnppjHq95T8sLl/OhS9Kk8irCBHAevX3fjXeQMBH5NZOFdsUR/zF
Tw1FAutjOzhP2M5LNEBBr69EJWJWJPisq9K2eFftdSqK6tXIew6m/zI7d5jLqVUyvrYLgVYefrCP
/nzT5KtPgJTYIfqqmgkFmc1EHJJEaGaajrlvEV/SYp6YhTawIANBGSyYYv+sC+aBHIP7/IuyX5Gt
86WuijfWbvNIXKbsirYyJ4fkHCRW/HFt2AhMivT6NdoL1w3rPX3klTGpVc37BWqZ7fLg2pq0uFqm
Bs3kRuWa4HIejMSeSFTEnARx5AsF89+44ZGBYmucpGMhkHu9oZHdMy4mRGFShYLISc7aygldV81h
r1GRUolyqCG/lkxJk1Rps5MeWv05mfel+B2ZuE1sUsllZ+6s/YM7QIwvdQwsxtKS2ndRtMjj9AAH
by9u68E19ilRj6s03c7/vkY7+ShQM4H/9j6gWgMI3K9a9ALBFLj7SFeJRaB1W0tM68P/8JXEVwXS
C0Ee9x5H8jI6xW6JooIY/z7j2/XMXYZNA8qDXbMmqmNgF8F4ASCGN3+2ddrUMFH1t1V0acOVUwwK
2i14gj52vKw33Mh00vdfLYWs59kZ01P547vi8Vad/aeadFm33RrTWCbSPFX9Zm8DXydB976uqqeU
9Oijbi77zOqRNw6bsKDVay/xaAFmNMvTf63awSfezsl1I5I3RsXnpiMoQ8tdotsevyFDcUofSAQt
/4IIqui3qU0PpxtbwWferlMMNLdCmyScmoD2yDEN+GW2kcijgQ6r3oabSpdkxVsdj0V5EQdZOwXh
mc/djcFTf8q8CD2m6SGWODbUGsxLNSHjtiezYtQUBdHTFiwqrUQ5dGLF6yPnr3KWoso5iOByWyYo
QuLrvfzdxVr9Nqqd5Pq3mYg89bl+ehuHHHNo2w96viXHBGE93ES2eu9Cp6F1nqDexzU+sPMVrIvh
Dy3eIAuu04sUva+gX9YrukjHWWe6Jwd9JhkRerLjb5xI+6ofESiTCSVgyCqbb8T6AcNjaPEBKUQ5
f4wV00pg0pi2krNClTXrjtlgTxwxOhvO0ApE6PpRbWE1U+tY4mGvFM1FZo25BhRLDMPiRCGgjdD5
6nWHJfJpr+CyTUqS+8tJrB+COQy1wxQby0QHjP6OHHce8aC89VTm58uTA6bno2t1C8QniQiDNRoW
6vMereQTIG7vumtwdUNMl/TC8/luT9sKSwAh+Ge61gKUu6qzfNBTKAHXvGBtyPSJDst3gitAJBZC
YGTyHK9j2ECyWHgsBVvRR1wYuVjSp6LW1OZVL/gMn93l+4vwwsCV0WpB3zMXwtuNNK3WBfNboIIy
KLlmW7rIdzGiApDSA5Pq83Ywf2EZ2rVVHJwHza70AJx5IK7Ohgikf6uGQFbzN6X+wniKawtmKQw1
MIG05BeUU/dJFeYlyAg3GMYVz0E47YOIkByx6X/gKDoOaAaRSuXhJV9DCLFAhEvkOAriZA5pSZ6v
yAZ7MlDOWzO/BFPhb/4acB1xyIV3Ny/bIMLLVbxpqDQFouiHSQ7h415rgjarRTd7ysf/z+HSM8Iu
biOhOcAFIIeJuwGhS000xAZz1wyGEgcSy0aZUNoHNcw6IeCnmB21dEPGWH36OAp1b4zaSOTTLSF2
wxVvhewKtAV/8l7ygd5/3GTEoQLUzmGOpIBTNZu2Mtywg7/WCc5ixRaTUPyn70ttrE2CsBo4u9xU
PDP9dViCmVMIGcnKfRz7FXLFI/u/+4KfN3k4OBqSLdEI2uC4MBvvCBLIcApqdZ3lRRaufBBsFH9E
OtX/ly4o8vcIw3hVWVEtaFoOBLCjJyfmePywnEY8/9GB1xR4QsHenKLG5d0EXxlDj7rSb8DPQuFb
4ysDRsRyvhOURalS0cboGz0bGiNpiRBjTJT1Zz1k4K05IlFGr4CYCA6aVdOoSXa14I6NzMX0bOv5
TwMwC6LtjjwxvMa4ZcBWZGebhQx4+QfvD8cHUWVjKqeV2T7tYWFp415nL46J7XfMYbl76I0OsoMz
uP540pZ8OT26MvCBxT7UamWvJTrnyCJMWKlR2F4QimsKslbkFyCaLott7uR7SFhF5RUEQ0Ddeem8
YR+69uvQa/IXM4FbV3dpEEZanpmg1fd/KKE8oDDV82BZm8obaQxBOgHh7NEXaGbZqI5jPGFgAstN
i6PyvJj5rb6pFugH5qjBmMfEixS/tgMFS+3MsaewuvanxJupFQbgidfSAljymlFZjnrCsor8pZRo
lVdiRWd1qUUOUYgXhixvt1aPzoDAKeqWgkwBZtvjpbob0eeniwLRyWVhVrp1CZxAlP7DKxATVnzq
x4rO0mecmO2ge38a3WvwNsGIsJ9W3i4lkT0+x6StdW8nn+0xjNudmOs6rhHJ8GO3tQjesxyWpGFp
bt5O/6d1gJIqaJ8GXU94x/QCxlYN+N5lDRLeOM5+XWsVaC7GMMWZRqC6dFpfLLSb68TzRdwDsz1A
E1gP44GxRCLUMJnF+bqB4kcbjxwbic+WiD8ppmO7Q/H/PDp6FyYCNmlY/R8si3QAMNF5PZs/OpVO
qkPcvjhJzqFe470Telx7en2ePqmvf8RJPDGbbzm7tKh8GjZMH4PA37kfU0HpszuPz469BEU8835W
heRPYhpbJN1F/M6QgT2fgAW36CmYh85Rwyj9WhzIDhkPuGnyU4xWeTv34CrISrFR5Q1S99vLdeuH
qU6hryzqI1v062osUVJU7s5fUNdgtHhK1JpFOciRm0/TokLc7tyswQw5lnc2OFY9he0I+fWJ97x1
7XAhcHMmxX+SuEO1F+KvMppNJYU598EhapndEKnKJCksuKjPC/un+iTkxDqMVUtaeIL2Fw6kg7xL
NtY6zjoZjDXCZm67RTvvIK6aizisrrrq3ohvHpG6X7NLy82xyuSWGVkNf6pUO8QQsFMJdRiFGAro
aZFB4aOzZBjuVpmaVPlGuH/0QFcBkvD0vGV5Wi4pXP7yvNggSbsHDED3UvNz9QvqYNBCFnAIKDoq
wqt3tORobfKWGx+Tl8OTI5XZpFkFdlsVj/yDLYphrVDxgqQTB1QSXiAqL5qssjlAXZ5Z0m9voIWz
vIiTOGuoS+RAq6P8/0yqU6yzbknMVSIbxTyCVLP4ivH1eeN0BCTw5KpL4ZW24Hc+L2qs0oT8TiII
7WkMv0LlkZ2tL437a4GgIZhXVh2putpIeSueE590OP+a218wO1M2nXrvGx5u1c2vU0BkjrWtcVL+
naXaPCqXgo3VybhgbMTAWPH1aFiPvOtxKat2CwvSSiHDQnstGo47krVK//40L4ggYaXs1eZv2WSQ
4m9nQzUQanKFuJCLBF+2SxrYW7H4bLoU/MdLeIM9gxnzeTI0lLQgTlIf9W9qQPlXunY2XDkyR8z+
HWILF4govEembJJHF3Tep+eT1skDslbzcOYpd4439daW0XgItLdxt0AfLne1Xd2pjRbDIbcUQVxi
DAsV8h8wfbIzmvpxhyB773MTms9Bx8Omm7iSDOLSvQop57Iio247BgnS85lJmk3xxt+y5kA3niBz
1DO82l5osC3SUqaqGe86jeXI5T1aS6/qfUdXHUCuCKenxLWAJaPMIKrX5+FUYlzOceL5GotBs+hA
C/Oan9jKc0WZjlGNtTo6N75+HjRew155IWxxrX+QBGghK8L/Nb/YgIAhC3Uyd04jH9aoGBibXUT9
1l4V30gWW6G98tVHa/itTlHqrQAye9Kkjnhp1wZgRthjrzuwIRzGspBs6IHNiNOYIKLeCMQ1B9s4
3lVqUV07zWdzKro/b0Y2h3nhPr4y1IWUkbJPnjC5jO5Pu/80scdQDJmSC4e11R3t5pKO4tZTu4uR
3yD9t2SYvC/vcyepJvY6Oe8X4KI1Drwim9HbzkIHUWed+GcV0KDs3HI9JzyLEyTqQ0Yp8MH4rsl4
uYU2LvdinYi6ypgnaQlNFgowGxh509kRmCR3hUS0bZw0YOhxJlokFktdrzTM1WAVgsT6gLydlY9f
Jl7Cppr9x1JCo58K85duemdqy4qvJw185TasIJeL9ZJiReq2D50gtirbE3UdWNB8Hc2OgFTwse/A
kl9rJYIfgUECGxPCYpZaQJ8ASDUqezHTmNduk43sCGBsPXPmgBi8BcpPLIT/vUIwahU1ObEiTIHB
vWfL3CudiEKW9Qat7DvagoYpnQ2PeSV7Is+lS+J8B9YwqjdBDiWticGYXZhkAR6EKRquvscL2xjg
jUysgdb4yhPueP3Q0irK7C3AVAKmJGH/HjsXe9bISa7KDweBy78pmWIs+/CWoAzSXXqlVtTnYIIw
gMY4hYbME2rRdPOqSi3IPq0G/+lJij5zkU1d+JD8ebU0K3XCkiCXBLSdu26V7ukFjZy19K+hatN1
WwjQns/pn3dzmc4QqUNznVnOT68w3f7dAYy6WTKqYskUXEycItNSRb3Nn+JAFRxcE8SdZ+LahlKr
Zq1XqNCELH7A0+fdr/wmt9WGvSYHfQVAzBUrezqK+pRy0bbqWTrU1yYCJHvkQYqr0t/oevCk4Uwv
4BFhX05TlOqTItbgJMLxHi2HEbc2ZqrVZ77KZo8GF+jd6ktuTfQI05JZ15zCjH1Ui7DOKYelt8XE
BAl6IQ+CJI7GaRHkwIVezDG65fnku2c/V8adqaFIdxWOXnfmYM3M1VTgM+weNgcb9NEUeodY5mWP
7co+4l1d3WBIO63wrNNRW3dgjOWGaqwSvEAdewxY3y0LhvBmVtMOLY/p77+ak1/oi1OqelANSnvm
qSyjTe417pKat1Ni5C433CwkeXVNVIl/L+js/F3i5lpcL8KGf+LPgdg4PbWHw2N8IzDNI4in7XC0
kR+JQ3VtfefQZQnNxXNhjTxHIVc3xylOWLyTMljMblnKv3oBYcG6VZe208QeGElpt5i42Acy94gA
KTBqctiQEBXgnOalsaTV6a0iz+fwiMHGd/cZ5xkcR+pkeIK4Rx+TiBqMupkENxlTtAaq+9Ru3339
72S/04NFQjc+D0C/pOOnRVVyjrxKVpeojz5j2FM7rcjA/XqhMrxreiBmg0FsMUtoeKvxPcpND+We
jtUl3My38L2GzoAPWSKbBbotU1ZaRgBNUMi71kMuOvWn7NNG8X89Hm62G5yXaPvq2PRtUGrCVj9A
91PesYFV3TTKGHCfWruie5aSQGOiVv0HEqxvg+1HJ3g3ekl5tetBncFmuaqf8Q2tn+VfjXS1rwvs
FzPxLkemqklDwlfPuXa+pAxgv/BSHkA7/bMpfs6Vzws+oOWd47cmpmn5l2TqiQxAsoXvlMdUXFXW
byi8oJZlhW3Zo7ilO/34mIYphprtAx4xyx02rKJd2IRVZdOl1eN7pHkYQwP+7gRSTymc2+Df2xt6
0QT/+Ak1XAyzY9tElJ6B5rVR2GWE9Y5OcpaSL0/Yh/0lxSk5fvNd//KuxF2qx9rSPa9voh9kcJ0F
CHEp8l48ajKZPofG5XECSeCj7VaSQokdfT7FMyc948Zw+aEjA2WtAnTR3pWCpybjpOEh8Cqb5MBM
t/+fp6oFHY3fc0FqZP8LS/ZyQH7s7XMGmejFnroo+d8Y+BPJWujaMP++9F4rYsP3jwSxmVitOzIX
jcPyWRFugOD+BLo+AGopx/yBiJSX8EWkcQkYHxltTNYsI3KPEJbt5OktAaTCLckauzVUnRLCq+b0
BBc0hQ/fPZAAmTPMBjn9q5sYsIER1opEs/sL/kN8QhabupFtpwOWAb6NUwRGdw4VTwbHmr7vPPUn
i/SD+bEFqH5fdZOMRgSaQ9vN2jStstjHCOP9LwSQBRqCitCmbgruXa7i4L6OYL53PF8qBVLeGE0g
I3hts63bELiyuWc+HuqK/rYMS+IshiY+ZXo24WgHlmg2T7YNgJLNVjaxFvQeD4jyWtG/UGsprKwn
RYqSdo2EjFjgxccbtnDrNgBPxWqTOi6EWRqSR5uYzX2fSEnkxhwxuYe863f3YcSYOCp6mJ4mMpg8
2T2+OTsuo5ZJ09Ic0NJO+SiXFScGZs5YpPWTRbYPANUv+MRFdW92lf/nwj8GR/lepb0MF5JKjOTp
SXbCUofYdtOO0kbEFoEXegfKbE1oPnBWuK23XCR6S1Honf1avIiXBzJmKh8d5GCwrNEYaxE7wwA9
xyHE8VS1TBpPpsunH2APyzm4ZaUfQZmPM9gTf2xH2HXL7x11vhZTq3txWF4rOvF3shXIykybxYz5
HFA13Rhyk5zhCxbiJMgCukIw2KOLZ62ly7oD2mj/Xd93IRzM4C7ItFRIt7IuLEdvph/wkLEPRdH5
/r7YrM5wPfZUt18wjI9vpN1aQzNhJPKMbptfW9bm4xJWoYAhtBa7BwOwaih54hZItiiIYxjaH2hF
3TYVhFl0AGPeBhThHKCtghgsF5Gops0IiF8KZ9/rPL5fKjzFvT4MqExiUw33aZUPlBkiJ0HdxQCe
c1WX9Ry3bP637p8KI4ABxE8gwy3L/tE6JuUViVn+xHm7Jy70H6vWfnzVZAmzZ8J4uomCDa6wsam0
QbMrSl+nO9WBGfJrqZ+0k2D8idv6aAAuZX/Mkv08+Xar9z/Zk7yJSNAMOuiG7F6AcT4am3UJunWx
otBbyuhsamVbBIZboCr5PAsHSCTVdniqR8FYqsQ151/MfC3uC6jZNESvMMCwuzBmtNiUh3EANglY
LXEsAx1O4oMJ99bK8+k1+UT+JHo3ks4jQSUlY0cVmTKKQzaU2fdB7VW+WgabUcpZ0EiTviBaJGfF
7QBsHKcd8VsRog81UVUVgumq/ONGAdmZWXzYAYHWlf5ZdLafNhWmRdJpxvLKdieg8mSMNf2ESeaM
AV0zWmFugvEYlOLB8dRdIbn/Gy4Cd0llvOujz6DSTW1i4WyJewcBwVQL1PjXzrVE+/dxeT41yLTv
JehuG9FbrlKKLntS/oCMCUb59pmtTtelavMtY+VznSpcwiMdWq3qeOA07Aaaud1dYi67OYlBlekS
kVs3c2ZDrLZKEFJZ37PPymnAhcqkTLnw5UkfBJ6BS8QwjhwPBZ3E81Q7klWeB/RGrqOxj7y6JPLN
XMjrSYs8pYIc2NZr1Qndm9vOun+FmgVk8ckVEVH4hZ4nJzxAjVXH6YBDrnq2biEAIxijZsGSUreG
3J5Nfeo/Yo6lIqoLIFiMP244ugZhUIYU8odsSGiNxvtbQDxTSgdR9wLzSF4mDEziqlT7asfCMOql
tio3qlPqsx5wFWPmjk+vHrqKLrDmlHi5564QGuBamuig+AYAwKZdte8QUugHHUPaI8FZdrw+KKW+
nHJ61QMN56HP/X475j4270HO2zupMGxNNuXzoonpqvmZWi4ujRDdLDu/bG4OFnbkJmawnO/dbSOZ
F8+VErlC1ltEr58+IQ76O5O7qtrl7R98OeThgNZ9OV+D2IDOMZtKCUTcGVrn49zLPXfZdm2Qn7ZI
JiA/91UXrGIAsp/Gi4knFUSjk1oB8kS9UCGs0sx/IHhQ+Uf6TkI8g8o6rlvjjC6uecka+xzTs+KC
rG8TF8ap/VuVwgLjWeSaXi1WM0Z4xhUz3cc8Tr7nhC9v5SMR4Xs0N0m7836XwWh4UtqvZ7wVowtH
fYEWEaUIMUfZUg2qD50b7HVDpXZBg4XioLR+RR0hObHah5W4La98QtaJ92KW4jejKWZtomPWDMaw
6iwC98opHpl8JKZifsdXnUF2Cz0JouFRhZxvvHx9hf2wfTNrSH8pk11I1A4DPQFy0W9vZ1zrCgky
Fo7jKxvBlyxaiTdF7qOViSU0Cy0edqFHfDGymN+jeYbnUFG87LhL9MJ+ZMrxyXAYWjhqAkh846su
I7/D4cDKeEQCp+BrHoYcdbRjU9fvtJD8GPhHa4hHMYweCqrXlrfAuYIr+5pbzxa4ktvC/ilK96ao
w8seiNHpv2sTllsB0lJJQlGxUJhHCcnfBCJW2PJhNxiu1R+OT97y1MkrOyVFzIvlCvJPVf69DcXr
N1BDk+7cr2daNNFlVh8d1wU1kr0r+Itpvz4576vwLopc4wN7oy/T6lLMm7y5FN8a6s7tQCzIX5qy
Ou4pPa65RLs3DaM4fFiw6wQTHQcraC8QgQgREXBifXBWmoAlqWXyfCDP2FeMX+8KTGaW7B6QWoaD
VUn28vQLMew8zXYP9ngBXaYBFDDepsHKRS3Fx4vQLn32GlcCg9rHQpqMoOeLK1dj4DmUFMFZO4jH
yLW76Kqf8Zc++uUk2UD6AxmyZM3NJWBzNdtxwD08cLyCNQbXrhoRukrcW+yfZJqGu2gRiCrMWnON
TJKHndqjbeazpnweQV+pxdbzneFuDreDM18VEbiCo24+I9oU/Hker2YZ/si6QcDIYI1tWuWhvg1J
lslIQ279827gcEZfOqdQVlva2q1lT4Duii1piIMc6cHU+RyGc2x4mTgY5Uy3UeLCmRTdehqFUDAD
N00rtOFFEOkmeWoZ0Lr9x/83y1aFvF50cbTrTGobQp/EWDKp+lNyLKgpxpTnQuL61Y6QPfRdyPuF
ieJ+H426lH+GCPdG9meWRm70g6/VJ7rKS+6g49Qg0He4kJf0uEgI/uWv5Rf65Vdyt34Wqup3pIKX
raBXtGoNG4wCkYZsoOIxKw6l/m2pf5Pm6AR6brdk2k7mvFahpsrYmZaHHxwqehfn8CTJEDAcbrTD
cQYwaUoGzhi+WcTpfsCpNXrb3uS0S7XvzieABtiKb8xkAusvhoTaejyuHvjNz6xV+7/skQOfGADX
WHFxrxwkwvoP/o2c1lMsvjv1xjS9I5dZcYCoNx36z4inf6AdHTJIa981umKPx8tRGmg2QYUndHIw
YJQOnYkABKO9QeZ/J5MIGFCskIiMqehuCJqZmyvdlqlkAcv6eHwcH3SekNozmRk6JePIL9vZ2eaK
jBx4541FAVjD/+RYQaxO6hwPutMnN7HfTSWhtWjtD5wvladrKigXJtE+MC3z4xevPlyv5PDvPY7W
bnuknMPX+Y3eD2QFLN/vYauqV5+NGGlgoBxT2u0qAFe5COGhT3h1Oq8MZS8cLICwiQl36KN7dyxL
GKc68tXTFOH6asWnXbIA04z6y4I7fFYhgE0WP0/hj5NeM85cd3SACSLU4ZdOeGIkpMGvR1svB5r+
CzULHKc48JmEWBV3LAkKSZtsM9fEUV/xRQQb2FX6S7b3Wls0v0FvzANHBydQ/bFxla+YCdg92SXY
7K07urjHgTYEJQWKYKAxFOpXBSjoBcI87y5CK1x9jOBEs1SblKsAXAqLd0SZ1GQUHEORV8Mh5SKl
IYR1IMQfyia0HJcU8fs5trlXcnI1/axBszxKAa3YI+I2GL0qPmI5SSXV5yJyhO+QATQhEVTKerwX
QNc6V1ggMHz0HlHyLZ6l0SdUSLx7kLge2J2ixOqsJlozYmlKc6ASv1w65HJF1CSZb5ZtRfL6QJGJ
vUVYBKhlaqZaJXmKz5AxyhCwHggmavkyZH5fvkUN+6Be4F+4dgWNMLgjEG0LhW0zyZ8DNnX8aaFy
PZyoxA/5tsv3gCZGR5gml3snHVBma5XaTT2xbtp9ezIuX5c2rBQ39/2g7knpgAV0RM/HKVl95ack
RDjfMUAU9SWXvdkvjZFqSGPWaYPLtyCio4GbE0o0v3F4YdP8pNlD1vsjk/e+beCBMDXir1bJyRJd
LvKXaC1xBXJxVMTXAXvE0euI0EoNfnbhvrxZRlhTJF0cL1QnXh1Pu95IMP0zf+nhZPHIwGIm0xAi
1vLj4HanvfDBAw3qyp7ok2j0Bo6S2azIs7kIXg5iM6sqZtHOSPfN8BkfD+MtKHMDTCP3MxTTGBMs
Fkho54IkPeKc6UcERWz7xKqf83oFIcKcX71Hc2QaaDH1uSRY5O0N3e1rWsY/kITOwFH7WjIoEf7Q
jollfnTX5S7yASBO9rLCEYA3yPaWMPcriQWpyD6xvHnAzina4GcB2X9CxHqHOzwAx+XBlrrTf4jl
B5GD6qWfvAKn26d27De1E/xoD6R8yt8Udz3dFFKvQFhSCoxNaS8sqST4oT6XblVfoUGXdMCVmB8K
ibdJM9cM5ivAKaQePWAKAVAmuS07YRnpk2yPVcV79eLCd3jWLSqPcmVMcrwr9dkCqsGI5ECdIF7X
eK7DNE+aKhPCOKK7yIrRSdBI0kUPYVrDx7sx+3akMXKXdXGJNA5uZdOvAkaAJT2rLl8rYvDv6bLx
+OZrTPkhPHBaKvLMMhoEryRmPrZISul6oaZlXF6IyJeyBgPzbxwuvu+TvYP1v9bfEbLeqCjltF6o
0N0hL1dnrP/eeQUHzBwUdmDnSJsYgAruka0yfBrisDWj9znyFmdJxyAKrFlIN+jRdFp1ywcs5VEA
ibzhA3dxiziNroQ/7urE9UTq3Q/yjBVIj9h0A8tz+XE2rwHHpMYQ0HCmvo07HqyxdlEDYicyrt2E
VVxfWEVVcU0pglW2M2auHDuOFvtXUF0fUqmAyicwNhRPeEZ+6tvWsLrx0jlCTLMF+rCxwyAZ/kjg
EsCQtz015sB4KO5Wwa1oG8n0vZDTAAH/JinoEPEZ44aib4vlq6pdZUDmV0hkHbdjEyvOGsVN6PvD
/R7FyEHNeXu0Kks2PVH9ZTBl+2OIbO29NUPPPWORXxHHKY/6qyPACXwKDCyDpmMsbbHcJY5t4ODV
wqXb+5cUJVrQ1FDk4WRm2+cSgApWt5V6SspTt/qj6AdOTtl3zRFZ+ek6+Gu2HpxFH9Ysm2JlL2xC
B7UhqT6+ahVw4is7D8YqmG0f2N49QOJDTi8ACZEnUxr47Y0H0jUXfTI2NmmI3ytEQMj02cGglZe4
kp5ixcZQU1CNWwNGUwcJrs//u3C4tdx+ewWIiqmRzMVdNL1Atvjri5un3V7Z5E7sb57AbJF0xCtx
ZbtOjeVm62zpMTuypeSE5GovM+NxkKITJR8hZra0MLlybKWCOkR2UltZ3FaVfX/fH5MajT88Np90
nz/m2RUDGBN5eyKvy/bLFm7BhnUEAdeNrtbSa+bQ4kg5FZHiLmFiwOd9xg0hDrU37EpyF+I0sgMO
49vDRJ8mRd5uFGqdDlb7PLeFllTx5DHbczlAU80D9UXempSf/73TZQnjUARC/+52CisClSIv3Ige
kpkRVU3XMJQ7e3JnizMhHDht2yKA25lwgquGhoj0VMljIqeMAkbkFs7ANqwMx087y2+4gb7FMeWe
jQjmheKP2U99DwEb8M4kirVLTSH1TnkKy2u4YWv0Nhjjq4ZRq4n/VIpBvqgsd27c1uexJ0YP/dis
+ZcbX++5Rm5jO8yLwUwA2YI2oLkDr6N0S/IZAKS+a4p/NzpZMdI3H2QIEVAzwhV0Zb2czOmgnrBm
wJ8enYWrYo5PjBp4NGF9MlW5+L7BWByAUuEul+0ARr5Ov/nkAXfV3PfIlX8u3gYL80gsjiSJzKzH
0Ridx9gd3aHXQ5r8zx/TV2c8JSJkPYShag+kFeY1w2R8LHL3rpTFsNBuQzZo6PxHwmDiaGkB0k2e
rer2P52UnoHfq9eIho9ZD//YGQlAuf0AO3HQyEQoFOcg2eQTL31ZcSMOGqpD+/OVH66gev6CRwK4
HEFoXy6wtW2TftZdfrUElud60f6ruQxMwTEniLjSgKLDg2kVVtT7N95jnUiYXUtF30gwPL9756Cv
l8+HrqtNIZTE17EwMsij5YrZC37v8dFt0lGhwFn76hxXpx8XP+ldg8kSqb871C/BhR8xpta7i2ls
cx3g3TjyDoDrU4Y8HLBjTG74Eu8H01rvyXEVmH8ul3NtPDvNIQqzHXm0rA2OC2V5lgxX7ykOS8UO
2SKBYAcmh+nqrdTfUidGm3AZup7TaKmLHP40lf6aCdA2CQ15b7rJrL40i3FNzuR11FZeEZz6yTHh
sn7JuQjB0u2nX6WffsLbCUUfkRDHMVn+TosZ2FSO4Q33Pem0eil4U0tr+WIFu2+BDRBH0uq5HAdA
+CC4U3sw12OeWB8MLkI/slZMJWkuojv5GjurJkBnqV+q1WQ/sskXbajaKJ9QpDxFdYQy4Kb/NW+l
cPpJUtUntYbHS/X3d+vsMrElZLN+XNDgXj1aUAgE+4krd4yYWOxKEhaM03r5tsIR1C80JuogbWM3
+pd+WqhqRa4YpBOw+fEmdeYb9HSYSLt+pMEha0cY8ldmaVp1qKIa6cDTHd58EcCj1y4/8xYtOA6a
RdzIbzqL3QvTOvpMw0c/IxJZfhEhCCD63PJDzSpFLotbR1Z8UC0Yv40NyOwGuoosv7QohNmml6m5
ARX73O5F/9i/xzEgrBv04yt9mobVpV3z0WdN6OsBIhyzcPMTVSoDaZkA9rS3cE0zv0VafAwLwcqT
FZFFlbUJ52LPrdzCqhohTUvvSUieFjjNOGsfGwsFzv/ybPb9agcRjQBXhQ/GWNl1xpqp1QvoAgsQ
VMh3LKOJzEjDD5pjevKBz+rwPL/IvACiki6+g9E0xLFyu9TOc+mJRM9O7hiFdTa7omZMUFHK2MD7
HOcuxqzC3k3eemsb2o7j320INPVlqYztOu/wwCZlMSXSRjLlOtUit+/mA8u+AuSdwCbOwlWuYH6k
awCB4iIkVDKFQ6s/brdes2FL5dGH0a/H6b0/iMSiou4ZXxSfD+T2Wk+ZM22uK3z42H2PTyAEsgca
g+tskEbRmnlYZTQoKIfFCS2Irp7NVlUSvwpjFyT6qW2v0+TN1JISbAvXU92YHqNKncv2dNs15/AC
ABNgxi3WD3xcHp0ccrkN8zJDwW8LpwtJjDdmDFKt2PVxsVo3ZLcBHXt3j7abo4Vn/sKQqtI+kNHV
KubDEEtbn0e+e258+YkB+/so1lojeN+vgNLnSezlBjPoKONHqeipviDXYHg4d8JZU1ERRTLc4c3E
jjKaM2R3uRpL5itpSBkDrGT7oWkH0nUoMQPzVQkJy0KU2918N3W9M8i4GgzrDjmck9ufQg7Ow0Y0
z/KbNha3zOUkFpTSWxftQIcfS/NNTGlpM05iZ3BJoVS/k9d4jKyyO22kweItHybTf+iU+0OPmNKI
Ag2gz9N1CdQN95KsN2QKHSN85bZ7ypqlDebNq6PRHe414aQw6yUQ1Xzxrn9n8Sk64ZVneCNxIVTl
lBfdY2K1S2lgLlekX5EgONgP7Zxn1y+GILZB2qGC5t5T0NUV07M8VYMQukLX15aZf8X230dhPoPJ
pYORxha/y7OlJctFhKBEQp4434IXn1WWRjnbQYnCS+1zxZTbpnBPypWgIvJUoD9peCJ88+XmkNDW
THy/zCGmYm0Lif96A2tC8YffldOXLKmxZijJh3asLA5FdDHxdLpx5eJnPLa6kGTk3SO0hSvcbLQE
l8TXIG9iRv6/UARYzUC56E35gFGjnV6GlXipxsNd9y7w23nl9VLVDZN29gZS5skDyofs5wq5q6bV
iEXwkM6zaNP3jJ7BI4ebAiqqqgkx0I59MOIRdF5IcrT+oPQg8EOiLobe3sicN/gbtQr6lSCzl8IW
3q4r3hTUsSVW8zO/1+mn3MkBnmwVhhQRM+m/EwgJ1J0Biet6ltjR5uSrfJU2G7oSRsW/+CRdlSMe
9UV45Y1nMJlZeDnzJ9ZXsqGAUvOjsPSHXsQKCDVhHcdzE2cstCYasKKwtJoVR1HUmeHJgCS7yKgV
MDV4/KzwYhfqTybZoCCKyN+EmqKPcGeVbXEWIcGOgHZUQebmwMsJKiEl+lWydfoFIFd5J19Oye3g
96TK5mjU6TXwh4ArPuSKkDFmFtvHKy9HOrpFmuegb8/KH7lBrG1vo/TYBM6w4U10wuuNRLZK6ICZ
GA4WQhWTTsxu4lNioEhKXDXxxpFJyKD3S0JbFmm9TwPoZkp+VZNVJJ36+xk4xaBVBzUFQxND40Q6
Ecnq82ab67m+qtk2XG68bMNHhmdsewqOaaMTP937lHeVwi/0hGmXn9TYzedmFW8P5QQhHrgovTWh
OXjX4VIfrY8ixHzclio4uKQbZ1LleH46IhaPEIf7SwTzlMmtBIx7+3syibNyRAwLyhs5QeEq+a+S
pqxWYvO1EckmfTzN/4oY9NnV574Kapzz4r5VN7af/gy2Sod9h565HqBGXH0LB0iyb29+F5N/vGGL
eLr5J3ybrUVqziqWLvwsFM+dYU/EqR6kHQeCC/m90drZVhHPklyrja2RY6pg9Xc2qxKce/QInIay
SiR5gHGD5kbaEi7Ktxi3HQMGPCeTnnBisY35sdwogbAm3kqKVlXwkgOSr0NgsufeGW290xxDsTep
HY2bLLjKEauW/rpFjLF2iXoSjE/F89bPWv2mbsSXpLPgVEGrmS+cXBmqd5OyxyGsk0JPSca/vF3U
z+DS/HNRJBd0gjd4DshcEmaZsuQT+6yN95VLhMY+ffQ2K8ql7bECSHXngqL5cB3pVZqqUEALK2FM
jevT+wajJ15hVjO2dTwFDBSO4gFNj+LLClDoo6c7mCgr1ktYJ0uFg60QkfxjAFrIGw59pKX6AQw5
00QTVpHpPi7plyiH8XCWoIYBEnZndKv4H6/7OWDjDxc5Z2EeRQtnDV4wLIGr7I46OV0mA3UrsNC/
AbZQmD3jy4KCai9sUaZrdrt8Jr/wqs2HfX9WnKNrfzymwC895e3c7u1Re+ZsfW5q6eB6Q6ORLJ5x
jX2n7fWZAkiIBavtEcWEuJUzq7keg8SuvXkHg9Jz7P2XnGsQI3qqjpb25CqTf7Du7HfxiUzRmIza
XzmZvEAxrxu9NVvcmv1HBHzO5LQFfs+7nI7yHiEDV3renyilbLpguPk01ZbJeb1qyyAnDi1MteNn
VEvPULp33nJ1X5RocCrKXsOIp6JSwmLJd7Nu+XvxHu39J3rAz3uAVwsVN/pClCuudISeeI90PJwI
Px4LbYKNuXAv/r4C8NB7v+jHLEMdUFDS+4xeoauCdut5CCtmSQ0jjnCeiCeBBsANTovspRjyZdb3
YF3z7b9l6HsrE2Dt5GH8ygYt0h7WVOOE6gEUMKpMZ9OopxpJ0hlxAOjxD2QX2bsdmVQzzo4ip73J
CgUTs5kEmu7eaTcUxPCTABbQKEEjydV+T9UBgtwrx7AjasBWojoK+TLjQA3iJ1Gb6h3QICUgpGWx
OtqnLR/YscjFsTzLhWPhS5AQUQdcixFjHiIILWU4yplsvFUNqQOY02+tp4sSx3/G3lxfhVhJ3KE8
zC2qW+tnY+kCw/R7aGWzWTQBL9wd0XBo1024u7v6ovQaW5FRPK8jQXIRDtXC5bTjbRo1wVEHjS1q
YcExLP4FrfIFpq0fRVG2UB0XAuO9MlwYycYjejrutPVTuwnu7SwMvIl8t2uXf+e1t74LjhMz0RAD
Vn4myrluAFzJUR0c2/QTMaz+rHF3PRPHq4UE2oY9Wuq4bVE1I4vM6tWFwudfj3Su6TO9SoWFtWbl
xXCMqSMJpWbRYvbhq82NB2hTwPy9cZMvopLy/77iQAVeMZ/txgIHSOwdvKvsZgVFUs1KBBBXfW2D
3013ZeWo39zQtk9QakC0QvsmjUZR5dlQqpQeF1JjNiM8n4/lwbdVdwqfBWtl3JDnDZKJlEnrjL9v
xSpMXdS6zluAyBt3YY30Uywwo76eWoXiGv69xKvCdp+MalOIUwfAjugID6qTOPpl3dxwfwbnQTW5
nOpFqIguZYHByDed0jPrCN3duxxd1bqkqwHGrYU0+xx2Ygi3JYV0VaWcijvW8yvq7tZq8KuSAdvo
YW6s7FgZxJh/O0h21Q9LRRas85weWZ8TLX24NearxgbY9SyS9un1xTbs1pMnQQRSm67JLe7hhZD6
ubbJ+YL1Z1kq8Hx0+TvGecXHZx1qBH+TiFXcfAPfrw0c4DHtxPbugqUzbtWbYMTxMyD/eCmOiTjc
nl6bVFmgb17KW+qp2iwC97c4yvNIXcEAdvOOHgNTHwHDpSCzMqKLstFtK1mOJH3SK7ZHpWuTRRh8
z3RcjuzDfq9JkReDTeSI/Y4tXg8IZCpc6d81Igid03nRvt8TrBbjn2O5h1LEx2u6xvTH68/PVkt3
RC4eSLEpyEe2UPd2Er4PzAyRN7FPGVLl0Yvw9K+qro39ZGr1ezyOR9PL85+PSVEJNiiKyLsSIs+P
rik6epaip3hBLd7Ysukqpm5/5dHm9Woy7HWpXxsjXPogPkKiqgbtow59X3WnTffr1qR1cOU6zFy+
qbw6Eyl+O7DCN7HiuRbPVv8nwX5A6TwGOGAUurcEEiDshH3d4aDsdS7t1jcSVzcYevvsaDoxvom6
5YOTw4ElvK656MkCbZhahHfiGIpQGYPibQiXc+XB5/DZkXGEZcnsCHzb085K8mwU6ur2Vb1zBWB8
203k/H7mrYEb2bjDigMCjWBZcYch4L8U1DMQIeVavRW8FE4zVypNZ/RQycC7oockIR95c/AbHS/y
fs8KHoZk0/FbGOKGdtlN9nlw5+tkSiCUM4sgxZgOtses1VCFC75qpdkZKWAB2UK4alo80LPePhYl
ZSFNtichtXlH6n7x/WGLhALk1kBzze4JgG3s1mYohdUellVrgmOXicXak3TKre0nMx+kD/7C5T5f
0XgdPixkb3J0Gx4K5wkIwE3e5sfyDDGuV+au7H6w5lLnYTb9LSTl5KBzpWz22whl7XvvOM8+541o
9yobvS5z6EFeaJ5Qc5CilLkOpEFpNhPd6tj46iALkYNDShjjmAgU0agCSk0eLOciGyu1xaVAk8jH
xt8PZNy5tchu/1baP0ltGJGSPFwOZwE97F5WH7JXwzN9DOuw4oZWjhHjP8xTC5Zw6Hv50WI0wsTg
Ucmyr8fRFeFT7GDSTZzrkGnFggIAuz1uz8raYndC9noT9zcxJyG/Nd9nmHNySj0+cvEW+CejcTqt
z6PEFWM6Mm5cXCKPMjItZzZgZjis3u65T7AsalpGs2dl5Zx/UqW4Qs21g8P7Pg4711BBfiIVLFVa
T+I/ofULdOpw/0Wtr/QBkJ9Lmsn7VkrRhQSc6Im7DkcREBxOCTl5J4lWMdiZkKA8fYicD9cK1pwV
bytSXigBMmDuz+qUZ6S3sNXI2aa30q3dqbFUG6upoFMduf0FZso8Ks4HkZqFT1/acdRlwxIOMD/q
LdQibRQar+AVckQIVBDaA3eFTZWUNxLWMHMIWtxTTL85yV8ciYBqa7Td11h7czLJ/Ja2HJ4cBWPF
hyN3gCiYWzOMD9ZFaehpP9UZQo+tROk+aGP6cNjlWqs70wtCtRMV9iT4PSNcL7jCAOUfsmRPBohq
2w8lLzAj7XxEmxsGTFy93RgDbJHSUGDGHfKy4XrjPb4PCGk2II1mg3oK5feFF6zL9GZkQb3RlOSl
fVqG6EGrdUCJAP66X/6OkJarxud0jdJo6NWjd66EAqkLwdTF0ZgyOIkY6++hf7SmOHSeCcmDSDCn
X6lJCxXkJVcSREI/z765uJcg2CWyc/FUda2RIz2J0ZiaG/FYAtbA39cB675ZuGLsygHNEQ81xvB6
YmtRKOR6veuRyqIrd16dJxp6PMTF31mliybtEyRihXaAgIcYKsx7wkWGSZ4LaD0aHrie36a3rT/K
YoND9V4Z5A0all/9+Rr/+SvRd9d9fgDe7HdcinSziYX+L7yvTeEJWju2NrLibb/UG4EZKceGml/u
QTkVTatgXlElFAPX7L6cklVRlY0Od1OyH0c5lw1VyEo4eKXm+9CPzk6Qp/OXfQyJIqiJXZZd36Qp
j2rsUjWviP0UpPwWSkBIXgqsdjWhEv8CyPdnxsGTgRDLlXKTCFhzzV4jJeI9C/MWeIdA3nEnogIl
QK73OyjdmaqfEl8SIBNwN2wlnJaOH76TTEnNN2tYwxgYPIZ8ppZ5TE7XWvpzeeGYYN808BcDze8X
rkG1/M0yFBmiKmAnlW1ycapNgSteVH1NMcfv/MoaNdrQKzbZztzzOVLcN39l8UvvabASHZGs2mvQ
6WZstRQt00N2ZjtH3iftSE35IZxJx+LZFAESxZgon/VrJXGyKCr98lapPX/dytFe6I1ug2aEQX8f
HWUTl4QmLEA6WmmswxAgkzQFephMBhXSPNslOcXE7S2iQFHDNNP1J04kiKd9x8i0dWnldW5H5tsY
6YjSiux3AnBvUXHpPeEgxq5r9FWhQehU/EBG/4Yz3mpH2Wv+At7KwI0zb8anoJSC7JKlKWaYi2lD
u7zQPMNl2y1uC5yIFIjuPNcoc80T/zmE7Qm0xA2UwgQPb/R5BYo5Yye6g2elzyglzswWoTcq0rbh
kkMEyx1eEXOJ4HDsCQ5H56UcT0NpPBlQd0K1ku1XxA9BUAfu9YSc70sCCfNVTw65bjZyxDTFYyjn
yVmxnN+CYDMAcSApi1B7FWV97uSZCwBoCf0ilLzC3Mhc6hr1tbviHMXvSY9LeJnWIirxl/g17Ayf
VW8wgbX9F7WdroFRN4wxiGlapw52dS9WT0asfj3bfI+TFnRJBatIq5BH6yEBfJdlDgiKHQjfN534
lr4l2LcN/XwfFerqLwDgFYibK3OlOFGVhPHfzVYm+27JBGxsRE4HIf9YzonJXNo2fIbXV9oTg50I
L+Pbsg2G38Zmm/vvGw51JCd+F/SaRchsT/7EVx8yyDVTNrowwIgfY56knI9NN5L5M5OKDQEA6Yh6
4N0BJBIrT+r2RtWkR08fV5wYciO4HEEsWFkHr36q8HuY2DDQgmQKJboCf9xMnSIRA9EcLgBb14eA
rwTDoX96jdJq/h0MJME/IRfl2au7fTbEF13WEnzy8ApqWStC03zJkNbkwmovh+hmNke0bgARoaYZ
ZK/OrDYbut6tEZHjrXPg40w5L8zuRmcvQOvt4tzTD5lJ7GHBNIaCwtl43I+G5hM3zMPR+Ho0dhk/
7fHS8mGBBFRNvHnKY/vVe23fN/adL+fLamGxy5Sr9UvOekKr3FHQWaufOTscogVyQAYH9n5H5ZbP
/RC/GVdDRXF/1wTVV6UFhnDn+EMNhwGtW3xEkV8NohW+PieVBfpK7FNOc0yDBo8Y64NP0zWNND8+
Mjx0JdXWCH2i6Fm0aMa4gMfFGZwvBFKm7wDeLRLycAlzmb5qtBVup34tX/jE/4Ft//bT3nJr9WJa
go4v1WOpTSa4EL5IMUVGo69Q9dteOL/0bj2gWDSLOne4eWUvWuwkIHdKq/+8iql9YTSUWctYuBVF
jlqkd28L8OTBmFz9skOimln7n0pfjZFuZULZdYXc2fWChuv8+4MYVXx72/UUK0V8wydQLdJuGFw0
PKKTbBbQBoNQ7PxUVHeNnwablwyia6usJiMGfrW+a40DwOdIQw9x6msK/Wfcy4O9/AuRoSbFGHVu
CIQ6L5RTMU6KSwGXagh6Cg6qZ8uMHRIda1BUenccQIGLOrgeoxYgGSZ8Sa9nUlLfn2YesacQpEnL
K51h1d9x41qdhrXqvto1z6jXvUeS6fSrz/syOc5tvNm8JtIdHCv0HXzorDi2JcydiTL7YjxXzi/M
kevITKxDq5gY1gX5LT8gCgvHgYTeMZCVCQ+uoyRrBlqPjAK0yabfJjl0a1fJYhOV76kPAV1lHVfZ
yisxKmoxVXvz5Hz1/xB1J52FrKD6QyNVI9ewEMLsd7oK25tIjWRwZheCuIg+Yn84x5CL1FQv7bEm
Gvhrv91hbGiMZ6AMdwkF7+SbAZUw5zMAtIxibsOxVa6KiuWDjUC3tIaJnLub4Ke2RFyjcf6q0iFB
dQyrCROSaSfeAZQGtA5AAnb5UZo38r2MOZeJosYcoOemKD+SVp2N/j8zNfrcGqQM6Xnu33vzxL4M
dbcCRvxnoeclDBxtXA00hx6mdlAQ++i1CSF5V9q/svFBQOgLzDGSsWHpCohrOLmRIHyUYAZ9k4YP
IEX8g5ukSdN3GjU6qwMvcUQrxU8YuWfw/JmMR0Hc5fchGe6WNd2xPD7x5p+gqvdIEFO3bEdF7VaH
29MMZbOkHFXffLLpLQ1gyraZQJJxMBNUKDGpwg2NL4N8rJE4lFaGFHLfmEzo19GOoplW83FsfIKk
sZ8MoTWk6ombKDB0WSVM41hMuf42Dfu3ZjCjnmxvbnfAKmgwhr8PxpCVthGHiEYC2FYOEACzOchq
D0cWEJhpl+tKiNhyINFHmHMB3SlmcagcySfc3mFfA/4z2lP6nCYC/pCtIEt36hv0pFL3NbLQe5NB
7jlNQtFOgUA1rH5t5S5wbz4XD20MvzBhmul7z1KUsdQQTsom6FJP6bWG30dDv9DizLFcUQN2DY6z
pQ5FgVG47gPpKHCzdjveyIPv0wMCcc2qfEeLf1zeKHKjRUoPir8Jj/tAmuQFZEgLEuiLxFn05Cfr
6tFvvK/qyXlQjS+BhFn9lHjI3fkSyafv1J7ZmwVtekEr/JNo/n4f36rlZFZLVC924tqbi90P13li
0kVj+T7MQDXzThhEScfc4xTUFsofbXiJDLmy8EAruheCHBO3DYvHUX6/ZG7pxl3cHGhxxtHMszTd
nA2rFlQ909Co6zYT6akbOy4NPPA1TyritZ+WYZlnMcQGfMM7dhY31usk1Vebx7BBidiwQHz3/rQO
vSmi1kKhA+/d99ToE7WI21s6EBcPDX/94X4HFZUSuXXkURJYTkKjRfQOJQxs0BxGQSEI6OwLpnoT
T1wg4VMv0g4CLUz2qWdL9V92Xrx1UnqNJspaZoJr1H/OyP53deH42B3Hg/obzwGz5afjbneZ+wtZ
eYXqC7Y5drtOOCHAi/c15md6GcAbr2uv9Om5x/LoOAWhWxCsuBnFeQGAuAzq1VFgkDZkFDevJDVi
0JJeTsyWsv07fq/oPxNo7txx35Uda3EyM3gk9xy7hEjL71BjE+JgX7qf6ARJ9oypEbAq9IrbRggi
pdUvAvdWqJ7KqB+PRrajXzl4lvyZfW+lBIpoIdPyVC3Uaqp1sgVhlUkghDyhjQ6WAHns9QXy+zWl
hVULz75+CIu1kr3RUJQ71ublTYihwQQhTECqs50GVvPbStTlJjK/ZlwT5sKQKeuCSJGiIV4Y7X1l
KtpL2B5uFS1k4Xz542ohiaKycIkZZpNHIZFlm4l8jWOnYeYD9qW+SCnfvqGKyS9Hi6BpBo3SRV3w
sZ3OvmNUoniPb7js0g2AtwlUNvxzosS/NtPvJuT14lRkAog3X1HglTJRu31hqJHomY0SYcXtNLJ0
IQFS2e/FW5cg6FpGveiQLyUjvE8cK8kP6Y/SHyrtLhuFPppnzsxI137mSDcDy+JrEuQlSe99dBy3
eCM7YzadQ1XtDNGDr85RVYPdRTQhDxiFlj/7XXymvXcJR3A1854nR/hF0yFf8s7DlQ/HmIdxr4y8
09XKHlGvNwQAfCFvS41fWvuxtoROg91iNnE2+EV2d0/db5sQeINW3Xm+xxq3tBbb4SSZbF2yvLm0
j3xzMhW7IqG/QzSNzQg2g046CrjOchPS0a4z9x2gw7hP7VXGfnOgojOnridNwnShHrYAH8cj6pF6
x61rMveID3IbjAVslHBbmWsUvk/IW3kaUyz490T115ZWBBm85kyU9vRXvNrzNLUXceA89xlxGKLJ
uqC5S+4Pph9lcH5oDa/ImAtyrKHV/oBPDSeCwzHXxQUwJEJEwMsL924lm378/zcvD0BqqBN3cgHp
nNjq9S4HAtwpm3p4OrK16OiJ9j4RLT+D8GupJg3dxgp7rcqLvRaIxF4DIX9PNIbRWrdvSEWUvjrQ
MGigxMc5eB/wCzYXFJtzg36bKdcSHmNIe/JUEtN+AwGgscvCGeMV9EeAxEZVsN20afru1Bl4ibEs
Hrd7FzkyUkncQ3KeAYdLD1iJjUA//vr3ryhmSCLL1dovvsgsncmLLaFNmMPm1XuAmt1DBMChrjrK
4SNI6XIAZzXL6cmvc7Nkq/trHbjPbkmfCl1by0QrrshBeK0UUXd5+Jm7eYh68tSmRiFCSrlIg55x
xH6av7OjJsdj5+Cc9kxTD1MCagiTrTRXT5rf8VOGWUFg+fLcES3Cw2SPoXnZMI6gXDPcuYyhj5Ru
G00SbOYcpFzsF5hlGa892Sv2kSD+E5+JMp+yhXLebr7o+PhwFDQ0QYkOLUI7sOOYZ7lc7wO6nqq/
Ha/Pr8eiSRXTiVg/a16AjY+SKR75e2sRrHnbrXOMX/61uZGx57g4TJf0hAyJsAHwQx+SxGSWXlUQ
AVP+QhNgVCnkQ7bOeXhnWUwT1b9VZBH9D+gKQSINEnn/ipXAwixa5Quq2LDubUP3gLWizSa5Pfgl
DpTrBCvRDRb3+HNEc/v+iGGAe9r/6IYSSS97iKlTM/7/snhYWmvnmBQ+l8QYrPmCiK/c7GBjwCmn
7znbPKyIX31Syug+fapQFzguDhL047V14shPmqcZc9Jo3Ven+QoX+dcmuGcZllJ2YOpTz6alX2lN
h6i4rc+C07lBSiOoIdgV3yn3LGOcfMfemjuZoJ7K8GheqpTpazXFuYY0CRUKFxI6iulcYE0yz+z5
IKSAX+lDI+F1BiDXJZSi8EnwUVLH3y7pA+LrbTiutZ3SSFok3OsCKW2AtMmZ2LYD/L/9ivzTYDNQ
P9unPds3Enkx3IjWrTaPLjHv5pCz3chvYzWtHcbTUxbmeXK9ADj6A7h0sOMjnC3SfTFavtm91eJA
J9oJFiJt0eBSGbntDpDqkngrEPpTXR2/zRYj6RAYuGPEp6k+YmzHiSjWPaTG0AntAZoh3e4E1RQv
gyJMdn4pjqThBB24LjJoxD9uMIzXEkdt74VULOgdoZjZqmePcwHi0uWnYEHgJ6qp9IkXjSnYjV3q
9s+LijOcnAo+0EsNWK8DVD96J2fMqRO9KgssN5cU4s/emeiiBQwzi6x0AGkYjUeHlbVJ+ggcsctP
Wui5I6lBoZvw0j/JUEpvdh91D/nVTO2t4SQPCPLgG0Lj9lGvYCUWtGRBKjxL6NZPYSmDMLgAD4Gq
AHdt6NreGc+b0AP7uNwuAWGddvwHjjFykVcAshNrvmMVLW/Fj6MAp+NBC6yD9TBwDXm6FbOqV+eu
77s+1a1qbo/GKw6VmX/sjosDsHOcvWHaB9LCfoa9ewy+2lsihdvgCQjR6AOCp2TlpowSrC5HVOBq
UTnDyFW78STJPRP/T0a03zRpUaWRtJUYHRtEeIYX8Q2/PtcDECEF3gaxEh6K0MyFYNI7bQXiG5+C
/eHFCkEeBKL1FDNBFeBnguBb6Ga6SS1JQea1z5gmmv+hR+I/jOCxfAmwCDsM/hZybFe5aDz1SQe7
pQx46pwbDMEGo2BUgpjq116IlV9YhRb+O0MGF/YThjNyJJbcwkWXaCdSeJ6KNFHTaouZPXo5bbGg
x1Cp3z+jNAhaEmv3lJgAQvsZzVyv+wDz0SmrSP+meMbWixgbsVNS1LJ7qH19MS/VwPbtLKAo0VOB
nWCjIv80/vwjntpKM8edEbodnQ5lvQiHA22D8hiww5XmiNljJdqo31dHxOakeKcagj3Crv7O2Ary
XaOnSaS4BEM+Gy5wsbIJgYy+snmU8MoK6zdt3V73dqvmAtwXeDjPAEnLSuc7APGdYyObEoOgoXu6
kS8noPr+4kpiEelVfKM815uJweLsGmIKxK/IbTxeN9n7vl8hUEiJu9Djr/YuQplNdcaHy+dfvE1+
6keC8EV9MlX0hV58Bae9ubUTEvvTaGCG271nkHVxvskVoULWCPgi0PNlb0eMSUs+ZYyGUOTfurma
PWLGWPw5IQxO1bV4pLZ8s2OIN29lqneFYxJBoWo5JH8zrHMD5W/wBEOycKvck56KuHdFaIg29We1
A0M+ftmu5DhKVxPNgjFHgIrRBKMUUo/Gy8f+VWcKjzx9veeYES7d3KMahBbDUIKrfYBbO+YRKTJq
3CpuMCgdjQatdbUlNStspjX2fxc7CjLb7o5PKlOnVoFOeJfbbhwyb2U0FQ/Jb8Girfx5SyGCNDZm
3IICQVJvBibJ8FvpeZ8/SdG6Tc5BDOSXogF43SG5I2/Delun0UvVILloppWm/4oNK0iqzHcV20EL
Af15LVoNsioMFn81reW/g/n7q/BGEBL63+zOs4G66wdrEe4N1DpQJGdS/zlLfI2Gt4VYdu8kOEPf
1tCNAdfMhMZpV+zPxYVZKrjv5dJYZEb7s++XHxTNduj7yhHo+W0Y4FGmGcUM/JeGvMXy6WV3xoDJ
3j6mfJ17BvyzDigb8igve5s9GveFCaeGTcoQiwmMqFlGJymVSj0Qjoc9xcNGSkbTZ0IT5Hr3M4ba
Ycgv3pNo/y2cf2odHY3mczro5uTSayMZgdVx/DyWdTubINTeKrsgzWRuhp8ZeZJ0ht0PsfHN8CQS
V/1tdejBQMRDJdhWJioZ+AXwycdeJsuiKgtK1EE5OCmzMhAFefY0cONGKRK7KmTc8t0BEtSYExZy
ocsgOqfQPNx6NsA+MozTmdu9K65Yu/isc6jz/btf2JeEsgNZn+ZPDCi5hPZ+cKVMb/vieOG3QpUX
186+BA1xNciGKGmciQwWqJWHaeKffUHdJuuWD8Ppkgz1EoYlRb22zZrQtacBrju9/Szi6bbaejpq
CyOLa9RFvQYLGRiuMQu4CfbcYzIDEWMVl/r1t84zhfVKO7beB1xexMnGNRUlIzcD/lwIG/jh7Eox
8CSY8BH2hAbV2QVCbhMk11xgX64OjrWESiIWmXZQ0+ErXUMi1AwGL9BKup3zF+LdRGXasRRQFSLQ
DKsQqgsfsK4o0qfY7NWHbveiQ75wFlTeml2QB0FqAhpQ0URtphFgPClPB/VQIdY8oi43/r1S0KaH
QEokDilo7Js1QcZgUtU/rymgKvkPbJDCMQmnHnKKYvnCT9dB24XTBZ8VgxOoTAMOupXTUi23d/iO
6AAWifJAKRFbxvUJXlcDwmgrhUAPFCTAfNQ5sFOP8B/8rYDO2hQnrwS8ZMHDQOmDnUc+K6cmxd4m
WsR0IT2J80ruFDmj8h8VXoNFJnfDbvwM2K/Rl7HEzI4LqCmagEu7ZdfSYTTUw2RMdWzTJFrYf4Bw
9Sp+4962Gn5HJ8/2wDsgSuC+UoE0idkBormONmDotwx9tKzIlJlpt8Q370ULPsICJLHBme70BYiP
dp1UJB6K810yaNe5jp3edBmbrVE/iy4WF+pOqra5wULU+XT77difb2ycNc9WertQh6FDnEugGsHQ
HsTrLELeR0xe4gNyaX+dGoqE4FUn2Yd5wXI55cJNU1WV809m5DlOaCrzux9dhNjPr078UIr/65sO
OySwry7I8FKttqWEzDJuiFLhMWnjadcbMvXMpf9dyNWzLWBLv+pa8dIJnnXiylWz2Q9spdMYAvbZ
JZmSuy7L2qX2rrjQ4eUsX19JmBvFxlOGubG4hvQQPRsgBlYZ4yx3/m7XGO+4Py90OrOZ0hF+bcHK
JrlZEAs92GswxrX45alYavcHIo+blZmg37EMAdgb/Kv77H2R7CyRaJdeXFz+5DLAvcvqY7q7IXYO
ACsgFS0aJ/j0zdVx7WUSa/sndDQ0DaQwmISiP1mAQlZDZQAYjMzr0zrUA/+HZbjHFVDt6PSZ2chf
QGNRK9/IL9jhIZFawvrt7KYAzORybpWXp/AY2pIduNWDBqwQrQbtF9++dCBZtzjpz9tqcm+Q2S4r
GACkMDtGe1/DeBYJQS7JMqbXInWOKweUkN4dzTB+zuzfNuFcXwk0GyuEVYVSEtpm3U+bqTzcVzLm
0ECcRYQ8pTYpmlPLCaM9XO0BMdSJjP9kgtJVUTgo89NWTj4qNLAkAdhSR2OFohJsemkQS9SCIs9I
O9IQqxPWdm1qX5WKajnDOlCl7mnUoEUsCtOWa8UoEYlS68QomCpNRwCfvor+8qgnff+pVHrYMREd
oQICO0dq/8CQZhQWTY6wqcM0lB38F8FmeY6wkJPj0T8gOju0CIY8O8hukTf4+FI+r228dFedX2eg
JqGJOdrvSqicjFn48exedh4GSw4UjADWdNrPn9yADI3EmAyDDstdOurr+WDlIY2s7SufuNZsb4Nf
Av7NVv/cYedlYFd2wLS4odFvgIz7E4T7oEsh5Dqf5VnrRPUW5b3IHuIeck7OwYVgUTQIh5z2bLDE
5auFOphdgT8YY8AGT/KF85n1TenAPRpYIzOuRMOwBsyFtlmdme494ylkWKtYlgoaPFz+mED5yYaP
IUskb5kmbH9iC0mu4mIW5AU3vsdjZr35emATP+7UF5uytDs3DAiAyTiwiA8nzBt5teS2ytHqUzLN
/n8q1OoCmfFLaaMtBcQR+shYZUVg+UawKjksnc7egiDdH/mDnj4xFokyPotQB+xrdpslTpBnsvPf
3eGAKzdRv2CP/7IeEYj7UUe7SZNWAHuz1q2OVF/FOcOHTQGIu6q5VfjQyrXjgXiFp31DL9mQBgaE
rc4675mDCJiZTRKdiwvFwv8lywZwyIfWFbxnbmBoBjD9tRoVeePYeSg/b9Avi2QRIoNpD0D/2nBd
5dQZfJGPVmuEJdanrK/68d27LRNtil3K2kV+VNH4H1+2wAbS+jHaUPz7ug6y72lLccDPt0Azpn19
ziGAiTubMPTqqY8MJhyBJ4j1ZsOulskQQ2nIeb216a+rhFlNNd9azuFvgnnHxooir5ZewgmqaJL8
mEwp827DD/d9yvaXm5WE0kyU6Y1zSfSt4zW5H0HOtxTDOerA/hJAWgFpeuf+G0k0RlGcFuv5MEJx
ETlKnHRTHl8dPYZoyDCzrRqDHrs3bpGYjACH+WsCfeH2T65xYYz0BpZERfk1p2FODD9gct+EufBv
D3RAiRWIkMQlcXoEyI0lTLpaboBoqiRzmfBG2Saa2g2RUqns4Es++3EYYc8vCX4TCp6hFm8zMkwp
zSmbdUVhL3SSToMpIAF9wyqNHq+uXBJANkYtEc9bQbCSd+mS/0b/QEDPTAkdww4ysLlyTwyl+i3a
VOC8s0HqTv5o51CPgDWLQ5kkYSGCWxnXPFFr98bpHHOgRg1PwFEInoNmp6VnXPljo2k9l/K53vZB
SvLp79e4ovR19YXY/Q3UgsHPjNpmM7RXEWwzvWYuW0shVBc39hXIdzTHMKiPnUUZG+WhDOd9AjOM
g+Xn5yPDPDtK5kzrJy4PQCmyGOeGBVAu/EYcP/W14b3MDdA/8+Y8M1L+kZet7WfuMvVxEsE23TaD
0815nufI4U89N9Crb3t29G52aG6ERXogxKRXYQjr/VLILhHL7OB3ivuxbr2m/oMzKrtMVObFoP/w
kc9U7wGVZg6IdbMKMOqkkfHwPYZyD6aqRq/7YOzLYrjfwSsbtXC5Xs4vjpc8evWY7+LdAZkn3eyN
FQGOJ0/lL2PeYfhQq1knOxQCJXbqIBndJ6M24BVucXzXtHyD/i/dJkYyuZKg1/4Y0cP0dY34QHXS
0S8LtLFghhoM000ANg+XafDR3E789XKv04MQ4hlMm27o/iL+x8lWiCzEU/bP9+ias1OzHhZmz3nP
aTRdLJK+BIlnT93XuSjvQ65XV6LUeeGpUrMx9XDEOA4Mik5mEZUhMEG3hHUl4Ieh3+wIcFwoFqbY
/Wyr0X2rIJ+Rb6bGNscdBbY52+TNmLb78F8YBjcqg0X1Vci9Iak1uueRMH45cU8KtWeWrqFluuIU
ph06Bl9HuzWa4ygXxOr7UziuWxo75CFX5U3fdLgIuRcN3YQ4xolNWtafYrEKZxbEifoG8acYySx+
9sZHrlQP9BLigazTEPh8xFmEaxLA+g8YdztPpgdHTRceDbMIZL60MbpMJXNCX8rL7yTN6WSMCqp0
SGTdhy8dPQEauq7ixu9SinVQ3TEUQySt8JR8hCPjwNqjoPOi3CWZ5AhfkjLQrF51v1DuzBwUNhqQ
CeJkNZt3eW6y7mCFcFM3UgwJi6YkT2t9l1WHuGHsGNOnjdup2GydRmX7nnyaDrdtUupWjXve5IBn
1odelN/Llwa1ENYNfjBH0WNygd1vp/Haz0b1OlVNNZ3UE11ycW8iCC6LZ6grrFB3lv1DKGku9rh4
iMnTQxXH7PnbJpd24JxK0NFZeK1jUs+aB4s2m+vf988WqzRov7CLKX0t5CEBT0ir85pmS0/k2haG
HTmp6HcmdjBYSpkOSI1hgQPdV0LkbjmzCxeVu56wCJJCMp2irGj7CX93ZB8oletcZsEhhiEOvBT6
6YSorwliBjX/yQQVaO19kmi/3kSegDpE4vM86/AnzK3QoN9H+Yw5DivrG+q47If4oLMzliKB3R4l
5g51t+076cFj5uZSZAWGI/4obAjXc4oCk1RrCgS2xb+dGyDuZo3onFkgtdhj/t9fL7WILvIY4fjO
bXg2ucGkE0QtaYfqbRr+OpKY+rmp9xW2X7QJTQxCIeuz0hikORI2L1I5Fw750FykermWAQJFFxxf
P440p0p/j0BurRuv24m+LoONd9aiIRzf42jdF2n5ZES0mXNVfZ7NQIgLY1CFRHyReDUdm2PP+jvk
fUEjD5j7Os65tzYavWxW5fBFQiz01DFUUYVmDIBRNhKXy0XEqhZNJszKoNnBCBK+vrq/gFueoDWK
gKe0jzQaCTnmJZC7QSx5lVwxhz2sbfiwZppF1Wan66Dys5uQsIHANnQDz/sR4HWbXifuY1FY8QW3
BUyUgYC/ay6uCNm4sYBCGGGL7eeKXwwxmn/8d77AuCAcb3XtrTdZbBTKVaLz5Rd09j09UrsBj6XC
Rs+jbP+w7wgAliKp5+8qXuVoRuSWkA6p+T1i+jtiiimMOBJLzK2ucPeCLG8WHXNx3XvwCQEPZyL6
d98pAsvGJPSr2/Gu1PuLEF8rA4fGEY/LoE/Pdh7pLpzhPPgElAev5JYw4YmCl3yFwJ1keTshCTtF
rWipbWzwB9rYDkc1Uiw9nZ2N+lJRYu1YNAnkkWHjQJ3eaS5nhljDLInQ1rPoB5KNi6YUirXq5tCV
EiSZdHMVV562L6Q+1rFcrnyJa7N3PTOQZgP0at/akLe5HfYFFAfXfr7LAZ9uPI0ZX8vROExFIQDL
eHUG4HXjFIe3ZUt/q62SjD3AblB3zpqaUK/ajRa9WHzyjNKQGjhp2X6Jrbz5+IAdAXyIJlZ8kqm/
ar4cFYH37V3oMwkCON3fYKaIfBX+OcugnH0IUkvF9LJLlsksE1EG2/a8sSGOLOW52YLBvGpdoMTb
8lffFrUhr9UqLLgVyXyo3kb8LYhRCN3Nd9voP29LjWiS4Vq21D2kTQ9q6hGPJ+UyHGTUtlMgXX+r
hhdVu7S/e2bUR81wqCt+iu2IAD2M6BDiorfN38TcF0QKfOl1muowzOFEJ/UKLa0pPg4OkzRjFO7l
P2VN+DNtWBwpGruVBV1oSwL5vrXdJU03mhN2Zz3j0XSkWngnMH3SuP5JMv7nnhSC5aWCqQzMxzPA
cGbNmsHXGi7jdpcC5trUUGowq7MeTu01dngY65NFWY8qxXE/kGlCCkO88rf8bHeTzmKyFvaRmIRd
OsPhdhygWVuE5eaU4JdjVjeSp6r31uZ/AQ2YB5MlxEr+2aGj+cO1iITB9t+84wgY/TQAFEPLVAZk
au/jUcnuv9z+Dp+/pTCz/xydOAad7wOWX7Gbvk9xgCKzTyTUvQ18ZEOSDW2HsFNUF6dYuM9tDQ8h
k/0yC8zkTpVx/Jx6DszzJri9mndwkYQSLYauOJS5pssenPTyWNBt2yKm+BCfiGAq2Nvpfi5cxPwm
2O2OBt2pd9KKJh2VZkl0EtHE1Kvs+HpOLDLyIm6EP01oDYKmf3lZ2hl+FXsEClnfCHpU170TEmuS
PVWu6IDqzLJpFo2Msd0HyWUFHAXCIuQMvxuZJ/hHLblpJ/vOX6VpLfo3TzN4Qj38dK+ZtGyxNJxN
c1WiEAT9RqmWukExL187qCij1OM1X8NEaDGNNmm6J0prSy0Ml24wSD8NYOciAjzhdGdwIgVcrcaj
sA9/KD6Z4gjoxQyB03lYcMMP9PZhHO5sodpC//AdJPh9Mw3dDPyoxQ5+lZm7GfRMtJe8z8mmRvW2
Lrg6R9uoFL1nvFUcF2JxyjnOC+NprWI5g1kePU2JGpRH7htBkets9rFXu1dqUHzysPD8c94HDSur
1epUj+jYhjSIDE2XopIoff6OvMzd5zIjfSSSlR3hnSYImjpKEIbl8xze/VPNKPzyc8OWZpjCSoOy
wYvQRyI2ztH9smoaSdEymWSogdLnw9QH4PcObZ0aBmGYVIRZ4C892+0W3RGSfkfjzdeZi5j9sfDW
jrljm2hcleuZ3nHDAOIxdeJeTp00sMGafx0uXdzUeAD/c66xIaCC+JnM+QIjWB6IJ9tZTFgxWLsz
847k2ZSc0JtOhSaNKfzelNIjX01YN19uWL3cU/2leMOoP5U1b5Gk4K7Wtdb8sC8l3Z/Y5QSHGZKD
TjmVIJKqe7bd8z/ZygulfqyKY2wCvILDhKYRC+aeHIE8y7pMJg01B2nRkNZUKYSeKA1U7tmsnAja
LVSeGvrkmnN/NHbx90eLFTJBgNItO6cy7aqinBT9tGx9Dy9iD3Da55oEGY4TlpEHYQoG9U1iQWez
GdQ8PPi3XsBuUPlQ57ZIE1cpBBE4ACrQNGQlpUtc6FfziLdmGbZaKYjFNANwcte9egG1jDWp6l+m
GM0KPTX2IK9JPOpic7VO0FOE8CWffEZT1eT7FH+9/X0A8rNyFm8R45LrXfrngn64XAqZGRJbYPs3
7SFQsq6tkj7uRsvvjpfk0NLtgP1oKP0RMoEBsTnDolY7EIz7DGGk6sQyJ/u1HsPpR6rxi5eg1o4f
KdZKwMYLmtkOBw8pfEbDZK0RM2g9x4l06FStq+jDHdYPbZDtm3fotf9UFTqiLzOZVuO/RF6QTZdR
HNmNvPq4izlYnZZIjDeYGtQnYIMbItIuGJsAdbfzBluFQO7Mp4CtngBFZ8AlaDn4lNjQNHS5LrDx
AgjkhoJV5AEsutADx+9NdjW4GGKMp0hMyRY64zd8PWAJ3MF8LNZnnOiJ14np60iECl8/oo8DEhvJ
xSkNat+uqmlIRSobXdJlSIACMcbtMWXynbfgeUmrIZy5YOjBYZJEdfORCMXi0nbgxfPnwzcnq2G4
mP7rqLTs6eIzViGJlUwV65bevntCvJj+lV2AxXdCtSZeuWJncQVcnQX6nZYN3EwEw4np5jn6+Cq8
sQgNiS9AhyAqSnliNIzmyV9fih99b5P2Bl1xMbNcChwSIATlsDUlxfj3ZqQhJWy7gZQUfWH09ocN
cPbHwCuoXYLgexrc6NQfEH8EPRzmXmHxceVyXGDkTFEqvq9/k3lDgng3hhGBzle3xomQJsvbjb+N
Xz3rzs/dBwaPOPjZTJU1qHUlBltZatLAPnOVKtRh9IIPdYlXcmE1SDvPCQq9s6sEIDvab9U9aY+Y
RShdqpn5riG4V8GK3vPo7aaP5aiBDKP36hD+3TIQ+ympRut0sDh/f0H9MIssMknIix/bGEPqOCLz
4sxaWtVLeViV1PGGp9tIjWuhsCNGnzkVQbIMUR48I5UKij4IBEvGNiExzRH0dBJbMxkzMR4+mHsh
hd1rEebWAMCJmJJRvfVfXy4u7V9tuvw5ELIjuoehKrp8guS4SV/7uEpaiB0aBrk1+JA6whGOD/Rk
C350LXyYt4WCNslsL1BTgINkN4QbqPMQahb3RfYGQmnLv2NjHUdDQbe5/6xmNzuw+tx1982XYNoX
o1TGWzZ/q8C/FywkFx15roq0OFZyVQ+CMI/iTN93Hh8S8ARiBG6T6EzBhQReslxeFMY9hZYwXuiq
tnifXg5+iLkRnxZvvG7V1dfnLXmn4+P6DfRdMuCBirVpJBZq7zQ9KUdq0hB5kqiSExbyHUPyRuBk
847uqUmT/VwUrvQgUb4qWn01yLPepkVTwgrra4xj0r5TW625rLBXXQah0LmbZJhahIR0wJCcLbg/
7qiffXlH4xA5PnbYlCip/g3qPR/DG8msHgjVTqpxFT4IZ87rhKEw/bN77wS3k0FpV/eGl39mekHv
PPkwljIbxosIO/AAopbyS8wJqNFdh7dW7KmT88AeRIm8bEZIArpu8v+8NlrFmRc1pBTLupdlyw21
AHlyblWoHbGbd3ejmOJklxakyPFd20DeV7tOXr2cKGz3d41mrVEF8luy5yySs5u4VSeAn32HyGz9
C7fRpxZdOp4nPXyzxEwY/06PODH9G8T8PQubWupn+9PF8qDnLOBLdxYbH8tCieJoALN/ZSBlrBOD
hwaLtUeZ/n9+iN2I+80TPc1fgKwHdocixcZ+myzG4A3G+9ha+B101mLxHxhCe7zcMakvRrL4tLG2
csn+Dvjt06tG7TzbJuMfutPDiOF9jUIDIzixEZPKOub1ERbfzCjENdUeTG4f1ZTLMXT6iSnTYGcP
M1MNgD2OC3NG8g4MdYDUMHGBW20uqZkSS2xMX8at1M+hLYBFZMSVNKeOM+ipEJKORyv8A2zzJhqu
3EqWQeT3cwS+MSogtboJonk4+hsNzNIGMbNmaKr/VJFCyJdUi0HIoO9GPPUl/y5TZthfyB7JP9zp
yT3OaNYnKt/7vMTrVw4KwnUEX1L4FX9NcHt2tL2oCUkreo+03eHietKexv1k4b5stxVHQlvf2wqs
7fdwWzypyg/OJJ8pVY3wCjPaULUvoJvvpVxarQidD29CsVmvmT8hCQMNVcrFS6yGh7OBDmD3LcaH
7euqw8rhrjJGOVAZeBk0dQ3XcgJQItLDOAbXqDRghObBH4WTi0re+q8xWn9RSsg5PTXjBEX5gCoE
61mFM/Dpzp9a14W8txEgRZswOabxUdL5wJhq86npbFozZJDKzyighJMLATFv3atmiRB9pwGDWVmI
11q94KGXB5urSnevcIo7yKxKIm8pTknIohq0gKJIxYfRzW6Ivsfta2NUhN6LkSBQ5O4OelmBwu5+
AO0euDDrPyqH/Om2d6WpB6GWQAawjNe+eY3LCy3K7mVb9YoakQPdkwalCE3hIFeCx7ptkw/s8w/b
P6TJaZzI5kvoP20dOrBGmdVLs9YwW+BGaTTgWSZy3EDv84vlmSV1qCDpJXw8/JFOYCaIZxdOYMUT
I6T4sjTJUj0tDCbQIml97o9OxjP/Mv3wjQyKOChQStHZYl4cEMmcf/P0jyRVJcdr2PqMt9EpoxNL
pqKBJeXeUSicEeR2EE9mT4lcxvGOZbZi9TfVl5W4BbPivSILpA8Zvov1NqDl+CnImC0F6RmsoBgQ
D8BgDhE0YhqIXyIvZCeWsasm42z4oDEoBEGIYLjGtHPO4bUf7NKQ2sDJR1Ts+qTrvXcqkResC8qs
8GMrKOA2+VrhxWruSPx+DVGV7FAhOnpRLmvFsFbRRNchU1YBGYxin2ynyYw6IfIK9YmDLGxlid90
YXwLoCEu0EAp+iJOYMzI9ttr6cZDyMamLukttY4sJz7Vw4RFZDnYvG8ZUuh7k4WicVTKNdo7A0F0
qSzN/pOQVn4ONZI/F5FGt51NEte2BdIV/YR5cYxkqPVRMnbg4iVF+oX678ZiFqZBPeurVF2J7xrR
UlCMykg/HFaR6IKAzY2HiXHKHLxEzU2a/ZAwpuZlONpPz97BPnQnTKe7MViQ8s/Jo1KoTKKmveok
LX9wTdBt8PSNLfXbdMVhYxPzLJneBhPTL2fqiV9OjQ8txc3U32NgGpZNkbxjEA4uZ1FKfD6J1ZzL
6KdrSVTjXCfzWlqt5mSsDg2BjanezFatMZhd3ry46eWzYgdG8VIlg1PGt+h3mtetGQ7UbCHMDPQc
SpnDqYaxOLjWfB9N4mcMgzIwywvjVhc6kps10MC1JHH8CYGry0VGoFT9tZWRESbyRHy/ZnfqnO2j
qiUzEFZk1SsFHGKBc5VhAexRYBXVRDFhBgmDHlxelNK82jDpn4S/lkvf1ESsojGMco/I1PMA4bLV
i1Saqnubq9kY9LJP7PiFy5E4/cakfcrd44WXjvulw5SoFDznrFL639rG14n5BaikfJruoJwIA4pv
l8dLxYlkq8WR64jkYiZlfrgli1nbcekA0/KxX3D6ldoIuoQsMyVEGwZrPxvMzpxF7EMm/xNW2OA0
rnqXTucyGz5SEhYe4T5JwC6YF2N6t6GF83IpzqmzZU5SHODRv8LWKo8ZmdShWpfeFGQ3GGVdsvFX
FPbCOfIyNSb5ba6hrDsH3QxLhS7ibUHQpCJfchm0Pg3phoa22oGjQQZFydl9M53Zqj1QXFcOc1EJ
TSeBV9Y+4vvWd9SrXSVByaRKVZenbEMzLobYdiL97qpRObgFSxyHLbcsUI3yXFp1wrdKwI7xQDFb
nQCplwBLDRGpqyWm5LWpkuWwDqIOHly7MjQso1ifyp+dUuBm41xzxStMJf72pTEMMaBxgyBNJ/FA
TdSVb7d+lYniU4GEsnRUCxdBtMzXDFAEKAy6SNt+zhl/eq/MuJdSd+HSgKEoB3UIasLQDZuZrlXI
5BPTnwk6Bcl+Axuo6zINXLACdW1Amo3xtaXwRbe0eKYof5YAhph0a3y9hb5dnzfGlgfusxR8+c5L
gXj5OjAyoF4rx8YcvYiZPj+l3cZm3+XqdvGwvRzWF5w5GSMt/M4Hm1XeMYMyMGCZmKUTGt50Es5O
OJr/sfKlztl01VBxT/RlTDfXP4XQwH2GDjQ6kYCcml5CsVJ9ttw0VR5/Er2hkoabP6U3BvRB/nMU
gGAW2eFQtFyqBs7TYM2d/GpCo2gj1xxYwB4BFfm7nsQLLJsIYWYdkHY9SOqa4CReNHepDKNhGO88
8pxFn3uyFO8tfuXDkWjn22QhatgQz5bdph1tzH/JG73Xmm2XqnXNprIvMdc5CYFmzfv0wDPej9bm
xbpZV7oPEeF3CppZecO4svKvDBzOuW104rZj6AYnkof/1MxHvJNBksnIeC2wz0GCbyXINqE40R0p
ewJucyvtn2/p8lHU7ma0akbLJIcO/BYBsGYgABwolEVhqo84SH4eFWhbQop3+PPKIJHCtmeDTBUq
l3XvZlhM3IJhAQmxS37cSLbaOQQcCExmM9AZLOp5QPoqWH3uvSE8E0L2zPlXV4YijGI76gn+7G5t
fetr1yINK+ErYgK+IedkGdkcgtaOD2qhkTr+K8kfapABuBTlLrVx/I5MeKUGlOLB1rMpw7pUfECe
RhyaZmp2W42s2Z6KVNP5SSCSYU4fIPQ1pG8wa/K3JQksFAk0J9K7BWjFfSWHz5wQzcHr+eUDlmNF
U5TTlTo4V8w4jbW/hOmbPyW0LaqZdWsrD6F4BWBO1len23W/8tOYMPSCNzVBMZTOBxIQXFx64GB7
JkLiMrlqSEeAsVG7RtkrAtwErnvyfZSHYHmWOciKAXR5bynrX2twRa8B9xBotlj6Ibw1Rq1ODJLP
1cqwXGgy/YliCz5mqfRHiUFhnKnv+YFdYdy8tqYYUWxWge+Oj8ODTXqTcc6WZmCd5ELtZliLf2ca
ROZyi2EWDnOaauFOxspbfr8ZGtOVjx3ft3MK2gXKpR5W0VIJTxkZa8l2CmqX1vePPVmcm7xJ2RHa
CTHhv4vuOvlwltDPsdmSILfbOGMZxikcykteqdUSqdWJhmdsiI+rN7BKljQ7ZbIEvATBRORLVZBH
4MB6cSca5pNF1VRHMszdglyBcOLGU7cBpe2qLfAiBOJTgMlO/FUQkKGLodeW1HrXroexEUdsxCYD
SLLnMZM2vIaObHdHOdQ1lxhLGtzKzZMEfIUSBERXd57pnpAyXcfYzqnPs/vELTBi75+c1M2cGbbA
eiWVa5ug3/x3dfo0+9e+blR7wYcBeiPRub+z/ZP8p76d9QrV4Igcf++7IgkKjD1rkamU9HqrEoHR
wTXV7AY8JB9Wo/IT6o2SInZDw6fZ+DHeAgOqj0FEdgwxh3rUyLUjcbSacYKrYuZkOEa+903yRTYT
C7IWblR8cRxv3W39p15wSA8gk06ZhdMjb1B9oVXB03MU1okQsXwWPYa2iMPdJRc8bsCBLqpxpwU8
ZmT+KLTlu2g+xUXWuClNsNJrwnAUog9P3czakg2GvvDL9h5NX3dymam435Hjurx6V1Y1yRaQLvGc
nJr5A0ctGWhEOlJ0tEXE9iAUPt+qGIvV4FoHb/fBfQQ4V7oVyZmQTyRdfup74Qsc1We/bhJVKyQ5
WsMpUrhXHxgqK3oKbK0R2HrYWVlCXVK4RS2JeuRx8aM247mwgaFQ0xtLnfaZvLMQp9fl9RE39tkR
083YBqEpQ2KrBasZx41JmphSbApmPn3VRJoCfMWHwokLgN7k+e8x1tmmSmzfzDL2RSTM6mVdej3H
0EUfEkd/JNhT6KixRMu3k0doDXiF2V0evry6227OAep098ISGHo0SUqLK3BxbHCXiyo4bwrhOlvl
hy2ksZLiw8loucy24v+j8yjlzA5CaPPOLOcB5PkS8sbiIsVnBAiXgCFJCU4bWdd1yimTiRjJmdeQ
H9pvzJnnbgLiCPolFP1xoeGUJH4n6UV/JHWz87VHj+JozIyPGYPS5luksV7DooJWuzhU8uU8OSMf
rQCwkc7ByyIXZwf2WsRC9SrKBUVrgivtT4D2Enq2NqPrshvAZ+7BWPmGqmP7rMPcDMA8r/w6D8z6
s8mM0GLBaLSeUNE0sW/Ygis7UKa4b0SalqbLIV2122dy197gI92pdVZYhtHdPrlyP/lDNoAr4YzE
cuSY4ORWkbwJtwnDVipLA60jSDFg8Run5bEL1LPOr+FA5s4si7urW8CO/JAwVXOh9kUS9XSVTKKw
F2WE/D2IdfnFfoyQmv0JCH5ymVK7+eXGagbjo6QluyMtwOPhsfwqBswlKEBR7h04l5t+6KxybZ1i
dl473aT/uY44NOdzmdMaAwKpce6O+9KSV4TXCEH1/xnMT2xguhcJip/xJqHKoeHSvFRm6yyHlkRH
EHVcMF96CgC0Q2ii98vf22Ml3qFE/zwc0OXnGA+XvCJBQzTTsM5SM0G/P7aGT/NEIU6LK2GxzOIa
4uj3VZqBlW4hAN06Xnsbqb18RXY6PoCI2wBBvcz+QNXFmKj7TfUeJHWLxP3Oo1RqNlmRapr6QWHh
PiGF1ykhkvkzzlgAFpVKKTQI45pVCy2VOr/ZmaUu8MPLGjXuqzWGM4IaObZbHjnzAvpWbNK2SalW
H4HKWM+/wRb8tua3Y/ffYjkxRAezx5fM2NtQIxx60cZyUQhLxJ91vAGiO13WaGKTQaLL5keEG15J
zn6NJvwpYqhIMmAL+eTWbRxH91fSL82hyg7gCZTkHiwk3Fzn/vsCy/xjrgoeWoZh+KWy07LAxi7o
fJM2F8PCed/3qXwSmroWcLE4cl42kHeO1GVcWy1DBb/Ib7KKNfDC6QfYJruSsVMv+uCnWogrF52O
edfU7it1M+2aney3EPBXfWvn9vDMyWYiZZ5c9N1hh3AKG6ftnp6frSJ/sVgm5yl10zc7XTwfElwb
+0QUUVQSdD+1/44juzdFawTIrU8OmjiVXIm43+hkF6TV5kf91THIiAcrykgkrRcPhtdqQUYVKx7r
p+FtFtEQOdgPkiG97JaJm831OK/XYIrGW5CxPWlis2nZbQeQFIlg9kB4U2Gd9Gx8Jwu/X0BKGIwI
yuE0s0qZXh7vDUj5LFWcet+72yyF4OqL8fO47pR4nQSWClh+QZXnoP1+zkwjhKF0qHUvnJe4KQ9U
E+GatmUAzQsDLpx38r2+16HtEELTpJqxLXtkAG08mEbLVXdni34pVZtq1rGtE53ikI0QTclbn6SL
sXbvKuPdcnts4/tyxVx0wsCBX3xN6Gde61itavVSfYf4RUABP3wdfLHM6oM8Us7h8KgEYJyGjWxc
XjyILXErLJEz7DsXDRGTAU8EauOM6cr2UJPLr2+XrTXcmVmq5lRF4CraaGT23jRSRbNt9H0qhulr
6WxX87mwomCoizfSbNRYLVb9hWzBjN5+VBV22wp7XIRzT8/lNR7/93Oc6ou1IP39ZFeeDO9wS+oq
n+1AS9QhxJMTmImzHL8HZE097YLBP55AlaEDKcslHUUlVS/aPKpoK5gyqIJoijCNE92k0zdCAmLd
ZyalRB04qVGbi4IZ121eHbuyBTZfFhUC0jLX97kIpPAM2sZrBfMG5e2VId336/Nh0pFLltvrvHwd
m2+Hx10/BzXuUhrWicgrET5g3VsSzK0wuD6Izv3c25AUQlV77HpSuxwFC9SPpO8S6fGzOpfnn2Ar
+kduyP8PFHYe98NXPHlizR4YfGCm7jcEi2eWd5N6/VlzJnps3yPSq7WLkBgNWSlx0g9opDSd4U1V
hQwr6/X0LCZBOM01XlVCrYeEpTZVkRf9ZhZ4y3o0/dksfxbj1yvHe5eAkGtzub5t/w+mN865UTw1
cHacjJcxiJfAZjc5zgwUfk5WJC7+YzGFAf/bCTmEwKMUxQL39tuFMdNoXvb8WeO5JxaS2x5ueYri
2rLagNAxyfFB2I0gGeAqeaK/fEw+UCa30WQiWkKY9k2qT7bS9BJJemM8Pb8YPsXSPUlQM0FlKRp/
/kSZxDsUicXrWzUGZ+RfVC6+hHeyUsuGR3xarLSI2rZ9Q0trqOnrrStONJz9vk5SsOSdqz69a87g
XVif2V0DQr67o5j39b8XzV3XfpEO0KwjlSJhJCrkTm80fO1nzvFhrLQnZWZ1lZfAOC6Px7GKDES7
XCSkFnwI6f2XOMO9kW6cIEymJTOF5ScjMWbDRMxALVNamrFkqy2TNhVMns8NBEhlFJ4iYTGOsZ3k
LEPBYELWziL4mzJnOFTwCN7Nn0oUuX3KvcA61TXK+99XJSGMMGcY4qI8DV1gi9XVRtdQqEVhrmC/
vjZihyjUfF+B3k6DEL8rJSXUbnT9fjzM+utBc0ENsRtFNhtP4mpFfp8ZNhrWaNizjOiku1VMpbq3
1bQCv+PoAZNf2+hGqAv8uq6g6o6QvTPY2/S2cdPvfU85vtBWAknA5E/qY3MofAcST7M52pXE15KV
5viJmSVUJC0naO9MNe4uVZ9FB+lDx85Kv3CYBDSm4T+jfvTN0pQliXVJ3xSO1EwOop5RP+qe2S6g
ssjpVXrWL8puzYCx6DHPT/OjOikjfd5QQdtWQnakc4jlghS2j9nfGvpN8pUCDbTuANE3wulAuPf+
24bc5CIjI7+7rztemU6wbW/URbjphAHPp2+Bj7ifNJVmz4LjfRkfWJ7hdyf2fT01TVKuDYdfXtpG
Y+99m5MdPi2HMvHJyY6AvzCF0YjDHX7Wg9ZeijnxflzoKKRxolBtLo8TaHGjBWcCi8jZWI3dKJA0
SWNZUd9c/kwi38rKRlBTHgi3Th80Lj5T49HWfLMMeTuuRRfYajAnTwz+7R6vNeZSJkG9eAqcra4a
Mxy0cr9uq/8MntSMIHHatt5kvjwOzJkT85l5iO+EC60tHh7FGODCa8VQaZowVEoBhfSIes/mhhSl
OSaz2Frxh4zRvolSonvszJYvAhzImyp765OrVX2zC5Db9u44zbYx5xPe+gLWHa85KPDYyy6EoGij
WgNH4bgM4H/vm5x74vl74hnI4VK4be1bHMEmbS/mNbQD917gDQyoazpNZJbmjqK1/kXLCIeeLmrT
yHP3xQRLy/VJ5MAfXF/XQGGYozdI6cCIHpl1chzlXYX/JixlKMZGPTxe6qD9Hc+vuL7+M/LaiEc9
h4YeFs8ijYycGduPYwCVZ2hFpSgxTDtirlvGmaB/MnVJstGNNBdnhQLhMqy881nbLhdIM+j4jv9w
MHoZrz9MkUejiTxSdIMVi6/4jXZTKA2wbMPVEXeqgXCx/00VscZMCKzKYq/kok6glfZ/r24rr2hL
+N18BJSRRzRIsEGUnFqp6+jSqSmY0v8tfUqYhPuwB94rxkCwLYVM1JTBFmQ0cZnhDDB/MoROCCJW
Ub35Aq3YcE47jcx9Fj3LcLxDSc7ca/Ynezpo2mAHpaXrT+GEyn0ev+9iLWQ3ijNaidSmML5iVLMO
12JXeRIIOHQ5xl+6Ym02GDX+U/I8mxLrsSIyYCIUcxvD2zJyvpC6cXMqfOf8caMv8cNVsxuCpi9e
jfUPQmB1tfjOGSe7Qa+qlKHYPxHRRHCUuOBkmh2YFKjqeE7ncCJYnCTLomS43ahHrJlnr3AXZ2AG
nn6F1bX4/y/pIUkBBQ+JRWXEJfSkPwxo9Y+5AwpjohbccvdgOSYsOCaGK/85ksMydwCGOzRvbJdx
njjTC8ZXlZt1MecJyhuxDwyUbDjT4aoGy71eo0OeIOo8Kj+JPUO0bE3GHzG/FOBlmiAIOxfK6waA
LByr8RO06ZSfFvJIuXDNeAIitwZ08X8wo6Niyuz+u6NqQhfKN70JbFG+3/YbSoAePFwimOpRPor5
E8+rJIWl61bkDbKDOKMEVWXD/2qa6H0b7zrU5Hv3vuAlegkidpB3AdQdg7N5IpGtndVwmEnVA02v
rR1ztFvQiF1myVaNpyyfCSlCWA84uoCr+AtjUpJtIq0bb3Ye49JstY6kd5G55uxSXSEFUk5eD37q
jy3ArgiiccgD2Wk46KHg4udSDrHVuiA5HB7+O+qVTFgmeJLXiiB1ogpSzU/fHoZQUjkt0g+XKM9R
tBf58oGDi63/EryIVgXJHm3Jgykej5LTCVnlNlR0vBmxi6c8D9eJ3KC2rCiCkk/YUizCpazqRHUZ
4acjGhXIpjYlngspAs4I/vE+sx/HRmb6v+6loYMb3AQTt1CPslg1Gj28YNWBbvjd5JaBYkNK38cl
DYWcJhyum2RQFmpRXuk0muA4vYyx5rkfkMrkiZ3wnpOnEB0Z5ZXAXQQ8V50G/hNj+vKR0flTK8Q9
QATli2RWgGOA7S1gdk3yS4TlJox0NaXmZiljdBD0/gXgvW7yLMW/Ej/4HIbS9K2yvVEHppfRdr0R
Ck+mjav1QYnDdauFD0BNDwUT3OPEiW++V6EITL7WYwUXUpWLNLwR5apVtwkeLRwCs5wHwEyGjKIj
hRDJT+wmNevosQw4G+ipgWZ49CSCvdJo3Cli641ehVLZl1UJSMFs9pbsKcwJ9ePPMEhYnS4WiCm5
KesFfZxnWgIr0RBPpex8Oh47Rz4254dJO2gFwONzS5dmA+h+RLir/ZCoTf7HL8O9I+x3nWLOCVOa
YWC6Kz2KYXfCsfhKgbCkUje+M+EDM2ofdymG0nFbHXwtGzvQ8LrjQr0Dx/NXumknm3wNhno2Crq+
e1MCKFzKaArdrLQVkhyPYA06HVixszjEOzJm1rBkgrlTCzuXRFFzM4f5Gf/rUNF1NgVOnOekb5oa
dWkkLiHLX+1jT1BFiKJAS2vOu3ULeBQS3FxPKCcYS2K66Jg1+yOGgFCTEqQ0srofIdyfyWJn9K+t
nKVEI6zQfz/Rg7FMJWxZuQ9GKdF0aBosacrQ2SFxo6qyETcfwWvi+pXlGf/M56ZlRAShkyH1bN1F
En/g1OW3td+x8NbGiYGFR3meB/D+K/9f2wyoctvOCZZmpvksxY8hGywweFusAhzkiAFSZW1eyg7m
yXqXJusCH2mI5B+Lmdz9/bxiRHwRMpwhcx+3GMU8q5TxLhctV/QOEA2PV0dU6FxvfOtxbJRpLzI9
zlIrewVVSMRi5s+mK6oFmYs9q7CjY8ZqGrSNXWrsFN38CHTw3R0eqNi0I2Gw65qU4Hwc8gBMDVF8
BBBhOigmSxwpxW8jT1H9G4owPjk/l/9NmanwVoIStrOATbMn8vz7VrHsPTRKrmKIDwLNpDG+FxJk
pNVIAYYUrblw5fiQAuX5RsOLyVaptDqC286gPY4BBNl2k/EF/AydmOaxZ/5tpKLgjKoqSFW1s/O5
RLShuR+0535LzqDLnQLfQcIR7F5eLqYYaxuRnkRJg2r7b1A5Xxf7LngIZgM0DCZabF628CGEwWtP
BeeneKmkpD4PUcedqEXK8Jk2rtXWXm8X6J5oVnOZJUgkUNXksE50sLWO3RGDlESjQFkLQ372Bp0k
SODRM7KB25wBOWmHL6bZtMqWmD4nf1XD6T/cD+TaZ0vcTv8YxpdjZ68XYq1lEAQktmcPmZq/qsJO
kGAwkmOFIf+KAWSnMfha9entiE0GWilC9AVWtkBHtoie8LIItivf4kadrY9wJ336qgV4DH2Si+Im
Hky/BWG/iZ8JPFyTSFqwMAwElJSQ9kULzTnSm97aoQjAIaDqIspRxKOQSGWHOa1IB0GhayAAc+eQ
C+rIZspskaCjF+LBccjrCA7+wg5/h7wX6dqJ9iQ7fYLGcZNrHfDaJeC3uJJU/fNlZs2o0RQBXNwX
BorQY7UC/qzPNBr6VZ+DH5GyfMZlbWU/DqqJLAy+4GTkaaWLWQoUsDb1fk9HFi0CbEU/DvX9/ntR
ucRvrsDpImg45x+gJzShHXejT7erNM4G0S4BWnGpedrI7URYsNp53KXx3lt0YyG6hfoCaJ0rk5Od
N8CAXh+5BiMsn3qMsqt0eS6/VH2TklFa94/nfokhWW7VYFafL9knqENpt28O5IvZpS6n+jpHMYgZ
zWXJCzh1wRV7VLt5Hhn76yYfohHPJzUUEQUOlD8BaLfiCAgGq/R9nhplDmfSUTQn8oflPRjUNx2j
ITivaEgYVnKqE/I0pPYCrb54+doG+0lIRfq4qputbHhdBkkXUMQ8PDzm8fOfvqHi5o4/zd0sd80y
MPzOc2LziFw72JGJbdVnKzo7M6INOlgTyyaJfq85aX3TJ0iE4wkAbqKMPDk87U1T+GHNY/wDB+Nd
ppUlCfG/WKKGYrQzIbuzFvOsQTsKu0UX8fzykRNcARGiPI+JnJhmRLIbHq0yeYfcG1h6oKFf4eFl
AR7dNRF5sEpF0d5BVIi5Pysa5iZzguwfxmU3JJt43hbnUNcTl1A7XU6IHN7JW7wLfxmd2C/0tADA
4gmKhK773Wh8F65xL/7us0xjG7pGYss2TsIA7TTgwyEzx8SO8QLjLo3tgqcj4w5SG05LSosmuMPH
KsKZ9Z/eNX92yJ2y0eFhWoYBUe93XsN4RBJ61jDHnNS3a3BO9hopwbzKsHRTjPhGOSqJdZiduhK5
/YNtRYCcDmf/W6DRribpuRJZMQ7MVV4VQqfZAXo0d/niBIh1x9mI4uD7PGXwjMB2VX/AlwPNGwkv
tR/dSYr8TyQE34LtRgZfhLfcl5b5phxsGE2w9KrFarLi2Hp692TM4J/x6Gn6hzBdddZd/Ga1/BRG
KnXwTzsAGG8hw7+qUGhWsKHrWe6u70PQNqLeucqnDE7C1oflQblIibN71hDeGuXIWDjFYoLv7K6a
tfDEWONC9eL9nWqeLJzwWdDq5S+DX9NROptNmxZMm64tUf2zbQj85Oh8YRZ22+75tfGiFY2scBzG
00n7K45jIwA39FT40vKsD9tGyED/YM3qin1pw21vAYHMg3llaGHLAke+oX2+9ksr5/HUFLbwBMHN
CNtandIOEUHFzjUsSV53DTp6UDno09ZyctMMLFEZ/hkJZJ931BFx+C/5k/3dlKrxBV9R3wGjKRAw
htrwBUDSeNYfoCfL79+yNumSUYBLnczW6SyEDpoXNckkSCNFVWVEAGiv8AlN2cDSDPY1HU3yCvde
fg39u3AtdXvbG0ZWF1JU+pDUBXfWaASE1idTRI+NHQckgSe1DAc/Y79xHYS/XBsF1/8pCZiHtts5
h0/3EHnM5NwpkYHr/7FXrSD1xOfWcFUhCHiR5VAaq4MqM5T3Z/h7CosuUYlz5JCTwy+0ZsAbbX5P
8qeMDDk+YJhWj+MCjxpa5Y4MsbPgLFcVE9uSLODg9gFgRvmSeeCQwcje6pfjZatiMt1U0ypAd4vh
MbEj5l1QQV3ZRe6M+I0pk7xb/qYaWXdaXp7XQnpMMX6Sh1Bf2goQ9pXLTyDcB5nbT4EWG4+4cCH3
Tpws42j950pfyrPTYzd95FL6qqKwZBUAMU+24GqvodX2GwSN3BQBgtwssQpmN6AKNVaI6WzE4YVj
rVpninGKGRlcCaD+A+PhGpTjTRfxT1LHjPF9xgcCLXNJHfCBRZXVK/ab4ve6JYakRAC4rSCzqZmU
n9zpNF4kIcDQHvfnUTX+jT8TKYfEea+BYipTRy9UjV2T18ZjWaIGRfkv6NaxIRzx+X1nB9fWh/q7
HCdeqOexw/XdwrxyB5MoWCsWOsc5F/4IFl5oxyEC6lvC/apgnY9yatregLzbyauIdTSY1fmsqeTJ
lFnO4iYGAA07EAWty2CHbqXnWHmLZ1mS6PgPFQtPt1zekdC1aCrlkNahwwrco0JMEpFL9S2GnPez
9Ua1PNeuEPciU61kALh08g6bGLOhNLHLk/F5geHNVMjLEwQ+BudgANzBtFAFh5dYfbUWtUWxwucX
YQmXABYzEN7o3p8LygzoM4MF4BFjo/RpmkBodTC0YcYUyRBJI5q+uhzfl5ZfgwC88EGK3CtP5l2T
umPgtqmjiTl7zq/hthRE8WqD/Q65XQFvwrAUqqGGPb8AGTsEdt7nKTotzYXhOaT7dTx7jrpEQsob
tZhNzMIrceZHv7UZq95nh4XPmXRc9+kh7liqYoY/bwiW/S8RGQxNlpM19gRQW3JWRSF7K8FtRXqf
C44Z8cW3FWZ4Mt2FgmJwZz0AOuUQE8vO5j+yWMtXC4Effhz1U/3OgKOdYygu/nLny0wEWYmbPEbI
pNYlDuSM1+srzvxfN3Cf1sf+Dn2e6PwKxpUnlmrAoyC6wLXDhxVQoF2QCXuCTYb4SJ19Rr+hYtWJ
JXzTawcdTJ2vKrxF69ghUZXQnQGUaXEUVRxZJQij4QpYy9+nEu43OMBHIw4hMOLGcREWwmoIacPH
QfrancywhO5KAE+BRLS+OcDjczFdVHuwCy+TWzwzWGdVteIlK/3G+IQeUnLGsSKOAEk+2Zw/aU6K
4rNV6/8T1vAPOMZMfC65fDc7bA6FJmq8XtHOp2mJGmfR2aR028izi7TRnMNGYmIWTEaCAn83olHr
o5OraABHyJGDPe0aPXdt3WiOCBLOtlRBTqJaI6PAp8azfHEcjG6zcZAdAwDyqA7qkcdxk6HMcWIT
Pha7quH4GO9PPtW1AJ3HoctMrGrv6o/JgR3LJrIVbdqyGUUiHjMBaJ30hFlKey6YHI1RMDU/Bgy4
VQr+SzkU3k9MSwNflG6AzAx5dk+4GO5/XsymELnVcF/R3xNzBL+OxftRUAE3FHTRDDCbZfaxHWl1
bGIq8qppZS8SrVThwkENXTSncbmqPLGEV2LOw+tm6W+iTSzffxUeppbkgZ2mVMDQ4AKduBRP7+cV
YCc3c/qH4sbShyYVszv3VPeqy053slaFk6m+nS6Nu3cwtRCmpQfVLOJ7uI1tPriLSoESpLJ3KT3y
T+0TB+ZvLek0lOGRE10TtKKyKNmZ4u8HoGhLcgRDakYGFNV3gq2BYTN7IjYjVVURxT1atk7F1UqO
bdVKb/vu9KnTYsoCjZwzUzkvakp4Db1U8er2h6lje+/iLxFnpX7X4EyLWmOiQI4B2bRLKyv9Is54
fJRXqfQr+erPYltx5VZ/BOK4h6Lymbx3g0qgrviZrz+UV3sDnd/piyVSlXCUB1sWM6n6wDqtAU7X
5Hk8p/3FLY54LUayYWmQst90emZIfyMbbuc9tzokZHH9KoLUlMGYJb2nX3Nvy0hpaBJtSu65CTRy
0KlGmB7t3fa5iY85p5hgdrtcYz3Wl6gV2Qj4MmGZObnYWl/XM07KLch9PIp4X8QmGjGwnfvsXIgb
l6Ygdtfv6ln6OSpbWNFyPYDa70/PMdpiUYVPwEpsATTKFYJBIlysMfEXOG/DO3zy7RRUs114kH7a
l2WfuEpEiXhaoA17r2+PdxdPvRzk1xtnYZs1QAMbNx6nj9s4hCJTP9iR7wlbwcJVqQ9iy+9U4nfb
V8NrWDuAAb7jsLOgnqb4VXBhs4brLLhoQuYOgLUXFAqEBT89kKk8w5yMdfASxiR0VuwHOdMhVb/N
uVVbAl3Wx4260eakD68C+qP1w2lCRv6cSnWFZzw3HmaYz59flc4rHRlmdThXWXvb/gO4ms7uKnMc
F5FkWCN/S7PxiR2497y+TnvetF+9fijIgYlP+VtBayDiYP+Y0eYwmUlhL8Oaeja+kg/As7M6w5Zp
eEYWeGoVG72uU7SrWFgRs8jwKqd2Ommy8OlJZu+yEDrsfi3ZQ/UtawNUGB5G6TQPTnfZs4TY4WEP
jNXIEOppx9IEjWS5CeoYs4cEl2gvqjev8Ge3d+FxtbOPhToSxtOn/YdlFteyN/XR3cykAIzwMLRz
alORjBxk76lzfOdRuyjxsgaMmCH3BVg411owJTwoyHNhVj5KWCS3bhrOcKA7FIPPzcxOW5kOfS7b
tesxvHW9Z5W4TLheP5cCvF2Bm5yuE9sJDbD7kEuXw72aK13GxR6vhAcJtMMcBXWzjDpKS5gzoSm0
n7SnzaQZRZP97coQJRDbAtpkmcXz+Hh/MHhsDOL2utxVcvMGfn7So0W4NQNbld4yoX2gp941aTny
Ajl3LO64ldn3AtP/RpwpnSCGCzVvDceHOSeN8qagjaGYgHhPHQLKqJa1qTBAbf3mBs7q0OEpX1lA
v0p084blevGrz7poQOrDTAhuFhi1mejH5yCm39GJVMir20is1/Um/ClO3pB8HzPdYtlqJiQ9BCpG
aNuaGzAci4rOm/ZQ2XQEzdmgZVCwgtw3ney5hPqryApNijoXAUh008nnvxmxHvJ04bg27n6awzIi
3IMElL2Bp5Os7IXtGaBWNVQEoQJP8QdwLEed57vB9BnLE+kBDXVPPWx5XM1/F+bY61alXveeG1Gv
EDGHade79QsgCha+lAx1CQr3Pm7aH+CZ+7aw2MZEJMgZm/ldHoc5WhBtOt55sEFDezNnzprwOMNQ
WEC/PK1ZztbnScs5TnmKwsPZaoaDKd1IU0arKiJlC2XzoYLU2XQOwY4GKUOO9qO/PeFBxZHNMgsf
qFzu+u8pnVEcyjNffo9fi2gIA5Xn/8qw/c0sk9O4DbE51suN7EpdjLj4wBq+LNc+pk/lc6x4pys0
2+kGBClf1slNUw7Y3gS8c7QPeYcJu2pZHekL9pRt+DgeaTfVe3023soDZPxpaaaygXgFGVOrGCsg
yrhasmgDTH+jfJXmbwuedQdR5szZoC4EaAkhB8wG39B8idxW3MDN6iI96pWBviNJuAWF5w/uUCbl
p8fJiv87lQn/kUxRAdillfj1PSbg8YupRq/IuX/KKQTBWw91lu6OfXQssu/Mk+d3zWPmKF1Y5M2b
Y1+iHbKRlKSpbaiapx+AAWjoQ++sZ/aM/wOLoROMT9yALzALxe1UTcS/ZIIF2xL7lLkTD0bKcaqH
x+oEsIuVbXk23TCVGvjuX0gMJO9doi8nOB0ojqB9qYNIKXQuvif+ALyQCnT8pXJZY0whajB2BIYq
m+01Rugh8pShVgcsrCzKgRHHlrNqqFv9JDGFQqD9gW4A7Sn/zVZgifvDeWcddL2kEGnY6IuqOo2y
/1i8N8TnXa1zaxPSFMvdeb058Jl9CCJK4jwUfGVTcKhzvgcpPoDvqH/WVVsyjlctgz/0I/GIFc/8
ZOcZN/HOa7GONQZifJQmCvLmr4Y77RySNGdNvGHVOmcCVTaCc2H/vpMcWzUgT1d4+a1uCyKuXbEq
JlICU+RiD05FIPFOI4PK7wRIQVoaX9ADFC9CXZVxHnodFUIpNfmANnosCSFgE2afi5d7BKpqe95E
TotGKj1IydU1Zx+lTClTl8HmkXITVQg2Gx8lq3jRi1ICppQZ9qjWLBYCXH26un04XQ2U9aPJfe94
H4/IjoJXLKSioSFWR5IonrPuTpBy57d2guys5e+ynYiRWBAYYEjkxjI9Zkmtp0BH1cr/DKSxJ062
3ci6EBoJKaiOhaKyXJrQ2T3koj4x4w1ppV33dw/yCL0OZp+LGsuC3W0lSrIit6eWdVM7JHVIbeIb
FptIFldAdA75WHCNhaT3PRsYKng7AJweDfaQdwRumOK2Dda8aidQhCMz6vAj97mVT03Eo0reMNmn
xElYPYSstvdj39C7mf1u1mtFIjeTk8cpqTt65X+xF5SfxHtAfRpr3ifPdVH2KZv15Hcd4V3xXFEU
QC841eyjrED1lPU+1SP6B8L5zU7D7hEeR2cYc8k4MCxmZXtNWrkOk31bAHMA9eWTd2ysYkhyUq62
qQ5xZPi53w260M5YkO7PPpqnUkdakaPbOMGnBzbjj/NOXMRSo/TfSCK0pQsR7lcuSBJz+4UWtwBj
yT4XEEScM43XzQ64v7xcS9LdTMUGh9astk9SlslZAEliLRUYWzSkTp/CLANwBqcPos5Td/QPCWNS
r3wylsHXGgtXgcTGe1xDaqUgYyBWNIRgXIraXm/To/pe6/ZXd9fhJt1Pi5bWAU3YRMi/oNocWStU
ibDumu2WoFiu0EsHxALd1Nd0ADSNs9rW2VF3/Bh2VeyQ3LkdNWulrCdhod86pu36UEkVkAd7sH3r
Th1oZ4FFa0S321k8wOaPxN3YYHoUFKOcwIIWLzu7+4neJC1FiXEJXmva7IczgYw3GFP1ZOR/O4WB
YT6bInAco8rteX1gJvTqTWHzKB6bzYwBm31TfC1PHANO79RirTylKafg1qar6iRGHGnHre2SVLZ6
5D+azEcw/OI2tvVjm8PzbWysqGSpSZ1HWbus8TUC7h0//qZrFiAjhrk/hCV1I+tSapkizCfywjNI
e59KPFI+ctLNc3eLN6Jm0iyAs7yJzjqnQS0Pk8gM2e+GUgAC7X/dJp6aVWy25jt6S/aVhYCBj55m
PlAblcpxF8iJn+KjhvFuiUFLGNW0j+2V/S4DcBm5yNHJ1FJbXFnTz79XgKBPPBKIvFv96Yn3La4g
xeOebfbP0MspjtpWJt+VBRnd+sPOAIgEjdxQTmx1uX1aKPqmJ45BOblVU27GaPsSAVpcOZv7fdkl
cESRjLFrui7XbVAqfJbEIr/xoKrlHTPi4IZgZtDIbR+SCMRWV6rDTaKFhCeKF9+vZ5qcwNytQT2R
Um7w2owwG4h/cYoGzfi8gbA9/FflfFrtgB22CnImv4r+zANzsPjdrrc9saPEV6x2OHWEfbGkYteS
DHFyGRVbmP/8cChDnfP0X/QLS+JJoxWXstRbi1l2EfcV2rA5O7GwMVm2a+sTw1hY0+0wj2RsEBYE
LfGEUybLEsQBXyK8wfZKIbIsC9N5CN/taroHmHBQIHVNGdle37axwDneEXSMrfSa+tglOzcxbhX0
RqKReFFMtAzKdjlwlbTABYMvvnwarKFsVziYl/BfjKCZonLWMdc9yuWvEu2LcqczZjjMbFnB5RAr
ksbhNgzItyx/HXK3PTlGtTwwafrW8IMn4ZiIAtDAir6ECFfihRz5knlsICeSoOiRhAZVhbWawuXm
AVA7bIGP+ACC0XpAoVMqOAAi1LPkkYmHw/VEc5uHVl/WiDVH3QXqIr4ANpy1Q/TFJae4cQLs+w+C
2kkidyo/WJzmDJoiCuRf8y+sPIJMuMGZ5m3CQWcJgq57PcqfBCCb1j8KbxlUAERYrvPvsDViryjo
UxzMj8imkL89dhfXiyuCNLR01m8PzkD2Xny6mDXN3ciKwLOX1YWXAMEZoCn+T5OGyA1nb7PGAbEI
4/hXnB2giNP6nKfAEeRrg/YS+fTh1S17EAz2L/8oktGROKw4PiPBLai3bsH5DTds53LUi0e1Wvok
4QQWYlRw8TirwFKF5/tev0f540sHl4I5GvMJpKTS2bNk6urpGZDlqMC+IxQEBq/Tht7jNc8Lj8zJ
6lWmuyjHtYIBc0P+q8HdsOtKEOLoFi0aOY+Gdy2Tuvu/aipBwvifqa0aGoeV6ybuYhb/pWxLA9p7
ClNBrZp7MdBnZ+r2sNDQ/cJFdFlDyY74xrygiTnPBY1AoT2ih941kmPmQfJtrZD3VlhhF7N/+RKM
Sc7qVjFgHHC8H/mOnzzr8ELOY2cagw0yMHdbv6bV4r7VOQts+X/1gu7KJHCg4FAwkjqUPFhgyst9
2HA2jy3Lo4N8UNWIhysHCyMF8aIgP7skNJVlLBlCT4AlZXeE1Kqm7eawt+iAUhXRnJ1xltsMf+vF
XP9QnS6EyiEXvygcuyF1utAE+KL/30O6M49NmNRnjIYNmc1fzoX9pmnvNklIOJL4Auz2fqK85pS5
mZaAqxHvUfEjH65AMK4hNFmoxY45jUZK2wAHvOQPf8bc8NZ3dILk0X3DLoMSG6o5WQQ0SIN9Yt1Q
uqdNfP+3F5EhXkCRqSaMQbJDLzC5PN5zFidM23x/dfpC+ggeMHyV61tO3Uml1b3WsFSkDV8PL/cD
obpsY8TBX7ZQfOrQHwjgvk1lhWVWR0s84AXMHg5Qd+bn+H2GLda4G1zEKAFqCaqZ3PjzOjy/eEp/
rITlMQyxxh1+CQNU8UC06d8/kE2lbwv5y+xjKyZQxJ0RR09au9eTq80xhV4+x54DpB5Cltxt1cAL
w6hWJknK17CYC80pct9C9rvMWCm7VaM6i+QOKxAD1RFO17LyKix/sJpkODVd5LN5RHVDv9vlGbAL
Sxrz0EZKn3iNMW8lpQb/RTn4PBiiKVoWLvsfLPXbdeF0yg5dcB/pNXBz8ighTdhhkVG2QqNaWVsL
FZWNP4Btf7J7aKWO4v+EmYMknFugMpvQSvxqD7A8J9rE9+BX/j+0n8fn/YgEG4BM1QoI5AjQ0lse
atUVaAiFLdRC8JLo3my1pl7w2u/zGNEIpY9vG0+XRD2er/Sg4FpsB4YPMb7bl/jg0jU390Nli5vU
VrPf5cvp1coo48Bk4RUrqdaqsdsAr+ymQDJ/0VsO6AibBWsQQ6EUWayZ/6nJPFIbyWCSeUnzuIIc
rBQHoqcioe8BccndA0Dpsk+P00MjI1goTFwpcUVoaKBpMTACOTmnMXWle6HUaWEDcNv+gFTghof0
Uo+OPIgS9Pajj4al78TLbBJy9hNstxq0tCX9Tx4N+yHJnTzL9H+XMPfiAdu7zzylg5VInTPZ7tEq
uiaO7YhD2KluaxrFpk8T1poCs+dQxfe4L3eOzwyNq1sq/9hDfa5YmNnd1LF6FUxeWySe4Xn9h8Sh
9EJGiC3v+AfMHTR7lpBsxljL+7LyZ/Bl/oBiEp29fJo1rRcCZDe/sv9nAfpukX87XGfVWD8dwhsH
96ntv/v/9jeLQvfCcqlI3QT8zPeBPwGj0Yd9cZiRusKXTsEQUkIrc2Z8f+YdSiEpGtgg7m/FIttX
xYD2uW5ORnvK8mlqMYJnMRO/DgP2Spjm5Tnb/Ee8g7mw2z7tSZHyFsqGaYCQQ7aRCx2bcx3XW/cq
XR+tM2dJw6CKa/Dm19pyg636w5UhU4lW6FVQxF9YDRVr+9cjOfz9MnaYrftGYHRRJil2ZrLxrJQM
Ww5dAG7X0hQBMIsQhC12weAybsstCwMwnv5chLilX/un7BS3mRkjfOvWHLH+FQxyczM3c2IODBgr
b/cF3gjm7jSZDsxjA7s53celoEUxZO+nj671yYVDDcKnycbkpTrC4LD+GboFjtkjj/wOvtUi9ZSg
XXYDbgdwPrxBRawg5CWV7s9amlAlXBYtOBs+bILxqIbzaUO1KNnaKC1tS8JmLSYmx+ykzImivUS0
7YPeUBTbveiG5OMivu+UEEd4lyGgUmWdvM2r8Odod5Niv+k6pX9FFzEdwrzKtwEmjPYoMhymhCVM
a3v5RIyVTurcta8bLJ5FeZsS9n4Au3r/rFi7FdMHDXPwtJC1f9/aVH8kqyLE/+VlXgzBJZTAi4fI
kO5dcVngimINigPuDxB+MyhvApAvnvCEsyp83mbNad/RE/cFyAekOhZxXz6pYEgjZVgHWht0nnyl
PHWUgbect2oXWkZ8wY/CNydpvSUcoUfwWXMFQixzogh7rIue1SNZM7qIePjfRWlABVmGjFXyXDBk
9olQukP2pe61jPGYBIDpKCCrmyn6HPBj6eRVRqEkZoB+WkTgyQzp0NY75gfFQ0+HFkdNa/JPcWFC
A/BsgOiiqENJoUXMPKXq3iVhpNCDPd/5VSTIuXPC4sI1r35wJZsUC++rkSok9Vg4sFqv58N/LMgt
sHpvEIP5Y5VSRXi1SHUSBdMnXrqdxVHgwCOZYgJQ/ritLFw+eD9wE+gyXLDmrmyloc5ZN5vIeMql
xRC4s7g/eKL4JdH1WWU+FgEfJPjnlv6Rle3kQmSfELGwjncs3xeMTLZgLmvMh7eQGlrhYswyhHZk
bOIBDmEJCj73IGouQy9BxmUUg9aY2dsRQPgflnXbJzQP9kD0zKhpA/oBBTXg6ZRRcsrv/g+caUur
eflPTmEtVnczQhlCcRz9awjIK9U22MvzRVw/lID2gliu9YDxDZpLp42z4jIQ3BZ19AyCh1SfoqkT
0yxzgUBDFxvIh3Rgsb2uTF6VOZ/SqG4kOtIOcCYpEZkd8w78wiRX8Tw0nfPJTcIHat86snnKtyOO
L5sm4eZVYyQAle7cYJMDY9ZwJhMYPVtSIcDPrmVNSeNlcawvfHkX+fMF/dNeHhcu/GebjOwgCRnn
q7Z0GjUj8agQRs9LFEDa2MFwyJH99X4izNQZszjCLAZasjt/O58NuAYOw9uoZl8yRvyZb0ij/GXL
BEY/wjwNMUF2dzYXLt/ABYN0LX/LI4gBAyPS70FIUZJC7g+W1gURuVP3KaM057s3tUrDx89rDE2l
fWs/rMMws8sd/F5TRDUUZqZbPWPhdK1cLu57hsMCFZL2RIvnVuMgG8nb/DeyNjiMzRD5XzXYvMbg
fwPgoeML81xCSujifvgx4gMOd4katy/DZvGrEU4KNNpb9E3fIec4yr0k1Q58q+o6lmcQ2pQLluIr
PGSVTm0P1B9rb11imH12nLHL6b3Q2mw7Cr83rsU9VGqyI8sw68EcoidLdQhthW2Wx9fl5xUiRcof
1bXRhMsYsIlqx1vrq2vphcanTE0UkLD58/VyUnbp0SERtP9NY+VQ5Owv0oCMtjn94Gcc6e+VHQlR
36iSUAxf63B5IYPA3enn3n8gO5fBd/WSQtxK7GqmfXfhy+WLJ9wQ6EuuHBDdK8B935kw/LP6OL23
EXc+ZVIrNKknt2V/wviYIHJfamEB57/e/FkWFd+Sm1R0ncHKOJFVraoMKYWjbrFOIfdFVOYp6t78
WIlb6Z9yDlKCpHHvN5j6YwVxc1xIJLGIFN3AW9DSCeaDW+NK0ELV0kPzJyAfulDXEgaH3DMhEx9A
6Bu7r9qmxNcZPYPPOF52Idiq/k1++gK+SjNQfMKUmGlxtPwrZAeXs0oUsz6Qf8hsTaVq+40J91i6
F7Ha7+PfPW7uAZ/xwKumvHQlvP9lu0+glGcbEEL53FEtoupmS8Hd2jdIsi4Ent9jeOQjWtvTjQiT
B2dGNQ799UtRi+VfzpS7//k/P+Sgsa5kfthEFC0fjZz3W+3g6tzB30m9b+5oYoeK9ClLrgAI5dJd
DItFlytlIxmMuDOiyh5xL8l2ilRZ1tILWImygIbcvDes78INHjf/R9E4odjAMFZqWy+FymkT+jYB
/4+SVqAWr3oaHxhaDNYxpQMCgyFmFfBf7QjEXoeqc9O3aD8fJWmrCRShqAZtop8wPjaLHQyA7pKG
QlgWn+tLKq+bF5hRiNr0OArgapmhMC9D0FvykqG6khRmBwsuZ9+TDcrsw2YY+eL5mUmR7Z4ay7Uo
9HmCSOHU+8JjyO6hqIlkLvFJRKLZRnwv7L3OKO4fwfHXY0/BEiWHen377DnuCxVUbZR/QKPrIJAE
tg+JI1WjStX+XlwbbhJm0q2zTxkrPtE99yIlTcQBKkStqATsp/s4YgaHD47q6tdq308luw53RxzN
0ilEigbljRVUGZWTT5EcJDOjO5DluAY6sWQpwWmj0/fOJFMkq25QGy/N0fUX8n9EzbLiZKQ3Wyz+
5jp/3DruYX8FZhdN42oakAHO0sHuw+XU+CpiYoICiDiSKjeu6SOZaC2WJcmIv7g6Vk4ONaLOoPVF
dV6FiRWFNZsHtMCCwWANMKwvoBh/it0/C+lLOvy9u02swoiKUa+f+O+pkP9HePdBk/jXu2+CSoL2
gnU8yMdDMP9KhEX/0fN20leg3pZEoLeAHo3Tujd1e2KhfkzPfxG0YWGUDw8Txagzpf+nT87CP1GQ
utWhwW6RRcMYCLzHiIrsc+TABBYXrOLWiMp3m1yeWf2+SSvEveJzTMov6sr1oEKqJVbD+yMweIsV
kRDVpMVFQd4rtEz+dU1x6oyvf99av2bSwEfcG/JLICKQX1yh2wvy7/oYNlk+TbTJNt28XwEVSIKp
mAytpY2I5xD1B9Zjk0SOGg/vTFOvmwEesZB85zlkMLFh8Tj+30z/ZAnrioj118pafXbf9oOCppw3
Qvm8nstyxsJOZqTj3JSRw1ZiXS3aavMAR9nCWSCI57za+rx+G8x83SowRoVBzssfM7xhVHHylX2g
KpOXOaABfl8fmKKB+TTccvPRFbDtQ7nW/W1JR8KqmtNLSjz+bEIIzj4fqfXF+gXwDTyuRCG2D0uf
08oqvYRS7LZmR2N7B4MBSrZRlbBPZZMCwACyOeNsrQDptS4BTZLC5mDYchgE3yP3ocSfE0k4kBkU
/X1c8+55lzPK+piXyu2VuqVDbjZtJNEsHh5kI40M/rEA4v8dkCAqdc5PLyYAfd5/ox+egS6QPDHA
YSuvlaiUAD10O1TIfoxb1WylI7317E1Qt1GAa4528koO2iq4YS+V7KVoICoI7vXymHmfnLR3xV4A
FadwPUqINPZZq/YMhatrjyhmempr8A4IFK11hI9RyAM4NpcTnfV4TGsd5S2sQK3dr7Keg7TsqANY
047lrpHIkEfXYGrTmPfe/M5bmyasQLgcbUR7I6NlN4ZShAdOJMIcBpnqYwwDpxcDyWbviiULd7Zd
QFVjOKseWYmeJxe6EmDv1iK+mUxX6E6+etERjNAUKnsmbNE/f9ESU9fgh7VQkIcek+q76W8AEIri
yH6yOJiWXo6WatIzCDMG2zxY7jbXTssz4/PpufgC2gzU1UR0NLjlrnuT70V5gFQMYWw3URmim9aG
iM79zAWT4kdoWsy/i5CW4a7qulXhqdiDzbJXJFKcFcrzIVRZJSMgCQJPtgyC3EgRF5RuvkipGZwJ
ZNcFEJEZja2jN4SwTqDpQ9/iBIUU4oS+Vq2CaW6O95RsQbO7Ypw0hHEWU7I07Ab6pXa9IvkPTubF
wYYxMaluYTvbDem4KQU41StMfPYGJmzGN61/9zBWU/sH+1AerbkslMEVY+pUW8ztAfjplRftrnw1
kAmNkVx0gVjxOr8l78gNuobIdlK/67s5/wD4LrsgTcprpEVPAxW3/RA58cQZANJjCxnRJPxQBAKQ
4u/hKQxVJ0KfFXulk1mZZOCyABKAdKk5m9TSphU2jaZMw5xE8vQihLpDVQkBLadgAlsH5jKH6+Iy
c4Gy1tA97ePKBJbrHyx2u8pIsCaVAMxJSCRvE/sx9M+Kj1M+AD/sFx0F5MqRcsh4bdFc6oResuA5
UJAeHlN9ys0vnrpvHYihILi1ua3IV/tn33loRtW0n2rmu+eYkqCplwfj5nVSP58FTUkQZFnRxF7A
+iUjUoha/sVL4A8cDLlq0uvzU/hYP/yUrZ+0YMPCBOQHKUmMjYQc05SiKYS2nUtzXlbzbe4diJoJ
2/1f9VAwcjuNuerZd5WUGh3dj/x42WF80foTJiD8eGx/n2T4sxZbx6/epuO00sfat0fK9OYCPhX2
Omsd7TWz2mFShH/TfWvnGyxZtShX9bU/PpFjRd3vL2OgVoEiHWQUe+uW1JZYcvVx/BePgAkWol+0
qRitueY2LCCTXy1x8ETkzQy4GxdtJ0dDevjIB8rTTH7I2daQQhGwuqZSpoFOhDsjub+Xc3V1/vcy
oO8z1B62B+m3UQdyMX+wUGnsplq0ExlibuHwZoU0KPDb9xMbHOsaOF3zLBFbdn4JwkT8UGlNRacG
tzqXtG48niyneMlt6oGHqZCh+/5xDm8nWG63QiXrJVxWDpoqUM0wytyLSO315ow+xBYxFEVz610t
42HVvdHIDlFVTmzv87Eddd4Lnoex/huVaQjlbPsM4FxPEilPjPNRjaXulBuW+tn2kOAIYC7eV9n/
Vez6NB+5qUvuXaDJtMImvc691V3uQDb6jVlVlsRxVrHMopcd8zpITXy37WsTeL9aKbxsjJ/YPHuZ
UOkjXDMls2ViCSLqV4vjrKtLmv2EbtDVVlyemnpw3Up5UWaIlmSzk4/x4xDU1TEmfwST9T17cc86
s3KqXNtD4Kk01XUZrQzdm3YY2FShBGmjDTW43Pe95p8yns1wYntpd3ljxvZjMOTr5uXCTVbBVDTN
NHV7lp5RYHZaOfYV1+/ep1rV0og774torC9G+lh35sE4UZ97LD6/AzE+vkvi6ujqJ816huWO9x2N
oKPIMY7xskuQzVDGibl3hXEp8GmgIHGz9N84OB0/Qph1yrcOvuB/nRz099xOP+iLZ9DHvw7Ksg0b
Wj1N7Cr4rnhGFer8MYe1dmfQgKdpfMkrKsNjXFYDUzQPed+ecicrY/G97PAEQ/M5B2S/vnkUU+Os
NutbT67RaotufNhP8aAX9T/wfcFMGnhjl7uXe1Ma1gFPbQnuzTufoLJ3BcOAdnydWVjL4UwMsBOA
+BzUpL0uUmaodl/fxzyLpoQrtTn7yzWPx2Jw4jV+RnGorSDbLAzGQ9sdGOGR3g9WbmdNJViVb/AE
9RsscPDRVgHPDNLISOrLCoYveKs1aL84U38zDhANr41wA4i2UlkyxVdJrjzHFjPH5eNqmilvo4Lp
YKiUiBLaBRJNL/0NkzrvKcpX6Op2gJduGm22q+shYWxp8i5DmkIR0myssW/AzBEk0Tl2x6zS2xea
SnMSanW5ut24D/rM4WlM7PS7yfyNEYKGvphcf+KZXo1N782AxWwErs33KDqFDRQw1SxwaWgbuMJu
Eo3lpRvO51NluPu35ZE3254WJIWqJXTxPZ0UA28WWmSVpcW36VLNE0Yah3UAaU2r5NF/wYvThGM7
bkHxoIpD3zEaiZRvukoP5+MKNOqjQEcIYAgxmh2pvVfR2Zv463vrrFBC5I2ILfQers6zb1UADz0b
9g5s9j6WOTETw/vtfwd1yLfUW/bQcBKwMaXX379Q2FhweuEfgRJmxotPlOeaMzwyvhCwK3yr18sw
1g1fUoV1X8IHrpgArdX4OG3Hm83bfnnMbWAyasjoqKBglcosq8xgiAp5QxpaAfwBHaohFMM9Bk+c
DcavWPd9LDFWj0Fyd0U8bmGJLEhSlavXIUGDVKY0BwkpOupntC4wcnGquySvcxo3FgP/tPZ9UJwx
F8mkxgSANR/HtclHzYF69wPxlFcHqkhzna/IeBQyP4ofAJvEeGU6Xd48WNM0xYMYad6bkw36ay/2
/zSgyWcfIqETTaEafW71xjtrfWSnLTyUGVQbr+uqQjFE5l3g3IssZrjY8l2biJ9iVYCMkQc2B8jC
RK/slmfzrj7y7Am9CtvgDx91W2u50oc01iANO/uRCbGaikO7avxNUX8kIerE/WHt/O4Q1GhHdf/k
gMxImbC5u4upIaV/bTbhNDpD2267HWncOwPVPIx0I6UIYwNgZ2m7fXPpTe/iti2c/UruCMXU+6gH
25t16LVqH2hSAoUTg7qsJzoouh7m35i5CcXK8gHbByKljMDafV6XNtVE4CeweWNAQb1Dk5tu6lAi
wjOhAkGwWGmk71KFQIN+aoqzeIuwsU0HQfZQDZNip6ybRhgD78kyY8UVVnA5zg5aE0nBIsZ34wCB
vVl8hJ04JY/gUy7ZqVmmM6J5l+SK3v96PtwAFWMu7jNcl08G7urWanGJjOaencZQEOBE/boOZyjy
71wmcmYkKB9Vsrt8zmySRNQYszHO7F6T2GxtiU/6R1DNdIm4Ml2ojc2nh946Wb+Zdy0TUHj+DsvH
z51HDyV0nVuVrDVznqTCJ5YjTHgVMC6PaaEjbq0302RR2Pcl3ZPrTjdo01j8wo0zo4vSxXnyWYW/
FkHGyySWLr/N4w8uAeF6EVL01hiQ6qXq2fPgAOzKjvHE3DoK3JGYLYxXkYQHw3k0Jl3Bn808pSiG
T+5PvoqUe6tkJVO8r1xwyaBiiCkMvH4jMLwwhM0zyMHTs48KESCW8XLoiv/eo2b4617cu8kgHM+5
zSRqi+qpHftzJl+ro4eoWoO3e83PeGnt9i4L3bDTwDSs/Pwa7qhqFxdR61PrwkNmdHiV6tgaMFu+
TbhoEGyJj2QgWr3mAbvONcK5iFGlfrEY5Gu3WCNYpg96fWFf6JItga7ZnbeDSo05E7Y2njBeWnyV
Ci4CXOINQYY+EAms7na33xmMPIRoBT+Wpij6h5YyRZ9Ifs48oji3JpuJPI3RsuT4d22SE5gnjv1L
8gdMaRVcc4yraAoore0jrYcUITJd6abdshIP8YyEt+8kONyKoXi161AmXKWbxZbA3j3HtVgy5qpo
5H+jk7xR0bAxrYPxvn35GBAYI1Ww1mIkt8WLc+GZFcGZcZuefsAuHWKT/ewnw9SPn19/zrZPlQyW
rZoX8rIjRDRCIDFhTJUxwkM+x2VQsaqgedsZq7bFyzpW13xufy9pP5/g30xN6dvLB7fQWaG5L1OM
iCTnGx2oic+98WXZHaiGaqWaK0Ef3SAsWU7ak4UnGrGFQb7nCWZNLoyblIRwUzLCYuG7U3qnOxm9
byCpE/m+wwyTloRU7CGP1LA0M1uY5/wN7taiXt9iijV7CklEbttvVXkxWfOy8kUetaa3CN2Y6Qje
HFBQhroQEW2HlqIZb0qeRmGCHNq5ABd9Lp2VRCvkXndsb6Q85XXd4q4fJq0UzvuflRgvNeCcrU6d
Y/WEisVEGCzzuzw9SOvQzwmX10QOuK3QuHgGRs9iS8n/dsI+9TRZ4YeWZSSzy/DMVMse539l6WzM
49zdP21H64IMJm03i/SHF0GilkP+T+Y24rw1T0CpkBj314fYoyVYyIvrg+TvI11IgKBWqwlr0tIa
hSP8rG4FRcZPQtdYtVJl1mpi4eysE2hjq8RUOj+SNSzmHnrwQPJYZ0ZIsgt1MDwmrsPTrWCfn9g4
PBl+WXywtfx7RpO9C7hIPRtTHHHti42S8syjaYEwJx9QuGyggChhKen7unH5gm8RlhINlEMkcUQn
FzpwFSinZiqBd6hPCB7SvnRt/ulxhfyV+4KTHuNpNNE2NPKBunE2iwBRhfVYtMo1x7JZEo6SGg6J
1l9OM5c4mjYX+ukdOMUqYXZqHMU8C/QdtP52McgNJdvo8nFnxXU7o/zRTeTncPt+P2WDvTEqnLqc
VISHRByC6I5i2buohNX4Ne/msmnemDoWlFypAGLsTjZYixn2nlOy9Lt+XkcqoXGNEUJ4T1x/xSCt
I99rc5FGP5p/30UeHEqSyUQpCf6HALXJ2SM+wHnUnD7oAeJl3gqTpBmOx8zP1pgFHotdzdL4sEWI
F2oeF65DTu6wKe+u0O32lwxk/GAqV+kOEaMrJFvgpFnB2iyW6QMTS2UqCXWMbIy8y5DA6vi7n7Pl
b4mvXonKBOyuMf65F/s53lJLMe7o1Y4qS6+3eLfJgvKMghm2+9WdUikY13afCbxCNDJeyq4EOlGS
GdqeomRTIBbZCopDLvYAVlZvvFc69HPk3zf/E4GB2gu0nAs74at7th7nyneD2jPM+YCRR1/lsSln
BxLdeQCFeiY7f4YTLegEGoFMR+6N6wZerz1aXDvsJe/NlxCmkrc8Ln2WZ3xFgYoorDotWD+LFR3t
ixsWU8rSDhl9yZMV2GPyN/0uKDrSO9OzUsMxJY9HwL+4pDmqxjvjFr+r8H8ruP2p6FwOAnGWrNA6
/ufpUFBKZHZsbu8k6GFkCCeTIS29ru1igvnRIcKUtKncwUaJDcExoEnXjq6fhtUv1fU9fx0FD3TJ
hMsi7wIZ3A1fXM9jz83lUZwINa4ah0l+acOA9dFJDwGoScOv/wQ3hVL1gK7oMo33T8gL4gcGeALa
H6sUULHMT+cSq7BPU+3TWYgRNJadeO7S1eJxgL8Y4nVMHE63aTy5g1Ei0z1azUWSx1mB2sKj64ox
FiuBoweq8UIO5VC3/S0a/cacO15668XhBOg0Z9Lq1mGTQ3mj6t1HTA6bHDzxLqn/VCr8A1W3vvNc
LZxifEL+P4eGLWXUeItnh1+3+c/gYMvpdp8qhVIGXhmayBg3xIp6BxTE+gWlbcuuldTLcNk+fyc0
yHF4MWPSMGRoo1pY1cP1XKdNYy2UCmvycla9GTyeP68dSt7ry+S4IliCnYOHzl5N0N0Vbcosx5tW
cuybfF3bpU4rIUW1mGNakcLnkzi0YTN3Mvfvmpf5ndcc2X3t6C2N937mNZhnXFkWNHq1wF+rdcQA
bgrJvpEdYLQ2UskGJQQxdmKdXMcc8WBDjXW85A92QqSFEmW12BWczc8vz2aIPCcUpsfqE6NanjI5
aWttlRgg6fmPit8i/QXuyRBIJsx7Dlj8a0X/cJfk4UnqNXW3YMGtiFQ8l90drIi+QguZIABsXRRm
jFSRHSYjd6bjPHk4lXoR6vPQ0sehtnhvb7XdwfdFWugdr5NKQ2b5i1jMEcWuPHwveZB05cSTR5qV
i3GUgjYhH89OAPkwvh5rRtbFoIrVaL6xOCg3a57vOHsqBkLrO66dIpuFDTV9AC2phmOfS2NwJvFc
zCskJ2du37e/g49ToyMTX5tLz1E6cM9QE8aiGMWphRfU4orwJhX1ZTyh5ax3wXkS7EY6S7nbGdKn
6ngT7Iil+9rd3sKi97vV75ZOo2SYLAkpn/BowXVxJVesjcl60r4jW1OU6BKTxfIfDlZ3NqFUpQ1v
wK/vY6jlB6Yvq1IY8SOukdjMLtOdJAgF3x/SGTS2Ykxz9PvjXUuW0ivBRq7BdKQlidgeG8wkbSTJ
/TZY+sGbS9k+iT2r3jYgXwLmhc4co5eP9aToknz0rOz8rDJioqpTkUpTsEtn1hVqea+VuQCrUxLl
iwm64nFwMenKGVK8brFn81LsnagwDL6BDq/14DHmWzdYzdihZ17CavwR7LmLqdI1RQISWBs7Rzom
/k8N5FCvO//VyK/eN1kP2hmpYksOrRNRKrzdwW02/GRcGKBmyCgWHI1S6jkVWusR/RXev4eTqvAZ
18+3NEKFXfuOaxaMOFJcUL94zIUBvO0VmED+iXZ0bTS8EKiXxUoa/A3mYOUCepzGObVXD98Vs9ED
ZIPH2pparAHvs8kn/EpillJg6+pPgEZtKEbJ/GSbV5feldEfWXL6cRoXC9rL4VdOP33oD/cycwGL
ue75ueE8/aFavQ3v1Od5+FbmYw+zdIy0f2e5omdBHGOlvTzR6r1urGInx0MPGDcPBI4Fb2NU4sKy
DT+yrmOAaDtzKi3i4uXoPv+4wdipENdwA03Tdt0Kc6rT7OxaaLFLZYiBGO095f33FUfLQgbtJ0bH
q7EZmCtFq0LXdlru1WraCUS2Vvr0nmeodjf7zuuh2PF3NPISwFqrHIAYUyEMEPcNGATfAq/PIg2S
uWSLfrh2t1cuVRBSm5lBUvq4hM32L1ue8VPPTkkEBowDhi49A6Pp7qzIeaRoaasuL3TytFeNA1xe
j7HwF6y4VdWTMY3mbwkUBVArvE4W4YgWXKUEv/iBpKaX7wNWMzTqqs4RqjouHHY/2gezsD7hGXx4
9sOTcA5ROsCph9JwP51OjjSd+uvqyYE/nhR2lSa5GBnwW43BzDinlrROvXN8hcebO17N0gbc3AWO
ffF+u3zdfW+AfSosknCZEiNXc9+Yq5QO6D/d/0v/EMhcHl+Q34XElbr0u5BSOScU7RhrMH3hlgeG
VVdF+O6p63AQh5aWuilxfRqln1WE+XhP/La3VyMEUsJEenaJ/B87ZoibSRvs3gZPVSeNyYi7so1v
yqrAQW9rKt//mhNTiPSHkko//n+LOLKb0rRd/BulLt61KcIojv1OPBroIy1rpsuHsmePU5wEagxS
cZ+ugkWBYzNpZ6J/XCvYo1QLM+mEa0biKHcZDfMOOVoFZMaZrjcpf0nAI3/vqVN4kXYZpbk7t2Px
ZdtSjqHkejnRuBCP29O2CKtYoWLn1Jm4fo3a8dqWIRf3nnRLuLUZk6Tyiq4FJXgQCUKmJXNJxzXD
5SQ2dtj+kmE3qxS5eZptPYFf6gQpRUX/BC/dLNF0d2APCPesvm7ZTWKKaDAe1ozdhv6Vt1ky8BC2
VVSTB4xTOCEosFeGxUCzZZFHc+co0AyCSlcgp9Wmmk3f9FJE/qzIpI6i7BLKzRcI96FeSctGC7jh
XiyyToBLYQloN/VDQhItpd7NOJBZf1aXTzlvFjgPEOhkgK2hz66Sxne84WS3hu1sTbVlb6jScTzu
c3VyfH9jbsDvSwg8+nyQji0xNGzZ8bKHwAN3n/KTj65c4iW8SVcd5mysVEPb/rnSEdUznASiHV6H
ZxBDcwU6U82ElxHSPdaUNVh2cRYHH05GNr5wddd1UpQB8Pb6Xjk21uvy8Lmqd2U5vNLcKLfGzEJq
Vzqeyjl0H72X2bzbfJ8nT8HCNscI7Y04KUNhht47SwwczuObNMC7l3Y2N/d3+Pw35VAku/oSjZ9X
W48cALJsR4Kg81Oe9vnLeZF0AAzdHhqpQ2T1wF2mIDwN97TPTFzIirJlYHo+58i8clVobUaptBW4
2v6z2pn7kFd+rqTOwKEqHmf49IF0KRuzRo8Gnj7dnVCVAdUdc6kHObhAMwAA7Opo337oEM3JHN8q
nuZCEnMIoL3wL8e5rpwAD/TJz3gEl1qZyeb2ijj9tf0P0+lW6FGbISxlClMQpOmPXNiYTIXPPGLS
foNI0E4Gjq+iryWh5SBwej72fDN9b5Dxvub+Pfl3PZl+FA/00jzwN2dcZKMIgaOZVQ2G1dh9KMSF
/vc5cYALWjaoAXK1yUwuXK+XQ7QntRWEKBo21eAYsY6LqOpVcqZP3gzQHc7eN8ruTVRFQwJ087Q8
7HwBFE96nYZjXjYmO91i0AwxsqjC4476aQ2nb3ZBeg3V/rLWUylD3+cobGwBFJIMYYPSlVEIqAor
PTKlPpgASk+hiNuss+X8Z+dPvspWI8ogB+H3UyFpRmMud+rCo5pEQds/EPZIFamoEV85cmSUtR4N
/FvdRGfFoSY5RUr+uSTWNSWXdnfQfIxG2xxGItFOUH45M0Ua3ADUoIM4S1IsZ0aye0iHJTe2AI6V
B1YPqgwbk14RyiFSNCd78ZqZL5l4Be8z+TI2dfzgJssoh88AVNlX90pAP7n97cnwmDU/QXimJV1c
1AJ3W4ktnHeoP4C7f4Ix/5CzttwaAheMdukk9lc7dIrFVTJGC5RfvWy7ixEmjtXq62BSfiwSR424
cXTbyK7OQBCAGtST/eyxPKFfAE4eYcSM37OYvcFSpef5Qv+7RRWrmd7NysvXrmDPfEWzpSYH5sdl
n5t+T0NiB7gA/u3PXH/1e+85/kwWZMIECOLeU8UfPOxXulUSY7VRYtOoPdwiKLbgL35K15wktzb6
lVD8prFCCbfe2oarXyknFNLbdEdoqnYCDEZlBv7BjiSlBVR6UyixKIWTCqoBOkHYZlPOwk0uqpGQ
3IjvQodlXnC4Z+64u+KW4YJpT95zeoMSZ1FSiy0YnLdbBm1kIku29HPxUea/IHPNmneNdgLnkAiB
OVflOv4EgLuhW61A69LG22K5HzdGi7zxyKkqY0v3BjDdCOiK+CSSzL8614ZccwRfZnRrm2TklEIE
aE7LO4u7OMrDHBR9iaM32aTV4VzJBqSJbdeBhI3C90ZzrXT/MJcTyPZz/dLM/ONssAkNWoY36g0H
tcnDC0CREoAR35ujjHbD6RXO6/hNzWaZwJt0DjZqF0JbUfeqrNS9I0NFtV80oDGFXNU5gYdc5Vse
Tat1FezAbVFlPgk2GZkiqjYomSSyByZfIA1UsP6W0ofgmfz29aVqHeuCpE+iDllEsisMIhy9pIQn
uQDGK5pT29jZmctNRO7fgzfqXcuQph2v231/IuLaWTD+sXHC04KB1N5GjS8IfvbOO0//XCj7dL1i
BHiLaqWjo1Eu5fF+jvd6WHuCmKVV4cXbppyHkOhFRDpBeBNlv+CWUhgUdPoCyf2l4S/PODcs1zhq
owpBl1CWaTiXP7sJ6SYMooVsTJLWdxUbEEwj+rGqYHShuXqvi/OLx5n+4dpfANPsV6NudQL7+Jt6
CodIpZDJOmwyHcUyG6juRsjXVix1xBlV4Y0kd7oDVhC2MIYNMdINdsFLD8HMSOvEUAgdS9YpO2PR
yZ9dv8IRFqkyva99Q9qOsCPFiRKk7xxPoyhmK0KG0u3mornqBHMXbZNJfJvHHzMmnPabNEYUIYkQ
s66HmqYJC0BqQs+cYtmJ61OPqfq3YLxY3o2QcwpP+08kfeKPeQ0IWmYhUEM28ctWpsyBtFcFhn1m
16miEiuM6mnl1fWlcoh/276H8FcKDX1/FqAsyvjpXtCF5KfHtvBElPtA06MJf2qz8FhdgCgvrUbq
3V08IJa/FXn9CmE6QPbDlHDOzHYkXR56Ws4ZFdBb/JagF9XD3Ddc2HHjGqRxN5oTqNgChIsR7ofj
0x6yiMol0/ePZreNZaIBdJPIcuy7CXWskWdBgdJGwdSfCr1VKSCffN/2CNpGDcOuotSAq7T4pISS
A0iTb6n9qPGEZaS4Znea0AyDw+6B3j50sQMQP2HwB2UQGSJEwwphOsPwoxerMozcVPvy4KTfdhQG
CL+LV5aLrMmGFODtoJOxvUorzCAWf6GTuVqPahpvN1ZqhMiccLT8y7awPc8zDI9UVpxfnYBYDygq
wir4HL2gg+SU7YzM8teflbo4NoYXN3uFQadUGOq2DH5LyxMCwtZzksdPEsQVal1e8Vng2eLfK9GU
b2jL6H64mZJSVBRih7Y7WMiO6u5lTRABYlcldleyP8SavLMlCRLgyHbnrspBsGGz5mMe1pXhJvmz
u2IxnduiocXpRvbicgUvxBHEycGDBiHdZ5VuGQhkYsSRnSOC/VTJYm3pECo96VOdmH/kfuEWE5Xe
Is4BYPgb6fqiSqeS7i1qLtnuadDjCQZjNOcwAVXSfzDNUtr+rIryyZg4xeWy3v74gHw/CcxsV/YH
R7ZSc5TzZ9x7Rhws06ntM6wBFuH6jfr2W8KXNBXm5/XMNcPAoCF8pociayVFKcXKj5WNezQObn9q
Y0z2T9IcB2eb1FpywhsftkN5QnNpB1Dvs18oZJK2lJ9/r8wMgxgpbdlSV1IcmCnMP38jujW+iY+a
MOGuMOMVDdcBhpJMMgQlnGsEEa84iW6zrG0CITBR1xJH8rvjRWl1x8pdlYsFDEzdnNNuAVpSp3Hh
C0ESIe/91J7eqdjC+gjgiY1DjBhtdg20ws8b9gL1v4ujgszLaHDkRbbfe9Pmdchtda/HVB8LxBho
R87FuYS1qadhnxmgAzdvplTE6KgxskDskh3d95PiHsnj0gsZ/MLsgIqBj85L34nYtGjrO61clNv6
/4jclPKCxzyHA2whJ8osbv3gWDld8Ockk5TperVzfjV29MKhDMG9EAKtSeoJdklPaDx6b7FMdr+P
lJ84c4LN2KZp0iIwnF2ql5N18RNvPlNlwsq8c+t+5lL9ZancJwufpGWadY7DN7/lC0JwGR6SiSVi
RwXeZ8dZ3cn7bkbXQoz26X9jWt+DMikptaVn2PdXaqq5D+pxIsJagdS318aTyuWmCY+QsWRIo3MI
p/lHmz0Gey5ePk9KtuD3XY0BrvW9KEONrpTw41Je0NnR2G7I4IBeS3oNkvIAjhLwdVMt/3Ry3Hfu
3sgb3q5f6VFodaBbogOdFAPB9EF1Tzo9SEpEaEtcRcpWSMIi7TLS27A1QbXZodpgf+Joo1oXJsmn
xyBHXVscnqnfmEZT7cXeqW1dKObGz720hQn23zSyBlUvG/OVDd+bzzdQonKoLi7QnveTS+DspjGO
GQ8/JiJ3em0vjGaErGSI3+UXXaz1t0620+FEGcA7oM7+evt44kI8q0+R6loQzPrevaXWXp9BneBt
AiiE3g0VoSr2kdRpqhWxRs17HR6Xv1wDmTOuNJLIg2wSBZzPAATyLtFJ127jGXnb35/vre4l843s
c9LCkg8jJ/uZGyEjBG6j7SRqYeRBj/FhtqGCEDABpclxpw5GDJGgayJCP4gLZMNJiDKwqbgOSdFO
GbI94WeB2IMRsp5g611DcIV3ZQR16R8K7R6owisK2mtuI3ELAOqtXeC1rHbwvy/+IoVGHBqhRHad
0IqNsf5gQ9Zaxk796G1PngvQbESUVphYbnjIOlfgTmPm/ruYpmNGl8WSm/zFOdZv1x5Y5j0dQPbW
XiU4i2RKPebxfrVp1MoVRec0rrhwG8qr43BhH+f3S/dcyKHCr9697Yhf/WgYQtg4fU9l6c4dhN4c
jJPJUkSisSumYYIgsj12prsvaCn2DH1W/uf7T7M9zkCk87Q7ltOWCHG64zIADyUEUb07EPX+QuR8
wsELujP9sFnBCSP7Y4ZuOABEdpmyG2K2u84ouep8yIJQe6RV20x6rkNk5ESkytlazvb9ED87vwjx
HgB4o92JlSpJ5qWJ+F0wrTSOWo7TD+oyMqvaKTc3xOaUvIsnIfUsEhfoqwraqngEzeWg5KHX6NF3
/Me8lmdIxXqkvY0UnRzVr5cuV6JiMB4RZOAeI+0tX+VtENkp21b9y2y60nq6/nx+EfkfpV10e+eL
fl4qvSLGKbDTe6I7rsM+47CHELXdsbnxieeDymQPg2mqP2yzHGwA4NxxHq43q8zzXHmA5+AFMJSR
sF4mvYfqR9WyOoUeGp76fFWoH6FeTrEYuurJqWXGu5S6qjhJH799ONVoN542nHsEiRYxfbZ9zWLX
CHSvR2jMbV6bsDfpIJ8TnLypJAM0tN/lqy9nAgbxRHJ6Hc6/Sfbe55JbJLeYGSeiAHsyfGW/rxJY
IM4ZavromWV9tXnMUbeVOxDu0ZXKtea7Y5thV3jEbFrm0h8QYT9p241dTpH4iE0skZj03hkaoKDh
a+5MAZxu1SedUywtTYVC5JBn3hTr4G+k/7NM3ZSTBtHxDoLoAIQTkqpjz1IbkE9Y1M2bEqnlWC/q
NTr+BP5q6JCpvimCSY5Nrrme6W1sJmVgyaz9mMaRjQAU86oJbmZRsZHL/iCk3WQWZGMXni6qHGZV
lCUA/7tJztYcNlylA+VnbBUKUmuwKiuJVJGvkHVADBuHBUcAuMdNOZUlzp2GyNJlvr7RjkzoNYHw
Was6RsluazKrki82pTZVfaQeppCFmSLkx9i9M+nURXmtHHzMVFujblLVbLNTAoBFDWggZMGX291Z
8AATE8dNDx5tlOjN4QUW/uWgbMiy86l+AbTeyNvjzaZy42xpU9PxxSs+uma21LBUowaEIq+HQ6ba
vYVpZlPsPC5ETdQtk1/hsatdXBfPHjkH59Ib2G9Y+PF7/9nA8+o3u2trgPmBv/mPI9bLz9J8ETrQ
DXPn4IZ/WFYiw1HlNml9QTxdzN14tRJQXOKafI72uKNQIXI6ItvXGibJ196fn+OZyGJzq8HMf+oG
JMzcovvxbl00DW3wLVFMIT9CL4tcJemrQV10gWLbtCTcHABmBx81UH9fdUX4ao6aowy7frbZpn95
RM0Ra4ZSZm9id+XP8hgkjO5QpotGcVI0kP2rphMgzhKtVuVLl7jJiDTbvaIdLDGl7yzaDearw2m5
2PEuTCRoGMIH6YcEZz7Pb7i2yjmRQ7roM/5pZ8ww+pwnXGptNcrOR4X4eqqDbtoP7rCWhYPvhAs7
MNJmOt6hdHEaFwiUy6905IK79ZFiJ7PbpXp5Jgj6Acn8lXva/sUJ1deHUfFPkUagdvgW5o8LrOew
gc3T1sMuj71bbd4vlxT/Zf25SWU7q8Znl+h4HgbDiKy+UPmudmfQPi1tzzg0JlJ2yc16nPGbZqCk
mrjkWpxBaO/MhS8+98VFTYIfpynCDk7QyljQexo7bET2o5m8hEHZali11PR8uN69esWhUImnr8B4
rS2OtcI2LrIVTh2ksKhhlRYL9jiu0G8EegxtCdQUoRgjNwio9VeOGh9vZpkZFEZo4bqc5ae6hXMR
AO9JrFHXkIwysVjjWsrs9Uz1puYG7Kb4AG8R5AX0TpbnH1sHc0BivLq8D8VeuL4ar1jVX/0Hwjse
C+zdP51SyTVrCCZ5fic/u7kNJhCX3kCvFxdIx3XyapgNtAHziGNnOtos8QXmSihSkLlErXhxMUFI
2vACHmnWdMzAYhitbc/j9w2OJGzQlMM2XLYHV6mFKccq9+G75GGRVs9l0oVY1I35Z2d3i9HXICxZ
T1bM/NCB9D1LqF9qqdrns99yigMl1M+xCXQhoY6Bhibx7ccnVPJwmwQZVxI/cln4KhUxBXHMHwUJ
gI23WibOBLDfxy6VY7GWckLaAMv/BQp5YG8VDSn1JjfnravJ09wtCK6oIplFz5TIkChB/1BGBLIU
5KoAtCx5GrHG7yzIya+KjQ+ASW+BuCvGb8RveVE6eju4ePx6Hv+9ylqvsFuCN6NB5B4ma+UtULNC
kI4ZB7gN7YOzr0nYl5ihMqo/x/uwQSMrfPGFBOYkR1lTdCxpr1AFJICt8sUgaNa0oIHxmc0BhkpS
otTYbJNwkcVoQ+Q0ioMs70zryj7KOwZDsz3k8BCJwnRCRijbGtWazn5BSeikhFQAv6BETHdbvJUz
/g9rLNSECo9Xu+cPyTP4CnbK1x54uSfeS48MBTsKA8gu/blUO6Ysnp/Iw+VBlLs/w8SQZmzd/nIo
7qSFVOCe+cZNT5qWeq3hgTmbAFSQCiBNd579aYWR3t1HF0exh6CS3Kbwa1TnWbtTAaeQmcDSzEt1
rzwLkaTHxORKRD6zqVxQecYb992Lsl1uT6BSDjoPYYJjfijpcJKAmC9x0KYX2F3yi7zOFfs59048
L8Hoxf4BVYRH235K5JGO23ngot3rM0QIC4ES5rxr0simhASQzH+VZ4JuqfuPbNkUxd5ZW74M+SDp
xcGihPPkVPv8tpIfY3g1YEPUpuvkG6KBfnk5ppV7TnNagF0FYDn8Cazm8z9ZnDdEatG87E36gYXe
y/43uMXw+pb60FQxiu1RS7VYH5AbMz7ON2n84t4gF+tOORJtSDp3O35vCjgf4fdMbWNsMClzwCkK
oDwKcQ+h9lT+C/hfLVmzizJWUG3vwcEXauIMNQGmKEA5SF7PMHRpaCSEkTh7RPuV2O+yGKkC5ESo
DF/CTkVUJo5e6+lsohA8Ln3JcfIntV4XNTAWuU+Y06eJYRt5juf11Cl+aBXp8hgM4b/QIScASV+Z
pRScKO6RIZHubS9QeUoIRWy0YwIb6kjSvIZ6Cn02JSyIcqvdtZpxwYknR7d2depr70oL/+6K1hbL
R7uC8SFP0CcXeylLQmlFaPxuzcCU6rahXHeX1uAHnXufxFxTiYbwQyiAajXvmwbVJU0EmSd8l1qI
DlvdfeYwU2qH7JB+WRJpGghWycUtRAum42zCJ+K/BV87kapP+krGvD2TFLkaxYNbawrLxyKOmoPq
qdP8diIiD+F41kW7KpNU3QHWMDvfPTsPcCqh9tx6ONxq5vqsdKQ30cJkmKKeI2Jw4VSBDR1ScR7c
Nm5N+UJf8VM1So6tcOYGQBmrYb2ijM3HroAmFUMfU61PYA3jum9P/b7SN2WY73rzPbP+KCDism6p
AdgZb3mDkUpaZva4miw6eifZzZ1ThVlI5Xboi7gjiVYZwJUD0iXrjqfHs+RvIQ3DiHFGjzaFfQjz
1MBbXfXpXdoKj2k2Falg/jdGqSArIOuH/FK1Pw0QXUULhzgXr+ZFCP8TGrEuxhk5yADjOwr7Vp8V
FZt9exslwO7/DejWcsp9UH+NFYmeEbwXzRcbaSORZ1EEOTLwDUf7V4hITzdAtdTmmaYyOL99EO7j
IrTFt42FXxRy2l66rYVmYrnfpiLNtzp5m6JUT55c0uNdjbE4wIjsdunI94QbvHklIY3F3FEdq+KL
y9/7f4UDwXO8OlIk7iZc6PBtm1HwSB3Gz8saSY3EFcxvE+Y8hqsScXCak1HxfEUC0fPfOThKWyA1
yZuUY3eMCv3aq9uflhs/epBUmmnU8iUUcEA/AIJwYrUv7WjWik7qhecA2UbjX+tHjV5/2ARzNsA+
fvanLPdgrdaIGSxOWhHgtNzoQCfM5rmFDmc0tfucK79No+n2xgC4/JuC8y4gDSJzeEQ7wsjdmRLq
Jh1qXCVeVhBnBjssvdFBeJSEe7ZvUFfULhdpdRWXJRblmOyzYDTD8n/7YgIP55gIwwJV5/b9+LiM
sKj1FMqHIbxdkilzv8L9onVciNtzDK1LCmaa1DqjUI5MCvA/klosjMbot/axB463xBBqsimYH5Lf
KaiYz4FDXa3dmTLBbfEMUSBMXxZeWKWpSX8Mr/ZzQwXWmShpTte5A2Yu5+0oTpKmd/KLx9lDnvw4
GBg8/P2dWUQGpvu5SoCu23OX+7qpe51c7+7XLALF0fGVA1txPIkmb97iBXrxuDsVEuEIHBmLTmCr
VFDEnGyfXS+48PRRix1yQoQgKQ2taBtTZ4ui76LRkFFP+bbdzkly1d4CUKfZPsEpKQYcHXLHZDnq
sAv6yMQ4YqpB7PUnUvwj7gbdQDMdcRv0Mo7nt/d6RBg9y3rgKSg7CoYql6xG5o8jiLUTE+yr6HUi
FsAZZqv+KKJj6S+O+Gp4lA9jPlChF2WoJ13PpczieWhm1yspWSBGe4LGA2sL6XITeajRuhrKq/xu
26I9SyCimOAX1Wi0gtw/UYwVas0HlcRkiY1QCe0/R1z0gFUBr7PR0UYzSIjTib4Mfah5f6GKYjHO
965+q08ujT8tbScS50LlR29Dx3eGEThdj7cRHj4reu6vcG7rijPRsxIl4984V5m4Oj4sf9umLfDD
xj4nVw47xPD4H0z0NbE47U+tYRo9v69+JlesBgNl/znW0plh++oOOVpzXlRQUt4cnxdXi0BF0smT
/U+84TiPWy6VJpmao2vz6zLUBUQSYpU8Y573IpGHnQ8tlh8DT7ohIXVWCpIqG/u66eVBmfwat2nt
IejXWDIR5PWz0M4VcqFcOL/0X+wnCbE1t/ikslSpVMXxAjGFC5so1JnPo0NhGAPvWV48Fcd/DuvE
yzaoeSn4DRJq/L7T0PxxnD8WU/Z6/7JbqLG1avYQ+CmBKRuIROQdezl0AbYZ5rna/u1HWuvZ38ag
F9nuxyNF8NyHQb0dbYM4DlEXO4ny24Z7PEbSUqHAYjQpbefcTl4vvHsVsjyoOoTR+GBVQDM+NUSb
wJNMluhjR1fTIKDYW+rBBW0uOVqLU6oZsJYcU29X5x9+l2Kv0SIqzSOjfsiAXmewu95OwOAt2rLt
jjfIDaPHhhJTuTYFalhhgW8DJ6ohvwPE2ZCmQJOrobQMt/YEpaEySjr//Pg2BeCAFQ+SCnRLlWci
9Am8jf6IEvVb9i553Kv2yvQnM+SeZ1wtFgjboBMi58FnyGyOo4NREZNE7B4ilKbPnWOkRHwyo4PL
Y2Q76gYIJK18JLdko3NIuH0AkPLX4fIPfCBXPJ/3tJFG1jeV3jB81LD/hsVy22KQSXvdNegjztMI
AyNk6IaewK4BVOxk69A3IFWZJkRbGMVj2dpHnXqc1LDW6X9OAhBMGWdk19BkHOv8+EgSlims3yr9
qT45XPwDUQprx23zyEq5EBdH3qRC8j3K+CzPTFiGCxgWEwueIu7dOBNwkWsDRnVssikZNCsoeeh2
Z7ZgCRm9h+EKiH2H3N+ygID7G4MGXZD+4ABw6mzijfvEOsUjAb6n15/zQXIaXEf3yeYrhu33eeXW
24R5cStLNrre9VgkjZi7OQHwUEVVGbuLgvIlgxOAKpeODIKycdspnLJWH2Bs//6KJIDAzMnK+o3Z
w2NKHmFx+9T+cknrf98GwRtKbJ9bKYYOtbzzwtD/PrdK+aQkTwqTKReekQvFVzyYC4HwDx4jb/Eo
a2o9qJQo8bPv1wqTKRCzKyKx67MksHc2U7Ds+U3hzZjmSYliauC3bJAA3/AaVeXBA3TMbVHn4w5d
mvOVcYxd3QrK84YDCZI3JaLW6cwWRHPR98vj8hXfL/OKX3mVpJlh5KXyUNePItr6nUX4RVxDBDdn
fndqpXFq0HkQsrx12YTxHDS4YaMC7MzqqEgAMr7EOUwDeVD5ai9c3A2qk38NI159JGHz0wn9d1cv
FvCy5ykqoRrCr9B7YnEOERoQh/3Lt3QAyLtOhUHYqsZ1AVvP/UjmxCg3PZg1SjAvraJvCjiZtHa0
NTen8Kakeh2vuzeH7wgwzNFNWlB86WD8MClC/LkDEPMoqCIS9iq+PUHo5GkCJXa6D9Tg/9tBj6AS
n5znhgBsP1dDI6zT5XzYidxXxXTtBbv8XdPJgkQUu4YQyKoNirwPFHsMozT9cAcmaJHrvz2VGGUO
mq7PHC8X+rxtyyM3vYV7EjEFzCHnAfVXJPYcBjPX7uJfPMFUg1skXfz04mj0B+LFMMcxlk5MPfkJ
pZXfo+cOQ1pZyXom7sxscnXFhrIW6EplHiDXQW+9fEtrxkNhAklwkTKdCQwiwA0N0/C8vUy/wpIx
LDY7Gq1zHjq9zhviWNowOIgEw0wAbJP3pY1I72dla/CZPGoGPghR540kOyx5YrsKeJBz4kd1k8/j
bUvOmL3TE0GDlsMzHVvoAWpNH7sozYpaimaDS5OXXefUAyRRzehdazuQ0I2A64k86L+Pnp+bcWQl
TyWjCHA772qxLjPiNR2Fu++ZkE5unrYjUiHXt6DLJWyWOnah/0MoUUvGU63JvtjURDwVbe2vP/GX
WF6DjdLy0VpO7tjgDR7MUrN2v4/zyU3lwszP37q+E5hMJmZjGn4nywnXQUtJPevwKmO/kl8hu1Dn
TMg+qym1NxaSCJxe9kXeUHkj1hQpsg3xjXPAJuTD7E9HJwx6XLhOMKEqW71xQoBkiWpPRzN0JMsf
XEFdxR4eI2R87XyQL72QqbXdVSNHDZKFaWUWF951sZ46mxhBWz+BgCEzOZV3YeTQksQY+qhFRXaR
tMz1I0xOu8i4UWGP6tb0SkBfhBpqGmP/UHNT+XeTNlyyoH2MHpHfxZi4ias95b2gbH3+oAUU89jA
BEIRSNlf4p4weYQ43LyNComefIAG/S2jsyjgVNQ+/utVAGNXtQjsyR5NGB+6ALRGY8djolMiKFoW
T8KbzSP6TGjaR3T4SgGgoFVk3DcZ3vlF0bcxmS9VFSXINnrl9vyYL8Zj14JKghqea2Z5bM9d/1X1
wiP5qb2PjrxGhyAAA8YrbtIxVyCT1QnuIj4qGgIZkRDwr68wy7FCNTM1R4LQ05GE60pPY7HsXtCV
gyr4Of5bvSx3Tz8MtEMaLWGiUf3H2wo0bJXjttc54dNARXjwt0izxfN7t6UeB3kRDnqVQ1mbjtjw
3q1Dz5ikQoYvEOJC/B3ibgnNymAPit1hR/5bzLDk0vmF6bQEWx1dDaICsFJsHZI6TZC4cUV47Kvu
qS9NaWsYRv1joB8xjCftXgk4i53uH58Ezez9HQLNda2hDNBodBAM0MCOIURDCr5mKa+Tv0d6uSDF
u1hQ0BJBGz2cZUUoG/vRExURaqZzHUc4pEPR9HRHLcvCWg7gGXkI+Knyu7jMsVRqC1on32KyL0el
zm+6d42p+QPyvKjZNEnMmcK5ARgnpDOFw5wQx8PqoDZqqfL/7N6ZMdBkJXlpw2C2hQc+5emYiCoX
zWY3nRxdCRMQO4s3e248a5tcbZwOitHFdCjey06NvsfdWGgAbEMMfAo2xwNDMLrJ0vNifzfznzwA
fSOzabiKgBPnhM2FDJo7wubeUZBwSGqaS53EeMB7Nr0YJE0GQV2xursKikBqmnTHTV1U/NvE57Q3
bn3OhZaGf89tZH6NWRWLeseHXiePPV3UubQ9Tx4q+6sicy+zHJzfARxnNxPlbaolomDUpWAGqAV6
JbqAmdFpBGqYznksi4KSHjJzGsx8ihRn0C9ouZiY8LQXlH4t3zROTsUsuKJLfSiE1RrdJuAcUVco
5KnYnYGd3NnNUTb5epDKA3tWVc0uxC+iiNzlb7eyjPi5NUlaBhQI7aAMLOLpE2HR13F43iLG0kvX
JeBJXFVLGoMlYLEwrXc925+4YzW+iRoin5VEBDsSszLfBvZFN6T6+TwVE5HfFAUk1x5JXypeH1s6
Q0TR2Dz3L5tc2FHoyPfovwnUAYYA4O3CuDcVJ5gGae6PVruSVd/DW4Bh5G7GxZvWraFd9m7Exbn7
UOsxM32MSnPxYaqDQ/Cj39PMNOFdELm5quNXLzSo0wiWrT9KLMh3hc+Bww5fNuhGk+6V6jbNnpRF
+pEa+y/AbuKED/61UtRFcsLTqZGblnOyO7E4UZPCXLhKkxGs2rSVTMTebxcaK6lf4rRsENId1IKU
Pwc3JxUZ3iJR3DgumYnLRWvf6jF8MxF9SGRDfUz2gdRNW8b/jaEc2t8ZQFcsQTkxPf4RUgqlVShB
NBi8Efo8fbZLWZ+qaqcZeRxV9C4Z7cDMpsWeSY3Vbw5JbsqKQr+OAAr73bzPE0VUcrnqKALP+shW
t2fwjvqHd+gVfi9HvsyS/jFVoFL1UcnWWJJPo0pNCJaDif60NVGrGpEOrRAoUFXuZtJk7UiTtcMS
ph/6tzyozaUtksliNdFg9Lwhsl6JJL+EsFdfKw7JOQE6lIX66R7kS00es/SeZj/lB5hWK0r5RoNG
i2Q2DH9gtc+PY9ke9Mk+9rXkNiDJ7AZfFUYcIPu0uXLGE32fZK/LvJGsipv6v+u3rj/PXEmzX5+d
P/erm7pFTdonLHmnBAU/9/I7Lm2vW5IlaD3KPaExLhUbRIDuAxjyPaAF1T7wrJuzEDKThmqWoOdj
tzIlFmM0nDVNvgcngWMNyLEOgHA93PHJZsNHbYxBWUYPaSD2coYk+OpNar7D1KRUO8+EzQpGWlxJ
bzPYMAmuiQjJJbtTbp5v0kzpxVXK/U9Ek9xqzrgWWzR2y26rGir6F0XHl8wAwjdW1uNWaU4yQASG
HhcWw4N3Mr2iJbJ7C8LeodIxZii7P6RnEpsJhs93WL4Da0ljbrtPt2mWgopYVHYMrkXR7KLZ+HkC
FJ7ntmJEp6ssWuQB8hkhN9NK7CVvAFZq3uG36paqwl5/Hzxq2z97VVNOrTfmBBmHhrUeatjJaiPZ
oVJCey6Fg/w/hotvGGxWvLS7VheiRTZ0YeFZWoKNO+NE4kdkjjq2kaLya9JOeUrfbPhnp30AwXJo
/KhlsvWJ5zWpab9te21j2761ApyiPK9F3CRLfjVCvsd7EWbYz6K4mYnv453CneeXgsNw1IzWBymD
o5ehiHXceDVdA0KXice+pyfFScyBPwgPoO0npg0QhS5X13YoDvVHxZ+xkPC9DSlIJ1nKu48sAPDn
ZZ5pNexu2Q8wwicCuwDfe+uelyO+WxR5vbGrwg8RXSywpz1/A1O9XjAO2Yupt2LzXBiz3ER0XcV9
d7N3qzXnouzbeHkHXS6LaLFm4vkpLhdgnq6Y9hocQYMFltBw4xALJRS2CZ1IGzYE2H3hCp3Cuypw
IkFBdvn3B/G/ElWQEe/BKQpqdOD0aN9YkCp+tsLhmw1WaQDxoO8GedXa7IN42Kp7mQUunbQJ8/N5
JFBQRuxyCqsVYc6rineYlR6g+Sh1aXn6fu7rILp2I6rSGx/lSzp69Gv8ZpeMOSJCrnTgDZpk1MbJ
tBjEVXXnNy7twRcSaigp6JYo2kVm4dQ2fG15DjC+1ORMWCikG7D4SBHw06MUTnAtoOQs/Ll9B/eW
xO3AYEyZ2mj1yVoPp9jvmCsr1t2Zl/YWYzlxoGhw4nYt6xbAgFpHQ7cqx0l9b7DoTmbX63UI3lRY
f5xM+13vF/svkaFRQKQlw/ahFmMDZQyJVUShil2bJFYCQ5YsZX0/B1JTlyZP+IE+2S5zWQ43up38
8M2Ntf/z/kZZdmswAp3cvJfYha0+DE1L5zxdhrWAj/zpukMmZp31EdltGr6OLvx8a8SkphGD7yJK
2ZYMOaP2pInVwMuB4jYLhxB9C8dRBapxEE8ylUpOLXHc2458IFfse6FOzdd+8L67YOQWPIhgPq6u
8oGKp837IfBZ5UGsyq09Q1OdMNOuAcLuX5R8zSUfSqzlHSuE7TaYv0YFSXHY+toQeibPFZ0bhja2
ZV94/bRpGttDj2/wdVmIZRJa4BGEwjgHalhWbEyz8b8mL2/OgUKc0RVVIvrGAJ9O6jIrCJmQm09V
raiQZcUcLrlmkRbScizj4SMKe/m89kuo/LgarzQZXWGStmuEy7KcXfWyo2Rqs/qFdrb8Tjddu8qK
yoKbCrpau5ioCLW2aRJcc/js8wbuGVBb4gqbdvR028KZ9uZWgt5pmaCz14yr1QFcfsgws5TTM5LY
bUgahT5IfWd8TQZ/QvBRP4bCIEj4QBBBHKAqUZtlG8uIPGHvkGDJDPtoWo3lW5Q0BZThzlRi0+VM
VmlevH54+js6vZL6BX9X/O1oBfoDqn6+vLK+aFsvfLk2+x6bhYmg0TU2Xbj2f/1EZkfy5ekpHJ6x
AYKZh2+VNRZGz9ITrtz1pfRFTxfp6UYmWaP16Bawjhfrio5UkNmt2zMd84Pzp4AIrN9BIu0avIqB
hluPGsjes8CdH10JocH+XolD12xKAgByxrUN6DHKXc72Lf6ZoJof0Ttm7Q5L4hNmFkkFzNHvRPYK
6BW9dl0dZHZDzcPFMSpL5F/2sfZeOQa7ks71DfoJCjUhoTdfo9hPYHzLmUG2oldqVx3ocEnIONdt
Z/HiJz8WjXX3HPNuFU92IEq1oR3abscEIWqgDt6fWg/2vNwD2SNZaR1M15z4xxBktqKfwDyi1nl/
729Nkeu/+xJEOWAfG6+LxVWR+E4ufTbOZcFnhpWVmvrbnNM72TLGXaVYsO1Oq7qTOsSWdG1eNJu1
0yzyXcjUrSBtjrmGVl9Hk8KEmQZw6TUN7CNXLycFEwNX3g6YexHxaI+poy6Vl8hvhCNtOQE4fGlG
deHKFRz3EfquqyFXloFimmMha/1EV+TGALCj/7io+P8sDu4z+kHCPF8K4vdVSTrI46/3Q7m+WMWb
SyKj5hz0Dy6qHUxtHXRzC09ER/71c2sT+tSsoDfMWeYFwKItRwEX+lBe12/Sr26+SqXzeG0h239p
vMQVW4DaTDAVSuXhwo1pCxgQOWa0osLxsGMFWN+/nvOSs+kcTzvsk+DJn6aih5KG1k9gFSS6AqBO
yI2NaQFClqdtBSLHIja34oqb6QVOrdsY4yVDlSuh+RTP5CfmKMDB98xYz0Q9dOsE3iqnOUaWb+qs
STT7j74mUwZQqKs1kBbuXH/GgFe+wFBh54Td9ABNYiHO06XMrjwPNo1WA17MveST2vm02ApnCSkE
l1eijneBuVp0i0ohTfZOXgtIoHoip3kfpxGuab5bqB3ZA10kxqiZ3wFFCsCfZxsGunjcaPgGtVzj
G7PGozVD4Jhlbzz8wR9HOiwFA3jAwVonWseUWgEAaaaFwh7pHE12AADAxchDkVt4OYIF6sAG6zha
9Kj/YJHlWUebNyOnoVVkma2aFQc6zk0ke/7yLYk9Qe/hiE2Cso9D5Uddcw8y/MjEdNql827DeyXm
lYQ8H057hkMOtLPkyeKw2hfr/yji2sGw6XOTyk2DhSBEIn6aD1VzmFOWaVn+eE710z0B3zs8u0pU
KJIiec99IcSuosS7hOW3xg577Ei+s35YEYq8Uypis1aI5iS1DMLuWhNuacCIVm50+nH637VTYj54
QAF7a85PoZp7VYz2LwLJXgMbczgTe4sFGrlCJZunjHKWt5CRINGkkeka2U/xGgflgBlcjVpIJ5rv
dmlSg3qKg4p4QmqN/MjQKE5U6duoOXznSayGfzYwP7BzCRRZaHyXO9AWpl6G9QuLOPojq0wCdXBH
jK1+6IlyXx2+900wu7C036iFJHmKPL0rUTqC662oEBEjnX1ebILp3+yIZN0sjPs6rz56pYNDx5W7
5ueohYWJMgJM6xm0BOnzOEHsofyUtlGcfE3Q0LomAwIUmm6j2kVnPkkr0k7V285ArqxArRkbBiv/
iVCR1eoXOTwg4Iv4x9o7RP5ER7YlPC+IVXCZAWEu7768UKmAOupNoqeKAHl2LYK0rcZKZLHkILKZ
a4YFQFE9AKu312Y6UCE6QdZcgzEPLzgtCZ3iDuLxOmzYBFcFNkGAEcfoRBLYRDagKnxQjgDWxTd6
0I7wZPQ95J66npIMV63guw1D3+Xtl3yjatF8AvghI+8vBepAZYo7fa4MsOTgw7cKp2c25LPNWCMX
ihfjGA3FTksQSzqXL3Q4FVYfmX3qgkHR9ewKxiVIOO5jciRQsK1a4W7wmvjnALE6dwVNeMHZRnBN
XZHhXeUqo1isaFL+aHCIPiKdzi719vQKhMQAwSE5aUXWPfVtdN7NBsOlj3NNynqE4IlOkIwec+Cj
AdK4LDku29G/ifjClCldCn/m3REGe1XKYgueBf1C1WXNALVtrVXlhVFZKk0PsyGLqkemc3ZEkO0L
lYu3iJ3lMthedabqizi1Tg8uslxrZGRwT+z8jAed0NtQXni9dPmY7r9hmLOBkE2g5MY1heEKfxs2
NauS2TDX5VZ7d3azZgtA7uUmjsVceEbW5Vn+DfGccjFprPQh+BMh2oSiQWWudC6U6nlg7rEg05aV
4iYoyHkMMSKK4rzm/sIW5yVfBAM/I1fYh8yHJk4DGvl+eJhhoxGzBY/u1mgFGiEqlWTQgh18qg13
GjQctRUKZNQN9q36Z9pjQIiZRaomk57FAZJVNJbI2G2H/YcA8Pfc0Vut9NWWLY4kv8kmlxqz88RS
bGsuHqBJs2SpFZTesYJAyGhyAUb92b37MAByzsZUPzYdgdYVC7uxkgg2xIuQt59TTtmjB0t0xk0J
2xi2czMgJkljDL5w/JKGqoeSMHm4UjBSnL18OOi8iyS8EV/o0McwUzuo4HUV865y5QCFpNylRBSm
q/yCntqIzpP2LUFyENbW7EFAF3sK7imR6cxBjp/thkSPyYDUVbhPXpRIexheqv0p1CAHsEnlFBZP
XQMd4rvEChKUxT+CMooc++xqVV5UV9wAIvcnyKrN61QilVXOKHvZDTT2JC+NuRWQr9kplo8v89/8
qWrg/SFOz+M10v9Da6sLik//2Z8sCh/P+yK7oxTWnhpaPiqreS8Ul32szI82DOE8eAZTkFPcYTNS
uoDZP45Q7m4Y+DLvk5DkWta2CgMrin0bvnK3+OteWEwd17ycJFDStK8cv1OjkqVHZE6dVYCJogNm
22wY8nTD0M/BcgskbUsoy3rMEPLZhwQhJyeJMHQVHAGOaok1oEpKMIOl/YAeELiHDPttumAseqc3
w9lGwm4UhsPCeXLTw6e9a1+j35cGphd7zB4z8/SYK8JyZ+bB/yH5ckx1sY5ucAi/Xt2yHDINoQgc
vKFFXv/OCsZctU6PBT5Q/vbDciAsZvIUNKITyqB4HhGePlmprJ3NNuhVjDXeVQKlUOjq2ubJ1nAn
ieE2MlWj4sbVKD1ToaWv+uIU1YCxZ7sT+Sw0nUTpS+TtvfzbeIqlDuyzvP1E1EShbPMcegVobeg1
CK6WWPrM0RbyCn2IN0eYTOLhco2RxqJ+Tu0ota48jhh5Gc4QpuvisLpSYebm9Ska0eJMDva9A8lC
eTI935Pg5xSu6aQQv9CZYalIfBkiFqLaczQAHNUYFtmzOZ6MI0iWclGsVL4ojP69gKVdQTA+Ls0N
3mjgv7ms66AaSCLTRzwJ3nltRuGxp1DS2e4E2F6nhABKkzqZK1K1gOny8qq5/CToNFOlnMpcb6ln
QPzb00sJNgXv/sR0InrXEM9qF8NeDdsPDzWjiYxP4oQMMrW7F0c+DNoWsJE5+Wb4T4tB0A66SKLv
erAiMB/W1dnZblx9LDTdF4Jn0WaZsQTg17fUX09zlj68XEZlpoAUQtvUoWCylzqXyMwpYzRiuv/N
dvI7q8fBhZ4V9nwaQJFIa9/fgWIcWRA0BiYnz3MaVI42c2X9mCoz5QZ/hhQolfuUjmZNoOCyYWQ+
KaKZNs1SlYYdapDzU4DNMOm10XmdZQBwwT2ztFN/61yVxjtdHUBK0MV/WAmIfigP18UVEcxgmvp8
U50q+QvOamAvqgLgDIAY5/p42zpcRTf41i3VfU3WmwYRlrjy9veTM8zxKfH67XiexCRj2RbIjVnY
NPD1fCWaykVsG8OuAoLicIzVBrUrS4geAxJK5KpSAHkuj+LrbM3hYk2ZL6NIyDVd8HCc+3djr/s9
dRJog/7PlYFZ4ykWHpl7mzEC17GzgxV529a3UeUOK0h7f7/zwGA8cA7S7SnJgNPDrglLjnRIH/dV
EtNWvL7oLNagorXI0a8k6w50Vgrx8Zrv6K2xM+cHKwqqmTxw0NRgebld8T6mGxA2HXS/9kcDaOIL
W65RkJOp/qh+9YUkipZ1xhBOwGxSPAJDy+AboNUg4QQ+AuYbYcd7nwkSnp/wguVhEWBHHobLBg2Z
J8EpUpQBV7+Ji3hRYnpA8MgEvPzp2x9UaAI/VCQpULu+6pSHuzMXVHeO51UTHDWYvNrLWe8vcq6E
o3lx8O4BVJ6z6Zb/dQpFr30YmcL3IZgojAwLd0J2SO/iMYQ9RqDyGfqqB3CCOg98zvyrkASGWeBb
G04+yJdmdoifBkyPatT47cOOS11oExu6E4wGWq/Oy64k6BZOrbgtNcRHQjJJpBA9IdRGHRmy+c//
PfGPNbU8OXcYK9NDZTc1fs2d170EGiA46YBjhYAqE8w+dN7Bwt9IpYylIgRx3M+Rivd0Xgfpvhsy
jfT5QmB7gUAtDDjFCQNm9A2C2t3VyRL1Mn2UeI7Nk+qQq7MUCDbZm1Wkzi4JWDeHJjpsg46kRGMT
hcuUkgeIsjzqbysvu9yqhbqs3xnmFuF9rduu1KuP4VIH4Fn6pUDbQBAC2+Hvo9e3pja8Pn5owlKu
6iBuzUBjC7jwIz2GbQCahVK/Nswq/ME7h1D27WfofYVUiPwkDkcIAHoEcUOnrFtuUEoXaLRC5vB5
cMhButcOI2PDKxYBwfOPFN2uleBWST1EKi8boQmqF0uovo/SX8hxGoSRsW+KQ9FTr+wQFWulV+xl
BjKnTlcXKwfF5sB4DIrP5+YVLJV/4Ez9Bu4RSJeitUO7X2E7C2Cm8Ztnt8x9uEj61HxeY/GylvBE
Hr6LpqI8Gj67vtdy6xtnywvtuKoWSz+x61+fyJSEZIq8Iwn/aAM5c12JpG6JuiXJ8wG5l7bho5Bo
AglqUGxrrDVD5bkcd+eY1pJ6nAl5rWBoD/v/cKFFeTDc744W2mOsb16MG7TQO2oyUCvYTT3kdGzi
hoxR5Z5T7cUgLfXQm7yubz7mGgl8V5GlaMUKs6E15Bn9DF1Gkw47intZrJV8qcdmv96ptQk6sh/q
veWzTuPBYdcb3+Awl8twViBXvvfuGv4/IHbN6wemDLZd4uE4n7fpmzNUyk+s7aKpRo30SJSx93N9
1J2AtbKkknm+Lf4kEWIpDPB7NmPJoVxHFwi7It95qi150MoCDZFeubBJgGnfg1x+rbklG7zo4h0f
QhDbpLFrfTOW1RVbH5nFYeYYI9ZYZzahEi2WyyleEupaznmHmoQ5P+U0JVz2lpY8aRC5flW6PRbm
XN8AG5MEsgZ8YBLFycoDPs88J8r7NRSkVt/G75ezz8VEuw67q6a7eBk2Y+tzBdFPQXzJVoNNfJaW
ultJM9/sExx0t2GlM3w8OPihnMlWXBiRfOQdYSvDZaWN+3+LKCQE0VO8l0qAQhII9hiYwWFTvYCQ
FTh8HfnA8P401mLeajO8bEeEV7Jn6dOiFuSL61XkifhmqQt7gKcPm22piNNzkIfOUlTo9jCuowB4
8Gx0d8e0CzFMZOy+n17HoKPFUepGBjexAIgWus3MAzdyx+MorSL8UC/0Va9tJCZz7TbEsrycAcic
WJ18/UbRgumUWXlWUI9am2rJQ9a3P3uRTCIIoMBbRL8pYSBIy3d3O2uyYzD9zZWORYHPgfP4RrsK
tlI5s6qFOLKWpH64LgiMkIzMF+AO7ENlMz9E2tjd4TVNzipCOdqAG2R4QUryQKcg8B3T6fDO0hP3
8u2+TJZCVeA9PPHMLgMzmPllsAl5qdOSZVza2RABzOEsFbkp7Qe23X7Qcx2S9K7wt1MgrMDSLCv6
28oBwL3yvd1vwmSoYBv7+BUaTf50NyHfKcbbUEu4BsHeFBe5HopPC1/N6eqHt/vahbVJlKoWM+Dw
wvc+0mAXwwHsQZeCuR+7mXpj5JnjQmJTdCEFPbW+1MP6ckVdNTVQOzG7Z1A4yrhIO8a71PLTUx5W
xKLSW9ySoCw00dBlUkxWGYzoFdb504MzF/kl19NdWkgVVs3mESXkfX5W/ZodzjxfvSKeFl8aDXuE
9fz+oLI7x3zHEwm/ka/pPYs2PB2QeMoIRJp5yEOSz/ot4JjSAOlmvjlCNel6jy8sndb2YoEWj8Sq
mhiVjMM554JAFsF1UvgKHdUL1Rh9QSQyYWM05ct3jq4mrcVU5o69fa5HwX8tFNS81QPMmzSY9ylA
wH2YSqv5g8SqMR5oiUN64Ggk/LjnEiUHbJ13Z6uvlSvJXf6goINIbO4haLuVL8SHsWSv63U/v0Ot
GBsOenYC7TwlckqCH9XsKbxL59Dd9XSIa/q6+RFKP3JAMAWQHnL6bMjRpLRurU795cdFtqEkLqtq
BuMG4jhBrhjJEtLzcDUgzu7feHWWdlxho3Ql2wfPl16+bHE/w7c1j/VF9s6PzkYRgxT7pAVcOOfu
CYJK7vZwsOzSaZfoP9h56jK28VYxHTmoePWr1WVS1YAhSyZgiMu6sYYn8yAiXVh6XQFGufdK/C9h
YkjsrPrd6HQUmuszSLz4NLZp9mgE1SzPaT8P/1Cjoq8vqd6dWVZraReWzaqK4i6xEGF8f79GVyjH
2iM3/m+d/m3VBJey86ICzaZm9bzWpwaTqo5j2jmsPw+hcLHpCVlW6vIat3Am8VSVRlUEM956J6bN
AGgwj24qvYK6eKQpA04MAoMzoysqxfHO7glI3LWgLXni/azdTlRlYrLNSmfvteFDoFTLV9+UO1sR
rAVX/cWiyeWP1ZP2GhfVdon7Ox065pEm+Rvh6Klyntu20f9ERrzF7zI7f6ELu4FCnK1/jb3W6mji
q+YEht9fG7IiW/PrNtPyddWiS68DmkKH/L1VC2gYKokgWubpjXwdQv6g1XpP33Tzh3RA2hfYystR
JqWQjjc8kYhTGF7JPI80fxFS3kP3f4HdTF9JA0ySL5409R5qau6FMlqz3zcojXze5g4gSXuJledB
mG8SoelwihIHFVncOABEtu09uuCII32ZAuBRYSuEHsdLgxd1iAaHxgZGJ1UbXeJrHW/Zyvm9ISl9
lXcWK+BZ/ZwGsF7ZFjOc04fZQc87ClwtPgNVq5KlAy2Fw0P0kmQeqW6FRLehmBmmk2JY2v/QkN/9
pk0xf/8jMMBg1zcP6cORsqMiJKsz26LQFEiLpyQB4kNqMtLUhrWE6NaYT5MksV4LS9zCFFOu+nKG
WkCqA+apeF4KSyY+orh/vGBfNAB+TlzLKd1Q/5r/56xRF4FKwKp84wdC1hg94H4vR+B+lmPtsABS
SNubEHXvhxxPd3Z7GmJ2qiby+Hy66uxUq9eEd0Uz1+hfspHnLUGp9mj1bZk/4CA79IjxFKuYwAB+
BNkqBmVLK0TTGY1/mRRQq1bdd9o0HMn4czwjnnZyUreSadKbvOSPNsXct0E0Mdh56N60ZmPdE9mm
PlrjkoTVqyddNFnp2ezsPPw/MclveY8l0b9P7PayvFDvFAyXR4xhG4UA4lX1c4S9tP2ZXmHLP4KI
pFzDBzy0tRIF6+PlQGqqTZ2961ENRHz9EtjEVH6do2j8xbnamb1D8lyXOut0XtXq/jxgdkA6R9Kv
AVMWCqgfMiW/C/4VjNiFV/Vo5XhEjDFspTDAV2rYCzhnzNO3OnJ9FezvGuMBTbXt7Mlt8PKuAvd0
bovjaPOR4Iem227jUo01QEORCXDYO348/+UvSq6B0aRxo3eM0mcdVtZpuV84GSVwPRobDfBuI+nd
bmCpJH04qgYamwbg2S+nPKwgctW2+fDIxI/4dNmVQ7WjcXmFVw9lq8Sbs4O7IBdXNmILZi4dhzA3
xa46vAMLhvlp7+mCmnAHcwBH+P0392I5/+VEPVh1idtYIw+6haCxpJJuq2e3AwhJbeMkDS9de0dz
5OlbqgTIOx+IEj83cVgORfdpv0Wfri+6tsjrM7Xu7XZ4DSm3gFmff2Z7bUVxGOwvs9X/PRpr492S
L2deuOmH8fRLp+S+01emi7fi7sBe+yTyFhgqPmOOH3VZB4FpQWxq9ulw9YxIeGWHB6RKNULMcaRV
kGhX3jyVhc7g/5PrC0bmTTPOjEEIf9xqFDSqVZiqTD1H3c+vr2arEaSBSyGz9V1w9+NG6SdfhpLU
psKT7vk8Qejwo3vAyB17ypfeytr5OQSowGSR63TE1UVxj3vyKzASKxtSqMGzS8Z/BBrbIshhdFUm
ixOuV8hm9ca0ecZ4t2r/EoQQQ3hm4oMluNIe7QtVoHOMZC3PojDA6RjSGPM3LGXcFgjdCEE8lgKg
yGFkIhP93dF19mZsQTuhiLgzoCP5kjpkNfn+ZXM2p1QAddMKzwWqqnBcun8yaMqs/LNgdvRxpoTg
QmUh7AxoKGu0r2KCXjcRtCqBSIo//H0V/PMywoPnYBEoEPCP3+mv1z1A0iqzds7EZOtrFv6jwsgh
AHTHr//6HIuG+obiWlB6NilBtVS0IDQPERqvNMVs/Nr/ENsDHJ6VdZHwZ5iGPMm4ldVyscTUZsOA
u85bGv3wNu3Ll5nfvjlvyqrmq7IY+f2nHfOHDZ5jnOAAwih5fErC2hsvqu+F8H/sqsC1YnATc169
5VbXzazNPLlG6e2lnQo7PQhEmWpahSeSdvB8xU4+1s3BU/u7ltuylkJHJvBXDFyHn2lx1iEfsZ5Y
FnxvRjxMOIYPaMwfJMzG37ofXfn6AfdmApMiiw4hxdRUQPOOrHjAVz5bubJxkZd2auFD7FHRh8B3
2sAuwFH20uuirq+WNbYy2++FPjyfftKlixA3yRuRLqT123c/NZ1jw6AZwabQxREmxotUZXliTTrA
uoSpsvDja6EdfcnAl2Von+TKMKxzWwx5qK94IoxNsjcHxo641Rsdj2Vkl2FdCuLQ07VFWD+sgV1m
YomFaQZUzLo8Ul1Bz23Ux8Xs+V8FHGmwV4PWeoeZF7hN3+iJsQBqm1IPr3bU7+kI9ZUv6x6XO/Nt
uStNA5bg1UkrLm9nQMXhi6xHUo/zB07V2ej2EV4tUczlVtUqhZcIkMeqjVu2ylhiXir9gaRNp4cO
IuGwbrzkfQ5K2htT/8AXXTzhTLDNcSVHLsK05MuPVW9PDiWzsZuxY88M2RcSXM4qxAKo7PJxgcPc
eSZHe4Kzgcx8jGpx0EdW7zBHPfPX2AULRR652CS1x30MnZ5gmojYK5j5tXy5Ttk4Iq4ba6Z+ZGDk
ouEtpuprmhwFx4rCNPZNd9XJ7hU4ZK//TyfIVEONL1jcXy+Oebq4kOkOjx9m7GNiDqoPBLt4UGpP
kXpITTUGLiUYwN9nJiWPu9b2SFE0lczxNpWHU7gzuZQAVysqD76ufMX5m60qc1P8z8JwhIRP9fub
2L0z/Uivmm+6e4mFqJGUoTuCxdcZaaC4k1Jl8RT25mVUfwtph/yk3AXFHvreTKJhAOeZpAY7j57M
E8zB7atdbPWhqn2xhmf/2mBjedXZ86Yf23Xxh5acXykQnfDjPZsynT1GXQ2lzg9sf6ACfRyGBCRd
yfd5ddP0rleU6DqVs2w46Ceom03MoFK0q0taQiuepMUEyVywglMgRFloEB1ojfl8k8GlPoKtD6Ng
yEg7NWuZj4sOBM7amuX4dpJZdqFcwfE67U71GbegCoRcxn2lw704d+Tnspg3WfUqIpddYD5Yb0Ya
BXElMQ3DD0Qe0G3DQT1jawX3fPS9xPzqWr63vFoDy+oB+vWj45cZ37l3OHvohH+E12IZqpjYik5j
XHUoWIhzu82PSkBALjdFTP1zhPz1uD3uXnwctloAGpnag930GQ/G/h6ue9x57WQOKZSNVajbLFxZ
YiELqAopjW0ANPsq3PWCgXt1aadVY4OjRP1gnRtgSATL0efh8TIdJUK2p7okC42NiLvdCeInt907
aGG0BwXdmIQ6JoKePBBuZaLuIkbuDweGpdDyovwMBeWuaCH73+PEr/hmDiKDMLcv/Q52IjZl1eth
K2G/o33llq5Z/tviHWPlHWfUzPikHl5Qcx/KHRW5qRIIGzA/XJoEeEJ2klm20SqXN12vy5E2Na6a
ISLCVog5dZNhItOoTbRkOEf2hyPhltsMaa+hkhVnBdA08GymKO8ItsXZGwgDn6vIlWCdDgiz2l+4
0xV2Puns2Ndwgy0bQxdtlCzsK2VK7ajYpuCVMGFYT14uHe0PZI7roMn8aMK5mwMH7IQGsw1Nzbzq
eFHZdoTgkH7k+eJkno2LaKLNN3JMJSJZT+CNSZFFwxmY1GunxpkuxU6cVVJcst9lRVXC9v3zpi7l
1L8Og2oxClw00vYdLgUaa6DmerWrOsHoVS1YrAeppkuvIEvCqmcsd2bwbxgq1nDMts9cJVPkKnuZ
WspVlhAFtkhpKf969jGpCuMIaI1g4cTLQchVFLG7eASppjsGZOYdlVurphLmxh0vfI0dYr6i5LLl
hF35BDi64UCh+9P+8q4UfqzMdsYjepE8P/zx1LZSAzZ1notd5pq2XMB+CduvRfkkadI3OtB7vgz0
7yWSJ2JNEuGqFgubUWwpMfALE/GZIIoLx2FkPUoucjThoBNPfALJg1hPC1U9Hbp58YVTL3EGL1wi
7IVs1EHdz4YSGg5G1Mb9JsVgjDevLVK/lVR6M3GV4o3/JRmmuetKqkEc4rknykvqVIOhawctXSFg
8Ck4L4nsZ+fvwCtB2zD3n9/yuYSTOeNGcpFDYK4Ls+wy0OpxC94+zf7ird1aji//W7eO6hDM7KwV
0ARWNOS2avaxq8Dx6UaK0xRVlWMAMHTHStpE/3dxvHKgxxmu7kcEAW36IfZjv8nGWBDX/tJlDqOO
0FdrxY0z41xFhQLsl2HIXAnctkN/hgKbeMiEfsojPWOQGazmfFCHh8IYTMDbsbA8OnHucFhLQ8dh
Y7Dc+Z10aq3swO9y6xJ7P5YyT6VWQiguevEMrP9l6ElQGjb40xqGA8LECHaUKIW9uvYR6aM7qpBW
QsGA7OVp0l+cROch0ZJB6P7HpX/xbYxunqFEq4UCCAl0p36Jyrr1UHnqrkzX/CgiiMa9Aq9AI+rp
XminLebLM5yrK6pbIRmfsRHoGuL5LCbsyE4+hKyliW25I8yPfEoWYp7Vw7Oqzjb6QE4Ae2MpXgIR
LVN1IWCHnUeANAYC87o08Fa9cspUMENbGAXFb1k8ZPeHm2GTFFDohuXJn17NPk0y+saW04p/AfCV
v9SZTZstvR6H6tUT6tSzKQnOGKDqDSmvyBnyvalz5dO4ucuCQTUTNgu4QVi9ItLlwSWFFmvWZBuk
8T9oIpqgyY4dpzZkoKZO3HcFmqxexd2UTqwBE+CuoiSOAJbKUhWnLF+voaqRUJUeYYDF9YJnvqxu
u3ZVZhoOJtBxaQ+Mbrp6WIrb+V6ffbFL9LIecDsGicCSP1rKvIQsFnSDqgfZ2L/RwnKlMlWOyZoa
hAL624tS6mMcXxtaFs5qhRvST/SdiTOCDuhPgSUT8AOm+NfHBu7Tcmm44A7x6Ozh1OQXbHiRU6gX
CZUAv0ZNBnifzLNYXT+DtZHDbyiQQrZ9oaV98JeRmSjcMnHu/mWh5aN+zJKTHLCiXpZh4A39r4BK
is5oywUjXD49+UtWq8is9KOIzyZUuvuhXLg5wb6KHPwGgOpqVwUpJHwHowDbJBVauW4jq6cELhZR
r1pej+mr1v2APCG2voFDeRBks9FuaRIWXyCVxnl0Qa4/byw+YMyidX2U+jAPAVLck+obsVG9IEin
N599WI/BXJbVjSdzX/qfTS/KrpyOEPckXALvqi8lgCEWpFdj1MgN4vJtlvVs4k2IPR8TRoxJTnwe
JZqAzb5T5TD3B3ID4xiooWTNF7JgL4rEgwqdSu/v1FTkCIRh4yQqTss7ArirSscpgj+k9nefgad0
8HE5YrKPC9mMhVEzTvvB4Sxs0kXJzI0ovoQrVCNyDZLAAriAJfsJH9mYl6KWWfqT00wcdu9tHovU
GKHr6gOvjzUYNS07/6fqBuRN7Qphige9/2BL2WHK3UlpshIYxavLUF56xQFIYJuT+PpUxUW6dMVO
nv2fR/oyND8FFJZUT+w21KXC6I0QyuY4/y15FnXnHb5EStDS52ZOmQww4ehptV5JH7Zp/DILuR9j
mbHY/2sYyWj6vrNK/hO3zh3n+0NxL+AWqQKh5SZ68j8f1C1cIDdaDDDB8Z473zr1aMqFCFbzsqxV
6wkQxxzKrdRazbfIVc9SMl0HNjJ2p6HgUJcJ9XwWP2HA4T19WgSseVZHRP8p8yAhP9T0SAYthR8X
YN7cVUKMy2pXagA6GqkAz+Hm8O26vTd1TLpdCKpX+8OuJiX4ux7d3KxlkIEY1LxaogBPqwSnjhAp
5H5fRUEQszejhLHK8aIh5SDJ+Vb6rDJRDppSw9Ol8U0JuTHl1t2Lg4NegkW/CSE/S0W2QzGGUk/W
7d6MdpAONkCt3PL+xZww4tRPvwpi9p0G8HTuUHsM8ZVOi99y/MSvPLtU5pdv6cXIV/Ll3uedMazA
B/O+XhHMMHUhFZGDP0OQbl60dtd68UvI+PPrl6MDIsWIAtU4EgJqPTNPxYOpaXm+vsUceO5v5rGt
KzxMzg+vmLI3xSDtBCTd6P7qejJ5xGPvTvFHInOupv4ByxkAS8xmtgn5FohUHm1nttD7A7Mkak/G
LUdO9JG8d7dWgQXanfv3bN2U2XVHmapuesJ4u23EL9r6TCqk7jbhKgMpHT0srByjDTRXCH5GgdzT
UaNlMXllDU3ttY+MZ60fvHKEpMQbKvk0I1EnzPpAI05D6ZbAgbFPDRMkkhYw1rbG+KnVl0I1fLwr
iDyvv8RUHhbs31+h32bh675WUPpmq218yZOwzV1yYOdkrNCAlokR+ZLLbHmx+RTWQPYBi5FvXi8E
d3otb3vqZt1/B2gb3mzEeWBk3RA0osgyWvWgOxdU9SB+SxebyDopvNDaSQN6c3/+5bYfwmOYWClR
6Yf+vE78Z+r0jESCgunKxgoe8GknEChsXiqCNdA2iLCCnohz4IcHQWhz6i8vKV3DEUmDvVWc37Xg
ttnMqdyHB51n5Zs109FqpSKX6GMW2mdZSdiEw3orfu+a1uGrkcO3PDt38etpGq3xLur5AlB7xVaZ
UcM0wW7Wus3bX8BQJunGVS68a5aCXTEfn5kjxzPfqqkkNZCBDGFSObvVP0STaHWEY2YHsJ9CQ4H1
tkO0kHeH8g6Ypi1WF3Z4ARNVgW3gQEiMJOxJlfuu+8eyGgPx9YLIFmmkWEwvc/D2Eu3+SdcMlOTI
hDwBD6IKvJiQdlEF+pjFea3NILltnNS/nNRyoEVu0tsRv1xl6IkXpRs6chm/AfGAjpmHxEDwxa0z
Z2Iyfaptq7FxKA1e0TPnz2wIVpKbuYfyWQyJbsnGrqF5P9xfJGj9Utta0AkIKIo/shc3hrvEZ773
ZFpSWxptMuF26uDC90SWJ56GEkRu7SevhfYwOgkueh3nPg1A84d7DEzvvmCzLxCnvnlXA+J5Mz13
UBdsaQrsw53NCidMS/HFNkARqHh3bDaVcSKxJ8ZiuV3NDcUsqDEP0sL1Cz55QJCL7CtsAQLoCipy
GkpuOL2RZqTf1jKmAJHn+T91xVBhqwwXnibtWI31JBcjDWC+jKdoQBnQqfId4sl/Y+tqzoRblLg8
smIvI9gnDsJvGyJKGcp1NpYja+DIdANDSJxn5QvQ0D81pPkJJacVaxJ4oBmqA7xZhHU0O2YByIiY
3IVAkMeU7JxgTH23fi2Yp/WTpUvovjRDY0CJX9OALTDedStKBBc1yU2iAF5lBBpTYq6SRtzl6uzv
VmR1f7pmaeH252nCH7PhsMDmVNAHCzQuTDkx+Et2o873pU++lEA/S6lVwUc/V4rkgNJ6DPoXjXBg
lYZcT5aL1avkkLJC4uovXjwuuyV3evvndiHqtDYeC7scacg84iCaDrXb+PYQ+DWPf/TGmlJpvDI1
byDrBt9Ns+M5c2FRUUZT8IwSuKgCmpNdBBZbPjWGH1iIqNBp5BGZwm8ernRTHZnGtM6sLzerHZz4
IixgwZfWLksdZdjj9NKbQeVZ/UDmu0m5P/LXVQMGhYtHuDNYMWe/f31nVJJvwsvzaX/d+dWeG40Z
AQpBqHku54zh1V0sZQYXFI9rRERj5UwD2kFRlVS6gx+vCQ/WuUK+2rz76BekFieGRQDLKtrDxKK5
+yiQMDFBdwN773lFesX8+8+zDzTy3LTpaNcE7MgP4TpKLT1I8vhX78Sej7GWy3iv7osSuuBK7ZAy
wknCnSEk2af0XzRNH9vfs0smR5CQ9HmlC4It3zGiY5Q5oYxcSjktnmtLYp3QF8o1NeZ17yDQ+fXL
xNlKcxNZaVlcq7xqQOBvG5LbqZZ7mtNNe7zMsorjMHfIO7okqGGHAVTaC0EldwxiquXhCRFrIG4G
xyhD1xXaOzkr/AHuMA3sv2qltrW5gGsEJLAwCgvEtzNg8xDxCLjpTm6dasyPeavYP8UAcxPJyvoP
vsB0hUa4gdti92G6tAphCWkPsKYhWogp54TROyCh1F3IPUVIUkaNPCadwARLAfi+R6MKM8I69CVM
q0NY5TBgWW/pMKg2ImhDJkBxc1HJlAL34us7Ri79ql8MaMisiJJpyo7ruuQ6MOmMfk2IX6M9I8jZ
AcDEDDXMviZx1Fsl9UHsUbEmsl85pCvIqzNxhZXwEXFv3G13VNMzOwOQxpUUbNquVhGcaNBLHBHJ
CcEBKxdSZ/og8ayJ2cJzzZqZniNgdc4subGX2FKKIlFQCTs7/oZohCaKf0vzjvYIBDfDz4MR0fTG
plKe4fHviVTGQS1iMl4kbrZpK4eGYTwb2XG6d00sWEpnj1fhuAq1RNHqv811ouAevA6S6c3FDe9C
KKIzcAJOBKRoyrx57Rc1+VHqgxSL+w7vaEXf5rnGP0Z8XUfGDnmplmP537mO3AfAANAwkUqBR7j7
ko2iYg00rMu5w29+b46esgiEVpg14bJ+kPvcBWUp5zan4enzuY5GansHqyihL6GrWur583e8pxcQ
6RwtUeCYnlA+7qjHLVarNJiRv4Vtbwk2JrPHH3MB7wJDWlDn/qVda0BbNorF2p6Hcor+OfUEZ5ra
pdnLRUB753tPTsf8ssprfNNQ4eZVQnOefn9iQpEm9447EDT3+iT9O06daxv/aA2lwvmZTJubN2Zd
ezNevUdbhcSfjnsN+uQXoVJFUCFNrHK9iQcpoDtO+rnqFDDrUdtNReD+7DJPW5uMJD1n7ev6CKA1
C1x9V4yywv+s23KUf0whqIQbLdhSUk55KJc5KC4Za54yvEbl9mLbog3h7wmQu89wwBbOnQFni0qc
5rnGXGiN5ATH0SYI3nCI+flOXDNhsqFhUaUs3+0Ag29WWFVGvUQlr0h5B43ZCK6duG+cIv8U4Dxs
eSv9A1uE85r8RICaLCDA9FCipQg/qCLUWO7t/J/I6poYqrfkBhPoh49nCw0oEcTpX9KtPkv8Z2xa
NBvsq6owABapdfAR7j4moqwPmC06f2KFJ7pqeEmE+R/0DoqxiPee7KCjcY/P5XbzPxBV4ndEefjY
IQNWwqTkRsf4LKeH1QiER2PPYo/tutjeCKB1DeBgsNdewsOpb75/sVXAPxvhQ2AwCFN6VrwEzUb0
myPvyI20xXKDO1FguFDxew4G8IPDeIDXTIgBC+KzwvbM5vnV8UyVADylHTCgUB9U1FQ0o7vuWjPr
T3klFxibOPwUXw/tGQB5WNqYmFtl+6mAbWHn/9zBjRJVOozLsUk2B14cP/mcfws/9zuSYqi3N3sU
FJ5WAspOQhL2SDstldDeut07ubFKnqZUbFkTpVxkpMF+sYiNOFc1dv6d16vjfgwN1xnQ8QYvDGtz
hY4twwVG1bOmIlKsb5zWlhf0qTw+EpMiHsoL7gwtMyr5M4wAWRHl0M6q6Nujh4dnozKS7cIx5/lK
hRwYiR/IAZDtEpuUnFWjKS9T2z0c+/TkDktjyU/+UJ4iG2/6vHCDW8HJGtG4OCMoqrq0s9Cxm8N9
7EtRr0A2DDGOU13uTR+hmbj1f30VgiIvjHNgcUpeqodkKLtgFBX0HUudtPGwalV+68ob7AyRG2Re
wfSXf3lKk/sdGCa7eQ/QO1yQsBejt/N11LG59Lo5mPUU2kKa+EXVBVW4BOH6kePlw18j94Z0pPNx
w3JgJpiYJL1gOBX8Dnxbvj4lOlH57p+tY17SliMYoxL77AjaEeTq98GVWilANw/7FCvEP7Ij3/I1
kijZfAs1uj2j+1u9Rr/OvC9R77b/Km39MB0rBzAbMeUM6kIl95q3YtBupIQgX+Fkf0gAvbbNyyD7
SUt7ZpF6oERFSAXUPmOm9+kKE0nDsFSUT2WyyFgUeXVHfz8vrYWL0jEpncfDRHMQu3nMSZFyFGYu
KXglSe111tNA69Cjyk4Ch+Ldk0aRnQraWHhGp/a9EbqLNdBazTkniUM4OxbJqQxW1HZmOeODSUTH
9KyH6XxNz9W7aX1soHX9So3CdCmJT1B7gH5X2yPn4ra1ORdpCgYXXPIShlFp66BOESdQiRmI05KM
yjKlyC5/6gJD6PoTGU5huTDNTuNvS60a9tjWV30rjIaLOyZn4AEBDm0x9A6HXIQ6cLQXY4qZ7VKl
odoOb7oDAUI3b4aHEz3oFlcf/ehvVDYbtp9fhNOj1fb/gGAvLeszm1XTbNUM9h5R19QcAXcoq2S2
c5H6dwm482rNGJ8Z6eZLwgKc/AsvWnZJidCCv3UEK8kb1bliYuOxL+H4ZymV8mntQBYcmb2ZP6nj
xSrX/2bS5eVGm6Gb3FzVwQT3bx6lW9ubIHO3s7t7kxGC2pJImADABA+oy5d/qMcnvECvyZDkO5p6
e1lY5/Vdf5INTXpwj70iP9uvLeXte/fbloa7W4syicEwnh2mYEFHv6W+J8Bd4qXcmQdE77Mi3na4
J0bXq0h1M1pLPccpAzd114CSCfIjkE0WhkZ4IfO9SchLGLxswbxKxkSzW408KLOmWhBLghek1HcP
uo8D/aiRwdirHqR7LVh5Fomgfq1Skp1oON+k22bF20BKsNy2lCG3rNnN6pczO0bpv4VKxEwsMY9e
n+QCGQV9fjzc2P0CsmIMZrw1C+qEuL0SX/awcw+/hbA3sApWpFT52fIRBS6E4j8OxJ8jsHjWRGtp
JfPM83ed55X0meiNRq2Yd9pk8Jbivu0ZDkCuo7khGg3Yz4frZ1jJhySZvEIO63YALDRQAVR9/1Br
9yVtbWkgCU8pTfOCrNvctuXBcEdeoJOQJaOPzQ1gv6/dNMlVCribtE/BadJZTFWfyJpnhHtAkqF1
LTJLHLCjKNW5MfkFQzWQeLInRSLRFrcLm4F3WWLyftb/iYDe5X5enUnAJK2tndw8bUIyDrHzRHFG
I6/Wx5w0KM79pfOANQjR1lyfjWlYrNC21n0e+F7nnwSH2RmIyH+Ykpi8E4nrO59nn3ddRZldRjt/
ANarAjX5GWvNAv65eomPqCg/VnrdLjff4vANdFDmqjJyK8XzBMSGuymjemHAkKmv9AeGpylfTbhe
Nl0KcxtqlOEzfbJZJRGHt1lDOcwdSu5f48CYazwwLrR4YUft1S3PXZsfQczAT7uTic+NxI5o/oTm
AkrKiMzpsxWr/ipNxN5DuBZwetUSKb+8+3vXm9weSX+usV6BWyJdRDorrr8F51RvSTRV+7bFi4Sq
+h6I+cYZeFrao8a2yJMMMY2zWAwIXmPxdWz7v3FTly8+bShrubI7r1wjBARAfNweZgmocQQJHnoP
egigGFrLbcLyqrIr6O3znh9QKzrb5TyTOislhKUgoGN6lMuHuPCwtxRgMuBo8ssR78Ah95WH7IAu
ISHNBO/toItu0cSeQ8azhcVLPakcLAGlGMsbV6zwH2n3F4KOmMb3pRflGTM1jOI0dMemfOvDMHxK
YKIp50t9qJqK0GNrURUDqmyShsPHkEPWn76OlCbiN2oMMc9JwxK/tm4ldgxzuXm9BN7qcDFEvL3Z
zh49kbhjxxLEIBjS8U+y6NoShLH8AojFBlDgOCn9cSLuNCCbIBJG2xwivIduFqkC1iqJsgQf9Cut
pPEC+caboB9VFVQr7EujVh7cEZzARfie/WF3zpnNVqtzqXaiUpS59f6ut9udxD8WZEmco3PjbFX+
iQChob7tpun2+ZoXHPdCvj6HFbLKNkAwCvGbPTrqoTa4hrSVr57nlLS3mQ9j/ZezQ+GjB4l50rPq
i3sCIfZnEZ85NxlV5Vhzsr7aczUKysSuVRthlv9kdi8tJoyhEh5DJ2i9alM1M5EwH0JLyT8SL4eQ
9jFqenMGBaMHfQ8tbojPMgeEK69YnFrAYQSLINByx89ixC/XjBWsqQbCalqA+UQjx9rDljusL63D
2LA1jjAYnqOfEErcUkFItLrh55cm7kVZ20Ephe16i+2nK/soYoGviE0OGFdCZiitusNwYcKzWalF
PqpLTYf5cF/nFprVhOWXbG8Y9aCj/jrZo40whndZOBCF8iynS/rKIUl1ZAOSPGTgqoE0pg93Uvnp
Q2M4t6LUcMDJwnIV6DgsV9qcQbnp+r6eRXfP48qP9eG1QyzlEOLfFEB7k/InYqgkcuR6YveLIFsz
Ka3VuX0qTmPssgZ1+kolz6M3/2be9xrDUo/8tuvKI3tdn+NP6VsG727BVOvWWE2K05xQdXl6a465
IWFWPa/m8evjA4kqbvpi9Sep6OYi4Z82jqSSONo1jYyqF25eyCkusUDhlsvZoxDOXeC8xxI136sA
N+TqBO5V9w0X6eydO6U9aHMMp/xMytVZ+eZtAOfuoh3LfZLyWOJXy0P+93YxO4dzIXHunINAg1qs
jiS7594NgZyDxOW9MbwBfuzRfOauUou1EG/2JGVjCFsvg5NRgY2QzwPrkPEi14mHnmWiPyX3Xaq8
PFMqxbRVf4b9HENggBpWWfS/uHkKDq8L3TzGCyiQ2+NrgSz4FdF1QVHJ9tli7AKYOw72J5n8HjeV
TfJk1mbb3RBmSKqjnwceaRRiR+ihMAob0q7gOVFVIu1+Sb/ccUvJ/BECeQnwbuO4+jp4KdCWDTf4
ug2NRLiNdVbxpN0KaolJtJmavhEMiI7o4ou8ugb7JWrV8kfIpXKCTAeiPmTGGCJ+er6FV9MWLeZk
wudRc/Qv3w98FuhsIhJxGuCYRm51G623dnjdSysQ9RA3b7VEHe2VN8jlB65B0YdmTe42JRLt7yrz
zIseu9mWS0+0H7wzWd6OxzOsPiXU7IagkIjqVM9puXoMld2DUbhr7QrLs5u5Ba7MuSGo63NY/wlu
w5OwDnfxL6q5tw+ZL0c0gB9MmyeR8SHmzdViZjZbiAsly8s401+nZGU+t3GO/n2zr1kMUoZubx9E
o8I8YsNcvkgP7UFMLFIRyTyKY2Mp7/wKfXXA7EG0quvQkWkx9/5Nda0uJbV3RwSTzSGSeR/tPa9Z
lgmI/ckgRDTU3Xw95q/d/R6tnq5Pqz+3SWHKoBgzajuRKy1ExHUfchsmSR9bwrtEJuIsSKCFTrB+
GdqGcY/74unekhFL3UMC/oiLGKh1tPouian6RPmeGWw0S/lJ4oZmf2B52Yn6wkpscpJenBsJBB1u
VSU9hqkqeNxE3b1trLC58dUOIp9BHJjfn5LSvPKlIGeOyJKD0zafkexPu2Y8ImQWr6Eq3u351/JV
8w26+tLTsgrltpdQd8BGYwr5tPUgrJJItdyDtX/tSjPOnxl4iMcpXt2FgYSOVjgfEBpxb/Dh5jFZ
YDD6AtgI6Y8hKyZSCZE22DjaqSidfsFsqFqevT1aMQ/bOBWmuEynVT8UqkCkZeKOoIsLxVtLqhBV
Tq12W+sxqxFqj4PeyAyftG0/cNCB4+CdunlDdSjvqGwU8YMqbFqaqL/peO1pjaCkro4LCU0bgixO
u3j5uXk+DkQJWkCaM0oIwm8Emh3OWUhO5rq4Cop7BZISjgyWeJMzoX6xpafkJvsmAwBK8sUkz5fh
AaOrg6nLARqJINe8u69jaIlTHPUgLmxb6aBQ9/3CNdKn2oSVukxu8Z53Zmu19p+JAMxyn1F0k+U0
RRdKboskKy4ra/HqmBeMUdGJxprc+2bEyFekO87FU2h7U8+EsRM54qlVNKZvWMuT2TuoERPQg1lW
7LS02em+UNs3lJbSbyHjaX2mskAfDR+XDMiHRHT3fnuokJ+zXcFYDtWeZpcUq/LLV+9Wq954zk3t
Pfw13t5TJuffG66Nv759+b7EfkC8hWEC8E1JCBSDL01Kuj+Wyd+WUtsxro4G3b/oA85Q+hrdVdaM
pkCNjVT4dMtjbXUlVUDG+BPMQh9EXBhCKUcrP3E+Wf0sxM5VWOBvFIngEjLnPyThZ1O4PItv0V0w
nOx8x4sJN+rudHtWsPS6wgVAeG7vaDsrqFzSxwPrCLgc4PrsPkB7Sen0PY0v7/PsYLElpbQjAy9S
5E1atu2W10Me/dR+I607XHL0y4kQmmJIZbosQz8lLz2G//EJcMdg/fBOYwda3NGzGs0y0cPgRMjA
jIWUK0hhc4db9sdPByJOQKL88YhJjv8ywVrCYDXoltG5t7CkznGMEjfrrt7hQAAevzQOSf1xIMIr
zBXrMZr1DRsDY73suaXxkkKDvFGnK28QdrJfSpdBM4mVeXxfDknggKR+aeDirPK6JB+xDImZMCS+
Y1d899IdMcYbPH7BHAEaJnTkmyH0BaBY9QPVsPI4WKt4QHHpY5cHHmNYofSnv3A4IyILIoLYDzDN
h30bcOiuCV5jCygUfVt2V5TAChFAK5a/yPOtqmciFTfQpA5BIyU1i8m88t7jVWEFWMLGEJrOGavP
6UHht14yWHIMT2qoZGao9Dq6Y1X+D3MBbPIKvt/RQungiWSlynilAxj5JMEtDclg3zqJSGj73rhc
s2cqrUqqwuC/IyzHCzGGguyqsa74vRbZ3jZLAtL9qWagU6CU47149/3qrN9QaNvf9NHuMUzG2WR5
ORqHG1aH4PoyC4fGQH5pNhosU7KX1UoqM0ek9RtTK7jZn2fx8qZSccc2vDn64D1pgeoeglw1raLB
4wd4lBrjSUWfo+GpgIhF58FfwtyjZckiiU2NOUBwmKY/Wlrc/sGj5dHGRTPXqenT/Y6fLPMxZSsA
80GaJYdU19wey7dZ60bhl2nVsyE9W+0SqWEoNwiH3zpW/5i8WRI7TaLKCx+k6eLwW4/xmvrRktcF
CzRMSDtq72arAJtiKpXOzKzOoZAF682dLfXp6BwCkAE3xLF57H7plhb+v3mM9+hjmqshMsEbTaFi
D5w+G8HBI2J6aDMXeDRYwfXPTDUAcF0WPdXrhGc5721PfE1Ccz08UEc0JUPIpVVWUPAlvUhJ6HUt
efqQdgldQjlA3Q4kPpYBma7meql4EgIf6JB6x72ygHfepXW4Qc7wAnD+XAAIXgt6nRQ6LDBn84Nw
/lZhilIvCrISd9TlF6M8gkrusiu52bSS42CJUbhdShCYTsUgboM+eE8+EV9Aq4AfFPoHncMC7zzP
ZGTKgW6o5QbvVzPK1zuyHP28GwwWaIDep5D1PdfsWRPnqijzDmNbKIBgUbyQnbeQSnhuM5eAN549
OxngfL3EMx05gNAw4W8BXbgsB4+sOHW3EK/MaIIpC2M7Y+Rzvvb6L5Z5UdMCJHJl6zwIcAiqYrae
u7habMrMkzf7MmWFAIyYWnY3iWkcUgPS2Uri/TFGut/5JX39XCYBmJarOeGpl/UjcFUpf+rNXgZm
z0ZSMGpM3cTbBlZ/99Hw7w2YYxyVUAHoyHvWIkU/qGSCeECVDEoAujKVhJBWfTuxkLSxpSTWgiJl
NZOqX6i6P+LMqCHak67D9UFSi7zJ3CjggUVBh8a1gO6O7GxLyZIFpRUA5OcbZLv8Z6hKd+B7zHYi
tePUxkGSiw1kNXjXF5vpsdAbO4RxYxdvkJWreH1hWN0+C6IkhUEoCdBnlOR38eKzcDqgtRKsjRdI
Nwdd27dq3jQlyrQK883ofwpvLMe9wAjWBhW2ey266nh3edgYyVcb5R/oPj1yk+tHXiWcN6bA9l0v
kda8cTTW3hq7uU+CHlcn1XLW5VTu+3zqzppC1yfziMYxcEz45BS6d3FdfErZWPHyO/6DAkMHNp4p
RTUfFYzHJK01znbTOJFgFHRlNhr07edSvjTDfoFnc7YU2T4ntYpx4TKVZDqif0pB4N0eELkFSEW+
xUWMeV0Fa22BUq9tuzq+sY+io2uE2dhySIAjhMlqWA1YdK9sYHvaGK7Xp+g/kNHoEZE4jUJPDwqS
b3mZ1+4HiN5is6eGKf/4aRLxzEBbFhXe0HhQX3RDq0CtgIyJE3Bc7tI2DG6+afdUu38pl5Dvr9KD
IFyY4mVP83g1kfU5b85jVt8P7HCP3h/TLW0tLKiJ/SHKuZI9TxpZsi6psrXXJ65OyZoaMj6Y1USn
spOYg4VGWJ9W6xyUtDD6hhdwogA3wWgtJw0p7wAhtZm/TkiydLy3jc4NRX++c2wedU0jlTL4rhG+
q2cRPcZsXH3p5/9xJxd6vpDOqheuRfj3UfpM4PwSDB3MDHUBaLi0TaWJLRKLRs8/59s1auvQbdFR
9MjP9q077gkIqrwa2c3dFvo+nfk7KUa0paZzqydliOsuJXlvD0gBXg33I46qkKmmPCqMKY3Xg3d5
QgoUJjiFY+UGQeUXkQghuaFRIFQHmO2VcTzcXWMViAXPu+sX5TJHxcr1581uMQHIihYrxguHSG5z
HtuR8yMOc2xiBEn3M458jyeER4zOKleIQG1tL9BXlKkUZpuY9Jk/rhZscm6hT6G69tNVLcmOw+9t
Nr5qRFd9RN9QO2EiZpNhbzEXn1HHBAxhnv5qQJwUBBKNxwZQ76Nq5qEjboPaxqUq3hd2Rpf4ESAE
yO+6lMckZcx5jWalyS3w8ubPD/DOjmjDOk8mRGVQxjKJsrZPRCiUR4fasjPwabPZ1EUWWldxu+uv
F3GjoOeSoQ8eGsr50Ln1xxRhNlnBNyIHMCDmLH3AxJmexsE4JOT+nPcWU5A1tXzLEvNmyz3XLUp4
mIefJ3Iir8YfpsbAeAYvTXxan6n7UXLMHt1Wx4vmGokdmNbUd/4k36JF/Niol5PVNnzUyJ5vjBGg
kXRm7oIJSTNMOz1K/dJOrnVBezpi1ZHX5Huwy3QUxu6TIqSWOQq6TLGqh4SY3sXMYDA7m1agMD3J
8lKf2B+JdUYxAvhFz3+D6V0nmdrNf8kkrX9myxAbN/RvM/32GzXII1va4wPknWX7CbLqy1n0Wjid
Rj+UQyTJy0mXqEZVnsGrJCPXt/Giu5912AzW1rLQz0+2w/PRuy02wxGr4mRIKh7VOAVPt0MZGYp1
C+0BBCEdVstaLRT7LCH89Xsnxcs+oBFDYBZlYmYSs8GeEv2/0WeJEf/NfFNOZX3j/z1yhXMvAQhE
vzPFUxrzh02VscvqAkihgX9V9gEb8hCVNglMBIVLJy2IOx7R5eBJmcEGSQqi7/7QSZvvsAMGyOtq
SvpYAnv7BeMJNNxGmnfMw5G/r3WZHcNgttElHMomb8BxoKbs4SpRNxN95tW3R5L2i6dS+J2PSUwK
+l4tjxK7Q3OuEjLFO6qq4cKjGDFlrxdwFQejeqUGx+UrGXkbIcMfoYFsdvKtkqTWgLgORi6B6eWE
hCG3AVgIpyuBSKMkEQulS+2GS+gDwyOV9f5iEoJpFT2iWZjTOpoR4lx8A70mXrnWsCnYHMK84VFh
vnJzNv3hZ0SDhgzW6yeCId0WBt3FN9qiiRPYie0mUr2sbuCdTDR2HLBymXj37vsOn9RjFf0v0Yt7
OUQCHWfVf8JOW2LjnWlCJW0opN0VnKxOBGePXRq0v8Q/z7A9+XMU1/IBff667Wj5m5oulL/xVZBH
TcolddOmV3LyyJ/RWWt9dmcCv57VgtWLJVV1EnNJ78BA5e9JqsaxGALXYPwtzxoxq6KIj5mg1VDD
ggFiILL95FgC8eHfQOgII3ZNP1Uax+ne0qFusQmdA+lOrbBsRLO2hs6UqfYyGiDesU2zF3LJfXwu
lN1pXk6dp9RwAiGhdVSuiTEsUJYE9tPNf7bdxthohJiRdfkIHg78sNtq1sDP/n3Nvv3UzUTV66T/
dA9yNUuzn5qpHByMpnieC0GjUa9B572Vvms0fME32a9LBRp8em5IcDRlvkxl3SOKTiwOuOcHkVcE
KRDRp4JthfojgbC+pItSLo8wE97AdYxEhJHQ9OwcjFPaP507jIPmLj1mn+Q9/2HFHC/1+N73b3XH
wBE5zbJ6umG+PWdlhKrsQLFndjikGuWojLOFGA1ZF8EsgsD8cjyRAN99SEvwN6h3a23zBNLdTLk1
8aekTbp4sE9EowqIRNkcmzO4QDWkq3HfbqEgTn2nIgbdmuO6nRq9Ft4dWb+4c5maTVtbNtBm/Rpd
rLfq2LbC2VU5+uGYodV0Qz5FWoeyxA+amw5odkkISvi18oDR6SD8HL4UkTPBU0ZxMhJKDPlaOunH
/yLWRKHcIEFF9nyhGb/DM0fYmC+IzQ6d2wSaYP8x9Yk8ycv/DCdd4rcziYrzIgN9BAhYs7S3hGr1
LwcvNNcvJeu1MZHw7Qa6VEhkYrGHS0kpMKDs0MV5cMjUghx8KCJ8Y7HdMmvs9SAz745u1jqxn7Ug
UI+3BnsvSuangnCjGTJHgcN5YW1USQCujFYiSVw+rPwiGS+SSKcA15dEuU6gJSyos54Kw5sLIVBs
HLxT41Z0VAHXqTBHoyNkHNC/mfWROS/Mslc+d0Vb4GPXgZBwzCVIHJ6A2zBY9X3dA3U6av6OTj6H
Tfc7l8GTLWXReE5plwG1W+jD9TCXB0MSHb5cxxok+ycIzKSWnHgi+FMjhjXwAdJCVB918BqhMJgE
4x+/S9+vSQ1ZItiGCVp+0WR3xh1KVUVcAltrsOx2Al4D8zdM4T6AfR8zW/tp3XQVxkyyxcEszjUu
z1IbIKYdtIsOeqvwwO+aQgn1DPTEYsQTuZsS8nI24Hicc6TyMVfc8TL1IaCsBaBFKThjESJrXPoF
IUpSFHPJ1SPLljgc+084dIUUK/cCeZsHR2eSHHyDK+1pzwIadKtQOsni/oDZzyoHmGDrcvcTwRpt
ViwHERlmta+9vlp3LC8VVFbzlQNy8VllYL1rtYA/r0Orgm2F2sNX7vHHd1Dy0MJd0r3ogi4a1JYO
Zi9XfwWpXp5pO8tHF7Me26LWHS2+ofTeAPiVf5hY8qk662UAoVLm/ZdVOE7HOdoJK0fvCLXTLuCO
5HNnqQXQHP5Bq9sC9UCxLXNHd0ZeelA1Mbi8h1Eket9MmQm6k/ooNNLSiHnZQdwd7RFCge0vhgYy
m/C6iIaA7kgDXTJTrF+JqDIlUp3qyjY1sop1N/ujNyDFScKmUUvpHhtB5oOTl5utKy9pYIFKnPJn
QKyA4lE48QHL79BYzu21m8hkDgUztnUPjzn/Sucp8g/G9uV1fkJ9hkP+mezfiTLc2cXPVzHlHiiZ
m7lkn08qCtpwbkj9yy98sanAUSa1g8DrbXtdVjQenDP+lOcdMthLk9B5d5+aNcCFKR9DoxgMEclx
LtW0uHuBbHIXB1jIRy9RQtnzNIHQl+FZsM7PyWviHJqXKe0BZyXrT3hb7uZgpMN14rTIUz6GVPkO
dGE5BDxR+8bMQX0/BsxHpnegKDia3oweEYI9kFv44XX15vawf6SPgz1vvUJf0Or9gZaYl5ncsc9q
Ic3XLflDjGpsVA6q/Ds3dhpO1al1mg+32tQ4xxWe+7G1//3VDYaMnW8/SpSBvYccGpzl1xw3n9vs
f6G0egkvpPMxrAir3sx1VKfKDoMmYh25NYRPiSbt0GiEeF2gFgNvh2ut/qCSUbzbAZn2z1bi8H1h
Tu/jzRz//411GmmppDMl/4aLO5kRvri7mVDXZ90pRlvfTCw+oke3wxGpxputIodi+8J01VfXhAzh
HjTUlkIec7iT6DhZET5FHZ3rnyR8pbN0DN08QxRRRdiYwgPp+hSy5ABapXFLuVijk94vpkJA5p9U
is/AlwPq5+Pze3dWMReFyzYnePRnWbbX6I5ghvhQlF42+Kki29EV6DMNgaOW9Zqr7+PChyIcIjNV
O2cVe4VOkWWPt91sjeqJJLkkn1RV07wjfquBXIc3mfa4t00PwgkKCfIjSv+s5Je0TXjN+sD2yLU+
084LXypkxSPvV6e/BSDIm4WnQBGbEOWuaAVR00jKqpk2prt9L3pW2dA9cqVSqdZXWu6O1hfT2JVB
gc7E/h0ZFYUW/XYYua1p+mwaPqaF9RtRRg5NCRQNBMIJIn2D1L1hVGyBW8R5lM6NP8tPFIlQ4WoW
bFwz9/6WjUvSCnL5ofiLv0Wl2Qir08oIbjiQ2owynL+LJe0j1B7xQ/nhOleqk1Or3vg1GVV5Y6Ty
qJCAWCrWBizy6+viuSA8jy8tExphNwt24IeuHsDXqn5siXryrQbW9FnvNaDJt8BeG/0G0N2Pec8u
XKJBICBmQT5AbLA6KAYIjauRDrWNfbUI5sWemXv+K/31GdgwU5Dte7dIKUJn2YzWekp3R0ZTKGAO
0sZ6B2fUaObmVblAmsN1Q4TW5HYfrigxG4fJZMfA5W7ule4aRLvRkrk/EMWYLC+4w9PSqp1PrOpR
s1UGiRLQcn5LXtQlPQZiKiSvovIYKx03EpQi2/uIKgP3b83vpuJM0NeMvs2BrINf9Aax4SvjNZCc
DrgtjTKJDXLAi5KY7L5EC3cMIxsvkkR6i6osDKDXOSdsF9qgLaovxo4FmoZ4xMt2x3Zl7pkQIG2v
5zKZREjImcvmBiinM90gw7LlFoDZ6jBa20VQr02yeolmLab46t1ZtKPRLCMDgHpSADyDV1A3Ouel
ILp2QyTMebaDbFVq9PokOBgVKiFPfKJE/NdzbVOZFllBcYX9GdpsfH7tk37d725s1q1cJCluMOxZ
C5nLQr7fj0VfCHbaI7B4tgcnmuVaKLIPanFOnMSBbunEaD3t2jsP148MvzBCBDHzJSMxtqt35K1Q
Nuccj5SMd1FktDwSCebvOzY2fgmxD8P61VpNMgTiFwjyeCYt5rNVQZHOL84J4vWw6LN8j1zpJXIj
YvTkM2W1XMlncaDVKtWyIBdBPUrMZQeAj8s+lKWnDNUSE6mcunxCCsNilMHzNjbRIpnPXXa6gG1O
7mYfSkLLOFdqaUOfhIef3ewpuEObmshevtAwaCelyp1x2Z5wH6NDGvrOcs7X0SEJdGai5SlQjOTh
Wyruo5sTG5cDZRtHjeA2kQF9WldL6pscbL2BTJYCH85DxpPvLkIKjI2y9iWTOt1EReb9e39y7LNx
wdirHmrvQlyiCbZj2N39V7ySMomxYU64M7qROJYtcuWug1pMbb28ZEAz6WQ2jII/JqbCCmjBd098
RokzrnEfAfWlIhfjPyZjnc/gFtuQwUBlAKjdO+m0cj3B++n3KEYdk9B6l4oE0BU86mPbTKPUaomh
Y3CWj4v4YURgY2/FJGKZjxhiQZdRUPSyRLawE0BtISQ9Sz94maN/+rn5O2Ne2EwN0txFb9mbU0G9
1m75e6A9RnJxozRDz50wlHrBecRyfHiHEWL8Z7eewIer1aOWjCtJUVCkAfghe2aWMStiUPL5ZLVN
K8oXfPA5NrbJ4AsX//qPihbHENwLkk63WSEc37LotGuf6ZaWq/aFHa5drOMgJ4w7dCjzZ72th/6g
7YhtmAdH88qCT8c6LE4JQJSp8cimTnBl9cSnk0lbEGrcoRu7Um1B0gZNfg1bKmaznxHhNmrgE+zQ
ezuuuEOv4fVZ+uADcTNm4WWXkK7nQ5h7UxeEhdPy5CD3QU89RfLxAttAg9VcidwhpHkkn33Y0TpH
fOsTxLOTtmrSIhAqcE+nm6NPiBVey5X2N7hbYJQ2dNbxtuPKrj+iVClu2ZzmnkOvh7ORL0P7qz4X
ZiibrJeT3xorea5/oNjsiDx1vyz6UO3bugMkWp3hZuZ6NB7ANGOvDtvHToJ64VzNX8Y3B82mLN9o
yPC4rRUx69q+KwxAqp4Nm4cM+jb5VqBZI6PTzSVzI5zWpSCPQAOXtp5jFheM9YqC75CewwIMXEXy
PvC8JwKxuLDF0XUU8pZF21gMqFnUQcai6wV/RcFteN2s+R8f8Wpf5s5zdsz55T3KgV2wrEuDqTiD
Z1YFDxkWsEdDKCJfoO0R+C1XsYoded1JC8fjslBDkN7OnlApMlEju8npEM6O/+6nauV9K3MKZ9dr
PNumrBJI1p0PBKo4+olckPyhMk8bWs3vLeO5zr10rrtALD54olDQcJK2KJmiZY8Rx3ctco8YUCKe
KoZ+ql/jhDHhtnEPp9Rd1eJFEUzcQC7bH1aJ+pDs1yUDyfdMMTWcTC1p1OwsnowTrz6/NhcXsRp9
JcECNeKoEjPAQopAWfhPq68nJJXdAS2qJB1MYNY+TtvPBaIya5Vd1lra6dhCfrOXLGNec/haBFGs
nyQs+/GE+GgKXR8MZvpWC7acNHZuneD4AdkpYqyo61ra0DI8WBtUASh5+9UgsKvSxxX2fGgJXrGe
b+4/om3v2vxZinrBkhI+Lztsc6H6b+XgW4eMqclFhjP4yJMKfb2K5eRwyeFvMTAjz9R2Jxui5+Lg
EQgQStHaFG9onBUgA2Yjo16eXhD55S49yzxm3DS70JYhDuF6/6N75CRcnFIAzRVJUJpzn0Zs4wba
Xl1gZS1BSpAjMg4L5nXohqpCo9ntJmrA959GuUHY/KTWI7rOTEIt3YEdzxFBZAuOigu01O6dpw8X
xpfWSHJ7Zxe2I98nF11maI4qMJyEQLangusFfl6kpGCy0qHpsjcQEo3YjztVWMP97jgbQ4QOm/ei
W5vt/2F2HTuejsCDQWkuqbPUBykPQNqmjk+zqRS4tjIyogPTOAS5bruRSLIhi6dI7Drk5hwH60TU
I3QHxMMgIJubkGO9YDxIiJ1uvmQ52OedK3KWW8lBMZkZIiRv6F8+SIhWifD/FreR5q5kNIeV9McQ
IjkAGFaolopvBnV4cyDaTbSaNUMLeD0DOwIPU3HBaY++cZ+JXW42xb2LVR7IjAGF5P7v4hHFDt6B
6l0i4MYtufrPciQa/9Y0MZVkw5G8rAPQslaM1NNjncKY3BUW1YrPe8LCw08dM4+eg630SbByYX9z
qNFXvETF8aKkSOY8ml0y/sHHqKcQMB8x6eS/bXvtQgnii78PWCxDg6NabTbQ6r1GMrxqMLSUjgeS
s4fGWQmvKPPsjiCBUu7XxnwzFhBaJHufiL9UoX8gk89Okp68fswABi4cP7qkTYXrr/TuGT0dMKJM
GH7R6fg6jYZYZ7OA+dXzMDgx6RbQ4Hi+v/BSXY+pV9iRU38f16PQtkYnB+cOUVt/E4ZQMuFGmXYP
FiotkuPyYR56us7oPizyl52yFf0A+ZEn9P5jxkPAmPseVV7t1auNwNs7e8A/3kYFOPHCYkcUvbNY
gqHusPq/DMtrwdcf8LDJVjlJUzxeknV32v5Udek31gGaRr5bpo9veLPvLnsKpxICevpicyu59lnz
LG3CvlSIii41CFWv5BNkyievENamPxmrz1emgA+YtvzGZa1umgmNkdoDecHoBKK//if9V0VAxuNT
qT75YfuGGJhdxV0ZtbUp3Zz0r06apv83vWG7xBQ5JiAxXFFltz+2OP92FUwWmoDgLxR3URGDnu8S
IzTuuous7sPFzwA+0F3Pet0qC5MABoBI/8CNKtl7nnMpJCAKJnFse53/b39eYJxw1msRmcLXaR68
4NRlXBQxM6Vg6Yo6yLnGNyLjMJ5UwXKwbWPXIt6EgWpnz+YG9+V5OLuen5D2En2OL1iDx6UgUCdK
kQJ1NBoimcKitubCEVo3pgx6aLejuwmO1hOC9LKkaHcFvkmkMuQxZ099c+yIhkCY4YZP74x/xZBt
APz9v71m+RR0Ow8+U6wnuxCkIPz2M4CLz1IeT4drEX93bNmA51zpZZMd5HwH0s9Ii7rIKeIhbbuz
ZcvAIjj9f9dtdQWtMa2CLu/K+x553ceL5+3BUa8UDPE7jW1T4wLFWsl1rIvT6YOQUFyx6DGQUHWA
bYRBr4Sa9G4T9N5uxw0rk78iarr1V7rfLeQvOTOYc/A3Khoxu5Wz03oiMhDilNN+GH6UE8YLcnpD
jSWNV0x9BNfl+zuU5Ft+isVFVnD9e1rMIJEIAMe3KZGfWDQOwfniMNkDDdBPV14l5bTRQRIWQ79b
dpB5MeXfuZsAXqwjbQqWBnOTWZv9L7Y94Nqbl1xdV3OjI18QDS/zyX8aeBpC1qh4f1azPpzb+ldU
7ZAOTZciaEI/V6DsRRQ1LLQl/+wX7OY2wNDGWmPFOZ36M7b0Pv/Ha9aW0iE0VgWF7BYQS/Luz5jP
MFIHZEeWh0aJhI9QSS3ysd7ZakjxTwpGaFYF4JLYQ1/0FMNoWgsLclbtksPdlLLoApgelq5ZsJ3o
M15dEQWBF+25JlN29aZVCYfaF7B+TF++4fA74PdevrU7xR+zM3K4H6SC+stQjZj1HYZvLe/L/GkO
0Q/N21zGhQfp8LIOrHNH5WQm3r+S5C+wgXzLZZujwllk6nTX/ez4mwHXABEUMn4/04glmzWdhJiH
llZ+5S1tlLjNMcGuoAAClX7q9SiRnEmR2OCNrtHevtCMbk/kCn9rQSDg/YbnOUI0V0O6GaBYfqgl
V+Lm0ZE23MwcUsXzYaO3jmsG+OiMEwDnsjeSV1Tg1cVYfjPT8iqDz07WTGoDsq+CX8oajerDpsrD
OBNBmuWoTJ8KVEvl4LPJApThBAzQEm4qbMXaXXuQDOo5oLCG041wx/g59rrNtBKMmcnRFIU62a7A
XFwjDsgNDyty18FznBcojrv5cAr84I4gCepAP+sHF9nrHqzH950GGrRQ566N4Y4MbORQI4SmIIHK
CUG2IftQBnY4PZe8vPE85lz+1TQlgBKHnolVg4vsdZ3B/n/NxXtv4yu4VICnWMAIrvrytBxyny5x
O7VNqIKAH5TJXKwa0ZZ2W3n7vGT94vehQe7EMj2kX/M3XWhA+bpGWphYBELSu/zL4mSpDMvWbKQT
wNaMFgkO4fe4x2eOM8B82bXk4kCIdaJisVi1N+ds+63f8qLwxgljWq93gE2Z0WVuhA4xxeSrv3Lf
I1k3Z382elSQI2FpjjzUGL05RBrVQdZ7BVRdEQm9ebVrXfRy8yfaa/+pONaMMnTCtTs0m450dOAT
By7MfQXZBQKgu7QRQqhpkiIWworn/DDotnSI/KXHRItDISlFXKErWNkebdM4Sf8mjukgQcTpE6fG
mtQWj5ncBhPruXlDM1HZxGSLyMKpxku3WU9RrfxMXKWWAHlRNU3c1Sj+aaECzzbQkRSm9GedVI5W
27fbsXigRzcP59m9QENxZH/oJrgTtEAVW/7malDJ39R6Nsht9TCLPb18EwL9shwOgfJJrwi9hR01
MRAh9FGZqtRV/h7gQuW6oq8LWUOI1bZHaC1VYAj36ezxb9OqhM1YpgT19KpnseXXr2ALXjrcSnm6
kiLk3MQBtyNg66qGw3HRYkYiJc/R1NiV/LWoxcomyHloMvN/Pgus6WYdTPaVh8WpC9kRmvyBphUe
2vM0reVdbyC7vc8ssLukRdnsLT8Xd3hEmvZq86muNBHjUaLOIVH0kX9LuoutFuONGi9Q5kexdJp+
movYczDwhHqP+HQThtlgTsCmf7nwbaPByDUc0hUVdqyQ8h36iRdxfbfjeb2VAT4iE7mZBLx5KyZ/
bBsjGgfkQfDEMKTwOlmW8l3h1NHuDuTwNt1+o0EdCZP12clCo7U6/X5VQPEth9DFmRAyF15JujH9
HJxCgJyZLRJBj/wRIE2iZ1S4+mA6AIwIkrpg5D8+pVPIbHfjhBcmf9qKmQ98ySETn9WI0GrdTR19
/Ntiog4G2nius6ONxClX3vMM4oPm89glEs1FkxeiX40bSig4ozO//WSEWYJrOeG+tePWR25QBztu
E90yG942vIWaXg3LN1XtUXWfEU8XkR3gbjhC5myBOiSpz0Y7KjkUj7ow0l3knSDayFlOthadDPKj
230jOtTQm46D0zWXCnkzEXHNHF4n1bDB7cywpDzoUs3jgWvQx3q92R/T1tGPQBg40U/UeJchNB+C
swVEBSrwFhVSCBETR5gU4oJ7OysLngBUL0XD45iDhde4iNPmpuQ9wMuho0gusE5koi85KjBo2Fnn
gMscjq1S3JJTwn8QGXSt7O3tLW0j/0W/gpEYCHsFU2wg9yiZshabmASPFUi3EuPCVAH/5wosG6WQ
aXOoYYzOccqPTxZ9yE1eCkla7vC5AhEiaWUKA3z4eZA94uczsOUcUbUvz4bJ+90y8PkFWTn8AYvZ
yuWtPOcmt38n+pdJBn7mDvyxypa23NMINk6xEubsqF6141g4utnp6zyUZ6eVQ8etP9TdqkGWmL/5
44MsdZruDXakMM4DkRdriqOALxP7rB4PcsuAqLUDxhqxILWm/5EWZpKElVgwwMcd412xrnked+jv
mCnmzOlxkU3iHTMAnl6HdypMv2hGjLAR+yXFVG9OmGq0+MgPaHXyLB3uLlQTsm/qFUtwrPvZo5j1
6OYE6M17O9YKqjTaUqbAxF9WXSMwoOU3PP7y12CIWmmgsUSpj1dLG/0XPtnBhY/p5FmwlmK/K3YR
8073nzDs9x7aqu2Oh4te2WB6jJlCK65a5ZiY94mVOIt1UEu+dgIV1pSlz77I3cX/hsNNc8NhT9zQ
t4Qa3yWDjVhC26y2uJBvbBDkuLUmObh5AjMwzYeY0VohVwDJj6ftgHMnzttqlesL//aEQvDG5A5y
iooREH8LfdxNK+Av+KJk0G6iZ4qvTaXq/XKYaIqcC2SVU1gy5DyL2sw3FVMNcDxfF19kura0ec0v
6HG5vCfc8GAO58X8YAavvy/iItnoEn1DghOqyNofJcOKCd7Abg3y14a6g0eHLqLYKvG+32/Lf7iB
JNP8SW7xCFi8kY7CBCqC5jpASLEWP2qy0epvQBaGC7yNBAPAJumfORC3XTNueY9/0LBYE8zn7OdM
rtfbjFEuFEYZPAXbSDUwXEKECamrgursZRYtgaqvbBOpaCB5eL7pjNOQiEW0u2cf9zERuzUVYEyK
jbKzRfVKxnhccvxSNq4GMVvuEg/47ZugctiXO11/nFBmgVY5hVbx7z5DHf8s1+rWMyBoQUz9Xx13
8uj3EgW9iWcnOrYkyJnYyV9uWVZd2ivaTexk2xUct9eoa9FKdutYNJyZpTzfo9/DMes3fgSLPjwr
5GPGq7qrnofI2Li5Z1XcwKaE/CW/en6IrUOLoXy6iyM109kSb6pAZqsJgBkNFZKiolpqrIWbDeak
z0Qg37VbxJZFUeLfWZw22mR3RaRBX72z14QcijAd8c6q2EIr2gOogevleGfWtuLwrUfh9nLJpq0+
+XmwWkInONR30vz78z6m283a348RabibZMNMzBIMUvpn+LOKd40XHtRTIYEVBBnx8M/FdK3/uNfA
K8TEwF3hO1J6HXlgGhU5k3GudL/gf1xAPs/c15D/rCxxffwkzi9iE6ba2Pvk2fllkx3Gn6G7NX2I
eVzwLdi5kwhV88ld1mgo/OG0R9/ooXU6E4rGKnrBkOU3ag2UZa9izbNf+cLbDQ6cYchSqQe4Tx2L
6UD8+NVr4DMPIHK3kSXPsoQKmDgQ6hfdabtUmCZTx4jsQSuocZ53mExV5xX7+4OQsGtbdGDDiQzM
Aat0KMMA09M8ot1hNijXhU0VPhTYA1/FbK0/TNwZhXcPnZkNdC7/0vdr+TbAKQN7+15pJari37za
Bt3kVqmCh5B1b2sZDjghsKn8SDIgpZi96ucMSE7cPIXgMVZ6YF7+Z21Ht6iFcZxTUqjbzsUScszq
rZLx4eNOD7WmsFJgNAzVM4NtQ5ZLe0BJmSCfc5xuMlFVqOn6dqq8hfzbZDWaZ1gkZ2XXWSdOhd1X
PFWbhhLXFrcd/tW4RtByqbR5yJPWxi0iQE+Vw83YmVlbuK38eddxXMYcB/khjpehDUIjZP0NuS7a
N59cLle3zsd2ajRmCQVn9WwaxCUrpjw93Ms8u4/BB+056GlEiLesLlivqdQasIYMIdWhSbPAV6y7
rF344VU7alfo6HvqRyrT8ykgRMAHDN59Y6sIEHh1YD/99Lt1imr9/yJVlbaq7sA19El3Ur4oulUc
KwuXgEwSfeyf4DWBov6fteyQlIbPK2NzrUr6EvQkq9buwvlZXUDpIn6LhC0lC/ucL31EKN29/fvg
J4hONxpnPNRm0sKvsCflbkuBPzuXVxuYcpa3D3H0HPa3XXlc6I+9C2KIwiNPf1m6Whyfg9StQfhx
2JVkTFo9Y0CbcUpJDupr/B6qNJjPw0T0vlycz/vVPOnNDY0BXtdZO9jELvKlhCwBbg55tBTmBe95
yybhdneTggJSxU76dhkulQfQ1M7d2yclWCFGaUf9S2N3ykg+OJT+Piokct677BVVs1Fyrh2y3SAs
B0dniKITsUX/JY6UniEQRvpvDJDSD36b1Gj8bJpFC5cvtfriwzxbOJoQRtpE+PBoC9t6AMh7baJU
7qsRWfO95USgJqv+JfRilBtA+8LtArXyy68cscZBewnG8mj9ztfhFHCEH0TrWnu/00fUQyrqlh6K
+BBWIb0zTLfSyjerHgFNjZOVFWhan1lgJ6ctZuGTfHmPlsWdiWlmuvfiiCuuESdj/YYyqqmuaHbr
wedTvBmxknBoXaGj0C/o/NssbFPvz6X0+xTXDkknO5SM7btCZzKAyYU/vSJFpGK6Hzxn+lFtIRib
ythdzZ94B5RLy4rN38T69jjWxWTZ5OouYNw12znoEhL0rzRxJnM9m81e1nr8My1c9Gm6wp5d9BVD
YITcYIJylkPguiQMk+c9KJCNW4Y+5iEvaf+/hZkKBcaWgDaXBM1H56+bGSENo+aJ/Gu62tzalg/9
+2AsQA/jiI5qEKDfTMvXqy3/4MeasfsyZHpyNFuxkfDCApHQG7NnE71ca+n8z7FAQzA7ylQwr2hK
t+LR4ikAw/ClDRg8lgtmm1TjT0X15ZXWjR17leRUDsQ/Q8gKqLOxo5hWaIbWW8kktlB5XzrPFNyQ
eOosH/LPMUKRPKP0ttoWg90sSBUqEt3LonArdilZNgWs5luFlVqrMGoA3xxUGbpjVSihpl+Si83O
ZWrGsmL0wAatdpZeiMYXsRIawNCrBlyQ2EtRR54Ce/iH6Mc2DZDG+s96H5GhJ6LzMpiRpKn37dZl
aQspmOMAdDkMOfGSYdRI26SqQVZ13cIIEliIDkXg4XMWv49C0vrj0APMntgxnfXW/mnccbRMPyzW
sp5b7u5TYs71UNi+ZWfELMw3oOt2XA4opdezKJxAFpkIZlasRfEXDRSRQggdUzmvFKkENMLA4N4J
PTXoPJU9TbP7NXcS4ogsT/LbmTlkLD6cw2RRb4em+0DNvqtF1mIWS5ZCkqHelsPcMbrWs07FBaDS
3O7XK1rX9oq6Lwi9GVV9IK+9Sq1xypiyZBDq7FV5aXYBhRzVkFAvi+1dU3KKwjpOnlfg2X8k+ocy
Oxb7epuXOA120+UnYFJ64NK1K1bIvqGQJTwWSN6R4uI/T6sKWtc5YrN1ylxhHUbaopJabGnVavw+
hTlVRjfNO0hU1u3RFAP0HUjhDGJvi96+jI4UllrXXMCAFbQFghTKZQrt1GSN9KdtGkqNGbM17fs/
EYNXPKgPKQ9t+rj/HL0CeKT5J/T+gK9WzZ7dGNDtq3JnrzZWlomMeJhM1UzL0H3+HhruVVWVuGN0
sZFhRWvu6u0igx73p0/AxvRQd0yUYRmqvgY0eTjNBRpiBblaWBYnfr6J2mJ1p3bVk1Io14xbneEH
b4lSkt13GUq5OZf1T8Pku0atq4OLoMIbYT+B7B9329ZCPbfk+jo5KoL38FCuBzmYxL3x4PaXsmjp
8aSedosMhT3s3SBoGX/sXOIbrQJPF+QL0jox/NDGIa2LK06stlxU4MRb407gHQrDyE2vZ0CcoT5M
2QZRk9mTSYg1bIlt1ANAebG9AjMTuMVzgnl7kR1wUI7gdrU16bxhli7/oPO/I7iVFcYC6A66PuR8
GelBaqeR7coKJI3sY4M0GNRrF0MaS0bG6OXFd2QFvrN/3ejwuWgiG/yX996lIxydwHklLf6mawNu
LYLYySBAPpz9fSC5mn0yEomn8wVQ2gOYigGGdwY4OLMjIX5nyo12G55K/GfgDt84ScX0eGqgc+uX
9HPWV3mthtOBA3YS1Oku5q2Tj7dKVRM37mYsFdx+GlfZbg+tCc50h8jM5EhWMi0lq+On7QMoSmWk
JJkBN2nhseBCyTlApBYJAT5ddiYWiH7BZR2j0C3uuH4wM13G8a5P9aqOhShz10y4EFJBwa99K93R
HsjIs6gqCFt48easJ/RVpZPGbLik+rSd0WMb3ujrSxmsa4ncYPXSg7zZnFq5KQUPE6ax+g6MLI2S
zwiyOsYoOn47PenYkhQtkD4XXEkU2nnp/uleTAbD7KudtsIyuEqhL/7kTQuBOolgjekDhQrBIPkz
4pM6RIxB9ftkTqA/pY70tup0tGaXs+DzRKSLB6syt/y9053k5sw1xG6bNm00t+s/F2ZNSiQegfnu
cm3UEgmOQsvUqGbo7za65pnKVtbNwEkOBdOwAR2ok7KBvAVHyIikbDfMAngmyXGgSnZRxYEP9Tws
p3kuOccfjZ4lKysVwO9nNsflMQc+YDFWiQrQTKvTgJdT12dP7LSy4YOwzev2N+gyVznHGNM3aQiz
EQL0s1V6b8fep66XevYJEeNQF5GqkSa21VMZqLruGsCKaZoX/CM2Fdy5NH/YVEV2HV/5a4pH5P6n
whpAGk2CB158SI28HN5SjQTKe7/ewnaNgmlIucikXvAszgd2+Ho+fZYEvOkOBau8kF0bxVvDX62C
R3IsOW8XU6GL9+Sq/o7/28fU0PhTWFESySeBCweMUJVr8p3GRezjO0lAKL4BAjmieq8C6cHFfRKZ
SkoCDtjC6XjcDagkob1ZFEfsjhNe6svhJXVFPP8E/n2CaVZ9RCN4TxJfmzhaPwz9EDL6VSQjntrd
LGN+tND2sv0KtUCThPgEhI4MiotD/7hkIPlkzGY97Y8iEUMh4K8Qap29hUGRsJoyGzi1SfIMBEB8
nXn7wNri+Y0oMIPSI/W1PHvFKXNs8knUlMketyCUiH018KdnZifYhm+iOcXoFWy58pZIeLdP+XGl
60Tc7A4mWGjheIGAwZYWt+fBj0/RQCKAiFUvC+WxRgknIgUXq82mSL8Jg+SePAPtRpvoeQDBpgQi
piJwEJkQLOaR4sdeIHnulsGkkkogHAtionhghcOtON2kLZqifcAMZiGZYI/CegiIwbyuv1vcb77i
5lCAY5QLldZb+4/6DE3Xq7PPX1Qw/ntljxD+wc7uY7WAQUn1D2d+0Z3a3bKFcdokRjeII7TYgjTW
VnNRRR1owp8lmBK7r5hShmZL3j/wFL+q/5VJBxGyM9wU+nGqhbWrqfw29cjP32BUz0BGyOQJf/Le
jh0+O9RqrfMDvLTChl4M6HGjR/FsiaJJRl2Jkd0bTZRHeksVCrX1+oN1Z1+v5Euh0HKPSUkfhl7A
HEkzlVgAIJW8KUGS8keqA76acHtMxPr4f7TOu+k7T32BdKFptneSl7XG+UxjMGSqmNmM6aXg4Jsd
Ry5wHkAOY4WlfxAOEZUu4cIyJOh9oJ/3ptjPKDfkcvPlI6BLca8mle0m9mKQJcZdPeQvY1tudWnW
rY4xmBbmA4wveL4ZAkB08h2wqGJHGBMRZGluhQV6mEuFvMObxC1/74HPXFp5ynSrcVjnjLXa1K8O
lqbk90YfhGKuOCIubC8KkpwsDxrcRLDfa0YRwiP7oCAxIp/1V/gpLkcj0xisswm2+P63Hmw89ip+
eJAB5KssSCTlseqYNf0vZlG5apqsl8qmPp0fv92Rd+te3wLUG1rrlO/QEpU2z6liDp3ugxXt9PZ7
Y14V66cPbNRH0GDt3e9lkJsUiHWkkGIwBF+QshmimWdNrOsVqCog0uPofKJjYzZARlgYIMeBsdJQ
Ns0ZdtJWph4TAf6EenKRUCMNGgtv0SLHCoNr64RPzkqNd9cqt7erFOZKQ43Cmj+I/fnRqUnMHCbF
cdw6cKwLtx7K50wdi/TKdeO6+koX4pIs7gcm5t1IbDvuvTI3K3Lt6wHov8dOY1lVBIwD+yFeU9xL
uEXdyC/xulhq/rhNiZPjlQXzfc0DPFG2HeBy/78ucOz8+uDOO9/Hw3+SB4bxE84gUuve18V9jbaR
SLBMUfYTZP+MVnuTiqk4dhjp37mI0tsGrWuQYjxzUBcZiBF6cT706TEB9yI91YkFY7ZROnLhb4Y1
519979//nZeSoccrijKAqoZQ162GOUvWmIXhvvw6MTWtn8RVBIbqm5Ua/gl2eUq4B3F05I/n8l1n
MTQDAf89v4CZQKLxwxVixx/q1RaNxDP9PN9jai19gfMEHkqiIO3MbV4V+/Oq1j6azeqvUNuLbUzE
RVtZOPxcchk7aea4PuF26rgiX0TUdqsrxjeWgOwyjrdwC6ctralGMf+8lIuO/gSB7n284y2P8AKB
9FjdpBD717OmTIwAf1btXJs4K7gWAOIUO6UlOUy/pZ2XYUrh+hkoMUcJDS/cqHYVMOZ5X39QV3of
JI2GK6nOTkybrCRsfEvPAVz+Pu7AyPtPudppKDc6e94SL5TZnPWvF84OUUMO3M7REv2Vt16F7UsA
gHYFi4kf8rKOrSupf1bHPDU8CTWgGsF39lCPKR0sdlS2BxFsiCtYViqjX+WlfHl64RRFjuF/Jkp5
Rx/lFyqvyXqZ6yCcCalABXHIaElc8Nja4P2L9V+W3dgQJbiVBf/Bw6wWjCe4nsTunE8Gkl9bsTRJ
rreUmcCGQ50kRK5hFwDZzzoXHpWQgFxs9yrfkzJekOpJY2K9Dd1Tb7g/EgnSk41ngPK44I0Xo1hm
sqO5DELh5Dol57ui7jMKf9qZPgKPGxaEzXn/GiBkhAtue93T3/E16AOqR8qddCAy+wPxidgtwnx3
pJmqvoAjKCCGvq1uZ4vgDqnvLyiSiQzAlzFGnQddsyIfSxGG/p3SceI+sXLSjBWDMp5QVramaJS5
UzBSfO2h3GKlDRjAGJBypupWbdiIi3j3Qzlg6fZQgneOMNFBRSE0Za6Y4GxCxulWjQlTaqj4x2PR
05ycBf4q27EHmSY+Fp7/uJxJoqvq2DcUQsghm1FzL1diI584rptfu7amos3WJEbTlkBYkTHR0UM3
ebv1zHsHfEvusKIUBon5PphXcyLoiOzvLO5ffBdR9MYiU3MaY9BlKWa1LWVwlAJhKnvWa4Ey8xqP
xslWtxYbPoqlDhb0Aog3z981054ZgBy+l5+v2jZO0zTEPa8zmgFn+3T20M8SVwlvztnCQNOl9ORA
Yzl8FmpwYafpUcntm+wTF4t4BNrUlJD0mnv8X7dZlAMPL0S2KqHkIiS1tp9n05LoxTSECtk6Zuz5
jUrMXkKiBaZxCS5m5EF18isZKGUGXwoZvObVHKf78d4HAFB0fSrz/cPOv29NWwfFkLSgBfGIEEbT
Bch95Q+uM1w6kDSCLu6YysJHNueL1loQuCF20x2hwMc8IJkm3XfkAFWWY7Fks1cd6jA7l3ZrPQzI
XkjItpxPCxg4Z6ZWSqPH5eaYa+Ee9Fkbr2hnrJZce1gEcoZuFCPRxQ3i3/InlIwdxPGh9UcHcNak
3HBEwMqMpTFy4TMW6ifd1610TF2i/qkqC62QO0Djq13OM4TE9Atgp+zF6yMJ4nSwP7LRGni/a1TA
zQ52GNLF41zD3Ads7wbdEsj3aL4oblea3kCDUEVFpZC1YLPnpfGVCgSlVAfSzeylZj96ZmQgE396
1p4v1BStpcLlsh+FGk4NyAUNJ/lnhaE9kLxQwzAsPDhH5ttwnZ6px8pIX5i3Fy41e0calv7ugR0p
wV9iLEyX+ACX5lTHMYftDUiOPek8PbKEBgf8lrq0MblQGjh5kcoy8cy3fMCvAMirqpGdAuVuG3ut
enA04YdHFEQ7qLXNKjevY+WCVCDAp3jrXH/lze1X0GyV2huSCytCLIPbeC8toNlOfZiaOiYX2frP
umrcp/f9XjF5URMD4NOQ7lDIb7Nmi4d9evc6Q+dVU7odoBaP05DrxQwPxqIBvs2Sx46WwtfNu00V
8qg+yiFcbJ6B4fdzP1v6l35JYn2NnewEgvZo3Htjndsq8JLGG+V/AHzhKjFf7W5j1x0RE+zOvHPE
mM/o3r6zc26aYtOxT+XeVjAti+4etxVXI1LdzAfGf8qzHEYB8rBjgWb/EvzA6SzpLBD3EnW6gdWI
eC78MN6gO6AHziMThm3a7JIvACK6Iu4um8TSz5BT+yCMThcymTdno5SWAQIEk4Dxfw/iMgG21TMx
yTzQhkvLz9vnh3BSSCUzt7tcS5DdDvVBFvcsThjdwCZAISvoxdyHN3rKio0BXWNJEvIqefK5F/rC
pFgtdqTuLnhNBylx5vtqYyjJzwZkIak/QRuG791+mJ1B9jrnIDzbubXhy3zClWah4D48ZlUl93+l
8hDCg98JK6yG4AEAyhdyOp9NOJQGiuEa2LYpHI73wBKdr5lOb1DkdtIdAt3FA12Y3Q+EZREEA4jG
VePSt+wzxrnjcHUulruRrEpERpuNVyy+T91IqckrCcxRGAvWDvgl//89swW2u9qEwoG409jCW/8S
QG8gfHzOUKUEWGsRSa6SczroFAvZ+PImg2ODjjZwcy+XRYh/2SVa8cVb3BVCrWWijO94Ik+wTAbG
crvEqMNt7M8k1tkaCIYHgrpDyKjJGoSwqbBWkOwp/4tQm7t6yzk4wwCnuxrYMSEvgRRlU/okdZz8
jBP7N+K/d0LkpVjvE9X/FWPFekZq3Kg5+kilhRKFRS3G3lx+v94hq1ZpzOPJiwNw81ntkei7jeLX
fIRxWfh9iMCiQiqEE4v3MCIDbEjjCRtftBtnN75YtTxjCHID5RrZ61USBVSg8ApoIzeqaKKJEYtu
3HdfJRc8uwDYVRsCWX0NOeR/RHUTmqi8lalL0ppmme9RATN90q17XHsb8l/06rs6xapWjZqrit+t
9vzIcOIvqk5Y3u23L0l+uQKX4JTLJrsGfL5UyzS3j3i1sd6SPts2E8hZPGzT2ubtDU3dzqk2GxBL
Yv1483NXUKZNDbYbLfXeSfz2rG+looF/RIMs8KwoMp6naEWvt9mKd+jOv7xL8Js4ZB1R77St7QML
1Zd7bo9fJuJTp4F8A7uPIeB4do8B7IR6E6bGkVXOCAliefFfoSOZkjc+H7pI7gL3RywrhqXDwfSF
P2EXz938H8FXoo/TDu0a4quW9894JewPgUECuu/RbIta+fIyXYHVV87bOZz5TjDTyVxZ7qQxqH8j
/y0L8vy26ERyky85CDZOIyx/dLVtrAfxBCz9MCjLQ71mHvT8K5hETLV3fOpqpaZUe1FuH37C2evL
Rbq1tLObwSIPvkghR3YihBrQFI2cluThtaDMAn1U2iEy2F+CPPpC8xSk9Yp5zaPQNtOeZZll2nmZ
CGnjUiPDL5oB7viuXL2SO5shJeE3QQ2/k+BFuQhCV0O5cP+LBSGrA4Cv72Zwi25kdRfBZ3ZTVv/P
Nux9cvEdjeg7I/QQh9gsRkijwVFOqD6wA7sf+JV982+h8pnvTvY8+RJlj17hu1b3f72kN1Ing2eG
Iw1NwelWCys6NiufNfjPO8kfGrIkjqPlSPSHg1cTYnLQWxHGNQqJor8xFqwRlf67k9ag8F+ZGozl
7rKTOU0WKAEiVBR6hUVZ/KcqBm4QKcEHRLvMXIAFQm0SuiHJoAmmtHhUDpzWgLEcKxhEt6vTvEzr
4xi6AVPAAoGqlqwzljFoM8BGCSyJY+47pducW5zwZq187JxDEoXTpyX/gME+4HtnaEH/Yu5B0V5W
6jqOzDGL7WRpbwmewqnu6O/+FnJ03wPIXbJuOOspMk/nrRp8sCFsulDbm+y2WT9Y8FnbUaKup/en
+qlgrGbqGwVroOFq6eCNsmjZYQkpogGnvnYw4xKkkosABZtsdJ7F83z8cAPSZIXUOu2HDcapDg5q
LYjb4FCrOl+lJkYw4ppIIlIBBIj9lZOpuSwsFgXXowWULE4Zni0hhrcg5SjqKnJAFW4mTFsj5a4H
084Whv+0MKn8wFxu6zuT5Vq0RNyq8ncr5ahRX1yLf8Aq6YJ26+tigS/JYn2AhpzxnFmwgE6zjCfx
yrOOYeM6XqlGEC/aRdNh0O/2PisXtr2x6xLluxqmdTbpW0rFMcmo0mm48a5WMba8H993dFnj0Nfh
3cZLUjHN1dEPgq1bQk7Wlso/OcZoP4CbKDl/lYZEtSb5VQeosKL5JZw0ZfjytpxRtRXi7v+1Tl3i
z/KsQOqQs6fAAHB2WrIHoxrqU02EKp+INT7f78zKvRi9zuXM0iVAW+u6ZxsAkgvzue9pMp/SzJJh
HmKgZH3MX9omRSQM0wc+143GxMkEFAttgPWDk3UlV2MerFdXrZy4MAH3nudzoU29tefjKi38LJuw
XGY0F0TdYvJe86uvB1ZJSMNBpkPriO8o+JXQHJY0WwRgbcpE2nDQv/RDS3VFLru2xNw4QgLfmE2X
3hCa7AAIBwfQjO3ImQbcZ3CZoYYpBP2Z31QDAhoAun/UinviTOQvbc7WT9KI0zd8KiiZrU7SIasZ
g61Dpkh+4JA3ize4YF1cJJ3ICGz5nRvAP5UifGLf1J/Cba/3plgZWqowvKOVIzg5hKnYZ3ajIrEW
PCWixR0Mg/qo2oREMKICSemzyuhpnVTBIRXp+z0/IIsCyD4bd4ywePcgdEnTASXz0VcGGVEn/kt5
riVx2uhCz+qCQTqvE31Mkz7XLPt1Zq3H3qn7pEv1duR61YLx46+Atg0cmQ+in62Ob6Rf4HFmmss/
H3TiZ/1iQTA/Boh2lNLJWERY3nO9WIG2YWUxrCqGGLCUqmMurpIGq7lixLeu15NRM5JCTe3vd53N
xFoT2LHZzSV2nXrtAUavFLOufbqY0xPo11zoEd3yxmyuHlALvw8XGFnmN8tgwqSD6TjmUMR6KRQS
BiXc1/dLEzWfyYSsHK7Ti+YzpDsk2jkwYLEJeTuagNugtnaUtD/TvgCHjHclwnMnXYS/SwntlhdV
MlonK0lLD79y0tVrMcoPLc+b6vx2cDNjYFuCjGc62T4BuDnUebmk17Cji4Bire/RdzFmX/mAlRub
Mmo7TZ1u9bI+D4f5QYlYLs932W0ShduJPCynUnsANYn53vfNGiOEdHL1cgAyxQADFxmdRxC0meuQ
yGR1fY9qWi7Vunm7KIoh6zdItKGq6RH/oMHSHNVGXKC3G2OFn4jx3U1Eobr7FMUR48b8aYB7NrDR
bOOkbIL4RvPYTT1bcS4O085mdZVTqdW4SFpeHZ6CeyZHx8LH/poNFQ3e+g1rrjYKVNBjHMJj+ktw
XnH1ovC2uDz4o/3Z8tgR/X5mEwaZtbdgjpb40z/cAm0EB/GkPu16hS2u1sfsrervLE1LC6C+Bybv
DVH2zx3YlV5XFFUp4s3rEpMijY5Zlo62T1hKzG35dSC6PbDKY1JiEUSl7P9Ja2/ak2DhHfNAZeao
CA3xa5OpsUujovpjk3doEyndk5BzpVXZXmJqjKKJZm0hgbRPT4/pjTXOg7jy1gdSBsdZUeEJoHWp
1VBAhb5yiLNmmojm+7OAqJ0R7v0lDRUV7RqicgZrEu40xMoCbPeJB6/NTye5P0pQdQxODfEic2ZE
fpxwQZ/pmVyi4aQKqsMn39NkwGTfxvwig6Z9W9tW26diq6CZ6VkjLzZRLHtCe9872GLkD71R8cQx
YtUxtnKts6vm+MlO3ypUMszV8M2mCWHRmUQsKl1MSur+5Zr5y9IfonS3JCUl6ZMKy+JP/XIBAhF2
77UxsVGNDJNkQJ9LLD6d1O6bPocnLoqy3NucDcWZPG72zjzDc66uWtEFBxpacaGCqbo3WIt0FSqo
Z6jN+1J1CdSU7u5Fl+EsVRCvMxICXEsEShNUXekFuUnYSNmXyZ2IXPMsqgyMfNrQv7lrFvDgDJGZ
5RxtphQV9xPD+y6ojPmWMNwEwII/HqIWRVkXlvcG5Ok+1QcTIuLvXK28OsPvJlk1IIPQATzJfy6p
ljUhsKrXEMTZEvuzjkPL2b2uOdNWyi4poylcBlZeAGGdXjKflci0k2YxRz1f88VMoMxPEl/cF+Br
dI7Xu7tZ0gJRB/RXn0gRnXT2NANFGaqw3y+MmJlHHLjzPD4ZIl45P5i0YxLAImrrXNZlxCiSmhKz
m9wD7LoD/dSne7f9Ai1RBkA3FfzYL1O6SS4Hmu8rZGbcmhCXHkG93XCVibeW0a/g1DLrcTCDlNBk
6bwaEAehY3a77mCASnRMpJAGQW/5Gi30Xu07+FAsvVTNvmz17d0wBn2kLQyKgwvdAmNrQSqb2RXJ
CLrFmrNIRRCsZaq6Pc63Ua6muYNkXTOCUqg25xvMR02zFOAV8G9ielpjIsaATAf+Vv+6zSSNMqzr
2i65oLjWDDD2f+92RV7APKe4NdMCHk+XSg9IqNf1uWxzdqD+iI8GbZM4kG41SK8TAYrUx7yWzC6J
cBpz/T45VXgHeIlpw8oZ3v/wC3yJ/Gt3BUYL6C8SZ0bwIXU5j9i2s95ACNZyMzX/bJq2mSojb6Gi
P+OyKvTQijmXXPIr8/a2UK3v1DGHVIHDXI03zWDItcC7LcVFYL6aoxA8S+OP0O2I9HBFIrfaTWHy
TA/XBc2XA8lKIR+83KT0nRxG+ur9d8bQXekxteXASfYSYQ1h13/3jqx9AZzqPn+G1aKuerdOOPaj
ZjSG45hhoJSVzJqjzyzXmD/hr3+GGIyHoB6+7a2BMWJ5ceUSyViO8Hkh8WJtC4LkOczffQ/ywIol
A7WkWZ4sCVOD1wd4jeQK1Kemoa3aI3kK1swToi+hLSTYZu+GQVC6A95cUG7XgbHu1bD1jTzywVih
vjjlRPPxWWvxBtrPX4LGTr4EuKDh7KKlAE+lBaxdrcOKN24N975bkXrjrAFK9RoLUCRvClPGMyMY
vnkEXIBzuY6RUtuywq2g4X8GHtHX1V52II7AHkDxmv/rfH1QgjUca3ryIdwCklyjndk91qpKGJHB
IcWpaFBOP3IeUqUbKWXG7ldexy3A5hjMMeruQfHM5jAuX1SPi4/4IbSCQ7YfbjRT835cZviXvCxf
UOq1W/Fj/hRaMSxctu8HHtxIZb/lKXzB0XK/UYl1uWUOedG61cBYn/rQCiSufl9VpdAZTaAzIYnd
nLQwjKaG3d/c1OZUmjyDdbCmJ1m3NDtUurBWSzsS4a3HtmxHnS7QoxgGqzQl8ObtQw9wxT7LpEAM
4f+cIaq/qXZmLuVslKDHzAAqa/FJFuW5zIqlNtILqPwRkwXIqqBTuFJ6f1p5nEoa2y26PPaEcfOi
rjaNnN9S2PnGjGxVqmkzc/B4dvhfCUpNDdqfNzUA1QS+yooHrJnwKQxfojK+SnqpMeeLjfIjtI+b
KnGmBtkrdZ9ChDgZeZxpTWx6knz72qyJ+kpcoAzSmCg4Zv21NMw8SAYZqOgpRCJArk6GMkmagy8f
9KPaxY5gpxIaobvIJ67mem1p5Sn5FIswn25+46y5uC4c2tR9bBfIZxylRyuQtgm+ez83pBsosIN2
Ac6VerwlJvUdB8PV2JWtHNEkaxiPafA4rGqO7mx+4A0fBCz6fm6wGcBvgN1kuU7qVFL89PpAmIAH
ZaNsQIAXrxx8WgiC1kE8G7RIyNLOKKuPGnHG1H9tf+HqQ2PzWBNWelTyuxfS4BLjqFNz/IzuayHh
G/zf3GFQ3+M3rXak8Q6bVdvgNJjlsRlSUrpONTmuvjLbtoFO/bgFUxnUb1zgPzHHfnef8AoN7rta
lUhPBGwNmhjzFqTT2GXtkbHFT0BOFVHNFC9ICx6jdi2DTVDWUNHKLwCvSjpJp2cmsgrY79fzuhn6
d5U92JKOTbRnjW3vMpPgKUel5gD7TI/MAEztmtKwwFa+IUQQvOCK6mqQ4r6xS0VgpAytE1pIciws
kiOIOlnfY1Rj/pkOvOeWPvyB/yN3Et7SfRCl/dS5waROctYFxi5Dl0YCn1/0dNTupIBjBbCtJE/D
oh62uUrPlcM0sBtuSfk8IC8i/4ESBH5oG/X9Oy3ZmGEHYds+2TJ9ccC6WoKNmPSxIhIhiFCF+QOI
MgWh/eqNg8ldkEUjwtd9Rac2Bs2ytdZTIqhfbSY1buwwek9hahnqNyy4z/YWuW/OUlbQcxAHCEY7
M3FXrtEUKZZyVzYJZtuapbhVoR/no8d7a8burgiy/K1nRkXkuJXw6X7Pky2VgCq9SjSAjcE/smCC
P4W/HgrvVlkVVWiWk2tuPBO/NYwk4aUaq6XnEts5h+rDXzYPD+EWEeHS9l8ZTa5R6N0xLDjWS1+J
r43WU/22ZCGsZ8N77F87rU/tqBBxbPUIMssfsIwA9tnWjxdlq6yfp3PQYy0Kcr/oho8SLrtjuzrx
zFc5g3G4A+3UHu8Lj1isLtzd3KbhToFrA/SPs98BB+U4kTjSpsYQL6IDA0TnCenFoveZo7GgPReF
wMpuI6V+q47WStJFctO8cyUTcPHDGpKbOdc4RJAJTu3pub+/W2pgyEgFIn0WGtsF3R6sr+5IKxhy
JONwBYIGVMcZSYUcjh3olM+OlZ4+2L0E6gx9m8PlVN48HubddjrhxNuwIpIq8FXx2pk8zoRqaaKZ
yE+UfGQqBVeTKjv2XNKXJvh8kQM+Ov46J7tw/wKNV68oN1zCIc42TcM7yKwgEhSxa8+tYqpSb04b
yo4ru8ExwRUH5000L+dftxUHh/9soSELFaaQ3+QIoMp3TyGeE5mNOpRL20DgxzvkXu5pvx0622ni
zVOkXftH/f/Vtrrk3GoiYThGbZnB/RywnNyUKXF4oGgG0r3KZCj6Inm4fKbu+mXfCwxvxfgVyDOZ
hDkcYlhJyWxqWljTCQOy/w7Bls2FwsDRwFdCuxF7qjNk0xDwWOgSooCWqRHBo7fAh2GGVmHHf2ng
0TDkGS1VmkFbe7ep8KvRIQB1tVbAJMtgRfSrG9BtGya/yyNkdC5DPbqFammpSQN/K9a10xewvEZP
VlV+Bc2j4Y9PHV5REyHL93t8MAQROyW+evSWhU9htrk0sCst9IUrFvnUy+A0h79yecerifNo4gP3
c5nH5Q4NjHfFWPMUU+3vwjzzM3JJ8Y7FrUUdIjMdH+Ha0WnexMPaZ7w9+IaA3kdIy5a4Z+1k/JJS
vWRzZLluz/u1Wemj4zcWScF1F3UU+RKMuQxdQWjxQoRdFFoWGlUhC6yBeC20j+LNifBq0RqTWvdu
q42V07z13O+MOz2GWjiB+hlh4M9UJ+wxwKzyenMT9LurNzv/oAHDOycoZcNEDvK2iV0E4nEV/mSA
Cc3sBjufKZq7moH9Q3RYWE3zdSSpJcU7khi0zIVotl3eRZp7QbKAK2OXpPvkhAu4n6UqFqluQVRv
00Qalv935ijasNiOLVfUWS5dc+hC4Rab2UZ4ddzYncgU+uJIIHIzo/X2yH1NBc7APU6afJ2rMatc
pJ+1bwvr+TPQGefq8QDvpBuXvimaIojK/HBYoZS8qGG10arRPkvwN7Hr6LNyeUhxS7o1V43oFU/9
VJTuAVwsJX5qlCefa+IAk8/xLyWG3j4Qs844CpK37SoWHGtPAwlG41034nuAROYswAy62IPRQaez
UBEK8hi6U2gZGA9BrdVDk+W5VXVehCaVn0RItUbxIyP8IKveUm05TzOxxl4j8FfoHnbdvtDmosIU
Q8Bf8WTgw+aNWRRoYznePIZ4Y5tUeoXRUy6MVDz0P9cZsZHOMfDVRP+EjvadSk+Mqz4jsMHOh2FW
8nimRbzTP0JlSu4lNUe8M+hJQtm+1pF1+kyJmF7j8PQjIeuiWYoL32VpFA9rLRFXqJi2hLrXQfbz
O/CQxoGK03ENW1tFUnxXyRWTD1shbRTKiha10WuOgWURH1dWNOj2bBo88DWE6kk/r3Fb0kVAhtRf
Oft+rB1sp64Xlkjj6zeGfRoGdA+62AQEVhY1lhkww2gDysJEul5jzkcvokkD5yRodnp+HpxLso19
YQFe/0zitRBHKVeM8tHP1CHJfx5f9a8Fti9H4OCX/zkud+Z4HPdZGTre3qQcyAoGIsUpgkSEFvuE
qOC5XQj5rX/P5sHrN2biosd+pfZcPicqjoo1FgHdsg8nrgtiJHZ4TMKbG7G2tZQ63XtJQC5pcPWe
TB5yFshSJ7YzBKFSSo6eyJKnF4W0vZtJDEPaZNeH9Zlrz7D5AcYz7UdoQzxb/xUCYVFjM+Q/ND1P
mPVN7RN3oAaCfmXmUP8b1iAU0EXe00WzLd/KBv6PgDpMzTyDvDxsuua2m0JmBep2onryngcND2bw
tLKMoRiqUtaqq00pU3osKh3/o8q6hcOpNaGXpqp5QLgx/Rkloja5UcRLSylfzUGpvVMi1hlw7vZQ
sXdZRRVlMsSDm2jrLyVWR1Ih6U3cSdhuEj7WE155LMLTSWdthjXFWsWUONrmNnCXz0x7yEOW0FQu
QskYfGRmLpShgaKiiApEgi67R40VIVKSoA8j69BbprPxew0lEntf507MzaiTlVK3VOe2tm02n8fY
eqsQcGcloZA3dSI28Agy9YyZGOeRQk09XfVqRfWjrZKuERBlM5kC6BifzfwS6SOvHqo7oPZycMzu
/KBvggLW2rAhqNpbkk3kVZiWfpbUdLVWJUIG0FkjBVDEKceRZHHxq7JAYl3Yskmyfq3XLNoHMroE
qGNZ10S5zCmacpX8TEwtCAjNG1zFt1wCts40dQxk8/RtcHiWnUHZn5IOORjlEwHHeB/ANl0v63Jp
/4lppbjjVG2hXXbuk+A6lgnTuvG+orqheoZxPEssc9PeOX2z3/vTSo73xoQbg2TegvSg0iw+sRYB
RH08Jokz1cr2iu4X4N2kUHDeR2KXAyfceejW4ufcjs+aPVi72If/HvPrLei1UxKIrNJQiF+D8kSw
RygQdlp2W4Tg3AvmNwVDITnCWT/Tuj9jO+pNE2NTCmbD0IBgc6W+0vzNDnB/A751JYTzypVIsa+U
oY/KJEG9Ti8KeM9OQrJ3/UzNXoXnOS2gMLJ+arJO0191UnO/2GKvDd63F8nEN2Yck+lRVpFgTZCp
a4gucpdkwNEKuqSOUkcHqtO59uO2b1ixSqDWZS4Vzd+Tbm01uiEOI0+9TN9s59elVDRCTkb1dA9d
51XSqRqTjD3dkkT902T8UeTKpJ0js36wU0JE7Fz/nX7c5OXrYh8dzR2CZFj8MGnm5087xoyHPXmT
YAId1CYBiBN/cSlsooIkuza0Z4I+GggnokplbSWAn1QQFVijpUNlnYQV6DdyNJOoqfMAUUibKq78
ocTvosJmCNWu9SDPhsmx6D1AlzrykjSMRD74xwAuM3GPGe+pXDrkUnmS2I1TsX92euFMIm2QyGwo
CmvrY60Zuc+wi00IUhvVVqHnDQwHR8LrdbeoCyxtDxe8V3G4qEb+oA8e6fGaTMwsS797K7mDQReV
iol7PFIY30+KGXvgq5JPobi3aldSKZv6zg8HdWhVRghka2JbTZegVtrDMYg0grJJfye2+FFrnGk5
FbDHC+tBU7d5vSoakdkUZSE7q5EArhN4HdDOieMZyi4hQCZhQKhzKKGmdSydlU7yIZtD2MH2Oy0m
+0cnUExF/z/yIMu8yaUHqTbreQCy4Jbwiz+IFCFEZDZ2T+KxtX3zhY/M/CPqMVoQAmuqXiJUJk4S
06jHtlgFa8U73lbnXkBGuOCqdMjqPhu+yk0/cskxi11cUeL0VVovGaGmHHL3mXTOUAlcGZMICnHB
LK4x/7QoyzHCSHcFV3jmMVvDG8dVog5J8fhllAMaDyEuZ46CjWARUYtds8fvHFueTPfB441XRjAy
qsxPjVEb7yVAQDaKfEbsBNw8fU3G6tPvmcB9cum0DalwnN726Dx8ayymHZTSZpp61B5+HUpjaWpb
Ms5G7nFAnrLJlR65vCwdZaipfxsgHKtXTzR1T1tlVLsBgNEqzEVUmNY/4hJRXR5Q/3PiUvjMTMY6
OO3ZGgSh240LIs3q9NJahGwAq0Q/TU/CHk2NVUzkE/Xjf2t2XjGdMCO9bNHbW6Q26Xab4btQWlMw
JqSh//D1O20brJxHP4i/sJqQTxIqPB//fjXQw6Uy7BKwRsgupUzNygsQEDpAb5VkiF+nZKEQnESi
ZlAErDWRKaVztN/PHRvQH4ILEK2rvX185Wuot94jcCAmWILbW1pDr39xJfPyJraTspR/t/e18gFF
VWyoRlEv88KCiDUbMI9qnlnVSuIJY/RM+7KklCLLTFWYwuwDWBDeJ3Wr238G5Pwk6aLEZr2EijEw
SOnRDBwggitkbEAG15c6RXUwTxgQmzwEqi4VTK+1E+AmN8NPuajHa9gIZ+BDMHqkDtCcgUdcVd0r
OpQdLYcMncvP16GeWUctnM2CaKU0FIdbaq1qCn3/CsDk3Vt+TwwFynLGxt8nBXGbCyhEu+vyeA9m
vegE05Rz79BeJbJBBaeIAnhMvwk7G/5eekq/TICnh62SSTZA9Q5eaAiiS28XBjW2jn+Q+lF2YfVb
P6Un9BROQia3rqSnBLIV0KQXyLkOHkpkk7VRb0Hcl9ZkKlTkoErEQMoy/s+hjLNTZFK6sgKiHk8z
BwV8Ymv3SCH5NhfvLFrJwogiPnJIKFFtRr/6o1MlIdnFnJDc99HzfIA38+LQhi4WekugGIdpV3Vp
dVR8nhJ7ui0t39WSfnilXVNEb2bKiYDDFC/kLXaPvLFCGX6BTDdMx3WU6I0ya73u8BKsU0r9QJsv
xwWMRCUMqeh/RhRkuETa7anWSLg2LrcHX4kChahUBRuy/tz6rUb56maXkpaOmAGITm5i9694RSF0
CSUEUjD+2U5bqSgdE3AFGpPfPbc0SFRz6DZYrb705bgkBqTxYe3mtgKgTp35h2/s9ujAwEZJBWOh
wINhk0LkqpLSzvGwyNIUuI3NbsZjKW83/8cxYEi+fTTyW3YBtJZbcMqP8ejhQr5Cxk9P9BV281GX
9BDpw1kuegPNaJ9sHVO+sIcQ+E45wrvREe/wnCrhJ0hNsiKBz/hn53lZUYcSSI3oGyckgQa6kPN9
z0RN+c4KqRmz6nVQiknkTLpN0vwDG6UfuZWr/nF1b1Acj05HpuFA8p5A+tkh1emZ79jBF82UvwUu
AhI4FDz4zpkr5TIRwsjZ5oFyii9NuphrrbLDYwGeGMPhrzVterPTNibakcaQP7Po//na9HJDDBxB
Ym6csYJlyT6qeEMyKzNQ3g8jWcS9fBZtUIWfSW2Mms0gOCOLO1gA5a9DH6ngh9xWDYDGjCtN/svD
1G1kqB9fyIvEtCvELCLbJUk/WugLPPHKZeYKNJfyQKGBZqPv+p8Vx421Z9bSTFnj+82rw29Z+x5W
FunKG65m857aDekPuEVbf8RpH6iQT6CwUwhQVoRGIfDbTo9BcbUNBM/mBqroZMW1VbXvsG8vJEYS
izEQhnbKadEzVIfV1Hld+HqDfDn2AI1k/A4EIAX3RPSXyn6tpNDXZUEKxBsjQwTtCIZQVhKN6E1O
w2uQf+BxMs30Y9vROlqeq+hQLskwPZrx8nEdTSRXYCvaLB46hpSKiN8U22cX/jHSDEvCKa+QAXi1
m/v3n7U6lGQMLTgTbDpJxJLEky3dRpvJaqP9r3Bn3L0sizNV0Fc8N2nBj2qlhpjW2qtusgs6HMZq
yxMXqWGzVnIeWdCLPxelwjWf26YIX9WEJky5Afk8p5yfVs3IlK4CRzx8HBn9kloJFvhvcIxmNmgR
io9gpczy2V81chXvlHoq9PQzgt9iZMi/x4LTz/I80jSQtU73P6HUeeOdU1UUwPYLWGfszv3TieaF
rJx91tYKNQ5yEBgDXFBKxst+SaSegPalYGnP2L94oZPaPog02Fx0qUXVMrFWA4iAgQgGlhmWpwaN
86vPM+4IysXHVVlYB3XN++VzLnNudjCbOlb8H0Fl+lxRhIdMske2JOXGVGGdxZojbq0vRA06rb3t
vXjKz0Nz951MnMEbGhNu2ylkKTF4/cxZub3drWp2CORrlTCEGS+dUxy1yjAvfbyZJI/VT1Sv9Vmn
Wl44rdIwXVphf933xawEuZ23wojjlXo6/p4mPaTY49sPZJIUsjZ/BjzhRgiCM30psYe2XL1zq8Uu
9UldfOUZhDnTi6MDwhULPQu/4aCu/fY9jqS6bEkiOhy8HMhSfsdTERDBUwI4enXfW+NyxQl9ilZC
DO61digXSNHPYQus5J5v5rPui9IH3kAt04p2OiQ8fXbkqv+o6Mf6kM0FBcE/zP4JFXXUPSi6H9IQ
/ga1m1gW7Y++lyPzW5ilAfNCahi5UK+mYoGBCY1LPTuAiTxR5TL4qbbSxQNqbn2n6GHt/JFHbge0
d+c+TUIn0jSauOxI74zFmGe8MmM0f1uTOItpdLjc3MhU7OGoNaHVJqUBIK1nVOQSkfQzqHGdWpCf
RBXS+bSG0D4Rs/Qz7V37+B7+jNh09XQ5dETpn8GatMt0CxBh0kuaFxNFiu3c1ZvUHHTc/bTZIzpZ
ctUZe1NeRbDY3bZ9de9W3SOLuOvxJ7l452YC9k7seKST0+qKvOI0DUQh4JOyj1MTYuHYdVpSm0Nw
WSKczZiYfVGhmW4VgC8EbQGeoOjG/pduhCdOKHwYGcTAvrJjsa75EPr3DQKxtgwUbbbvIV69y/Ty
9MGDXQaYDXKEi4aEhTlHmDlrz566bCQW39MsHb6+ZUsb3+HC1NpIzCZvwaaWY588rQDJn3Oes7gz
usF9efVk41avVIJ9Lt8/vYtoYoRaPDxTcD1MWFbECGTjzi6cyREtCv3kSd3EsNulKSmP1GLPxd8d
e1I3Yr6QyIIMCVHj7psXT5ckfsHNOaGJnYqr0/Owzog+6tVGAH+Rjl45u+XXRaK4YnFG2uXOPToB
PNwOuvVPw9gyOcV0a/wKN0WNbyR6Z9QFfacP9s4pqMh1ekJCpggmC2polVIcpyYQUOF/6NaOjOkC
em0m23HzBYg3u0dxg1hDvcmfKp/M55G5+45juWwjAdG/shIwuY6Wpy6gxQtMrzW7GB//j/jzzhAZ
k0ZFzMTlW62rUt19Tlo8AlljlEfuo+uEjp+7qhDz25ImU+r3WjyxB8WiQyKMVdOIMo+pccTwfnpt
2RMQAtk0uzWtWBRnz/lhmnRKQsGt8LX1JlXIdKBQ8fzCnHo+wkiicd96eDs4bf+vf2rBKkuk5zvY
XTklffYDNac//NwwHEYotoXLn33XUXho/wqpuhNpAQnLVOx2dkqJpd9eYI5VIGwv5XSdrCpQrxq8
J+lJxb40B6sx3Qu2HQ1eTmmJHiZXKq4DJfj3TzmL/cNZ52FG+J2kvn7jUdMhfhtLRMl4OhWiotq2
TpXwjqhDNf5ek30ClANZL+T/n6uECQrKUfZkfT12dJXupKBArBXNKqq2R6H2PTmh8FhDbZBLEaqS
Uxx0UVN1NVa8zxiJEpt6yLkzf86cm5Dr8JdI3oCSVkrTTiKOyyqBSMDMmSe/t3JKoif3/kokWLsM
jz6dWpmQWZc0GDvsX+C0i9UZyQ2K9XleDvZHsD37hcZvbV9a46iuqZjSDgPVPmf8gO02fEpd3TJP
qCOTyZ2yGYDfabwq+eUr9g8jYspaIU4E0w3IkH+OCE0sT3SUST9GdWz0egBj1yHZr/zNlIQXKDQQ
Bx21VkMd3i7+odR2NzhNdfHZpZNaMbgzH+YocBDJZf7anUDgFLkc63do00mLZxjxozEoTdR4zxAG
CwN0lodIA9lcjB6IW7kxT3x47QJE3FR+hTzxvLkDgMIwU093X4LBAH+X4Xnk8U76162m+61a5Owf
XwJgzMibd8ek+4MnOaNyN89ad4EntZLuiGkoJjSbvd2WRVL8UmUnXpzT2u4AC4A940FQhayODW6K
dH90kju8Yx5ahivYOLTP2eHzurLSSyAV2kX7KeoMwoSZbvDZZv4roNMO3dViCCQTctoYOU71oRoS
NguUbHm2mVAAnZC+sAsHxHE2sCnjNdkfvTAcv2zxTa9nIZ/BYGIvzupXQOxdz2clTUsrLMMIo94n
RvaG+nlBcZrHjI1tf45Ud82XhLDK8RVRVH49pA886+NDmDicpu9sFUQuPB0RQ0MRSm66vB9Tm7+9
W/8QRbPY4j+mBXlPyKfiiLTv+3eRYEN7br4ncyWQ9lxexXe2kUXWobATSu1N9uQqb8eEThO7meZQ
tvEPz9YaoI4qHV/6pRzGB22kvTSbxZgIm2EDz+kXNTNWuv+GSqa9kcNhpUlgI24MIXCP69FVyUC/
lua2OhYR7UgS8xnQMoOyOqKb4ijsy9pL7zB0WuZsd3ywrrtvQXVVXt9gCWL4Z/vJW4WeqAD1z/Hp
Vp3jaADQ+VDgVS8oZCa/3wNeBbD7t1UQYaHGCXgR/WOmPQ2Gr+bYXrJ9oceq0LECZmk0WXbSS4kk
eAnF2TyPAylU7hsd2h2VPSK8XkoCWRZSGGeww5wkHR/gu3Aw7XXkBlWlfGedU/3bmj9PrsoB/GJ0
cLm2AuCKeOWf8yiBDLCRUGnEl8/ZUFlWe2BTMOE61QdbJlj/Y+dCRsPNJs6YZhJ+6lZxjbW+awOl
RPWC4Kajqpy0LjtQQlAbcTZDnNJ4EZjcIKGrtdqkc6BChjhzSacdyLQbeJycKxczzJlL4PqGvkJ/
pgk9BziCf1aFcnWZBPTW+vvPTGRpwpfkfizS2mD9YLi0ISekz5AYNaRSgcfWRx4m9H4zpWczRyGq
Q8zFYQHfJ/hwlD9nfLH4h0iVNGOxvGqRmBHuk5/FxVpiAWfAwq2JAIPH/5IepDrs6XxgEm8caqQR
3MsDktiNiDR3pKU5OHPziLAFVY7K2pcc6ONCXh/XHIiZUsIBWxqTyOSMsLqmO36OTWxc6Dem9fp+
DhxfVnMmkKfL8pduHU2wHj9ltYyuj4z4ZLylrTmnsbvLeqUleL5PEhkTsdJ4K7fpesZ5xIrT2XB5
2YF/KV44Vn5mLQG2SUrxnG7YfFWPHUVb9Kqc7Nj9i/ny+M41PGOrs25aW70c89LNTIdPXeK1/4/Z
QYG5h3uptDA6exWJtRP/W3zh6taJde95BfLx8c8VahXWUuZsZsod+zONEvOUyAcTSuguNNGFXhAV
4UqkMLF0WdhtsUI1IkBk0iXXMTnDGdrC7N0WOBhRsGBjPIDSztgCHUUGlcpLf97cT1za9p0FlQX5
w0dnHnjkLPHWgDYxQjeWqhGlbkhGQeK/Kdty61KsfuQA06AvMKXJEH+d69SDwrO+HnRfoEuUcFkA
4J9p9WQAbRmgPEsLSWBYrS01JoyFmxxlbsUEdMQXfBYbnZvmRUJKeZRT4UPPgZFIUig+/QiI9kpj
87Woygh4eOb3gRK2MK+ijJGNt/yH2p4gdjaG2N54DBWyOn7oXqmsVCwOQVMMSpZBxhFcS3cLi4ug
6Kt1dUkY5Mm1gUBabbRltdKTWmxuMpTwIuLbZCn3luUGana6jqdItj0wYXW4wVjWhlwDR4NK1mnM
Cp0ScS8IrITJpa+w0+QeDO1pEnviW4nDWxi55lOHB0/tGh4IqrAhJ9SgO86vtT8uJjmxahOoIvNq
GsLwpRD9hX0OOz99cl+kCosR1FJzGKd6On/uq4ovy3gFOU56RyhExGQ+7Wjt3F/hOwOmoTxNnjUx
PSXhQsIM3JhQ4r1cwWdkOQDdbdCdNXo9W236/WJGhF64frghom0AaZtyULk3BqvsGU/7/D2LqfJM
oe5loNfuWjDMC1iQyikJfeMOM/UaW89wwmWT0JV55ipbLE2yxurn0fukfSxv8me9DM2/NKLrVW5+
JGfzhsxBYbziw7JEmJ6jxpqRLFkQargq7ty2bNICsLubVDveO5b2yoZVy6uMh3b/9dM1x897b8bm
6Oroobcojs/sdivBoqBvpcbt5JNLVYgPps8yAIfRtUFfL+ZWvfo7SX3OU2IGNi0o52AXotgNSRem
Rgzc2IRDyiYkJ6WilFecXm9CjOMarndH5MUMnS9WR1YKwnFtxZCLxZDb/fBKloYpOKwZYyJ4Y8HI
yqnNvavUM1Cd0hzsYiK6q2UEwdwOAe8d6tiq8LFjT7TENZQXAIeUW0PPIFpq1PqNm2AVE+ndkdDl
mhvroJ5itEI4CjYdT3sGO0QX/V5ECb1qsBgdb/Egt83jqS3E2ghgmZHL1GSCk5VRKEXDKLpCxsgl
CWs6TqmLB3D1j1FzqXSaQ4PVpASU2EGFbTmJ6JCv7hB0EpRYjGcqegrCMYzB0U4/vHeLIyZzgkIg
DYg5feW9g70d872pHC8YsTq/4OzDEk+gPKtDCCKwW72gcXDwZM098u14hz2G3pDoLt/vtm+tC76K
AIOevSdAVF4FfZkZRUrlapdFRbInTxIBcdQknzll8kjwRIDG8+iE+kjbFsHtHWPa3A1p3gXIOmZP
rMm+AaHSAK+CLo4QlAPSEWF/u76zWZik088kxqAY6GYdPVDwuCdXTHH/S2ZMp1SGuaMwFohUuEcI
Ehc2tRP4A5sL73SL0Y7t28eV9eFIzQmzjh+lo/LQpseHjN4bx4sO2dhutc7Ci03zMXUA4CcvzSNP
jDenNjN6/2a0GYQ53HJciTDeV2MGoEOvrPxk2xUJ2sfnuebkSaKprEodRv5lYFftLuWS+0LQuZ9b
tqO3/E3w1+NE+tYI9lzClfLv6OJr5Oa2I6GBWqAOTocBmwQNT9o5brE+ZndGR7ExuiB5q+QYsYSp
IoE4sQP6aBNVHFVW1wyJqz5VekeoA67AikkQgbn/cSV+aWW2itOx/sZRbIh0vLGKiAf9WQQ+F18c
BDiCRjFQ3sDOLP9Zz3JkO6iizqhGRRpW78WpL9ws83piG14HlbCWgiA+VDEoAWffUQnsAjmiCKPU
/k6xTJlAQzoYqWkdYhYwshIP9ScQAs0ys2vSKqCVnC1IPWS5d4V488en5yzAEopHw9HxrkPRtnhO
u2JYcoGeLe5pxFpXVcqIeVTTs8vSNqtWe/V4AMa9GheBjHefIT+9RoIcubCobbW27qZ+EExOYCYA
Fy628Z/TrCUA59Uo2pUABi4gos3X3u2nHPfN2RX+efooi+JYVFakRXUApOvSn+NSPHSg7tOh4irs
Joi3/kGu1c+PP+vYiWWwMVzLj+GVcHqwpsZjiY5WYysCWEwpCczTAW9Vw62z34pFFpHDF0qZe+Ur
jTwNakEDQxKbMtfyzOf1KmA47hBAQE/c1CiyTu9a2uU+WNXD5UNtLyDSu7hLHkjiGxWDT03YzBuB
YwpZsHX8+lBFW1TrOaRH7eUbnihbkVVofBxFvzajYIjmTpUBNibuNp/BotMYGRxfVO8+8RlaIUNK
FN9d/meKA9aFbPtdi08WP7RvMtlBLFgLpSDsNQrHWOK30biD1NiHbPS6q+maaKaLfM0OGTCFanmr
j1+Lkq2jwli5E/YTW3NAYK2q4bBZxvo6NWoYlMiH/ri8yNZHb6G43GQ10Q8I/LYOJJscQQX6lK/r
OMleytTChORFL1i6Bu7cH16nx/m0Cdzfyfe7lfwCcR/tdtH9BL4++5VneyXHrxlGUSzcf9HfaClK
Swb7U9X8QQLQBt6jlTLKY3sJ75L+JEyJ5ONMbTQGiwDqzJLjjho3/CKFcjx06fOKrCUngcoaRclj
7f8sBNMQvYzKi71FUuS8BgQp6i0bsTWoBX2EXPM0P59IhJjC6R0BoC1MaQEklOCezTk3yw7YuwWD
H02JZMRVUbino/pjX0mkCY6btdSaMcCBi5Li+9ken+fvJmOii9MNeF8gOVuaV+lAuQVOoNNfJ3JW
8lClasG8NWBdJCTjpZ7/P8zOvFi1LMHbyXq3UtvQqPeTUSayXUOygSEbfuSOBsv+iK+08n5FXubE
/fsTMPfGgWMGLy7lhMx+FxFofkG13ab5Xm00pr36ADMynMVKjifn6HVwS+w48kSn43MH4b/aZGRT
+b6NUEPAVPMYxfwwceKY7unnAXExzOkb9qgX7++5iJ0BEjp1nY5fJrmQPUVpdliRqlkpjp0LtcN0
aWOU6Cta/F0fQe7kioocuYlvdSCA5X5z8WJexHai7kwLdWmhBJ6pJB+KG38a2baOpnTX/HzfofUI
NUVwFZ8kEEH0cUTVIiSmwE7gFRkma+PkJPjZ8wZBu6NS26T3X/djhdC0ddYY3/cQ85xZVWrrMZfv
reMWO75nUQpkVwGKGv347gb9JXEXx4DOx0DQJtwwsa7Od4EmKSWarsVieOdowZzN8gnokvR6fBMC
aaY0qInKJnoobcpKi3mukjhKwVF6ScYszCug8MFfqrlcUwGzjksTMjRu+5wlYGrVu2Km86a5uG7a
gEM0NAugid8s6ruC5BrJZkzORbzde7VjyapOKgZ6LKD1gXI3LrfEQYsIPDBgLhFjftLVeLFo1ujQ
oBvw4SDDzrBVn+6FKvRfiiPDVIbcIk8CNYxviDi4RCu2H/ndMh7o7Ae5denaJv+eDUFrvrH0W6/Q
SrTX5pSrIx2VSdncBoLC/sO4ovG8yDs5df/C8682kCEBYLg+//1G6XRLNRJsCUq+7mSkXRTzceCM
myg9q0aUu+6h7974cgZbIvsl1I8VfDxAS1yiR2d4U8JjotLSg11zcEA+NeAxOa6Rk3663cFMkknU
Rys8srbm+kWXIgJf+/AalbytgzmiGr5hUhPBHDeBjcH4uPz9CICm70jvdswRk/ZvJvyW9zDJme5F
PTGeCciAR+k7dfgUXH3Kx10sSQLcKmymtXPuDYhV+8UutFE0fITgqBu7ZvGGiotzGbO8lQgHFA7E
4eLKaXTYbmdK2fy1INtqvcv/kxVRh11OGO/G2Ce7kH/NVHv0hlZbj+KWJ9nIaBdBLuTURSAD9ylm
bZHUFlFVTvPknuR75Pxe8LLNRgsgZGrfNY+uhjZ0XkS+l+/7aFYuJSIbWuoqpCY8URTG0BXpysaW
1XWNqhdKQI9++w+08LZlP+WdLwR5sqwlCQ0olRTmxaYafIsb958conxXqAJQ5UZfh0+YI1a9MolX
HcCZ+ugPcueSw4sgounUZp+Ama6Ff9ynGPsPbxSDslADDSyZ6cRgp93l0AlgRdD+ZT/QDnnp4wus
ahxbHTV/zm0U629D6OyLLusstXm8jdH3gj3sfPzIZzLlgpI71mFygsiXa0vPf0Od2RF/221vNZZI
4Vsod3ZvFoARkq2eXd81vjkJDtR7rovdCFJDXwPzDN4hnWciOiDJSnELkgwsFYqM0xEjuzjDtho0
DfOlo9hcjf3oc/7H6k0UAONV37Gqv1QKVsF+UwZJx3BKVR9Cdxts1cBAaIW4CielDfqH0LqKWGsc
dZIcIBI7Ed4SZPIH49CTstpNno0xvcZ6jGyi+ZDCVO8pBYX17+15UM/nPgTyuAwWwozagEi5/smY
bYrwIQE3idNcEt4Rxe43igoXiGgRtJ3JGBqdws7ueDshFT3V8uYnekVwklMEeRy46o7i/bADR359
yr26m5cfxz5bn4ubrvHTipwu0uZrBxL88goUSLC7ZkcUdzHowT7I/AvwjHt5b1Z/T1sfjs+6jdcl
Q2axvcpRGdCMD163qaiZIzuRbCr05iB3VsGm8bM8B4SHTM5YU8QK7QZA6k5ivxi+BWdJirVkygOs
Tywq0JszfE9LGdhvRKAU/oGbybMdgUe1zZB8PyFtRTPlngII4OmzSqSbHwRUt3DsFwFXOLqpy9eO
lDC7QlZuDpjgZa72XJc5bGk9fqI42owLgzjA1iYaeEWG9GF4AF4UA0+L6Ww/Xeyde837YYwXO96a
hLYXLXckZIhouIVIs8p8AJM4waVdkzwgeEegZO8fUk7L72r1w5lwyaEJS+A0YejHDAqyCwDsZeja
sfwceEeIEgnYZa+PGbnhCtyGlJiR7lJ0FlEvmLj5TNKM3EsxZbsvM6y04LgGw44tUzGq9nMRSxni
8fRWq+wOwIqxOZSoTJAAwbrj8IyYIG1NNRdIwLPGLkajtsC1v1+oI38WGbkKAQvN9EG+fRA9WnD9
RYOorXtjMM4AfJJRFeRUJnHil7asK8lDgQAZFZnwSa+ELiF+cmy6VEnuIZ4UneindIHoGwelSw8f
hHtmOO4IlNxWhL6dlRIy5ZOGabtp1MYcdSpWH7Tx7v9PR1Mit9AVJGj49HXEVXuU3AGhab/K4xAC
d0/OTUw7N5+M8nD/6f7MDXBxI/+vlkVSL6LEldj0GCxDong19oq4NiDa5ryHsfHIos1wvVsX7HVX
jbGYak9yw68ZKw36JinpcJeENlP27ZYNpHy+3DcaZz/M9K51KNeBvjqS8evhtyznytiw/z2n0AeO
22gjD9Ewu3WiOZgF65rWSwPw5f+3DUsMw0Ns0obLTPt2h/3rHLXTyJfIzaBhQ6NsQR4IOaIY7BQK
u6GSQLxz161ojGmGhTmllUPpvLvu5voiuIfL2DV+O6/Wz3rM76nW9WeXwi6rRvDkqOyUZ6uSXbox
WNZjNsErvGn3KJEnMHC4hXxmmsKPgmjKRnIRD2zRgxVtdMRQEZ/E/YHXuRxSCCpBMlNg7wuB0huZ
sQN0JdxFY/0rndyMaKNwuYJtHobR2NIO/9to5d0xAAwfiqYGESAVM1ypFSLZH/VHfPewX4WDhH4h
mmH88mY1i6nwJ0Ow9VDewwRSv1wUkm1xbtgpXN7SrD/Mf3EoQvXrqhNsR0mBtq/OKRvThutUC1ft
GGM/8Q8X+E4ZnNhtAlP1K/XAxjWkXEpol3v5y/I+jlhVRNvQPP2kTglM2wlbVxgvwdd4yKAdZBhi
qYw5rcV6JitefHgk4tMdx7V6uS57E+/wxBOnRNYjmlUOOgMQwKdf5jeg/nLKyg7N1zUzqn6wb8vH
QDtds0Y72Y95pTK57KDmJ0/FX0rC+J/fuLq0Ddvfl03JCuo5biL3vjZWBRGPbpYDidBxGirJeOSW
aRKHH4ie+VIcasgGVtkbrjN+XRq4Bt2n2CJHoY8o6Ym5KMGn81HY1s/3gwPv4ZuoiJhUhoEaGgBg
orBpUeqHwebmFwgyEMvvHccSxZKmQ3/jbYFuxZP5LVq/Gk0ZLA1qWtrM35vpu85Ss0vHv6o6WdBN
3XW8SwvhNBbJyh3uVBaFdG88JDZwutjGUCYIMvae8cmVrzw8rsscBk63mIa9P5Dd732GqscgQIjv
nfwi4rw0L27TLE+l8HK5XeGlhYpkuihUJaOaBVZ3F8iNM1YE81Uh5gOXycEnuHWK++CTFojZXztE
lDf85xyn6BurUQjAOr9ZgAv15bvzolICw9iXS6r9n7705OoEOkJx1Bg17DRj3pjy1HEty/JBviVQ
cDa20AQ28c/qexeHnEirHGs3igy0c8TsUp3BEWGZBMcl+kVrNTPwkur1mw7uffGlsgIKqjx/fPnP
xH+FsScNGv43SmLj0ojruoSSsENd/idDrQwv0gBi8A87I0w3IaDHuQ6lwmmci+vs1VgcVcsxHkxn
N0w079nNv3hPU1+XjEq0Eua9h3QOKSIKQne6J3ZDn8Y0YqNz5b94A+vaBsTpaT+vNWJxTDLmAnjv
ICVrywPqVvys0rws7HNiXOPxy4ptbF2HXfjwFd3bDRvvgWR1XPh/Pk1K2XJ1iKiqpyuo7/rC6pV2
3ZH2yu63S5bpADVV3Cmwj+B+Ss7gYjyO/oBuYuYjeabiV17elV9w81dQO3WotImBRPhWEe+gj2z0
8YUA4b+Z6SrYBW2fJ2S/WiB89iu267q21e8rDNLSUYpp/lAZS3aL46syy1iFGA1+iEwiRXV+2kJh
t6EXEEngANCWX3cfGjpXoljqIl5rsMEtwVxMvoeN1IPcmYfxLI4N2szu0nnLG3Ck3zLwLKGINlod
sOKKlMbt+fe0NJTI7ABEujJPDpL7OC31uwbH3iCVLPN7NyURc6UuRf7hBI16jlW2eGuaYzGebZEJ
WKsAGOqysqe7tHgBdZwxOCTwzc140EArrt7TsiAcfEpm6jqrH8xarHTzoRt9ijblsj6BUgqIsglr
7lPzo8xsDp2AGez9YcB6deRdQlBcl5PY3jBMGe4wxKAbmGuPC7SHGezQHCY4pa/Meqh3lMNV4deE
EzpCmpnV882lLFknOcSM2lbh/g8rP6zCaQ3p5VnJJzt56uWjoXB3DLxP7anR6hkN88ouOhL/Ypds
2dMpwp9rcmD/TJ9Tc2YjqHD4Y3cN5nNa80M48fO8Giz3D376eenbi+egkx0VMRL1iiEs7CF/YaL6
ERRC3CyyWGQLZb1yW080nv4JK+vcAQNMBxjGu/VoU5pEEtbBZ4X3IAv2pnsCHYsgqmuXLQXFyn2C
fgPQW3BUr/FAUJgLnOk6M2SN3OKmRHXepImsV47Es+NlbA93KN3eaH1zm7gb59z36cQlVsUl7AZt
nQaJbuPeAliUqkFTw3wz80c33I0dOf5xoiEMGk3gQFyVleZsqFmRsJA99spDNEvSY/YuYztcukYj
vNrq1zZuyraXTSCHsyRNfMXTp/RQEIl4hkbBd4ZCi9cFTUqbeW778ikmJfBc5vkCLtGbMaQpZDU4
0TXdiPRM2NFz/QFHmw5TGFdPvPL9KY47H8UDvzztWjFgti3rj8YteIWBxJ2yDdHVKYjQS2L7M7Px
gScyakSJ6tjgSF8ji9vXOtAnZ+tBwxTcI+HieC/bQvkT1FYAFBx1i5qJlxy1y7ecNCSQMJvVRQO6
eH0MbWWXVS3YMc5ThG3NKl1iHnoMYy49jxEi+QX2+asPBLNY99zHfsGqZUNpu6u6ygMVt3kkItEK
3rmf4PiHq3h0slfVyj4nLI2V/Tpq1Qhy/h2Ez01lW7i5xGJCJIXXfmAJXYN2N6cRw9z65aweNgeo
UkDEDD+d7gTMpTW6zfJqnzi2122AX1Vdp4ohnqZRmryYDrut/JZcuNQ2hZKF/dR/znELTNSv2bZZ
fH8wlrFDP8rv/5Ndi9N/MXtA7uEcDyPlldQdVxW+fRZs0cV4wVDxcsnRbEVRff1W7MvQSwvHgeo3
/RaOJuDbYL9RsVpakAKeCXikt7ZJjSpm3AVWnQZk8TB/ijvSZ13hV27q4jg7OAkgWhPHumRCyurD
q642DdYZRHMBILoppMPnj89B+T8TJwuZTR8W56eAIMV3TOMtBGDTNDdqhDzFHWcp5LVFvUNopEX7
cTQNAhFXpx/BP3DIEb9Gq48fvUzjhtONqYq0MH92Esw/b2jdoafpUfTxa+MkQcgxI3jbuduChT+w
QPKWokrqhXMAbG4bBQNP53A/WX2zMWdeCQkqidKW5puXvefx4V8H8csBW2iQ7LpbGM3S94P2e52e
d+EvzK8542I8Z+BEOU9CzDckw77XRa37AAecbEquGPkA/GRxoMk8ZpQabGa0xhrUKxAuf99p7C2s
HWgbUdWD7cNZfeePK8WIudeKddqT6I6Sv9irJEmwlm832Dk/NgdrIHI2ZtZ2A52ftBcUS6HSZGi/
Pkfurwlw7nO0dwxEPdd6X1ypGEmwvp6ccWP28JPLdLZ25NLKwa5ko5z7c18IbCJD51DNzAUSwy/j
kWHTZLWn5ZULhXHZBPyQZXRGMWxV+CVNpyJUBNxPPpcjGwrti++jdYw12wcsG3wKiZbg3uce5UyW
LysjDoNDf5u83uZ521YUvVv4IXw5z88iVCbi8nvaZ/bD8YLSHlM4SsLm2YMQXykg6hxf63r7ckMm
yojdzCgpYaX4hBawwRzfnB3x5rdM/1Hq7gbyhixg/SUz9ML9JJULfa994Tq1NhNd3ROZ2sn+RkVO
wx62Q4B3IzFhcq+YLDraI2r/ACfO8cEcGzMFtF7QbC/aqh7vAe78NtglbVU+D/7Xm504/PYyf5sP
aPj/e6wfUK3VA4xpXmXMHJ9HMs/dJghNKHDslJ/Yxsndgx+4pNCAUYTHDfcrLfo1lYXUuZz97abh
I7Up/XMlrA7H8D6tnTDNVXykgkdLAw4G2F8YlUNcqU9d4h3XuEVl3yPsTQupATP9suBujqsoE9Vb
/XXGpmUCySsgmYXTiscexT2cYD7naRMOtMzsGC6kGi3lI+3V2n9MefNx7YPdM106R/5ZL9i4t/Oq
ZUv2JHQk5IvHmLkknMbNVQDsK2ub7kBM278H9jJSDpJFT//aoj7oCnGO2a9glVCzz3sb3eJABjrS
XjpEIrw6RpDSK0BQG8yVDDdiHLUtNkj26UuBJOLmCHUpMx2LB+YpZSWYlnbanem8l31l6ETGSPhM
j0AmWXHXkLsJq7KUx0bOXWDo5N4potxCELG2+DAH0V937TadWn1kcsTZQX+41vZriDBfOaC46hAO
o8S2rs2hHAKXE/wMGEX94lr+747DO50CQotgY4pbih17Hnv/8ezOqlhekgJ6Qxg/NRSky7ICG3nF
g5CPY6NQBFd0550J71FydSX5C4ldYn8/RxN05T82yBA9DbQ+HGM88hXfEBTVeQEbVK4I9awk1XrQ
ORtR03gGuwCOFoEmhXczGeWWmOOdJR24StDWJMbgUF3zT+pTXEq8bBT+qMw4U8oh81ieNOTuWyHC
OHKKaZ1a94EuJgDSizKF9gwTH7CmbKVlgYq12rHGvuOmMklsN6UfnBSFzfJD7TxLho0juexxOVqd
SEzrF5AgNqmpE6p1Qa1i/VSrzSVkPh1lfWESzR+fsKa8Y151Ou4gqPYfxC3DcbG3oE6QRZODxQKK
ipNT1OjkU7PGD9JZyE6UAU+BL6Jq3FvSr/Wx8RkwOr3h3Yt/LtS00kloYNPAjR1qrkTjxikskYz8
A2hGhj4OMSLvTJaa70SGWoiupctv0kzuAoRpPV6WYd8QlpqqXOyQNckOFa4gD7+L2HKkOtL4VO4c
UjRei/0VyA2r412/EyWG0JDFrBzstlyGOP93IxrNAlvnZ89twGxsS01yChQqEV1lgwiMGZi/MEyt
ShdIcLjJcg+5GHz1A+BfqAQP/pao9meCnRU+K7pdxruWoOYZfBLoI0TMRhjG60tFjJBmo3jT/wwL
JI+RNqC6wgpcmHKc/eIA5/MaDMW/F0YlX2jjhjszIhsMLzrkd2neY1Tw/T2fR7CNDAyXiyQQtZyE
Doz5vFzS+WAiXbtEfJOnVaLC3R8NpxXE9VRm80lb1YRpbsDI7h646X/6+YOQRx+cQZ/LxRcM1ROh
WedP62bLe7omksbtjSkb6L0NNSIukH+d5rIi66TH+RDVi1AqlRubbhBQzNPG1eWejgtd7yvLoHiP
PkVpkx6GnA9smNM8O9GJlblplBPvZ66o7yzxEE4Mn+1+GFqawtdCTivlHOMY3hXgItlM08pWxTmR
z633jaE94Oe1qWgLQq73P4psqdgwDvq40ldiRQGLt5qPp038cytNZXbc28I9WYwm16rmT45i8H0Z
R3uLb3Qh4if+5hnOmneuHqTdGoJjs63ZIJ5RDhOUa+liD3IVQyQpPv2O896XpaPqJrOSLOAT7Eo1
De/sON+QHbaZX8oUwVLcYBfJXPro94EyOlRK3MT4IBOb2A7TMJ/86TE7+T3faGzsa22Kxhk6IEfC
S1FHhxUyH7x+ZoKhh8YG7XLMhTk1RgJC2/OPEyvffSXJjfmnfw1VmExo79iRH37xUWBh9hRZTwDS
chI1UWbQqQdNH6/XFsGsKhsfzX2iabV54gFKSxNXEPGqfCfW/zFhs5hX1+VYOEI+1eZLyfWZUXBN
eosgJQggJvd1CsusVfdU+8AdLE/ON2FAADScKAxiPz2TSjV753g5TzMo9MH7fSgScItlMdVmBIX6
LuQ90+UbkKmCQKEUVmSMz2/Rdr7O30F3Y+57XbQPj9vUpyTCdUG7q2yXOR5H2dMLYWSVqnArqRwO
DWJWmJWps/MUtjFhaVBXrNH586h2mT+xr0nVSslPKbQyuVAL2bxbpWwi5ddIVIydy9WRlBoAAXz8
6mVHV1IwZuYz0z7KIYIoHLBGNvB9a7J0emg76xwJeZw2HD5sQGq69DvUD/QN8719m6qnSDnOuHx1
hfSI0TEyn4a/MR9YPHx5h8a5fqD3UjGEAOHjpkzqhtVgFo9MFgezypsqgijWFTJOZp/+tX89aPQh
2yfiSnxGou8q+v7UpS3RNOQ58i85sykxmabcdvMMO1rsI0cd5tuufMBjlBIidrudB53sDJB75cyH
f56D1GGJDOGp3O/meXrDa89hBJV3K/fKgXZFvUds9QHoG6trhkWkVvPnYF/q7NRAUzOixgFUqk/L
MAbbwnlV8XX2i2F9jJZnXXXn5Ycy+FVcJIacyKRYoKCjiLZXeEoNoPTPUxpOO54Zs+H6zwUTn2Cf
eoa5Bd6xQ6aBC0sWT51XoqM6GNxVlIsAZKu6eeylKXSHFM6kBhHF4EUrm7hXkuPOY009z/cgtJLV
Nooum1b3JyC5qL2PWAZ46cvLoqvIvk4dL+h/kFDblsWnLhvOM75DmA6caGdOpYyY9v87Xanw/fh2
ag0Y7kbXlKpV2tqyvI0PvLonKAnyffnjckOVm0zQRkZAsG5h5oFQfJFkqnMDAeW2uBHvQZawrYWF
vHGJyKQ+ossA3e7Je4V2S76vel8CyZEuTNcvHQ9DzPY3Oq8Pa4QTOM1DfXuI2gxuAbmvqwqCLFFi
cFRihkP+B8az5YMbOVwoDLIXiKfl8v0CWbnjSJkg7hIWMoojIDaeksK25X9UH8h9EkywnnfA8a/k
eppCQcI3GuLyGChez0acbrucUFVs+S5cxzNYyDvFbdH2FJMmW4lixLjTl40/Kdi2Dp5BVDSsnNOf
CXYfuVyAazeZXI3wiCpvXW0TFSIjBlvkybZH2Ntbidzo/ActJXQM3ftQnRIUgCXeGYQPf8d3aY9C
cyGpjR9ADE0zH4gy0yRhjS0kPElI4fexV/HVrlEphaYvXAA5NEJZuVEmE+zOu6YrsvXgNGHZmz1W
qqr6oGr7MCxcnA2zv/G6f3vzLEzC4QriEYOR4bVI6PBSNXS4BWxd7wvynqllpG0RqEt3JVKFiEzw
1LIOAYKFbwVBwR0MQht3XVv/bBHcnJhhP6rv9svOe0NLhI4OJhyxlce1JmbVrJXZEf21i2FwZK8B
CpARB9asE+jEcAV4Q7Xf9Mnhe8ABtrsq5FqNoYfhbkb5I7R5stPFncOV+8/IpeYWIEg9y355FaWT
Av8D++fi1piPy2UYPje+I8yIhWD1CTuAREkV0YCekvAdWnbu+SfzNzc3cK62lgsbtCI+dSqiWufI
iSv3sWuHQAk5CLRElznczM1jmT1ZZlpM5m52tpV6PVCYKSqTQQtJCxE7ege4ehYl0FDh5SYAu6SX
+PwQ+b0SCtHR3o5yUFW+r6pCKaoBQ1lj116OEvikXPo9rHMYggTMYlY/4EId6RqbkTa3rkBnKvhf
Lh7djZFHSFhYzrQ1E2q2CUUx9A8skt39Gle3W9a9HTbWHK6lH0go3uxhDa9YBAwa9YN8CK7UHhiQ
5GuBei8SY6Wm2fFGa4tjjwxgYzdANwDNfI+TqRuBrjgszqGOBY2U4r/hn7Zr/H31q4z1DpvYXXi+
uYCQ5W8ZzacI2iWQTWNLMJ4utOEj8mLEvLE8lM5n9kGxIFc/tdFOXEypzVx3cBoHVJeyAtJAaEdd
mhbqu9+wd3GVre336r/xHyDJjozmfg8t9UGsNHYUpRbmEE8HL4GS29KBsfPLqYELC4PpllXj9ix8
EV5U/0JWXXLUehLLNMHZWsx7/S/tbdzO9Q8GAAUs37Dd51X+wDosFbpXUSbf61iJBdtraL95HlIV
qrxaDlaZNzrVrlAsv/K51rYFhyKbc349zp2ePOqPSejpraZloQGHCmx8wWpU8PIjc+ey9qWAALFD
7EVLujRGf0mywpmMjsj84gWnKCqzf/6SVY6bSThJL5IQFP3LJ/ELTBT7pOAQDxLg8uGECsg8ZOgq
wg9AjkVa5QxUzMGPjoR3JqpO8VnpuOb/mR7gMf3sZZWnxbKO64/V8UhNonFzRqmazms8nE/QH7J2
qrp7zJiiGgKFUSJmabqmm4sdHLVeyyqqxYt5C4Je9/o/uzTEoqQzNGv4FvGqoZN4MAkJ0ceF6W0w
iHdGY/5nHPMlOEbnlGCKsmk50xScPSUvlWvwOxIYtkcrSWWT1q2casiqHq/fYb6CxAuM/UjAUFwe
JAgkaxcpuXN5bRQ9lnHdKxHiCPNYbyHsTHmyMIUnh1SA0j4y+hcLV6EI3Jf/yqywIVkvBRgiGmQ8
ZS+wpyfAptJn+b97zWg5u5ZA+Zqx6vlqDtPoKDcObc5/F0O50x7MXkOViwdU31OPYsHvtYSN0sKp
L0G684DfVCzj15483qINdHvl/lka08ldEk1D5ZNU96CzGk1tGKfnawa/Okjt2aVPTSz1adBIKFPc
g1LHU5gugc0U3cY42gFjdnt0mC2IEl+l8AA5mEXl80oA0MXD22y/LMFP89Q0O1AcwE50pmOwqnOX
ZkV7Fh1EYckyE/JSxLkXyh+yZaSg9IdWy5eZ/zUestuNxkt/KU9tkdVrnA1XIkOmqlEfAp0RB7qf
13UbFWCO8y7x2etzNWnT4r6MGr3EX2RYNHOyC1tGezWxEushxFE834Gc+KMyn+BOYJrrt8QftSsF
21vc3PF1uRsIBZ/CkS23Objg9mz4wHl69caXw3YJZd4XZb7Zn/tSh6JdsFWVfLeqZAOchxfkdEnu
yq3V0qUJ7sHRF4K8JnutKPrjn4H1huEalthrmbjiOqY9xD4APoPohJCWHFeQEXTWqvoLlTLj5cta
MTuU2g5Xc79oPSwm+yIQ+tcyJViZbkVZfJ6SyHHgKIR7/SqhFNHn4csdGVfIRqVYtY//2ya2bdOg
/CHZO95SKMbtU79nxx18gBrCpjeEio6jLSDM3Gn13mj2j51VJj4xCPYJ69SNDb8sYGferbEeAiXf
zFZWg6NMZYLG8Ko4AmYne96BCDPdZq1AKWt2igJzfiis+jTNpirUqypVU+ptR+BBbYCyHpoFpOaW
hcnoHsppPTOnWdHECQtIobEB9aK9IQ21VP0em9x8LncdSFyUabm5GsvjYVNe0a1K9WJp4mCG19DF
fsxsVYfUlBIxZDxGxi5tNd5F19yBGEdYLqiamRkXdXNktm3wgR4qLm47rjmWnm+7OjIa7wl3Ftb7
w30QVyv0nOa5xeg2+NKRcQ649Y5ft/Ir9VKUWHJ7/F+7TjS3Uzjgtyt3AsiVnkWF3zon9/+EMaL+
nt6O3hIt1T/QBR9ka9ewAbi63UBCgqs83i2BuMXm54S9bRB372G2u+nlNHVP0s9KKK2ik1FfsBNP
ytSbh5iHdSclTZorKfD+U4VASqyJHf/X3EgXHxFRu2wu7/Z9VnZV34+Ug1bKMwyd86GVRIW41snW
27jdwh+/8iooRglAG59Ef+Ljaj9lZkSF/6vxOBrTTyNiwQq/VU2XDLfcmSP3P7LMdS/TEocU18AO
QhGi0bEvdOc4AvZWLIR7YddA4NQE1n+311gdkImD3iKox2qBeaKpq0mjtH+zfv1rUDjo9PchVcy4
xkh6vRv6wQq8w7dDtVsV7wQDLoqJulgUpSKZWTnJXmJ7PJ+diiORo84b9DhrBVYieteqj7TEFzlD
UAPXUwJbzADhA8w7mMhAeVGTP0KAGZRiBS3LkPEZUVNhwNzdCwP5vqPaLCugeNnHv5yktIkXR9YN
AOBW9PaRS/UZDElPCLsUFLXmm/ZE75glSvnNBF4RoEDJqMrOFDJBOee5wxJceXVNX23O+deIrgjz
l98KFgzPxm1y0dcpXek/Sz9+o2gnFhJtY8o9B3l6OkC+i6ib3AGA7V2S2C8Ra4n+UHIZwQjQwVHp
lfVEvVYt0fYH+x9uBzHDx1tLVrDy8NPj15/esiad18mRMEfSjickRiJ8SZaI4i87eucZZ2ToMpjn
Nrz51nEo91iHCNMgNpWS2XeYKPce6P7kOctfP2dteC8ee+QDTfE344vHEBcCWei+Hq8Y9/OmUpDv
T/B8L2ZIIDguvk5+wLcQaK7A+9eK5MjZLNbn2+xE9J5B98YjTjFGvWXbUEumxvgLxkBsSNNkTVp6
r3y6PYZxjQbn1cs/ifSv3ybb/JDIj0W3je1wWHfBiDdlVp3qSp+CDKLwHPsgbmWqUbk4jydzuIxs
2JEWDtMjjO+VOC8tkqeR1tOLzb1MuGPJewwMA5v5W1KIpVuFo2dZdZcCVOMbmZ3ush2fvKrRgA1k
v588JfoafO/c55VVgnsJls+Dnk1rXmjGkVyJBrlIsGJw/MB1HScUcMZCr/YOSjkLBovn8qLMuWW/
X94s6fzLV5lJ3rrXq+Ujmda1ceez4TShdWaDAMVSLIqJUKuF2u8W10xcLKalPwrs8ff5SEroNZA/
NzwtiIXKSxEP69ov774XCnnupv5fqN/Fv90FUg1OvyJsjZhoa1XfOV41kEdWMZNJ6n36CZgUq7n+
FVRUeF7/xQK6oM9v3UkKC9LwPTbpEjTtsyGKAEwIDny2flelkI8qFrKpmwXYFUh5su3mJW46s1V6
HqVkezwNS/UGvQ7nps/Ycndowyiz4Mtbv2rM98zfhQcx3yhew7uYChqzeGNPZeGF/LntApzKjNFR
C+XDcbwPDlTOAxxYDgGLWz6HBIm3JvvT9MwDktLdNika9Ubxts+foCCAkIgGKx32zQpJ0gvBLTdm
ld80QUB7+MscsP2QBuHAnpmJzjHVBKcl8wNJRpFon93Vk+NwTBs0fqyYb6z6OpzVsKPXjWdcP4KO
i8QtfBqws5uR6QwmI4w3xsjOJTed9+apACxoxuuAeKOryww8o5LtGWoVPn4Ycw9gMR0pVm+rqL0D
m4VUgUdN1IfZcTEpxM+iErzDZZ+sIp5d/a7mIonnR4Lu4vs1oUnS+azwOtIoGX8T7hYE9H5LFl13
C5RPmjUuEC6dCZ8f3G2mcjeOHwSrO2E6TmvaY/DF0KlI3ziruwTGCKeP7n4eqdAAN2rGqekjAOik
jb3pammM3S/0Oy1zVzI84L4PTPklIHt6rxr3pQZoT9T2ggL77ttSObjmjJXDRFy22MdCnplrv4ST
IKQknbv0m0W0TcF8iwBxboGp4z5CHBxSkVkPfa/7W6znYWVTK3ATgQAqY6zTvSdRjUscMjVtAy1b
6WgLLCxqh0pBjWGeULITpHDtIb5W6OnMDz6vc5AYP1Nc7s33+vThvcCEiwKybo2Ucgyiv8DZq6q+
Yt5xxR+AjIStI75tjtSl2qiE3B8SkLVzobLO9LbJYKj8FfWHndNxUw7XtqDzcfiS+JOPZIFffsmG
YIAPMZgLwJTb/C6cmsfLb/7naswHCmXnHgkFWuQMMMYyse8e+4z0kZt/MkNeCXaxt8LbvHT6PbJu
H7lJsNWE/K/UdMXfBqO5D4FtJhaVXVotjwa+TdMaOUCAt8ORHizhc8fifhdqI3adhnLKq3czOicl
G8Bm0Go7OgLFfYa8dFBdaaSGw/Of3XlnNYksom6Zp2P0drXvYrJmrIk4BqXgmr3UMJ6UjUbZ5M7G
iFcefow1oD2WcQAMfZHGUEyoFVUYC5U096s/xza0qTFXCdEH4yLYsfece8qCBitaUGTojeSEqLFV
UndmFdV/iVbGl9Q/2uUIpDkeq7heLmh5/S9zXNsUKXw+S05NR8gJCOtmr48zhS95wbZRpomL45fB
0CNInpFD5GluseYuk0Mc4kWSMD+RrDbNuSAm0/i7jI+9uRjto7sr72aZ6OwrXFSlngeUh1MLor9x
2QdJ/kArXO3DUsO0mx1QRlbXisp3ELLqdl8VQ/lpONifVrt0MNCGNDkWUDQUO0ZpfHxQKGuYJl0+
fRVEEykP7wMhU2PtXdlHKNkTpBids5F96Dnf6Tm4aHy//2pat+5slRJsiQnGTOI/3rLU084DHnwS
sEL+iN9czaxG+mhVleQqYWjhIfJjKz+21TW6Rb11KlavE2v4Ib4WZrAaWtPiobR1JdD9Z0Z+8BQk
QymJabT7YnG9D2VjhhR45LSl9O2FRvggEFl6s2QezYcuSV/gyLDFOClKZ0iRPE2a+05S4GNk3X39
lS9nldWSbnJtR7gFrBUWioGyyz4/4fROCO+wkjA6dHDugKx0ZabxSopMiBq5+Wl+UQ9e+AGzoBXA
9IjCe+Iw6n8rSq1qdhl8FwjuF9Kgpp0TQdL+CCpDORAaFrPBe2NDj/L2OuBdf1AQqpv6lsoY7Mcx
eWPhEFF3gplSNoQxpmCrVT+AjOWFvztcF/C2px3HisiqvqaP5xocEroDaK8w4mx8bNXeiPHJqDA+
RXIgBEr6SJsZaJevTEV1JBeOzuJ3x+L61yx8wJ+sjvSXTC6GKQEeQ/4K2yPvwZEz9h3gYe9+PgnN
tX4U9YaOBYcy0S8Fbm7+yY9ntP6CVuW2SpgLGy/hqS/nvd/96NMG7ePDhAeuOBRktaqLcGUOV9SV
tfx4eiCPSC9AY/4VBwsFA8m+8gCyMuPQwMwSAPBAaHsZahbAGF1iUJvzWhRAJ6ivogDn9qDRYdIs
17uxfGWQor7j9PQFSh8wDDdhkEuWWgkUK0stvGZsSPlgRusSkVDjXGz2XLZ5v4khUw55k5ToeuAt
+Q7AtE5A7tyuo1fjLPj+38v1c2kVSmbKrOVoL35FWoJbmmBlSe77Sjq+sYzH105fkE2oE19du555
f78nd701WA0sfJ/c67vAQXeNQyrBET4W8xOzKMCDLIBPDkJ1cKfXpyjsmEvH+VxLewiSp3i090a3
YkSLpkiLUeWasxFD6vtASppWf0yWXmaoVJHLdsPYgu/Ht+rkjPUj2OseWivSrcHg0ZP8DYrzes9T
26zv/KfKotOksUsGY0wzhrxmdR929MKOEZcKSP/YBkz/vSqcg4h0tI0ci2dbn+5wJ+YPqckiV2Yk
cUI9Y86wcDG/mtbVABBUPa0G/V8erXvjZCW6foZZYYtg+tNScVaLkdILRqVIUD9lm3OjZyWu2vHY
8qNw4H13jEPlkt05JQLnrDz0dqBdtK4LDVPP1L+9p1tdoN45Onwmh8rEmUGXXwOb9LLm0gsamIGj
URQNGK8pczVAbPckeF3set5k/KptUNKTRVU06fEvOCyCw99IoOZGa/ZJcVoCJqatu9oGG0LBUYAS
lkle/X/sdOd5WSjOzdYHMQ24iaiRTfWiWLXCpnYV5Lqyi0/4vFwh8BU5NC1xQL21EMjZ3Hr3IThB
XLHsrp6ZvZU1MIjaf+Bj6oKjrbTCqfmAkk/A6IK6IB0fXgqUFyq9G5R2N2BzS1TNxc0Zj50+X+ci
o2KOyQYTQgV4zPT/jUWRTrQYjUw/FSDiwuyXVkp0atMrbWMHR/5SHtGUkHOIWlfNenGcKbH9vaq4
yL6NkTR9dXLWco3N7i4w1GnCfDxIJuQnRlB5/LzzeRB5VOYDEAHhlbwl1YAgz/ycnJjzuWebiMTn
ln/NbWWF5XSW9RAfkNItdGPjsvy078S8zELNEUYzoD3rOpxJ7lENTsQUAS3pg0ryASiWzK7aeDza
DfiRuZwTWgjuuwSyrrcvQRcmyY/yuCYTr+vqZ4bFG/aN4isI2OFm0LiBnJKmjvNdBGQKs6tBCDXB
KyS++rZir3pKl4Z7VPqB0FqqMF27W04V1z8oZ37ebN6LhaYnhTuwtXqQPAVePmQKkMIFpLQqEdR1
awiGSuOGgdAJ5WyhRw5Tz2y0/hMCrYR8qq5hH6CYwGAeLHyna953kUJ0+K8Nbo8mk3ow03/f/g5K
jnQSTB7AJJvvILQ8JEa8aHvul8bbV5FqFSaLDdi5I7PMyPFY2eHSC4tM0r8d7zHxm3MQb8cInJtB
rtyptWKcIHwC2W7PI7Cb/98G3hOJbPzGOyr+l9Ud3TavBAjNcjLrZ9n2iShuAmOP7wrJw4VMmtDq
55uYfem4Cnkqy/n9ZIjISqAD2UtZOKuoAUNc9wgzcAy/IwFy77WGLcrYInCibjrvk2adgSkmRz0q
uUI+UDRZ0WbHEFoVrZxkLC8MZISvSq9FdFRP7UkJqwb+SGJRzV96Gf6TfL2GxI4jQNDWgpGmrRIs
Uu4h5IzCBGpTcZL0Rd+qm0WELg4BiUS2ZxbDM6NWxDJ4zTAFIe1Wzs3kjuSQfgPgqpADUPP01iM5
XIv5zH3AYLcSCzwdHWUMCjB8O7mTlWgNtzZrsX+32wtIBOBxG/4gnUeqNQEPv1+XjaXSAPNvF0U+
7CsMq0nDicZuwxkUHiGxgoJ7QqzAErQVgzq1hfs0h0OQdSLR6YVF1J7tqTTGjMkiVpq/z0FkopZj
PjDYD93YptaDgIZUi4tF0beWZEtyOwho1RADmCAyYe5WgrOjInPuykFtOSk1F4egU+rUFdDO+vzt
25h5M2yvI8lN/s/PkuwDKXSiEbmJoipYoIcLoCuBNTcqdB/3bN1nqBpdcyie5Qjy1hEP0D1m+lGS
eDvf0EXFm8kbtN+qw4nBlj0Zh52Kb87EGDPBCDYqgu98iiAlXa66TR4W278uxZYP6Ef2824WeJ6w
dwlnklHwR5v9YV8MJ/V8FGyqEYj7/jfDlAhkTf1H+3Y32VcG/dKD1EkS1Fa0B3uNUKIQPHexDUm/
vgVxwhC1ycDxrak2aoXr93UDvtgSa+LUAIOtDdARJQh7h0t6vbRW9g/mnwRJlErRiDeb5IEVa8Y5
Anb7tOuFkGkz8+VGxDeO+PEH0/5+4Yq9zrTbC+Ng8p3FH6fnAL4U2g/w8JE6HsWjlKWtmGx6z4/I
Vm9yEBaZ386r1ETpX83EfGXT8Ku0stlLMCChMRA6oqiad/jlQ5cescvm3FaNXzK5BoWgbGJWmB/T
5Mw7rJH9cCY089j4vL7va3UgGUgBm53uBs4Lx7L2U+NDvYfF1xf8D0cQYJuUFNMogAAQmDxFb0v9
oCMhTh3Q4l54AUjqcygXV86pG6vLo0DCwywrmM1F58CImJ/NN4RB6lWegTF9virbXeehnibXx5sO
MuByfJ2Tpd4luBHWJIiGFQnWKupwf9bmEvVlEa9Q5GC05WMX0hDHiiXcGKgIK6XyEfTLd5spunB+
RxnSNHkpZNWuS93aFXde/0TamQvZqKTefnbiX/TCN7iPH1YhpOTSuyISEbpIQiO/yy/DkHrmtI8V
4Nl10aDuRvp6+6gUBJLPNVDM3KhGc9paZmDuIYUgsBRY3eKF7zpOLHcJLheqChDIZLQyfRmb2PNQ
7BM8+vEdjWE3caABiM4K2fN+pPYxPrQrom/+jrvor6izKYqxuT4/00oxmhH6yoMhSiztgBqOgjDW
jcIIkQ7IcUIjlXFqaPi4xHvxWGoWEzcHC5MPf+KzN2sJW8yhSh1J6G1qzD5dlGyMObUaSNnPXMGt
zLC6FCOE0ifE7WVBlBEkOQXv8pPd3uP/0cUhpQnETERduh5zN8Rxl+yDkpGJ89jtj/3RQpdx6A6M
8qVGKVqNxwhd08qcnfAF4Kmq4mI8dWqh0e1xkK8BuvJqQPUJWUKdEzkzahOKtMRj/dcGsrwRYaz/
TK2WOEo2QVuW370jU8BBS0n8XrjViS8ok2QRb3UUFY0tTwKqNZV5Tk1Fk+At3W/Qe6ayvs4CSfUH
3R6Fnz0ROOSsexdJA/HqqyF3miAt1TyI3c6sBvvXE1PfAF5zZ64efqjbvtQSfR8MoLLRSBJJBLqs
/+M1R1c7FxCaWrP3fZG+QNwq7Ze0q4FJKx6dJN3SR+K64Sejs0DitZ8tIuNLbDbmjE7sr68L3W8P
zJP8HjzcksLiBTJr05W8k5OzCJeqNlDyCVAbXDCZ4hdLnPAbab3Fhf0Av2J/CMmJD9vbjoe8G9R2
a5djibiHVasONWpEnhKpGZmYYXjOawL5wrvLCXA4lLJ7UsMtjFpKKG08ZnTq/r3Gw57L1SGinCYz
JPhLBU8a3DsIInslR87sA5KkLUh/hYAIJM9EfAPPkah6Py4oimfE/JQOXq7ZvGKumqc8n1xQTDfa
oixRWSRsWPUOdRDV1LiUr/NgQmVL+zB25ZK8+c5LXWvq5R5TayVfYNXm0UKf1dhZkchxB0uYDpTD
n5p/1NHcCJgDytHDxKdC1YsCwfOT7LBC5befNk6XF4uEHFo0UCgL0iWKzs+HMUVafP0w201MHTCq
jW8kG35+AA6HWhXNi+0SiIxg80Cyqm5lEo4LdMSPX75Ip+2fOyOgvaSxRBSiqbfMxzdgN5pfu5oO
r9ID1J24RviviPdr1N//uz2g80GqbCO71UDlKJLFlhS98/tlgs/q+7DKbOIYQSw00pqysf1bZ/Rf
QI0RnJX0vabY9bXx03Qfw0jj7gwtGb/lV6HvdqHohyWAbHYLQ/K84M+NkSUvBGSkMZAhkqqg4d1+
npnGDATkNlVXYipbM/uRTG5rF406YAMpNRtboOb/wxHcTEYZTff8pHhkZEj8WxAMGrlW8vET604b
6kDqZBP/OMYAEzdQDWVhXjT519MhbCQ9tiygO8hXue8JD27Gtj1v25dW7+KtObN4XUli0uxNXXky
QXoRWeOS2bKY54wbptPS2N2FgpnZPiueWKVhXSH1JiAdrK0sIqlMGCOPL4+ijRI46rr8C3OYEdtG
XJKce6feUNBsziK4ZDGLlt3LulYzNxtEKs2rA36uo32JgvQYORk0U/gzMf8HgRSjNwPB70+9oLGi
04wtO13lY/165A2l2VeKYSkG7soqYcfkIt1zgPBIk08bSIKXXkFQXquNNPmopRMiPtISzRdGK4Di
7HEbmVsOxKunmLSBnW2tAJTWW6LERyZ+BhS+15vdVmtbAx3PGHtslvVNkyWdT8qKeB7gwOJgsyeI
SrpBxyTiWoUwEIrrfefxiMG5VH0KOROh9I1oI7xNi+O3vvy5rJzbcMZmjIxTI0DB+6wmLCqqfabM
mT+wUSkEQmmAaacaSV+hg/bhySxsa82X4xxGMETjrV8UNONWnAGNzH+0IAilwy395xJ8vd6Ae9aq
v3IONvYbk6G4XrrujHoDflcRfTMoeFnUm1IBvWw2H8tet3NMTvUddnkMmJgQUL/VQtHqcB48jZch
qD56ItBeSEVqHzkGJjmS9dy7icechLrDwOwy5sgZobxwkUPoQn7shRNj4fNPMudXe2QeTKgtU/NJ
N96Vt3jkRX0WhiVY10fq0LMtCouGS+0MD61hLMY9WtjmJjLe5zMHBUPvv++qkriyF6k3Uq33gYQI
4v7pK+7BjmWtahAfgg0Pm0vmyOBADJFCv4GBv8m7Xbh6K42PX0sWVKAIuI3KCDlvO3h3FelMp3XC
fVCnjQJY+Kuu3z9KYkisnfpQ3hcMHKGDb2Il0uXOS+vzz5etTqWOKXHZO0QK0DieFc8AzTV3wjvD
8pXEed0pPvRjVOKdEik9Mrt55e9fRETlB2avAjlnc+ZZlC1MEuPLGHM71y3PioBfg2eWBdZAFefo
LugiSKtc5ue8LAkISFT/GCyXxQFF8BFfnToEE1aQtlg9EeuWgczWnkTGZhUWVGg9eengBX9VaYTN
yPO8VwL2KLmONGuQg/y2WfcJsjFfJjQLpFMry82Ueqzpk60pvCyd7kzWN2+KwfpNEszztPGM3HFl
C4QtdMo6+pFMMV4DwNZRVlrIXz37/kcOrjJdrzqbL7cvoQAPCL+IXgKQaCAGXbYFEthTFnT8utkp
WZV4CxfbI3FDnq8RHaAAaEcUgAgA8MgkdrRoDwCLxSh0C77g61sNtRR9jWqQKHt+Uz+DHxVd0kOG
SKYzbq6F5+PyF0q9W55LsJBUgx7evkyn514GR0jbKEhalNHuinwCITRd7f57ccLZCO7ypgOR+6zJ
zoHfYNCkycShvZMBb1+l3X1Acjt8SScRGWkMZ2BVhC+Vb/8IWfZZGf6Cr01DExrj+0Tnzmtnjx8b
+X0rbPj93b8W9Sa2PsWzr/CrHnOJ7okJ9C1+JbpMje2VJ3npxb/GlAQXnP5QYC0Svf8DqwJAEpTx
Am13SHWTNfFlEC3PvkzH9sdRsMiJpaug/QM4F0W7alh2dyD+XuUL0AJI4bgxfJwk0dKOi0i9lMCc
HBiAWZ9ICswKz9DHG8B89zsulTuOWB+SJIbgmEGTVRa/gxTikmSuVZhye4L0kyBduPfoxTMfjPom
Pe1x1eukqBCUphfjs42NYtpNIrrLEQ0v+O1Gjkn5+HZqu+4MUAUMCU4FXJnjQGO6QtfU/Gs7KrD0
aYFrGMPb+LE31hg5qf/CoQOboYu6CZrMzSaVBU6CEMzGgUyuPy/r3VoGs7HIS71hOCSTq3TXdG4N
q3nwG+Bdhb5xJwHmMPXDF+oAiRRoUxD5LLiJWkWPOM9XZRWGI2HX0hLfR8lwjzyHgKgkW52tFiYy
lZ7J7q6Di+ZGylxY2jrP/Akbgpx0c5+AfkbA4IBzF/EMVtv0MmNpesd0/yk38mc32AuRAtcgMVfQ
kLmq92NwHGAUI29tEsydmNRLHNLhlIabgaIOaforK1J1bCEAwBn1FXaXLAPM09wJgh291eJ6MRCf
Ps26j3dmIy6IiWrBZ4M3tqVsCfa5ZlynQgQHiC7q9B6UKjlK3F2lC8ICTZNI08YPAGxC1KKtnZOq
msrIJl9o2S1WqwgcTxDv7hC7RH88w8nrTi/CpygBuL9YbuD4YxHaoZEdiaBfJaW6B3QpC6pBGpnw
X7xvd4XB24Dj6Cq2p1/glBpOcp4E7v3VW19fQ5m4V86jAF+4FsdHJNz4fc/FzT4tXtv3RxDh2rQR
8Gzdsyd7pot2My+oyOREDhn2rXK5eG7yM42grhqIh2iUYtFScpbl38njxCKxgUusGHylzcbYRbvJ
fSX99MW/NeLs4t//nUGiR4qqMJGZilLukBCGTxXnFDcfzRRcbQZA/rM4+T+aTJXQaheKpX7fWUrG
Wtlef3jgtoXMqlTUCgFEZNaxeeRehz3FEXBxiIsJuJHAn+A8P6IVIdccngc7JPalSddGgYkpD1+b
YXW83VC7MAHXKrpu+Jzgod0wSBIJrDV4YJQizo0W7JYqerSlcCOxWi3N+29UX8ar1v2y3YkGnn8R
nZ/zrhpnA249UygQLfE6OFG/QKUgbDNQoUsOJtyw571mDUCStWztf/Wwxo8ElNlA1v9DMY7U9Dqo
UVwaDeWeHH3r+HpY4NAzU4XkskWo8kwYBhV3paKiwyGtjME/r0bME3XcnDpTNsLKm871pkBf71Wd
b4Xp/9KRLUSTfoRBwanCo86m3yWICuoc7Gmzvkbkk2gj2Qd3Ob/bN4P+MU3YE76+kWDFjmeSDk0y
62oajsONrputWq0/AOx2EFjZtp1B9NhdK/MHx+ZWmG6YZ54AvPK0q3RgXTfk8m1aBAQOPhikEave
5m730MqVlJ/aCNR4lXHRjWa1E8+tn17DkJm9UPPi1UsuTcQT+mIaFk7LS6Eho0iyNTQkVCuNOnyg
ZJWsXzS5QDANkW1qVzHXPUk06Skoja/69NMWHyQRkEm8RizZYkz9pLTmcosgdOa1L54d1QGpmihH
s6tOVxFseZ7GIopgWXcwqwMl72T/EwqU21QBOaaQDYnE73Yo9UaEfoUg8pYlDCuVDSGjpLWwq/kG
J8FeSr6LG7rQNZXygPI6ZBz6iKc6Gn4txnKEUOny6FUWT9D6R4rrr25jgIcaGHegIm5g4BqiyYtP
nZiSx4ZVstwDI5qSav9jR1ObzLu/BQtyqMfRwElXYshcOoqt6N6pW32EYm70OlOnTaK6mwZ+bAK0
+Mih4YcQCNzbWeha2UY7Hj2E0Is61wm86OKE2McUlpWBpSWy8pvQSwAFgXn0a6iSn8Ol/wtlPDuc
/TVwbbtItLSj9y2BqQM2JH0wh1Ei56zXIuXEWpPN8y9+VELL6yvrbqu9uld26waAguL7aKeXqMR5
mzmmgLVb/pADnwWROx7SvuqTHFfu/5ygkINXMxma56rKU/LRSWeZU5FHcsWmC/p0GU6o1dNeN+Uv
qrZefaKM05Y4IivN67xFtcMdt2BORElokWFGsSAQvueOHyU9c6JDaFAmzImT6JC134Qsv1wImXvP
R26YTOtu1Wy+uK3b621SSYZ8h1H0ujEQAibTgrrylqtVRv6yyovGS4+nqizdCQcKaXzo4gh8muj0
Afxj+84pPd/uVndhRj34LDFZtcA+a5Uob5jmf1ZaHd+1JG4KBqpVqg12wil0PZYVmUWzXIpjC1xe
JI+umba6C0PXYfzMSFwScTi+7/ysUZQcs7mQYQujHAOvCevCK6YW1m9nfGOSS8WCFiLFOmmqiAii
wOO0/TWMxWlVjDDLy3EDc/3MHeHQfF7njDBgtMhY5WCZb1QuySJImE1BvUXqtNZTeJdrJkn4JhRJ
49u0yvupG4y3sX5uQpbl08do6Duj7knAZgEJqdyAK4eWcoSf27AR1N0qB5Tfw334pJlW93nrlxDd
IA+60tXRywOQ6dz/IuI0DXmgacrV+RefR4w1jSYuUrqhcGRXCgefpEyIwLsnrqYnGsQxsmsqOEAK
NmaIRH1UnftU32OV+4WdibqCtqVkeAsHVaHATsKaLEcRS0+d5bW2yfwCDSB/xS0TJppw2+n7LH8e
3yssfPSa3hAhohRE6L4vYvgsjLUb1D0dQAQYfyJX+ozOPuAqG3TrDYw/XDQ3ZhFeeKKUOBLSu+7i
Ts/0qJilY0Gdr2sOjdb0MVKRy6JOYkuIrkPCKND7ugrD6E6iGcSVDPD4DFpiSMavcPUuPqZPZsFC
gu2qAZkm2PIN0noeXRzVIIYBbw/t25XVXnfK87HPnpT7KwnP8U6m6NS3iWFimKqYgEek8Eje1GiG
R8QVcPo/XOPqpBiqly/op05Tpu2QQ0sEz4DOzxUwgCGXy1X9tEDdj+R9b3raadgSyKFR40HPEzb0
cII+LJzZpwg8pXeAHI3FXZn6DNQsp7/ed9CPjHdMsNkzWlqfSTiL14cDDJi84yNj66BbvZumJC1z
OBMp4xOZYYlQ+W1tW4sM65tHkkz+rspzOhr6Gb/MNxVyJX1nrE3mFN3N16JdiBK086kJFrwIF7Q2
77hI0j6WEzoKGasQtjpKcVM8UCpKKOmoIKOV2DvV7mGirJTgkFBSNVhiXI2FhMuQCBVZVi1UCxrp
0zleIP8OMZg74ZB9apS1E7Qv5Y0Va4TiGzCDgFO5B6AGfqr/lHpe4Dfv6lr0YNz0AkUFQj3cQt1y
INyoUmPc2ACg6PD4MxAAVczrCFH8r7OYQkXvpnfwr/KZ8K2PszdluyeJYkK/w76JyIiCD0KNJ7Ax
R6TXx+iVgIKJSzukPR+e0XSl1ykc5EukrP2igvcAoYtqWP1oyvcZJQZlTXrDoTO/YQHUDdeLOKfe
w1Knr8odnq//w8wkAUf+Kl1SU3wld4WL0M6kbaeKLf7d/iup+QeTEdoiQQHdnhjpwRdib8RR/Lgh
BaRUo3y4XP0Q58b9D0fN5yxCTcBdK+iQbeWHkXg6M7J4NcxTyBzvvjPJahWoevt3QCldqGV7z8C/
mH383ME/wSfdzHW8pCbf2R1drPSlCXWHE5MRYQCFPOWgBVMRefgbyvO/XYRf41oX6QTD3GFcV+Ug
Sf6YwW5IBxkSlV1twRzNOkOvKFChTxbGBg0lj5lMqfaaZC35qCYAxeCmSSFQFD4XDf2jnKuWSHky
H9+WQ3xggPoDmz+pHrc7zwAlyqhFdGxSzZaHl2SDRAFQsE+C0L8+085CsBtgD78GLPxrUCOXbDJZ
B9/RrxyakeVjLihic8S2/SLIcUfBN6KBaADN3IBUZ8ZbgEzg1v71AeiZgIax/Jv0ZyIYFsghcpUz
HJviy+Sa1RVnBz8klLsjdC675jCebD1rBMINAHcuq6HQRGq5T9I46jDLSyF5UdfGZsak4IVTxwux
lY84OEwgGrm8yPlJaC+rMDXpZO3txurp4UhloMfYvvMGQSv6LfEGE9v7daKgfZDyyN6UNAcbsH4D
hT37KoUJBHWOPmx72awp3R1H9UclgZU2PjzsVEuUP198kIfXDKDVqi60XKYxoe2r5dpP5WRskFij
sQaUDGPlbrZ00BX2/knk1fh77oWqK2ShcTAfF5gMytHK+aoLxMMieSe0Xz62Sb9/Y5M+1zMd7Atf
d2D0GTxLoVSpgSLtCGfNcH72dBxuxyG+D/S8G6LfkqEKACRLaGiH6tkLIK17JYJnDCDbK0xU64F8
5X7Ye3DhHGEvHEt4vdqdjSl6ZBrjFQpVcEkDBvFlfhomcl9gQVAa41pM/pRYzNG+9Xi/pfQEHwTh
8adZEg6GIdiynF2f/rtJ8oqVRpnHIxIRFcAx60taFe7yop9Sx3G4fSbjtoMwk4BIZhobJJ9gay+c
yZ77iCXFfAhPSMCgW12hmDJHJ0S0b6KltFRe6clB9lW0Nn2u1u+dXjYDAD3oifr5+9Jv+ycXCEkR
tLlYXOssNk7QPEJBbSgXhDi10i0o08n7M+mcZLDogX3ymJZ5KgKxn8H2q/BFG1W1HSb62BrQYilk
2Pmukc+zEUPcjZu7ETR/+yqPutRfqKCc6daaLMxivLAGp2L6Lce6w1FlI7bdmQHNjCRoSB0AQlSM
xWAor7KWlktYHL7iatGNkKN90pqTrNVCN8YtomVtJ7ySg9/uohqigk8mZobplBI26eZwrVTPOQ+f
/ZWcsrVT/azi+uRys7dTt/7WHmgHfwO/y5dJ1pFs1G3qK+6VgyVLOIa3WD8L5G3hkvItiTEh8exg
Zw5A20WsdBSNiWc7Wt218fIxT4f4MKFBZTTQfTiLW5xN+x70CPllu0yni6kPE/ikGH6gZlX7IcTj
v4jtKOrRn8dp3O9DJ/k8buFzuv80uywxngDH6woAjasmmRRW0f9z609nHYUXaphAliOE/IwuAAZt
Zj3XBr7ZoTuGeZQ6BTgV0qgT4rtnqGjSAWoMN5oXULUDKN6Oi5zcnX/r8BKgwmW5SZqDgEk/WaMq
gkK0VilxtCh9wNcDg3YL40OSyBytvvVnxj1vwxFxTMTk6Ab/AwGtK+KO2Ub3mIXSJZUoc6wmNvTz
O9h7m+Bb9akwq6c87G09AXzonFO0u+gZc5GAW2lwYxEwKN+jREOLCbUdQx8KvCQpw5DMM6jAI7jR
poJ4AtUHyFLitMVdg8JWoCk2cLx5OgMQBhF5594//Qv4YT3rCV8BiCOsXB433chuNfYK1HeAcdAo
fqj/RqLEgOO/AlejRmmBYD5KH7IyoPGdmRN4fV/pZiewiVg6jinWjp4ohHzygaXfnY90oC0OG0uw
zFu70gE6Qw523Pa5zSMDJOiHSPJb7c3rOUQMpyqVH/YLU0C28L8CbE3M/sawI48/Clfkth/JOTFA
pizkSMXliX3Fu+8fvhlwGMCHEGKCHa3SYYKfvFMPuhKDZkrhG4Rt5/Rv3s7vZemnTLFMcn8dU3/J
mW4nxJYfzbJa5e67iM8OCtrS+olEim5SG3lXcXuN+iXAQWwPbtqEfS95yiIjUjccxKYZFgZL5tcs
tOiZF371F0C9VRAxDdAPFN0j936a5Nx7n9Vb8gPbvrsUv56EX4N2dNetVh4uzhS5FjWEiXt3PWRV
wK4WudbJlICrv8Q2zlM/ymVd1i5+sxhb7sMBG6XTZudYe+HeICIj3B/mEiVHDgNKT/VLojQY3v1B
FLXeK1eTmPZUf/whl7Y2zDa+k8wqQWeTLKLXYSg4tat0IGzsyM2S9ix+J5ifjrgIlBEpL0GDyLfx
oS6x2XK6JzVveHoXPSSvAngAL+SP0dUWK5iIzZfv2YmD41Vtz312M8+hKzwvioVUG7SVJoJGBOUd
JaHx1s3raaq+jcbyC9+aHadpfmt4ojlf/iIczAcOgIVZz1TlGJ7iMOPeIawcJ+ZbgTVkPDRlLpm9
KJpcTP4zyo8GVDL7IhGDoL4Czog4nYfMXAzKedUdYv9ONM47LzqKqi/JpnPQfBHaPhr2ZTwaTfn8
TLMQNWUcolWO19yUXT3XVjiBPERpICsYKttT7UFbUPMprhmxI9WS9B4xvHLRGQlZhnQuedW9slUZ
R2Wsm+t9Zyoqy/JFDUckV0MTWjCKIY1MZvAiicExPYlj9/VyA3YxTpqTfBSREmZm6CQnx22MF3bC
rQlRflAv0ZYuXKfm+Z9Qa3xCNSqK3FFtkgTal2dWjOETudTtmNSc6+2eljEMVK0hz9dDaUgtLibV
l4Au5RXK89waS3EG0jF8ctQ+U4m9IJbs8hIWBF8EzsfMy0FdG5ghg/2f04dyv/c6jGPy/OjEgTep
aKfUZkBUWurMXpeJ0aDFH1IhMtVk1JyPO6HL7A1CCLc8oljjSwBWdZt/uhJbkR0dr6NYbKH+PaUL
Fz+r8UGKJa0dUpbcqHeASFaM5vYh1kpuY/zMD/r9iOLFk16l0j5sdqxHVDRHgRmg1Xn1GjIrrqPj
EErB6r649CF0yQvEKwSpfZJsMvzzwnKL6v92yrZNgs5FMr1DShS7GeCMEhx93+lDColjl/vfYxZG
AfJkqmhWQc56Dc5+JDsZNuxPIN2xUHFOfJjrysQoJzk+YXlnIWiZpxUkCyfw+8/qMLaMuboFeEX2
ZMuxeSZy7fiPePMqOM59ZjhlnZ1km96z1fdbO910MZyYqe5XAfqH5Z+T3DLhu3I4tIXN9zGFslYd
6Hydbrammo2XlCbwKN/IQdgZtdYDuAnLdM0Wb8MfAZWyjCoJXTiLMGIURjN9YayRqJd5qaIuD/O9
hz0u7DM2yB4G9EXyLECBnCgdqKhomb7859UzRLm/1hUoahX6E06z6R/6HEvLW49oCzAG8pAbRc9W
x7Gz/YhkawQiyN/ez56gUS6RlzJ91EkA8klI2qBI/3pls//Y8CXbX8FEXauo9kH4JyMFu5u96Y0i
hwBf0WsiufqpxJdtNpXe4doLss1ge311XOWBw13pwDNKuvE5XSkZSIictheVjU05jk1XmJOd7kUZ
BgfnU1pIjgW5X01arzkWC0rUW2jsYOqOreGRbRIa+0mLbV6nHG1iMlXup6aFbOshgLT+MruBcJGw
OyoEc3PQLCl9nzwjsmHphY1wtRybm506w/tbiKnf3Q3KevckhMNxYs1w/jS05ktmrGlkeDxOJ3mP
x02UobOomxAMuQxCFBOCM7OdOlFuMAALEIyaL2YXhnumg5pme4L1owk1nMXfMb/s7iSoLYZXuFpR
u4W6dlfLJGicY7WfIt7c3eAnkyBJNBjMr2tkpqnTafQtBeZoZ/nebtpvy6cwBZF6m+F3D/8/AaDm
xq72kDelUCUBAtEfadDWbD5sDVopBzVVwseDEpN6walFym2ooSwLmShakxPoHDtjvffiIauXH/L5
woMZSSbbTQWG0pvc/v2MHFUltsTfeonAzIvPsJlyNErZZ9vxnSz2uSEYUuXP7caxNT+kFywc8Iw/
h+kVQ/xe2oIX9k3KGr91INSPv3PQlxSVYWh4JUVm/TjJEaVWpJmIztNNK+pUyynj0IkZyXL+cw72
2+onV/Gi95PncqIFYs1m5nMkmbX8Wa8njB0m7c9I1usHgh4GOl0srLANJgmrynQIcvLZUmgWsje9
mOJfRxkL/gux2IAqexQYZ0n5CjDx0zu14WITS7NAVgHnj43vRFpqsHVwmOcho6VJlMNnOomNHYU5
+kTVwgqftJYVWndegE8kxbJusVAZDrElCZUIT6WM5maNrrvqZ5NzPcR9ME92gvhUWorGvb44d8Uc
KAApTvfI9onMjFumeNAjPTEJED68pcR3C+SPRilhuJmyuQNw6ZIZElmkUcl/5ZEbwMZ2B96e6qEe
omiTtXl02cEyrOkbLs8znvtwOgKPCmaO1tCFTKai7sq4ch5IPgzfhpKyiaLVXrbKqFCfsjzeQRh0
XW3phqMFe+ljwv1KShgN4xnSy86/dt6VLP9Nu6QB9oYSvaUHIT01xSWBB3fhBzsdO5HNcwnbWast
YPTcFkbip6OYlozFdQLpJh3VzCG8qcLk6MX/EtibYTnbjCeXR593vbMX90d+CCOzK7WszZhb44ku
Wr7LXYPYEgbdi2LBUZaNycIVlfY0D0ytBTQ9vrv5f8QfZXKy2Owtb6iy6JLRM6nFrfS4YmAepoGR
9jlthrLue3AipQnQQqhn/h15GOxQ2aFtip14m1idCiD0CesTHeBDMXokYJA5bQqHtg0YPMD5U7jQ
/2s6u3Wrhrp8pBnRpn+uxoRV9LYrFCj3HlBOrVNvitHZpIQQu2BfMT6ze/QVSduj7XixCVUvAXHc
D2jXBB1UKZElGgZKv9a/bCRHKWoX+rOo8gdvJQnRSfZK2D4+HExOc8uBbsPVXQW+ogMBcUYMdHWR
lcrKmoOPODfknJX+zNwTSYFa4i8c203i/gRHtAD49urRTXGaODMaVt9cbRW2SY1h6bOM2MDmOgUw
pajaTOIBm5hsW8oqm5Z0uR+hukWugaeGIOJJNwk/4cfjvNLvAcheOebTnX0zps1kEeobw0tJQkQu
smQodQ0ritElNXRxJTUYwInjvXXfgCYTTZ9pXbNxbmY6+56J8ByWAHRIZmo68LZ6bf3BUfXjRFEB
h6YXS0mhgrbneL1pAQ1ZUXs1jcfCs+CNYyDEQZPP+0JcpwI/LoQCE2c4pwUdCihn2NvnD/c5gxLI
NUI93iD2t7CscZZGwKgxiq5x55UB7K78InEF+FhXA1JLphrZ9edIMNs6zevDmv6MahB+XfEGWMDL
Ck8HHWI1LEcE0fPtFQBQ+oXZ3v8lHe4y4Ra543s+M+6sGFfa5Qm21+J+bTtV/O5kn97Ur/yn1zGy
dn5i7iF2fw6Vzzr7vBFSn2jdHjQzOClWpgIWqYtpEvL9QIy79c8FkuOt0/6fDDCKDn2GZVAbB26j
w+l7AQy7yPK2FyPW111dCgBwIlTxnQSzDJad1t5fvKhpk6KWS+TG4cR9ClyoTak9pnxrCfMb4sP/
EVyjYssXNBPCgwAAtCPInaoyjjqhICmRsca+6F3b+0Dss0OS0hCOJDcO6VymZSBC/+2La+lJXgGH
3XCfqVtCK/SVrrH1IGwJJDFlkE/9M6SvZsyXnLVT3ASuMzpxyygmPFdSVHU1ITRd/b6C6aEbJdh+
wfkcBHoNIWAt5h9zPV9WhzWxGyTEMoodlxFmc6duZNl3TSw1Ml+Q87cT4j1P3tUyXGdKCLsUUKkg
lhIAUrnLcYUIUX20ku/nRaPA8fXzy5xXOJKDmiqExu9CkzgjzPtgIimiQImsbXbBzRYwhekKqV/Y
sX5393k8ovX063wKaV2xkQOJ4hReDQoStMVBFYM7c1SRF2rvldZ1OFZYSs7DwwK4ykoGBBT1Pk17
Xk7ekk/onGtQKteOoHmBKc14XD/4CkAYt6Or2PFKZz+5PADh6HXz/lDIJT3ob1DqAHiT56KHFD0q
0hzaT/zR7dSvjUfsVIE4C7WV9/lPSxwqrdz1ScSYKy0dTIMSJbd4ZTEjf44+DRWARMNNzvo2tqb2
2LdG7layPgCNd1uvtx1LU62ZbGNsOX4SK3K6Tz3X+IKpGogZQrrDLlyPh8aLvg5hoqX85pSWq4id
xr8gEhvFHvd7PqPQGCvRJxNqurBoVZISRlYjQe4FtBPOza7B/tuLVwrK0Cbi7QhHctIQ3L4KZOup
iuuh37N3aOxpUr4WSpEp2/VlyWtWkuhBpFBfYsFOCwupAeZuvmUFgtkqEZg649hq/BtHF+OPDsb6
MMntwTi92RYfsS+BfBvSh4e82lz2qlVmU1/H45gAVruKtglGWo1K/lBYztqdwNi0N6GOHXjqkuxj
d/pUQDxY+x8y5APg4zMJzniCzl9+5/rl2GE7RO3fNcAlkd1SQIjXOGDXVTzRqhANMoe4xaOXQSTk
RaIWzSe+xFu+ZHgkN0/nPGR+zj4vzpd60utYjom4KHzcOGlfwVibkB5hUPmwR6zKnVUFgCHpKgIC
LgpOjg2H9x7NrYwiH6mTx+TYCh9sOdiTdFe9IhRI5rDE/ZtEu93jEA4Xn+nGzh0d/FVX67sh5+BK
LER5p72edG1/zLqwHlX4hVNMQyFqr5AYYmJ/kKgBeqnGaHBWtBZj4wlaP4yB0HNtMaVWLpaDPmdz
kekUfZ2nVZgxONQjjrxtStaPUzYFYGhEdSDRqpYo30KWWBy1I3XKb+65Gfxq1vZkZ3g5lUdVapJM
1n1VY3nwrqDAZG/tjKaABqfh3mIELapvznWkCR5hzZ1/zOVSvZUc4X7NTYB4GV/OJZyTYJ7hPvfU
mzDQ1rdR+XLzWFh7m1U4aRlJktjjX8ovENzUFyp4TkJxMTF7Nlx7I79S+4GsEKs3dJuLeEiYl/r3
oB2ffVVIjeqq16yL9JVx6MST7FAXY5TrUpWE8D/OuHXnM9Q31hfusx9S778OGpQZviuXgTeadkYf
KOs3BfnPXM4rfZW0bnkmRf3CIegCAmFxVMgWLTtJzZz9C2tc1FZbuYTLz4uJWimDCN1QjM+lIG1U
1e2Wn1jcWjNaeNmU4kkgFCHX9lGY/By/8bVotq42SpWJT8ucT1nJQxCLojYfzc81sVk+dxgBnsAJ
dl5pTCn4QAJrCQE=
`protect end_protected
