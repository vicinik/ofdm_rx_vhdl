��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���,�Ô���h�Mk;wjj��em	f�3�ON�蕮�t(�н�r)͡��y��O�.���J0/b3�g��`)��*�n!�?h��nV-�RR��q�E����Z�-<=~-޼������ 2�
[�6����_F�s%�'��Z��kXg:'�]����E0r��2lh�]��UQ�l��$�1�����U���� �J@����^�31�ٿ�tOAE,�I��m&���^B�s�V�����M����8�2�R'}h��P�[0<�y�P�HGWE3ͯ��!��Q�Y��m��_��U*���^���0��T�Ó�b6f8cq�MdǳQ���H^�����H_C�	/�V�lC{��5H⣜>jl�$�Q	V�w:u@�ײ�݅ԉ�^$����r�C�A��FQ�E"�0��>���X9}�G�����j	���Q[F���i|��Ņ����֮w+&k�?���D�p��S��q��m�S���,7�l��5[���%-H�X��wu��C��0JND�zXs������o2�dŷ�����j�$�h��W3��֛&�/Ǝ56�AZ���q�F�A��KG�˛mt�Q��'P'�����$��u��j�χ9�0��P�)��H�%A�B���E)q��#9>��4�*I����R�2�;^0'�n�q@)��Oob�%I���U+@���iP��i�VI���g��2�
٢����v6��B�
��0���q�У��U�h����#�S�����5�-"�q�H�W���'Q�ˈrk�����a	�����������}m:g�	H�mMQ<�>y)R�|�`�F;@Ф��E�(�gq�b�ui �<��=]0 Eߥ݊Ry�$F�V��"�*ж3�9�xP�� �ed7i�YC��+1a�W�)������U��U1�Y�W9N27�H�<��C�a��N�u,�N�؀�N����u��S�+���Q�:���kɷ1J���h�g���N�$pxP���]%��M⍸U���,����I���@$�4Fz�V��ЮPo �p�p���
�ᨘ�}I::�9�ĸ7�|��Ӑ�� F�*��I�M����0Ң�Uh 퐐|��h�䛘L<�BBkV$�>�_���������o��\ٸ�d�TX&�:l�"�Z|
1�����1�!�Ȧ�WYq�A�Fp1���ǽ#	�����9M}�O½*�s,�t��$��(腼��Q,�R�Y�.OHuN��8V�����/��.��?{�d�~��&2�KJ�-���?i'�4�Կ +�ܸ���8�)�2�0"��  ?���P�@�]y�^T��𽟵k�Y�al�
��X��O�W�]�5:�a=��8�-x@��G�E���kˮ�$��޽��+�k@�����$j1E)فKvt7�,�O����^w���G���w �/O[.y d#��$��P��9Ryf����XqΈ��kK���*u��ݰ��
�t+�#;#��a9��BH.��x����ےʌ��Z�O���"�%T��1��8�'R"I�9*�����a��hn�nt�Y<��08����M������!Z����['y�U�p!7PJ���]��jX/���Skf��~����D��F]��]/+��4-��T(��L��=�]r|x�մ/��g[�;7�b�*�d@N��Ŧ
؈�8�Z�Y<�p�T�M� ���h��Ƨ3��r�n�{~n��sF��:fU��N�g��%�!7	�<߱.�D.����NY�{�
�2o��x��~�`�6��X���z��TS���M�I5�G7m�KL�f��O�#��Z�bi-(b8_bЯ���k��B�<�DE"�XV���i��e��oP��_=�4��束w�������2\�uo>��ַC~̏�ɐ�h �w�*G$鸈�k�_�E<�>��(����.�w��%�~{e�\3(S�,}0�܏�O81{mˁ?ê�iN����H�G��ߝ��e��(�0O��_���/l�e�`=3��ؒ-���ߌ���`�����#g���K{MH���B*�)����E�17zP;���j	D�uJݨ� ����-kS��;-iT�������9P"���MH���V*g9b��� Q�