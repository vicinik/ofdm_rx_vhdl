��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�E	��ȧ,c��Y��Hߤ�/����Vt���+�q��ӕ���$����#�����W�΄`��g-H���;��Eפ��?)✪��rgƽ�߁���$��[U�-S}��p�p��m�N��/��t��*��|#��aO^%MG1[�{�m�oI�S�3�}�C~�ށ1�
4<��.Y���,��#en���C���Q-'�G����Pw+����xf��Pp[Ș��rB`��#�P�Iƫ�Y�L����z�X 8�Y^�������;��^Q���a@���-̴�J�Wxd5}���ى�\%�ޡ���PBl���l��!{c�����l���Oa���G�����|�8�8�~2�CW����
�B� � Z��#�XC�q�V�
{��R�]a��1�� @��&�6G� 	O���0B?}�p�#97w�n+��#$FD�okM:�$umYL�(�?v�!$�u����.�aΝv���p���k(�T&4Bt)��#�9�#���+bQ%���{2N'h^�\z?IQ$��5���h���x���
����"(կ��ߛk��,�$&����w�ԩ]=Xx��P��Շ��K
gh1^wo�ܯ�'M�Whe���2�x͆�O�g����4��m�u10k?�' 9K���'��T���g�(Ǥ�����a�_ ?>3C,m0��v349ǚ"!��/XF�M ���\��L!�:�����F��.߉q�����I�T�J�%��!�Q�b~��ɫ��� n_��N�j6h{5;�o�pv��3A�XJB�p�~�|T���c���$S,&&0g�D��fDl��x�v�ZV�(T=YNBEs��/3�`a9���=��5Ý�*����?�4'ELx�>,��R8���\�xѣ�G��]�:7 ���c�;5rd�NP�kD�m����Ը5A����F����	�
(�eb��@����l!i"G�_4
�ۋ�cY���yےi/

'u<�Rx.�m���Ǩ[��5�Y߳Ym�^3�:8xy����5�B�zx֜�r������*u��86�e�F�j�R����R�Z��C,eӦ�M�hz��=���zu���>��@��=&����0�(=�!"�3��Ooo����Ak��?�=�C�y�qзj!�>r�f\7nc�`狙~�1oxE�lO����:mV�9j1q�7�\��)�v�]��+J�1�"����ڣҢC�,I,f � YTj�W����,Lu�uz�O����΀P`�pYơ(��O��~�S���
�%(Q,�o������:Y�H��iLUO�9��&�m�����v���y�w��ӄ�/�i���`�,���.ȱԻ^Tg��l�^���_fґX̛^��N+�h|зp��f�FI{ڊ���>�ɼ�Q�|)q~/�����O����m��=�l����.����{f`�T�H���OpX��5|�*�˜��f�]�y��,�a5{�ɷ��e����>�n�%Nz]��l������(�b��H�u�s��0J;|��˷C�!�����is��,_`ϛ��{�g,3\\�\7��`>Fβ� N�3°�o}m]]R�w\e�)���H�Pͬ�V��Y��M�>j������S�� Nc�M���96Pj+C��u`�|�}����Ii��Rn�oV��Hΰ�xH��<����u�JU��n�bξ;��SH���D`���;6�3��ü�w�/\��>�8Ud���&��g���c���gCkN���3`�۩<���Q��@f�E�R��8_(�z�0���]:O[-��6;�.�^��v�ԗ�ʋæVMb����y���������Cm�ZO� �0{	�܄M�x߆�r��}�ee���@�Ĭ�9���G�6��vc���kEA�wb��fc:i6L�$i�Z,U�3^{@1���9�]b������_ģ̕�������k�^�	p^2��T��l:�H�0��ݲ���q�ֻ�濙��n`���{���H���p�5 ].���A�w�F�ֱ>�V�kj�0YnO��o1�z�C>Ъ��K�;�~�%��$1�Io"�eR"�u����b����Ó�&7��dD����<d� �&c���|/`��(E�2;7�54j:<X�J�!��k@D$��X�	=�����%��#�d��q!>vg����$�N"i{��E�=�o�h�^��z�M�^�B*��r:u��U+A^8j�@�pL��B�|Z�#g͟�ڥM���1M����.��7`�d�	��Ee�q�C<�\�(;#�fÔ�z���vh)����y����	r:�:�B�b%n��)�&9��Ů,�w��m�D��P\F��]�zK �L1�/#QGs����U;?6Ա�'�9P`o]��B�$=�ce���Ӷi{~t����k�p��?b�1	�����?��@:!ݓ:z(Q�$�~am�Y�H���xP�Ac��F�'����e����0�H��Q��:a�-�;��s+���D��)P$��a�`�,g���G�E�G�j�W���A�DRޏ�p�i��'�1��$B~XY�X������9��6n� 6��GRz*�~�px��u�( cTMq�%�Q9ݳ�9�*��ƽ��3�`����I����i�yb�I9�uuN�ƈgT2c��u�?��� �����UU���tay��vm~F���FJ4�2yQ��Q�3J���%�+�G��2M0����	�o*�z�
���$���n�Y$���MU�wk�;��?���8J�E�8�S?�~�kן�3���]��@̡uVp;�N�f����feW�Gb�w��`�w�5\��Ho���� /�ˠ�p�tkҥb���D��B�0�Rd�&�K�X��{)Ȼ���$� +c΅���ץ�B�9'�87�Я� O��"��P��잌dp88�֚���wn\�|̾��2����-���l�ƣ2��Av���kB'����Rl�F��@~�5(m(�#̧�Uߗ�2M����Gj��/m����o�����?��Ҋ�D�ύ��P�G1�g#�f
^^�0ߩ���
���E�{�ҧ��HV"���f�ʶn狼h���BZ�1����{�6�"ۀ����������黶�L�������<��4�^-�l���Ap��A;�G�Ps�RN\�ֳ2s��@zI�AɾoW��jJ��q��0����/Ќ	��R�8�ga��.$�q;~��ھ�?>��+�#fC��t�Ӡl1|���R��=A�P�����q�q��Uv�F�#1��}Z�NeVن�I��O�EN�&�5S	0�_��C����%�[�q�^�(w�;Eb���фA�`�bk�Lߢ���a�w�eJ�_�4^W<���{q�vڭ�>Eְ1���"����&�U�y��4�{U�F��a��r�NcM��7ǬW$���6�y�>�Iµ?��C� 6�|�a��P3]�O����3bI%��;�*|֑[[��ZY�)N��B�\�Y�c���g�%��-�l�J+���ش[rʻ2t	�bNF�}y�J��
ܯ�Ո��Hv��� �t�1�8��|� ����_1T9$pz��'J�b|��� -|{��Q'�2��i6����yoo���������5"������E8�	bqe�
l5��~�޸�X�`*��T�d���=Fвr���2Q��h��]���NF���bӎ�o�k�S��x[�I9N0�7��'��`*$���3Ax�O�an�2L���|*���͈ss����0	"�W3;L�~���b�d�;�Ħ��1�P����U�".;�H��o4�}{
����[�A/��C�&�s�Е�\�����\|�,�t-x��@}t�b�� �v��w]փ��jXՉb�
q@x��(��ؾr��݈�9k\ۺu73jXr���"X�����H�85��
M������t.�G�D"[d8�!^�k>��Vڪ�_�:"�)	O̺B�&$� P:��ꉦ7��|�lͩ5���k�N��s	�a���]��NF�,��!Y� �L���|��G���B��ѓ@�;ϸ�\4zTc���Z�P˥��֊p�av���#Id�6��thdULo}.�!��P)��>c��¿��%?h�)�ˍ��@fI�Ou�]Eh�\,�������E��hR;]B-GiJ,�r�!����QW��Gm�JQ�)�o�� �u��:����>4�|���r�9G�d�����fv�l�]@TlΝ�I�5Vl���+�k�y�h
h�Ҷ��}�4�j�"�y����2B�X�d�UT"qF����R2�����BN�aZӜm�7�H*4�|����<�|���8������cݷy���>�m�;���>([�9V�9��O�rY�i
��F8�.�?+(?86���Y����y�|-�y���{���� R�t����+���b��T*�2����Q�������V+2sњ�:�X�z��U�y��U���e�����;�ל�Q��g%	Q:x�>��lJdr)r���Kh���iz�J�_�h�S��E(��|�Iq�'��l�� L�v�ܺ�H���o����8��"�kL]ʽq�J�~�\�-�Z�>�'��{gW�g�ehctJf��N���F;��{�ݶ �K5=��a�y�.T�1_�q��!';���#�V���A��d����d�7���v@�g׸7�p��U邏��o�-�=L}$�{oͣ�
mP�㰌�4�;A�4�嗓��5�2b	�Y^P�X����;{b`�X�6�S�c�T��<р~�!4P�h���4#ц�aC�f�zW�ɬ�ἂ����	�[%��3�T�yN��a�����|�dh�������&� ���� Y�	k���Z�e�����cA�59�B0Z�w?a�ˍ֔��#�a�����+�v%,ϙ3���w�u]�ɟ��7���ڛH��}���e`y)��^<gBU�;���f*#a����.����`e�ҧ�qa��Ֆsk��zvC�[v�m'AW3{y�Kff���V�k3d��K(�w�[d`AC!Rܧ�� ^�ݿ�y_�}���o:W$u��(�B���?�[Îi�\ї'��_�j� �� T!}���ɀ)��0Ќ�(�(g _�c:�f�r����4�Q������\�>����{�Ԉ?�e�q#]��M�֕o������g5�7^â��c.c� k�_�Cg��ک�}���C���g�9/,N㊝V�R#�e��j3բ�-3@K
(����g�~P�aȰO��Ms �)���Y4?�;E����Ӫk\������T�� ;S��A/4��F_�"���\�~�"��6���Wq��]L?IS��Ѩ��� �i(%e�V�z&�ί��"��@zFH��y��h�G']U�t<����R�#h�J'����m�b.>�="����h\H>kjAa�	&X�D�挠WX��G �&Pש�t(tp6%+��Q��C\�}����;��dn"l�9���� ����h�ơӃMpmT.��[�cB��:�b�
2����v�A�����܇4�ck �Xm�fN���s��b�¿F/���k�ݭJH9����Q�B�<�u`�U�F(g]7�U��;��9X48���[��7'��=6�#GU����r����cD��Ӝ��#;Œꔘ��=d�mZW���f�������R���7��B�ŷ���:f}6䫉�}X��R��}L�8�t��@!�@��ס�Yx��fQ�Oс��9'rюm�n�uY��7����g��֌;����.���|�c��B�;&x����e�Ǔ���'7�$�0���� � �Ǫ�Y�l�҇�o0��+��lko�굓!f����-5(�3��} ��sI�����[�-���.�&�����  ��]�)v�1RR!���Փ�������_w�J*���QLi�q�6V�l�5*�p%�7M���桂�s���L�_�@�������`x-�N0F\f�AD�RE��K������D�k�C�[���[T�f6��w���o�9��<a����0�ş~�\Ƕ0uI:w�P������OU@��^�I1_�]#�8�ٝ�(�Ϳ��=���fԚ�A}QB_$!%�;�G�����g��HJm�z�T�/�J��ϙHmoFA{Ϫ�P�Ǒ��,��h�_����b
L̈����b�@D*-����?Q��i������C}وiٺ�xsӑ	p���C㧇�r����K�)+n�u�w#>�v�f���.a߻��\"���o�0�DQ�D� �?E}���p�ml�{�Z�8>�RЮ;~R}�m?����������ߺHj�<���ٍ��� ����Ę�� x)�c6�-@Q��z�Y|4�A�(�R,-3s�}�c�^ۦ��K��wpG�q�g7҉OU���n��E;Ѝ������<ж1|!�wիb��_�����7RB����NF:7�	�_�Op;��d��̮�sW�.���5�c)����TU��)I�~�s��8���W磩�wtc����2�)�;��4X��O[ԉ�h!(ϺF����$X$	*�8�;ĜD�:�������a�y�Fn{pW����B�:td�>��l�2&	�dUk��F��7�˝����k^CI�<��~b�����V�w4�/D��˲s%��T��2�ϑ�-�n�ʦY�}��ِ^��������<�~Kov�<�t����.l���<����`QE]���E��M�����g�ȟ�xg���R������oR�Th=/=��W�h1x�)�l)8_�Z�W�`���N�qZ|�;�����u��o�M��@�PGSHb�.߫e
e�s��/Ջ%"����SJ���4�ĐR/���%m������I|w��w�	K๾}��`�z'$�Q�؀�[�1܆�Ħ��<�Y��x�m4o�"���>�X��1�<��Et�Ut�n�[?E�M_���ܚ�|[;��Q
�J�`�	K���-ڞ�Q8$�?�60z5H&w*o#3�uǇ�Q6�L����r��+�8�;S�ڷ����s%�t������̽��Y��(�y�4���.�_h�~��jM�?px`7�4θ[d��F��WЂ� �4���k��%djJ7�*�����G�'��ɉ����\�ܶ;������\7d�N�Oa:��^n��Zu�*}V�_��Z)�2�3�k) �vq#���I��D���K89��$+SB��u�}���zӸ{���#lmإ�;�%���Pn��:s��%�C(ܳ�()��!-� �h�Om[^9�1�N��ֶ��0�F�����.�9���;�=3Wױ�ʎ�1J_Si���З�散2�x�F8s�yoL��W6��i"�p.��|������m����tju4L�j�����@���0b��ٶ-Y�E:@�U�t���^z��DR�<wh�؜QS�Q�6]���f�kC���WA8+��Q1ᖕC���-0�m�]�ؖx7\eWd�H��X���'��/���E��՛z���ə4�C�:c�ƐŊ��`$��.�{�a��:0�A=�������b���/���MK!1�؛;����(�Z�Uf�t��V�,J�b4ٿ��6N�B��~�[��'���	 �5H��G�'���w����w���S��^AF����LS6�EQơ�����AT�gg^����X6Xp�d���1H���{hz��&(�L�Ǭ7h��"���OuV�k�$�� �M��mn�&m�����U�n	�Ȫ�ة�ْs�%��kk���c�U0�� =�c�.����!��%Su}��j��t9av���y�"����O<RG�%�=S�D�
a��6�#`D��`$��5aE��D�(��{0@Kz�k�ɞ�ǦUP]Y���Xxs���1~a<&����^�~��<ҝ�������ۜ�Y�Q����/xG���$Ks��@�,0����rf����H�@ٿ�@
� ȑ�&�I�Jǥ��PE�P%o��pT���m�"%���1.�7�:���}���`+i4o�����?0�k�d\�:5����î�<C��E������z�.���r�o�A3<�+3�I�z	Ms�ƎD�'����V=��!�F�@~���<{�a�����2z��Td��O-O�%��}yia��]Á��脊WC!6��&S�����Ce�3�����y�y,�1خaH[6����vY��N!v��6�����SqWGp6�Z�g�e�=��C�+[�M��4�R���7�|y����@����ejW�6_pZ���5�<�L����3JQ� �F��}��vZ��XdCu@rqt�6��!������@�V�H\�h�ZG�8Q#p�	�G1�Ҝ���#�FQ�q��������|԰}n�k!Z+k�p��uqxi(ӭ��1���W��:YԺ���9�Ntn��(<������E�V�	9@�����NJ=tn��M�-*Y�<0���,�b`�J����VgäE����6׆/b���&'��_����}
�3�ێ�i�#�F8��1A� %"yݟ^�/�}d�c��	��Շ��M�|=8�l9�{ w('9̜�,1��ߙV¦`p�R�aO"�بX��59���\�R��y�;������u�����g�8߅�?���^ {�20�����,Ny��R4_`��3GhZ��y����#���4��Z����a�)��n�_!h��ثA����.̓�qk�p�a���ԭ�}���H�Qғw�#Ol�����]��3x-=��d��WHN����;ᶷY��I��D��ɸ�oyai�쾬Ȯ۩�!&g\�1��jW.��Q�N���v���H��]�iP#� H�ID��M9��K;EJѱ�d�u�v����������
��G�=�q5�騎8�oF������{��~��ϋ`��/�XT*�쳀�g��--���������V %�t���]�J��Y<�W�s�!r~�}�
���$B�Gp�8�}�E�x'Q1�G��Ya�n�7I�P!5ݜ|Ҹ>)���?��)���؁��� ���:e?�F�:o����q<�<�N��&�l��aC��jo�
'�z�	�\�z�M��sBr)�ǅm�cOt&�eT�pf�Z&b�C��Rh:��<��7=�7Bn�kD�9�Q� }�,�r�F������ɬ!�?+�x!�8.J4�b�"G���;W���E���J�๟0&בE(P�`[¼�4��$4߽�J���77�ǐ�����닩�Z� �����=���74t.�/#I<6;��w��N`j�Pd�-�ƣĈ�B�sKc���I��\%���)� �w����V��)�֊�9d�����I1����^3�O�B�:E�<�b��8%N�{|m�Xͳ1��8Ϫ��w�"[;bB"�\'�o��O�t�x����'j72���j�p�7X�k����_�=����%7��[��������.A�Lى"HӖ#{=�������C��f��^	�"��N�X_Y��8=� ���у�b���O�$�!��U��g�Y�7.��K�WV�?��D�?j{&`X�e2U��u��r%��٘�r��H�L^�v�Y�Fok̊�%h	E���X���9�V1!>A��Q��mIfT�m�-��Bʌ7]㉪,� �s���lOT�'`��fc��W��M�;�*@��ZF���u��_�)�2���{�r=P�E�hk����o �U���W2���Vb���:���YC�}�SP�x�����諃RC�-��Wh��ۼ�6<`.�'B��S�I��c�+K�����pL	��}�Q��-O���e�M*O�Qb0+8��t�;���?#�I����	Dx'Գ�+F��
�];� ��g�/���>�vߠBz�g���Y�hs���d�~Τ�!�?esJ����p"��F�����J���JJ�+_'@c*�Faj[���n~�G���K�F��u�UQ�����6]��y��=�4�'�"Ajp����f�6�W9�:�����LW��f���gԭ�ѡ�x�>t���i��fzҡ�?����Q	����⩗-��˧Y1��զ����ez��#��xV�9j[h����v��������~5��΂Q�F�\svn?�������6��-}r�M�%�5cx݄t�'�-�����[��=���
Y�B+[lG��t���ZlW7J|"){hO���~�D�,���M�K�z�a���w�A(�[`9�MБ��7���&f�s�.��A�C1F/���N�8Y�0u6����Yj�<3 k���-hqG%��U�'���Z�0�QAh�N�ޢ�����o#{����T��)�.[��g�`L�a%�/�ށ��D�R����7�c1�)��t����f-0��C����R �+�t�%������������UR�ƃ�G��S|Q��}�e�+y�I�.GS�M{�9�2z�r�\UÐ�j��3V9�-}�?�%�tۿE��`͉nne��ҙ�"�G�,x�;�	�ż�I����+˳nbkc�U���-B'0S��n��+���T}���~�<U��;��x�����v�5�4�N���ф�3m-FN�9�x��Na}0��c}ڊ �������Fǅ��m}�_������6I5T� ���\[������[�s�M	��9�[���:m�?la��}>�a�[{�ZB���W�$��X�7��>�#w�j��'ϙ�4JwbloH�6��%x��p�y4�����`��b�Iۆɣ���4�c�]���Ό��ڈ���`0����3�:N���Jn�r�ꖣE��:3B��v]S{�'��@���9��Kh���-]�5��v����O�fy�5���N.8'3���=�Gx�kT�MN�I_��8��c��:�e���ӥ�^E�L��@�-~ʌ�dܕ�|5uTKffK�`+мN��Hn�"�e6��M\M��V�Ž`��Ǵ�P����M�.PӒ�uZw&���w��I�C<zu�t��Aȇ�v�4�Q�S�������p�Rg�M;�kW�pP�u�ch���L�0z���� �H
:;��vS��އp��#� <�� �j@��H������U7-�����sk���l'If���Q�iۚ�I����@RF�聳�Q"��I�f����ߜh��Pq�V`��b���@ǟ����.�����[T���-:t#���a���Ȉ���0X+��	Q����[aN�Mm{����]�Qe�������<A�@�V�C��7l�� ��x�S3{iH��Y�Cc�R�I)v�F�&e�V�J��仺�4q��Ph{E
�_�y��A���I�%���ɀ�ӳ�ðV%���{I��9�8i�3�"^P�C@ߠ�(><t'vKD��"xW��p�RL:�ƹ_�'����Gx��H��񑵽�`I%�N�ԏ����PG �3�ai��Oe����ʉ|��=Xl���jڒ5
5[��I�q�JZ��v��$���-_W��MM[�8�l��lt�T(d���*�%2��_j%�j�i�	��)N{P�%�-cٲ�AR؅M��5Ǩ��R�����JI����c[}���4�'��dⵚ%��l����KU�� |x�=A���7�2�n"*k����U��eC,%����co'�$�����C��S��ك�bv�/�h ��,��ʫ���d~8��u=��S|�)B��#�������cL���ߖʟ�:����#^}N��ʣɺYf�t��A������������Ku��A �٥����0{���\�P�S����W��A�"_1(�a� ��R��0�[p+��l]5%��)(=�r���j&�A�wZ��<���,�E�=C;�mvR}�h
��5�"IQ�T�4W�'�$#�����~���?p4�򍓰-%��i��y
�-�kM�|�6Z��[C$ӳ\���� �u8��j�\��K<� ��#�6�t{�k_`��en o����AgW7�v]m�1��|��ܡNA���%$��N��q'k��8��G��y��<^�p	��g)}����ǆBJ���������e雳=�h� .`�D�h����t[�}�w��޾���"�����R{m�іp���"\�^V�:���3TS�-��)e��-�8k�Л��DK�[�1�B�U�]h�������98�jp֍??���RRq���´��]�L�-v�0PW��5�2�rsr���Ƥ��W���~�����	��q�2��K�	z0JeL���?���"�1/���g�� �͂�D�<�J��!�е�-3�8�VɜؗW]=>J��콎>���}z�	����ۊ,D��'��i�D��|gm�sj!S��`�M����Y�7��N2N�(C<g�"�5�\�$���������_��;Xu��CS���>s�Ʃu�LC��]e���|(_�'k��e�z��կ-�=Q'p���N=K:kD��]ۜ���0����� �(j�� �wn�ⵌ����U�O���VPkC��� ���j]�*z�A����܆��[�ȘK�Qu&4�e�'��w
�iƘ#]�?�%��#@ߩ*]ż8(3y��^�31�>��B���Y�ge�rga�N'q+7���fp����iwK��M�[W�U%��,�����P�.˽��E��baL���{{�l�>��4��X�"X�*��a=/�V|��@y1��@s�Gفp���>U���k��S��s$gg�$_�2������
"- X$�bA�e��>|�z�1oΊ��S��=E`��͊�1C�j���G�?<�L��	�Ìg�{[��Ť���2�4ZOȖ�NS�g+z����͟~"�O�U���Od	���3; �C�Zɺ$��{�"'�$� /␄��'m�"^t�<�s���Z��mٹ�U�d��؁)�OU��Z�}o�&&�c�b�ś{�~=6m��Cl��^��'��� n���P��w���
��V^�ْ��VR�B5�"kݬ �̉ �:�p�����Ԛ)�w�}a�fK���='�K'V�oʋā�ڶ{��;��^�
m�X��.�W�v�E(!{����������쥞��u:�T|���G���\η93H9UX-�$��M�a�{̩�)aZ�����u��z{�����Y�����:rD��k$�D֜3�X�"k[-�n������r<p�R�=C)��y����)�}hO�3��5 "K����]#�(^�ƶL~���X`yr!G�c�#�N��0���o>�[�c�Ff���ۦ��R@2�LY!�ͧa'�]Ŭ~M�1B�S}�U�^_v�VSz2����LG����y�%�m�� �j�y�-f�9j��d�r(��&b����:��F$z�

�i���Hi����l��?�^��g����#z�\��@�.|��2�4ܘs����Yɜ8�BE�����z������'{2�i�XD�,��":���X�,�:֘�]&�E�n��ȓ�bV>]���wd�x�ct�6�XZ.b����"�@(������yҀC��N����"�|,�{�� _9g���~_�Є����0�����D��}���y�O�|�_#Q��\"�����yx���I"�`�Kq:P�=�JK�����>*$�(����v��ZǊ�䐰U�e�:�	�o��/�T��Q6L��V9ZjE��7L��[��6ۓ�]���w��p\�� ���]G��s�R�:���K:]�Z�K��+\�Z���xg�R8A-��Qm�&B��z�+a��E$�l�u��(9�1䣼F�ۮ�x���;P_A;�@FqLZ8�L�eߴV�΂ڧ�Yo��i��p;Ž�M��HB��`�7��#n2�����f_&3���1�u;y�� e����5��H�!I�G�
M�2��쮔#�-�1�zI��7���a)��M�L׾>�5f&ܘyP;�������;f�f	Y߾��l�ĉ��_]���/aȜl�]h_�k���T���>��P�w�HS � wuF|��C���֪�m�Ci����3sKǱ����-I)��T��Z_$u#`O��f�`z����W!����a9O�l�V��@�������ϲ`�K�z��J������C�3����BC;)g_����� X+�p�Sh�4�Iu�E$�Z�l�F&h��-
�(0�"r��#}��f�oxdǁج�Q�<���LK_�������D3I���Oa�N=��+H�Ӧ�f��H0�$o4����7�kE���rx��e8#	�a�N[�f{�
��q�.��C�-���Ő(�}�(��M���#eꈳޡs0�4�"�҉b�¿Zr$r:�Y�����w��@cE�̪ʘ�q��詛���PqWR���V@�71���H�A���<�p�E� ���48��
�r�	+.&i?�h5j9⼴����߰�H�)�H�� B}�9}�G�%G���*�K�T�9�!����Y@a��y�n�:8�YڑC(ӵ�8�GJðB�pk��7)%9}�!��G�[�X,��3�Ȁ�.��5A��G��P�1<x��S`5�k��v�h�������>������$t��<M忍z\r��P�9���MV�ӻ�{G@'Y�Ōy_�8<ð}BS{M�.����}�����Z�k���~��c��)�H֣Z傯0f�@ŧl-K��xH�m؅�v�a,ֻ�9�A��m?{]��&�|��8F�⧈r7��I�/��?�	��=_U_h��_2_�����Ӟ�8MX~�lP G��q�����^��������9{�'΁�w�0X�y�i�n�������������a��2"os��`�Y^�i��S5� �B���n�QL�^�8��#��r+�9�V���9�a�����-7���j=����$*��,N6 z�\3��b��(i�s/�@5������XO��̬���1��U3��X��X�K8><��6>jҾ�Y�Æ����/�,�˝�/�w*��5�=�~�OcK�(]o�,s6�z�T���R�3mJ�pH�7�BKNq\#�%�yp�,̏7����.ګ ,K��KS7�Eĕ�/���G�#�5y�P���AJF��(N�j�$E�F�7iZKQ��<���`}�b��3P&�Z/��3�r+��O{�F��0PK�#� w�䵈�G-r�Q:��;��ǤFg�J��<N"���5좫"����}&,O4T�۶�0IFؙͰ�m�|�0�h�:7�X�[y߾�p���X�e�؋^��<v�FM�<$��)	Ժ-z��n�M�'���t�2jT���������DW\�g��+ �@V�~Zt�x=�}��x]�.]�[�qc{�#2~����
N�6�vq@�����G�7�ԃ�.��~3!����'r �h�*l����N�E��Ȝ��n	%Ε��2w	�N`q�E�� �(j�f�F�GO�b?T���%r�0�u�dO;���}B�0�c�w(�n~ʵuo���YF&�Z��g#��.J�x�Ŝ^(`���5�y?2ڎ�J5�A�n���S�n�ф�z�L�K`�T=@�:���R��х�]�wa��e:t��@۶KO,�3�z}}S	�]�Y=�h�����3x��R��B@���O5�פT*~T����,M�G)`�Bl7PT��D~h��d�ն���,ǆM���꿡|5?k�m[���r�я$�kX�q�mxz��!�p4�H,NgV:����8��ǖ���Z���"�f0g�*��hO� ����	�3:�C�8�H���{�ŧa�T%�kY �'Rj!E�96 ��b�K:����%<0)m�?�m�YnM:C�|7��K�0Z�a������2D���ڮ<���-�S�Z�V]-٤FEiW+O@#_�k
w��q�f�[~]ŗE���k5>�;.=}�АL<���O��_�����h��HV{[�knG�ww1��1���{�����B4��~;���
Pk����s��'�i_�*.7gT���J��3��R��	q��3��&��C��J�Q�cÃ�C�+XDw��Yf}�;.�<5��*�n��b��O�!b���Z`�a��_ �e�6����:�ln%����M�6�T�{�r���B���(�����k��cO��iqVtk�:V�����[��� 7����}F��?t�{��� �����/%H�m����8�_-@]q7
�%���|�6�wkgb�0�d�J���$��Fl�jOи�:�%�E����!Bw�K�Rw�L��'�o��y7Գ���88M�����l����س�6ĊL���w��-�J��VgX�p]ǵD��R�;�zi	�Rf��B��ꌐ��<tT��3s�x�g��tڦb��P���u���䓞
��p����ྖ�I5n��?��M��8���%Jv�xHa��8�]�ay�vi�O���� ��^��߅d=`�a$�s��'q<.�)�q�D�"�"{�a��m�V^�K���0�)F���x��2RS]Vs-��\)if0`ie�h)��1%*=O� l��b������J����b����V6�wa. �Z�����'�Z�x��d��Ӂ�)Z��}��ތz����N�5>~�5��[�Ov7K��Rn�xO�~�F����Q��yU�w���G��}�� �]����u��2JS�a y�K��㾋y��c|1B�,�<�D$	�ws��h�'�-���%K�y�Dn?>�I��R���*E�3e����5J����a�K3~�{*��J3ؓ�GbY:�`�����-6�j27��>D.��}������-�*� -�-߉�1YZ�NS�ԤxMՖ	�m�'��Jcm�?�Xy�9d�#n�nɗ?���fs�!����ffɊ��Z"������h�[�]4h���
9���2��m�#|�3��L����~;��jl�c'�#���{)���3XF��t���o��l�}���x@��2�M�E��m?��zb]l�g���^v��%V�R���G���"�IߐtrI!ݮc��
�ŷ���| mI�����ԍ��~�2��Jc�|��4!c�n����	���h���zPc�&*rTǉ��UN���
Ꮞ$+"莿g"݈<���� A[�5��w���s2��"	���'% ;������2e��؃��@��V��U$�d�Ur!_��F���2:�r�a�Xt�P4�Hp��k�r��z��Dӓ��@�5�֞|���᤾�)m��P�S�xW��YG����}E�ۚ	P �b�/Kj��8��)R=h8�WD�H.;/u}ށ���\K^
ŉj�h�8!U�7��I��R�`3}'��	�1vw��L��6�x�KE�2����+�E0�$��ua�"/�	�#(�Ϭ7ߒ�-�Z&-k�Ia*�`������
�SF|���p�
�~�Q&���&�(KI�^�����	kl��z�<Ũ�����ʳ�����y荄gXQ�g^��~	~6�Y�N�������`���p�������W��EӾm�(zt���%� ͈�%wo�~��n~�
&EN���7/�|����,�8��{lS�_�V����Ga�g �mY����]�~����fX]Kn��5���3�EE���'H��FP���os���˗ [���,t����d�����S�45�&�Ul��
�v0����Xl�����+L?�-��b6���ֹ�@���Pv�2�c����c���/�J �pV�,��h/'��V��ȨyI���<�KhO���o(��^�����l^%��w�l�LA��CYn6�?��qȀ��ED_���m��4����M�L�p���ff�&!�܉<�ōgjG3K�xs�Y!;�ԫe�%؝U`�
�g��鴐�5h�]��b�+F?ԛ�:B�)c<)c��)�>|�f��o��HH��xa� �ڥ���3�������5�#�8��a�f&/������=��'�R����$6uI��K�lPՒ�������q5xeL4/��Jh��,�ll>?{g�H���`ƾ��
���;�qg"�y*PM�m�j�.-�����B6�++zeCϽ�C���We���8v�y�mL9���!�	�@p���9e����k��G�2-�Em��9��V	����*m�]j���{�m�[}���� NxM���*����Τ����n���H�Q��n+�Fx����j��I��3~��o�ھ�I�}ؙ�Ő�Aٟ��,ژ»S�����_$ʵE̼���Gk��W�S8��޿��5�ޯ�ߞ(!@�}��ٛBT"Ø����1�����;x�*ӹ�x1@��f���e"���AC3�W�-�j���� �ӟk:�Vݥ>�]g3YOP)����PkPYyC����8�o8#�8K�ʺ��V,r!'.�]=��������*!6@F�d�>�A�c�\NF�����E�)��P=e�0��/��0�Ч
��(2��Y�����X�x�&n��=?2�%E>�S��!j�������y�X�@[��t��o����=����k���g9.W�O��i7�����d��z�@���3�E�v���U��:Y�K����p�q�%���(�7���5�����tu ��PUnt��ֈr�����r��@����K��&ս!S�t��(r`����[�$�V��Yq�*���m{�5�%y��8ƪa&��g`j7.+�qʪ�a���\!ƇZ�q��9���:9�/:����VO���}#���!��
;T�I���0sy\������C�Ws�X|�]�j�]�^�\�^[�N�Ԥ���&�H��)��PX�Nsm�6A���!e.���D7���E*���[�)���&}�
3�2j'l�
�k��Vp�%+t�x�� ��0�eVġ7��g�����\��/�>l9��o�.�Q��y���@����q �AY���M���AX�v��-,`�E�\�4��R��f��(X<mv�8F_k�H�W頖�+8�HB��U�����q�Љw�T{�r��Ȍ%~W���ar�=ęf� ���I���fR��D�攽��oXr'Պ����3%��~�������}�4��~��Q"��c׍�9͛��(��+�_=�ͧ�V�K��^���J��8i'ˢ����^��L��k0ت�Ob	w���gn�"@W?�p<�<M4� �-b���Et��X��S��|�A�\f���Ȝ~�(�kG�RY\sُy�[����ɺ�Q� �`vU����)�T:�X��&==�ń�a�J�� I���l��P�6��O��=��6?M�t�q�G�,���L�?'+fa��X'�n�5o�������1��G	\�^��_4�[_+�&ߏ��R���FW@�����1V�����)�U=��1��U������j �W�����͗&#�(��Ab)0���@dS�z�q)���J�Q`���@��'SNC������1�$��TH���@�#|�qN��7w�7���M2���H4��'���RhB�0ä�9/�kކ*��*�ԪU��OZN�}�m��/KJ�feEe�$;�z�G�����Ra1��|�Z��pA+�hK��eHߩ��7����,W��@�W�\�ƣ�[�{a�!�o3i9�/l�ͻ}+�%�X����qcN\��#�-g#�ӹ���/�1N;d�'����������hvXdAk9߀>Ϲ$e�����-����rX��k\��c����g۶<F|&�f���;�+�<�?�����t�������_U8��=x� ULϐ��|�k��z�+F����7���&ȣ��kB8ұ�v���Uy�z%�[ɳaj �1J�_V��%��� ���95 ͞�"������.=DG��#�ҳ���MR~�.E��l9��������������4��a�Q0"��_�����9�����u�OI.�ی���MRv���U��R�Fv_��wdz������aC1g���D�T��f�Hh����C�z��W/%�� 뎶�"������`�E]۬Uk:������s�t�t�̂�\��\i�u�6��؄�=���ښ_����e��P�T�F�*)�V��sBv����g�IȕC�vU���<Gnߢ��V�}(�ސ�`�Hm��L��U������@�g#��?U"M7_��.?��QD�r�}�
�ױ��9����.�yȁh6�r�l�)��[ �pQ���8U�團Sl=��i>$!��?]��zq�<�j	���S��S�����F?�c�c��R�6��
���S��mPJ�����7hP����ɽ
�Yv[U���z� �5R�t� �g)􀈯�_�A+:�2���e�e����/A��T�����qN�M"��#U��3<���ز��G�	^��f�-��/�N郾r,-�s�-�Y���Æb�� �,ېN�M������x�YM��<�=���Ƞ��$���b8�]}����<�cƲ�Fq����P�+��L[d�m�wE���'��F7Mlƹ���8:`9R!k[�e_����� �����59T�Eb3���Z�p�FV��A��o
Qf9�S0�Z�Q#��
��Sh�c��󜣯��R����y-�()�@�0��z���P�L�����0`º�9�p�zΊ,iv��Aaw���Y��(_���T�/T�%�T�cUaz��]P�6���X2(�~<��:#a��ߤ��b�"��I{2<&y�h��;�BD�d���$B%mw7�B�v���/�X����'�(VŜr���=�*�tn�plG��d�i��N#���o��9����+u����.;A����~�^	��i݈x�́*�{L�������������5��!w7�XU��@�pO��1�vA�`��$����T=�;�W;���h� -���7�(�J��h��@x�z�A/�M"�-\D&�^�O���he�-�'�3o����PD�:���3Ǳ?�^�������!7�o���D$9���*<a��2��'P��Y+Jx��S�k�̽"l��{I����е��X�Gw@�r��[�$�C۴�N�յ"����YI�H.B|��@��׾��Ǔ��ST!�4�Rn��F�u�4ӓI�l��*�mߊ}AD���>^.Á�����+��C��$3��5���X<�����J��|�?�9�K��
,����̑$Qd2����T��˼�� 2��U���-Lg,����j��ɺ��;����<Fũ�̩C�a��۸���&�o��deȾ��	���af���-��ɦ���� }��L�C��tDlx��tW%�|w9�3'���+����ϣ/�ꚑ�{Jd��}�p�����cm���׌^2�G/�x!l2`�!�P���Dc���O��ƀ��{�0ڒ� a7r�B�0�m��N���Z,(�\����^��7͛N��ؚ���޷ż$$����0�������Mv���E�0Z��MEݔ�7t2�./@!�:��2{�ŭ�%��$�}FO�McU�,���M�ad]}�ty^��V�a��$��>W�gb�����+�90Hr�� �xԹ �/E��M1CL@d���>�,��'z��|�rR�%��6>ڥTR"��[��~���<q륕���8�{<���	�8jݵhE^N<�T��oU
��9pc���h�c�=tX�B�4~��Y@��4���'x�x��A��"�:��cA4�d��ң�M�TZ�s/q2�|1�
�,`�rc�=�w�[���@DP��w�u�p�<�GK
w�ί���N�$�m	#�z�4�{`�0��Wj1��5��[�5;�R�J�4�X���J#�[��#R����v�#���� xQF������%8���DN�ۄ�/[�e�%��������(�uFͺ������D�`,̈́�>�*#B�V��������>N�W�P�a�	�w��VHX� ƞ�IemEF�v�sꇈ.l8�?�����ujv�d)�^U�����)��9�يf��G�D0�8�˥	��S���&�0�Ϗ�y �X_�R@c�0?R��jN�1�����Ů��ds��$��lb���,�P�!5v��#���Up������,�	C}i����^�V���qfMb�#<����o��� ���*���������՞� ���)!KK׏DЮ���ɥ��Y���_�<� ��hjY��£��ԉE�N�-b��Bb��M�"��W)�h�ؙ7�P:���/<���oPԀ_��w�c)��R�I� �S�͊����c��Ħ��'�
��(����=�QƠ����x��ޠ㪽./��5
��{�4㜷�9~*~f=��V~��8qk�sMg�ܒ�<��� ��b�v#��髽|m+�#TE&�
�N�@|4�d?B����F�4����<E�LmS��gc�%��i���}4�0'����FS]z���e�e)���iu�B���cB��Rk�?�и*K�#i�3�R���j��mv6����7��RV�8�ֽ�s����i��4�ne�j�s2Rɣu�C9/��r�r�\ *���=J�q��R�?�)�۾�b�(.��y�H�H��~��L1�P��n����`�Jd�Q&ʕ*t{��͕�)�͎�I�
j��{�`(�jX���U����cﲊp䤒��_��B�~�V{ZO.�q�#n +j�^A���RRM����o�maL�U힁�*��<�]d�Ax7Mn�J�k{u/�u�T�0�ܯ���Z���Fg�c�	 ��*�l���?
�smya�>M���pDa�n
b��Ȩ���ԝ,t��*�tn�L^��@	�+	8�[�Ef�
�ZET6�z���}�?����-�(U������O}���x;�*ᰏ�2��"��,�?�,.��#��s<�|���x��X�@��v�;��E���c�zo����
?�I�5�����0�Օ�pӃ��~U����4�t�Jp�u�Ǚ��1�6��!z�<�uy0�W��mԦ�{nVE�dQUp��ؓ�rT�^���[���i��҆�n�k�ھ����)��?���(Z ���������Y�����6n|nѩ�_ۮa�J�����8�l�D�o�\`ܲI鋫�ə%�݃���}��׃�
�����:!��df�K;��/.�������$�<�"��D	GW��H�r���:�?
����'��]���""@�����faF��k���$3
��=��n��}7��lY��3T#ds�oi��v��S�'�+��S^!^h�^�F�)��0̐�7�m>�xJ��>{O�ǻ+`dz�����O��C?�#���'(��w�P�^;!��׏�)=�"�+��W��
=Z~ z� [����-W�?�&2� gP"*ѹ��3�;�D~�@�璄r��^��D��*I�t�,.��ě[ͥ�z^PO�}C�v��@�55�����Pֶ�h CVF�v9�^l�	���0օ�ӻʩ�l} }lw+��i�]E9,�����3�R�Zs�)d��qD )���r�,��d)���8����1b�����?�/��?5�c���������%��:%/������j���g��������-�[�A���RU�����b�p����Ɵ�3w��q�W�O�A{�{��*Ź��a��Ba7tm�Z@���]������7�����j����IR@�Ӳ�a/��n����P���V��z�DZ4���Ėa�����Gno��c��f(���YW��v�s-��W=�tbi�,ݭIt�^�/Gn{�g������}4-炢��a�wq�@2dL&Ĥ��ࣺp~*ݿ�ů5;��5����$�V��^jY��k����$�V�Y1�+e��L4|CX}M��O%�S�Ȃ;ڝ�������]��BR>�"(7�G;�\�_=$l���}%({�Y�#&�޻3m��=�y�9� �'w�(���8�@&�eW��ݼ��\��]򚕁*�L�%aԴ�jf{q����d��>���m(}�h9��g��x*�"�M�G���*r1�� ��W~�6rO<k��/���z0QT8i���ïO�gy����jͺ��(�Jn5���+�<�xYU��-�����3��?s(U�˜�d�c����oD�R����?1*V練�e�.��Q��N�7YUv��X�j�����ʯg�B�}�M�������M��01��M?{e�(U^1Q宝O��oS�	[��m�:��NW#j3���Yķ�f��^��K����q�
#"�iQ9 éw�N�Ps�R���ݢ�nP�����Hƍ)���i���W��Z�P�)�jcJ�N��M�G�+���4#���p��Ͼ����s���עĀV�l`�s�W����U��U>�z$��լ��C��'����Z������k:�Z���=��F��=S��d�pČ���C���wZn�g�R�.���Ӗ��&�,v7Y�f�{��#�� 1�J��x��<hr��$�N��L#ؼ����.�G��H�|�JD[�,'3d�h�\q����!���q��$��f@��f��gOSN�V��V��R��o��\�T�����H�5�xs�Ȑ�-G_�z��I\��z2v�i�8���)'��*n{�_��,1���# �zz0�z�HXI�+���ff\�ƹ|�.�h�?�:�M5���QJ�k�w��LV��ޅ���иR��Vъ|�[���N�sRɏ����/8%��ȩ5�MZ�{}�bl�YWӑ_���V������)>�G@�
��S�6���%X��m��#פ��pc
mKk��4�L�'�G��w9�k��|p�S���H2R24b .��c��X��>td�$�2&�O0�r�$	$�0�^Q��P���r��=�>8	6IJG��N�D�d%�È���gt��Ѧ��$�\����_ӏ��m�f�����:|޼��B��BT+t�_�����,�ժ����r�r�"/�
i�\���/z�*{*��Dfm`���	�d&�v���1"|�T�ߩ�QeE��poG�m#�XaZ�Z�����Q��PpK��E���9���Vg��a�zm���=�Ԋ��6����m�,���օ������O��v�s�"��S�>��d�XV��x�7�U!H �@4L^S+ya.Ą�VR-��(Ryd�rBd�jFu�V�s�9i�A8��&�J�a���R% t�:���B�Vr�tí��YK���(�)���*>��o��*��`�d�#���5yD*�Ёm.� ��-��@`���S���V�����My�dLG�JF��b�u��"3=����VG�,�ݎ���S���y^eG�B�"�(a�~��v|��� ���+Ni�W��n������RJ���+�:.-���FU��񕸫y���9��YC���%$C>�wE��v��$O�pY�6�0q{Ay[[|a��5rDr5;+#����M.l��
��9��`n/��J  �G�����H��p����\=7f3)�r�W���w������$��|��[�(���"Zp_u�nJ:S��ٛ��o!	V��좫�`�{+`r���E�صeFپ��mK�ؕ[�]Cݮ��&��|�e��!����Ƅg��"yϬh���e��m]/nF�����4���lr>��Ӹ��I���]�� 9�����A���f�@|܂��{�S�z��C�y8��1���_bN�άcXm/�V0��F��aZI��}I�^�ک�C����eÖG8�֦ۆ���l��ŷ��؀
���qX��*$�<F�as	��J��CX�V�v�<5����<~b�Ȥx�XLA�VVʮG��\[~�j��8�|LT�^���#J|�!O���D��ԅ][?F�y��x<��۱{�-Z��;�l�=d<����H�Zf��(݁_������k�&@�J��4q7�t�N)�,�Td�d��8#29C�[}��-L��o��6��2��^���m�,��8֌4w^#fC�d�SY���p�b��Jd����y';�S���ql�|63ͷ� 庝>YJ�����8Q�[Ȃ|�G��6J�jSZi/�	�x#��|J��tX�`U�؛�������C��F�3�c�����9ނE�P�FS��s�H�8��;L�{]���42�ؽ�"<^�C��!�f�r�����1�֌£Y�gSXv	�N����u��&uqw���1��l�e�#n!��	���q�K2�8%�Ȩ�ʑP�MnE��X��	'�^,V�s�ыR�������p�}��!D@����0�D�����q��t^7�Q⧵�i�6Ղ��/r���N@�Ҳ�扂��s�(I�{�y��������_Kг��@|*��f�l��wv�6���Y��7�F���Y�mj	[��������z�Ԁ�_��D*}�<Ʌ+���GūO/�]���9�C~%�1C��� (h-5\�qiQ5�V���i?�9d� q�1-�
�glz�c@��3���4� �M�a�"	^Yi
�1�8[�2�}��ve:s����V����)�dʄ�b�L�{�",k��,�M���<�3o�ԋMY� �6�P��=����A���^{�xi�H)<K����ؤ��8�ڥ�_ �ASU���w��k���G��ͣ�S�	B���A̭�W�L�?��J��N|�]��yD�;�\u�����>���G���v�7;;��*��
33.��R�z��#����[�r����a���83ޯ;��U&�:6��*�H�(Z�v�t�ouT3(������bh� �ؔ˭��2�,)ao�0sA٤^��d��{�M
�+�������0��$����9b>�|*��g�� �S��!Zk�D؅����~�.��M.h)�h�NQ��+c�)⣄���:���v�p)ע�Lwb#5M�jQY�K`f�/���ܓ`�7�ݵH���ga�%3nA*l�TM��ð@m�*����nr�ьI�f�J���7��C�J�̢���
N���#�.U��^�U=�La�=g����w(�;�M%�ۇ2O��_��G�wC�ڸ𯻷䝟��n���2��,�l��r0T��H���Y�:�@p;�`t�j�S�i������X7�1�k�ȧx侢6�4��TcG���e��r4��n���<jXl��h �d�ꨤ�M��b����)r�:�y`��ԛ�E��>=Q��F�l`�����&��������
䀠����M��u�MOu�?LB>������)a�L��|<]�Y����]
an�a��;�>�dI�@��c��	3Ҿ�G��e�4�[u��� ������nǮV��@������2AV�K��-�x�/o���pd\ �����m�i�L����8��E��{�����V-" M�k_��0�;��hO�
n��v$�&����}. +Z}~�"�:��hc�ùj�?+?��?�o�S�����a|�+[��x��i���z��Wś��q�]L�z��j���3.i��S��֊x�7v1D�D�g���`�L������/`�_�QJ�.D�9Vt_n���\2�SӦ&ǵ�su�T������]�6��� v*3\�(!���K�=�/���}-+jӈ�v	����?}�)s�L�C����&�/����/�U�^����%�<��8�;58�Xe(��$[S�_�1��F&�����n� Ŭۖ��!��=g'�*t^�ؗ��f�[�i�C�z�<���*�ְ�@g�šEH8�˲b� .oO�a&���[Y�,߼�G?�\��;�J2 %C<J��'֣Nq��r
O��� ��<�dZ�M�&i��1�g`�4��,D^WȔil,�I!| �$Ë�=���{�43�f>?�#�'�ՍSR��#���^�v%�%�5iX9���K�-��*��9f�2!���A��Eفdb�z��!���*�'N���Y_M�,7Kk�}�V��TH�%�.�b�E;�w<�ͫ0u.x���w>�r�y�~�������hl��l�(}�3��'O�P]w������P	8�F�9���<�|��-m#��]ަ�
�bߡ9���<�f��������ƶ����";������Af�	���ϥ����`�����>���e��%��0�C���c��M�@�7��������uS&P���g��o0�W�?��Y�	�1���:z�S�ϟ?x�MH7�b1��R������ɱ�,��>�!ǩGf���L�y�R,�,'Bu���^����LQ���M;��gp��#���a��`���g:C����4����h�Б2!XY#9\D���N*�A���I8dL��=H�)�윚��x9�h��/�v���r�s��d��~��/C�Ï0ڞ�2�� v�����DHб#��1;�b��O�c�ë����ܕ!L:r�IJ`^UC�E\�b�0�|<C��8�5@�dѶ�#��Fy������=��cg�  2����4����\���Хg���o�mĝ�G씟���1<	�����zݢqٹ9�����2*�ٛ�3���v7?`��|#G(�{�B[j����c}�eR�T�G�7@?J��)Q�����-����!�n�{�ی� `W�eΫ�f��`���˄�Hm4���-,t2j�"���c�x$Sξui%�/n_Ƃ^I�{av^�*��)������ڦ,��f+��c�W\>D�.`VgE�=�[FEX���p�a����;��q4u�\WWw�a�}�W9z�X!i���u��Z&{ù���b���'�t� 8U5���nC<��0�ׇ	���N�w�0�vF�`��l��.G�.�[�u[��XA����L�@�<L=�L]��h���W�㶾]/D���N��74�}~�_����]&x��D!୍�tny�1��,,b��%西��gs������T�v�T�Nw�8d��^����U��u��"I�X�E�E�q9��(����(r�$Z�jK)����96�����J7�Ho�����C���6yrw��K���6�3 k#\�j�m�.?|϶�H�9���|��y�j�q���f[�V��<�.D\�T�����F����ܵ�,��TwhC ���ֺ����=X�~2,�o��̔�|l``����WC�r�6��߿]�W@���s�#JuN�����1�G����p�%_��2!�//��پ��E+@g����(�fJ(Q<&��{�Q�
T>U���XF�T褅���\B��T��P��"a�o3��/A��2���ٛEڳ��A�R��c�9�1 �gl�BuY{�F=v�#r���m�x��z����{�$�=`i ����;�b��+�D�[��
5�z�����V&]��_���i� �#1���h��L�%V�����+��c�!X���J��[A�4Ga0�cgu�/{��z��LI�P���\�W��B���R�kwl]�k���|:�^�`�ut���_��/��KO�������?ՇZ��_(����󓷏P`��n�؊�/J�k��-��
�F����1vz��qO�nLk�fEdfX��avb=�|�F\��i�q�?u2V|5<�݀�fg�� ?���^�↔&��Ή������ܬT��R�~ƳUl��W7z0V�x��1z]:.�+Z��)�rw�?�[�#�m`��b���T0��@l��Y�F.��
�n�F����c�����`�N<59��(�_᭗N�:6�f!QC��A��ƥ:�Ro����-By�6c��������D�}9�\ar I�_Z�E�E)uR�E�����-@p�w-p
��=��<\���xK�?G;'Y�h����K�pD�Ъ�yٍM����b�nWf���#���~�����1�������Y	���+>�Q�}�H�[�>l�D���#x���O= ����	���,�(xLF���q7��q�pk9�~���&O� ����z�<S�:��]J�ۆ\w��Q3Z����O�.���@q�>�乱�dG_/��=ba���Ɠi�5]?"�9vՎl�`�X�	TT�1D~���_�GX	)��!�0��I�D�Uϗ�͆������C�/u���\����x4޵��y�2�۪�)�4x$ab�0hkOY�� ��J�2���/;�*N�J/�`abĉ4�`dx���} ��!�"��犁|u��;�0We��j~�T���sgb�7�������n4D ������j�5�W<<�G~!s�9��#��'m������m�ھ%v�&��U���j�1��������N��Z��g}[��o��l����Ϟ�����s��`g��8��-��4�P����ܬ[�*�@��|��\�A��=�(�����뺯!�>��z��
I�-���Iˣ�ʏN))�u�H')���r�aT��+;c+@^�4���<\�w/�8��_\�Z3���\��k�}��p܆)���~1;Y�#ɬ��^]�Pа�a錓zI1�"o���uNm?�'��ύ���[�U׿����rW�Vj�(B�1�h���A��C��a&FEO���0����oE����-�:���5/���5�5NWa��4NՏ5�mn/7��m d�O!_����4M(����бa�"����/�@!i���F�\��8��c���e����f��#0�` 8�hI�d��HP>RɻS�����&��gb֪S��Gy�s;)ʹ�
KAW��|�K�]8�[�sǋs�N^!�䞁n��� 1TB��_#�~�C���UF�󬀉��(����Q_-=f{��s�j�h���E��\կ�=Ks(�A�\Y�5�(�C� ��v���=�~AAp�d�!5�����8�<����rt�
/]��l9iI�6�
/�ͣ�;�6�{�*�a_��n��<�_�$q�����'�oO�2oW�1t�_)Cf��+s�rރW$����L������C���ٍTܟa9�|n3��Cq՚�Úz���Rt8��R����}�'��P �Y�Ks4�Tv�UX;߶t����aIvw/_m�?����o����"�~;٭�E�o��To��ē9Z��!AV�R���oY����3��;3.D��)M.\�)�>-ى�&Xse�"�B������� L��F��e:TK�sˏq���5�??���$����҆���5��,ك�W���=��w>�i�R������ha�(�AW�����<At�^�$�=����1Yzә���Y�.��}�/Ǽo��Qo�Ytl�o7���@rEWLNra�|;5cU�7 ,B�M3��]ĝ�޲=0��X��2ڒ*.��E;�4��/��yP�98fL`T�]�p��-�>�L��Q�8R�O?<<y��o�!w�"�f�X+?L: ��Y�%�ת�+�n�%�[�����h|P�`C�κU ^#�
Lf�=����$僕ʛs�U�n"�J�~�D�����ڇ!y?g}�s~#Q(~x�A�A���m�a <M6��nWb�Éqј�E2�W�_$����iX��ܓ�e�ٰ����rE�V�=�W�9��r*��N��f�GiYВniҵ��>V�󽁝6ӆ�
�bc�謱�r����;��6�w�٧�
j��d���������Vˮ���Fw�� 7R~��u�?v�]�r���ux;Sj�MUnk~j �v��3#Q��S�nza��V?���Y�V��-:�0��C*/r��Ea��J��z_�L~ٚ}N?�����ђǩN^~���w�Q�2���t�ˣ�v�*r�~�X�{��E(�~l+{�_���<BP�|y����f�jf�b��2��72NқD����<%� �Io`���h{��8�v]�w���%��0��A3֬D�;��~0����)�*���^���{8�ΡdRe���A��]�FTb�jWF��q�1,s���EQZ�>��μ��Ԛ���ֲQ+�"����9��f��L`u���
`�>ټ+(ɠ|z��*öN��K?�,x��(j@�67^7����v�� �lb3��@i����f}�O@�B�L�ϖv�6<�W@.��JlD������ʌ�19e�s��G�/(�c39�$�{��|�.��z&�II@(@��כ��D��&��PJ�?��-�&����&�y�7�-}��oϫě���H1����r$�]�D�i�W�^*�c���|�=�Oε��-�q��(�2����۰'��}3n��J_�x��;�F�!Å�cآ�W,��\(c�טYO��۴eI�����[��kζpe���X��9�|�
{0z�i�S|���O �-��z���:�-:�Ie�;���\A|� ��)ƕ1����ا����h|����ޯ;/2��ӵ����A�a�^N�19N���<��Xo�9]�"���h/pV�WCE�`߻7%���3U���/�;�������'K��͏�X`�I�g��C8o�d˔�.[��j���]s{j�A����U�B�vhjr�5k�՘ֵ���>є�5?�	�ă���b��?�ɺ���ꊟg�x-B�Č��ы�O��IYhA9#��ϑ��w�E�wg}<�o�9�-�s�SDפ=tEj�}A?2���>���g���8����| ˸S�K%�RΝz���Z�Q��P� ``����P^1�ȸ�
fZp����Aha�B��4o�ﺋ6]NOi����?(!P'T�5/ICN΍.��쀄(Q�h?q��(=��fte/�*8�Z��o{�Ix�*�C�;�yz8�n��?(S�G��S���^BSpʏQ�׎�/�~,*vqr%�'�J��~[����RH�\��{ړ������EQ��L�UL	���/VO���D�wL���=�̸"5�լ�i��)G1ƈe2C��2˻EL*�z5�h ؟���%Hl鼝pL�!*7>6v��:�W�ݫr���s>�Y��1,�b�h�@ji��'����9�:���������y�.ᵫh�	�K��W����젵�w�!�y-V҅�}3(����? S�a<�q_p�-Q㜠�WKS���?�S\�	�����j�6؝CX�R�R͉�ʖ��nn�,_���M�����P��%a�iy��]>�:H�1��:��3j"�� ��3�>�y��P�ѧ�~��'�f�miL���7BS��������$���Ȝ��`���u���a'@����a�y%�q1�E;S��G6q2���pg�{��ԕ�}��p=����L۪ſh��S�27�@ʊ�E�r���״l�$K�`5�"��O��`B��� �E��?�ڞ�Y�<x��?�Bf�N�U6))��3����p6�(�t�i�@�� ��d�	;V�����N�AT���禕��ȲW5�[�OQLX��T "$)�E|�V,���&ah�eC���<�>Ea?�'h ����s��nwX���e�@đGN�xTǔK.�;M�CU�Ԃ$v���xӾmh�r~j e��,x�]m�"����l�DL����O�Z��y3�]�-�|�O!_�C�� ;�_��l���>��U��m&˜�q*3z�R�]�qA�/�k�L�r~�2'$S`���X���v��?!�C2�}��c:�EZ)מ����SS�d� �T�Ù����|oTz!_�{@��I��`�u�����������&�O��'���S��.xuO=h��r��ϡd���?��"`�:���� ׺���q}����.i#���V%�o��Ӗ:rŃ�Vل����_]1��v΍xA��<���=
E1a��;����7�[�8�~�W�J�A���l[��zd��u\	p,�!�E!7>Tn��ک��@_�.#w�w������V����I��MWn� =�46���m64��E��K�8=��!~�|�O4�<�L9%)���p ��*�(�u4&�o����E��_e�Evj�I�c﫷�L��	 P#o;:?�^�/*���4s/�u߉�~�g%O��¸���#��]�mhGd�tb�l��R�l37͑�N�5�	���½l��6���(�����wRp�H�ꌊ�̺a���s�a��Z;�� f\_iF���ˌ�R�!�7hW��QB�-+h,cr�u�j���w`��H�Z��i'B�O��~�I�1��?��1:=�K[s��q�ؤ]�Y�]g�JCV�f�h��Q�#_�c��i:�@���x��:��H��n�P܍�Eg4b'Z\R�1���x�e�u!���\��2������o�%{�����$c�B�:���pR�#��d���a�Єe��fTH>T({�	p�zc��%�v Mϸj�!� ~�(n��0n�"��KI5�E�i?����Pe-G�z.��mO��䊞��O�P�v�6������f��0���Ӧk��YF+d��	�J��
�ʚOO�M(�S�쬂h҄�T��>.�YZdx%��q�p�T�px6�-۸x-4��׬%�����g�>J
·�J'����d���p�a�$�@ ���{->Zo@�|G��V���2�u�~�����Ss�vp6/0��~�<~�6��E�N� ��Ik���^f5�Y<���$������w�?[n��z��+�w��I�Ƕ 1����7@�,`k$zw4=���4C���E�G�]���;  ��+>l���:z�b>�������x�i��}�}��*���*M��w�x�"��%ۅ�>���P`cs�b6���rm���Q|8�gK@p���2WV��k��5'���T�A��ݺ����DX�Q��y�����U��r�D{H�~�f��[}9�_e�ki�=��X�
X+��T�|��I�'�������H�q�G	R]g�s��!�]�Ơ-
��.	u�/ჼ����I�ٶ�:����r%R��P�#6����IS=�´���F����f��(V�i[�Li���25���^���ry+b�X��H����2��{���B(>��$�t���N��}�R�<\!�:~1J���s�U�5:?>� ���<Wԉd����`��&��!���Ϻ܂�b�V�j4�,�_o3�|��˱�;�(ߤ�W"��#�*�!�������jFY������E,j��o�����,X>I����R�s����pKY�]�ء�Eޭ�,��u��	�&��Ԉ�/�)���y
z;P/#'� _0���7���wS�i��3���\$��$D���{B� ��ڞp�CɇG��sv�p�g����?�Td�"��,~M�,����zq���{�a��������R.�p��nSy����tv������4�Yh�G��YJYPd/�a�ړ*g�5�(�s�Ĺ��/##�C�����
M�b��Hv�d���m�|>�!�M���X\�<U�C��l{J�W����2_��:�lQBk�!p�p3��A��m����c�>;�J���|_��:_�����6p�˖�R����;��D��n������a2�L�)ǰv�����g�����{���M[;בI��fRL�碑�Đ��Y�n�h3���L�d�I��U,g(dW��N��m�1FQ�&&��L�h�y7|����Mm�@ae�y� ��ׇ �T��=�/�)�ǻ�%7�����ߚd�ET�Е�f�f�Tߚ�&!G�Re4��ɶ,Vc��T����tV�|������J�]�=��"��^N�e���@Xþ���[y�9D��-�����טA�@`jm}ٵ˝��q�t�-��:<��z���ӅRђ=��\����o���%��9e_ڤeXt?��B�d�ت��g���HO�DZżʩ����qc�����WNd7oo}L}OCw�"S${��B�{3�5?"���ȩ� O��Kݽ|.8�P�1�*kڸ�i���-�j慘^�1)���OJ��o��S�T��0@]��f)�)N��Umi�����!fV����R<�hr\ú�+��+��g{^�)U�M�ƨ��*vJ�
�L��S�5 �)z4�ĩ�����O�u��ɧ�;A'<PU�Qߟ0��+�;�W�-��}���^�w�������@��Ơdn�Q�S��%ۨ+SKW32˖�ꑚ̹ ��4��Tk�b����L��6��I�^WD�KU�c�27�Mf<���=��v�H�>�1�;�>~XD�!����-�&V��$���:��kb����4^���Ea�Ƙr���JE�W:��ii�fd��$,
�iVis?Df�=��B��{�*(�v��J�4���__,�%�/;��T�,u��-�������mu8eIM�i�s�#t��o���U8��'W����[O_��"z|��g�,'�D��o�9��H�W��C��&"in?�m�i����Z�sIQ�K5Q:4��,�DE6��K�x�(���*})ρp�'my�Bm�D�ޤo�nϞ}4�u�<���̳�#Z����� r7�]꣼�x1���%}o�O�]���/�2�^��6I?�{��c�l�S�;wZ��v)��pO���<�tT��l�$�4پɆ�%�T���{i�;�M:�8�a��q��ߤpW�ԉ��P�xSȩ�|����"���d�@���R����?Z����y�"3��ᜧ���]��<�㲎��b��*~MR �b�E�EL�����Et�-�vq�w�����]��[N�R4Y�<Å��f��ݺ����K�J[��t����)S8�Ls1r�e��.M�啷�n�,�q����U}.�0�d���e���ID2TR>�-.�VC�1����3�����l��`J8~ĨF����*ILz��a�D�rSx�Yq7����c�����r<ӺT��)�dNC�����<�_����sTXb`#�M�g(}H���婫h�qFY=���ԄP�����`Cm�q{��2��` �Q��r��&���ے�[$v�����l���4���v�nj�yt��e~��S�2qVI�7`E�_&Rkv3��!B+��U*���� �-���|>�'�����Z�5z�Q�Ҧ��w��]�̏��b�@�@����5�Uq�ھ�ҡzX�j��W�к�"��(��G�{[[��!�����k.P6\hs�Ҧ؀1`�p�bzn>�� Ǯ�1�Ɛe�h�f�ڏ���C�~y�L��_�V�`�b��?|��-~v�]="��GnL�Z��'K��.�B2� �@6��[�L�&�x������<�iq�ʅ�/��C�LU�����;���0F>y��e䲑	���"cq��jf�����-�FaF�%��9��,ٮ��`-�p����f����Z��i�̉�{��!�[䖄�����	F��N:�6�Z�P?6�1���~1Y��9�̬�g���5�{)�me�m'�8Qi���
�ň��Da9�E�x�R鐣T}Ef�/�m�/[͊ߓ�����
�Q�M�� �o=�:�Z�v�g/�I�y��d5LXi����2�2=ZOz�J��x��
D4ա�p�s�h�����H��K�"-K�������^Р�Wo�! 6M*Uɟ�b��z�ɗP4��Ȱ����!w3����P���=إ�!�ɏТ�/�Ů|�j1�:Br%����S�z�k
דZ����gDR��"R��*�4�q��8�7��^KB6+��G�}�VC�ؒR��
�03�]�n���ᮋ���ԙ�L׮Ύia0�����;)R�z���õ�6z�rp�u��u��5.�-�O�n�w[������Í�2������s0��q�BR�;���7K��?M��+��F|u-ꖵ�h�%w�	��:?T����?O��>���_�1(��S����0z<Y]��@1o����+�Ԓ�ƫNm
�����e?�n68a���������V�t '�\��H��4�'	m~���)$D&��˙���<�'=���iΡ;��\�d��)��V���;��&��2EA���z�����K���uМ*�`%=��S֝�OQ?;M/�>]<X�g'b'����Q�U�[v�V��]$���zB$-b�:4�(���=�Q����-%p�(7E�1��Q����n��(��j1�B�CA��b���1�z�KvK#��r��݊HAIDxqś���A\N����	��3��_z��n]����� ��dYUh�����>��nA��imq�}� �/T���W�)E��WC~��$��K(�U�>��Wؽ��\c�9ˊ@�p�f�PmM�s�"E���1�҇$�i��.�q�.T9f�� ����a1��|AM,4�T 3\����c��k���2
��5Bp`O�hFD�^YD�T�j�	�A!������L$qFA���#��
�	U�����r�\��`�՚��7����UK��3=נ��ohVyH2N#l~G�D�>!6gdz�`��(�)I�,T}��ےb�K�:y�s��D;�z���W%��=�<�6���7�H����J�P����ة�dk���#�&�>O�\������0�!�|���:�>�o���I9��m��qj7Y[1��E��4%T�c�_ݠ�����\ۙ��5�D��N�����<j0����|�u���F������a;v��;����Y�xPX�%��޽`w�Ì�+̂w��U;m�>�� ș��5X� D4u���p�8F������^��>6���a���U��wW�GC��0����{6���"z����Г��喒��+�M�X���爝�xJᝪ���q��V��8h%�BZ�X�~z�J�ڻ
�D�ؙq較�|6���uw�oC�g���b�"���js_��[d��n�$XOۏ�w����<����Hœ��� ��M�^�<:]c�Ĥ���PB����h����,�S��"UE���0��oE-��B#D���n��^�m�r,�QON�jL>v���P��R9�kO&O۝ݏ]ܦ�bV4����K�7��qz��o�����D=ɠ�����f8qK���Z$��WfO�Uq���ɝ�i+�WvTel`�����5w��{�4[U��������+��&.�˔x�S�g��Y,��;�D�g��=����l���V��W-��I�i����K4ڄ�d�u�n���-��i�]�~`%'�� m�e<	@���鍟_;Jg�i2���b���b;�wTI��$�T�[R��Q�hgg
��p������?�U��Z`��\�@*��s�1m!i!xӟ?Hv�#�J�A<<oM������+r
�݅��73�V;?v�3nKQ�nI&�k(��s��p{ĕ�i���~o�����2�7Cʚ�"ʩ+�A#����%�Y�N�A��٪��0<��(�_�=�IX�^)p�+��X��Սۘe0aѰ�Ēٖ�i�΁9T럄�<	�Z)P�;�)Ȥ�ly�@��iB�F����;Q�����B5�޵�=�T���!]�z	�N�3lD���&*|�KY�\�����S�`��ϰ��e*n�F<lfk�����w��^A�O;c� ��(.��g�?�KH�jW�6/��%�I����Z� w���[Q4�@�@ݓ'P�~�y�#ߴ���U ���_�HlB*�)S�M�z�g���M���ʛ#ui��H�:a��((t n�?Gp.�<�η H�H&ß�N�b�G�c�vW	��Q�B���+�p���+��C��Ը2���b���G�ƚ�H<�i�7�9$��bK��]�<m�V�#�/V0o�s�3����������Z���%��(+֪���R�U����8o[xoV��?�0}ꅀ�	��݄�t�������X鈤A�k;�� �cA)
����͔9ա:u���f�{ϕ�S��m�#�
_��U�@!�.�1^J�J���z�q�V�*���b�X{��w⨸r�-�<@P7�S�\�H>Z;�7�1�:�^%޴�/W�@P �q�;��&��̔>~�dC#�ǦPݠ�bPSٞ�K�i��s~ ��k!���\�|��%r$�;ԇݑ�r}.�� ���(�OEUytXڨ��\/�f1V�V ��k����S���!�Τ��Ȝ����H��$/�7�-��e�I�=B��#K�z����iXVw.�(��ǼS�r)$��g4��	q��5�C����*D����/@S�ք��M`�g�0H�ձ6��6'�i�0�X��v-�����H�h���9�<gW��T����z�'�AƆ��˯pP&���o�7+���$��38�rS�YgS�\�ܸ�$x֋���~�T�@Y�Ŷ�����R�]����?}�04�!-g�{�p���s!�eI)i
�sn��� x�x�w>|ۼ�]=��ի�MW�Q�*L��,���Yf�=�໢dW˶)��O��ߌ~a=���@6S�5�V�{�~>@�S�>��zO�ȼ]	R�}�%:��G�����wn����/1�r#:Nz[�4{�M��k�H\�;��z����+I�
����/�n��̙�BV:��Y�M�iM>��c��:��or�`{�p��P I���W��%O�.ô���������~-�|E�l+=�3��U`x���tz*�P�`��^\���B�e#CX�ρ���$�����*˚fN���ho�����_S��]��ۆ�
�Ao	M��qvM�$*�*��0����hj�`A<�a�%��ë,����XV�q��o�,=�/Q�8	��k_�ʑy/�׹e��[Nv���m�0f%(�Yi�Y�(	銱�T	._�G���Ym�
�p-�[uI��&)ز֑��p�Ύ5o;�Ig����E���դӹ�Tڀ$j\�,#���@z���kx�K��'=�F�M� �<��Q��o;���ř6�GHh���u(X� ^L=�D���68|�����O�vRoo~
~>1��}*\�\�hO�C�t"�:�M�wx5��Za;er�y��Wad�Gb�����<��) �=ڷ*#駸��u�&{L��Bu��6�]7��VB4�/<�6Qm0�	K��RQ���w\#�&�N�9d�^�U�'�����{n��U�4N�D*0�P���P�z5�Z<�YI�A�f��U+`<^��8}j�Tl�GTtj�)���-=]a8	$-��.�$�/�1��߄A�)�R4�@����f�UQO�rԹ�����}�i
��JÁHq���r%̕��!��.F�O��#�u�=E!$���u����3B�VgZ�
v2�ߐ��S ��l�PX�R_J��e�̇��녺��N	�k���ގ��lj����7���FȆ�����폏	N�e��5~������>�����ȟdѰX�"��{GA	x�UУ>��V���R��y��縉�)�� e�8�,{yNG^v��� �b4I���1�c��ٍ[u�+_�>@����7?^�����TOi?���T����흿c&"ʒ^4��7��%�n�8n�k A��&�p2k,O�{�;�kݼ�3m_�j!��"�GZ���k苂�k��k G�'L"�4��$�j9o���)�c�Cp� H�����~`rf��t��yr����ם�p_-Z�]�ڰ�:����|��P|�A&��27��P���B˻}��:��� �����������һ�I�W���M� -)i	�٢�\S���������XH���0�d�s-Wj�)���-/�̤�{��jZ7��z�*�� �����4������SS6X�r݌�cnޓ	y��5*=jS�Y��`M�B�	���@2�3�t�T[is�KUa���x-���'0f�Y�Cm���-�Td7�Y���A�ߣ��<�@���hjp���b�s�
��g���j���>�v��`.`E�H�4�kBd&XQ_D��8K��ʷh���*A�JM|��8=��!,k4J�{����S1j��' �ݳ	�Aԇd�*諏�����	
8������u4����#��`�#�mI�T���4�9U�χ�M�'���/v�::cU�f�rG=�,o���B�\/���Z*����l��d3���yH�!��q��̊��)���h���+ck�����Gw~lc�J����䭈�T���x���%���#���U z��\V�6l���0�h���u�9�ט�xJ�<�h����
�tH����g ix͂��:�����I8�a�+�oB6D%��F��v�[爗^�e�@s�fY��`S��y��EX �ˣ�0��d�D�N(�?H��Xy��
v�]�(��4�J(�I`| ����M��nQ(ub��M!�8A�����z N���@�&k��X�'/�/E��T���%JK�9�:�0��	~�R�fI�#�z�p�_R0L�x�e4,�$�G��8�?t����|��'�&��j�g�z�uR���ޓ�=�P����@:��7%��P�͗)T\�v�2K�hN�y����DRsf�0f��H��K���3e/��Sp�H����,�[�|]h-X��-ހh"��c�N�;HN\�U��Ij��`C�_������_�}lW�B#'�]�����2�!�S@3]��"�����ё8�1�r��=�FX�<�������ۚ5.=��;&c�M�O�w�ɍ��V)'P�c�T�?��
gl@-8sV����������J-Yw�u�jn������=F��M�E�)GV��Ia�L|�G�]����i�Z���������?����(���%��X��+@�,�����H�ي>��`�qs�f��� �t���R�M��K�%p�6�M�$�����Tb�Gp��ˑi�I�yJ�zV?X�J�+����b��1Cs��YӰ�\%6��Y�<jt���[wB ����'	�e���Y�Ӂ�ʷ�#L]����W��␝V��[�x�Rn�#�}m�"Ez�%�.!W�����oP�t(
$_-����������V5�ؚF~\@1D�8�S�#+��þ<�틼2�~���{��g�S���u%�K�$Wӽ���q�R�'��s��a~'ڍ��)���d�{ᅸ�����Yn q��O�2&`��Os�MG��P
�}h]2~�z��7l�@���K~zc��"���sl̩��l��9��;�L���u-�:w��߰�q����a���=��������%'^�_�l�j��盧jz���g獦��ߨ/.�2wy��;�7��bC]�i�j��<8ġ����[qs$��)���ڿ>�SM��R#2��v(�������
y�ψӑL`�5���]�G3-�Ѽ@��ҧ~��!��:�� D#��Y��:{^0f�Z�
D;�e���/o�s��E�c���^�1��/�*-M<��%�V,���?,����*�*A�3ｺ�@{����J�|�Z @�F72v҈HuN��P��A�v�E��|�f������9��`�c�H��c�C��~S�U��P�ƸET`�[O%
a�DŊ ��s<5J7��r 	�S�E<q/jӥ�u�:����՗s���ζ�w�Ŵ#!��0.���1��ݳc���@P &o�h��:M̱3����e;��8�a-=�O��2N�Tp�k�>���y	 �����t!J��7∵G|����C� �6*\�� �,�P�2�>�8��>4�OUO}3�}� �O乳�I�
y�6�Q(8.wu�Y����v�����;yNM����茀C40�����[�n��M�^�����:������x@T���s�i��RN�㿈S;C��H��7j*nE�h��7S���P4C�e0Þ1�N�z�Zn}Z�}i�0S*�@��x뮶|"��b(�ЯX���6�ݪ�籍Gܺ쾵��W��8K
�u���Hc��Ꞹo���$���~pR��yĠ�� �����>��z=�]П	����?���|yhT������h6}�L�I�<<�� �����jv���������A���a��2K_/`�.�D�Cx�ь�/�K�h�eh�i����TJ�Gt���7�vr� �Y ~����"T�R�5��Q�Hg���\î=���V��hÇ���{�8:���L3p�S+�J��0��w,nւ���_���;Ƿ,6��r���MY���P$_ �^��'�~6��G�k���>l�Jƃ����>� `S�':� ��.�����w�oU�VtZ�PqC�&�:W|�I��W�eT)�fjX���آ�,5CE�0{G��|��Y�� ��8�H�(��p^�i����y��h�hj{�>�y2�}7`j+��;�i�W�[�y�4A��mq���sG��`ϵM�D!VJc�|�mƌ�݉rr�6�k�
�����jZ�o�{��I49N�C�7����-\9ջ���*#��u��m��!��p��W�M��1-��1�9��f1>������"��0�P2O�3�L}Q1>Ƿ�o�W +j�ʁ* 'x�4�k{2���y�:��_�=((�>��V��LSj�f������%�iH6�Cم�N9�_A9�W:�w�{G�=�0t 7�=}B@�� sF��El�ϐ6gɓbY��>h�)h�͒B�$4#"���b�pw��Ƽ������,�a������^l� ��f�捓��"�ob�J~Mfb�[���P/�(�7<0M�ܚ�C^�Q .7�[sbq:\Q0���+�A�i���f�4��Bz���o~CkB�(�l)h��"�g�Gxu�C5��Ρ�ju�]�`|��䑆l���S��;.͝:S'=���h��r�g:a��[L{K`T&,�JR`��j%^�7Dc�T�냿C��oH��[����8]�Z؛ʍi^³-'߁�z;�4����Сh=_��#��W�E9��īj9�E,`��k�kʲ�'c��-Ų5�F�}ʂUzr�6u����O��/�v ʖD�W�Mv�<�g�Q:��%	��g��a<�߆�F����n����+�Ń�e%����1E�X
h���L�k�+�̜ eG���< b��C�C$sz]�A��%B-�_�ً�9H/�]d?�q Gè}b�o�����A��؞��Q};.eP�4\��dnQԪ�e��>���룩�$��:J��D%a%�2�ꑋ�3�.�޽#>��.S��G�UX)��9��vy���^�t�z���FA��*t�5ߚV���n�lN�\|(K���(�|p��6��s��!�b���d�NR�t}k��U~�v�Z;++,'@���� �=`~�`����Kn��Ls�,��������]]P3���t�Es�������zA�w�yԼ��P�-f~vrE��H|�$�}�������_�)�"�Ѓ�q��)iʿ�8 ��"������/<�y���K�%aho�l�Y� 7iB��Nu�0WU�	g�'ܓ��d{�g��QO�Ņ.up���zEl��A%�ެ��%�ξ����ޟ.���y��=�è�����Z�K�L2u��lAA;���Ա%ubo��]��T��r�"u�<�tH�X�]�ڍv?��J�L=X�3�-Tb�Գ��b",�Mt�2^��ۯ����&����b|꜃g}�|W��s~QA$;�W�*����Vm/���F�[*4���>E�n��d���)L��� ����Kx&� <R&p/��q%���13��ھ���BT��/�w{L�Q��	9s_�q��KTƨ-C#��cG:��áa�tZo
J��2mPRSmۙ��GV��U��?��MS�;Ժdk�?|��BF��K�Y����by���ި�sz$�#X�QnY��%��?�۫�E�~��A�u��3��!��� �U��&���%�;���pP�-8rnԕU���lČʺ툑��ڝUw���b�N���un~�R��v���`L�.ʠʺ�����У+<�pIP� �����xt?�
D-���B��z�ÐO��2�t>���ї�n׿R�@0�Ƈ��g�CE����ϫx =6M�j����)�φ`\��+�g:��B ��r�A��8�fm�|�Ƀ�
��r�E���;�U�r*�������&bS:�<�G�;�k��d��8�M���̡��֑5'�/ՈL�fb�N;��G����g�`�f5�.���-1���$��k�y%GB6�X�8UtVEp���Xv寻�%�y(��v��2�{�w̄*uSL��(U�ŷ� H���:�m�LdFk�m���W�.����1�*�YM|~<.�H;�����UP@�$:/��t�NNEm)3 ���A;S�7 ڣ��\�zu��0�w`�"7�0ؾ�U�El�U_=M9RE#�.��#F��gش_���o~����������5ʏU,�d� G�'�f�y����6���Ȝ#vHC"��~��I#�_ZN�S������m��W�\X��MrR4
���eҪZ &�
�.a�~���W�3z��ĩ�1�$Tz6��P)�K;��31L�$���fZl5���=�X�eDvb���o�_s}{혻n�K�:<F�Ǝ��/ԢpQ���e�o�]9#��*vs�pR8ةgf��t�qa<���M_��^+6�*oѼ��.ݓWպ�g��y���2ѺJ�xs�D�,QA�(8w��s�=�iI��#���6�9� �NU�ls:�>�Pp�����N���b3�*�-1p�HA.�d:/k�$�D������J��!Ϟ('X�2 /�w�����ώ5����R�����jd]|�޳� ����8�&ɵ]��pU�����$��%�@"3�׀�36���ʶ>E,�BO	��W��yKi�˹���*�gV�9�`^��fBw�6������hl��ik˩�`�4���� W�_vN�w��q
(\7��qc�q`눷�N+��F���*�����KH�3�ۻB����|���{V�KyQ����eޫ	�y�~�K���W톳v���Tj��ʩv�,���s����n����W(_ 
�,������O���&��V�Y��O�J��p�?yo�E�琅�Kf]�~U-p~ :���"��}z��~l��q}�ȥ<g(4zإ̦Y1���u�y��Z�zyW�#����c��b,��݅���N��XN�6���Pg��X,�#P�c��K�KN)�[B�λ�g���ؑ��n�?��&�`4�&��-s�/Ƀ7�H��0�`П����[�A#��=h9�Y1.ۦ�\�oy��YN���ڳz�._�_Bw�Cց~h�M�ݪY�G� 淠t�����i��^5X��i���rrSTzoÆ����Û<��i1����tdWFn����R�P�i%�u�^���t��ǿ��ecI|.��"6�W�9"�mӠ�h���Κ�SǶW��qJ���OV!�☂�e�G<Q�j$,�:P����X}b�Y\����bT�݈��M��/�8<�$,�/��ʎ\�7���؅��gF����nnA����]���l9m��c�-p�<=�Eթ�$���ʲΘ�1ytWIh��ȃ��_U�S�H|�)�UW*���[�`�ޞŖ�˖w���~��*,Ե1�1��z������ˣ�S�;�Rm��z?���Z����0�y(��GZ'*�;�w�h�SO�����8�i�\�3vl0B�&��J� ���}%�:+bO81YU�������) X��uku��"����癢��Q$�%pZ4�xk�M'|��~��xu� �c�/TCm�t��;&�!�0�r��t�O�l*�L8�e9��^nvݽ�IP�Bmo^YN-A:�S]<���<k?���"�%a��7�U��y�b�ȸ*YY/������YSd�Y��W�'E�����Z�	C����Qb?�NcL��R��)�W�W��YT�n�a�ᇆ�.W���"X�*�u'�~gi;f�8i4Hn��W	�s����K�\��p(�t��׬�����!u�W�|�YnPf��^��� �fn-D��W�<�QO�>�m{5C��:������ܤ�3
2z�y��Ò�����L�le�P���fV�r�� �:����nvޫ��e�ᚶˬ��V���]g��������,��N�m?J�t�t�����1��@"����"�1x��q��V��gL��xl�Pt��3,g���ͼ���R�=6���&�G(�P,�NwH���������_[�yI>L��>Q���Iߗ�CxF^
+�0���mu��t)�Ed3�H�����DZ��l�n/����_�us&�]�f��)�	',�Oncwl�{�u\Ե?d��Y-dY����Sz���"w�"��8D�[7k�p2^*��$yƁ��S�������
�P/��2Ű'"�*#j��"�p�,pN�^�RՅ�^�"#�?/|�|��:֊e_TR��)�9����^�1�`�[QϮ����tq�M����&h����yWaYiE�v��B��_*�#KA�4�4��:�a��~�'�	|i0��}��w��P�ں��p_�\������>i]�rI�E1��}A�a�bL�5�|q��':6�w�=��&�"��L�C���ֆ�؜�\�y�a�D\�5�7�EQ5� ���&|��B���,�v���>���bV����E��M5�,�I�ŋI�.�/�Ю�82��G ��$��\nR�L<w���
c�z�*QI�O�n&�|�-%��#i������Ul�2��Pn��s�k��=�Js�,%`��*Qm~�����73�Fɑ�~�.0#��G���K�Yw����5kH�,j�w�Gzo�� "����q����j,$����~�����?��y�b$�}a�u�|�-��i��e��Ք�^`�MY*=�q.��-q	7O�{��	���BI�y����Fx�q|�>���U�	泔���S�RCy���,B���Q���^N|ӝ��l�u{�v�`�.�����B
�1�NN	t��,�R�8�1�+�W���C�b���}6��_U{q���#5\n�6�HW���~��E.����!�U��$by�RgQ�U�+��" (�F/�y��a�=�h��su���T�joJM�_�1,#��Km�`!#l��8&��3�H Ud��h�º��ɑ�ݟ2��9���(�zbWu��!��c���6�Z�����J(���=@�}6\��X�H
�Σy7R"��-��x�ҷR�A��CB�Gk<H4~E����+xBZ�400;��R�ulc�3`�ӡO;�ti��^ؘ������*c�e=��Μ\�����Y�u�G�ܲu�F��Va�"�xN{)��s�|N�鲉� d�rlׂ���..8A�k�ƛ;	�$��������>�QhL��	�~�g�)k��=�����uj��CJ$99r�3m�1���0*�o�ڟ�r((��˴�5�C���C_�aU�v(lrP*��ߓ�e��V���B/������sp��Uү`s���H]+Ze�"�J���h{rܥ��5�!��E���[#�h����eB��bڕD@�SoR��7�ݰ\�:{CPj9<���Z4�2wd�i����{@�V}&��m��IF�Q%�.m�9��ST�ay%��>Ә�ץ��tm�v�k7}�B���^T$��QՖ\�ˠ���snq7ߦy�ɁKF}�g�Qb�ȑ���/���`%v��gB�8#�^GN��2^���w�a�F�o7TH�Q���,F5Q���E�9�^(�ϧ�����7��
Ɩ˷��e�1��1�#S�;�=�2��h�����E�^�(xuА����m C˕W��&��=�7xs���}����W�o��"�>�=l��;̞����i0��~���r�sߛ�,0�\�(�Е��-8oM�fN���1t���l�+����|-�~��A~����rո$<�w����#��8�im���R9�)���:���V�C&���'"v����M��u�@Y|RN=�l��%ƺa��e�0)�H�W�e���r�hry�1��ɉ��:�8��<e��6t!�Q�C�,�2R��3Ҝ�[��ȽpK�n����5���k�7Ĉ�^	�5�s�Ђ"��#Y�[�`Qxvv�y#�m��O��bŔt@�t�Pq�ڀn��͞�y2p�G���uW�U-��5��� tLv�$�Y�=���k�	�]��eT��TW�yOy�=�dR�/�g�;�
�3 Z�]��R��VI�B�=�2��c))�NSP擖�y"O�������YC���I�Q��z���:�Ɛ���m���b��Y �%C�В���s���E�Oi��ȯG����d�d�t�L�����m1]V��h���I�z&JD�^ �Ɗ6���F.��DX���1�bS�=�S����[;B�@�xZd��=�	GR��0�����T�BB��+�
�uJm��}��L�� k�x���ܰH~ǹ3P��4�5�������7��ۆ���^��R�7�^���� ;��nf���=P�=#��qӢ|�_ԀeS����T`��0�~����=�����+�*}�LJ�x�!j���vf�Oe$��''=�3"��i�*	�P�+7^���`�4�<���{�$X\?(%s��ي��T̊\93螂H��C�#u�yv�ﱪkJ��	;Iφ��d�g��2ƃB2����d�x����3:��7R��#��D.)��f��`*���b$�g}*���a�}�hk�����'%�5+����[��%]�_VG����GlR�_�3l�1���8�0y"]O�U�1HOnT��Խ
+g�T��da�v�n^�/�Z�h.�N�6���X
[!m�V��`�9��X9���q�T����`�b0�x4�'�y���!�T���g���㽘h��uLMt�|��p��:����P>nF��a��E���-���;_p�-ʜR�z� rk���=݅"]�	�) ��j�\LS�xzv���4B5�����w�� J��㘎�DOA2�'��id�6b��h������,�gj򜨃\�[ܲ1�2�*f�E�=��C}�B �C�|d��/L�(��x!w5�����c���b֠��V6��"�-:i�rK ���p�/B`!4���V�m��&��HLA �?x���O��)`0�31� �V�7.k��&Y��\��*�Y�*�Ej*X�Jk�3d����|�o_�n@,?H��b�P=N�P0� ��N�_���d>��Ķ�������im	;K�[.BȚJkC� !_�	qMpF�@p H5�c��\�I<��*����L��F�.RS2����p ��{"�]�-���	y<&�55��D���1"r���9UY0�Jg�k�.7٧�=�ځ�ٍN�`���d2M�M�L\u-���/�0�tg�LT+���E2�xRӯ�Z�
�$�o�I�� 3̑48�w���r>Z�V �Fw@3��R_��&u|8�����&����Q��aSJ��{{�n	�l#��9S�dq1���^�lDg6%�;��h��J9��x���&0$h)�|������D�sl����U���̺���g>t�no��iB��6�ci
�)͹�f�a��e7���z���� A��5X�d%���������S�p���ù�Ʃ�vR����dD��C����ru���
'XMy�������W������)��1QfIj)�K��n�	�K�9�Y�d
@E��M��C���2�b�e�����ֵYy�M0��]=�In	��-4�����/r��r�Z�@1ק��7cv�Vn�x�ɬ|8��H>�ޝJT!ܱ̺���O����{'�Gw��)O �Q'M�O���?�9)�?P,3��t��0n�s����*��{�6�K��u ��%!�Y)�ua0Ԝ�۩����S'��I�}����"����ѳ�_��1ڽR��z��,T�w_Ƒ�'��/S�ߒ���)�M�]��<��.���$���F�Oi�|fH��vD��-�Ԯꖗ���ۺW�*���?�b���v�з��"*�tB�<�_2��4M�`�Ye��<U���w#t��������l�3j���nC����BT����� �7�#�,d�UDC���
�]��7s���)�$��\�����E0d��&����D�2[�q��Pʶ��4��!���8���L�Mm4�؇{�ǜ���	�x��5 �X���5�_����+scsj�3�6bD}��D.z�n��U��A����BB��3ܓ͠VhRc�@bk|�Q̟�W�`F8+�j	dR*^�X�[Q��M@\��M7iBӺ ��"tڜZ��p)��a=g�h�^���A��_2T�,&�L��wЫ_/�|�w"҉P���