��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P��4(��-���W�J��3�R$M�����	��0����;n�>�Ҡ�X����r<^�+��l��㚼Z�\$g��@Ȱxi�c��U@����Z���Ȏ��+�����V�f��\�.�^Q��5Z	�\s���^<�]��4YP�>h������j�p��,"".Pܬ-Ja���m��q��{O.Nx*�����)��x1�|�Y�+%��q�PG߿DU�c]�6 ��Vw��f54&F��Z��߿���_W�'�y�[�<4�̠WL��!�}N;��[آ�<��T�d��
�ߡ0i�\~��Tf��4pk��Դ��`��y�[7�N�!�7S�rEz\���˕p@l[�",�9j"��#�0%�)'bI=� �]�9z�x~���X2�dž4v��+[F�3/�<�3��v)�L� ���c/�Pܦ��.����<�}��L�;{�a�'������ ^�$��l�m����RqQ����4���ܚ?i��~aj����T�|qWc�Y�E�
���Z%zb��Z�lgw�X����H9�m�<�G��u�Tt8,�Rr�\������$�3��I ��ԃr)�,B{
1u�orr��:]��"R����p˝hޖ/���U�@ʺo�(a��� ���[�]9s�95nϮ�&'��iN/�#�r�Y���g�?��I]��aG��:Q�}u(T����%���oU��2�`��\@���!�Ά��|�E.0�Gē�,��h�m��b��R�M�K!�N3f���s�Y��"�28�*%�5=[�og�.�~��0{�AQ;�M?��qg�ѽ��F��}�&ĝ7��!a��\�]�#"�e@1G����]<��T�썫i������>��'��z(��;��S0O���U�4��η�A�WF���;}�G�O!^n�V"�2�<X>7�ꓐ"��Z�Q"��sV#i�5 �t+i���f ��Q����+��
G��"�!;��2b;`��	�Vd~8����OѶqdУe�D�O���b���q��V��y�c�.���9>I���oD���]�M����[����j��s�_��ű,�)�}~�1�=1N=�)@��]3޼���ӑl�	/��*�\�y%+��$	��?`�)����a��g��8����VD���n3�#|m�]�Ӹl�~�(������r��������ד�I�����~q<cH'`�Am�j����D����Бω�u�n��Ƴ���f&�ĺ�����w�_���C��I�U�0����!��|��9�̓]�b֘L�g?`ޒ�q3h?�r�7���i�<���G�se�}�����}��͸v�>G����HR���h�����/�eFB�Ǽ��Ʌ�q�q�D�����S�1'j �2�ט	>hٚ�2p�ꫨ��k]c���>���f�3��9�Ȗl����vl@�9��K�.=6ĸ蕛8rJ@ͷ�/�B����c�w��[�[WĴ��8ޭ�H�э?�ޕ+��j�?FZ�V����_W֮e���0Q���}�,CC��4̹87�۲�����8>9�I��_�l-̞i����L�1G�f���?w�2o�Ҡ��LL�#��S~���?t��|��R�R����L��i���fN�!,�RP�Hso��}"���'�}ژo���-c�2�+{��`��]i E(J�.�zT��}��<�=j�c'�c=v}������q �$!��ˁ�����5ˈw�Te�HG��`��}1x&몳��Fk��2��yx���n���*o`��ikH�K�܀$ma $�B����`�k�;@:����,?�J�r�\C�-�&>(G��q�ҭ�����+�DUr{����^��oP�}���BE3�P+ٴ�y&��ý�+!�K���(���Gڮ4Ϟ[vc��J��KN��G��u%K
8���$Y�|�R5_*�JG�Y��p�m�#w��d� a���֤���m.Rj��.3i�+D�V"'�Q�f���U�ą?'3jM��mX��R��e�5{;� �!�	����@I�$kʞڝY7q�jg�D�"�|⥋b^I��_�����8�\9Y_�����M���?2~eń�@��n�Y8��kO=��|,]B$e�|8	���b�H��R�p��Zoɩ�$���^>�S������ ��MBiع�G%h�=J��9�F`vhj�D�^/��*r�	�U�!�G�L�`;��K�������:'��l�����A"9�'��`7�+���ٟ����/����T���~�\�%@o)l�b �p���(��B��aq#�H �^NU)�uvӣ�@U��eh�oƠy�|�(��@#�`+\r�V]��Vf|�z�D��-���)ƈd��Q.;q`��H�؂+�L�%p�����Wk��M�
ւOuD O)V��9����L�������>�H�'��1��6�����,	�ܰ`��0�$l�N�o���F�C�o��ew�Q��Ii�$Upf���w�R�?�FR��2�s���iJ%��*'�I�/S ���2)ʰҟA�v%�!�ys�EO�U��"ɡ�az7$�qv�LV���j?4Z�����>�F��=(T��d�]��s/�u��tQ�+�3Fb�����b���m!@�c&+�:1��y�5ѳ�Ðm��ƻ�B�O��(����r�0�� ���fS�:v��y�L%%��7�gޖ�WD7T��f"p-�d�uV�RH�����Sy �=��#�����y�>!޽3�����8n��� #U_7�����oER\S~�$l$T�)��ݐ��(a�uv��ˌ�îa��n��}��P��w�����U���������/� ��4�b��:��S�y�͜���>�� ���R�8�ׄl�a�՜�r�P���I�	��*_��%��?�N��V��v��i8_wu�˫�1Fm�(1�AS$�}��v_c6%�S|f���,|%64�QH�V?�O/_���t���e�HV�Ī@�5����&β�?aH�w�p�?��<�w�Mv7�w��nZo��/K�at\+���{�ȫ��5�s_���`�aۋ�ǂ�)�O��n�ފN��m1��an�3zyjj����*�\!�]�6�I�<�t��=��8k׹�S-&�g�d����	���7"߀�QB����@���L�+ubr?j��gzn��uXFLM�H�~���:��Z�����y���a�,%NLPAʄs#��<F���r�,������MU�,s���d�h��hO��2�B�����eRBOb=�O~���Ä��Oa�W���tOumLz�p�h��"�����1?��媝�m�Q׈tP<V�5i%I������V)�d
Ns�`a��9���x&�3)o\B��>&�� �6������ n�Y����h��KډJ����4���`���0h� ��6�	�C_�kf�1��uR����N��R"��q���-��/|��ʿ�,~]-׻eC�v_y�+��%\���6�ڡVA#����3�Q/�f�a�������k^���ʯ�TJ����jF�4~�Ү��t�+�<��9#�Jj0T��=Hd՚�	Y�8�Nzvso�Au������X�.ߏj����#*�E-���2[��*�3X~�*�������/���h:�jڱ!9�=;'�5:)�C So[���JZ�(E��h�~�
`�ՙ��,�������͒���7����E�p����[�s�t�l�z��9�=lF$.i���[81ؽ�wĐ�����=����a�$��$\��E�	��W珌���	%�&���|Ӝu�AE�7���,c��|I�H��қ�X�G�}�u�&0�Q%����C�S,���;�d=��.$�UF�;����f�cr������t]���#hAs���9��iּ�z�E�#���gpmd��`��Wg���ՙ�u0�s�����:�J�A�jp�Z[R�t�,8\'�^l6#�?�NV���}%3\���� �6U���Umk+�oR��4���u�����F�nt�-�R�S��vI��#���igB� ~݄`�۔A4��z���JGјNi�6���43��p[5�0����:sK�r%ts�&\d�go��ܗ��&C�/ʢMo�� pڼ�æ|!+���n���$��D̔���٨���a? ��c<��N���d��;�^�*���FK��/;�
�k\*�C2j�P'���9Q��۶�p���tƎ�q�^f���&.�S�u|���Ѻ�H?��<{%�)Bap��v�s&bȅ�Lq��|ı!x�c
|��g!Wj�I�S���s����V�6�N�MZ����ɓb� ��h�������YH����8�`�
V-����}\���4!�� [ ��yB�T�v��u�`��Aa��}��԰�vyvU��}�w�ߓ����1�ˢ0[���J��#��8I?i���U�	/���Ig�xS�z@�E=U'S�1����r^�Hm4Q� ���d�3m��T�l�0T�G�?7���~N��\���y��#�\�n�����tZ���ۗ�2�M��+���fӘ*'���!*��)���!ؘ��Z�o���ǅӌ(Ҽ��n�P�E@5q�=��JO���Ξ�Eo`
7'2�����ɂ߼�}���8��/�m�>N�ƈ�X�?E>/�w���4�{�ȼ<�}�"��xR�S�@�O�b���	���*���IFC���[DV�H�]����Q��Z8)[�v=d�!7"��4}s,7Z���E�T�oM���k�zvU"ڟ��������*�fT�[���z`9?�T*u���NN�7�ـ��p���T���U��s��m�&�6�?� �$����Wo�w�y��t�N�ؠ&���
�
�w���j�t�=���'�0�]d�dh�ov�@�y7z�O�"��mmcv󎩱IV������S�N��®av> pK���C�ȓ'J،�&[8�cSe�LFo�4�3�W�D`%)�W���|я����"�� /ԭ��&l�4��a#g�П��W���EA����߉���;q����\��[��L*9^�56��~=�yq�<ޥJ\s>C���F�D��u��I��H�/�/�Ӈ��&؊�ih�uw�
cE���+�����e-JJ}��څ �{U0&������/=�������U	}����(��}J*ZV�T'[�}a�K�����O���rf����	����>��u�W���D�!��P��0�Rw������.&��-m��P�k�h%Is�98*�Qlj1\k}\�۾�D�S��@���~9O���
�\s��dn�O��y]�`�k��S9�;E�P�2#�fM���O���V�17�ng�K�j��2����e�A�u�d��tE�V�O{�ʤO��D$� ��q��b8�[p�G��ز���9Iё"�˳%�2��Ȭ2.��1���d�-m����6�����T8Q#﯋���k���zt�R�[D6�A+@ci��}�x��CV`��k���PѢE �ָh_{��-��F�������5�����"Y��F��J���m��'K��
� գl���m؟	���C��*Fou���s���5�D������z�{l=��7hj�y��I���Џ������f}oD�A��I#&X)�6���dFy(�obf�н]�C��.K���;�+�����@�J�Y�_�\-u�8�\�����Qg�AG9�S���c�q�1���\�XO�0!�N���b��a>�L(hQ�Få�l��$i�H�3N��e熎�"@��.�p��=�?�c�g6~��o?�dǁ1�l��`o;��ՁS��<�r©qB%5�D6Z�s*2�?�?�3Ow�]�:={8(r��Ng/�e=�y�C���(B���l��W���<�K�q^�nrw���a�D	�3�Y�zs�jR�&U��6�w�a+�?�]��Ӊ�}hG�7&c芜�`��p��sr�CڠG/m8m�N�3߯Ƕ-��CJ��e�8�
d?�"�	&���Ͳ���7Oͫ��J�����&��Ţ|�Iۢ�hV�O7Y��i�V�E6���P������͠Rߋ��V���"3�4dxU���G�v�r`����>�(Ѿ���P�b{�����\b-��g��a��)��*ݫ�c-�I5��Sɧ�-%�]�M~�@%VDOa�fU������ ���#�
���.ԩ1({�k�/��h����r A?֌��g�R��C��Э�%|����~c�u��Q^����u������*nZ_��зA��b ���AE���j>���H�z�B�o�3}�L���m�̨'L�
A����V�j�i�o��~")���Yp}�h?�n�=$J2�H����%��r�J�j���X����2��7h�Y�>�XG�X�`aF�p]q����ȟ��U>r.8|�dzZ��&�i��a��`A�VL�����f��N��qM�0�� CB}"نm����0�eIq,�8&��Tʹ�A8_ͤ�م�_b���Y���(�}�=j00|��L�>�������R@��:y��S��r��C_�9Gp�Z1��C�A!|r�&%3ؿn���]Zu�������2��̞ˤTE�5�ĂB,�Z�D�8p��	c�9r�|���ǸO��~5���p����}�<��0)	�|&���MR
�J4�?%���=8�LAȻN�g@�}}�[-( ����F�3~*����GW�7��O��8vҽ�]�ő�[n�5c�v	N�m�&��d�9B.f2�$e�T�=C_����Y3��D�fSu!m!X�n���+��t;��E���GO�����j;�Dv(L6�����:�o����p�� ��a���nP�~�X�Q=	;d� �Ą^�2p��x�lD(�Du�������f�����d;�#Our7璵[!a١�D���K������=��qd&#���0�%V�:N"��7"BY�)aw�����5yJI�����6W�)"�թ"��
?��O��()�( �l�:J�T�S�?<kM���_�Al��Y�+���٘�g�L"M��5����H��L�Q8�qr��b;�)��&���|ҟ�[j�,��)�ӹ{�&��g��1^���ע�bi��*L*�0�X3�1�cP��2�����8il�.��[�U	Y��o���h˾�x]�m�2� ���!����M��*���K���^	�lI��=�V�F>� ��'#��������s^q����R��h�j�o������BE��'z=|�H����!�PI�fK2儽e04kg|�07Q�k6�o�]f�*�_o��e>�H���5Y4����--����k�Y�Ɩ�_Ն��:�ΖTJ�"�TU.��y�tq��B�ܰVR��2�jYQ���w@��6GC���=ς[��o���ІHz������ɻW��Q=V,��Xa����[g�R��Q�`tb��SP��!_��Di��MB�����D޳zB�$���~��g8�e|ϟ5I��g��#�^���w�-q�CG��B�QL���f}F��~�����٢��p���;�@}]V��[�GG ӕ�mA��I�W��H��|�^�;�����L-��|�ד���e��]N'�8�ͦ�����-��-z�*O������$cf�}�;���M��cn�������`�XXP�C�NخN9	��U{�*���3}VY��p�]Pp\���@k�	��l��#���C͌�!�Ba
����N�}�
�4o���x�	�X���GtW��@4��Ѕ^���k0�ޙ��D�<}��D�Rr�[�؅0;9�vJ�(#t�!��k�0fD�ٲnCUA2�Y*�}���tB�;�m������5�����I���yB��m,Ӵ������
��R�����/c)A~�|_w,�L��QN��	�ۑ��At�hS�Z�妖6n�)�mh�5Sj�t�-�>*V���YC�^�g���!Ȱ;`�}�~�G����w8������t_�;��5E���	�j��ЩP����|��.����^|��tʀi4ȉo2��
��3�)�-Rh7k�h5��O;BX�ֶ��}����I�ʤ��4 �{T�_����!ױO.���mV\i�h[�]$���w��V�����>s�IM����]�s���e�b|@2ߓ��W��G`��ä��������,L|��v}��&��Ss�0Z}���J�bƿ�\��8ZI� �eAB�szgT_9��aO'���Ltˏ�|�`O�b��T!M=?���b��XL�r0m�Ň*N��=�
f|� �a���S�ti��E�
X.� :��T���l�'�f�g�k�ɐ��M]���������/k�/����2~��4)+�OZcȵ��z���'�Z�+�v�׊��o
�� ������F򮗰#2[����+��F4 ��y�����K����h�<��1���~t|��l�b�z�}���ầ~�1o��r6�1�����&Ⱥ�\�zI\l��Ѳf��$[�U��Ӭ<>�Ƒ�Z��6���)��h�4��i3<��PA�J��q���V��_���ţ�آ5
-bmѺ��z4��~g�Q��\�aZh� ��AƢ�>����̏p������z�C���[v���v�K�=�o�H��m�+ۄha��P3�N�k�%,��_O�����r��-�lT(�R�+X>+�CjV=�OF#k������D\Z�=`DC�pFۮ�O�osj[WJr�3�.��_?�ax � ��������VO� �+�}�д�5S�}���/`��Bm}����%��[�$�Z����[lPI����)�l߃�Yʧ�|w?w��h6�sS����֛�e�\L����S��n��hwHE���5����#�g�*�'��n/����|�1��:0���i;�Pݱ�|}(W�> g�7��@Fc�Wb�>o,�q��b���-�q*�C�YsH�+I~Z� ��5���)s��iT�I�P�3h�o"["�L�؂��\��z�p�FS�)c]ʷم#��'?#�T�x	�l�\h����g��d����A.z%�28���2�ǩ.$�P��(0]Q���e	TM�N�j�.�Ɯ`�݂f.�
=��NH��6�P� �{"[S��^�$�l��㲕j�h『w>̮L��N.!a��EM��t�����i�H�nb��-=��fz��
� ���#�d�P���X?���*�7�Ͱk���2gv�u�;������L�p�M�pwX!v\�E����n�Ļ��3CA:�6V~����}E�1ɋ/�X�Pat��������!����G�*���Y���ާRB�z��z�������<�_��"���$�] �5��?�_Oe <�}�Y�C*{V?���b�9�O����ζ��
��Tɍ8	��67F�Y�㔍��BE��O$����sit	��e�EPD홃�aI{8!�:�qa�,y�Gzz��x%��T��ϸ���{��0����"����SŶO��Gk��A�[�yd�F���ױ���R� �)�F��EʪT�+�������pp�9)b�Z:^��p�ޠC/�]R4�$��j�s=D�X����P+��-���c~G
Od������U�[wP���=KǺ��}�
S�Bsd2��R�r�E(��0&8�����c��G���^���P� T֊�"��\�M�H�!��/��Q"�{����iB)���@�1f�+C"b�'�=4�xm��������W��mU+,x��S��|\��-c�6�]!n���+ָ�g���$���H��M��>$P�����L.����ɘ�?�Jfɛ_���
��`GL�.���3i"T�>B�R26�lRuƵ�����&�g�.�ւ��@hG8'x���;h9}UB@ *|-fæR���?�ȵul�����fe[-p�׸.�⽧+��o� ����F�X	6����{��U��t�[��GN�"KG���D����~�ߞ�0�v�$Ղ�����lJ�������B�~�@������\wL�|]���SXU����,������g�p��XqZ�^��2�����=|�OQw����le)B�X���U8X��sl/.v�\T�>5��+�y����#��)VX�M���g��� �&r�1yA�w��#���׭/��ِ<XaH$ �K�_JW�+��B���2��j�m�="&"�º*�ب�J�yc6*�*��5eS�
�i�ǁ��;n˾|: �]hJ^��+�r�!
S4-��t��"�
�Q~\g����qŀ��ԅ�Ǿ�=��g4"*���G�-��=$�-�
C7q�i�=M~��U3p�9��&2Ub	���-�c��4��[s�d�oH��6_)X�犧R�q����u��T�W�����Z_�� �