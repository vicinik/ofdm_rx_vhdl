��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�#���[(��x�o�!F�\ܔT���A�mK�y������=�
�1�ge�b�F�Fk���5��L��.�o�N­L ~lt�{���]Z9�W_)J���8�#Lɖ���&?��=��D[�p�o���"+~�]M�j}�ɨC�SD:���iѕh95oVlQF��E� �+I,��K�tx*A�mJRx�т?�?�J���}�!4�=��]����cA+zf���N�Rwٗ���H؏E��VEaZ��׊ ���Q*��z14�CU[x�PxW]��2��]/��BvЪ?U�QzMo��w���>�i�U�n�鞠Jxufb�b)4}Bi��#�7%���smn�/h
1_8������u�?-Av�G�xF� ,�gΓ��E�[�!������Qvz���dPĂ�Ϯ����|>����`u�J@�{�G_e�\�/:4��͚�6[�v�����N�7Λ�,���򓃯C>��}I�t���Xw*����d
q�L��?1?�թ��б|�h�������!�R�M��͕8��h�Yt���v����n�&cKd��N �m�e`#y�F[�&����Ԁb������Ums.�]�3}o���_�L�u�r�<���>��/A��HJE��>1�
�VDe�Y��\�yQ�H��[
7l��M�{&͝�!���3�4�&.8_߶�ȕ��I
��y�\5 }��w���[c�u�
������In�5�OmM'�[�QOrsNLN80 �KJ�ڏ,���/�*��h��FE68�}z(��>sN1���"��W��bT tW�*00px7X)���o���C릶ӝ6$f,CE	�b�<����F$����z��M��kG�Xɰ��O����RN}��"�S�8!\�I�M-`�n��'n�F/�{� ��r�>1�B�sH�/-��K*���둼�T��>Z��Lԗ�$����leT�,��][����;9.⿷ʒ�����b��4Ă��*$��ŭ���>�k�*�xB�2�E'_�n�H^�:qD�Z/XӦ��C�٤�X�ne��"���Y8Oۻ��}R^Ǚ
 :�8�}��D}Uת�э,Ą��K?/ə}L�b2 ��J�&͑�l��Z����Dd�ޓ����o���>��i�K6h�  פ�Y�lm#�$M0���fXϢ�ی���FF���k1��(\�'��ev�X"}X&�+p=)�`U2���jl�Ѹc�(�@1�~%0�۠Kc@���}�y���#����&D��ፉL	ζoD�֨��PH�'�sm�7��Vs����R��-UZ�߲͛��Tҥ�I��ϭ;��V+�մ��3FQ�)�{�_i|�� X
�����j��5��+��Q7D��O���0�d1f����L�E2�|�ғ-���/�M��e=|#��?�(	�nO��y���Q�[�&���|�p6�.&���a�"�~��"��5>�_�bg�HRؐ�������`�Q�E��Lj,m�Y�9�)oq#)�IL��)�*PO������#\��/!,�c*6��2�I�zOu�ݖ�u�`�੶p�#�#���.䙟ݶ�6����Kl	���߃�>�?٢�/�J���}AbA=Nh�:�.�*.���2ͩ�FfcQ9���W%�Dɘf��b�i�'��NPQy�(t��$�h<.����&���-��Z4���0q�-�>�pq0�|��_��Aʎ�y���Z5"2k� #B�K�iLg�'�02(�$�І�`���uIRv��X�ϊ��8$Н����D�M��'m�5O T�l1��)w\�H�ޔ��K�q�s�;�:t�!?|	�d�m/��Rڢ�T�In�L��'_����
]��_�r�d���� �Z�_���m�����3�Ud�{���S ��~Gis� C���@�B���ꩽ�~N�(�:M\��0�耉:N'����.5�;f���Ș@r��#Zy�� ��
اð�M%C������=���'	iP:����߼O�s;!�,Й�~Vy\Zt�B�����xf�[\�zZ[-.��R���/#Е����S�v��絔Q1	��dxE�<>����b�o֩�����I���K�~Jĉ{�r�q"a��t�T��FW�@sF^��ޑx��ZB���]j�c�b���>S#����}�yP.���Ы�)��;ʐ$��:�E�"�����������ßL��+�z�B���Kn%���kJ�P�6̿"\"�[�=n�ĕ�;i8}+e��՘:(5�O��,�U�kR&	��~��R\��;�0�s�?n,���Ro�K��݃;�^�?�A�9��B3J�_8�{*ԋ�3E���*iODɞ�s��e�t����	��W<j�v��1�s�\ԓΝ(�����}�
q-�nf�z��$)��'B���QI�#�Ť���~�������y�G��!��
1vF+���3��ձ+�F�&&���%%D�J��fO�.nS�`�N$�N��ے��ͦ��MT�G�u$Tb0��D+�O�z��
�57�f��.T�~`� �N��=I����G8>]g�Ϝ�@���jLg�n�a&�W�rȓ�Z7���Q1��獏��M�ee�n/���<�\�YW��� �n�f�7���n�p����UX�}�f�+Z"ys�E�
*��e	�Hī�;΍ַ��*%-���s��9a�#��A�c���[=�^�C��G�	ɚ���:��y÷��eMU';�!�����i�{�]^Y&n����Q�4P6@ik�,������H�Y��{*1���	�� ;�e_����~�w[�Zj0��ezG��M�2�/�e��z�!��4a���fg%W���g��Y��&\�@�^�gzύ�Rx�\
�'&$������:el#�.w����)�7M�4P�ho|�"$5�fM9��y��ʉŐ�N[��ţײ=���Gޛ[&���ƛ�{o���,H��H�S�mO`+R�}�FL���B�ӝ����=
�����-��������L��4y��#k����<b�@dʜ[;�d�j��%�:t�(�T��H٠�@�D0p!*�[_��d-��d+�pb3�Q
�9�G�֮��h���>s���5?�ܮ�
Nl���4f�4����J*�a���o���$����P)���r2��7�*�8�ъQ��ݐ��C��:R�}@��.�0�[�uH�\��/����_E
X�L�$V��#H�dk�%A���ؘI��2@;�l�̶�������G<�!;�C�k�[zT�q�a	퟽g��V��?r���
��х�/inw�t2QT�Nc`���A��Ct`;���hn��[�$��Y�3�$zfM����D����
+�9R�|/����9kQG{h�di����6*�
���Fc�Ы��C ��NS������m�D�f}�㥬�7���F*G��h�b���E_��`�S��y	1����>}�0lV?\�:�j�,[�ӫiӓ蔲�mD���R�/r`���Z�H�*���A� ��|oZ�Uv1���{q��W����˗`��ߣ�u�i'�nv����m	ѧ��[��� uϞ)h�h4�ޣ�K{-�]��cI'�%�����֦
CJ����}�m����fwO#臅1�@�Jը(Aw7�/�[�-��/$���{G�"�q2���T`�0�-n�h;�f��Ў#(�-c�G�3'j�����
帄�,����Y��hܪ�d���<*���}�"U,��m�?��{U>�ǒA�x�_*�@h�1dU�=�3��w�J-����o���Qy�zr4}�t0ė�#��P��tW�/;��K2�B��4?�Ĉ�`d����k��)O�G+��������.!��!1�a`t�e,(���|lbJ
���vQ��1�Gy����%^״*d�/q.91K���[)$���Z�_W����g��5���:7�Q�E�C�<��G#��p����coa�N$�V��y��h��/$��:���4��d^�Wu�����F�^��l�|Z1��i+���{�V4@&���ʹ��DT���p�E��x�������7������%lT��E����"}��Pw��� �/ǘm�)��Xa�I�χ�:��)���ļ֣��*�ŏ<��,
=@N�����Fp'>�Ŵ�ˮ&�-����@�����q��n�yl�f\WSwH�jR�Z�G����f�ٮ�wH�S���	S�`�#���|}�14�I��/Y��nބ45��@��Y�y�E�Iscr����]>��F�젦��� ����
�� �"������g���>��pfI/W�*>r:&1��rG���I�Pr��۴X�k�lX�e�w"�D���;�n���=�ys88b�j��(�^q.2o4�^6�1�Ib�h#�l}ǂݵ	OGDm�]�¤�/h f7H�n������x���s��Ԯ��jT�5� �$n������n�=���??�V��C���~ݸ?���D�N߀��Y� �\f3���&����7�LcT