��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��I��Ј�r���a�=��sM�O��tOZI�`���dW��L��7z<('G�a�Q:���d.�Z�Aè�� d�=�l:��k?��^�<>��$QԧB��\ +jv����̑Ϙ�h�v����ؗ|��Q�ֹ���X�H<9/}.S~(4��6kv�Vq�.��̇3,�-w�d<�=LA�������h�fM�-]�F�/B$$�$��!����cb�ʫ�ʃ%�`z��请ec9�B#�7>՗�f�x�W>�MO;��"�����q�h�֨���-\I��$�c�-���>�q�/&H4�}����J��V��u��vs*���
sQx���YƼ���O��1��.���@�98�@��T���4��T�K(P��U���"z����;joZ�=���F
�]S�T�T�K���Ķ���Уe����K���o]�+E30	�����t�����%����N�!<ȏ�S9�ẁU!�`<-H���G �����x�#��H�S}mf_��_!�a�㣒�GL������R�th�ZE�uX���Vw��U���r�6�EH+B���y5��⎥��'���Z���fY�u�5Ƙ���ܻ�:j������h ����.��������u��ʊ۹I~F5��`^;��W��<͌�ѽ�a��
r����m����_���}�Nn��+��m�T����p���K���a����I{��vD��ˌ�W1���E4��^3��ɭ�@�y��נ���[[
ʟЀgqN�Kia�i�,F��/����p����P b3�p�lP?)��n�7�R�=%����49Y����*y��Ώ7�3Y��2�m/�.r�ݕ��m
���_�<���#��^L�m|s�S歡<�R�>g;��+��CN2��+��!�D{�'���U�� �S蓸(��L;���GsC��'7���&�����u�ɇ%<ېM2>�@��y������,���+x|�6]�EO�0F��=O����j���f��k,hy!.��|C�l���KK`e�%�����(u
+�9���B��ݨ�D-`\��� ��>�ً�Z��J����Q8� �́@�� *ݭ�"q'CO�@��Rt��+|)�]�v3�����6�Pa���4l9K^/���I3"�"H��P�,.'/�׾��Y��}��x�9k�(��/ј��3R�/{�����2ͪs�^�A0U��J��B�[��#�Ph�q�ώ� cB3»�%+$"I|(d�C0JK�uĦi�E���^	*T��r�8�:��I�����|s��7�aq�"�w�(0V�j�,�6�g ��w2��?/�}ޤ����i�:��)�H�� ¾:4�A��ܣ|b����yI���	8���Q��󳗌��K�@u�6�>t=/OE"���X�z�e�Y�-l1�d��� ��"4߱�tI[��mt�H��M��eьd��L��I�Y��J�{=@JM�*_Xt�Q�??�Е��P%�iHW1�/���]�V^�h��9�P�sҵ�W����uj�NOh�۫F
c��0��3sf�kT�m��R�b3=|�hW�,z�ŝŅ���V�l�J�GT���u�"�Ҧ�.ױP��\��(��]�^Wġ	?��=���m'�c3�|~���7q�4�^��/3v-�FbK�	v��"^N�oӟ. bU���"�>�q\~�b�Ӷf��ј�xo����Q�e�Y��F�'�^,��ˁS�/_�Ň��Y|P/f��
ANkOB`F���]�U��u��ǿ��AR���O3�d���r��ͯ�XL�S�3D��h\_��z�C�>6x� �"�LU_���<��3wX+�/��s£ЂǏ�������ooz�X!=�_A� �����D7*��mff�/��
��A$2O@.�'U1L��SΈ|�'gkJm����~~�LR��97Oŭ�c�mp�~]�U�LP;�Q ��'���c} s��#�
����oM�I�ٔd#����m	���̘ެ�:�.�"/uR�i�X3��� 5.�6�1��X)5tT�n+~��G�߻�A�Rl�lgx����Ȁ�Q{z(ə�3BҶ�-ý�-��ga��(��i=����T��1�Y��b��3�s��]�4���wP�̬��P.��	~�p!���B$�<lr�k����aj�� � ��i�`�~*�_����z����
ӡ�����X�#�~Qm��Q�lc �:��\lV2y���,�,��aa(X_��b1���$␷4"E��1_(W�yA��R��`|ߋ'������a����N�p�n���S�0,i�ǒ�!?F���?-���f �5�i������Qg�h�Ys�	g9+9N,o�HS!��<��qlP��jJ {�K�@?�un?K�Ӧ�ؾ��l@���F��xd�=�`�ÿż�	#�*�U_<�+s���n�_�Q�@�;�����Q�'C�O�JG5&#aQ.w�X�__��q��sbܯD�JvQJ��t� <
(�� t�6Ͼw/��E��3ю�Ô�ך�XW�[Ӛ���0%n.�0c:���v���+r,���xg��KO�|.�g6�j��;�X��z2��f�zr���;�>��,a:%%��	�r�!��n��]�0�hlY/�Eu���
�C�]�9j"��@�Zz����r~��v�"�ˬz�>1�t��"L�*\�l"�#����D#���_,�������}���zԺ��t�U,\s��G �V��Ez�LB}7x�a\����>��������'v�2F���m��{�/��x|��6&3�CUb\��R�&=���! ۧ���0�� F�p6P�(p����P���n1s��#�����F��0���ڿ>�ټSc^I�n�LoV�d�V�a�ē��<!�E�\\.��w��հ��42+Ciڔ,#��ڥ�b9/��!���s�P�C{�=��G;v�4_�:�o�W9����	+^ƞ�Q.��Q��������rs" �R���GX��4L�����(�-�N�N�'���:�/�~�k�Q��-Jſ��+Z����iX9R�ȈP��qhr��x�y�w����V�d�SQR���)�8�����Қg��P�`��J��L* �d/�I�8�ї}"�bA���k�G����B1s]�w�&9��5�Z����s�0��ɜS*�ɫ����U���N����#�%��B/��Y���0��ҋ��
�a�nuuQ52-bh����f(�^]��(4�OvVO8v�N�.����S?i�����\�Շ��"�]-�,�D"�v��=�*1RI�q��L
���'���% �P��*p�D��&,�f/w_B���*�f�*�-M��ug�5m���J��]K�-��E��@7#������8tr}̇ ٲW�����-��E��yw�����B6!T��Vl��{<jW(Q�־2�$o&����.��e@<g����%�!�t8PE67�k�r�bY��YF;�����<�P^J�]��~�ب��!eObJ��?Md��r��Q᎒�)�-�\�����D�w3�P2�>ߺ��9�����ć%68���8p��YP�C�#8m�(*�X��~'N��Z����˓X{N��E �j�{t����/�b:�4�u��ʇ�gN2O�p�zj3+\h�6Ҝϔ·4�ضՌx%�0�¾:����g3�#�+�x�@#YVbf�gg��4"m��9��0�V"�͖��7����V��+��:������$z�0<N���M�Xߚ��w��}��r~A~y���Dp�>u֮�
8���4$�Lj|�:��ۭ����~z�&����j^٣��[^=��
1�,s�[���`>��`M�~����4���ާ��(MW?�zV$B�*!�AM��@Ƚ5d- E�p�|��Z/�+,
�C���TW���E ��l[�ݤ�O��mxo<���=�u����{lNtSٰ�a�:�
\�ۅ-�m{����}b�5fפ�u�ʥ�
�Q�G:7�}��&��{s];r�4�#�2�J�'6)1���n�c��ڼY��8�]�]"%�}ȄR�Q�8D��: �У8só�����\�Ȁ	�f��"HHP���S&�|73���0�ϊ1,t�j
21�䀕9���`��)^~[<�%��y��h-W�cU0���x�1m��E.ը/M����T�TW�ݸ�/@�#k)�#W����ρ��Ko}�v�$�)������I3Qpm��|z�'f-� <C����l^Ѥ�W�P�2iT��%�;8�y��k���.��z�uF_��V���$�4����E
�9"-��VDx3��N�LƐ9��v�G�{ޝot��K Z/}���M@J� !��/�_��8C�_�����$k�[�K}�kZͰ���N�V���d*�3[;��oK.aIא�//	t�N\k��Q�>Is����%����-F"��g���a�$M�shi��;��
�C�ľ.|�5*�@��-�U��6\��9��EI�������r�N�0�T�詩z�湢!W�&mq��9�T*��Y��P.��F���'���u���f��I�.��:ٟ���q����CE��^ܔ.=l�9��(k�R�w��'�>Cߵ~��p���#��c�χ����]*S�@���Wb���j#�y�Gh���#=ێ#�U�J5�`H�F��J��NR8�;CBY,�e� �4�H��d �\ɴ�%�@�|�&= G�I+�����H���K<�']�)3PbZo��>*l>R��;�ǫ�><
��T��5,�D"�6Ca�ƕ~8�P3U�Y�Ҩ<�f�ON2���'w#u��hRuĸ���n)f_�;��l}p�3fA*��\n��Ue�Y��;߈�n���<�M ��J,�tl��ZU���h��
�JK�8+e\^�;��4���k[��"~������Vy��|�B�����:�a�햬8���ur�Z%*4�O��]�i:�`��pGhL`��y�-�@bY|Y	��`rZ�r�����������jA�����$U�"�A68Ra����ǆ��g���^'�	���W�R��m,�D�}]�[	�]!��W�5�v��-�=p�L9f@���R��?��L�������tt��V$�<+/�S��������ژ�6rhh���|iU�_*�����-d�A�������ˊ�_��簅�0�>n�P�C;���{h4������|R6#���~�`H�i�8P���kƵ$J̏ԭ
~9� �"n��s�EN�t/|�(�E�,C��g�9� ��T�3�iЩ�Hs(V�ԕ�^�1�	||�'B>n9 ���#/��3я�(
�f�������j�Oq��C��d"�D��	##2�]b�in�W�j�ZC�b]bD:�J��,^$��YJ���q.�Բ�u�"�$3�\z❰v�ޓG�#z	Df�Y��,�s���x�*Sxm�|��E7]pZ�����+IƮ���߃��v/�>�*~^�ć�-*X��n[iE���}9:�'"�����n�[�U�������ӷ��/���Q!#���1����v�f*����Ͻ:=��ܤR���?�y;���)b�F.��3����I
�s���*��gۭ�9�u)Nީ#CM4dn�MZ����F��4�?tT[2B]�p̽�`^�`��U%���O~��fc�F�6�uȯ�#�H���?V�6
M6$�����ϧDּb���"wSt����xך��C^dxah�Ip�3�#˺��բh�(�0�0�0JwYo��	�]��G�շ��NMɮ����y��MNEl2v·��EDG��xz�P�N;g�{����1Im�,�Yi����ш�k���|J�/E�ApQe�Y2�I3�R��22���bwO��J��ҧ
��g�E��e�@R�UL$m���+Z+��b�n�,]?-��(�v�Y�<�]C
��C=����[�unT����p�����"�̯-��KQ�rB��<A���[���~,�SZ�|�ǆ}f�@�ŏ��J �������K�|r�{�_Z�)y쉰���x���׿�oS��:�
߰���7�#Ԋ��+]��udBR\w����}��:���򩹓���?��'�Hi����3H�.*��X~H1����"5ǿ���o��C���V�uY����<�Ƭ+��h��E&&��WW��M��A��7ͳ)�%��~aΙWut��!S7�����$� X������ugj��>{�[76ڍ^))��|cFlq�=V{�Үjx�/��lByRߴqp)d�u�@���8����|�i^;t�p�u��N������w��4��ytu�LW�ř#���Xҩ��u$�7�?uXi��+��Q],I3K�� ��#�VCu����-֖���D����� 2*h�O�K���t�����r� !jg�U_�F�A����w�^�
<^Kfi6��J�(�r P[�oȦ��A1�V�h��.:}LYa*0��������؃dGoBR*�� ���G|�s��9w�� 粲�nGr�"o�%ma6�C�����lS3�y:��XX�'%I08R���wwZƐ7�K�BA�o��;'+ľhDg�Ia{x8Ezk�����v����Z����Y�g��(�����<�*8�G�$Ôk���Z��$7�+H��ݫ2@��7��^Q�՛1���`��9������C����'�e��KTc{�3��!�@"����<��%��>��}�F�[�$:�s���cZ�=F�h 1]Tr�E7>�J� (����a�;{w����67r���FE�o=��P�����"+���'���I�Gg�#������v��8�a��/�?�na�$T�L?"���ɏd��e��<<4�3i�B)�r6i\pӗ0|�ȍ��l�ڡ�����B����Qj�3[���^��d�Q7�ہ{�Cq/���e4�b%K��Oؼ�����0C�x��'�!��&� �_l�ud�q !�kګ�m�i#�D��5~RHU��t��JS~!z�J��!�{S��gR}�	r~Z��0�u�-m��-�B���G���r��l�kKDe�%Q��KX1§����(C���ZAE���}�;��W���9����@0�I�oŬ&�<��jK	S�C��/O�pB�j8NT+����1�E�t@�K��^��)!�}���f�ͣKiZLw��1�{���J�5}��]}��<��ύ�W�]q��	H���:�v��hY�� �W9؄�SC�`Ф2�I$E�?��2�G�������I,b#�1!:k���^GL�҆u���A�>�5
�?'�&h$i���!������Bi�s�és���9�x�����o��"sɣ>��+�;<9��8�R�Q9\��ewx�m����z�O��w|��F78!����ڌ�z�T�uG�A8Wo�����DSe闐����.�"��^����F�q��Y��2B�)a~"����`f Oo�A@0c� �q��][a�D�n�����Эl6{�u�<�Hb#B����b������UBP��՞i��?$��/��u��5�:-!�-��P`�J�r�w.�����x\���6P��hi�z�I��j��"�� �j�(f����9���@��H�FR��D6�y/�;})�~/Fs��R}X�ւnX�M^
L�I!���ůe�j�҅��^��Ը~ʱ�
��y����
��K�U�����k�}5X��Y7�_x=�-���V���_!ōu.��``�<�B��w�C���̝��ȌBO��*�0Ɉ)|��	��ϊfc�ı�;JRx ���i��r���7H����1�4�yH�0�
�J7QF�!�̒b;G��-�
�F6�"�䦪�p�p�Bm�b�ʀWf�e����Ϋ�p�&W�t>��,#O�g���q�=k���%ng7i��g��?Cq�o4��^����L�ඪ����V�L��bH�|Y����pr|��{�M�o(#mPL���e�bW�2��S��ًi���b�����A��\'���ӧ6wg˱*;���c�]���apU"e���:��r�FE�v�}��N��!{IAO·�-��"���\�ˆ�<�U�T<���Y�ljV�3Gb?���,�k{㷍��eR����s�-~�؜�<�(�pr�hl�
�=n��Jܐ�i�
�,�)M���d|%՝�Ϙʲ��@����7N��*-͑���&>��}�yE�2pOؗc��01�U�T}��my���3�3i'�H�J���c:�	�ԷK6@��E�VI*/v�<?��#$P*�L@�/��ve�?>�D��_~�C��jo�׀5�����2	��y�q]����0�,�%���Y�����ٵق�����!Џx鲌�V�������WZ��m8U����\5%vdU�8���D~�� �)/;s�&��ݓ>����]�ҋ��'.�5��=��/���3���%�#�?MQfF�m�[�iJci>�׉H
�s��⎎�/��*�#U��q�Ԁ �I�W�9	�7�.0{a��[96I/D�p�IW���"?F�w2�/��J��|u��phbfs�p�xa��8��	^z@�� sY�J�,��� ���H}^�x��~���J0���RC��JyR����YP�ʓ7iG�儵Q�UF�+F,$�B {�^ڡO>1F���үN�̗�?����hx�-�/Bv
p��\�̪eL���-kaH�H]L�a��'����Q������d��C�K�-�r�:��c{�1�+X��L~��&��Q��?���?�Ã�SV��e�;��DS*_�¯�t��38������F���\ptR���38>֧
6N9 ���P�ߦ���C��X�L�"��f��z�>�u +���5�^��� ���V��?�nr~ϧ}B��8d�o��fW(T��-����̆�=��V3�,�#���OP�6��[��X�����W��M�U7L��;I��Q#��A�����(�\�j�PL�̦�0���^��}�ʃ@��9/��:eI�rԚ�N�#EJWp�_Z0���x
)���Zwo�?Y�"Iب{K�X��:N.�_!��t�O���8�` �7�х4@���#�%t�Ro����-�*�hL�� [̧�WiU3����T�h��}�#��	'ԊʀR��ԕ���Ȍ�b�Q�����
qe��~�ԉ*x�I�3��u��u��,�W�y'�Ej-��h��| ���{�-�!j�� �i���j/J)��A*�go,�7>$�S@M��f�2@'������+���aȗ��5�&\��4��R��X�_��e���L� �pX�6���1�_��.R�u���Ey��g�ْ���ܬO�Qf�@}(�(�*��ꢕ�qպ=�5�2/R���]glx��k�� *2�
̉�EtaU� &��E��utuH��4xn��a��@�pl����ȔЯ�w��2�qq9��]hל��C��D3�)�݁D�5�~�<��tZ��Q��b�<,��OV��Y7áss�>
��J`�C�4ޔ�P$�]Z��)�sq�q��1&������	Zc�r�E%�Z�U�+����iw��3��T#�<�"%�J���6��E�z����Ð�ՊP�����H���B,�@a�=6�k�M��Ma��ܗ�E�W�^HK�x�k���cN�}�+�H�T���[Xs�ީ�=q
���J.e����&� x�v��d�]�6q	�0��]aU#�x��%ϸ{(��d�t���Š:���a]Cq�Ⱥ�"A�)p�%����1,Ct���V�@R��
:�,E�{��yy.�A��)�D�>j�S\�<���9�o��p*�$��`yia����O�]��S�F�%�+����_'�_l�җ�n��PE��1 ��H�k�M�Y�R�A��j��W��UW'�@];��7��$��q6���&v^�q�]�s)�3�����`1��U�����2�:.��G����Փ��+�y�y?u���XA�ҁ	�%?�ہ"	�en�G�l�$�����t�+��-��eWL��p9�#2�a��C%���"���
T���'�<ڄ���9/�I��n�+�[׌Ω`T����X�*�$��nX�H3!,�����y'������yF�yS^B>X&�p{���o��}*Id]*iV:nfizG;��OzG�(�Ad��!+��a�����%��L�Ot��b�h(6���P)�j��_ƈ�H����s���9���96&@��켍�x"�6�p�G�����nC���\ӢH�8s���,U�����Nx��n����:�˫{���L��n�sO�Y{T[���Ք��2 #B�X�y�K-7�����Q8�����1+[}+3|���C���m7��%� ���eu�T�B��%���G����gMK����b������1�Z�v��������'�ʚ��,/s��,�4�X��#[�R5�c�H�X��V�֮}7����e5�wF��G\ؑ_W�.��5����8��rQ\[�cg�mG$\���5
ݥ�!V4�q�_�ʥ��]�X�"�ˁe��Y��]jO�W5tE5�t6L#�彴��e������K��"�^xq���c�����B�"�F�jR�p���nxc�G'�K�˝�t1�Rm}#	"7x\\�l�[��$`.x�m���s���q��� �"��y�^�]UL�[k
�ٽ�e�F<�1�\���w�I��e1�� e��DY�}�Eҕ6bS���i�
@��{�vTm#ݕ�A;s�W-��@ib�r3������
r�n���Sn����Q�G�wv����P�'�
 u_��t��U�7��p�����&�P�tc�m �,yA^��6��Q�����,[�l��|:��O5-��Le2���eb��k�<���������-���pc�������aW���?��;W�^�[\�5)=XO��+AB�>\Bj�$Iơ6���(���l	ې8!SP�8�@��sB,jg0a���m�����h���g����ll!{�Bd8�#��m�J����)�!��H��f��e;G�J���|J� ��P���(�����Xl`�:KG���Y}��m��DcڻB�Ƚ#��g��߫2�������g��3x�x.����%��\σ���2�����0�pD����@�;��t�*�Uʶ;���4���8b���W!����8�o���|]d��Љ ��P�m�l��m�'��Ul����M�G/��1�W�b5��C���I0̛�c�-��[��"-�/��+������s��/hV�GD)p� `������3�	=�"�/���f�9䅎�_����"�鹤����٬;Ó��B���@���~>�����\�:�F��}�=�q�pKC�������ڰ6����g8�Q�O'`�r�4A냤r�_�� SD��_��NQoT�AI�����G�q��cKr��5��M8E24�cE3�u/�+��͏�(�@|��(lr���N�*X{�������Ԧ�P �����6B'�r��hS�i�~�킱�:��������(Hi��w�H8��@ȹ(�:�9�A�]���I����M�'�>��|���r<Q@|>�N����)���/9L�����Z��w��W'��PzUy��h]u�?
��
5��4��B���NK� 'Q���/`�M6I{�|��%4�U�� NYJ�QKEd�oY�����O��7\�q��|'����8�E��ʋ�����_a��[��י�F{���;C��:�o�d���Y��<3D�-:5��C�V&��u���`ň@���V����3�J]/s;���*-'z�ۤ�������.��t{�>����5b�෹��Z��vG��r)�3�m��-�a@�~�42l�:��g?W]���B�+=Xm6.M��W`�R��8AQ�Q�G�MuOI��wo��QLPNq��M�P���5i�~u�t^o��y4��vԦ@A��]��G��e�%\M �V�M�^R�H>{�.
TF��D		�"#2���W����0�L3���#�!�QPa�e�k_x�&a�Y����Gy��Yn䁦�z�a�>�}/����ꖭ�:���sf������`��Y���iކ�����'RD�X�����"�:�qa���[]P�;������5 �_�.o$20ϖ�Ͷ�w�H+j`|ĸoU�cՂ����B��*;E��"��^;3��խ�O���Ӂ�J��F�Y���%gw��6eߧ�J�m����w��eEEο��&�����	:I�֢m&�vI&.�6kλ$6)�J�~O}7��YH�С�u�{-+[-Z�� �0����x�5�H�	� [�qr"�ڧf�8�O&��rKEѢ#o�R�7%���q��>��:�-��w����а6��|�'�����^�_9��||���||�F���,�A/�sn�*��{�=�%a�^�/G`.�4+�H�u%Z(J�nb�BBD�q�`V1�@Z!Nq�Pj���uY�͋�s��/~�^����/��5uU
��h�A剽Z�8x��N��Fi��脈��@`E:�R�8�WCF�F@��\c�:���&C\M��@~�ѡ\��ϝ�|�Fno���,�Zd��CoU��ZJ9J
��_.�v؇އ�+ꏒ��zj��&%ؒ�����꜆0�f[�ɮ�&Oj�c�[�6a;�[�4�Sst������u#���6ryУ�K.��t�*��(����D�k�b���\^E3h$��nu.k�*kP�ԇ풂Qٹ&0�5I��A
���sܭ�|m��}҂��4��(���۰?- ���g���pO�&�=`�T��J��{nJ�~����Z�y?����1������>�)�r?�jr(�l�����r��h�_މ���)3(W����#�b�����⚂�^I��I��TT�t�f,γwS� �5w|Kb
���}
���Of�L	��0���P�}���!�(����Cى�F$_�Z�	�����G���0�=lih��n�tq~�G�IWq��*��Т��p������؏��qߙӞ�:"���Y�b������5�q��j�ܮ�d���?ʬD�%8%"nr7����sѬ��-�l�vrS�7lGyF y�~�6���V�ן�\twGS�F�7O��}�h%�0�m�%�g	,ZgW;:���Q][�|k�����4p��F��J�l��5.{.���q1�W��J��_�㜆�ӴO����Xb������e�'�<��b���$C�5�}���� �/Ǝ_��u���<ա�k�fƞ�.����k$�^*��x9
g�_�1� o�:潖����-ݳ����0&��Ӆep�2P����|��i7F���EP��z\0�
��\h��Y����+b:#��z��^�=���dM�P����CwE�e��h;��(�{�e���6�'�K���N���֗&L��-	�G �����[�t�'
Z�s�	��~E�f�\�)�Í{���Bߺ������zo³��)f�O��|��W��͞��;,���E@��"��]��{]2$�K�Ҭ�ꁳ�?۶��*�iW֜&��c�~�����#�Z����qc"�i���� �XJ����mk/���~q7���tb8�Rϻj�Z#�.r�����D�"��0J�V$��x��� Ww��;��F!�a3�1{�~���;4?�
���۟���\�;�׾�J���uH����c���q��Nk���g�ư�R������=X�;b�Y�5��e�_�\Ρ�Y���9�C�%ݤ#g�@W:�r*�?;��4�dy�Ŧ/��^�b�V���y|�N��TS���0�Z��l�0����p�A ���oԺ�����������N���(X\���Y�0x?:ґ/2YK)`��wZBhݗ��&�$E';H�,����mQ2��Jx�6Ë�_���<j �㔐~r�Fc�w�F�,�T�D6�$~M��Y�#�q[��(�օn(��(�8��y�1�M��n���.T(����}�+zϜ~W��]��N2��;����Č��#��|����h�gP@�'SA�����{�[gÙPo�wG'\��ue� ~YC��m���x��К�Ioo�v��� �������f7������,�g�̨y�QT����<}"�G�!�����D�ڌ%����h�6�����5�~+;��ݢ;� C�_�S��̶G)�L�ќ�: U�v�5Z޵�˸D���9��t��]6�%5�ʬl�%���jIg�@=�q������٦�=�$͖���k���� U{c�����7�#�|`a����^���k�⮟7qЋ����q��c� r��%�`����cHhMQυ�'X���i𦞎�(�*?/fwfR�EP}���#��- Y�Ԉ�i?���l�qNa@@Ǧ��({��dD;V����!¤�8��]���Op��m�Z�N�8O�E�����b�^DXs�}��X�%�� "0#��w� Y-YP�B��)�E�	�LH $�w�(� �������.�j�x�>������\v�k�kQ�(S���/'%=�:w��|w�T��|A�����[b��5���\���ȥ%�e*�������<�>@-�����$x(AR@�v����e4��B�4�=1J�����}͡t��υ(8�aL��ҩ:��i��z��򶖪�������nK�ߞ?�̹GJ-~%���Iio8㋂+�5��㾐s>q�IK���"O�Fk�0�6�L����s�9�y��r���W�D-x���x3�"�l���k%�V��!y��V(�E��gP���ɡ{n��X�,ܞ����y���nw���2a��S+����f��3ts�}) Q����n�\�\������i���w��n�m-�}j��}����K՛i9E��\M֖�̑�A^��lYy�|Jq��k��ku�Eh
ǲ�*�r�U�؉^z��w��tLw��!K��r(��`�s�%I�׬p�<�@�h�-o�Ҡ4�K��)�C �"�f��z�ҝ�o(J<�5q��	;K�bNc5R��L��P�����	���PgĔaO�l^
��N�.��&�)��?
�ja�?֓��j���
�x���xmM��	�K��˴6��L�kW��o[V�#x\�����>�Yj��$
;^�ZF���!	Q��;��PzEB#��������8W�m�Qy���e89���+x̌IV�h�nD�nY!b���58�MIO��0�?�`��(`B���j�[��m����D��155���B�yX�\a;:��z�����>�?�)��ܲf�ڨ�I�J7{���!�\r��!���1�M��h��>�2�6��<�8�E1sEˆW��r��P(7�Z��o�N,���o1G��np:�4���|��ͮ���\��6�X*�����zY?*��_yW��]��y��;v%��B�A;���O��[��͋z���P H�\=�x�s�u�|�Z,Uv�$.�Z�2@,I������\�ϗ��ۜD�ʣC���$��,6��ϣ�6�'9����PC���G$�Ȅ�WO�L��dف����s��>}Z�_.7T�$�v���|��7ǭ:?J�@�M>v�
��[\)�=xL%��:.faG�<5���#��V�D����*���h�s�^��i�Gy���e���͌(�]���%msYy�s�Yr.#�H�因9h���)�dw��2��*�(]2?�{o�7��S��r$IJ�VW!'N9��#yH�U��[?b�PXs�\��7%ٞ�Ҩ�6�ͣE��=�xC늇�YE|��a��e	U�p��9QAB��o(�����z-�J�O�[Y� ����)u�����#�9�D���[Kv~�໙���~�O�e�I+������#��h�<߸�4ǆ���T�[��r�4�Sd�*��۵��? �8��^�V/��(PUeܫ`�a~Vm+A��#z .���Oq��"�Aq�lЋ�"���!yP��.l����⶷Ai�#��U�)�8��{"v�LZ����E ���������6���O��~<�+�\fI������zM[�j��4a��֔_MJ̢Y���`�/	���Xq�O�t����loYk5����b��H�z6�t�Ӄ~]H���K�9����G��Ā��I8S�[|�.�JLqH���b���AtĿɁ,3V�1�����̽T����c~��Ŧ��)�m��^"m�%��$/�o�2S����N%�#�n͟e)yJ�ӪKw]E5��\�J�=n&4r�J��s����]��)o����@b�J��²�����
�f�o$x��{e�*&9����VO�,�?8&�7�AWk�W;v�mZu�)��'��f����0���	�����Q{�p���>w�T���R�������Ĝ��ϗ�d3,�?s�ʑ�����8{9]yA���+}��j����^�� �T��tG/%x��h�2��)t%��&/�7p��}� �4�F��+��ɤ��A��-7T
�����԰0Ϸ}<���B�> ����ؾ��l"Q��=�h����cψ��0KVm���o������Òa�Q�J�	a����v�/�q�3ТB"��љ��CY�;y�����Eq��d����C♙"�����?SP0���'��=�Z�6�Q@oXz�}�1\���n�)���^�]c*c5V�6��m��5G^M_�e���1�������y�.~����A�����Pӻ�А.��ָ�f"dx��v��-��X��lˣFN�/'���Y�8_�MD��T3������x��U�Y[�PM��l���2��n}s�>y������e�f�2�{*usݒ��`D5W�q��� �b$��f�C<V���>.�p,u+���N�����z~ݱ~Z��`���w�ܴ�"]��Ո�.�Zw^�-�+�
�G�3��g���`P��:�	�pn�%<�����5�eS�`⑨NRo�,"��hO�UXlvIgVh��mtI(�����>;�
%r󦷎�ho��B�Ib=UQϡ�_���F>�X�K��&���*����5��ѿ�A���k�cR^ ��T�]e�e�7�[`���?�G՘
o�g1�.�m��D-{㛅H�@7���)c�Tt��Qb_=�c$d���t�k
rRٰs5�0�E��{O[ѭ�Z�Dƭ ߢ�De��L��KMT%��PS��e���I\����e�!�ٲ�ּ3�
�s�E�d�P���ٳ��.��"�T��#�4�ʲG
��Y�H	[������&!ש^��&�l���S��>��#�K��O���r��N�I�/9��� ���0�f�vH.�0�Gg8� ��BpFZoM��i�P .�Cf�x�Fg�mV(n�5�j|�E�"�*���;��/^D�b�։ N:t)�yP	;:|��6�8���8��,� �9����+C`����Zz_�U�Ⱦ� �h朁S-`�BR�zߠ��=���#3c)�Y���\��y���'e��T�'��/?%J�%�ϥ�+tϣ�Y�Dj��-�s���mi��rWӚ�F}8*'E�N7I{�р��@��z��['�ѽ���W���Z�~�k�Mz�{�머צm��1�B�!v�.����(v�$[\ �wg6���Ӟ��ۉq-d}��\lsӎ��h�E���� 7t�le�Ԫ9%� ���SK�+#�DRJSǫ9t�������Z X~��d^~��Uh�	1+��"g5_/��z#X��xiE4������I����@{7�RfN��eرcu�(���|�Qje����a|��-�������S�(N�U�	/3���D
n}*�]�u�t�x!�x���x�c�ɗd���� ѯ4��;:S���9��<$Kku�{���Ε�!�@Pyoк4A�Ԥ��gR~�Jmf0�T�`�%4��0�61b�f�-�?5�e+�ci�I�<���9	�@� Zjr�5�����k��he����brn�u���Hq�%�8��͜,�\w�׊�%�s�9)=��*�#5�f)�V�s�G��傴m���2as�.��뎂S4*
�1E�_]&N�QkeD��J�3I[��3SreT�'9�fԨCݧ�!J���df�`~�Sf��v���vS�M3�XَS��IeI>�~d� \�C6�p��gr)WA�y�XzC�J�"����W&Vũb,�l2_H���C.��%�N���ZļH�5�n�E,J�B��x�ƙ�-�M	s�d]H�>�&�����1S��P<��;�ܢ�E�i S�JH��H��Hd�i�e��\ߪ����o�ud0!�<y��Zs����C'$扽F�VY����O�ǜ`ç��cd�b��6�w$Q hc�M9�����Rz-Pjn���`'3�%�ڪ���w<��}���/���r"s�����{�Hw���=���b�.��`�ږ�s�[��,���p��'I�nҢt�ԦE9���R��OÍ�h�렻�ۀ3�����;�&�0�.Di�x��6<�^��G�z<���R&��Q�*!C|t�`'�m��bP8�o�E9�N�q*�$h0(��vwB��ck�Z_��3H��ӐE��ρɘ^�TzN*�/��5C�^�4hE�K���D�aB�w���k��-�7��8�R��K%��љ�>���U�m`�np���{�j�|戊�p��T���Ҋ�uUm�XwC"c�<o��Y����� ����s��#�wTt��_��Yt���ZtfvH��-m�����%ȳ/�xțw�J�C�,�2Ʋ<�ɓ\$���V߱�KO�p$�Ft�j�B^%�Зϔ�S8��J�ew�C>�$Dl�b{e�NW�m��ݖ���6(�D�PΫ��7	�kγ�K9G�-ȇw؉���)0���*�T���F�O�Kǌ��|���U��B����?����?{���Ӡ���Q]T�]e$z[�����n���-Z����vb�K��P[{j{��!�U rk��U�F$.�߿2���ہ�n{�R�~�$�$�pS_�$L�x*d��n�b��X��;�Xnq�=F<~_�����6�������FS'4��<���Ͷ=f����߮�Y	��Z����U�Z�|�R�o1�?���du�����ji�:u-_+e�k3V�&0���&Z���M��8$=�L�y'Е3���G]ynÜ��T_�T5�r�m>�ҏ�#g���3�W�5�����$��Mā"���1�-�x����k累M�l��������8����@ k��HIJn��xΛU?�����}Z��-؏ȗL�#b�`�=z�W�}����������}�H���FDE��5َ�}�)k���~��ڴt�Y�.}H"��v9A�����q�I��r�"I�N�k��I�����B&�}8]^��0���u�<�7N��Xt8	���-�6/��F��1�3>\�Y�PS�=.�!����4����*��*g\`�� "B�By�f��1)p�·�y�
 o�x8�;�n+Jfw��|�^�T�PyW��Ɣϖ$N�Bt��44��%>D�q�&�hkB�t���vΫr�	˄|�w��N�M����T�=�l�E�-�""���P���tQ����q+�%.b좮����vL��f�U�����<Ni����Ը��D��V�:0|g�$����������:%X;>R=���n�ʸ�� P�����P�Z(�Na���0Ѩo�5��0�ՖV�1��c���:<c���v��@��5�#Y���Lt���`0Q�c�g�"r�Y�kbkj�8�G����'�7��>��g����F�/�4�߻�>Jyj�~�KyQmX�P d��
 �K��uȪ\\B�$u��p|-?��tq_�QA��G��-�٘*��j�X�C)�����zp�F^wY"]l��v;�q�c�)h�������!��"�X��#�k��5v����u=�L���O�~���U8��n�Ԫ�x��v���O�2JьBsp_@�a��"��ƾ@#���t.�Ր���b�Uk���nZ���@Ȓi�T��b�K�|��|����"��l��R$�D�ӕ.}���t�q�� i:P��2��]�}�O�����S���?��9�$i�&��$`��tȅc�#�f�߮9o}�]�|a�~i#�H˓��n���|��%�N�,$q<e�?��{���4ڈ3!���x���"�n`ˤ6X������z
'����p۵m-g����]�V�˫���c���{���FгE�`��-9��Ǎ<Bt�h��Ta{�b��'��옮�WZ�с�ws<<KXA�=�=Brj�O )��^0��\W����!^�!�]Y� �5J����b!���L�rG�Ѿ���-�X)9ƕP%H50(�___��Z���Qv�%d�!��:�m���i���cº�ݒ�>�@������cg�P��l�m���wJ�����d�����A���|'n�g=�ҏh�E_-{*�Ƙl$u�!�lR������'���?X��?C���������û���������)!̵H�1�eɵ;E\?�-|D_H9R6���V%+��鲤��]�+����D����h�?/qVḚ�����ƁD""��&48�_�}��M��ܩ�]F��C�ëd>?ٷ��p��~\q�{cO�U����!��Ɗ���f�֎�аj*R�v�����ɼE�7���;)PM����\����� ���7s�����6,'��ࣘ�/��O������Nv^p#��ǩ�}f��aU��6�uCOc�[9Q�($?�`�KT������y���fk�m�ɝyw���am>>�9	�>�,����ؖ�H��G���,q,��A�V��$���"9,$w�tN��z�ȫ���z����=duv��"�r�y���"L�,!p\g�d]AZ�)�[N����ɓ3�F=��j��U����π�����E/�,ړo��(�w�g��9 ��yZ-j�;O>��osd�܊|!�q�j-0൷�'��'e��z���� z]��Ӛ�\[a#�)r�"���0I[I9��Y���I��~lm����멛w�*�.���
���&X�Z���΅=�5�m!dkӦ�>��~���^uP����
�.�����?<���,8��;tria��5����u�pV�q)u�4L���欖ѥht4�.0���O�Y�Z�J4�5��v���G@��\��w�Q�rm`�K��������Jo]�'|d���T>�u�����ԏ�O߷x������Nmի��x����֛֓TS�ȶ�}���WC%U���^'�k�Ϝ1�`�&R��q��_�TQ�4�R%���}q�+��C'��FML�&���5����2�@4rPq�(���71�;������g���"�%Ve��gv�R���Y卑.A�{ E�NK`+}�`D�lɸiov��f���D��/�E]��,��y�����uѾ��96ad�I5�J6�4��.�ڿOx�X��S���i�'@?�>�Îw�~��������������C�* A2^l�]�a`�Ķ(��z2'�l����Q�9Q�|$���3���!�����P8n{JR�)�yVjPS��!w�+��s�4!�P�\B'鍀?��8�aM�$f\��R���h%	_OC_�n��������#�h֑Y�:��Wd�\}RW"�p�}��a����W�/V���ʇ!WJN�e&V�X�u9����eS��֦?9U���Y���;����I�AAPC鱰�L�0싨�+�ȕ'2up:l�SNʙ7�	b����i��G������ s�Y��O'Bm���3)��meWV�B�IO�N�$�/�/o���RΙtKǙX_�U3Yq�ϻ��9H�~\�k�}��~� ���0��G> ��O��^4&ۢ�Yx����vju�a�"�Q]�F�+�&���/�a0�#@f����srq���d\�����zF�/]����ψ�,m����g�]҈���`�Ⱦ2��F�wG0Cg�Gy�3�N�������jٿ*<L�23cx����/]�úk�;��2����>y�ư�{�I��?b04�e������ܙ��h)m\�@<V>��9��ξ��7�|�GГ���-nW=1˞�:ӛ-���WJ�����{�0t��.��=cl�R���д�$C���fP�H��L6}�p���%�0%�9�-`tȢSI1*��� ��H�G�,�����P��oNi��Ϊ���-���J�ãp�-J�b�H"�is�K�JA�MoR��L��s�|�l���Ni���V]��0����s����r	0���+�������W�y���k_�=�qδ�J��b6���G��!�U���o?|f�r<�$�\�KptHT�֮����1�Q������AkxXE&�U�S���N�D���5� Zr�z��ן+3u�[(ܰ!�����'"��f+}�Z�� <nO�|�%�x���+ˑ��~r�Rr{���/H$�����4��]s�!p���y��V+|�N��]��v�����((�
{�%����n�����H/���;֫1����_ydd@�:����,���e%1Xj�_��KR��9)o�eA���qK��H�� �=�iZ�����;5( �e��;lb�(�����ChA&O{\B,"-�`��4��\ ߠۜ6�$t����_��Q}E5�I�yqQ��.���@
q���F�p;'5��%��]t���}"R!
�Qn/���w��fz���(�k>�?��`r��	H�&��4�/�7ٝ�T���g��%�e��q3���>�c�c�Yn6�������Q���M%p�r���͆��<D3���q���\Ȗ���&�2($5$%����fq�
��ӳ_n�D�L�5�gH� h���L�D=|F��?�n�S��Qo�G��Ь��;��eܞ �K�e���D�H~ǡUSxbAֽ�ac�GU��G߿{��!�TmC�"��C��}�qjP�0�~4�YT�Tq�� ʆ���+o�4���6�Y�]���R��k����Dj-��)s��7�8�
�:�1-g�L]c��)m��ȯ{g�}�	���˱�-Z�ܜ���W[�~�垠b�\9�'f�%ӽwܽ�65=\-^%
o�1k0:��ӳ�:�I���֫��W�٘{pd�]�G�K� <#a �C0K��b�#k+\,Q��K|"�P~���	�t_��е��1J��K"�ij�c��q���ˆ���;��AZ),�M	�0ho쳡c\��k&��^���pi�n�5)�G���q�����~ڴ@Y�)�+9S_�Mf����%+��۫4�)�H���m����,�M.�!��$����h�u���5=��@�����
bԑ����Q��M��2��0K�{&��^��c��h(n,��������)�q4���bG��8K��3*l6 ��T�DE�W)d��.��1M�G-�qI �����t�G6�,�tJ�T�;����"O߾��`�V��˵1Gܺ��GLhG�����=p?W{˓��xOwH kJUUMo
N��F_�_�����8�cfLTa`�``������*?��~�?��������DV1"��0"�{��d�hv�>\�;c}���@����d-o���^?Y������	m��N���d|&����
O{{`7�/M����B��c�M\���({�gf6��� 2~���0���,0���Mx"_�in��w�2H�W?�<�F�]�|��V���1e ���(E}FNߎ-�Q�o|�@�V���u�Y|@�ٛr&~X��k`�(��ph��Z#���[��
g�@�ix���0O��©�I*勋ˣ��?Ui��(؂g=YFW�Ik�fbs���Y�$���k�f���~-v���5dr�$cb�����{[U4ɖ����AH�]�C����4��r�"+?LZ��l�IĨ��9VK#�jm]�/jKw�_/�i�a~��E)Tึ==4j����{�	^�%������2�?����}�^��0Y޶�If/�5�"�;�!U%=`^+��݅��
��cT�)�k��a>�����OMa3���_��/fZE�A$��Xb�����ŗ�����N�ڿL����W;�Y~=���5�f��}ۣ�ªa��?�)�K7ņ�؏���:�D��:n�w��I70��%�Y��7��(��y=�_g�c@4��h�^�X �(���Ǻ�.�1>ŭq�DD;�X"f�n ��Pq���.2}BY?\���1���h������_�PB�F'���^�_�0�Jf��dg"����_�F�1�� s���\f ���Z	���-���olp��F{����9�O��U{(��F,����jz�_�N����;����ܴG�jϜ��Q��'�	�.$�E�܌06�C����J��Owl��2b�E��d��&L,�㝾!	�?/��9M��X��u�Xc�h��SBw��<�`АR#D���P����:'��S�3����1rTֈ=�B�զ�2��C8����0[���ɦ���0^���D2� �תMY��U+:inW����;��"�jmP�~��z�/	xh|�otg�r �xdB��V��7l��(���-uTB �>4ȳ�^�z�Q�`�N"������"��R���3����FK�_5=Q��mWX1HP���c�:.y���J���U� �2IEb�%�D��c�ZxV2�h#������"=��
�V�,��`���'4��^���WS�� iaA�1�_��:���J3X/dJp�ETB��\{<ś�c���>E��:�9"P�1!�WeG�}�����ڃ%Z�!p��hؑ�GB����^�N]TZ�X�����Z׀ �1MH�I,9g�ɦ<,ˇ%��6#Es:.���Ŵki	���O�L��'b.����&!�i�M.bg7!��U��bd�m�ʯ
�ǅ��jrY��dvՇ@Z���\	��%��@��9g�6��ei=eO�X9PL�!�W�W��p������*}��h�Y����o|�t=�V������U�z��Ք_&w)_*�te�f$v�
��ZD=L��a!�ϓ]Wύ�0\_�>������E���;{��p�r`��1|�H�0�Ά�~5\��=T<8#xt�c%U}"Q�&Җ:Ї2�hdo {c��Hޠy��TK>��ac
v���R�#��
��ބ�%���ɨ�=��~4�:�7�@��1�m&�9���y�h�Y�]U5��e������>�Ҿ�۶;��GW����u�a�	v���C9�M[�y�dJ���B\�M"*����J]���8R����Q�����U�$M�5��:F 5��~m�Z�s�	XWz�9�M���˽��eQǪ)��&U4k�tǰ�ʊd��
	e�:-��^�'.��UM�������­���k�.�يde6�H��n5�$17@V>��u|u�'C��ҟ�2���1��nS8%�P:��� �3�M��|(���A�T�`�f��a5cd�����o[�R�˨�a���~�0�x��7��5��HN��G]�3�pA��%�!k��d�����a��NZW��0����=C��I� ��&����e[tmui^݊6^@Mχ�p�����r�Y����]����]��{�Ȃ�8�<(f6�"n�Qs�Kl/�erO3�l�&�X���]e�n�=��<��)������y��{�o�B�h�򣍹�_V=�"lZ&��Z��&$���%��ј3}��>�tP�,מ���k�e�{���A씸_�j!ηy��h鐇�dT ��{���A�>`>Sa#�x�MK!�%����_�C5�ZC����Qi�vd�;7�Q�^�*q�sT�#4�x��euN�����Or��cA��ZX�o�'�π�� ���Ҩ�)�G�IW�����_��z�[ݠ'e�A&K|����fL��`+!\˗햋�{@��t���e�ِT[��R�S����~�O6jwr�0@�|�C֚�p-2��i�}��r&K�v�(����|����e��O��Fi�� �Цt�ВG�@�U][L�Y�햲|�n�'���,�`�j��>�nWL5�������[�C�܌w5I����;q�bN+ͨ��5�"(uv�A����)�i�O����<��z��R���Ї��Z�eS���|�����([�8���Co{$<�}��	[�4�w�CI읁�&�����[��C�P�R|e*�0�xU��*%{4?� �C*|Y!��jX�a��BP���l��EU4B_^bX���cq�@��c�!V���"SO��C!�H�?�I���#�]*�D�]Y�GM&�2��Cc��u�G�A^��R��w��������+��7����U6���S`�<�#�=���m5=ބ�ɾ��4���=�k��?�Aw��,u:lT�m�ZQ����R¯0�83�\�(1��3� ��e�k%&�0��K�*�f )��E�@����ڝN���Aux��$f��=Vq?�D�G+�hL��
�7ٕ�k�YK�`�\:(��qOQ\��Vpߘ'����.N��*@�!~a����U� �Es��)D��~um�\?��jŹ��J�;���{y8���u��͉�̔�o���~�c�)3J�~\��M�:<}�Dg�>�~PVţ��y*�0RRm��S�p���!g
��B�A��A���1z�W��0��ƊL�����Ck��8]���:��i������a�*�4�k���@>_�bA��XF�nt[���L���K���K� � Y�C���mO�ԃ��ͪD{���o�Ճ�/�
E���C
ZTu?ڗ �-�D����#����mщ'
%�{��������W<�b�@�Go�Q�Z{.�̌��N&J'@f﹃h�3�S ���d�*ϭ������A�y2�^Z�V��n9�J��V�����`6�N� ����C�,10���q��'9���/�/R�-���nӅ�����,��&��K�-�>�{�RI��oA�k�A��}��k��Q���������9����d�	��P��Ժ�#�4y~+�4r��8;�<�����ʑn�q��`Z�r����*#%�y����31�FO�����x�2E��Q��	`�f���*��s�x��"�>QX +�i��,�Xn�?�����~l��2�+IG���<�om�ϱ[ɏ$���,,��6����T�ڞ�9a�㩁չo���/I�Ts0�`)��ۦ-�t;�'����y����|�(�����s!�-�$�NT),\�vԪ��[_�0�#b�8��l��FH��1�w�f���,?�P�!g�9��(@ڤ��E��A�[��lr����'�gv�@�^�0� m�+]�,Tq�eC�m%��=҃��dU=�P�j�`�F��*������qj����\�CP��9�>�^H�R}��i�b�?{\�y+�"���1(��j�mJa��O�����ʬ;�þ�d�[�m,��;C,���Y[��68tj㪴a�I� ����jޠ,����\�r���W��3�Y�������zg���n"���3��wsn�r�����%�nG搋�;|���k�T#��,��K!T��������4߻�X%lટWM��##����rLx�{�X�8��VOzM^ɵ[���as���*a
R�������\�-�P��qN�um��3j8K����h�S�Q16���q
�ւ%�]3�������XhR��{Q��C� ��l����3?w�IC,D%�+N)1� �m�c��$�����eN�Q-�Nǈe�9�e���@b�����_	7y?�Kl%ȧi�T������,���cpY<�ϵ�������nn1�L�f3fE��?Ke�ȇ��E�P& U9��UG.�l_�C�D��i��8-�j#���$����C�8�ĸ�M�G>|��ݼ^d�|�ļ�j�� #�u��˅��g�����G���@>�F]7`��V�v�:��΁6z]t�[-5!ɫf嘝^�=k�<��̚�>k)�����f��	�������G˲	��vu�7�[qq�,\���Q�FYdz��xїz/F��#�~ޘ�C�I��+� � �����B�	�J�SVɿR]<�ʣ�7��ڈř�r����*z5Os��>�ǈH���DҼV9No?�`.h�;�[4S�g��%���p�R���.ȷq�6��4`�^���� ��0[i�h��XS�dF����U��-�I�y��x�%vo��`y�����g�A�=�$���wh�RA�I.�1S��]��d|3��E�v���fccb�4�$bj?U	��|�x��U�Z^׻f_���'�X���d
���̠d~�d�fɃ@��+[&�6�dEm\7 =��@�tifO�vŐ��I�q�V�\PC�O�v�����y?{��u��j�B�DG���+[�j�w�Q*g���d���d�
�q9w�Z�Md���um�D��ʳ�ّ���	���uR{M�x�>�`)�hUZ�E��8��^Q�3�Y��o���YF2�М@��xʋ���I}U���@�ҼP�#�PΔEß׃��_i��́�z�(h���^����������$ӳ������c���������N� �P�0͡7b7۰)&�E �V,Qs�.ʭuAQ��������,�A�	��#"�� ��-�ګ�]���Dg��A ��N���%��v�C-"-�R�慨� 1Ծu�\����\�QQ!B��I�QF)5xe��~ΑR��������k��Ţt]W[ܾ"�X���f4�,`��hX���$D8�eWk�Z����o�؅�V������	8\�q��J��c ��*��c�lC��@�^���H�"p磱�a��ˋ	����K��0]�Đ��ˁT;]��i�/��q5�H���t`�z��]��ˌ�-9ȟ�o�6��]�� �WES��e^D�]���3���lG����.:���T-짬�c�.:��w���Dc5�Zh�s���	��{�_?�R${+��(ԓ��B~�*0fl�v���
��ψu\�UT��\��vĞL䄄��o�g�J̶Fd��$u�݇AtD�_}�?ﳦձ�b1��%ީȭ_��l׵3\�2Q�Z_�3�ؐ�ĊXm��I�3]j2rZi>�b��J$�Q��W���;'�K���υ
n�����>Y6�XH ���+�F���Ci���d'�l�'�Y�kqV�eE�����(/�0������!�P�<ݙ�T�����U���#'!B͈����FƊ�����	DC����jknh^�~9Pv ��7婃�-h��*I�݄�@����\/��D_�Ϸ�"�<�x; �0�~Rc���"qZ���d>��@Q�`�a#��^GG�
������� Q�&��ҍVab���� �,�[\����9��*���X���4eD���(�2�wbX��������g�h�:;�e�聧���Z*��+����>��r�I��U{=�T�����~R��Y�W�QɅ��?�X�e�:&ŝ�ܬ�_����ׯ_+0�Kn��,>oG���!�@�7����59'6��6�����&u[%�&)I�;BV��39s�-�̅V-�)֕+ �#��i��P�$�	�rkL^�1
�9z<�iUq�w����RZ��T��]!'��|�Ldt� �կ�>�1��=wV*@1�p�xs��@��R�g�X����H�WE%x��P�ta���O��u�\��
�{�	K�+�$�4���u�[5!�iSG4�{&,��d�v[ �-w��Z����,C���/��V�C�xj�� c�M��r���t����(B٭���(�t����pN��gc7rh���)\�V��"�Z���n��S�����1�l�Ӹ �$^�h���e�ؐy�чb|���M�~`��r3a��5���|'�'�u���H ��`�V�\��r��?a]�P/<��z��
�C9*��x���F� ��C��F�����1y����YGSU��w�C�&���g���E�Lg�>�y�&��!G�C���6-{��*�h�Л��PE�ԀSx�?�kD�Z����
41�7��*}=>�2�.q�E�Q.82{�m'1��n�Z#[HB��t(TT� ���#��mxpg�/�"D"+�������T��B
�N��~Xg}*�Ӣ-��$
1��J"׉���>��C�'��e$FS��zl-�S��=�є;Vx�lK��g�c}�k¡��}>��EU��M����'�2��γ ���%��zNFn{.���)��9f��=�`�̓ܵ*�����7K�2J��lA���8n�.� 0��o�Y$�iOY�؇�=�Oa&@�����C�=i2`H�U�b�h���`w���f�Y�v�h�SǨ���S��6e쟣�`D�hp�z�2v>�*�W>���T5��L̞X�� av�z�ū���?������mSP�V72���Φ�W�5�I��;Y��ߗ�G������:AL嶶N��p�.����� ��r��� �iȍ��	0 ,*�{��(I*�_��e�O�W��m3 �n�f�A[�Q�ap��O��4����1�4�KV;�2��H�%{�w��&1�z<�����`��*tp��/��tT�k�؀O,߲؃r�X�����|$ބ?��uF%t�9K��O�����St�,��K�g�55��;HAS9]���F����mh8�~��u������x�K�z�X�! ��xM�@�_%�=E[	q�Tq��+��ۍ�xZ_�K&Pji��zH��9�x+'����ut�(ׇ�v�f��YM�r�૝fa���d�~
Jd3����pX� ��4K䗿x�n3�r
D��Vt� w������ϼ,KO�u���,�������r���Y�\m�~ͦ����M%���/vjj�qN׫$�y�b_��[�ŽVn�ػ;���_���qU� ���ϲN9��:a���ޘ��g:Ӂ� _�Ͼ�fc�EQ/�'+(ڲ����%EZ�S�#p���&]C�y@�7hu��8KZX��eC-x�;��-�!�	
 ��n\���۱�o)��]�߳�����Y4�T�Y7�'	�Y�&��=�5YM`�H��[���h��2gڭ��%%�A���5���a��WG:�N��1U<!b_����g�j˂�T��ێ!�SdO����ڗX�4��z������hLk~���F�z��02�vR��-c	���l�>TN9��|��"Mj��d������ s�m���*����[�C*�E�RA�:���V+��ޅ�[`A�E�<E��� �R��!�b���Zχ�3�ל��F����0&�}����I��d�7���J���pVtD%���=d'��<��r7�;��](�ia]a/9Y	m�aH���L�'+Y�x��=�qH�P\�DX�����W��b�GvX�`˹<l�Kۤ�� 2s��,�^g�<	8'>���+�ӌ˦�7r(��ХRS�� �@̓a�o0�����ۿaK],V"�At�e�b��^�𰪒,t����~p��?.!	ˬ+����3���j��z�M�����e:�v�.F���Y�"����(���m���Mő�EHY�4P���n����}�Dq#g�`A�q��R`͊�n���0����p�c1��pT�ld�B��7��Znx��'k´������u�/�>m뀩d�_�ϣ����"�"��qVt`��M���.J���x>� �:;Ui��B�V��*3��d]qD�YR8S�ښy�ZZ ����k4�П*%��w��j�Lq����p���o�c7F�F9���	�덀��������vM�L�e˒0!�[F�-+vϹ6�b���'AS�OM(K^��*��^��:�z�����Si��3BE���1���sY��b0s���6�{�*�1����h��X(c�$���)���nn��$E� ��Qb��鳪Ǜ��+�fH�J&�[P�i��9%�m!�X�T�WJe���"����
�8S&�h�6��pQ.X���c����
Ȋ��^5�:���Hk*���!��i���c`��]_����6�� �Ej���r�"���2��v.NHtr����!{�8���tg}C�t�+�?��s����~"�ǫ��,�K��Q�;��Ӈ�^��"?�j���rd����G��sv������0o�#ʠ%߯���r�Ϙ�7�Ӵ���j�NS۴r���&/���K,�n��	�h��%G�%�r4�թa��BS�.��
H�
<��/.�5S�%8��=�3�53䴽]ÍCH���!tEd������F���<f�?���R���"3��[YH��Ȅ1����	q��?�N>�h �%�Y�u�[���,ɭ}��W+@Ъb1�Rw���Y�{J�O�M|��no9���j��~w�[wBmҷF�izU^�σ�f�Go��6��;|��W��A�r2��$
ڴ&>H�O�t�>�]�����a(�|��Ā�%I�^�4\��z��6����X�u�+��R��{��� ���q<�:�p����ğ�ň-g�\�>����S�\���!�Eu�w�@��ڤo��!���M2Y%�=��*�KUP^�m7�m��Ő�Pi��p}�d��2�G�)*<܍U|	?���O����c��7�.��,�H4x]�����}-�]��!�$4Fli��5єh6�os�5��Q���e��2N��5l0�������y�U�X�<�d���;�<.�ǁGIY��:��%Ż/QJ�qD�{k����9��mk��,��	}bF]����43��
�u�G&C�\�.i��ĳ[S~����w\ܔ����z7CPo �4S+������y�U6j��=t���s�&�b$�}�p��'؆c�@�Y-���G�
�_"�5�Gi���==�#��И�*�m��WjR6}��(I��Y"=�*��k����4��?��x� e^��gQ�����(�X��|N�3�Q�A�n ���k����Y���|�K���������J�;tS��?�F�i�K��bU?����Go���[�$���d��|�B�T-|T�p͓�ꅭCbHt�����o��^�Y�c�[m�e�!�ӆ�L^gR���\�J[Δj�����	FB! ����{WU5��]ݎ�=��)zs��z&��Ň�P���kB^}MP������gG�a�$��@�,��R��׃��Fn$`��<cd(�v���	��0��e3�?�P��,�𥌁 &���9�֮Ln㯉����p-�@:� + �j���kH��g�/�fz���(".q'�����B����y����Qw�Xy7��Y��LMRwG��d�^��uh�>�:F��8�����ۋu�y?��[Ϛ�����&�Q�H�(QI���څ�j+1��a��N�$#�����T�6����2̅����Y��v	XD�n��B i)���AG��;�uu�f��1(��~�dl4����Q��-�R�G?����yd����g况� #�>��Y~'N{s�uM3��ay�ȥ.ن)u���e���A^k��=�VS�W��/��Ѵ���>V��YS�g�(��t=��,Lp���@����@d6
AT�%�ի5df�)Q����4�mEÔL9	2�izZ�������UL��ǳ-��D���N��	�ǹ0(@ƪ�3�O�w�t �ZkY0�m�ɫ��a��E�p�d�U0ͣp��o;_h�(KPq������RM�n�z8#�Wd�Ө�s}w��A�iC�}qQ(�z��>>�d@Y���^,�RPk��Xӱz䦐�����-e�ћj��̩�i[F�z vA��b�U�ʤ"���ۏ�a�����eb���!"p`~+]���c���3w�7҃�5��XيKȱ����
:�=��.� �>f�_�7�pU?�}��vM��=�F��-�}�)�я�|����:��A�z}J�7�t`��_���9q�B�åm��_h=�`�0��!��Ш�<��;�p�שAF;��>zd�>�'HO9��Y�4���OV_rE~�t��[~M3��1|c�E
ڮ�B4%C�sQ7���W)����(s��eǩ�:=��>���sg���P��'�a�H��v7y��Z�Ƌ*�B"���Z�v3i+����Vp�D�LV%����3�4&�Ap��:ep]O����t��k��gҕ���)��2QPi��q��G�;p�_vm�g������8��1UM=���C����"�خ�H{�pgWeיv�/Kf��T�^�z*Nn}�����,��CU�)�V����կ�%x���0�N��HIs��9Ⱦ҉�խƗ�@�Y5�c��Hꪚ�
E�� E��Cd��i�pbgR�>b��^(��t*�C7�&�;7��d���j�T2�ź}�NOxv��?:�xk�j%��/VT^ylCd�]:��������
{���l�b"X�w��:�`k����G�ȓf
�e�D���Sa�����`ܻB�flc� ~3��::з�t���`�FH��ާn��X�����-�ǘ����c�Ah��<������?7�U1���^�
���D~<���l�~���1���&m�!����lp��SRcC���y<!�ͪ����f<M�r39�ӡq
A�ִ�M�(y���w��p�\Q;aLb"�oM�_Vaq�]�����(�aiG<�{�dH���6�ZM�{IA���P�hzMST���8��T�s|������b�L�8K4�T�#�	��,!��K�p6K/�N���&҅��X�yA�~|T�nn�y&��g��s�~?k����'R�e��n���kP��6F�m`���������(f����$-����T���Dy%~A��G�8��Kre#����I�vuZR�R��n��v�.�N��?B5�?p��@��?LF?~D|qq��1*O�B8YA&!.�b1�#Ǝ�ε� Q&��r˨��H�,�� ���2_�g	rb)�Hd>�a�7
���E�(]��Θڞ dwjWe��>�n�T�L�@���W���ay� �g�Ǣ�G�LF��z�da�gxA�JD��Rj&#]��A���߮C���o�jt�i
�cxH��I`�U��G�]oh�W���B�	[ݤ,
�u�u��k�k1���1xؕ>� 7�?�0��S�=u0!����l3��q�dq��+8�BR��a(Q�ywU�g�$�z��{��UA8�΄���V?O��.�tR�;TSW����������*!�t�Ê�g�6�>��ơ����J�؎��k;LA�s��۽�vו�z�S��{�3o���?r�nQ��G0��~���M�j`�![��dr����0<���rD�X#ߧ�?�ɇ�g6�\��Q^�� �b�>ٌ�x�C��͑��}<���\��t��@��9f?p�"a~��d(����:��D�f%�[CΞ;��^VP�`����:\�'�-l��K����[����>R��fj?��Ѥ��'ɿ�{4'�k��G�OQZ�zƢ��F��=X��f]�̏+N2v���so�9g����#Au7]�G� ى|N&��6,�[�F�vi��{�@��z���� Δ�عDV~���Պ1�����ĕ(��Ru�D7�YqTCݒ �d("_����.���D��͑�0�Z��k���!�+�T�m��w'��gXV�C�*rFz\����<�d�CH��Ɛ� Y�B�:H ��G�0�V&��OW���c�*z5Ѷ�-��LJ}x0�n�£@)2S�[�pu��/��QZ\#/�<}��
��e�t�[�x7�~����S1�PX�3��9�>�`i\k���I �R�DE�ǀ\���O-m��;4���={���2��6⢱�04�|2����ݕZ�d���_�hWh��Y/	]�E�G� ������Q�nF����L�[T%��P��r�ik9GII	�o���\��cZr:W���
��o�(������������饺���j}�y{�|��&�w
|0.m5���� �Ʋu�Qa�"�#��<� ��^LAX�u�����X^%T���w#��o�Z
���u��A�Fz^������3�D��b��g��0-��H�����k\e��fDq������c��Ney(��D[��HG������g[w�S �晱e��p�gg[���˱�J���+"�6��>��_��@�U�A!���1���3��e�qA�:f�)�C���I�)8��]�iz�KJI����ks
�,��<�F��R����1��T���q�#d�p��w+���1��@��	�^�?�!-}=�l$�@�l�nHb��@M�族(�q�5O$��D �0嚺Z��C�*Y�统��-��.E���0���ca���� љ�p4~���!a�(�v	Lž0����	� �ڷ�B����
�9K���NA��B�[���'��6���R�^���/���o����Y�t���Ǽ�$R�v��o�2OX��g�墎�.�����ra�n_���ڦ��@y�>��y0�	]I3�_�]`�؟[Vb���)@�����9�PФ���^�uݓ���`���D�? ̪�?�/�&n�p]��M��i �)iV�d�GrPƫY8X��5�W�6:A�Nb>H��vц�A ��*����=�9�~ =bǥ��� x��O�g�ڻ4��ܴζLCb���ڸ6?~M@0]����v��&G
3��\E��t��M_��`����ώT�En~z�����b#X)fڬo��Fv<�r��0�!�	�$e��|2���/Ff"�ź)�Yiy�6��ʺ��n�'�c�Ţ����#)\Ύ�+�:u�̛���cؿ/x�UW�����`�I$�47y�s�ޭ�hp�j����9�"�Jc@��+�hd]ހl(��[���7i$N:���u��q�*4�Q7/��49�f滙,����z5�J�t\U��S컌
67��u`��"Z�LG�!ӹ0�A��������Q��#w�!}�'5�5�h���Pz���T�ڥ+߉�N?�%�l�Q4�@:����v��,�-�I��.ܝF��ژD�T���&�1���t�BX�o��G sh)�p:
���c6'o�����瞁Al�Nj �N�����/�7z�n�g��;��:���_WIb\��g��S�w�ee�A�::����S�%�R��Y��n�(��#�[8���X�X<`���vt�l��z;^��hv�.Z'�$#_AbӮ~�W���%U���g���?�_���Z��Չ ��oa�^�����su���],4��Ґ�V�"R�a��`��FU��1�O�D\��an����>s�[�2���.��y+�Ʃ����rT���ϤP��x��Z�1g���1�+QZ���S���S���Gd�:ކ������&����6ݹO�+Z��MB]2��Nɸe�S��2�@+A�e�Ҭ��9d�_�yl�m��@���V����";\X�@ڮ{�s0�(
S�ະ�+���L�fz��v���Z���Ћ��N.��ځb�^��tMx�Y�#�+� ܠb��w!9
����U����?}�em��*��	l(��gğ�=..?���N[��
���n��_��e}����D4V����Y��xW�5j�1���5W��R�cWF5a	�8	���� �i�	K�sU?���*,��Ǘ��W,!5�C�0��j��֓��{=PyM Q;H��c�LPN�
�8.	t_�9!�>�x^N���UQ�r���Fີ��.�w-�/�Y�n���"t%~�"�\�Sz-(G�
���h4���f��w�1�uZh���(����2ױg����O����Q���S��|R��ڳL1������������k������B�bT��]אq���"��"'����ɨ�Z ;w ���� I8��ggGȒi>�U-��÷����J��y?�8�o^�"D��!�yV��؁��7��I���ߊP���TP-�fr�m���X��**�{�;D����_mkh�1B=4��<!C%�����Py�i��Oj=]�O朾�㗞��?[R�AmM6��~��ZW==L/�æZ�N��L�Ԙ��<�7*1��aTt(O��)�H<#�i�U��~?:�^K��Ge�O�雏n�85N��A��JO��X�x�N+�%Ěq�;�M���&��n�ux����[�����ϩ�.4�t� � ��i�AB: �TR�l�eҗ$v���$�7����i�~�Y-zM�~P ��6p�H�̒�D,�U�𒶭^���XЗ��
�.ɻ��ӫr�od9C��k���bV�s������j��(zH���)߶�b��p�,]�l�47HGz�,��R �\��B a��yc��P6R`�ɖ�h�����0����#�
b�\��_a�'�*_��7�H"z���+#,�p.aͪ!�>��"�@ђr>^[Bzಌ\���~>b�՘0C
x��,��tQ35uUjPX�`@'!����gKs����A�(��݇9s��-=�g!�L���+�7��y�tGʴ�����p�&�4u}��##Pɳ*�]���n��Yw�@p����LO������y$�FKh��� ��ȋi� �>2s��r�%�g�0��kiA��'��g/ӵ�9�א<�kV��F�h=�q�3��%K�?��迦��/��G�h2uk�L���T����i��6RM���@/[X�yV���q��@"��=y���KB^����q�a��IЎ"�ՙtu���i�i�,tc	NQ���E���͏H�]MѠ��
r�G�����`D�\<� ��P�v�+M�*M�_X�ʶ�]�Q�a�F�^Cr\�r��.`���5#3�R�F��j�O̙�ޗ�a�¯֚i���r�4���r]u����+�����?UCjaH�����H�?M�0n�$��S~gQjp�kbG����s��E��6	��P睘ۢ*��
�	_'��u�˄�$�^0*T���ն	�^T��P�_��#��w�N��&�-����!�?����D��;��0λ�~���e)F;u�D��OoΙg�q��=��,H��&'�9Ҷ�-�`��wΥ1��Ć������t!��4�%'����=2�MPB$iPJ@�,韙����a�G|�ƌx}9o��d�l>�W���ZA��Q�P3Q|U��	hK�78e�d�	�^�[[B�9�M��ԜX��`��Delr?�E)��f�\��2y�{4K���vy�E>y���h��۫d��5bO��JX4o�U+������-�EYFGv�aܧ�ٯc�r��ga>���U^}���v�#A�vL��V�C�8��$+!\m�G����!��f�
�����*��K}1�Q���,��KB��=%t�7�7�?`���I`U�O8���d R��&�P�29U+N$�ٓj�����m����� Ѓ�85�}+L�xn�X5��@8 �y�l|hAQ���
�tw
�Ս�1�Ƞ�8x�5�� =���l�
��yU|*��Im[�d�_xB{��HQDȩ*>l?U�S��ȟ��P8*T��h�P����`M��?�Rg��ҽ���B�Eu�E���x"UW꿷�8)7K"���p��M��#��[+��w�)����G��ɏ�qwD-�h��(��7}��T��G��nP-9�,t�ݷnk�-&;��~>��VGrI�?�,��`).w�̀B���v�E�AD���Ę�ZZQ��n��Sڲj�@Y��'��)3�l�&�g"��i��n�K��Z|]x��`�D��T��*!��kq�Q����Z;��(�p"�P�[��m��T��iK�PD]O>vU�������e��3���J�M���%H� IX.�!A�Š�����}��7�Q���e���1�4�E�v1`�0(�����苄{����9���A����ನ
w�<��__��g�z�����
.�%Rf����]Y�;v9�d���@�դu0>ڌp�,�s�o`B���[
�A�����d�bk��Wa�uh�I
��<�@��m�s�3|Q�����;�����
�i�ѽ�)�������[v���:����}R��q�f�����~6p��C�{�;� e)m;�j�P�ķ�!g#��X��h������&W �'��|�{ ����WM�":�I��q��P"Y '���&v����s웎4����Ph�۶��ܷ'B� m�杜��=B9Xmu�����?��X������{%� 4���o�$YR��k�d��MzW��t6(N�CR��Ps ���ѷX}$�0#I�
�d�櫛iF�ͽ���h��
<f��9s���y����8�D��~�ِ�vy��<$O�8�v'�1y�c�T5B9$��Ԝ��v��c�w(m�%�c�8�F(�`I�fE�/&�b֍(�!�U1r���F������@�+tL�R}L�i@BߕL>^��6|�W��F��k`<�f!jHy�U�
�s>��*�&�卮�$f�G��{N���˫���1��Ҭ�
ƀ���/�}��զ��&P����a1J8�;�Z�T����K�d���0+�x�u�C�Np�P�.<:N;%lN��2�&��b$��|�����%pH��S�����N>Ma������KQhT�1DY�?+)�1b�F L\[E�aD��O�N<X���l�ilVYb_RD��w#μ���?����%�dB�qg����6�Bd��"��?�š�����(զ����v�xHЅT?����%]��@Z�nc�¡�0�
��/���l��gxv�eNg�W��օ���]�SL<�n�sh���X!i_kS�A'�B������M�j$C����m�iW��f�fЖ�\�g��rG�֜�Ɋ��>Y_�-���T6n�h�{��ё�;�*s�R���,�����4 �:����s��^ӎ  R����G$�/A�}f��reJș�r m�D����H=׭
���!��{t������%�Ws��$�UX���0_*=Dwc��W��������2#	�T�"�����\�w�"�*(ec6���2�_��1����f�9)`=
�E�X�z��=�ȧ��%�z�N��<~�w��äT7R�֙��jE�҇�An����,�r��|7��'+�m�_� ��C��'���50Y���`� ��lk(z:Q�L�������>˚A9x��@%����L�F��a�Q�;^�9mn��|qnI$1Q�:�����'u��7R�z�������
�X ꐠ���?���+$�N�t-2B�3G �x�@���!��t��W:j����z�h�V@��� �:w{mtW��I���uFv��'#92�5�|���`�׺LFJ�gf�.�PvS��L�tȝ��٪U�]������$@F�!-�H���N�՝}��i��e����S-��*��x!h�%tm"K�~��zq!Y���捻r�&�:&暊��s�t���R��R6�d9��y�����x��Ư��;�:��2c?���A�_�r!z˵@�~g�o�{���Zo �|)nXOm�ЉI%_Uj؄�آ̙ړ��݂��x@&�ø�1g���Y"�Z�
I����쫩���G��v^���E�J���R+)�1��LN�`�!"[�c��,~R����J̥������ǥ�$3ݜ�m�[@!/�JFY�G�j���BB�H*�ӯk|�hșA�-*j��Pd{!#�9B����,��r�pr��{&�IB��2��%P�#�8���:�Ԍ1��VbpG�8U��F��9��L��M�ˤ֪`~����?��S dm7����"�٩��o�+#t������?��S�����Y�"01�O�m�S�yH8w���(�>X��٥(�'���d+T���p} ��_��jy���$��4�v���K5.����_Z�M�W#��xz�DҢ#&*﬋�=��$��B@�h�G���E��Q�P{i�N�6`�H�|Ι���D�-�\�����[pk�`�ǘ/�{�S�*b��)�1t4
:�0��Z��īH���;ރl"�@Pk��,;8�V",�ݡ�2|Y]y�a��4	mTd��]�?V��H�(%���F/.}��YiT$"z�@��[�Z�f�UG�*���XzK�e律<�)U��!]^|	�pֶ֡���l�|���z,I����%6�hm��h`�;�y4��VW���;����3��"F�=��S��iʴ�%�.[���pϕzx�(���Dx�
%�q�![R�sK��r��QtR�'�,�(ui�d�N��vbFTt�$�ϛ����=���0kV�j��i�%��E��i��Y��k�C�z�77n}
)EѦ�xVW��D�߱>/9��LZ
`�9k�.��	/y�!�2�ת`���I�H]��U���[�/��/�|ǜ��V�L�
��+A�$�㲗�fԢ�7f�T�"�V��0�i�
H���;�:Z<y#��D����%��"���,��g=f��F@�-��u�Ef��s�{W\xEl�>���2�|�:j`m�I˓�0�z�̃���)�{MU���^� ��J��Tk]�,( dQ�#�M�=�{s�8ڌ19���w�5�vܔ����ĹE��6@_NS�����w��;�r�j�-4�:����ݯݨ@�X]���S�5D��7(;<���.cXK��_�<o�{��؛�+ψ�q[���[Xl�x����W}�h	
��w�99G���B�������&���e��1�����U���t^��;�`�co��h��f+79N^%�;k�!�υr���߮��=�E� �Fف���"� �]�tO���r���Dd�\�@j�)��h��bPX6��\�����~U1T,N�yH۩��2��@���uX$!$��m��$E�U���I;L�몗6�~�*EΛ,A� ���D���nk��t&@��L�b�G���ۍ��7��kҋ�an0�cj��*���C&���y0'�P�2�P]m������Xr��ކ$�_j�1��h���op[i��E�]�E������#v�8�pD$�|�K9gʸ��F��G�Cdy�x}�h��?���<bt/~X�
~����.s��JcJ��,[�������^��wAM�(�[�����Va�
�I�=k��?;�
�o.A��`hkX�jF�E;|��=E��G�,�e���3~n.VIb��:��9��X�K�h﫯c���YGLm9���� ��N~,�΀.�QW]�!�b�^=}�)�N+5R��ި[�����S�"5G�,��B@u�������4O:���͡���m���􃂑[FYx0r����EոU�<۰�Gҝ�1?_��[��d=9��w��_�q�Q�SWH��Lk���=!�����܎x4��	{�r	�	?������B8�μ�
��Y���Mv�d��D�\Ph�����6�P���Dq<���Ο7@�[�-%�	y�9V7w{�W�l���(Q�S�B�O�$ �rɀ���ɂ,�ݠbi��o�B�Egq�����K��Z�)����ņ3KY�m�#�'�@Փ�gFʵ��H��j��}#I�_u ��T�'�@�z��!_"�u�Kn��D��l�5���$��.��z�Q(vѪ��	<��y�Ç>F�:XA{�B��Z��j &sON�6�_���]PSSEx&���)fKz☜��̓0W�CkO �E7܅�b�I�{=I{��YB��r@s3@�0�#������F.��$o&k2FqQ��ZҞ���`RG+�x��t=D�8��v]��U�r����
;$湟��Ԍ<wV�J>��gmsk"�(�%xk�,�k4u?���=]u?�تlƕ-��
�ЅBl]p3�
h=q%wH�j)��^w�kI=%�\���%h��DaW�/P��ޞ^��vE:K��x� g��c��� ��v������ l\��d+M~	۽d�\�R�hȇ;$$�f�̹����ev^�P��&�՞r��䅒|�S�t�Iv�E��Vl�P�W�uF��q���}�D�>@p�\r ppɮ��HAw��@��+���U)����QRL����`��]�}�G1.3e̀�+��:�>�a� ������M|�����1�f�i�5v=-�
覃��l)F��
 ,.:�:Q�O��t�7;(#��H����T�l�戎��{���]��yo���|������f����YR��=�
G�Cz@�����~�T�%F��� `O��3=�z������}�ގ�~�M��bG�pr/�3�0ny\o�5}�v�Ԏ�y��P�)4�׷�	���m�:֮&��%5���D�Y�����l]==�EyJ_��J��P3�f9lF��5�"mZ-t?♆�"\�j޲]�U��%Lȴ8'۱�ބi]zY�����d��#���sʬ���3�����IM�!R �̞�h�y��NR0�i���c��8������*���Ԭ����0u EÊ�'\�lu��p��5,�7ʴ����J%��$4�τ�|(UCr�`� Yw�y�F�ƒsYUL�f�n8P�t�� ��G9 �u�Nc�?|��
�u�O�6L��u F���-�(�K�pI5#�?/0�}NK���~�K���~P7@���v��E.�E׸�����S1�I�;��Z���-���0��}�"�}�`�$���]C��u0o5������C@2���+kS]Hs���X���զ1c��d��ׯ�ޡi��MrN���2�[�G�赬�Xv�y?�`ی���VoAK��<K��������ht�� @�pE���3� i(L��Dk3T��mʧ��7#�)�(&�\������*�j�({�w���Q��;��g�K,l<�W%��u8�i`.�y�D�V���NX���2G}�5�>Z��h����e�wuTZ�pb�
�6��XX���ͳ�L��쬡��^N��2z=���(���q�,�P>�t:,�jU�
)L�BL6l�*��p�f� �b�����U1��\�1�n A��Æ�H�˃|U���r���$&M��╦��*�κ��t�E�C,`�y�G�G���K}fM�{#���ʘ��5!�"�b�7o0��&�Nv���:���uG4tL��d�ً��~nΰ��I:b��:���4	9���D�u�Q��x\�MzN
篸�*ʖi��};ğG!.�@��<T�<햖~V�Rk��C�6k���%t�b�j�Rd�������a3>9JF�	��&%P2�{��HP�W>8s�C'����Ϊz4�fQ���ϋ	M!�xnB����,��1� 
�כ�0��{/O=%�1�QU �a������2k�d�fq�y�Z^K��e��d�0W� � ������C�TZ*[e���9���@�5 �0N4��"c���ؼ3tp(����VQ�,�}Z����t�s�m9��xG������D�L� [�1wip�V3���Ѓ��g1?�OT[��눈=H}����^X�)�}������L>F���I�������J�I;}�B�Ď�,�;�B�=�|�:�	2�H
J}X O�g��n���`��<wTGWX4FRs ;(�t/����a�ޝ6���=�� n[�r�E���L���1����c~EV���e)�4C��pn�᠖!��hu8�>9�Ī��9C/Y��;��2�|[��˽����*, ��?��Z+{M��?԰Mx�]Y�Ǻ|�mNGj]r�a$վ�4��Ri�OSAW��5М�Ϩ��	�U�Vp�-\�k����u^�eؗ4'��Y���&�x��x{n��L�9}��Cu=��2�%�����Y&��!���(_��prf��h�u[t���;R���/��c1st�/��$r9�Ͻ�7W-���{��#��)j�g��մ0��|����"�3�)ԍ��q�Ew�\�{7�B�����I��Kw�0 �����ʰٶu�������J�尥����9�8"��L���GU�@��ϑ����د���j	�Xf)�&}D�r{H" �,$�Z�������p DI�9��[+Y�C�� ��+݌3Բ��i��i&�1i`�-'�*��I��<���������e���c�rd9����7��������(f�q�e�t>�z�mU� �Yl�©�=V�<- 5�ל �\�-�GR����q��bw��|�ξӌJ�a}e�Z�L��%[��.�C�,3K+('���ՙ��#A�Y1��^0'���[�U��!A@�B�QQS��~*�v�4˓!�$�;�5�X#<�GNN�(��Y�D�ʤO墳�,N��� �q���7+�y�Z���^8���7�e�D�Y'��1(���T�S�ڂ�f�n��~fn�v�j��_/߸���#��˲�>�6�O^�TMXG�t��+˫F50�X��B�z�V`�DL�5*��i��{��vf9U˄!��'�R�gX�:�;

5Ot�:��$�?okJy�k4�K&m���D����[��7�gD%Z��s��w��c�������r]002a��b�q��ΰ��F�h�r�Pb��g���}1��[���S�p]Y��  �mͧu�: ��^�����bڋry5;�-��W��7BGמ1�X�.$�_���pǔ$�n\p�Z%�%�Ҡ�z��
9�7��(�}�C���S�KZ�p��0"�����R�PaX-�N�B�d&5!����*
�=�䔼�d���b�J9�H^�#Pu]x���Q�q��5��|�yb��t+���H>��G4�h���c+��ZFP����{p���%�u�ÕlfY��'⦱ӊ��?+r�(I�A���wJvo�i�O2�Ds��s�6B�s�K�k!��oN'wC@Z�@%�=���۹󣾗݌���7I���n_7jfQ��W���ˈԯ$��!'�A!��&���;&�V߅��0C>�t�3|�Y;`�+y�I`�Db��I�.� D�?l)��� ��&��W!ZxT��~^3���7B�\���:�j<,�}K2��O�ո�E:B[��-�C�?p)C���bix,C	/��@j�j�囏�0d�����KR��&6����q\��8�&���\r0�B�ã����}���b�^��ͯrd���	�"kfa��B^s�y��f��z�:?�^ݛj�J�'c�Dg�����K���X�V��I� P:��o`C�R�>��̋�d&f�l����o44���o��GB8}k�b%��P�"��3ӿB���Bп�(�R��~�ގaІ��!{l�-R;~1yz,aB�8�Ūk�� um� 	x�t��d�<����>F�*ɂ1
�%3�C����`$9�5i��L����@`�ȇ減��>S:��#��UE�+8��OfX�0� M3�4Fq/�q��oGi�W.�M=)'���-�4��d�U^$�Z����T��,�&Չ�cl��9nYC��'J�{�4��F!,�?E��@�^L�2�w�&ll��w�K	�i��=�ϼ�+T�m߫��Eov������V�[&��0f�r�����]���K��$�L�v��is.�E 6!�/
���j3\CHև�"��0��Ґn�=Ь*���cwF�GH#�M2�g���♺^3�(�e�qxk�#� t�5K���LD�s1�oa{v�O�K�v�U�"�+K/��nZ� s���^�e��<���یX����<ٚ+sޢ�l�>�G�fF�D�*�|,,-�j��8�Йa��>�U0�S`��G��1/��&��屮�2��#�s�;�=�98�� TZ,_����M	]ǫ�g%�F|>�K�Ƣ�
���M,�����b�}�(�"/��9$D�P�
}�S]����#��ݛ[y)�%�#P������K���B�|�^�F��=�۸4�C ��%9aD:
Hxa>�/�Lvǲ�������M2::!ť���.�p�L�����"�WB�ɘ2����}Y��#z#��r�����G��w���$c%�;sܓ��Oj�-ֳ*���w
sp�D�4>�b?�l�{'�K�Roq� �R!mN���+`�	g�E�B+ş)�>�>S�п�^X>��n�D��;O"p��+	�D�3[ɔ�����͜��\�4�2��v�w��;� YS/D��U־T�o����U�r�/ye�~�?r�ݙkd���z�ӜnZ7�Ç--'(�����-�ui�[?���h�p0�ġu��~
���r��\js�kZ��z)�5�(
e�9]�U~�9��F-y��I�g�)��-}�xgc�s�K��4��k&[�#����w��z&FK+��v%̳w߄p�(e�z̰{�*��u�y8A	F��n��q9��>�)K܂��N�_�|���s�(ߝh��O
�F*7ϖ�j	ŕL�.莩�����d$�n<e�˃f��~u���/���5~2X~
fĠyDi��08JÙ�D[��¹��(3'��������Jy(�.	�%{;�@pM[.�kYQ������{��_lg�q�f�pB���		���E�h!g�Ԗ�.Φ8so�!�4�x�q;;�W(����	[���. '��d+�H!��8 ��7E�vW�'�E��	,:�z<��޺+����<+#VO�3>��#[���D��'�ESg�JL����FKOO2	��aQר^��d�7�;.��䌀I��&"U�V�[��/�؄�FX`���k���T���(:�d�Q�II��_�Н,�>�
Ymnsa�ϫ��Ft�>h�*����0�*6���������b��!V�n1X>>�̉��9w�XC�@�^�A����ETpH�_.�j"���E��*�i��D�gЈ�M�҈a���z ȏ1x���·�S�w*�_�@�d?��_:"eb�4듻�e��<�EE?�������.+��%y�fŜ5F�Y<��0��e{�R�䃒��L[��t��S% �d���$d�8C"��2obb�u[�ҪFW	N�߿��4��m�/��]�҆���0��H���y��b�9�W���)b���e`��@Ln���D�[$��������ҫ�7�7<3�)5A�D��S�3���@�zWW�T����8�/V\��ķ�e����B�v�=�v�[���m��8�BKK�0�+��&P�N���yh�c�o̬[�G�Y�O�Tv����sM12B��cm�qg|�Q�}  "�aYj��a`���v�����P��S3��V?A��E���>��L������m��x�:خ<$��I����͞�D�a�������a��jќ�2h��x�J�{Eea���Qjӌ$�߄	 ��	���Ar���[�EY��1rw�8����`3&�e��i!"d-��L\�{�lO��Kb	)\�(*2����D��^�N���z��[�1$�0x�\5���Q��-N��7_�#���� �đ	jc�`�X�j����{}�\�~d�Ϧ"s���W�T�8'�9�*/��r�
{K���a����-[���F�m�������[U����D1=����o����MWå���3Z��>����@)���O?�[��4:wE+��ɴ��/|B���(hxI9ρY&�k�O⚓װ4}+��q�"�v�C�яZ�/8h'�� 4%��Y��\��q��|�����p���p��W�r��@,`��ڜ������OXvGut�[���fuW�]�K$��K8����u�~!�����|<e�����0�sˢ�΄�\Y`�Ϲ൰��ICKtI�� z���g���V>�O" _�E�/�M7&L\��.�>$��}�Lr3قXft[&�'�팫��p�=c�t��;{:[d�����!M+_2W�fhF]���J�(�>BU���~~)��v�kF���
��P��0����5.K:N�2�G�A��$`V�S8�T��qm�y�Q�/�9����!j���Iβ��A�`(��(�@��4"�☝ɱZ1���ac�B.�"�af�,�Pz�ci���������u'��C���^;��I1��l�g0�#v��&�,gJ��|�0<�L%�G�pv�����|��V�/mz��v�^��_O�5��/�,x�/>���pN|�-EN�&*���W���U��a�;���V��/��Zm����_S��i�%��8�X/B{Am�"�ub6v�*����F�B�5��IЭ��Ȭ��
LTP���%�t�����d3ͣ� ��{����)<���~�է���<�J`�Z� M��!��Q!�e_p\ �h[�B�'��Λ��3�1�tz`��_[y[��Ç=�&�����c�h!��M�l{s]?�Y=^Fx��u�&�BI������a�Ɔ����   ��5DA�2�165�g�+�ppZĆC�������~C::°`�=��$�sXA�czb�w�1�s(�T�m�Ɉ����$��?
��>�7�(���F����܀nf�z6�Y�>�5���Pj �0Mԋ����RI�ɰ���G����U�4B��cg�@r��>�����A�жb���w�O.|�nޔ�Q"���(�VZC����-��8��G�e�j���Y�3sl��b[����52��I {!�#܌���k(ޕQC��ў��k�ۘ
���fhd6gLq�MsЈ���k�{�(���x�Rx\iz}�Q��̊K��F�ǏÑ�T	$�N~��~)M�7�/�kl[�!S�l�����R.�A��,���1&�_��Y��>�ȎM�H��΁�e�L���#-ݜp����1��<!Mԋ{λ�OH6��N�NB~��p�I}T	#��|�A,1��6?��~X#�^Py�kpʵ��H䭧��i+�'i4����
��w�k��
�WbUOu_�q{T�K�'e��ޤ�ęz��6�/��%ƭ�R
w��	(y�]�?.��f��3�l;���n07�~��x��mO��%v`|^�u"zU6��W�G�с���|b�%d���. ����mqnE����7#����ZR�'�ٺ//�p�{�m�{z�� O���WH��-��R�%M�
�'(ZVCL�.���K�� ��v���4r��Br���h̕������0O�}��3`00�I�"A�-z1W��'��Q?{0��E[�����{��� �m�b��q������l�ؚ�`�#8��o�F���C�A@ԙ8P�?_f�Y!�WC����oU�'�����;C�����{lv�7�=k܋��k_p^U�%��rg��C�@�>ͤ5#~P�h
8�P���n'�y �%|`c�4"�*;�j]���lƙ^%`��d'�.�|xntdN�~r{nR��}�׊ ��}�y�æ6�� Z���>�8)�&J����[ܨ+��
���R*œ��XP~ށ�g�	�V���ܓ��0�%û�j�t�j:XG��J�רi,+�������m��63+K̏Pf�*��R.lﶀw+��;�؈���kz>�zվR*K�����6�U�tc��	��$�{?7M���y(�J��Ԭ�����*28�	պ���	������Ds�=��}��Y�
�bs(|҈C�iQ^���������������A�K-�1M5ü�����pl�w~<�1<"��ƚ$tey�c5��W�C�;�qm�=���na����uQ�e��Lɶ�B!�>�2�pT��~R��c�}i�&�x��I\�^�=�+�'p�&e�N"��Y���"E_B���ANG#�v�b4[���Y�>,��`7�����P}�}`j�#K��:�~�o����+%b�y�����ss��OJ�q��خyh���h��F��;��X���r�w��īū��D��bo]�.���p��n���rۮwN�K�bAy9.l����y��;� ��(uQs����1��xx�F�C��7g����R5���*�q	��|�P9�#��n�HıWx�'7��SUc|��wYC�����_��MY�?3�D\��ǒ��S_�)�����$�_�s;�9-0Q]��j~��ˣ��!��W���V�M_����P��E��z�;�-��j`i�w�cF�W��T� �K(�V +��� ��HY%V�u8)���N�ވ��k��s�21�(I�����\���J���@�9�,�ɯY�1�bK6G���G�g�y��=ۙm�f@ ��$�Xrr�[k��)�h%\X'���	JaQ�v�
�?o��e6Y�����u|����ݖPd\p�_�DDr�l��êNHa�Ə0.�=������g[x���aл� <��]CQ;nQ�IH&8���eҬ�J#V&R*�#�lDt4��l2q�+�pu�Q�e���nO1�pr��wqf�k!���_��up�_a�=h^��h��J�ڷXY<Ot�櫳�܍�OU��#��8�m���C���h�x��r5+�`ң��]Fz\>��2#��������+N���[=�X���\�_k�������]^۔р�=��>��\"�-�")Ah>msi��{��#��c������޷_8ʟX��H�I��t`f�F|!��d�}SebV���f��u՚��}|G]���>+���DJ@��DO@�)H����*	���gLI�a��#��
H�z��1�x�jR7lO	�_*�X�d�x��������)������D�[v�mw=�T��O���R�|���=��ڡ�ծ�U3�l����R��*ι�(�h�(���4��E|���[ W[x�f��j��&k1I�B_=�<�]Q�`�3�����f�>3] �����*�[&��V��0m�W�����9*d�h��[�o}6�ċ�h�ګ�ħ�{�OBb�v^�!�Z��x�V��*�]�����������O	�D3k�gb���\�l4�]<^�>FJ��-�����C��	7��X�7?Y�~7Е�X�_�3�rq�#�z�-z��(,A��N�ᠹ�U* �]�`7%	�P'l�` G�hvWh�6�'9�)����u��*۹<C;-�2�*f#��z��9y��Z#;���[�s2����W��~M��do CF��a^oB�#���}������PG}��`�[�B=l$�K��O����N���w��%u��ʤ�gS5��<�(��x�A����U&��u��{�O��W&�����TN�m��!?W��W��q��5M3g:r��?v�_*¥�*��j;��������W*H�Ǽq�����<��hX�1��/��7�����Z�dMX���4c\�~��҅�~^4� !zZ>�'F06�.���}��_,�)�7�gݻ��[��n3�`	��43�*?Ʈ�1&C�~��}ϧG~��$�V�SF���g��L7��H�;�o)�ސ$}�����Į� 7y�Xh��5��	E�RX\�y0Ѷg� ;9$�;A�w��fJCژ]1��������-�\E-܉V��v��%i�}}�\Rc�#Z���(��Ƽ�kt�����g}aΊ%��=���K�Ȏ�ŝ�G��7��.��J��e�W������%>`��SnxfR����9��2�:P/�fܡ����B��v�H�-|b��D���_]���o���CC�(�����VpÞrG�@.���iIO�k9V���M�"������^B�m��58�
���vO�oO�ShFa_iNO�n-�#p���E��^�h���V��ȳ6IW���10�r0{+L����p�1�P�AD]%��s�q�m��=.ўjpյ�p��-�p�����}F��#������@�M�Em����#��C�^�Y���?A�P1<�B��<����Tq[�Yʶzi��SCЇ����z?��5��~[��ӜJ���9��\��� �z*��
S���uL�t�X���lo5�nK��y��Y����fՌ6^S8,I�� ���@3�
\ �;�Z�Hw��0��s7`҆0x�#馑��>p����j햀�ڇ�2�?����@�:��.X��N�������o=W�/)O�����p����r#dn%��#�Zؠ�YW�q4�9�S/�6}�h&F���v �8����A~	� �L��vyZӇԇG�W\�8yn���YI�@�H�33�tǒ��^r�)�Vq�������9�xP����u�(���{��;H~�Q1����h��m��6q�-��i���С먩uq�G��|��m�Y%�4�v�M�[[H�R��B�B�����Sq_r|�-�����\T6�yH�ϝ{,9��nI",��̳�U?���Dp�'���B~rh�tT�F0�&ۖG��/$�o.8H���:��_yu�*^���- �|�=��AH|����a}�Ԙ�.q�ޒp���wQ>�m���`����+�j����Y�l׽�% �k���4�ooi n�60v����z��hlw���Pկ��0��Nk��N���&A�dSk֮at�أ7E��4��qBL���U�h��٠�e��؜��_�v<  ,�B�c⇿����T}��~���hMr�n"���/�s��!��4SX4�i�F��ڰ=qT����\l��)J� �r��ÅV"Y1o2L��G��7�F+O���lö���L�'@3@T��X\��?S�#p: ȡg��t<����&��E�V��bAu��`K��%/��%!���`2�-GJ�_�$��f�<1���bX���O.bMP6i��M9,�cIK�[��g��MX0rm,����@J�N��xjT4��Օp���0c!�ʑ�O�c���J�W�,V���<�C�,w����T�-R'��)N�����\;�f���A��� �>�g#XB��2�	̀�|���]ɆP�G��ʧ`��� ugJ���Nx�w��i͊jO�O�]�ջ�G���9u`	��575�?PK��$͋Ie�
J�Ƽ"�<i^s�k
��K)��(7۔U�N����(��Xu��2"a��v��v��h��Xg)��B��O��;H��x!��q����I�IҹE�
b�p��������,���u�[�ŕX}ic��F�7	�qv��r�E�پ�F~샆�s���q�+��dKH�i͜�U��Ғj�I��yw��� �þ`0+b�p~�[�E����n7%.�T�}��S�b�(WT�7���mF'��#����r���>������@e��~6S4eR��J�n�[G@��>��0�[�{�Et�<$��j�І��=��x\�]*����N�\��9:?�u�B-U���ꜻ�坠ZN�K���yl�c�B�*'�@r=�@�����]�W��O��֒p��Q(˩�	P�Ȼ���ɢ�	kqW&!2{֜2�2�XB�G?OW��/W���'úz��^\U��X(}�$���;�Ǝ�چ%�q1|��wju��3��q��ɍ���Mo�'pAdP�x�ٽ��U;&O`����
�K��&W�-Y5��hE�8{U�E�Eg�Zb5 4[pM.�%���k�궖ln��E�%+��g�|srI�5Jʲ�U�E\!����9�帽���cg�0}���/!�[v�ۻ��@����9d���eҁk��aYڲ&�s����u�V!ng�d(j�Y�(^8�Tp
<8�f�"�60��b,����Q�����w |_ֵ���T�DK8� ��B� �8��f����=e�QtAR�DS�dg�il�*����G7�q�xrN��#�U�h���/epqsm��$��;.7��s�g����F:a/��0ݐB�0�lil��9�����������~��ۖA�U���f��.�?���"ƛ�@|8F��4�w�T�vi�'�&ᯏJ�E��X8$�L�.��yʢX���Mږ���<;z�_O���>⇫7����(��,s])3�I]�L�*1��� �J�~mA�n��w�s� ��P_�"��-��^��ah������~^d(�}yH�����k5����#�?)������=�=Lс�60jx{�o$j��O�c�'�/�$3R%� \���P�ǹ���S1�>�GL�-���ԍ�9�r1�c=��\8���陦`�we}-#��5]��F�T�P�����e�{�~3<Ǌ�d�'�`
��\3�����kp�1a�*fm�ՑC�+ i�3,�����ݡ�n<Rc����4����IR���1W�"=�I;%o"Z�.����Nt��z��6�uJ�]7�ڞ�&Z9��`~f����g�T;e
ō3�1	��x>��R�'=�P�5aR���E�%Ϧ�����XZ��PV���Ҽ�;�ж�]���{�ܼ��RZl�(LBf�}������8�Sn�[{��x��b�n"�!b����Q���JsٯlqQ�i�'X�F[����sv���)v��Q$$~�l�9��8�ڇ�ԇ�B�����p'��ۍ,��+�w!k�;_�!�'���C�"���n��+�,R���V(��ڌ yp�4S1�\�^rBg�����I��Rg�
��Js��h��bT 3�����iE��d���=Ȩ{�fy�X�cq"Ժ�gr]��U97A�"����i�A�^��&w�����#<g'1���i�t���Gs2�CN�mR�:2���&��8dx�5�#��_�<���=��pFN7����$'�6W�m�kM>��R���_<�ӎ�b���_�{��J��z."!�Z�H�[�A�J�x���k������4�.�iNp q�xm�f����l��nd=���,���;YR>g�M<D���C�?�}ℓ=$F��.��:������it�~.ri��L1�$�h�L6r�W�*�O$�Rm����ݡJH,U�a����JPZ���[�6�m��_S�T�M�����'9S�,%*�F�Wrv��L���T���θ;m�@~(T��$�jt�5sֶ�M{�'_�}!��T=��@�?�n0�L3�(Sך+3A�H�6;�I����(�E˝���k�?��50������~ڞG�������a�ţ!�}P�� ���'�F8E'�)GUG�mAS�4�~�������@P*�<�kz�M�j��50_��W�K���_<[noԏ�9�?��ʦk{�R�5�r��j#θ�З���4�d��5�:5S�Ljؕѯ�B���B?׎���`1��s�+�$�0�dq�b�(�ȯCS�����%�n��v�b�0�R���1ڝ�/voP�W�O�i!����Z֚�����v�G���W}��h��B�1q,"�5E�:y&����bZ�a�T4��=���>�@��|�}h�[n9<�]���qa�؉Q)�pI��KS`5����jA��v�+���?�P(�5`@p9L�!\N��8�T��r	:�!Ǚ¬#�r�v{�2����Q@��-�$�����~�7��3��D)��~�^���`�/]D���o�N^���p�rn��]�������_{�5u��ۋ� �(�dq ۝pT�fu���=M�C ķ RW�[���Ii�F_��Q�'4s��Փ�i�~�o:��!���,��G����͛����u2=D�&O��S�I��=Tn^S��������)��*�q�;m�f���M��U�]��$����í��t�M�r%a��"N_>{?kG��)���"�K�"kݵ�IaO�KI]�6����s��1rL��
}�;5�d���.�q�K51͑��(v���5�7W�kkz@s���<y1j��T��O����E2uߒ\�����ͷ�򪉡l��vտ~`S��/,�"~Z[B߸=V����{꛷64nS�;�����n����ba	����aۭ|:����[y�_����05{�_����t;Em���a�\�:�l�7�˽��l��|FD����� "0�z�5-�G����%3���%�~ �B-N�AHva��M܌�MJ����Qۊ	���������Ċ��J���v�n`^���z�F�B�
�%"G�����hI�?r�8HZ��{ |�_R�wY(d�l�b�(��7D�昃¡���Yȷ>����G��B���H�0�����)����#��~iF�فv�R!:�5�DRA�ؘ�𩇄o ���4�85&_�U��n'��@p3 ��ɨ�P@j��\�3��$�})�J����٦�B��X�?���p�����b��;e@�����{���c6-�G@�5?��3���C�δLFh�ML>8�g��ե�#�s��&pgY3�)��� ��b\��n]�~5\=�D���5F"�������E'$�.E���,H�A�=����<
���fK��#�d;����(,D<������m�ꍖ3����'�z��v�\�O15	3W g�	H�&����Xe��M�;Dׅ�si�����`cvV�B����BC��"е�Z���M��?�Tx_u���aF��nП� Jf�d��P�e�X|	mv��.�;�T��`ɩ��;'���	�+\���d��[ݬ1���x�,V4qg��� jB����֬�U:��f�T�A�z��̖_.���_��~
����,0if��\���|�V���Z�֐G��Iǳ~�H�R�1��(�F����l��*�!,��#�3�7ݕ�j�LNs���w��C��;,P�)PR'z:2uzI�C��Eĉ�`���^��U�}|sjg1NHO0�B��8�:h�ƇW��Q��*ڼ�:��H��L�<����B��W0���$qz�؅nyIF�+�o[���j��P؆���蹕X�/ѠJ@�~�Wf`�
W��'�
�H65�	������odW؄�M'��@�yh=��$�宷`�E��@7cj0N�h 63h۰�إaP��Y�� Ԯ�b�Hc; w�Dkj�#�2�Vf!�jg]�S������`E �;��*M�B��\��tއ���zX6Oa���y3���.͑;�}7:��!k�A��u�Uچ�'�w�m`Dk�����o0$�B��e\��Ɋ=��﨧��x
ٽ"���&F^y��e�̺��i%V��+/:SdN
���Ё�,}��?N��@�l\�O���k�!�i�ʜH���c�-U=��b*� ��7)j��|�q-s�;L���iIp\�k �:��W0 ��R��ٽ�����m8%3��uW�L^
�ﴄ 
�5��FL[��rŰL�լ���I,��:�J����"e9s�U1~�" =$f�&gAw��rB)�~�J`��bjIn�b/�E1[L��g�aA²��-�hP�![���Nz�y��@MĳC��1�/��ً�Z�=>�e�B��@��)���y�z��1>������gpcs+����}Bu� ����`��-�!�(��_�ֈ)��x�tF-F4=m�H2P�������$`ȥ���ҫ��?�w%�bػ�ku�엕#�L"�	N�� qdɦD�[e�볞�(�qUr�H�eZ�=���T*m�&�f�v�]Is����5{Ԁ^��2+����8��fZ�%�y����_Aǰ�F��1��ƍ�a�$��Yv1<F�s( �
�i�$�j��0�9�������#
����|k��.�;`�̍r��9k(���]ӟ.�{�@݌�A<��.���*�B�'2´�ʋ�Tā����A!�u?����b��b@9{~�:�c~5���Z)wG�n�*-4���˂�K���-�w hwuO� �� ���O��ԏKV�ޜy����r��Y+N��>�(p*��v	C��e>�:�ڶ?(��������!�(���'�/��5x�ۄ�΁��ϩ��Uw��e�!Ӆ�rI
i]ISn'��]^���(SԠ���ax������D����0�	yG�L��tz��c����y�ۡ��X�|�]�����o�y:%2@` 	j�a�ܻ����h�ɨ>�K\��L�"M�S{��n>N p�u��%��i��d���S�J�Ӧ�)+����ĜW��WS/�wN�hN��RW�t8�*�|ƛи�0J.9�ڨk�	��xQ�ң�YQ�����
N�}��)��Д�/$�&q�gK4�S�hA�����B:+�-X~�P�9_Z�K�?ߟg�.ʹ�8@*=�x�coi��B��K����X?)�h[:�h���^�!�w��as�����5��~4�c8t��EB��E%����
��E����s��Bo]����_���g]:Vb��9�W������W(�`��9��8���l`�{=~�H��[V3��DЫ�"}"�����_��bE�{�s䪺�P�Eؚ�rx%1$�(��W�>����\b�`��VQP�8Q��(Q$�jY�b��Q���/��3��ԐG�Y3��숺��B! �'Q�!�'��/1~�b�L'h���2�p�³D�$�C݈M�`���U��::).�d��K�v��'�'�Ǳ�''fz:��u-lT�p�ڜ�����>�c�O�c��s�{�
��-T]G�A�5��r��x�ۥ�[�H�æVJp���ڟLj�ա��0̓細��P�EWz��,z7J�q�eK<dpTr�7�z��HS�����jG����t����R,�h5�m�#�c�⾕�9�F��I &9a�$���?	�v��b��>��m��rBm�	�q�Q�P@�&I��0V�0�q�j�sv[���ǚ날�8�r�5�����]�~>�`xe�"����!�	;��\pn��{7!8E��/ZgO@��Y6�7^��4�#O ?߇��%����e���Fǘ�����TrrЋ "���̏�BO�U��q�5�af�:�"$�7��������$��إ�X�
�<�y�.��2�����G�@��H&�WΑ�D
ao^H]�'\�p5�'�Q�8'��+��8�[��{Dl��v�����= i^.B9����i}O��El��PmY9=������
�?��LV�B|ʝ�NH�'��X��6tW��;�@��<�6/�nmU���y�v���@u��֧wf�����c�]�� !O��	[���q��,��~������tP��R��o�0t&%Ԑ�Nw�s��F�ϲc<�d*����҃D�%�b��{�w��ae�)̻x���4�"�W�({�Z���b=$�Е^�|r�
�?�Y�5j�(�R�]���	�{. \�B97���
�[��w�$��y�zC���"$y��P�I,���6�iCZ(�(�6�;nx_bÂBT��Ƀ\�%�!@m}�R��n�׫��}�v�L-�z���-��1��MS"��_�נ�bᚺ	��|a���ܴ��P:���F�6��<��x��)�R��h�F{��h�S�S����f����?����_�*��F`��dL�z��Lv��8�Ɔ@�,K ���
��ES:�=z�s�(sP��*���2�ʹ�2���re��yXҟ�0�)�M@"�.��oxԫ"籘�my�z^����:쌍��X���魻�O�uĖv�3��]�f����C������il�2#��2�*�)��+=Yg����vCl��\�Pj!�*�dmY~��y��H��u[�
xp\�Wo����Y�?���j��!�gUYտTx`f�Sa�X��?\L�9�z7(��ߩm����K���i�ă��d4F�f����ҕ��4ݺ��49E�ANw0�~��y7�9��Lx��]VV_���N)f{��+���#x��^k������@[~�� 8P��9w'�X%�P�T�1�1d�+`�vtw2M�5����C6��Y���񑩼r�@Q�P7�M�q$��-�m����bk|����mJQ�aQ}�|s��|���?�OԹ�4L5\T �?^�`�؁11�G�P���e��I��E��o���ːe�(�ı�9\o�L3B�Ue����%��UAowC�$e��za&��|%�K����xڟ��_��ҲVE�Y2j�ө���~��}�S�9	�bG��F����
R�+�yqҸW�-
�Y��sZ:�x���4���.��=r6v�P�]B�_�B~������L��Tt�2��E��}��}M������>�g��X �	WX�-�V�E�g����>�&XֹۗHk��2'�}PU��_������bk��3Fi�6.Y-�؉�I�QW��F��tl�CU�V��V��oZ֒�`��pʪwv�h�Dz
r����4eZ��+��1�H�A7L��i�c��|4�����x:�5j.xJ��N�
��8q�ƍ�F}����, %?�Ѐ���YTH,��:��H�q�#X'�+�C�h�`�66xU���M�2G�&���d���j����.�� �P�k�#TC��Ъ�����%�~F1�	Z���pݷFOS�AFCOZx�F�x���Սnz��-������y^;������s�H���D��{�fV"���H��Yyx�I���b`p�UG1����&1[.B�4"�ʊQ�AX�>j�T7��L�&H"Fٳ#V�١�˪Z��D�)�	&���+d��{�C��_�	�ȵ=js���#�絽�����o��v5`A�<LwhD��t4h�v����K���<��lW�iW��-`���wm��qRfλo��]D9 �?������)�{6/z�^���f�Ŝv6`-�KW�+>�H@�D�ڣ��׵wzy8c1+B0�R�QZ����s��1�ܓ�m���U������d\����T��� ;�̦1�0��4�T'���=��A�pN��#&��(U��,�w�u�r�ީ��ܾB���*�e7�/��$�8�.zލ�H����=I���m�Y.�]�:)43�U��nBz����N��r�}�i��D�g������u���W۶��.t���솴�W�4/��\��pI���2AbX6��q�-4경-���H�h�:����╃�C��]B%cO���%P86+���E_<@;�xR�q��Ι.��f��7+�������<u<kG��� N��@�'�i�]��n��#�Ɉ����T��)���g;!�d�zh��D���0�b��A���u�l`�X��wW7���h�=�
����#-����{!����q��߶h(�tQ'��!�VqE Pk26뷙�-v����鈉i#���&�uX���� ]	��p"��nؽ
4�+��|i�xI`!ߥ
�S5ǝNHIQ�a���F*�n.�o��y���� P�z�&����}��=O^�H� $q00+�0sҍ�u��I� �(��8.0(���zƫP~qr`=Nr�~��7��:J	����d�=�|i�/12�7������������nT�,u�b$������?��ᤎ%l������;��n����(���V��\��X˘QVT{	z!	�Pn���\��]�ҷ�I��uh�x1A'V���Uew�2$iS�NYE{������?�,~�/I(4��T�M�\Gn����
��g<��[)u�8=h����b]4����\���n'�4?�"+���~HN�z8Yu���Ü�@���Y�R�L���-<KP��0e3i��iJ|J%})6Z���;�[S��[t��'V�]���%{��_a�(7SY4*�.�a����lrL2���L��Z�e1�&�"���F�K۪��
�#��T�({*%�P�&�\�Q~�|�U��I�[E�C�%ڨk#�t�Y�K$"��G��n��($�Z�q��s�X&ֻ`��0c�TV�l?�;֚����%G�S����Y�CA���we%K;4�FP�k��<4�.٭�V?�͊���a�h*�<��������Ƈ��1���B7?j�J-�Vtɚ�T&Kg���w��]{��݃�3�����-�=�.ұ2)1UmX�k���)�)�C2�)(20x�_�)$3�T�lFK�a;0L�ݔ����2��P��*PN�%�ڔ�zSv�����U}��X_�����r\���Z(�|)U*��v*u��{�Cz�U3p;z�*hZ���s�Dr�/��l�$�(�qB�T�$�3�8'�݁^Ϊ�!��ה�W�����f��>��.�6�}$�
��v��x�7�Wr�����d�����b��6��H}1�͸��|
b�_)���O� %��;%Nl���[�C>8$�����Az�ϒ!��6w����R�&��EҎ��M�����*)i6I2��!6`&&��4�C��wwZ���+� W�R@�Y�S9���8��3锚Y�q�3�R�~�J��8-��Z�ִ�(��!�%Ԓ�#`�ڵ{Ym�>��9)�j#�������y����N/ ����A���`(�(~3q<$�C�r���u`]�{�/Z�	4	,��r12��n��vM�6���i��~�lOZ	 Kn��������T6�e ��G���������S<t�s���
U������{w:P̥��D�-=&`�B"=F�}Z��	�Ws������qb�+��5d�A7�֪H �&��Ǐ��:��U�'y5���4k�n���B��t�Un��R �a9j�F��c��ꄣ�V�'�oʬs����t� ����m�#RX,�S��VR�hRE#�����hg�l	��+�r嬰�>�q���
}����>����by�/ߡ�ߥQ��$	���]8L���eg�q�� <Xf�2̙dl�N5X�l�d0BD}V,���9�K:K1��|U������3��Yg�Z�C%[o��2<����vD�yAV�!�_!�xzi."�F�&���v��^��v�n!�J
܇�N�kH�MF*��6Ü����H@q��޷��5
�Ǜ���
����,)���;��k1�I�P�d�n
�]
����)e�<�t¸���$`(h7��bA��s�=�2f��/H�� X������t�r�*HȢ���I��?[|�p��w4�+�]ױN����A�F���8��m䉬�H/ �Ӽ�&�ڀJH6v*F���u$����;���n��f��.�e$&v��^�e��ХZ��x|�ҢL�w�j�+�.��1�C�U��>/c��&��m�����Si�%��Q�|A���[=g.�w����Fsl�څjf{z��D�]����r&}޾ClPx\�>u%ŏP�U�m���Q�x��0zh �P�zE&��>lG�d���~~���ȴ^���|�C��σ����u�RHk �x+HՠN-\���v ��MG������,vk?�1jF�P��c�����iNVG�� � ��dҞ���]�;��vZ�\&O�b���39A��C.�ʅR���%� I���bIs��,\�o�g�"gF���g����¥�=�A��(,�Ya_�����\D��3��fL�(�y�̛W ?I�aKk�˨��fvŉa��)�1�[��{���sA���o ]�~�5P_Sߺv������e|�{�S`���]L'+��Eu��G��$�
f+W�2�2Iʴ�M�py���2����v7l��EZ�d	II�r#�k̙	�,t\�7�ߙS ��/N	bt�T@�A��9���'jsz�^���pv��!g�u8�[��c�F����HV��$��6�Sn&I���������/A���,9e���	��S�?[�t%}�!Tt�� ��x���q?O�([�7; ����6�,�VΉC�+��ˇN	�4��Qxg"m���[���p�q#h*���v��nw&�)D6�(�Pàg��^7�B*<0�lʃiv�G?�lz�d��q	�G�Л���N���iT`hT�d椽'oN�8��r�� _��RLX�N`񵠋 ,�j2�=xY����;�ن�(60U�%��S�*5����2��|{B������u$��̪F�qj��T�~�#O�	�Hšq$�)gXG�۪`�7�P�r(R�6��N�5�U�~TO���L�JmIwZ�^t�i�O���1l�������w����»rg��m+�)�D!@��5�����sE����|_�Ʈ�(�����[c4�1��6L�[%�1��Tr��6��[�M'W�$��c���!��Ex���Zcj��F�#4��C�	����X�X�<�zs�SWT��>M.T9�~M��`~���5}�y4+	���2�Y3q3v�����ax��À�z�s@���n@�QW(�x]LٵDW �k�p$`l��x�hs3x�:\��ެ��‖�K��'���B<�SD��嗃F�������Ŷ�L����y�^=�J/t�̵�T��������'���u�Ȫ�����}���=�ʋ�&{}�dj�(q�Җ!��q輘������/h���^���yQD��m^�j��A��+���vkQ)dN-�xAA�t���/�C�|!<�2�1c�����*��6L��DB2w��MT�Y��i�����PX�4$�����od�*C3Z���~�)GY#��2�bԡ�y'8��
�zfh��tXI��P����~F;]B� ㆇ@q�E�pT��i�f�Ҙ
� �q���֢�� ���zV��!?J���?ƶ]��� KD��
	Z|g��͆� Q#��F0Ne�B I]�j��	賅�pu��$h�cDf�H��'��!�͘��i���-����:�З�K�����Ư�ԏ��$-Ч%"�yo�F詞��l�l��j�.����o����%�g����Ł�z_��W���^,K�"�y���Y[�	&b��S�@����<tnN�X��1b �s�r���$�X����>݂s�@U�o�{�/���;����� ���b�@8��;��.���S"~�/����/���W�][=�]_��/cM��8N
�e�Xr�Ƀ�Y�Fjcl7걢P�TYe��{ۆz_��U*�����l�St� j����b��Yd�q.�9`��VN��
��ff�q}*���V����V��B"0������8�]値�M��8e��(�1BH�����8<������)��8�7Շ|E�����5��{A��A�_$�yp{H����xE���1���ݺ}�V>8�6��p�˳Ђ�H�*��w��x�@%��N��I4��_!	�x[з�"�*HM�O?�y���� ��)i�Ϝ����s���Ix*v��g�d��]���\`�I���4�ok,v>���>8s�;p�@��.�b�]����,
�G�"E���Z�������@�ɼ܅,7���f�m뼟�^��[4[)\�R�j�H��R�d��Eɑۘ�(YS�ɵ.�bp�����W_{�\Z�$�+�A:e�E2N�1	՞�#�V����-@D�,j����lA}�0_=<w����w[�r=�O`��>l�GtMR,�I�rP3��TJ8�k�2^��}�gE��j�����[���h����*��SPl�_�N�[/?F�y���񸰂m fCM�	�h�T%]-t�+p�����|����%t` �Y�(�\�P������� �w��e��&!u��Ȼ|��Tn8����.��75>�Ff4�Ԝ�q���w���S}���\���d���^
��:�a���X�Aã�x����?6Հg�'���T��%����<���S,r�nH��U���GZb�HZU�a&M3�>�U�2��m}�%Q�*���x�{�J��M�dFnR
��lDn$�a�G�?7�\��4���}�<D��I�OM� -}��4z�xe{E�&�ˇ�	\�Ϝ$<��I�9��'��jG�g�Ǩ�����'9<��q��"%��@	�"����m����U��hH6�j��+c�ْ�K���`*@ۓf��E�9c����J�s��2oB�i��Ya3%i�&�7z&x\M:���6oR���6"�"�B]�I9�kkkt���Sӛ�U�ٔ���$�c���W��PFk����O�����	��ҿfߙ�'�l�d%�a@F1�D�s�4�}�<+�-p�����a�U1��o�M������1^��h�A!�����@�@������ �EDzöUf�`9�(��Rż�訯
���B���>B��dJb�<�m���3Ϋ��Y�������g°٥3��R,��30�E��u�+�O���S�>�F4�G�$l7���1�d��$hKD�Im�ѩ	�u0���.�[=B��|^�Twzp�� ���GXa�HE-/C!��+P��sb�Y~��#��J�EK��ڶ�p�F-��{����Il�ε(m�꫟O��6��kEKT�_X��N�TV���l��e�0`�g��ӡ�st}�{<�l*��Y�?��{�jߎO�=$�&�-�%�f�b���{P ��i/��%/�K���Y��k���
Θn��v`�[��ŀK�﯐�O��a1��0P�>�r�c����ں�:�}��̰͚�bF4�k�=��J#�Q��5��L�%wB-�<͉���+C:`����D��INH����^�.�m��+([(�q�RL�a��=ʘ��W�O
r��JN����"�j�] Xպ<v2��Oq��X�NX%)-�&�ϧ��D�X���������4U�R�!�Շ L��8N)�O��#?�A9�Z�Qc�}��uh�|)����M�����f�u"�>�'}w_� ה���+�U��|���cn�Rp�������%꧈����iI�>s�ImOF3Ŏ��iVaa�|ӛ����q8��J/�L��/dK�2H�eS�P	��Rry�HlF�>��?֊(a�ʉ�\�8�;ê���#����Qw���o��%��^�x�����f�"�qdl�ſn�������	_4��Wc:��F�G��m� hH���/,ً�;�J_E�Y���u�0���@'[\U��+�2x�e*�W��y-�>���_ؗh��a�r�{�Q�ʄ�NN��F� xW5�'���
u4���$�]L8*R������|�7�h�����G.qj�I9��G|��wl�K�Tve�` �iO��𓕰��'��4��N����Ĉgbs��#�%c8�G���;q5�4��g�.I���fW����<��	��$�N^Q�%`XA�!�����v���&���!��sQ�~^k�J��� �2���w�.��|�՞u����0��5�!��Cjʖ>����	6׳km
�����m�#�M�=@L+0]�$N����T�v�3��;�PӪŻ�@��¶d�ݗ�&BW���x��[��cik��O!jb�������zj45`>[ė�W�c�}K[)R���n0�%��db���,�]�?���W{��\�
�CAR���D���r�����o$�����t�!��Y}��{���`��8��d�z>�;�,ZkG��/Kp�7��IC��u�rI���B�ՠ���a�8���Y�k�3�L�}��<V��'Oe=f���"n��Օ�����y��Όu蛮(+���2��7��Md�YM��lse�`�y��O:iz���S��]ݍ'��S�zq�6V�� :��������p�Y�Z��݄��_.�O�[�۲�U����ƺf�_ lH�0 )Tm��l`�;�w���D��` )S��������.Z�d�j�h�F��(���&`�8Y���E&��Er��KF��_sߝ�Av�#������l=�A�P��yY �j�~�%��P ��~���h,����mu��ƍٜFR�Z�ɫ>l�(��A�����*?Ӑ,������5�f(�3�k#i] �:P\�K�M�INﰴ�t4nV��ɏzZF���
�>~~���<1�V��k#+�C�	c�R02�8�cf��Ȏ��e���V$Y�w ����~"�*����d9q���S�omj��3��h���T8��9�1((�F�ۛ�. �P��C�%N���??���{ X���ͻp�8qַ5�4:K�6��c(��M32y� 6��T� "t�����C��'�q�9<��$U���>{���j���"�`�.���=��I��[�N�SG�b\>��-�nv[����/�]�0�{E���tn��15.|NC2�n���<�y��ږn�#X����
ᮖ+jh^�	M�	D{��$�3\�G�� }$ge�$���M�x\�y�*��vAo����R_����bä��V}Al��T��� )t-��ֹ*+tz�w������X��D��}5x f`C������(�y\�����"�E$;li��
,~.�Q��M��~�tP=n�WdK��`_5�g)5G5��B��G�˱��t���Jނ�ÇAj�@���]/�$>A��N��"�a��f��ăs|�3\�P�����?{st��#|p8��~f�S5:�
�W�A��y@#�D�s�h�.Pf��e2F�棵���I34�NW/BO&��ˡ| ��KN;���Ƕ�(6��r9��G�j�{3��ݛ?���~����zf_RDD��!C��-P���;G�S_N��5���i��X[�خ7fE����P��A�q�vG�mO����ja�g����eWH�pA�U vhH�#N���S�28CQ�`�8�t�z��\�/�W.S���,�i� Y���;�����b�q��ꡐ#KvzGNk����!E!'����SU�4��vǁ#�ɚk��UD|^�XU-����o�5M��0)"���^.�M�$�����Q%k�u��;YF��Sr��[S-#>Kvxi�}����E�=�t���l.<�PWko����l�aT����v���k~x���'�v��)�%N�!���<��.���2C��k��us�%"4���wzS5]Qi_]ƒ��HT�F5m�).���+�����g!���R�Us�n��=����+�P��K�}�����~n e&��P����`��])����uT'��)�����j��D���PV�b���8���\��.tH�dT�!�|s���Ee����'��c����8�K�(��}̭�w�W�!˗8̇\�
�r��UF��Fd�yVl�_~�ǌP���pՁ�@�p�1mnI��lQGnE�z>}ǍE*Q3�Ƿx�KY����ʡ��=|W-nVyU�w���W������)Fo=V������zR����l�'Ha��%������k��cΨ���9se�b�eߊ��u��/��)�Α��v�,�����k�~՞��z��h+�G�m|�4�OR9;�Y����R�����V/ �P]�֜�O{7e-�$�pe���-�ƥWX��C��ܹ�yO��_4P!�Z�AN����$�@P�R����As���bCc���zZ T9�̦�'v���I���y�m��Y�i"H9N	��ہ��3��á��9�b5�\�&h!�M�O�6M>��/��B{�����6'_����m��A�H�����t���)�l�:6/��ve�e������ܟ��o�v�t�C�H1h��`�����2�1k���ǽ�4Ϛ���R�kB=~I���݇r���f�L��+O��zm��4j��=����vq���&�]@X��5Ԥ-s�:CRF��	?ad����-��-�qj�9R��.�l��ݶ�+ka6��͌<���]K��O����B镼�}���KQ�Ϊ:4�-�1�t��AܼUu �s�$���'y��r}$^_�U�� 5s�Zv�$	�"dǛ4��;6�Ph]�N쨤D�ݳ����y0�ޗ�ń���p4Gr���Y������Z��\ݳt:L����	a��ܕ%�_}w'�(-I(�y㒰
,��k�6�x�f��ն������?80K�s�6��'�s0���>��Yg@����󔷣��#zD篹�e ��#qT���'�`��_�S�Gxi]�v!��smף
�aq��m�s�vzE�F�0;��UPX������j��d���<���f�4pjM�D`/ť:��<�c���h��`u�0��η����w�@�r<�����n�O&ɽ�}<M]Cّ�2tQ-��qX5ga3�m�N�9ξ��7G7+'>�i�M�(<݋�/鿼mE�O�Q�u�U�i������NB�5�w"a�\ |wh˥�I��XW0�em`�Aq'�8ڣla1���`
YP�!�0�.Ӫ�+�T�_7�ʁ�Z����X��}�~�^���R��a)������"���s���̝�����נ,�ĉBv�n�-)��G��fm �m�pP��[.$���ڱS�3��ڱr`����lE�b���oK�� X����5xC�вEҋ!�Ό([��r�a=��[�y����"С�˟�$خ��z`����5H3Ƒ��/I�h�JA*�2�%�u��n�wZ_���%d�*�`��(J��E.D)0�����n]o���n��w��	+�c��E���U�1L}����.�Xq���)W�Z�R&c�M��.rJ�c����FAY�o�-�&�7�9S����R&��/�"�I�Yz�*[�F&��PHgZv̴�@M�=��a�)��E�j0'y�nI�@�!�`�X��,�w�f�B�6wӃ�H��e���g�Azp���	B��ƴ'[���^���l�b=�P��i6X���9����W�ɼ�6���U��}�Q-�IZ�Y�i�Z�����5���uƜ~=-��r���"r��Ew��-�ru�����A<�ٮͩ?l�e|-}������^^���4ܔ��Q;�H�����+{��rb_�4����~xM:(��x6�	�;D2B.+(������X��KfܶtN]k��M��a�]`ٟ̗�^�+����AM�c��H�x⇭oQt�>P�{�Q �02<�QE�Ky5@�q����tQZ��9v�6%���ɴ^��o-ݏ�W�U9�SR�J��ʁ���қ�aN�:���v@�u$��|��C4�����sW�W1��'�:�$#��*/,
�[U�Mb��:��M[1z��5��K ��\1��c�����s���W�7g�~{#�sf9J�F��Xś/MٲV</�u�讵�{�	uv����~�B	خ�}��Ǔ��"�ߴg� I�����m1ӥO�9��Od�0���j��r뺃��d����� �vǎG���J���Mp���;�?�>¦�����4�ڿOgd�h�lCܽ�84O���y����k���Ė�5����XDxLO���U\�)|�_@#��?��pO4`�> ���͔a
���+�;9����sg��p�g n\�jn6�������]c�x��n�b�����7>�rue�E|F�t����6��݆��	z1n�}F�S�7)X�LU͢L���,�'�Xh�r��=MZR-!���EC�Ԏ)�ŭ2��� z�)C��tYj�X�N�	�xk$���Z���i"�6}{2�*��2�&W��6G�h8m�u�9��8�F�zB��n����5,pu���ƻ(�5����^A�G��=�Ø-���ٮ���֞�=�z�.5��#�+-�C�Q���>��!���C6�g�|]��V
N�-TY���8cur�J�&�QS~����OZ<^����i��\8,�j�����\�Q$���#�w���C�(�3͐eJ�\�ѹ�&��$�4�,�n~�����\@meL+=L���1��-=���&[�4[�"�`MP���%��ɚ<�p��E��%,F�\>��}"��}-�3����;�N��^����tǙ���5�m��i=��C�����H3��ԅ�F��#V	������z�O$
�AG�a�e�AJ2��ۊ��� Y��F���@86$���@�E7��ŋȄ �3�QvK+�i�>��ԑ�g�5�.3fo�����ǆ��Ct�����9>��bqP�G1xm2���zY�R��l^�[�@�����E6�Q�;-��9aÍD�:S�&���Tq�V8\vu���ːB�T��W�p�'U1(GՓ`��P<5A��rp�eg�ğ��Q'��%�m�TR��r�!*C;��U!X��k����c�O�MW�/�rR��zn;�E�G~f����p�~�]��j�8�E��j�xB��9l̩�6P~�z-�N����\;�n�@s��T�@����8�d�.���B���%����e�4a�V��q>_q|"�`�/W�voz9���or��� ��c&�5�8j��Pө=�1@
x���RB��;M���~C��1m�v�E�S�D�c7�������f��X��Q�m�[m�;�w��ߌ�M�B2v���&�RM��N�1�y��Xr9.P׎Y*v�J܇�T����Y��Y��������+])�ذ�˾6h��=Z�`"[ĄY�8_��W��<6X�n�5~h�5IA}�:J
�M�xC�
|��$)]��?6t������1�ѧ��07�y�$�m�ޘ֛��& +���Lx���-eXcUC���0.Bh�B&H�x,�Q�QGY1O\�+=���
#�����$5����*�a/t��=&�~^�R�}Y	y0;6��Eѥ7P"E+"J��o!�#O'
����K�߰ގW�!٩
9�풬��HN�Zw��2���L�w+��bj���E�=_$��TD�l��� �ͳ/W>�2�<[V7�l�8*N��X0�bzKB=o�֋K����]�"C�c(�2���(=��M�)��ZeƏ��dt#z��a	�/�T��!
��#J7|v��K3Q�qO�8S*���OX�X��]�����T�"���=ȉ��og�������I��Ę�k�UweO���[�2X��x7D���2IԐ\H��5�f4O��RX��T��tE�.2����X�S�.�����_/5��me�oiKyXkj�,�N�M$�~�C��V��#��So^2�ǆ�q�HByb���O
�����𱕉�R��<P��5�� GLs���1��6������񖔇����N��؍��\{Z�LS���Ӈm;�)����ɹ���*F��F�?��O)~�i�Mk ��PW�'�DQ��C�����W3����ec
�L!$������ɥ�A,TC�� \�H�ɵ[B��ې�T�WT�.`���)��?�9`�
���h�eW_e���Yl=�<�y��g�t�&��Ak�~F�[����w�D���*���&��j�#s�ҭ���xanJBn��7�ް�Cu�Rl�6����#(�5�H��$��j�毪�8� 5����1�#y"�m�x���̱��w9��A�PV�<\9B�*�����&o�����L�gHAɂmz4���`>�S���·�_@��d������|��D�4�M�2�D|���p&eS��.�EX?�����A��4��A����v���"Evӄ�Py�S���0��30�W"1_�ez�r�p 8����B<���M`ع�U�r�킩Y�4�68n�ڻ�Ty�/Y����k�c�1��A�I�u2)�O��bρ5a$��h�3_X<�3N��d��ʑ�5�j;A��H��ڗ���%�Q-�\������+����E(����|}l{m���3�o���؇�)��C���r��j2��y�P���5�O>R���to/]0����ҡ�i��-R{6�p��xj��%km�^�~O�.�L�G����ϯl��/���( <��~.��fc�"�{�T��"�˗I��;�9�!�r�:�a�} �-�Fk�G�x}e%�I�!a��\��&b���7��U>�K���_?�WNl�]����aJ8S8u��g ���$�����;�(&�l�>�[��tp�Q;�3��=�J�c(�ƌ@jP����Z�{�VH�2����P]����1nԠ�����l��9j��=�#.ke)���@����l���y�g�I����u/I��獏#���xL"A(ј�U=/#M�r���5I��!@F�]z1Θ������\��*�%C� �6�8~V^�/`}T��8Q=%QS����|�������l�!ԓ<T�G�M���We�S�VƟ���|_����g$	���s?k���Q3H\��ֱy�v32�3.,Y�qg�PB~��n��HFA���|�'��7���ϛXr��7�&��M31J��G�oWڄת�	q'5�mL���5�7Ei�4e�DpK��ش�g�/81���F]_�J��[���F�ڧ�p���hl�.v�>f�*r�����M���X��Z:ҙ7H�0e"Hi�P܍).~�7V�	z�_�fby��T�1��>q�b���u�o�{�М\��dZQz{�������z�ZeX py(�E!���w�E	�k��]��/��#"��J�'���� �{����
'W�7��{q�u�F/8�$a�r-�3�@���8ʰ^Y��t'r	¯s'�/7k̵Iɗ|���n1�Liċ��d9;�X��M�V<K�A\j�}�8�&��qӧ�şl�<�	!	�بl�^0�1+JMP���<f>j���"�r�W��o�P��z��B���^*�bk�U�#om�� a�0C �r��M@, � �|N�����'����UO]6h��WÐ�����E((�I�tf@nWtۚ��d$���t6�kH�E#k�}�7�+h���27�oS�e}�;�'4����OK�;��y���Ha˻�fH�n�7�0�֞��~�Zj���Vq!Ϡ7l�Q��z�p`��Ɂ��V��[���7E��j�um^K�Ir;��l�H��E(D���݋8���,�w��'���	1�y�@C�wG�4>����-�!%�$m��hׂ6tp����%�^�5��~�G��e��;��_o_�(ßS!ד�����4|C��!�d���:-�&�&('��P�� �+�;\]S 5��wi�ɷ���x�4�E��'�J���jHe�\'��a�O�0d�c���bɔ�.m'y�^��X�a�����!�����r5sZ5v���ۍ�ӝ��$ߺWE�z��y�������7	?��K9������q��P9uۅ��0i��S��-Xt{=����.#�SQ����`z���|!���hI�b��Z8�G3�W�7�fY�o�%�4���!��@��Z%0.${am�_��e�+�9���*sF�ǻ�w�0���g(_�70�F���S�o{P>��M�K��x+m�߬c�1#�1��l4�:[�j��m%�l��؊�ub��7�B3u����ؘp��kQ���6���A��m�	 �����b�:G�/�O7L�PZ���3 4љ�#�^L�J=Q[�y�Cq��@딄�+�c���6����[�.�`��РZMY��+%SRUl��_	���������zJ<u㽩��^�a"�vN0���9�e����O�#T�`��f?�z �V�
�mP,T���	2*rDj� �.�8Z�sH�5D���	����<6�=u�c��\	T�9�f��
�Jt�T8�c�k輯�Q(Q.m�[m�[rnO�-v��Ś�Zl���_2��!�\��xMR殃}�o.K�އC��˒V~��XU�'Y��xE�^m('E��W�}F;L�P���7+�"��q$��.kٯ�S����ywS��[�?W�f��17�p�u�F:b��j^P5
!�'Ͷܽ��t�e���K���{�(Ku�ju#�7R����{���k�'��L�R֢<c��m=�5���n��yA��usHA��(�3�l�f#���X���=��b�j�4��|�@Y�y6�}�7�:�{ش�p& �!`����f�L����[(޼���[�(a+0�Fi�� �g�Q��á�󘪳�,m���f�	|�O��W�=pŵ�*�����$�}���*�����^i����lC��K�;�8l��N���G�������o��wGQ#��[���V����؞�v������� �[��SD�7�W�?,?�4nE�(ĪlA�Ε:%1mSA�(�Pl��$.1>a��z�ư�o�p�K��y�J����
�P~�J�5j���kf����I�|��Dm5���8�߸��.�[e���ص#Q�f��h���x+��4Mb ��qeϔ�ja0�������7v�Z�Fë�f�O6:M�U�0b[z mA*��-�޵�TSk��Ts�݂e�֖�i�Ѕb���־7e"g�h|��_}��ي�R��a�:M�m��u��I�t���B�e�d��Rm����[([R�kn�3F�"-�����M���̬�n��:�c7]�yI��uԔe��`�̓�^1M3BC�E�����K�*��"y�t��ۖ��U�n2?)�ʡ��=��ߏ_����c�_ǔ����\�������ڤ�N�G^�I[�2�>�o?��`�!�tJ}~ꈵ��&7e��5yo�?��=�Les�te��jy)}�C�������Q���T6�5q�i0�8��7�c����a���/v.#-6"b� 2�a/�d*��{���<>�L�n�[0߱��� s���5�,܁�����}t'���n���L�3���?���Q�s�c�.��5��|��o�b�']i}���+�Rߏ�ғ�8b|��5h��Kª�j?���7�<` ��9�<�f�L>�!ӫ:�j����JN��~���-^z���TT^���^�O��'��P��������_�꧘���xLL-�S����S�׎B	��#9C8}�J!��G<�n�E4�O�ۮ���5xП�ª<
�q~5�-�,E�)L���Q�V����=.:��2����"O�*�N��<��
��_�/1�	S.����<g5XY����t���w��p]�������W����B߭Zc�t�q;f�l
@*��Ei������I4tɪÛdn\��5����L��Mm�5N��;�C,e���"��g��u����ۄ�m�xK�X;��L��8�?�J0�r�����}c_���0���k���^�&�d]�mH�~��a@T�5z/�;G�Tx/�"quP��b��r撒sX�S�c���d�>������R��kr;�bm�t�ܟT��?��è�a� �=�|��<�d��2"9�_��S�O
��Y��ۏF��t�/�{��SڕS�42�@X�^;4����z+n�>���x�����̓,�Ӕ���
3|���g���:��o��Vc�3���h.�K�g�th~#�o$�J]m��!�,�+~!���}�.8e��1�����i1�xM1��?2�nmZ�o���	���������W���e���ЊX	]���p��p-�@&qh�´#A�RSkEˮ��bp���E���w�vn>Z�p_���ަ�=������AeI!p�ǇA�>� ��c�=x��s�u�4��)�j�u@id-;=��2E �����Q#np3]���,.��z��R����;�\f�XI܇�8���ٗ�뼬yx�}�1R�ϧI�O��lS�G��
�r:9E#g�l�.�����h �.�q^v�e����.����Б�B�+؈�8�*�<���8��ښ��0
��!�����|��D������enG�z��S�Y�_4�߅U�Z�Nv��uÎ�r(,�z1E��~��j΋�;�6F ���f���1и��Ջ�����ЍT�&X�1���#����.�x�}!y=��^�'���+���ͫבK6�Ag�R�Sᴩ�����;��O��3e8i�ow�>^_J���e�c,��8�:�sG��AL����骾]N�0����5�}B���³�������} �PA�w�� ��)5�{t�ز��@,�>����NB��ҿjX�c|ɚ`YWGPKAH=Wd"����!jt'n!���I,D0c�	�(���ϖҵN-ٔ,������'�D������d����iB��!�����jOcx�0�uP��D#�H+��$!��6������@Mo*P$�!��J�Z�>����z?19'�$�z��`���?=�2�v ��r�uDG{����R���C�ё6϶x����vY�7}�pZ`\�h��9���U)9�I������ٳ�p�잣~X�O+�>-E���K=�ӝ&�[� &:��DnA��l��\��YU,ېv�B��_껩N�����ʘ����)�t�/�%�iO�P�Ǒ�Z�@�k����F�bq�L�PU���)Uة���e:�
����sf]�Y=����EaV��iW�ӢNK[���	�@���9-|Y�C�<f�cg%zЛ�5	\e8<ԙ����g%0������R��B��X�LP�LW�����X���/�d���O<��Z������J��A*Y4w�v�ې�ʭ�~䑼v�n|1�EYI;K����x�f7�L�N.�W�"����2�83���:i�(*(�6c�B� ��Ɣ�CtǪ��Ҁ�;�sZ�	1�J+�����T�(�z'��ɮ�`���`?{���1G:��\`��|�킕׭qd(�{nw�P(�Q��M���f)0��<��Xп�9�m�أ�bU��4b^^Ξ-��5���X��#�Tl�y����;l&G��]ʴŜmR�ݩ 9v4st-�j.[^���K&a��*�Kce�_��^e�=LXϰ@�B��7F���� �D����=� �:e����U
%n�kܱcX�]��[���]H�V�1o�t�g $n��i�mKtjMAᶶ�n::�mH���z�c�fIoA5&G�����SZ�$�d~�e�%��q�Dm�L��H�#�Xoh�
��Le-W�iW)'�c�^�gټ����^^Ϫ#� $��J�}�o;�J��o���1������ɛ"zo��!��i�܌f�T�[ŽQθ������~N,@�j�[��ҝeq�n��1w�O-��I[���� pdG;�^r�fR�ʌ�4m�����V�(` �z&��gb��<��7g��Ι�R�g&_��<�#��]l��8͏z�	�c�%��he�Ev�ӿ!���6!��H0�3��p��[��xg�%�
�dJ�M�K�I� ���r�ݩT��q`)Lb�"�!�]�=�x�����h:�Z%\\�j���٩��*+l+�p��v���Eni>�ɥª�G?�C�xJ�.Ʉu�R���D��*)&#��
f��.������Q�9�I�O &$��A=k+_��hNk�j�u�vX�q�vZ�|,��0��W$�W΁�  ����l�*�`P��|� `�t�UH��,Pp���fx�v��������g��,F���1�#$lT4��s��ß?:���tH����"[zާ���s�?�ڭ�w��>��P�#g5�z���U��V���Bb'�=�/�����w��L�RC��� ��:���7�2eG�=�'��s�� ��⾌W�G�ED�$�:�%��F��?h�	D�[P�_�E61�B�_�KQw��#*0��=Q�GW~M�����0P`b�_���֟J-��r	
G�7����u��.��_�\����vN�]~u����w[mk�������0���, ����H�ӡ"=�"�Ȝ��V&�f�S�*֍�LHl�~"��!g�i�}���dI��:�^l�RX��'���zQA���nۦSRb�p�e���cH(�0��t;����h!���|���������Q�&�5�zl,vS/u����h5�#�H��|}ͫn!0�&�^I�AB����jZ�F�?�l&p�	��r�?��h��e�g��K�%횩W ����Ճ��������?T�y�ǣ��-��I�\tz� � �ޯ�;�E(a3z�t��������ekNձ6��L��N�iN6"t��[u���K��d��^t�j�Gf�,�s��	U�(Q*��Q��O�JL� 'd���DӖ0�7��U�û<����}H���M��z�L�'�tR-e��@�?�4I�#��Ƌ�1����o��<<���c9�[�������*�2�~8��Ƨ����A�`r�F,§ӆg/�}v���65��K٤2�����b_����ܘ��&|B�ؠBL�̽�7��W�(�4�H������6�yL��r����S���K�-XHfS���L��"��	I���6ѥ��8����3N{����h����b�Y�^�Õ߃��U%�H��)�˳P�ޒy�WPSe��+�y�:Zܝ�^~sgr��fº�׀4�ղO�Tl�/�n�,\���.���(8����{�+w`��R���C8��k̑F������L ���$��y�����-= �)_�ݗ�I�p���p�e5�2�|0ƃ;e7>$n	%��h�xȈ�҄܆��AZTD��X�t"�������
z�j_O�������"��Y4���xzӰ����9�rEz䪦D8K:`������#A
��|�tx��tr'&A�I�� ��3ѲmIU]����T�ܮG��&����j������m��H��X-:����M䞪��ȋ\����|B	~�4S�^�9v�qi�SIL�~�GF5�DQ�h�ְ��M/MU��;%�<���8���B4N���^�qOa��Â�{0�o%q?ܔ ���=`�`|��~R/[5��:��d��W���Q��FK��Ok߯�mn�� t2
|ӈ��ݧ��{��;C����P�cn?��Y�-n������݁r�mY��=����d��`Sz�y�)�]�?Z�K��!͵���+�
c��xp��F MDmƾ���-ɽ{r�=h5Q�>��3�"����{
3�*	��ˁL�z�샪���.�n�^H�0+�n©���IA��Cx �� �\I(␣���B��d|'��5u����TX]��:�S���j��Y�I��
�L�8&��UbC�%���g�X-���g��w�L�
�"��!�9����3e#w�Tٽ��4"ec;������g!��$V[Э���,f� C�+z@�ڧ,
 y�A����c�+|T�;3s{�2��@�����+�;�r[�x� �_S�qb�ƶ��a����빾L��X?�LJ��B��t#��׳P|�HSY6��(F|��3��^jd���W�Y��{Y�L��M��Vx�}>�<����;�:X_�v��T�� A�W
p�y<L�!��
��5<ɇ6�#(;V�7��a��}��U��?7K�!�jM��(#Lz@����:��7C�N3�mtr����2�J}�I��Յ�lk`HA��GC�ܷ�m5���A�p�OEh��IF��5�讚r�<O�7�s*�c�g�5O�F���
�G\oZ!f1��iB�Us�M��
!]�d6t���]��]s��K����D�|����cK�R�T������ʚ�؏�絧v
C�dN�A~6FO��=c6�W��ˈ���@��	����wZ�G����S]��%�-��p]�t����ۍc�}�����Ϥ {�hO��P6�����6�{��E��~�D���[X��vS�n�� �=�J���i�j[�v�
�c /���Bc�����ޏ[d����F��m���E�hEݏ�#<y#W��J��xt��uq�b��np)�����H��G�J�j��@P�d����`�v<A�������!n���Z���d�v��+9���w�S�_Eim��I��_7�b�<,��a��27��]QDZ�~FN=�~Ok�il�y(*:Ru^�z�:����?�Y�5��U-��5~�߅�8�PD�Ĺ��J�����}]���|1~���+�����7E�ٛ8t�xb��e���J���P���6��p"L�:���;��A�'�M��@G;��]EV_��)�?ϼ�w�����zĊ����ƶ&��@����B�5��������Tv��H䒄е�~�������:]#ʆť-52�5��Pc+c�Y#�.������(5��h��n�fm��Q9�ZT�G���3~�a=p��� �[	`��%7������)�C?4{�5�{����Se\�ގӄ�'�E���;�C�}D���� P�?O�ak��۵��yl����\�y�f{��N}T
���ŊJ�Q�"1�D���n�p$b���y3�?�ט��[a������`�vX�fPA���%}�\�Q6�.�ⳫXoPz�������Hmw�3ܸ�L��t�?�Ƃ�O�O�K�܂7]F6$�1L����q��N��J�#����t��kv^�8_�r���I���[r�,ꉫ�8�^E�e4�Y�쾀=�f36EPbM�%2�qM������a��C^go��4�u�r�/��i���\�eN�,��i�l�[~�\�ᇤ����(��f�۠��5�R�H���{�	b�T�,��Ǳ��2�.F�)�J��h�YND��>�K���}\>�X@�;\�����������S·�Ӕ�#v���D5e���ME�D��qNrlE�xjd����2��/9T!����F�&]��>�B�^_��;�p���֒���#���{<F R@*�S�u�&����dc�!�**�R�M������h����>W��+�	����#d{�hSl��:��CX�[��X%���%G|��@��܇f�-��D�M9��}_py:2����w����P[�	��������(���]7{�����T�=W�W3� ��	>�s#�͊�
]���-��7�	�b�P����I���'=������41�}���(ܷp}�[��fд��LԬ=,'ۯBD8#�<(vmR2P���mw1\#-"b>EA`����
7Pl҃]g���Q+�(&o�g�>��Bڗ�lJ��SOkM�.�c}�uz8�h*��KB*���^X�e��e�_~z=��Rh��<@��r�$U���iX��
)woJ�'���O�.�H��e��'8��=m'��#A*��|L�J��z~�2G&i��c"���!�P�&i��t�V�2�-�[�4@��c$:��5Jk/6]f�C�d�0�i��U,��*�d��*%��d�V�KT�bw��)O�0��������XYv�0W��	�I�y4T���Q�0tcT���ۂ�p����.=&d��^R���˝�N�a�,	f��2N��rT������R^�dN6}5p`SW�D�ܟ���#o�m³ցOs��j� ���o03���@��b����K]|�B�-�[���D+��s�}��������{HI㎡Q�R��iW�v?�B�8��X<7�!���$7LZ��(�Z�-�e�[�FNcl�~Z��Z�$�ک�C�����(��$:��	��^��H͊�Z�;(��8��׌AGpN�A�p3�?ᖧ=�)�戳gd�M��-��O��p�T�xZ���pN������uZ-W����C�Uu܆ʏ�FX�"$Uo�O���³���n��=��C�m4�0�Ԯ�$%P��l���Aq��ܿm|��)��([�*L�㔵D�s�;�A=��y��'��>[�qJm�;sh��U�h7����?.��=��面�ܭ�ҭ s9���w�F1[�ЏC�J{��
2`s�[����$�󋄢��9��x	�@m�,��=@(fVC����:H��U�����?�W�JƤ"ptM.��z�7��.�]�� ���a0l��?���!|�'�X0�.���UۂN��G8����K�j�v�GZ4����	���_)��]ip�J�8y^b���y� M6oO�P��O�H�)��9����T��y��Y�J�ғbhxۚ?��Q%������i�!?�g$j�]�R,�D8K��n��5N.8B{Ǔ�.��S@3)ǜ&V� ��ޛ U%ͱ\^7��^�*�=s���1�D���-�)~XzQ�m�$#)����wX�n���c°�&rm24Ƈ�}����5ӳ�#"�C�!o��S?No�\��w��2ǪԜ�q�$Yc�x���������8u��q)������[
��� �iáp�L����R"���u�b�|���pn΅w�%[����ƪ��T�Ϧ�d��� P0����Ѳo��	:|���<�,�G獻�E4��,#p�(�)/=7�0�,�����a�^�U�ӛcH���E��eH;ze@�S���_,^���(C�*�y�f����ߐH�%���I�ft5-
4�ϼ@�Z��A�D=Z'��|��/�	�%+ f����$��wo'�3���U����l�:�'��3���9��K�ۈ)��X)}y=̓)���w�k[U��w�wn~${���$�N�{�(&����H�x�N��!V�O�51�.��M��?  :��d�������b�ʮ�:�������H�OTg/_!)z�GX1?-J6ڥ����H�v���\j�Ou^�ȓ�G��p;�6�y �#��;`����2bR΄�����"��.�j״l1O�Uv��(La_l�.���3R�OÐ�K��쳻dOMR����<�^��hEo-��j���l�K��o���(ek�0����z��0��̺�5� ���b�q���G�x>�C�#f���Šb(e��iZ�g_��'���[�$OF�o:4���~%��gJ�i�1o5�G�U�o�3��./�.ü[��|o<��Ц�e"U�&�K�z��b[R�7�q�nR�V�[ֆ���E_	Vrr��R�;É�0��)��;`�!Oo_�h������X}H��%Z��*ߔ�!�hh'�g�8�����g��v�º�O�@���`B,d��!�c%h&PC��x=�5�8#z+V5�n�&pɥ�M�	� s��)�G��Α�
5�F��d|�����Yp���x;���=yC��~����e�������a� ��c�k�Hr���)ݙ��IZ�e�9�3D����5[�I���.^�hF:l��Q�`c��4H���4_!�&�?|	��+`��pu�;,�%�c�u�&�|-;9��2��w��+L�[�.�lr
_�C���KH�N��kK8�{׻e�;�v��p�r�%L�}u��.��b�Yq>o������h_�y��&���L� @�jø��,��VW��Ҫ��O�|Or�ì<$|��MR�B�geE��A�y|]���qw��e^~����C����"��)/V��p�89�텶��n�t�Z�vh6A5@���F1ٯ�2��*�D:��@~��~-��Ny����ݹY+7L%Cp��aΧ�'�(���� uJ�V2_U�v~��3"i�_#�C�1�¬�F�X��ʾjX�����q+�=�Gd��߀	_o^M���K��s�{P�]-B�רFm*�O��C���E�q���!�I���`Ͷ�3���ԓٳ��������:M��&�6�)�>})"q$���s���|�4�D����⊓��+���Tq$g2����{a���jh��o��9��?�䭹?;��Snw�
D:5D�P�Q�O:�����F%�D�&��J�O���/HxJ2��;*�Yq:���t��LZ�ց
 �H!�\�[��J B#
�9���]���V�.I�W���t "�#Й,�
������V�\�5��)~���JZɮ_��gD��
#�`%;�قh�Șm��y�5R��^N�i}��Q��,,E�p�ʓ8W��C�ɧ2�j]�_閚R`F9~}8��͹�"(|}�;b������$ھ�6.�j�/++�~F^5u(זZ	��G���>y&m�ѐ����V�ܸ����,vl���R�.}�	Z7���G+,���!���?ntT��M�rE�o� 0ڠ�B$�}�^.����8����A�Sf��骆1�7B��I�OI{��z寵H�涢L���B)��lݔL�;{�3ɾ�Y�CR�j#��/��q�������J>-�,�-�J`�������<FqA�N����q`�(�Y|N���/�G^�*���`NG}&T���g/��逆Yp|z�cȐ��[�N����B5#���R���1m`JѶ�c܁B 	���MM���ʷ8Y���N=��W��495KF�A��]@ҮA�%|������6��!z�FWc��&�?����V�~�v��.Ut�7%}�ff2�ꅃ�Md�1�������(�4ʬ�)�����q��V+�]C4����q�g��!$����Qj���z�J+��}q����H� ��&�u@g$���DP�~:D�~Ӻ���>���Pb�:�.�%s���
QI
�ۤ�h�:,4W�]�V�#�'h?R�6`�k��]~�ǩS�8N���%@���-=t^��>z�<R,2���+2�
�5�7݉�M���s��U�1L*L�Ɯ��D�/���g�d̘(��3��_&G�+#�*w�:��]�JP�����k���k$3a~;�_
\���CQK��}��Ơ�b�5���/�@HՇ4Xt7~�J]�MZ Ќ[,��1S(����� L�a#!P�Ĵ�h	�/��%ٓ�)E���1�շ�{"6���gG��.�x��0�97��`Y���%n���W����0C8����Ä���^ͺ��~�#�qdN�l��/��. �Vvz[}ԃK�V;�=Y;4.n�=I{�0?o(�-�*)߂nWG\�$!ہ�ht)��i�:]�A����LVu�r��B��$R9E^+�:��)t�>C8��7�ӡd�ŭ�D���7ZW�t��A�W����S�qNl4�!���8LiU�<�b=��t
�a��Z�y�VQ\�-}iY��{�q��'�6��#�����6(�A�(x\�L*����NM^FD�Ч�E�����"�������B,�4�|i}�4EDTm�[lh����0���r��k�o4k 8_����[e���R\�Y?I,���wk(�PJ�;��X���E_hZ�R�@��l�DM����y��d#E{F��T�5�����f8-��m����и{\L|���o�ZҖ��������4�z9c~ʙ/+�9s�Ofu3��R���R)���ALt�s�R!v췱��"/���]P��<?-)�5������U���Z|����n�=��4�n�ý�d^!�qJ����(8
���\Sy�L�\R���v�ɋ�t�/�������&�D�9tG�����84�s�w`*#?j1�b��kH��~qI����QQ{��vl�+`�d[9��������\H�'�pa�ĨE��_�F�$�Rm���GD�,f�z"?|�>e���	�� ��8	�,�ˆ�Er?x��5ﯤ��f��xI'h6�w�F�����HG�jyߤ�KS��kb�&�-��C1צ�	����o����s��3�~q����o�iTz����t�8��櫱Wb�h�̟�F�����5
�G��n�׬ܪ,*t��m��u9�����|�ۍ0`�J��'�lp�9��;�ӥ���K�:�M�4�����˾O�#�����l30�j
T󰌌���|��-c��%"�{wϨ��jv(<d蚺�W���&F5ܒp���zi��ה&3�7T]�	��̚=�ϳ^v&(�v��B�������|�Vs��ӓo��>���u��|
�C���ueL�b��f �Ï��0U��-�z���¯�\�hk��z�Rbǒ�]C�:{���,�]�̧x�V}�$��w��eA�%�
0E7ɹ�7�{�uy�LK�zg��I������=�!�uQ）~�Ҋ�B,>U��DyU���T�e��2�"���Z���ͤ-��%�̔�=̞�5��|�c���ԶP�{�Ĵq�2����V`���̛���D_�V�Iͤ��e6���������@�0�8��QO�Z)�%�0 �x�>��m;	�4��ۢc4�AyC�:����u��L'��׏N�� �0У�+���>�!.gCF�_�4�`}1�TV�}��{nhB^�/ߩ�a�\�%Eq�#а�Ĝ\L�����b[�:%z���_
F�V@���ܭ�Z�m>�ش��7�(���I!ȉ�V���a��)ęm'.�8w��-4��x�]���%s�9�1���{��'����yk-j�~J��ä	>�2��sv�J��=B�s��	��2g�4ūS��8���Tm��܊Y��w�$Q�l��BN�����-� �:��5a��XW
e8-m�S�s�c�؃�P��mg�}�G�b��(�g�zY ��{��-��F��2��%/"�ӧ��@a��O�ݷ��]����WTE���YZk��&j%%���1���U�8�3_C�E�V�{�Ζ���M	4����Z��}[36�ISjšA�PuGK�ZWk�n���?b}�$*���({炁���0�	a��N	>�?m�gU~�I&�q�h�X� f��F������Th��>@��v�Kw�o̓@K�>X	��\g�#��pjβ�839��3��ۻ��@Z��W�\�c�ל7�D�u\��.ǫ&���g_;0w�=<BBv��I_��C,�.6��OI�pص�l?Xi�$�����DV�\�:�0�(ID��N���W8��^a/4��s5b��;	0�6=���o�j.a��-�@<YK�}͍Î�t���zV(�ޡ��鯶�#y���(w�1H/����0+u}�?��:=\(�2������Q��2���o;Ԩ���[6�an�OѼ�.�|��_p�����~����F��kF_�]=�aS蜮�=�"x���~�n�&���_@$c�]�{�Y�����������M1ּ��\&��҂�R�#��H�%�^f�ADl�㪪����?i� E7|y��K ��^[x�A�b����*��I睽�f9���/�މ2�CI<6�5���ˮ.�F�:o��h����8m�q}�C�<��#3��1%��s,�iJb����;"�;��)��<��7�c|���(�˼TI׾�M8����6��O,�	��.�H%63UA{�ău0QNǐ�Bkk�����D̬�fNηл�r�ϧ̠-Ơ˨�_"�����C"��˖��xF�&pc�iE�����R�b��2��;,�x7B@��Z|�K`�&U�L��mu4���F�G[R� ���
1L���rpɽu�ކ�_b=����2�>��z�uT
��8�R��x�VX�ŧ��D����]E����߱8.}���<���O �%�>
��\&P���@.m\���qn�/ى(��;E���'�]<�N���a]�\Vs���gJdJ7�2ܯ+�7�ozD8E�ym:�����}W	�i���1.��&�UZ2EN�iR�6�����	_{2>)o�ko�F��N��X	�<`�s�z�K_x����~G��2d�����H����2�g�u�kE̥$���	��I������^��}޷�K��u,���%��1�Е��}1�&���@]��u���-��v����Q��>�+aGV�p�k:#�N��a�R"aY��4A8*���R��>�fc��L�FE�.hm�k�i����� �L�TW^v�(�M�#\���nܞC��T�4W�_\hƷ�ğ��⺬��@��<����*�'����45���*{��F�4��ٙI�2������L�>}���^B�R���$XUTt������^0Yc����Q�C���l�|�֙�Z�R��1�P��vz�z�� $�]�.T�x�t�0�X����R���ȕ
yy^��*}��A3N�#�>r2C�\����?$� �|<6���9_H7MA��/�l�4Dф��)RŘBd��!~Pɞ���O�D�t�R�R�ѹ-�Ճ��"��*Tc�@�\X f'���\���W��Hļk[L&��.���ج�G�
�l��\ww�=�qF����T���'�&���l%��h-&GT*�(
�ǐ`�OI���y������;)�k���b6�ا�nOO�'J�v�)��J{��[]�L�<��@
]��b�֍�ٻ�`�d��=� {�dt�/P���9B�0/���6�(�)�3I�+���!T��ыb�;C��K�� �׷�'ip�����O�������Z�����5�8c�8��p/W��ס����Ok��>�I�������c��Y!�b��n,j�_N�5�l�❥���
����>*�i�.���"�@�;��O�E�6g�X��O>���A-4s܎�u���r���FT�x|=�HNd�xK���ur_y�&���:���(q�*�vp���ы֧�Qdp�L�h��������+��:�p� $O��Zj�S�e_g@&�Q�:S�� fw��l�4�+�)�	q⳿�W�싪�sX\}e�0�k�}�m�8��Ũߍ=w/��\��A3S�/'at�Rl�Vo�� �
� �-%q蟃2c�Ѓ�{z�$�!PR������B�9��ɛD�x\�dE�
"Cr����ec����,���w��qN�ڟ���^*ss��1�����!�(���qo1�İ\����eqS�3$-�rCC�<a��m �-� '�^�Ы���[��J��D�W�<��Q��)3BOY\e˽>��7�z��/�w���F�B�V���I���h�ZK�O`���~b���b��)��m�U8�#����W(����j��U�f@�.$ ɣ^_��*��{�i��#i��9�dK�l���]2תYv�e�ң{�4�2Z]�T3=M|d���T�^�����[0>.B
��$q�4=5)��RY��W�WbX��tܾ�ԟ�1C��9p����cR��7 ��G����XLd�0o�7����Y��d��$4 �_��%S-�J�I�)J.To`4��Z~p�qINg�v(�Q�$���`u���}��/U`|9x��!����f����Z�YJ��!�]s7Ҿ�$��\7P���;�%�Z�7{v�:Fo�s�)��Auc������!B	� �݊�"�^�����gS��m����w�}Z3\���1��1�U�U26UP��8��k���7�G��)-��Wd���5E1�%�>�0�S9�� D_�Ī��J��?Y�!:�QWhQ]ʹt&	*+���E��`��� �
Ȍ~\�Op�{��/�Q��^�B���i u��@p���#���I��J�]���bδo�_�R*� ���q����Ӳ�*��Q|tȜi��a<�%`jl�SY�r( \�Ư����#�zH|�T������K��N,���ն)Mw�#XYQn�mHP�0]���ū!+k�m�l�z�ۮS�zF���80��q�P���۴�~jѶ�M�� .�jq�fA�$�Y�i�v2Y���˞EK{
0����D0�b2�I������J�z���oj��DyT��d,�}
ӈ����t��u��>rS�Ӡ�z3VJU�ӱ;HjD�@��&Fv��{Ht�����R�o��A�N��l��F�"��x������@������	��'�'A���]�c�����o��.��[��Sg���plL�_9 <z3�zȅ 1mU2i�
�ʪ���^ùxCaʹ3
�~�\�e��k�=��|�����HdY���۲I��F��##I��ة�E	B��zS�&>9��0:�pL��]ɗE�\5�7Wvc5����i�B X���}%�{�~S|���D����N%���|�<7��N3�����#�@ؤV~IΒij2/ �U:� wS�����Gp���A���X�8��3�4��b�������2�qk��ܸ^:����1�-|t�(�B!IK��$�=G�ҕ���x��C&�'Zƈ�j�S�$M뮐����?�@�a|C��(8w� _�]���n���l�ւȳ����*v��a�℁��(�wغGw#�ED$
ܤ��g�ѻ��W�}�J�o�Al��a:����$4�Q���ѕ2;ʦ��M��+6gX�7��*�n�� �`<�Pӆ>�;��z�+r�%-쐼�@Gan��'��O�%��қ?���VFτ��/P'������tt[�P �p�wm�v�M���O���O?k˪�O����{+7�_ZJkQ�$Hc�C�[�'�R5��⿟�H����qG�s��8�B����"�M3���4eD;|?I��}�ԉ �q���Cz����Y��wk�b3ȣ���[�4����!M�?�p�ED����zI�m9�*!�P���j_-ZDw�yG�V���.�Zyϓ��?�������H�(��m�專�.���֕)Yɺ��n�����Y����j�׃�R�B���`���u�i�����זg�/*��&/�6�A6�FOAx�� ��ؔ����#T�|��K��͉�ĭ�K���ޞ/^����ąO��Ǵ֘0a[�{��deM���f�����]���0q�-�u+��f�a�pl��n���, 1< ��B1F�+�%� t��YE���y`�ϖ{��Ǯyà�%7��R�nA`��.uI��D���J�N�s�e��B�;� �L���%H�78z�Dv��D�i,�.>!�C-x���׫��M�箿�dU���77N��Ƀ�&^/�Wdq�c�$3q�s��L�Ǖj�<X\Y6��] O�l�@������*t�ֆ(>@��k�_]G��VI�>#|��n/r#4�
�P�x�<X���E(����������Xʐ��=�������nX擌<k��	#��Q��Cb׃)�Q`����XB�8ٽ�eZ�L@��ޛ�e��mE�,xA!����VB=���B�� Ru�m���os��n=��\@{K%�o҂4�����I���V��_�"G:���c�5琑|�Y�5��L�*Gzڷ@���|�\��5P�����D����X<q5�kg��ؒ}˒�${�a�}�Fh���,���B��ǌ��P�'I�B���Q��G�=���qͯ�
X�T�Q�?� �p�5��"��s�7�cC�� ��j��lhՄC�8,O͟�`K��+���9 ����s� A0�&J`QjbYA?y��h��<c�<=b�Q�g�o7O���u1
%�-�zaR<��T���ϠV&���񒓖��aӄ�R(�5��䫉y1\5�#���˛cY������*��?�H/�8Vq{�u��+3G��	�����*V�ep�YD[�&z]�S���JW��:jZ7��y��z=qt�P:�DX#�ݍ���4z�FT��96��Rk�ϒa��3�������S����a	�z�����?�@t�����y����Y��k�j��JEp�T�������֏r�8��F�0�v�Ź`�V�Ũ���pe��߽K6�|-�|�iOi4�\*�ܳ�̩s�R쳐/^�Tj�-7D��k�4��h�f��-O�l�-�������<(+���� K�?��^Q�'�5�3�H�֘�q��B~:unP|���%5�9�4lB��
�R�}�'��'�,�>�)PK+W�Kʟ��؆60�`��	����0]3cG���m����{�i����	&*&��b)P�!��ϧ����c+�I��(�S�|�2Z�qv��I��{4XE��lA��<���:i赜�;����Axh����D4��A8�#*3�ݢ6W>�������Hx�i�RK$9�v[����I.z�6�w�����<ӗ��O�B<��B����a��6nF�p,�wT��ˈ쳫�"��Umn�'��{�ᱤ��c92q>��-��"��~�[�h#x>���[4 �Qf!`�%j�+��Ml��C�4"���Y�BC+�=i�������Tvʜ�f�A�&�Ĉڨ��	7�&"�A��}<�D� 1l��nEk%�F��GrЯz ]=���xu�C�_�I�=��0������un��~dT�e������ә�ߊ���|J��{m�3U␠��vn�t�5��ۤ �/�]t �g-+h���C��i@4�X��H��T�;�+��̋���5��vN�V�d'^պ9'	Beh�I����4��b�'�L�`�,*�j�/�or�l{�*B�K�2t�S\;�ͶE�e���D'^���D~���|l���H��e�j!q�YY�u-H+6��UcD#_��+���i�FB۫���,O _��x���U_�o)uC�T���%���
����Ʀa$� 3���ܜ���8j�'d �:�zkˍ�!��E=Kr�X�A� �׼�yi�wx�� �����)w;J D9���ҷt9��p��:��k��6s8V��1���'�ЬT�m�H����-��PO��i�5��R~��:	*���P����-n����]�m}��	$`p:�`�Z�8�S��	86��
��?V��}Y!��������n.p2���g|o"|I~��b��J ��˝�Ds���%���C�8�繘ͥ5��c�U�X�&�h�ճ�O�)	W�@y+·Qz҅�Q�����/�p��'�\t
N蹾���	��Jz3��T�xӛ�4���L���,�'&U:�>P��^�!�b�Kzf�fH��Kj��سTVAD�]1S��"��V�I!B���,���(�e�^!/���@]S's�G�$�u���Є�|�9�J���������Dk�f���U��D�����2n%�k�n�d�
]Ѝ�pN+�������z��.�a[��!�<�H��I��p��C��L���DF���&����B�X�����������x��e]N�/򪒽��A�<�º$*�l�+��祢<2��\���VZ������A!]�ђ�e���8��Ėw�&���a1����Ӊ���k���@W�fe���P�ǝ�z=͊K7@yLÊ@,\4!��`>f�"�إ�ފu��,��e��]��Z��gM\v�'�7L�򬀿���<�q%���7���W\�K~I��?�l}��I�?�������_0�ND��:`����=���$LR̍���&z�J/ �[4��?�z4Op(�As�	R� �b�au"��o�XLV`UaW�}� >M�f,��`��<�����5�F| 4 �CIߴ�f���dA�zϢ���i|����2O!7�.�I�c��/~qO=?晱9�H�",�	��Sxh�ol|��;ʮ�6��%!L ��B�&���i�=�Ͷ��X���/��F���i�ma��
	����d^������{��rLs�)�9�4����c��>3�uL-�h�����uv\,�e~��7�Q��r��k������l%�:�����4r�2���4��V�h�	�c��0]����^�`ٷ$�1ī��֛��)���Eu�h��X���cݒʝ�<�역�g�L�@�\�xR0�*=
ec�+7�t�00��DA�2�1�� �йd	�{�m�g�*A�92gn���D���͗��kl0�۰�#�!{f�ݨr���G~BKy��T��.�m�����l��+���z�C�G^�X�� #����QS:���W���p'Q4d��7绰�@�W����"���X�U(��5Tcv$��"��.���w	?ȉ�N��Cz`wM������hˍ�]0}.��镱)��:���o�}�̻��j�)�����X݇�j���=�0�,,aQ�X��?�g.��ϋ���2���ݚ�$R'��-�l�A���u�NUO~�j�)���@ѵ�r8�$5�6�
s19�{%�L?�q$N\:2���(/�e X�7v��z]��q�٭��ϑ ��;�1�Rwf6|�������N�}̎�Y+�J15�c'�Ζ@��{x��hm��$~VF�rs@�dĻdo��K�)p��w'�1rf$}C38m<i��-1�撍�?T�� c�Ij��	��bU���.���w9T�#E�_&pI�ڨYt���NE۷�����t0��E������Ж��v��Y?��5�R�Ū�����1��N"L:S3�*ewkLb|8�V��>~bΞ�ND,�vM��"�	���ۋ,����1��S����ʿ]���a�Z�����&�az�J#�D�l�[�-�tr�	�T5v�!w0������-w쏒�ò�a�J��d�rf>���M��R#{{Z�eV�!���Hם�`���4x�0��{׃����s	ݓ��S�F���[h��g�6��< .�a��G~ �n�����M�����5&�nL�����s�:��^���}��(_?�B�i��}��=M��d�)����U� �IbYS��<H4Hr ��[�����OP��mV�?}F�ï�º��됨�%��A:�n��J�x���2N�TK�k�B%�8�)A�G
»��X읯���bނ�^L;i�,�HHVFkKr�ZM�<M}B��j$��O;�o��y �$sA�}�Q�����=XrڒyQ����Mg���f�­(�jq�3U�/��Y�EՋZP;L5�C�%�^�6��Y����U���B���l���C���L �07-�W�ml�S���8�0 �a2���d�ĹJ�u�������#�%kF#R�p��l�!K�X�TFhN5$�;�m�:F2���2������t~�m�JDe�)��ÈQ'T��0�$.��f�#�r�l'�1���eZ寊�`���}�`�kt�P�*��m�@�X6a{�=C���Q+HR������2�p:�T��&�;)�,����T�Y 4�5��/���<��H��z�~`�*M��z���z�}��鐱/��6��Ȳ�W�+�_� �Pj�Y����V��SX�����ka�e�B�",J���p��g��ť(���P���%&���iK`�{r�"v�V�ž"��7ۗ��$���a�R��i}��)E�~74��H>��qu��&�S����f���dxn3.�&� �X"bgh�LId�`=��pJ����2�gE-D%T�����4_�P����49��=�H�m��j��]<r��wzJ��i� �<	�<i��j@�հd�{�� b�����V�0����
.�������R��fƥDa��`�f),2��(j���Zߚ�|���]�:�Ơp���|��P�$~���\�1��k�p��D^*�i?yEf���8���=�PE��>h��@�Q�I����?O�ML�b�����e\Қfuݤ)2��Ӎ���$����M�E,�^P���T3��%3��"�XE�i���]+�~�
�(=�𸗓�P��O�Xb����Ո���q�#��	��+-\�n��5��]�8L���,;��gug��������$�����g{vY]���d�d�8��
jI�Ѵ�7d�u��|�r +ݯ�EB�a���޽����p喟\������("��*y9B�@ǥ�p�y�1q�Xd7�I)nF9��v(��I"��h�	3�F�H����10��뉣�<�i����5��~S�}�%5L���6�
\aD��GЍ�<&v��E������l�a��^��j����q�&He��g�M���C9���|�&q6��4U��&�m��D͡?���dw�^�M��+9�+����3��<~p�_��Mf�7$��KX������BX����m�M�Kt����q�k�֥Z�Ce��Qp��'�'�(`��i����
�k�w)����g����L�3
�Fc�"yZ�8�U��%�Ku�Ď�#U���[ r�&��Hr���vMQ��G� m(�q)n6������"Bg�.Mv�T۸�(_)=`�5)�1)Hf,߅в��Gf����)*S�;��<��%%$�'��<P"
�G2e�Ȩ !��?C�c:QL/�4��Bᶒ}��<{j�rnkݍ�V�:/��y =)��g�`\H���Xy+L�%���v�غ���?�;�%�#f����\��h�����	�؛p�����k�QiM���3���.ż�I�����|��AO��y�-5;^;a��5�7Q�a�#Iwf��S���
r�@����aC����iȝ5�~��^���RG�;��?r�4l"�Z;�XaJ�	>� MZF��e�7�Jw�|���ኦ�:�O.M0%M��d�Sa
��c�:��v'8Y���Z�$B�Ɯ�@��۫nT��D�>�����%�mA�^�Q.��|��:%p���o+�6P�ݲ���7�B�T��j�De[��{n�1����#<5`���Qڠ6����~�����J���mɗ����� �Ѽ�������I���	�!aR`��;g��N��(�`m<�1Bt0'�v�\Ih�_%浘��'�Y�̣�5�*�^��+2���!��4�W��c�&�U��P�����]YI526S!���l���`Q�_�8������������Vh��bq�Hg��A�drfh�](젆��S�P+�~��3���3R��?�5�����I%]�Q�(��=vh�^���<�:��3�]�&�L�i�,}�1M��{t�7w���Ko\�0���v����Ur��®�[�tJ�ew������݁[�*ye&WD�	����ˍP�����{��S�u�3�»P�_a�3����A�f� a���d�o��������$ð@|,aK,���g���(r�7�'+��q�-�Y	*�)SP�F�io��|�3�$�N�#��{��ZL���Է֫^cǕ	5��+�Z�T�Cݾ|�F���ɶ@$[��N�mwr����S�x�5�TC�+i*�ے�(��d[�W�{�b��5q�R�Zg���-$��Ą��!����cznұ���� o�g�u���&��K�4�[q��6��
-�:�n���<��O�%#H��_�u�v�[o�3&�(PL<�דAҊ��H�@\Z�9���p�M�7��`Qጒ�ۭ�f<�$6N����ΜܿZu��;mg��j�t`K�E��4 ��c���M��j�I���6�Oq/�HZZ���ѡ��;<K2�v��8-|ᵘb:�8��֑�pr������
M�=6��ǐn��&5J�}o���Q�K��j`��c�ѢF4����7W�Sv���ڽBn�!WB"[m������&�L��@ZN�����]�W�8w-q�#ϩB7��ݳ�`|"��3tм���gu�nm9��=[<B�/��x�\�5��1]IjQ�~�LN��Ue_< ��='�_��b�?3���*�*4��a�ys筆��z1 :��pH�$#�]&�����&%������t�=?&8�;}�gW����E��\���#��ᲣE�[�ܮ��]_�B8C@�?�U����J�-���*+_~��6[�I�_Ϳ,�D��	s\O/-���\F+�D_Bwf�I���%�nY�d|���_���I���4��7Q(g=V�Ϻ;�@���0�(���fU��-���sgPK�\�l�7��z�"m]`WQ��o����T�p���pfv8�'��L�wtN*/2��h�t|%�E��wۣKx����Ч!`)��"OmEM���}K����ϭkM�z&��ܴ������WsR( H����j�_P��#]��T�#ySPXA\g�ށ��	��4�xIN��;_��O�'D��c	n��\uT�d�yJ��3\�_��ӰY��g�An����kn:��1�&dBV�K�����x���:�|�}�~=�c�U����Q3s�

<��T4v���	:�(x>�ޭ�b�`m�G/~F�Oc�Sφ{�~�kq9RPA}�d5w*�<�L,��{�Ԯ��\���V��j����y(Ɏ�CPXL��D��E���s!�=ߚ-bF,xE��T񙅃b4�y�TLS�r_�f+�	��8[�����P�e�f�\.'�$d
�<�%Lk���.d��]��� WN<��qo����ף(_œ��?ٸ5~&ej���vW"���?��;!-���_�D��> z�2-1 �2���,W(����$��������S��,��}o���ݧ�������l/�8�^���YՑ������ڞ�=!}�\�t)�CF§��Y�� ��e�B�$?�{m��|WUn�881N:L{��gl�Δ.F���<l��MQ�|�î�q%� ���M�Ec�5��W�vM�m�����MVP�&�H���$_;<aGG�Cr�J���Fm������n� @)�ed�ʬA�g~ۨ6�{��,�=p��^�dP֧��~\����c�+�I����g��������@o���qР�sE�z2 ��>�6��-�A����Z��9�/|]�Z��A���	R��^.�;��ȑ��)��b�U��𾇼�Jv��"[�Փ��������M]��G�hV\�|�R�#b�8�T3!C K�(���E��8:jZ�m�ܱ��1Jg�v�{�|��)D��4~�zM�����d��⨄b�gps~@z.�&D�%,A1������Ȝ��D aUV���+vv�h>.u
>{���	�^�<�j�wW�aU�h�J�v|�ù��xP ��Ǝ��D��@
�b#6����y(D)�{$��BX�����.�JL��� ����� �x����Zœc�м>��oi��pl9[L�1_�i��p�3v��ii��)�<��A��f^�Ԕ��9z�	�5�DJ�qu�|?�N-�Qڍ���V�;�k�����\W,��сm�{�����$�A߮�T�`�u;�q.�y�a@T�ǁ��XW����iʈ�f�afb`#?D(�����:�~7���� i��Z���M2	M¿_��HFrC7�Y�`Q�pҠGn�A�k��UK@R�3��/���_�l �<J뻷z���TaS�`2��~ƿ��v/u�w���P/�!` 2l˫���D��s;���{��Y���,���T����lU_�!����:(0RY���y��s '.1���������+����M3a�5�.$�l3>������Y4
�V�*�����i��Id��آ���A�a��fh=�[�s�l�}^����Cz�]w����(=�m��e�o�=�z��{�[8n|ܦ�/��<���x���� \(���1D��H����g�,�6�G�S|�Oa;�7͗����yĭ�$���9���0�<a���hU���za�,*��A�zuf$<�������c6-��:D��z2�E����~����3P��rؾ��3�As������L{a*����cE���S�|�Ln��s)��&��q[�������o�	ܾA,��VN�>�i���4H;X4�,�6ٷG��h�wJKI�-j5Ϸ������c�X�CLd�+W�Ɗ�4d*7)���'���$5���G�/
y�t���t�v�!��O�A�Ȉ�U6��lH��\58R)s�$p\p)�HAk�x-�E�����%A���N���K&����E�V	?6t��w������8Dt���)�Pu�r�����.��N��E꛳�8 ��B��^�?��!��g�Zr��.��\UIY��\�,�ý���WTk�;xᣄ��BC,I�#�	t�+q7�
|B����6u|sԞ�k���ϸNR <*Ǩ�2��+�վ?�^!-e��^T�v MѲ�%KR���ߔ�S�\�=}�;�\a�^�FS�ֆS����P�|Ds���u-n��\�l�Ch�C�4Ӹ\Q�Iҋ�Rjr��TJ�r!���sfC���V�az��C6����?&9�*�Z��0C �"�#P�� Í�8p�3�a��:�B��@���.�%��O=5��x4����e	�F+���.�c�g�z��<{�I�Q�����]u`gH�Z��n?��K��B��~�zY�:�~kH�H���y���e�^�T���Ǯ��
)i�6�S{f���:h�_�z� O�Y�@Dyz�t��Ƭ�>7�aE����0|�F?�� qLq|�K;,�.��W.$N��=������}����Flg*�=q��%�e�6���|���@�:�-��.9�.��{���?Lu�9X�$���������c��\�Խ��K����+��0\���%�7/���LGl/��<�V�ƿ/b�,]ׂ~ۚ�G[�٭�D��e�,����'Cp]�C��l��R֊�B`a��� �C���;6�;��;@ʂ����FL�	!�؜>@�7�0��t����G�k�hhh	 �UU�E9�˿!�a��*%sQ7�le"��W���[�o���p��B@�pٱ������rIÌ�/�7�S�I�bʺ�����b�dC�;AL���O2PD����~r�a��=OY=��J*+r��E|��(X\8���P�V�������Zh��k����ixc�`Y��.�T����0 ExYO/5������+��M�����{��Rt�L�gR>pe�a�G��.�S���S��l��ҝ��P� @�Wo�F��r���>^[i��{��k�y=ulРC�����A���F�"y�7k�Ĝ�_�����.Mp�ur�^�&뗐��kϸ۱A�&D}�w��p�vH�th�	eϽ8�$,c���] �U��ҕ(0��v0�&\�3\2�C)c$(m�m/\z�b�\�hF�3yv�Ǥ�r��-�e6�P,i�Ni>D�DDtJ�M>А��_ �
;������+O�LM%��*�/T7�C�-�.8+�U��Ţy��o�G�Dsy-��~�yӅ���wt�$�)�+~]�_�[뾸����@���T���}4��L�"mE[~�0��z
�Δ��y��R�h��>ޔ@9�`�a	��Y�^g�����!r΃��NN��d����3M!�U�Ƨ̶��P�t��e�@�Mͼ�����#��fC�l���b�E��gn�l#)W�`�t!�P�#����۶pVN��xF����xW�i\��nw�r$�"�-�� ���&����P*�����}�|u�����R�Շ(oj��#���R���`���� �v쪄�HﯹA�"���N�A�q���;��ss�G/��e%���)Ѧ�L�k~�����������q%/�Ϭ�j�!�?�������鍔�_�!��d�ż���B��*'FH�ģFѼ�A�l&�%�b�=�������/m	NN߽D4W�]yM�������z��R�ַL��5�<E�E�}	q��w
i��ٶ�!��r'��k����H+�|�v��Ň��#=j����ݿ�j�(׆9��i)�m�PSW}]���X��\��4�}fK�1������I�4�(%���&����JG�2H����?}x����m%��<�����%�3�r��Wwx?ُ0��N�.H�Z*�yH�a�<����)�X��!q�Y�i/�"S���@�8��K�񔋢U�����/�H�?KZ
��)��ڜ)�sHg��qH�e.[�q������F넨8�����������������_�K��"�O�d�VvR�>-��J��vP�����P�~�ˁ	�B�i�eh�ǶxiB<�V�5���מ;�
�J��b<�ԬVE,t�\�`��i75rl���� +CXMG���)��~YSX5-��a���M�)�f߫��q��hJv�9p�K�!k�1\��iO�Z�O�r�n�N�(�l�3./*�
� zWPm�:R�f} ��&JfT�й#=�F�z��:�lC&흵?�e��5}O�UCJ5��R�i��_#�x_��Ì̻.�~r�e��u�5�J<��&�m^Cf�<�m�����WI�'�����Ct�0��G�Go�ٳ�U�R!�斣t.N�D��MIy�%W`�����r�0ٷ.�wճ�����Q^F����7���ڨ�ſY�¯����tz9e;�^���%�hf�[�b�K��`�J�k��į�f[�^�t�ERf���i�+���j�S����
��*-��9�]m�9/��y��v�GI���R�[h�A�*3Eȩu<���F��d�$��DX���"䣙OK`�5;|g��F{��L�p��}M]pDo������85�w��a�	�,�F"l~%�&�k[N�e䛹tE����	��6�h���l���Wx:�Lc���	9����+G���@�Q��+�����*�L��H�/9�ٱ�b�gs�����*(*��L:�r9�����������w���_�<vϩ�L�_�m�?���eE�{z�c�������s��B��
F�}�����ݜ��[,��&)9d���M����z�.Yg������*�;�F�;&��Ɏ��d�bH�-1���͌�U���Y��HQU��J/ �_xǾ����	�@�A� �V�X�ԯ����W�E��)� _)�=��R��^NϽ���0z��=�4Kɭ�>	"��g(��K�^������,�2p8��~xŷ�qۥ��%�*��x�E�18�${\y�
Kϸ�N��Q<�<����j)����O��Ʋ������0t0)N�授�pѿ�x_�ˉCP��%�\�=��������y �T���s��W���y�E��.��}���\/j�z�kzem���.�a�gS�V�?;>KnW<&9�y���M&3Q��҅�lmCg����b[�<ӓ<u��ZX��!�%�E=��GP�'�����
�às��y/�߇��dII�4�I�"��
{�k�#��<�W�����|%'��Jo���y<|�LٶhFzdt���JӢA�[ǋ.&g)g��Z!Sf��8���)��ec�0Q��B���"�`��ȗ/[��ao�J:|���vBج���=� "WF����?���[3��p1M]�)��Ud���R<�����k����m0��ė�S	�Dp�8�ĄeQI�U�Ӭ��hR�D�hSz�FCf����Pp멮C'Fq+����W��/���>##��C����
�&5ZC�[(�R-�{�#����h��N���t)�����$5ϵm0n\��e��4~��=E4�{	&+*b�"Q\��36҂���r=�/ڝ_5���~e�vc�y�U�����f�;UR�*�@����Gw"���"ٌ^m9�m�b�p]ScꤨX�9�~mS�8!E�n<�� ��|���]�h��(�ǫ��xw�����K�`	:1��QZސӀj�����V��X�)h��i]<�#75�@�M�G"Ÿ�k6"��p)��M�"�C�цmW��婕���d1aw���+r���أr0i�׋ֳ�Y�d��D�f������u.����'G�hX�?0vM�.C�ޠG;D��5Ĩ��S��U���w0����8��Pj`�m�	����H�l~��V�8�xjz+4�G��2
�~ab��*�b�!*'�Ai�R����D#��C%�o�ͻ� <ߖ�<�#��?��K�i���v�-Aѵ�W��h�]K����7rL�
X,T�+�C�	���-X�G-�M[��m -�-�F�S�`�./[2'�Xʞ%�ec_LA|�N���!_��"�3)���#�����;��R���yI����"�y�H=��((��!|�k�h�����hf�!��zΈ�!a�����'r)�ְ���������Q#�,����q�A
���Σ�qu���b���5/I�!z�#<�󡑼t������{��4�~V��͈���f��M�Ӫ�3!s[��4��d�*���c� �{�t c�d����I��0��ͼ�0M��f�%�\s7f7�^az�8SBm�;��_��^��� ���w�Ƣ���Q��`�C,d�ď��J3��O8���<�$�wuU,���'Ѥ��2ƴ��
��h���j�}��|���S��M�I#�T��qL�٪8B�i(6=�q��m��6�����cs
�\��I���I�0�;��Y�� @+�<Ǉ!�_gc=<<+�^,R�<�
�^r�<)�SO�����F���*s0�~�H�i6p_�¬�) ۜ�)��Òp�̏�R� #5����ȟ���X�"�c(\ʍ�y�)��,�wo�^e�R��.~��GP�G��D!g��D���7L4r%YT=��?�������1��g�Ⱦ?_3ҭ�8ά��|,�AYު?�'����_�ޮU��HB�fM·zO��Om�_�k��d	�	�c���lXm� J(lL�X?V�)�ϕ�[P�m�2���,�,2錴$y�A�Հ���z]�i�'=����):��CV�}9�ħn�j��t�Y��-*=]��.Ik	���'�.jH�6sO�Zl/��؎y�}�`YD��h�����?����B��"e����(����7G,	�*[r�"���)�M��w��+�F���L�/���32ܦ{��v=��Z���7_�Y��o'Q�����s�sT��������'ǵ�R�j��1Xp5ʏ[&r�}��W���y�լĘZd�G�Bqo�qo_����Ĕ�E�j�b�ᢋ�aN�ms�Dn!O�����*��"��c�h�ri5KWc� P�>R�@ɸ���z#!�Ur��Y����'R�27S�N�<�������Z��`��=-�H��#(wQ�3u�d������N�6i'�3��N=�j��bK��5�2��zy�n^R��\�5�:_��͛�u|�^A���_�|��Q#Me�A�M��3���	f�����M"kt�:V ^�)S\Z�����Ts�K�b�K��5q�$r�`��������gih��ͥ׎��y��7n�͇��D�R�/��fP`$c�bkҗ�$ tNE��T�˝��{����{����Ui�;��iкjScڔz���@M5���9�~���yJgI'����T�zS��(��S/L�O.냯_���C�Ш�8 6C;�
�`S��M�3=���Ƅ��x+a��$���v�`������$>���f�
W�����Q�7'�7�$n��V���,�tyyŏ�s��
aDP�]o���>9�6X?_�9��.Mɸ�}v�O�#9�lطD�tLhT��?����WR� 	��E�[�H���n�Or�00+�u�@����a_�쟲� .eA���"�~�LwA�:��t�D��#���9��t��}`��}d�����||\J�^�7�Y}-��ëVE$�fj�h���'P��V%f�/��ͥ��3C�\� [��y3�>9��mQ�8�S#�
1;ɅNL����xj���*p҃�P�Ѝ��Oys���O��  ��:-��.�M�@���4� w�ć��*�M����nW�� ו�j|t�ɿUȣ���>��Z����'0��mq�Wn��/����÷B'���W���f(*Z��`΢'�'���sȏ�\�j�G�#7µ͈�
���g>˺
�QL5��?��$n��� �2�՟�>&#! k<$BU���{f}!5��E!��j�����zq��}!�?V��n⬓����#�A�����#���ݳZ�o��QRY8/�|,-vm�^���Q�G2�������W���¹�.�G(T��鎬T�T�$r���Ҫ�G5\Dƈ���Y�<�s��xr}O^�>�QC]٩uɄ�[9��#��eGב��*#�1�z�i(L�d/��Q�G��a���[v�0�oz���'
�1�iuC*b�`�_��K���GtB6|��sw��(N���\��L�6�{�Tg n�0f��|,��F��G��Y��/Cr��"6?6�ء�zƸ���c$�7�wp�i�;�;S	T�$S׳o=�]s�*�R#G�2'KV��<į�m �![P�|hS"cMJ��e�6b&4��Ǚ$�tB���|��@��AJ��⧵��փ��ʆJа�j��#�,�r��]��
�����y����'�б��?izQ W����js���VO_�4�E$�D�һ���%�G|u��eUo�z�t �����H�>�e�q��fA�����+����{�ύ�G��5i��wEx���=��r�J|s�aQ_	�<���R|m����9%�Ƞ^C]�3``�X��tV%wL���K�Ok���-���*���l�S8�|�\�1W��#�U�C1��.;�R�ɠ��6�J�f�ms�W6z����h����;�.�ڊs�����R�7�w��̘�A�( G�����U�rS:�|��Syw]xX�P��:�T�ژ�)j����=��Ĝ�*�bq�:�n�a�R�\�!�r��:1��)����D:}�:�>}L�j�U
@Q��U+�����`�Th�H2�ZhP�%�23(∾�AC��/�b�k`?��ƣ��	6 ��ߟ&3"T�!iԿ"^�?�_��؈�KM-���a���8�w�p�t+T(!�Te�}�Q[غi�a[@���s��w��^ެs��^^ь�s�cV�./As�*��kC% ���^Yd������Ve��6�V���׍��;�	�{��j�������
��P4I?��_���Ҕ=�:������/�l�l�g��2�eT�u�e���<D�3�� ��_�/��f3�dq̹U��\.?C�������ݤ�;*��Ε��̜m���mX�NV#@F�u�Rnp`*�I�~qB��T`���}@&j2`�����,c��	0'Vhl԰U0�l�3��X)��{�\Z05�"*-0�8�ϟZ����]����LoAh(L�)?���-Ǔ���rM�bp�(��Ptr���,d_�s�#�Y~iY�{�oǿ�9j)֐�����0-��c��V]�y��4���,�LF�t�|��j=M�ƌ�"��X| Rv������e"K:���c����'�z,�"���H��6�M;Lx�z�V��w��2֜H �H�17�}6��S�-�e����"9h��4�֍`��~���h��62y���`|R��Ef���*`I7�6r�g�X��U��Kݨ�߱=^9ކ���Y����/�����1fG��5M�ʬ�u�1"��#�2��VʟFܯ
>���5|>Q�b���r|�Zw�����{Q�@��Ƞ�������?��O��x�~K�J������תI��H��4�`z����/��β�zH���m�\s��[�O�0�)���$�A�*�7�pZȉ6W�kIX-[5nȎhvg�4Z`g����9���It��3�L8�1����e��)\���$�/BÖR}?�+u�ȹ�H��B��r��Ǫ1A����G�%>��
��\5Y<�p��ܲ-���J��}2iR�uT����#x�+E�ѭrꭷ���O{<n�r�o-��\ja�jy���턧�y�YV������/^K�B����Wt����ȒU.�4൪�pa�Vy#���z���D���~Tx�*��h����t�c�$�}��br �63��IsE��� j�-�o��h+���M���u�Cҵ��h]�X�;���N��vq�ý�7s%!	����p��&*c�<�;���3Ҍ<�nç���̆��
^រ�@ q	#���}�
�agc0�o�H�Z<(L*�8薆x�.\{±�	<�����;�"t>R!�BO����D�t��//���`=Ї�b��Ϊ��&�.4�/��	!i����M�#��8���3d}}��A7�iƑ"�|����5;�@�",9��}�q؋�~�ʷ� �6_w���������Gi>}�X�:+}���%zg2]���f�
B��('z���5	N`��f̩�Yqs��Ƿ��0��4t�n�m����>;�W��a.U�u��-L��ea[�Q�Vk���m[����~G�CwyT}*��`�8{~�Rɣ��,��Q���o�ꁘrY�,�op��`�5��l��Y�9NZӘC;,:ȋ����[4�٦�R��@V���:[��KO��Fb��)��+�z�5�&����M:f8���*���N FbX��A��1��/�P��32<�����e�}��I͑l0��%����;]du �q[��]ZX�%�	�z%���;m��gz�d<,�#������>��&�5<lP�PKN��=hg%�!���|N���GAO��f�e��ҙ}��N����n�|-
��|��)���6��s�,w�0�n�,p��)�6\ť�a�l�䧍����4h��/�A�gN��sE���׃�-y��Q��L�:N�>��m�X�/Q&xʋ�K.�OC8���ԧs�3��ȰS&��Ӑ.�Q:�����ƕ>�Z�,�:���a9ORQ�-O��sh��?=(DH��5�c���iq��"w��fY�QygE�X����r�jU0�L�}�Hؠ����GImx(ӳwVj�y{�m7�plPa�v���&1OZ�vs@�	9=ɨ�c�]��4���n�Փ �BOӎ:�r+�gR�٘Kd'+y07�x������jڝ�'�]�*��z��j\՝X��r���z`�l�Qj0�'����q���(g�bRl��e�c�LTs��#O��xk�9����U=A���`*vsIM�2ɿV�G�I�vm��r_k��@�Bj�&g2�����ʐ�D��z���z�`���
��.�]bi�$�wr_��=sx��NY�0���	��B�X�_h�p��*|Á����ެ��Dx�ȥ�&�0��R��}F�ӈ�gBvZA��{���ySV� ��\Vl9D�д�.�b�ڌcɕ�>��^l�0��D-)LBۭ��j�Uy��,�"5<^�m��؍���UN��tԕ���ؤ��ħ�[s�z�H�g#��y#����>;��,���֩�B:	��i�5�	�O�k;�w�!�q� �:I��I�|i��Hi1�n=��`J�S<����ti6T��C����O��pӕui�5�Ϝv���)Sٷ��߅[���}�nI,��IQc����H����vz��q�%۝9q���u��Y��ݿr��%���&;�v�����CJ/��k�tL|��U�-BBT53m����F%��p�<�<o�Uj���?�:����% �T3�ܖ	"#i�i���G؟����KC A�����7Љ%q
��vn�������S���'��L�;�	�jO�z�	�Aʾ��!��N��`��.*K(F�����C���U�׌���#J����rbb�
��8��{*o�yϼ��fR�1���?�Ρ%�=��dN.3����F,b�a
�hۆgsb̦@�eD*�^��g=�ى���(JY(�*�)��b�Ւ$�� TW��.>$Yv������-b2����A�9���$�B��Қ�]�0m7�U\~A��|�nI�G��:J|�R*��&�Ƹ��NX`���yv��� ]�?��A��<p�f=��H�:p[DpY빤��ؘhXs�@^R��v�}��ն9Fi0�"G�.�*&f�54L�.�G�j��4p)�^���6�{S��9�O�)"������[��������܆W�,��̜���«��mo�|�)V�BNHh��68����|v@:��%5x�Nr�JߕьG4��.�z�������j0�4:�`W�����֢�]�դ���OY�0�zw���5[=��,��ք����� {�!��c�l]9u�K=D�G�D���t���F���v���r8r�F�9�����0<�1,'ڏQ`��������)ZG4=��k���g�q���؎�����������}Ê�����0QT��Y^?���Zs��+����m������o��9��]�m��v2���H+K��5�?QЪ�3,��l���wQ=�Z����P?BI���'���#e�_A�q8��b�p�O������|ֈ���\��O�8*�W�:*P��9l�j���=bT1�7Tu�ԥs�U�M����g=}GaV�׸c���<]�H!����i�	i�PKͣʟ�*���u*T�)C�s*|�{>�'�o�un;��sp"���G,�eK��JK���[�~�R���ղ@�I��v����p�F���?��yw�ԁtg\?�4'
���f:}Ӱ�ʜ����W�Z�Q\"����tQ��;Z�G&�?)�E�X���8z�d�ևjg���#`�V�|����DȢGWQ�NL�M=F��Y�M��Qt���
�dw	y�]S�^��OSgft8�c>zϋ0M��R��w@T�����D���o�45%��ƌ��XWv'd�*��I�<�~�K�ʕ�_���?��?�w��{�Ą�������/C��[^B`��l� ���T=�
ۚL�/ S�����T�����	��R~�a��*T�5!SԔ����Nq��K��P��ҎVFl���'jZ(\���ҭ3��"�ۜn��1�X�4)��+ɖ��{���C���~3���2D��o�W�'�9Z��N����ޑ�|+��M���RK�7%H�9r�|TT�X�n�U����|�s�AV�L�Ä���/�I(�
����רxZ
_�Z�%:�k8%0�.4t�^s��\sG�e��+-7�=��v����ҷњ���d���.d;����G$������ү!����Г��;U��s|g=t2UłI�^Uݘ^�3�4:5G�"�]�/*�6�Nv�tL{	]���t�ڕ7mD8pU����p�'^ |���f��CU�,��P�w�S�E/�E�^��ǯ�,F08F;�܅��I(���^�L�Z$p�Q�U��.�gk�.��Ǔ�����'V��x�Q�'R�2����e�W���=g}��?'s�o �R*bs�>��YDA	��߉��*C(�_QʕF�dy�)�9��R��V��m��bM8�љo��C�����4H��@�q�e��	�#Phi�ϰ/���� �-�4?H����z_��Ag ��Kb�m�a%b�$WI��ŏ�n~|�6'�ENA���%�E��/�D��=�w�$�}C=�}�����������ܪ�wn��\;������2�ٛ�-�u_�oZ����+V�~sO��c�}���G�ӛ�L{�ѵ]���vv=�UU�2�����ћ?�p%����.�@n,�"�.8*�R�#Xkrs^'�b�
�����T]�.Z��1�v!�d����F>��c?��B�,��TF�������&-�S`g�������g��tn�k��Y��&��]4#��`�W`��!@�Ў�������D2s#P]��DB(~#�
~cG���< �,�Z�r8�*��IW��Q�h=H  M}��z4A�SM�l�Pm}��������	{�4�=&û�
˲�U���[K�W��6B�w`�� /H�Y�3x��o��w�U��,q��Ej���Y/�f�fj�uy1�6�]y#M�>���y�K�+ ��ݵm��q�1��x�o�kL��h�d���k�M43.���p�6����{�ߩb"�]@9��lT� j��%Z?3}7s��.��7u����)L���ZG'�#� 7�on��	1~�&S����P�^B��Bfa��Y��YiUk����y�^k��I�#;]��!Y��Gk��I=&��dͼ�������Fc�rC17��u�&������B-vn�#��Q����
 �᫻ !� 3�$�:� g�_�bv�a����*Q��E'��i��;٥ɕ����%hL�p �׀����3U$��-7J����l�^7��r���w&x�SZ�.�c���qCU�1]
����܎�r]`��$:��؞@�����Z4�J��dln�G%�	,&������n�}ݣJ(C's��9�^�^�b��	��kB̜v�k�M���默Z�ȐE��j���4��m���o�D�ܬ�z���ۥ��?�O_:'S�����5���ٲul�!��C�vA0�;��Y���U�h��<���y�'2����?�>���i���b;�� �#u�r�t@��R\@�w���i�t��O�����w���������	l� �8��/�}=C1�ҥ"Nl�7�x��h�J�p���i�K�_5B��#c�;�A�g��2��DM@����$1E�%7Ar�h09��Q��h>��U�IS�k�^�������'�"7.b����*��+/�e����On[�j�&��V<��X�.�}��L��_CA¦�q6b�B)@<����"v��j�ٗ��%poa�w���D$��VL�V��A�4'T����-,���^�1�#���?ܫ�&2Mx�������P�Ww<����uZ��c�f����D�"w�8BF��
����׫Z��w��*r�j�9���no��5`�_�����+�_��\9���7�u�_O��wS�B��&I���F�^��5Qp�~�s��]�"�<B�Dތ��b|�IA�3����3�t׎{-[P��o�yxi�`InK�pB�@.Y��#���*�������ޜ=�MS_E�F�� �ȶ���Fү�V�g���%��.��( q>���tB7X�!�|*��]ז��ٞ�X:��v�5�z�����-}�0�R�|�D\��R3��N�N`�~� eo�-L�iyN,���]ҙ9h�p��=Y������b�v8/2�c�
I�h|�����%��}vP�5���>�7��p�r
yn')v%�� z/ibN�/�}���Q�8��8>��!Ȍ.�2Rf�3c��:�0JZ�o�ͬ�XxV[�F�!J�!PD�\��	n��I�W�)��jQ�,���A_����]�vvUP`��m���A�9�Y�P�TZ����u�46��4�K����ZjY��Fҏ��-�y��o�`Υ�9�l˘���yB"	�w�+�� $�7@���ڴG���с��EB��2|D>>��cr\�|�]#�=�HX�E~GE�Xf�P=n#��(�l�#��d�B3^����q�i�\�w�K0V��������� :q.��V捾�h�H���<��0�7�G5N�;u����=Z��M�W#;�����gPÙ3/���(rZ+�7���VaT����S�ִ�~՛���=eL�ڰn�ل��z��50�د�|I���|4����:P?i9,�1YR�i�;-J�R�u��F�p|q$D�Y�Γ��ɀ�C�U�>����|�A��ˈ�����r�P���~�V����/jj���4F`O�����f�޸�3C;d�9�ʂ�/���8ڡ�D;��"6`*v�fA�W�@�<�� �ۢ�����$�VV��]��-��D(��R�ڴB@c��G*��IŜ^&�Ӄ���I����́�썸�%ˁ�k�I< ʃe>e�����7�����ԑ�m�܁5��.���5'7�<|�nۭlY/X��0��Oq?��k��B�%i�Z�88%�ޣR0��8��<%�'䷸I؀���>�gHg��T���&�N�䶎���8}pĉ3ן���R�4@��D9�����OJ�Z��j�����E��k��p)�]IT l��]�� %�S�X���l��f�y[}C~�H�nY��ub(��ۀl�`�v���
w)`|A�К7K/�]<�g�O��<'��	[@FdѲu��r��'����5i����Z���aV��G^�({�^.U�m,��be�8?b(����A�)�F��̯�[��l���uƲJ��^.OR��	ؼ��y�%u��J�ݿ�4�a�<@���U�������o�=���)��d;�^Ù��[�QZ)��ZPMy��.�n����ة��c:~�uXJBj*Ac�54��
H������r{`}Ag�2���a� .2a�ОmQw��ӫ�up����+j�v��S��
N'�Z��r�IN箼��!xb:U�m��l��w���G
3�]mD b����5k�a�{��ě�辞�����&��%��8/+��͹Bԝ�;�[fl�����Q�Z�z�n<h"�9������]�o�ɭN�&|6s
o�ᆒhеT��C�����sE���L��D;"�r ����%�sʥg�>�X:	�&��S�mM����n�e	X{������|�]]>A�I�#�h2���8\���>��ox��'�IHr���.ͷ�9T7w����m�1	|����i$E����!���U��«��=d.�m=}Tf۸̂�����ǧ�:6���SZY�����$���.�s�`�O�+�T[䨸��Ӈok�+����p� �&��'�)_)B�9�w�|݆LL-��H�9 ���u�T�r폰w�A�/��n<�� U����<SfUt;�̗�#f�9s9W����db��c�Dk�
A����A�z�-BS�6�vWNa��	�T4I�J)S��j,ƚ����i;k�-x�o����a�8��q�h6v�A��C�~�f���mBd�5R���{��أ	�_���_~w��Gj ³�c�,����o��Y3]N��z��9��Y�2�f���� ��{\���r�TB�����j9�޿�����r�`�+Ƹ�m�����/�~�_�]Г�S��><CM�Ϗ� �<�i�<�Wa��
�� �����}`��ꗬ�sY��YX;�,�52Wb�h���*�����+��3��0��l�0��"~�B=`��s�:� /'B�]pmٳ��g�X\OP�)�l�����i�*�V�����V��I��ma����&�z�O?