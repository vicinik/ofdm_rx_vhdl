��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P����3�T'N%w��d!Q1%�7̬�ONMς+���u�'" ��)�4�.��R��L�0*��vX���Y��EY�U�R ة`����Iʘ{�Y*�b>����4�*}y�:$��i��-7��C�I�QPdN���� m��3��=K!�3 2��H�l�8F|��w����5�i؎���"�^�EX���m!�W����Z�:��:�=8%��@���h"P+������J��<d��	���J~�-��I���l�5{����Wa�W���T���w�})G�2H�p��z;��-��D|���z83�8�,�
����:��A�|���}5�;�0)9��K};e�]H��Bjp�{l/x]�)������zlY�6��Ɩ3c?��-�����KV��~W��w| �(�l=�
�"�wD�	��zq��1�����\�'�I���������FHH���N�W}X#kn�8vX0�>�K��69��k��u�1������'/ )2=PT~-@[1(^I�G,�5b�D�Q6s�I�����gl�w�AK�G|�P1�B��v�x$����s�F�0X�M'E�������d�xR�/�����~�{b�À�f5�"R�p�X����Y���ˀ�uNa��Qmt�|��r[t rw��	����+�r��Z�q���"��v�����l�h�d�`>:���m>m�z|��M�g6|����~W%� fB���}�ڲƂ#���� �V+}�7ׂ۩3 �*��%���=;N�Ӫ<���e{��� �����u��!�)+G�g�����_�P�{�.��B��֏W]K���D���Ҙ�v�{� �+���9�o�% ��ֻ2<-{Eg�^c���n�҄�?1N��Ð�m�b�d�֟V��˹g8�����l�$M�f"�(M�W���p�̕���p�>����zB?��k=ǸXo.���������?��� by\��9K�]�o�wd��,�i��D����a�0W�&y��� ����<X�w��]}�Q�Y`�]M����hr��mf� 4B����@�ë6��
B��׌%����x���]h�����)C/�_AS7�۞IY��;9�o�Izw�a���@��]�1�5j`���_�h$���у#N��̓97^p������_<� �n����.$���8��V���\>6�}��e;
���t���$*������^G�I?,�஋�8��}v���;�!��\8�Zz;w�"��a�a�2~C`�_���!Ӗ�5�Q��]�:���&�{���<�-�98x�)A�10���@�/P��zX
۠�E���Hh�~c�>�]Ǽd���5&m2�t�&�FǸ�\>X[>�=����(@U��̧ƞ���plZld4x�6��ң������	��cv�}[,k�G9y���#<��r1<��ZC<\�����)���V����'�QC>S����ޮ1��`�*�>�bH*��|��:���\`k�t��D~C ��5��@�;᝜���.a�(�Z��n���)3�%�#
;6}r���`��՝u����9�Y�C�����7�j�^'KJP_D]��� ��(O�(!
�@�Z�?NOn/s{�]�20_����_:(8N�/j�5|�a'�eձ�2�K��d�onhýj�
�H`�R
�i:q�������^���_��ǵd��w��;lr���0<pe}�p���%$Ne�,�1��}��Yt���������Ѡ�6$��H�J%���`�8�=ˀq��ޱ������]=:�Ui;QӬO&��՜ȑNzTV��!&�d�$�r�ؤMI6:ɶx������r|�ѸV�"ߒ�S.�Ĳ��uw(2L�?��m���lt�˦� �2y� ���8�׸ޥ`����5������$XŸM�Ŷi���)I��h�^��ܧgݽ��>7���l���Z��[��׫�0����j�7��R>5�
Ԥ��fo��>�Ѐc%��[U9�7�'sLeE��ɻ�&1�)�AQd�I�=�g��G�vFi�Ί���uA;�N���kHO�=�C n���������"��~Ǝ�y����Q^v�Mj�X.o����9�k���.H��M�c�P���ղpU��K��)b&��};����^���֋hm�6 lӽ=�N�_)M	x�b'���xAl��Op��q2(5҂�ܰ�'�rPa����!��s�O��c�k #�jm�	���1x{�*���AԈmB*!wt��A
3��h+�A|a�X��*��f)ٿ���z���a��7���*�9W��]b�zn3���
��k���y�s+&6*����m�Kݘd�HH�]�!| 
`*k���[���g$�c����-�k�;E��h	`ؓ�i�iz�CU)�<�v�:���:�#
�x�4C�,[��(I�E��I�!מ �!���l�t����tqE�ȐlN	���U�=b�\q�Q<O��B����i=�(�>�u���vqW���dS���>,�ӄ�R�=,[t��H�޵i����N�F��n@2�_��2!N��;)�ӈ(c�0��WϪS�}.d�7�z��I�?��v��[�D�/bR��N��wx*�	l�?<j(�eR�	E@4�yw��Km�bzy�W���=���պ�(Ƹ�;�P��q2��=
$g�)n�8�h��Jxnۯ�r�/� ���{l���@��p���9���G��2�E�.��E�I1����ؾ*��1��I��n���E���y}u!�;)��z������O�;'12<���K�n���>�E�N�{�4��YI�-�8M�Կ�O����;�P�j�<�ҹ�"�n����!{���i��&?S�4�o�Fq^�
�C�X����)J%�zc�XO��Ɗ�=p�aC��q��J��C6�p���)S�A�=#��
\ mWS��G.��3&x���H�R��*�j�Dl�}� l����sUH����lY�8��^y4Ӛ�xH��"�7�oJ3�]�}l��E?Jf� �����03Q֑�V2\�5O�[ 9��nUR��[>�~٪O��!��`(X�f��ٶ��c������D���u��*���cz?�y�T'�k���/�,��%l�'ʽc#
�����-�IԂ>�Vx� ?��\#���y�-�����>�~P�[���H�2;7��<5'&A4:02#G��(�K\���xءՠx�0�@A��>�'^,�w�&3�̼c��.$�
�힢��-Äo�H�a�p��dG�_c!#�>^�H����WF�!�8/L2��X9/;zT��(��8����)(,`�4�����!Ŝ3w�aq�����L%i�3�L��{n�2��q�,��R��{3�~$��6,�Ƚ���:X=&�[cng��ȕ��5tp����[�y���3	�Wf�i�j#v���Gs�����:���vy�1M��.��q6H�:���˿=���Br�8ϼ��oL���o ��D#�7"hЀz+Op��Y~I��Cʨӝ�c�&��D�����.����Eҟ�֮	����� ��]ʣNj+qG�.g0Y�z�.�Rp]���>�������8�E���h{��HNŷPg�R3��hq[4\�/UZ5�%o�7ҙ�etH1 �"��?��t�=�ĪtPQ��H_��P����jx3�5�ꂾ�+��dOz+���+��6I�c�7�1E������8�Ѓ���lLwG!�m�'6.�Mn<x���vJ�<�����G������˿%� o��l�D������<�Y-��@���quc� f/?{���RG��6�*�[XT"�{�a'����2��}0�[r���o�ZLy��;g�"�ĥ�A���j�Ⱦ���"�)ރ�p����;�JMWɩH`5ڹ@�<[�fq%�����[	��Խv�b	V��B���F�h}�H�)��oU�]hA���B����S�9o��?�����b��)��� %�'��_��7f�pR@���.|r����[���F|~�r@h'���-ǧ٨Mo����uW
D�����t����9��ݻ�6.��p@�@�W5�k���a 4R7��`Q��y���pR���s�+��<@se�����^<���'�>�Dk�S	GJF5��hnI$$��������K�%Tj��e�"��?�\�$�`��V��t�#�i{И�hZ7.��:o�>�_��J>��p���'姯�|^����SE�$�� pT;�b��7�]l���̩�O,]÷���-x��6e���L~G���+��)�����ڣ��UI��;([(��zE�}H0�{8�Cv^(�����}�ɰG�sA���ܶx�덱LWLb��c$9���f4E7u���6�봚�����u��	QD�eL�F!�*7�N��z�� ��mc�<��EJr�90��k6S�{f,�j��r�9�3Ʀ��4���qT_��wS���*
��f�E[�k�"T��\ز������z|-^�^�?�g���_�%�O!ؗ��PRB4i��7��\{R�n��iv==�m��r��T�ާ��vs�����iq�L��,^�L�[�%��p@\��"�0I�|ks��bq��-�颰u�p�T���
O�*D3B5=}��a���FPL��bb�_� 
Ǖl��a��;�]�4ۈ�j�2O��5�Z��y=���	EMT�GEnX�|hѢ�l��� ��c�	>]8�"Q�=�1z���(�l-y�\ӄ?�:��
�Iд�9P0�t�A�.�MZ̽qs $T�7�>f��}#[�	,YW��	�a׹��JlFf�x��n�~�Z�n�{"cgm��fdWL�_g�*�g�D���xL��/�6��P����.��ȑw�L���(	$Cܙ$��!�����B�����ߎ�K^�L�!:N��3RGx(��\�E��˕~co�bݾv$<�&U1��EB��c: �v��� 6��͕�������5�y_>��G��b�+T@3�����u!��z=��Uc�MQ��H0��&5�����,w�<���]f��uMQq�5�Z��mr��cE��X����M��CA+�b�9�+*��@��djh��4��@|�0���;�M"�L<_�Q[z6���f�=+;�����՛S4)���9���j^s��-�&G\5�J���ӱP�I�p��NM�>x�v�|3L�N�\_GinK;�a�;4�ѭ@`�!�c�i&��D����Ȣ	�AikY� L�)z��έ�>�]�ǽM솰f�&R�!5��V
���u�0$E�@F�O���Ev=[`uIN,�@������av��k��n�0Q���։��a��L���g�Q��:�K�|����36�3��Du�,n3���莘L?V�ģ#[{� ��="΋�����Ҭ��/,Ӎp�EI�����ub��6�{'Њ�)g��O�������V����+�A|�U
M]�jX,'NϞt��8#��j��%�H<-�>�L���Q�hۄ������s�Ԇ���%ԩ0E�M���1}\�K����O��nr��@j`�4`�6��������M�� \ҳ����Vr$�_c���,�vpg�-	���x���,���8��d���֭�b��t�J�Ð��O��Ԙ�C�������y�β����h��|�i������w�����c1��O��%��z�oz�DI|Y�������6%����v?u�?���޲>��=h�_?�g��fM�N�%x)�q��>�Y�z�JQPM�J�ܺ$QPp~,�'<�f�SZU7Nc&�;���D�h^�`}�7]_n���|T�����t�t���v�7��>�����=r��\�i��$.�����90��F��$��1��G;+�o�ڝ�D�s�}4^QD�7�>�PI*���ˏ:nYS~u��|�^�u�#���)i����c��LV:
��k0�~�=MT��Q� �0*�핅J@&Y*��l�@��\�:����n���?,f���Jk-wu�Mn&�T��u�{,iO�'r��C�`k�'h��d�	XF�<h�8������y7ogq�,�6�A!���=57k�����m������]	" hRUhfD�`�Gܝ���C&*#�����o���t�'�zQe\p4Y;#F'N��H���Ѽ$����I��>����N)P5R2�x��.`Dwk��Q0�l^��7���-K�Ԑ��[�cڞ.��c�w���9W:p�V|�|��[sY�Y�R7�}lxL{	K�b�7u�2�-:��&Ŋ��ht;���u���M��7����)�Ny�ܞ�Q(<g�Cp�>璘� Za��"<.
������f��~�&q$���=�	�`?�1�̯����Mw�M��;�6��o�n4q��{���z*�C��K����X����t|�8�4̸$�(<�����)<�[�ܚ�ȽFqͯzڎ���T��Z4Ib��S��g����&^10L(l
�vq`
Q�e���Wɦ�a`#�EI��@�ȵ�ͭ+�0���A�h��PR�k{��j4ҙ{��D��1�4�x�hxs����J�T�.�y)J-i:x܈�N)��F�*��H�4��]�{"α�������[�'4v�EOw�����vd��b�g/s/�`��[mkqP�b9�K��ή3'?�*��s"���`���"�+�oE��u��n*7�-}<�h�ȸ#�3r�}��.��������O�zj���!�Ί�>�BɃ�v�L�֔�F�3���tU<�G��0`rڌ�����O,�&_�ڍ,���!jT~���:{����֖��a���6h:ȳ��j��c/�`̢����u'g�-�C���=$?�8}�ȡ������jI�0��F��mp�<�jw�&�4G��i�<%C��r�>	h�@�Q:P�)T5�VׄȎ��t�}�'D��Z�-�+��?�&�0�����)P���/ԓ�u!���S���?ćICH�B�����gCnۋӚOj��z5�,ޕ��x@�����zC�Xb$&�)���e�
�Cs! ��7���̦�/m�����3C��po�1s�0M��AV'N����φoD=0_�~8M�x�b�k��C�@����ݰzy�����Z�IL!'�rС��Ͻ�]�	qR��7�"����rIB�d���(�F����L3����2-����b���}$���~�֘]�y&�@*k��uN�링}S�멿�}�c�(�1.x�����Z�H[C�[c?@59�^痎|�$cU�35�sP�'8'u�ct�#
��k:�Rk�)�~N��g��ʩ�f[���Y�z�A��^��.>�B뿅�5��ܙiK�"��U0��ԓ��o�wUB�Y.����=o'�u���-��=Qt�bD���	/S%���Y�!��I�2�~_z���7NS����3��\�m½5��$0Uğ�,Ȇp��q�x{&�o[*z꿵YU2�ѱr�ee�tCK��~U9�>��f�l��F���@��w������*'����ɤ?�߬1��lo�&�vn3d�in���Wr�m�ɉ���&A �=�� 4��6�]=������.1�q�<��54�Հ�_H�l���������#��8TG�^?4�M�d�}*�W�9���$*g�x�6����T-�W$H�� ��- �B��S�]�@�N���㿕��Z��id�z#?�%
i}�"}1w��.�M:H��[mZ��" ;���-�Ѫ��X�����M-bχ��Y.L�V�x�;�v�a5Yc���q�4�9�w�ɴ�wզ�b�Gq�֦�q������p��m�5�54P�,B=�m�H���U���۩%��ٌ&m���)L�ҝU�4c�mܢ\_p�ê��,�/$X'�<r��z��KL࠭�m���h���Fa�h.��f������ւ�Ӭ)7<���ڃ�F�G!DIURa|y.E@��G1;Uއ�U�&lS9(n�T�Q`0疫�u�=��R�p�(����Y�S�Y���N=��C�?�4�Џ��`]f^�X����i/�3�^���`^�f���"j=N�����"^ܳ�〮��~��N��^:�,3�s��p+I��Ǣ�3Y��!����4!)-�NF�D���m���8� {��3R��D��2�e�uw��2]�L����0y:�?�'�޿�K��y��`1���i��o��[�
�d�XM����k�k�h�̓TUb$S�6�����A�섴Ên���e� !�H���h	���*g���:�ǆǙ��*�R.i�2_5���9U��O*2Vsp����\!���&ȻZ�裆��a |bw��{�o {T���UM��h#2ڿ(��{�!��=9q�7꨾�h�W��N��и�ʮ��q�{?m��=�5�;�/8ʊ�_�Фk�Ϯ��W�G6��� ��W�ii��w���xO�$�G�Z�M��� c4¡u��@�Wf�o��F,Imjw$��%�	�H?��@X׼�Z��N�0Imv�/y�N8���y��J`2��,��~�)�~�ֽ�b���u6�dt�xWLw)�&�� ��vO���R����uj��N�M[@��c3D�n�-�e���BLf���}d�h�����!4���
������(Í��R�S �����3xw��X��y����8<���q��W?�n-���-#���_�X፩3
�h.�=Z~��ay�=�N�jܡ��S�W���Ѓ�����	�0Ǫ�'L�:n��] V��8�#r��VDJ�N)���p�w����;�R�H�������8��m@��B�/�g~խH�h�t1R�i�:�i��Ҿ�O�ݗ���6{OO�gal���u{fLPg�1���lS(��<��B�y/i�4b�D5�>arl�c�m�+�&-0ʲ�yUpd	SB��z����CR0��T�q%08��r�*֟E���M E?��dn3��-��ٖ�Ѓ�Z���Gs�d��c�M��m�{��5tkr
1+�e06����S>��:����b�\�B�w��,&�`ת�I�]#�"���k8��G��`uk��p��I�>��W�j4��_�2��B7�r�r��<�Y�~�\�u~�i��E����`Ɖ�V�_y�&[�m��\�E�ࢵ���u�i����k�v�V���Гe6�%h����-�98���(3 ����Ӓe��n;�J��1�p�?�m4*�[�II"|x��+��."
Qo�~�ǜ����[n�b���ɀ�/�W.ǜk���t-��L�ga�R�Hel�>Bc�k�a��xڬM����Xd[I�2��vq�slC�Hhƴ��f<�Pѫ�S�:-�OI�uʹ�I�y��@�Uڮ��z^��z��b5)�
0NRk����Uk��#4>ZM����Z����Tb$���5� 6��Z��m�z	�B]��T�VqL�)F�D����]~����4�,@�7=�� {>U.�j2������d݆�(Y��_�W�_��z��� 45S^�	@5�	���M��~n�Є��G|\�s��(�iVF��̃���:��t�ͣ�!��I�˕HP��5�"AX��<�ڢ�L0$@~1�,�����6�B� 2�����R����nQ���}�a
rW�Ja'_��s_n�V�U<���Le�I�1Ȳ��9V�\�%�d_��am��>`�2+4�����ܡD9D����bl+��������ɱ�o�c��ֆ�jD'5��5r_Ca������~ty���kl�O�Y7��%CK�Yo@��Ғ^�6j�abY9`.�Aے������u���w���uZA�
�zh�	�}�(m���s������@��_�և#UI�5���@�ڕyʾ�G=