��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�#���[(W��4.�E��q��/��v)S�a��)G���U{���W-`u|Z�Ⅱl?���	P�sALf�h���0�����𖛰�}|l�w�O Ƨ5[��2_�@�UI;憙��Լʐ�b�:���P��^�^x*�݅[@���"Ŧ�x���������D���m��y�����?2�\m�P��S[��9���߰�q�lrt�RƤ�"�8$F��4�+3��Ff�dM��9=��e.�~����Z��#}Ԃ�����|�WИ-+%�
,��6�Y^*.�6B��4 .�bJ.X��~OWS��h��]M��mr�UO?�J;ajw�k_�B!B��*��]�l�<)�:%���!���{�z\�&Ln��`Bd4����ɢ!"&�Q��	�s�=��R��X�Zf㸝��1��";#������n��i��^>�����m���Gh�_l	f��>&[1l~�]����3��GN�|�P��J�y~�N�#�YO��]
h�R�3c����_͹��\�蹋�Z��4�q�=b�3S�
&l:�o7�T����ί�����d���s�$}myq=�g畣E �~I��/��L]��T�I�0!m�5;@$W�'�B�c��06Zv(�b�=��C͠�����3�k�� =g�g24 �"��)�Ֆ�c�e�J�Z�AO��c�[PR���W �u�L�-o�ʑG�����=������3��ӕft[�5��qU������9C����/ܜ]:�y_��-��ٞBʧ���g�� l�)�T7���9��v����tY�Ȯ ?�AP����Bs����C��\��ښ�04����
�_�aE���s�W�R��RA�<����<J���w���HSvt�:���&�J��=#�ʸ�c�7)<�:�h�b$���43��3|H� �Ǵ�S�s�uT���u{=��O��Η�kR�Q��0�-�V|�
�_����b��YrF���E�?�|�_$�V�	�n���h�ƃ��&�d԰���e���J���z�_��4�\&��W�N�L���O�.��k�~u��}�q�g|n�H�N���4PLI��c�G萾+��-M4��+�y_.������T��������O���������QT\P���DRo �|�����h�~d��ƕ��)8g��g��L.������PFԌ-�|�K�W�7h�UЁ�񑂣 s�)�~R��t1`�o[9ǋ��{U�L(���kA !]3�73pq��\U��!&������!۩�j4���"���������(�p�w�|�wiFP�q9��7{�߉^e�ZQw��&UĢ��"�fwTK��"�6-܈�늂<d@�%T�;n,ZVM��0v6����[����4���Q�=F�z��]�N�]:
t.�~�k����奡�S��z{L�w�΅����߭���`��E�q��F'���Ǐ~?��FDf�/�O��G����ŕ�1�Rס�P��s|0)@$�=GO��g��t�;�g�;� #M�������ͣ���*(f��oN�-�V�7�c���^r���P��)�~:E��L ���U��|@m~FC���Yy�a��b`��+���;�Q�d�sV������T8
��v�\A�QG�n�t<[?h�����&��:f���qg@�t��/����Pg�O�>����V��{�u.;B�g�eJfK�#�^R�]ƈ�������oG���H8����@�
y��Tח��M9�z�i'@�([�K�T3h�#��Q˙��ܥ�h���w���n��"�N�
=	�2�V(K���ξ��N����kE��ʩ* FbF�Zr�k� .:	� �\q83�V�'��>���#�� �8!v �(����^������ <Hb�$��������1p����J�Du��"�jgS��,�E�?�s����>
�	��Xk�cv�9K�>�m�������6Kd9��lg�a�j��s0��b�Ф�
�J*�V-T�Hl%n�BM���?�x�Blv'&�~��S��O:ꥇK9���j�������m��K�5LES�8D��y|�%t��=g�N����ݫt+Ϯ���B�� ��B`���\̝��M{Α�m�_�b����%��_I}Jg�`��m�iO�\�#�KѬ���@�{�Q��I̐�.�$(�Y�ջ�)�|BZJ�K{�_J���G��}�T�7~A<4�ĝ���ג�!r�w�^wS$~`��o9��=���Sf�� �L_������2-:cFW	��l�`��9&qQw_y�~�̢ӝ(\OUe��Qa+m��{��ȣfby8J�<T7 /���8֯�������U�	Wo���@���˟�Y���!�������>��X7���Ց���֩&�_��.���:���?WVw5��>�4DQ=�<!q��!���<5J駯�kH�t�z�(�;���LLq�9��7QU��	t��j�Ѧr�W7Խ�"B�]�_�"0��5/�����̷�
�j6'���	�C�Ȝ3��@�V����1;[0�i���m�>�~��8����V`h<5����g�2k&\vA�-�k<P|�Z)F�ʅ�[������T�1�kͱG�^p��P�z��$��x}*�ɒ$�����0�W`�TB݆W�c|�y���)���Y%R��T�j��`'C���#��q��<����?9&�h���͝�:���"Y��r�xz1k�<!zyC>��[�$���2���}�� �Ww%��~a��e�Ҽ;���oO��n
�m^��j��T�[�dd���n;ܯD�;��?s�<����=Ӗ�a��c���9���
^6Ά���BBDrP_���eH��McGT��[�aᇛ9��Z���ś�y$YT�J.F���ɮh�1�&����b�	��3��0Gf-~�H"�/9R����Iܧ��֮�<�fY��C��|��8��=�$m���_��P���n�ߓ�U���ڲ\=�]��+�
Uw�����t_��]��US�?:q=""\K��X����V��/�3����9���i|�2�>+x�zB�\
��%� �)��Ud�����+h�C �E�a�|���w~�^��U��>%���3B �1��:W���e0K�BQ���K6Ϝ����{�Bb��Vc���!�3�4{^Ǿ�{H[��L7�f�%r��?����!� A��o��+h��|�!��j5?h����ʮ����V��I�#���]D��>*Y���̙�r�����	�}+�m~����+4�t$ӷQGl&��.���N�4����K�%)�ds�N���[�e�.�@��%44ǬN�??lr��|>A�9����)BC��3r2x_.(�0�����)������m񿻰 �Qr�yT��w���R�k�h�Qϔ\���M��)�:�H�Cc-�O���d|�F��A��>�戓�������k�K�`-I]C�>)�b��3&��/y��(����T��1t"2�p�*����UD�ol�tu:c04z�a���3sp�4��k&������	�V����j���}ةNe��`ws
�҂������ykև�>� ������}J~�69���7��P2�䂊#Ցr�c�����|��������R�P����{�O�`d�.�v �t��E7_*W�W��в�&���{�fL��俿H΅�������n��{l���xMm�Q��8�0�6�@Ͽ2�*;ɓ��P�ӞF��1!/(������(������$���؀Jqr5�BP��~Y����焓�VR�ҟ������>Cî�&Hf�)�=�@����S��
�l~�8a�)�4 �}K��.PR+.f=_?R2�P̰Y�6.�K�Y�5v���
T˒m��a��VKhtYOC#��	�Z8Bjɳ�j'��H�$�X���*~@,v�)����S(Ճ�H_��"iK�{w���(�y��M
�Wz�|k�
�ö�<�Ah�[�����.���)oqԁ��,��/d��.#ةB��)�=I��͛D�B�m��	�\o;d�a���_a%�#WbՃ�v*<������_��eT����� Mh���ڪ�����l`!�Qɥo�Rb=}���]I���,�z�v��M���lrwAl%��\4�s��I�%t:+��{�t�pD�|Џx���Rr�����ɴ�i�;r�uM�HY��Suћ���\1���=iT��Ϧf]�����#+���D?ڰfu���Q_�Toi����\L��V���=N@���Tt$L���>�Z~����?�� �}���Z�^1���*k�� ���|�������pjr>�V=�����5@r�a�Z��>�݈'����Ё��'���<���:���	j��61�g�prE��MM�4c\���^OE T�>���0���J;*!�Nh��F���ԃ��}��/Y#��I���W)��]�|�,�5�,�^PօS:n��@��Ô1N/W�v4^��b� S4l�vo9�DL$)�^A-2�5��)��ɜ'��_|(��wD�o���i�Ii¤�-.Tr�1.���	�F��)wJ��pS0��P�:Q��#�����&5G�.!��o	��ܱ��@O�!�x�Z��GyЕl���G�n0|:����[쵰�qg�#������P�t���fpԱ76s�o����Y
9�1n �.l�`��.���.Fh6�Τ[M1�;T+v�U)��J���k���fJ�B��:kJ�my1�$6&��P
���)!Z��*KO��Z:i�$�Oc%!2��!
�a�E�c��j�\B	�^A�$��� ��s%����)�F2:Z1w\���Z.O1*��7��F��r���ut��U$��DA}&<Q�HݟYD���2M�X�ʇ���F���q�#V�����řCg?�� ǫUL�m}kZb`v[��zVh׀��*D�� m}��a�`7 �F
�)������P
�)�2I�p�͋y1^�c�@YR���/GMCާ����a~��a����8ժ>����|��z�0�d \���9�a��9�ȓC4��pӷ�(S��e�#���d�ĝ��6�S��e��G*�����q/J�[P�}����#��0ߐ�Qo�D9Ɠ�Yxy���n�~|��Eg���VH��yn���5$���-H�ĬS�*������W{wH{K��A��h0ʑ@k-��2)�B�^3Ta������E_rqgԪ�id�`�[C�ؿ-{.��D5fC)Ʒ�\�6����D!r��n%�h����v>��Ӽ0Z��<�?wq��ʦ��1K�Y*B�����O'����8���Q�D�uT��h�T�AJJa�>�>���x��ܰl��*����9z��):�;XF�|��`�l>vw� Q�����F_(�Q�����X�ko�ҡ.���N�P��6b�l ��*ߍYb�V8FO������Xd! ˀO[�)P̀��M�c������"� ��՞�Vκ�H�&��7Й�Ӈ�c y��8���E�c:����,�
%��i����Tr��&�C�������Xx��9\� y½#IH���ύ�9�����'Zc���}d�kD�}��\>ݘq�z[h�3L���Q`#I�͝ؤ�-\�y���>�TA����f���@%��p��} �s�ţ7c�J�Dy�q8�B�^ji���?P�"��L$G��N���%_���� ,��1z ����itj����J@6�:�-:��!P�2z����?�R�-tH��5G4�y�S���X=x�w|De�dx���H����wy(�2QOf�4�j�=^<azY�0��t��9�bb��q��nD�(�@��u^>ߗ�M]m�bd��6��۷��:<�˪�Z��򊂑��h�?�6�
���H���G�>�TЛ	�Y`RU������:�Ā�ޯ�TDlN의q|�D��V0�D�e<�1��j�t���	�͒T�P� ����V��K��W�Z+��߱|�5�Ө�ٱv���k�%	O�|�X�^-ĸ<�0v�Hzv'�aY��H����i:��+��ג��S��EYx���]��ą�j���!Փ�3��-�6�,���^9c������?N��MD�����k�+��0y&�=�*�5��9��hJ
8$����홊+��uM:y�p�T<��gq~w>��u��4�&
�L����Y�מ`�9Y,��f��^p���|�&3�=V�8rvra�	.�*�?[�2R�� [�7���������_ng� ���9+���Kzl���;�9�l���W��k��4�g2uE�l�ag��!ۡ��B�J�z�֭xQ��aS�̩�ӎ&(��|��p°K{r6,W��;���&إr�{)������X��f���e
EVN�k��K���-�_�C9�e8+b�*�;%��y�"�D
�y,��k%[��hi�O��/��/� ��ډ@kݾk;k�83A��@�I�][�1��-w/
�@����_��X�v��Ĉ��݇N"K61]#d�6��ri� u�����	�5,$}LB�	J��)��t �i>��T����k$C�`�|�n���Eʣ���Og���`q񀋘�- ���S�c�ށ!o�@�����Z�y]�O��,˅�����#���9�rԽD���b���5*��ɉd'���i%��@������;ȑBԭ�6�����*���c�Nϝێ,�Yy��p�[+�
���O��֬|P,_~�t?���D��p�{P��+����A`� &-Z|����U�TI�R������\����қ!�b��O.K�vV*F>�H$�gC��D ϖg�G��%HBb,�d$l��X��fcG�2���Tw�߽3h��n���OQ�8r�fW>������*�XO3�,���d6��#�=�A�͹�?�A�=st�@KvL�>��jl57N�P�Ikl�GȒ��jE&)k�b��3R?M�x����G~lj�@��0%�T5+���`(7`�Hk��D�Tc�OA��B�� ;g���ŐR�Um�2�({h*NYZHȷ'z���j|��aZ���r�Ǔ�����P���sKIB,,����v �B��Vb����,~g����Z��h˥4�H���V�:.���B�Yz��l���N��-�t�Z���^|pD�|��s��c���Jͫ`2�[�"�C)πƻ�����D���֛~,�B�g��[��>8w�]qQ��(A}]�?�;�ey�A釂�o�9�l�iS+�֊�:7'�.�0j��Y��:+�N��ƴ�������`+���/��^���<�&�h��׷��Ŗ'�/A����K�����
�3�<i�Ǖ3��1}8�~���C;R?�0�@�˾;��[y\���E�u��F�R:ᆻG
dC��/~���A$M�,{~9������m\�Qps@Σ�Ģ�gVq^�_ge�'d���� O{��G�~U\U�|KݐF5����r�>J�@�%�1J�klBJ�^�
%~���i�{9�p��|)N���6v�QkMH�f/�=U�v�1_�U�Qj��
	�6��;H=�oY���K6�M�xtBu�
�MSf'�����I�}�ê��Q�)�6�a�������$�&�KzC�l#��\�|󋎕,�q��;b�Z�Qj�WNB�i0�)�էo��Ɲ-��I� @|ڎU��_���x\��=��ƻ��@�̞�������1�y����m��|��#-7�������0j�R��\��h]�t�š�Q�&~��as�v�>5*a��_�ԾbS�G�z�ؚ�٧���\�����=;z��j�8�_xo��SP<�_+Qo��A����N�"|�wD;:��PdkN^Lk��q#|w|i_D��A��Y�O-�h,?�����"���z�Z��6��>_��U�y�V���y#g	��Gl�L��1��؊}0�~�V"Q�րac:��L+
�7a�g�o۱�t��U��F�t��#n���?�}�PK��9������?go=b�[�,W_�kc�#��9v��:����õ�e~�4N� Z���� o�Q>��QzÔ�B<mLuϺ=�.��4b"��#Q�K�c�W��~'b$k9q�v5�D���@�7C�U@�68��p�@e0RD0��Q��+Ҕ%��"˟|v�v*�I��/9D��i;k����m��#�#��'ц��R���˪��m8����*�U�&`;��,|w2���t�=Nh⫷�� ]��;��b�./8ՠ�+��X��U'Y�SR2�������sO���95ו�����n5f�5�y>�����
I�۰�A���	7�h�SQ��d7G����ʷ�r=��#�9�0ņX�C�b��k���8�/�&*�:1W�q�+��VHL��ɷ�� ʣ�9.m���}����M��Ǩ��?�Do5�Aa6�X��M�ủvc$���_�ڵ�oA��։�Ӳ�g���L��̦�Z�x++u'Y@�42	.��1�n��Z��	%SO}Xr�x��\h�i$+{L�:�g��р5MJ���S.S_�K),0�V���U6%��>�����F�-Go�e��֊��r�iH����e�lؗ>���a=!xf�2<LA�l��({��6�/ /�v41E���zB�O�H���{cWҴ�÷�H�K�i��A��6.<pS��L9�ȋ0L�)�<0�a���& @��?����