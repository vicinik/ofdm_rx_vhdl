��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�@�9ڇY{���c���2����H�/�7�IG�ף6�Z_c�z���M5.{�5�<44?���k�N8b>Ic���Y)��ؘrbx�A���
'�����h0���T0�F��&�_E�	!Q��N�ELθ幽b�?�"bH��ˬ&�3�[�s;x��<����>$�e�k�Dv�U���{��eA<����� }�$��-���3? -ẖ#m��]~�G~F���261/�Lc5�n t�c<nP�����S��i��T��M�UK>����>e�D�r��� $�<����y�ڣ���K������!ǇG�5��cB��!vղ׃G��&Ǐ���Ճ0��B-߳͏�WҔ���S�tg�C>j�@�f��FSghH$�O<��ˇ=4�Fq,���%D%]>������n��Fx�M��dxx�3��%P.��`��"3J�{RcJ�JQ��s�i��TE��Fdy�Y���8�r��r������w!�~+�|����d�v-���4:��9t[����Y}�g�!ģ�ھ�����0���깨�<�h2w l+-�s�^����(�aك�!���}ˊ5��^��F+�\VHN'����h�	��<�.�k�N�ؿa�P�s��5����J.藈9��L��
h��~� v��@̫�����m����^���o}{��	��Og��ņ��N������S;HMn>���~�\���8]�",At=��iZ���Br�v)�O��֑��y+T��\�T���ؠ8;B^}C'/s����>�:X-ő��Ғ �o�L>I��ۼ�\�r�jht�{"��n�o��=�d�ñ;{bY�����}\���u^!�A&ŷt]�m'�l?u�\�  �̕ت�dI94	�~��ltP��"��C�	��^�]��ss~��]H��UW�(�mv�9�U���V�I���5�,|�(<\�U�p����{$1��G����ӄv[�_7���۶}CtL
l�4D�ndl��Z\s=���2��q��r�0@���� �h�]9ڇ{���bB�on1�(p���=Bq�RJ8M������+��+c�2����G��9�i�K�4����a)#5í��D�V9�uF.7C�<ۥD�D�沝В��d��������vq���<�#�+D;�����wo����BA�HX�j�!�)�im�:�{���UYCrOc�׻�ApA���f�K���(̢�fg�e2!+tUNܮp���L��W�;\��V���~��"����Mڎ>V�]\'�|�r��HS�����&�p�Ąt���{F��3JR]�� �b������ �м,���\�'g'?y������C���lqD��� �t��_;Qʡ��P^�xm��?�|�E�d�BA�t+���8{e!?ˏm�(&��k��j6P�����|3�A�	#�(�ڝ!��0|Q�"44O�9{!����B�=��@ ��g�O��A�#܏ 2C�;K��~brr<�
�]˓d�E>w����^̸�.$�`.�+���/h���=!���ͯ������6����M�.y�ަ��&q$7�|"�U�!��	��e��	yt.��G��F�rE�He��f��3��J.�I�%Q�
�E�Ή��� ;T��e����b׊.�<^��9���3j:���`�;��7���߬m}<�׾��D�J������eZ��O��V[��de޽����k�U��D�2ZC�?:=�<�l�iJB4��Sf!�m��@i��>?����A\�3��ѓ�#�ޕ���m�֢)7B��m���� �0�2�빯l��dc֕`b�84y���X��.��0�`Nu'lJ<
el��i�h7�Z=�?܊%k��S�s����"dt2p�q*�2�}�u~R4z��yJ�:�?��a����؝��hQ�k�7sz�,�Şy����w�B=��Ȭ�:���/74J`c���T�	��.�狀43o㭵��YI�h�����P�K� !H��j����E1��"��C�e��\Sҵ����Af4Ϳ�y�{�K������Iv�OB+� ���3F�Hfma�ʔS7d8�AM��h��-*�.��N�ʔ�P������G�f)'�3�R�R
�R��_�w'W��b�l���/�����S����-���P��{����X'�v־�m-WޔdnT�$�����u� yc�z�6��U\��J�����Sg�����<��Q�!��?MGKJ�F��q>Q2HR�s+��Ծ��I)������>�ZV��sĽ|������iv�S������@��I6�R�\��(�T�!�o��t�N���үdʉd�^z�jy��+�]�o����@����^Y�����������$eVR0OoZ���XC���GS�#b���9 �C=���t۵>�QϢg�E{��>�� �YK�P���Qs�Py��uS�6�.�u�E���0��u
�4�%fY)�f��j�
��-�1 ����{^uw� :Fz����K�s����t�b���o!S_�3���O�	�P���}_�
4��$�؆jB4
�b�57��f�	BxCx�L������|EKR�/ȪG��|��=Wͯ���ܭ�íMc�)S�d�b���&�mq�̸I{�����`
�˔�W������s���7��B��D!�I9;2������ o�/L����v��>��/��� 6^R��H���4=&�z7%� +����Ð4[�$K|�!y}E"a�F�;zD�j�t��\�מ��v�h�E^�J*i����9�1���g���JOVˎ$��;~���cJ?e�@��Q@;-Tæ�s��e�������E�q6F2����|�%�2iR$X�?77���pYQh�m��W=�ɛ��j*��R���ʌ,6S��DS��ݮe�0�hA�
qyţ�' �����3�z�C}	�o1���GqM�֖\>Ȼ�x���,�z"���l�B�w����0���9���.�Z->���*��Fr�wΠ��#����D�[��u�V�b�?u���P�� <�A,�o}o�����Y���t&^��U��4���F��,v~\�Qdg��OL�R�>0�̜O���&����EO����v����)�Vu�m*��$���D����ES+�	��M5��5��x=2:P��	F"G%���X�����ƞ�s7F��I{M�\�ݚzoN�	�p��G��/�?���b�Hp�b�����d��z<�^&�ޞ��N���������C8���.$����_��P�Hh����M5&� pDҮvHl)j���'��;2��3�vk2Y�{&���Y�o�����ʃƝ5$��l�|t�7f�wO��*����T7-�;Ӻ�%;���]>���쉶�����rO.�b�(����>}S ����B~M��	٢|n�3s��[tZZF�$�X�#��R�u(lA����@��7 �+�&�˘�0iuu�g�20�����ݏgȶ�I�/���y�����:a�ږy�Q64~��' �1����`���i�����1����髵��o���_d���;��v+�+�E8YY�T����\'�&��tyhB�c� ��!���4ΈƐZ]g�3E7���cw��E{(q��# ��/V&�_�}r�����-�&���p�ZZ�4��d\Ę��� W�z}.Ŵv�bۨ�S5'�w��(@�sGn8\d:kLj;��*���jD7�I3�9�_Faњj!fh9O�c�}q�8KV���sH������儽����C����d�����T1���7ⲃ��Fb��|?a&a-��0a�m^�כ����$��/\�f���Y��X�J^��J��3�٣N!�%�</}I6�v��=�N4l�i��F��Q����=}���%�SX��Tv;�8p3hf�P\Jå��n�)��G�{$U1GcqM(��
/9X��V�)5ݸtr*J�C��1*���;V��m�:�l/_�"�E�&������@Qg�$�}�\�z򽠶�<��gx���
�چ�	'�P�=-��s@��f$�ˬb�mB�I�@`��Lu�G�nᤀN�*d)����O5�6���V�W��qQ�9��Ma��ls��gd֠�}� ��la>f{��c\?��,��ԁ���X�s����w�h�d�_N8v��p��5�:�����n��+!���q�V�m�rG�l?�x�����%��Q����!�O]�:[�3����`���2��t*�ځ
%���I7�Eo>]��8N�k+�`�v&~��Y��A��`I�\ !��q�r�m��%�MNHo�-l�a˭Vd?�Y�9i�|���޶�48��+JO��P�~I��/���p7M�L� �۽_A�$�a�t[�%}�]�)��7�o�]����A�نa6+����?'�.�T���_֟�߶w(d��#�,����<K��H�r��
�U`IK��B�[bJ��:J��� Z�K��[yG9��`�C��H�>�n6K�Y �N�(	�v%�!q!)9��KRf�����\&��6�^��X���)�AGl��YE���9m�1��y��{�'l��2��'���p��f1�}N�;�hM��Լ�`�|�LP?�l���~�����
J%�*��	Q�LJ�
��R�t>n
�֟�INW�G[�mxC��HV0첸~P��ycY���aϾ]�1'�Rm�I��qH�!	���g�8$^������-�C߶x^9-�0~�����:���/�|���(B��(�T)������og�6fC�]��1&������Q8��3ӽ�Bγts��s*L���?=��+<���|^Mg�����Q[^�ԣ�7�Έ��� n�iwMT[��j���Κ�=@G�|��Uc�m�j�B�,��~y5/��Y�=Ĭ|߉���D�{�������	�c���F�C�`x���Ax#_/"���.Hd���cz����� ����S�LZ��*_�Z��,���u�2��f��]D�;}{]�ZҔc1���+�WS�I��(����Ŋv���TMB��.�9/4�-���~��{ȹK���(YE��&�;/:��]�%�SΟn�bͪ�H�9*G�ꃰBC�
�D���A�X�ЇȌ˯l��tՖ��f�1d�q���|�wl�`O1�j$y�p��.��J��/y��Tn���y�C�����o�kt4��z@��þn4������j*����=&������v�"�a��R�;����n�㛙
	���b�<�?ꓪ�|#|f�_�8ѰS#��#�]�O���>��Qr#ծ`1�	p}ƞ���zT��"ۖU�c}�r�0��x�>H��^���),Qڋ�Ӈ]M!7'nf����NKf�$cS)�ǭ#ȻR��!�A��n��ޤ�M�§3~�%[���c%�g[D�|_aN�0��=�_�B7#FQg���CvDmB��\.�ʌb�T�S��gl��2�	j9�G�ܙO�һ ko��k�AҀ��<��w춷yo�(H55�ӑ�>�E�ɋ�R�b۳�Q=\�mn��vV��	ʕ����a`�M�l�V����$cZd��A���+�֐�.��ø�D��y����׀�D��VT��is>F�R`���7���P��5䇙���$�>��pg&�w��*���������Ѭ-,^�kEzk�����s��oE˗�B1�O���tT�Rڇ$���u%:�K��c�lՑ�|�`^/!A�|�U���V�-���L�%z�2��y�kx*��
�?9l0� �m4�i��#8☵E"��L�sf�^�#�n]XK%�U��P��w˺TBoVB��.8a,A�CY=7�J�����H�ۇ<���3D�x�3�݂98y]�z�H�6EK������خ�U��%�A�Ƽ�z��C捸��m��<��F0�m��Ż�甋�"ݮ1�݌�g�8a��I�:�z.#x�O��K�SqZ�T���0�nMS�$p��S����(5$���ѻnYY�X
�u�>���q'UT��؛t��iB~h�n]L�"V^��8L�9zݲ��<�p�+�NÀ�Y���\��M:�"��{mR��N��жm�&���H�O��"Õ�ȍ�1xwx����p� ��Ẩ��@=�3�5�їE� 'E�L��1��2�}���Ĝt.��B$!�6Ⱦ����"�
n?z״�RF̚�e�LVGhM<�x��3O�vyx���{�_	���Ɍ���Y�/��ו�ie�9����U�A���a0a�X_v��zZ4�pSU������TW)���@����l2��L�P-��i]�E��7���n��ۥ���۩2�w�����lr�m�@l/~3>��"T��]��	b�\��E���S�������/	�]QM��f`��t���ռ�o���i��T|� i�S�#�^~�u~�%�"�~��J]�s��q}�ŵx<��7,޶��ҙiT�g���`M��?��P��c�6�hn�����~z��Ft�䰹�"�4����g�)��S���VP�w��t8 &�1Ը�����'	r��D�R�p�_������� ��u-�&ڎ:�Z�:w_P6&��,V+��U��I��g�w��~�Ӟ��γT��d
��TA���M���L�+��$��#]��@�����e�Z=6�7�u�W�-p' p ��Lq{�
^��06�=o	$YWaN�9��yH�_]�Y�ZC��\q��b�#E7�OƴHV�Q.�D�.����C�� |��?0��Q�L`��@.�j�5�zN~��n��(������3�/�.g�o��Q�Za�C��v��R�@�q,g�딌V��7� � �k��t�����lh�b�.Ns�2�3j�����Co���笔Fn�AP6�^c�Z��[g�w�CP��s_5-��#�Ye�B��V�Y��dp���e4����]��sl������`�C����D"��e�h$wyWȠ���R�"��qu�e����]���
8A�y�o��_А�����;�${�?1��ImǪ4����s1���_ w6! [��FA�]H����7����?��� �EL�%�~���x?Z��~wUBBb<�!n�ͣenw���E���%�Z1�#��M�FW@+��ɣ,Ǩ����h��qC����C<���y�؝����9@����L�_�tmBܡ���m�A��,@�B8A�䢩N. �!��Rxd]�屢V|�ٙ����� Q���$ᾣ/�Q�qdDNuH�ܿ�Ћ(Ǌ�����3������6�����e�Ş��6,�n���ClV��+�����闾�ǽ�%� �g�ԀC)JhϬ��6��6��*կ��֋����&�X��K�G&�|޺%�r�����5t�-F^7�ǅ
S+圕P��
d�by��TP�w������߼2t��G{� �v�b�uGZ����t��1�k��c��X1��Z��C��ݑy�c͏r��h`NB��܃[s��ǇA��7�B���6�Q��oaw�#)Kn�\�����P#��V|4n����QA&+�D�Re���_[Pß�^�t�M5���\�`6��̂��1qj�5u�s�S��M�� �Kڛu�2WՇR�ї��|�R�C�0�v�
�m�tک�疞���� &���JH)�T��t�0��&c:>�2N]ׂ����?3��\�F�ӵ���`�xǍ~��c���k�Ƥ�/{��ě��=���!?Pn?;�H����$:�|�=6� fW�Av�k;&x�*.�M�Q�$/}r��B28�-y�����h�Ĺ�
[7xz���qV3Viv�0_@|p��X/ 7�b��%���ɵOH0�$��9�����3$��N��vS�ҏW��mu��h�#B�\3P���'����0�/[�����ѦŖD��P�>������dH�,���jYH�����Z]:B]�F��CMI�����#��!V����mo��L����@5&��CJ;��9I0-��)I�0�NN~ ~\��I��v��#���~Y\��׈�g�_=�f�5���c�P��*��8 /�{�(�h%���)�0��+I<����1eߨ&��5^{o���ZEOC:-% S�� ����|�S�(5|mrO��_D�k'�V����
�Ac__{�\W�@&��|ѧ�t(l��pG�>aVS�6��p���ު��4h������֟W���F�����C�鍳U`�,�ۆ%�����b�џ$�{,h5�<N<�㵙�/�?3�p�"�)��Z�B��50É�)�aI$���DV�D�y�����'R��2	G�G�� (-O�����0,r\q���_�ESX�Ǯcd�_d�o������y�+{�z�ߛf焸V����N�.��|gU"C���2��dװe�т�I�*���B����ߝ��ǯ�@����\�=(��'��w�7�����0�YV�'���GMv6"�M�;3B5V{:	�����?��1���+�]��`jƙ�y��^bt��#k����m�*�C%=�º��<�,��l�8QuT� Qs�Q
���¸�� |*�ΏY\X>�]&_�#��-̌����c�an�
�y=rVf��!��sq�P�p�	
���^�4�����c�����1D1��L�+zb_���y_�M���R�U�h��|s�����