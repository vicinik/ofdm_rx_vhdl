-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KtaXdWB1jBlEyzGS9894gdflAI/ebUCBEix+Np6k69OwLp3yFEiXvKAR5vsDngOItat2k66tw0ZY
sIAUEjeHtOmk6y2iLQCO6BJfLNw60bXxDt7ftitUooPyvFUC6QiwUlyh56wWDskWjqDH1HkUyskB
0k6DGUVWr0oqB9Yn3NFE9yS39Va+CXDScT/9veaDI16B3f1aCMJldmlAIGyl4jEXN3BCfiiGMdhF
miQjCUTkZnXY0lk+5pflzRtLFIWOZ8hT7u/mBtwjQPwqY0YP6kYnO3tWuzq66pnOw3kSLoS/lC5B
nV+qDPme2Sp8kK4aiZWDXN0lPbpV+nqgZDQP2g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23888)
`protect data_block
yh3KibTTPWNVN87MrJ7vU6e7cOAb4uqnnH4rV/KiVyeDhgpRRPHXVLOGLqLgT+XSR+wttqJc7jeD
7/pVFniO6Qlwma/WOc/JtCUWqhoZnNE4hSTkChiHQMVO7p8bVivUtQUjXybTJifJ/QLf1sOKJY+i
2fD/gGq0rcmNEUvFg5co+472AJvfPs4909QJM6n5eo8Xp0J0wi60csD2JC/SA52oyWk2uzm/vQEy
PixFFMKPgy6qVrv453J6VszPewr+RtWG76OC/d9lBLw7WpuORzBE88J4wLGWOlCTP87+rkKQCjct
yrgOr8doCkrQDlDF76K9V3FkOKFriGBGdKWtV8+PexatNE47OLd5LzQPGjlioypxEaVlhYheky2C
xrdMIcS2e/OPvCiINGpswl5JTzoJmdmpctcrZwrXUwtvvvDPkC0KnuWtxDwkgb7zL9ly+G6p0HTA
SLvHIM4rn4S+iME8ds0EoPvpq8fXFKfbyAwg3PbPlu42eTRmPQuGMwWyhqLNrh/q2C9wA6u8kQp1
mHOnb5dE8C/fQL0iugLQAk4EEkKleUCbUsRsdoqbu7ga1PMQF0CqENF89/i9vFCgRyDDb6osgkYz
swLaFD4GVcRuZFh5LZZEBzQaZCe73xebIiiVxM45nnTqfXhPbfoltI4Dcfpls+EwtYLK6d/+hVcP
RJeHJ5jkX+Iq243NZ7ItkSLw/Y4xEhahGZt+FHH2187K90WNwZ2ggsH4fkwYy3amyzbZXbvPaF/H
2RBS3Ao76HFPiiyCh7k21YDR6QEAP35oBwgNzwdxuQpsenut3cT/1xDWMROUL5mY7XIgyQHHw6AC
pZ0+2CTjEbAyrFyFtUPTrUCjkT/InSX4YXv1BtGUwKHPWJi1qZUO8T42qP9qG+TDspiz5RdBxvDu
GbztLnJX9ALyxcuFuQZwsMbrC2rd5iDs80j7ct9vEtRtIkVShH+C+lxoFIVwd4titEk66ZNbSroR
NCtf0nVcqdncm7abfUZnVkBqr79bbq8eeQ27I4RFgBmUUBPJ0r0hikrOn+m+jsn6woCshBKECghL
/VfPSizD7A9/Li/O8TX3FdrKvkJ/ASd4FJfTzm/3tOYMquvML8eXX9qtLSgIn+ld3Va6bNOZe6lu
uSJUcs/8W27xMZegXFItO4DoJF8oc5TIt5+2tV3mpnxMZgnkuow3+hjP33crubPyXjpr+lBgOKkE
8I7992RQ6cqRMU3+hZbrfflikLoio6kIFCgozEgzVVHJLru9RiFdGfyAYfEyTazyaSGn66Qco7ed
9YkA3/g9l8PfRLMfXhzudRp5sx3VstCdoz/WALdEdhj6crsXdEPkh5Gz8+SwS+6nBRuf6yD5MVPL
pa20REm3pR6vcy9QEn/IdtGAfydIMf9FVX8vs2SudeO/ifRxrU7vZhmVkgg6TmKh6zFnEA9ShwF5
LrCOmPOrhY0ZFHjko2YBaea1vVVT4HPVXaKOtD0mmC77TCpWJaIR9fnf+7Ej7y1q8nVPQ96/D/3n
wHLteVY1xnGq1pcvh7L+lkhG2NJRy/3Tivii35pp0ofgy3u//b7XwwW28z1e3Nl4AsRCbO9oAl3W
GzHlHI6F2XNesADIue5Xt96RRKRZyBLJr/ib9dq8CC7G4AQ5VdUMrf6EzIVsZAiYjTdD6IabBrcY
5DSPEsb1VbPMQygcpYdi0I46xcvk+wgWxxmOG9i5oHbjO26RFYXMilQvkG2Kqqd+m5l4cOMR7suZ
bTmGik7Xa7yfnwTIOwybtyjNFvsGlWzE4EAhNcKUEM2sq3UKcb+t0JPjf3fa/DHShuAVNgNmhQ7I
m+UitprePKlJ8UkxorxnwT/XfEvuNNXte1R9SpIh0Xr/WG+chaL8Pxw5p7v9dt41Vh89iCrwcZK3
gdlG5CJpXJl+g0yPW1ihFtjxHtV8dOhei+UkrwmYCw40C5j1t30yvrBzFFQ0q4L+v081rGjDcoi7
Z/FTcBCjxxTmHrJh0S33YwEBSZPxXJiG3tPMCFuq5RjPsBCJptTXpHS6pBFScZtHvQTHY3FbygfB
il385MYk0197VHYyzg7KNTdqa/FCZo4nIPOwFB06GmZO+ecmZHogzRQ2QHCTcoQHO19Auqme+Rd5
+J9vHgRBJi2EVluTa8iDpEgstoKEa9iZ3Yy6wHGZ8ANflfpqhdHk6gxv309SiVBw5+9hpxq5y1Ji
iR/uGiPvJOAx+yzxLXXohwhD/2AzQSD9Zj12ib0mtm+5bECA3IL1nBO+nPP72fvxTMZg1kAaNx4L
oTct0yi8+SalFnr4A/d9KRyrxVkZHzQ2CuuPO80bG8lxnpmWAmiasFl2+6EttDerdqTRiXC+T0i1
AXFGJeoH2rsVzGlC+wKhPdRWIp+F7biW5OqnsH3pr9/kwXs3Ux5liVdtNFLNFBYAXW8hGJ6zXQLj
V8upDyMOn/hDPfCbtK9f/nr/TOsy22Gul+szBhsaBtOJ24hpYlS9PygqOPZLN+xdT4eP/ENlq6RT
FrHxcInJD0CZLAt6L9QpZzetDiwySplWNgrqBEogfJ5Jhr/zFbTDkE3tV0N+JiMTyewysJKg39ap
Io35lEwx8YhfT0ZZLjiha0WNkr0BibHifzPYPcA+PtXzVaJPK5AlQhFZ+ik7tZN0z0W1WHLeKTbJ
mpuJFwO6gFoOgyIDijluBQ1HOEodjk/+gDOufPb3ZoncY7VbRTDmQwKYPfvn8TXDjEIhQDQ/Mkc3
eXNh9FSJBOokhDuI19CnQ5/00Wd1i073eMaa3R2eGoelHOx1RE0MzxHCpFw7MkpFXs9/KW1beEx6
usBe05Cb8TkI69bQhelBTcW8FnWv3pJ0YgSVl73HTB/pldzhAOkSUgD/jEHjtK1XGEKY539JRPQU
pYiuK/U2+kZgT/feOXocDl9SyGgGRsaNF+Se2ZUP8xrEwgQ3ylGzkkerZBf06nDEHo15mUYWNhPb
jCEOcbMwGQLN/DlvOlCiJJG1owhu+q/PXG+pks8I3YDB4I1oYMgANOXdjfvXiihwqpnWIfwe7Guf
K7WxMpSy1qUbVK0WFb4OrVL40VNrfVPSyGp2PcahSjVqdkJR3QEZ3WY02N2klBzQM2St7Nh1GJs8
ZjdBytR+0L5E37CvYrLXbkrdTFwVDFWHPEW72NWyahwFS0l/Rtmbsk7kguySxEP1d3QViskz0VoM
IBFcqq00xcT4GVtDz++NCKDFtYdsrqODIAYIwHkJvXylrGUov9MHO0kSVja5ozMv0dOLvA2LXNI3
bJfohVbeM+RjLCotacJ8buG+7Re4HjyFBZPWMp4jmRXUSMH66SWtvrrnlq5TZa66UKHjJ6P5NzYf
i3nBbR7//3z7n5lLCJjgPeWcmP5Imeqo6mnToUNkSrXYV14Sur9HCwSg7apmGL32ctXh/zhE41Iy
cgEhUrpTKhfAEQ6J+FQBx0l/E+vrYzUxEZ3Ajc3y+XFyMMIZji0+4kTjdWE7C6m404T8+hAVPdiC
dQYhCWfJnXdGOLDol8HqifS38i0sQ9gkhft0Csg0s8DPuOn3yIJKKrMvweFLokV6jHuJ5zfapVcI
qhG3Nw99W0VWSIpEsEsZugFBdhpGqIClmvEgu0Z+RjVAgcPyJ5luSJ3/3C9EVRpBHRM4gj/RSpYG
sgD6iZh0sIDkFxtlu+5WikiMbNCnYYDlBW2UMT9qMoP+ytq1go4cFAhQpdfJleOleEo2yTPRVsMI
28O3NnLgmEXf1SRXcQ+miZxi/JX63Kzwji2y40Iry/cgMyVs3RvlC3VfuBx9gcFzpz9fGI8/y3rR
H1AE6DHUppw69Cw1n/b0yG61N9SvCfHx8zfiEh0ezBbPr9wQ21KplB1f+aKvMNZGWsWKG+FqW0SD
BYvlh2/fJIp0C9g6HJtrEXnlcCkqaVjCCOvSCGqn3Yfk+ZvWdGHIKWLQSbXCyWZ3ibt/OwThZXLd
ThubAOqS1GwP0L+LV0x11YAAJGw61N7S97iSqPk2/Wf1RzGZ1BwfZry+3pptuPkJUwr+I1y78AUW
IZXtYOQwClTO9QJIHzMY6+wr05lUgwD/xWc7rVOrd3ikdVwgtAuTcplabUJ8OZYVjNeyAuXBjZ1q
oAUJeP3+zMabVdJg0r+nt9nrhaUXdtT7CISKvcAyMQU5cglkZowhd/ye0Oh4g9xTwDzMjjAZwu5Y
AQ34BaiBxpd7SMBL/MzfVlsF5Ecqq3HE+3sKu3AAFYoDqvgu3Q5AgpzD9Yt2yUTKrhzzA1m5LuVD
pRZKSW1ipo9+gtWnH+JPGtzRPNZ0wnqNctsUeaAjGkrSmQjKttcygNdcRyXNiJ8gd/klnIeOBhMC
Jz03kCQHwdtSS0vAf1IvgSU/srgHieaInVDx6OFua1O2SGsTR2zPaLeBP3iiabwiGODf56eay9fM
h7ivwPLhTZaiHMQMy3YCKA3vdmF1lf6deMYsJw5Oixa5Yr7Hj0tap/juCxhga0QCHNzUcG4GZUIf
bNstDH5RgCwoWm2iZ17WYj3tWfrKDNNQvQeWwuoiKjSmaJMAVwSSKVoXqnc9H0MTu71HgV2W5Ak+
zgluU4qhTpNUCyD8rZWIFXuwvx94hyziRHGWPIeZy7JuBcunr1pQWmzyF4sVEOW1oFJqfy4F9m+e
faNRaYiLA9HMfwCZYrVOE3d09mkMsSCgfD6cK5qQF1lNmmbFIoDlatKbXqJU5Zaet1zPUBkpV1X1
Bt4qS0DmyH5l1k/uGbj47kKiv8HxP85aO9ZO5DIdGu/hAJLzZONG0mRi3XeYOWwCrq3YjuCC62ey
gZC1xCwAAMqltNPwNCr3kWPthW/Z0Hn9XdMS8LtRRUq5zGlKU9QjVzsIVUtMAsS83qyIVe2O8uff
3Y6tHLvJmeoRaLyoiQor9iva5cWRcMnrxcdLz09709wum3Yb7QueaBjAyb63N+7tXPeGxPD3qMJR
NuIc8fM6LryBD3Q/8bMsoyRg9wB7BILk5XUq+qfUzOnb0dZ+ir+JfTP9VGMLxCNb552UX0JwGL5F
TmATo9FfZ7Wck4CSJt2UpXFkZHF+3wLgCoBsUXjdP0JcKpCkmRZ46EkQGrAioQWXcMBqZFtznIkq
4ZlDXYdWyEp3VIgV9Nq2KeZPq23e3cMG7cNpIvmz0GFgP5SO9qCqI6xyp+XA1g3tguNMdTgx11Wp
4Q3AH38WxC379C4zeoThBohxyIca+ZRsPL2XXeNkDs9br2tFAgCHcUTz9taN+TH6msG/Qa4uFhi6
1wkv1a5LIU9LkHQhYP0cbZB8vd8EOZsja4jBBY6EDv1j09f14EF9q8gczDbr6D3O+ajH9v3Zp0ss
eTFbvM/B/D9hnQxhLz5/jT+pOU6WFqqFtsI+Bq3bPEMXZGfc/Ha2J8uryKeaLMYHI2Bw+2maPiwT
1EhwAj9NvM/vvyQWFXA+boDqgsEo7gF9pLMKZ8infonxy+GZwzUfaAMTX5/a9vwrrf9wttyIahKj
MxoMpZEECVFOWu30WbeORcPPD+3Gj3q118XHpzt0AEJljJaf6X3dwTXJNvvH+ssfUWtd2Ti6n7YX
jP0dSPrlSFBGyJTBpnvCMmBiudueGb4SM/DApKwMmuZ164g+MoeySUiKDibK002BIeAk0BgnLYM4
Uq/8P0TVNcFB7P9/edaF6sIjdpQETOVZOCQ5uYyH5pkhtNwniK8Ki7Kxa7RjBPh5byziTv24t42w
RNl9zkM3NfT66Y0VA/lzHgWcFoFRWcDGUPBRIWdyEpMnz1xFllraSR/4LEX4B/do5T6CoSzrMetT
4631GpXPQDa6/KtI/JFZw0lpL9qSGjPZztSAxB7v0lgAK7XX97x7ejmPOlOlkPX+Cjp6ok1Sw3iN
ZeMmFnKdVAq3qOEXjq102ipWXLCdrVM5LzpxpSA//llUcx3Z5NHnG/0DiPHfkI0CSd4V3/oaML7L
qe89I0lNv0naJ71zW0qs0wuFg6K56l8jOegUhModt1buYYHAwziz2Nvyf8Ydfpol6fVfjHy4tIDl
wgidu+hH5rSak8Oc1Ik/PbsE+HzYpioKkZppvSwaPtP9mWOMRzI1o+0OP0ZJ/mVFM7wDKva6ta5U
jx2QC1SwRncRjKURvIaO5Yg+R+pXcTzbFIQ0KCXkwa9hkTisgo7SoeYLcmcQHjNMB3YJJw/tLuW1
9Lk0cfjCVRAA8nU4FnxmwnwTpKDwVm//VIdkgyqa826IEyJoQIbrkwId79brherfqiJaOd2ujcTF
fl17RgQnns+oARnQyjXRtYrgDReeMfXbInSA824vo2RqB+JujX7y8JARiz+jynCLxXflS9uxfKmY
TKM6tzUzHTePVFHYHq0R13Qj1jpq7oz24jNVIJ+nYzfiTp71c/ZPf74YDRGYsH8pW0BSzuKD/U2M
+4UmNNKG99ODf7DFF+ae7kwQZLW/piEG7FeKfSxds26927me0iGSsrghmqZLzdLKFLqFBQFwvINe
JyvFLmuSy7Iv6oMcnCPG8pS8K4JXqb1OyPFLWr9w5J7kD6jHWko2KHVpLh+H6NxyZy8Rj+5qSM9X
nB4reOAzzFwrNSpM3i01CEHLPS7A1du92DYqRsfPQAugTlcXQdRulXvqlmch6lfxSKTm8xvw6C1S
DhXH1yAeGcln6+iMnhyv5q2nSPQKPuubjtPcroLrrsxXxEum8l1U2RHurWJUsFR4++WlZZGXMLuy
XQOsV+K6kBmrTPtAFbDcaraS2xi4T17H1JSNLnzMbzUWMhNRn8M3dcQFXmRFTHNNxdYxksRmW+57
LYVI+TWumzR9TVLMdoPkXsXKdnmdba+TJK08vxiuKBODb+rulbzmsJKL0WwedToiCH63U4lgwEoZ
I6FXzXdZEXPJDLUHrsFOAyImGCtCczrvzke2nnZBWpeFgIYZoGgC7It5SsUqSyXVuS9RhxNVshMp
LsAoarfSN+TO6Xo2rkZOYslOSznrYR5ehpzaqrb3cOF24vK2LtskpjbW5hywSAFM0RwESroeNz0L
JQic+BVZM48Cws+W6mQU5eXD6JtjU2y7J6cAPKyxzx804H9qUx8UZx2YBvtEz78PZ+clo4o0pHy6
0eFPXp+9nRj4z7QOfqd9HhmhE49Ufm0+j7GVeRiFrDR4KIT4VceCMubwz/5/V8iK1/KaDpOgkLIP
8XbPT9S9KPxG27SFIhSOJR44Rm21MS/dAgS5c3Yk8s0u5br1ai4QT5lbWFGOkg6OLaZL90+7JThY
5SvUDAVavQ02mB+VE5j4neBqltByKWpNB/m75Bu5hS8KGln9C4OEI4XfHWaZUsOVMiM1wRCR75ut
U+uNYM04x302aF7YAihFgNlk04v4Gesj/24UZO6q8klPg9RYGk0Y8C1I3O5rv8riw/GpNseWKzYr
jnkVF5rWtJqYX/7xgDLbdl/G4V1+M9aqV4dB6eqdGsJtCeUTdZvt1/ous71+VLdw+PmGcZOQKQOp
5NK6qtJ3Nr2hqHMGlFLexMGHwKce5zqe2mBTrKS4OtN/rwWsDqSOZKt00ZHXgJaXxiE6oe+3b3hl
4hFS/Ig/EkEEspXC9vv9cSbTZGm7KeRyV2fLe8kVR7gwiXsHJ/lnMHXOJSqzPnH54nW/yi+BkbAV
kg0guC8jDDA3Be2L3aZFdLpprsTQxlySuVZBJtsgHbbvbZQc5wmik8VUBYS1N4PjetIjLzlpRd0u
Sd8H/cbrGTNf655HsRLrG5v5oHjsm60jPdEs1Clx1qBHG4/7w43RAzTUxHwFdQhd9OU8YpYf6wCA
+hHIYbhpUvlsQdkVPf2/SU+08QFPOkEKC4VZPKmUucJsT0sZ+1JntySNGO2ORRG3IGlLflIAGtk4
A+i2F+9N0wfWLMICO+7YMJOREMlZ3bTbsTEB0H3h7CqiIAMEPf9lw/ildXYDLUUuR8GAvpzAZQN9
hBl0hfevZDOd1avNEjo5fhE2gyX4asnjlNq9PUo4O2Omsw/+Nb7VeGxe2JiSWxCQc0MTq8xwIV7r
Tz1YZJJLGV7Tov+F3AhsHSEFhPJvMhmzoHTAkD+1CHvlNmKpgVbIj7g0wpMOjIfuMtNV9zVoELYk
wjtMnKYwQYqiTRahuhmiOIciru+ukVjjCsNTmm5U39eOBqvXmKVdINEEPlE2sebQhw4etESL6oQJ
b5vRnFSSSRo34R9utQbwb7AV8BWrtTvrscEhGCspS7GWtTA96LYLXs6soHKHXlzsu5d/fYq8FWSd
io1xPV5M968e+3JZvpPLJ4ycPYcYJWAYQ+PqEnyvVObii9vtmEGxOmyZy0Ovdden4D7na0ltXcGY
8Dq1XYr/J34YeLNSdGzQOzZv1I8mIav5t08mHHQV1BIBQHzk2zNOjA7bYs/RcV48J0h3m4Nvik6E
OixiQgQ7AtQBBjVix3xSH98nKqxTqL58OrPi1D/uIwfcw+gB3QjpSls1tXA01J1fYfc3qjPTJUBF
wxp4GdzLhbhmii6aVuILVt/BVYSMK20nRlacipCAAYYWCpEiH5BRiOHsjR3mpoDSNFbS9Mn3nJjJ
yfaZR3OHMjXN7sgcOQ7rQURJfBLrih4OBIeP28KnqZg0vPvaKAXRHScTaq0cmYk1Aajh1ZGyDFr7
79T18tAlssOLmsgPJjrgqN+5y2TKoqnFMkJD1oEDlIrTRt8hptAYKWKHnCZRVGg61fjHbYJluH3B
21hzl9pnPQQB74tViPAcAefy2tJw3i3qDivzbhXWS50oZRv5XjaMA+loa5YowoNB843EIg5oaCQA
n40dngOCpcBjED2wAk4203qhiBItMK/0EJ+Z2aQ2IE+/udb3ekPq92aRj/49aOXX/FKRpyyD2GIf
D967o3YSEPxE0WHP5OM2PsA6NvJU71hza52gmzCobs/HSuOwiY6uSR1iKFMTlFZh2rWdlMMimlYt
92lzvJkTyUt0n0w4XJT9WI2zaTpq51NlKoJXREy3MavH6eE+0PbrY92e0gg5AVi8zfUizFKR9fwv
ylzk2Jq6In9FKkmpIceGbqu4U2ctiIKT1I0Mgr00mz6rEGrHAZ2TO3eGx1SXpqpMiWU49Fg7WmOw
6son4Bhe114lm5Jev/+6WT2ohGTaiMiRmcq4J5SaoOsP3eGad8EgI8H64CXBj5KHn/W/LJTgjRbq
Bj0W9hl4wOR09ZSZ2tFj/idm18MmCBaJlh8aL2npU5me4jcGY8gy8ocolKzqTkxP0gQdsDfRKSi0
evMWmeK5Z1SZ5g0hpFTDbLO2Oh9V9inEeZXSPTG9ZZWHdur1Wz7TtVj+o0vImBzljEN6VwXIu0A3
YnIvv+xFNwuYjIVlMjvP0TOQPrS9MKzOw15tvkdQdf6erAmF/mitRaW917OGdhnqH/veCqCVtwiZ
xIZ2kV9CrCUO0nCSV71TKXx0Bn9PSEViZ8zVH5A17E2D9xuNzNUlXRoz3Y55p80mf1sF2psBvlCJ
WzbQel44nyLWKQL64LEax6RMhp9LRWooGxS1a5Zno2twN+oCTsOUjI1RdlHvaxpvv8S60xt4czfl
A1Br/hFnvPvs8cr65IWNqOP+eQRa2FayriuEJ4mxHDlxQC0QE6qvLFiEvzy/NqVJQKsjEhJc6T6/
evTpd98akd/ICp55R/uyKdcC5iFwl4YZ2XtFhrsJwBgO2z/738hZH99qTaSuGJhnwwU7ybeO3mQd
YF7Lm1OLJzXkRcO77mgyHrUrqfFn3Ie64x6K691EyES1ufE00wMofR8A1wcEjeOMjPJzhI7fdf8z
ABIOZcBU7Wb5UZIDpHwcXmUPc1jfdvuBb6214U1fTt4/TxawGHystrxr5vCCpVP1vAgantSCE0ra
VA6Yyg4LGxK91uqpm32+YBvNNqx8a7bsxTyMBllPFG9JVl0M1XIAetrJ5KkIBFbjlOqvidZ+po/Q
tGqtqp/I3RFi7QClg8ZIJY1bZOgDcl4hsod+nnLpRD0c0bgxZqrPvK4deV+PPcK0f/CJ9XQcNDJL
DTw8TfrDLfWmMqgBH331Wy6N0l9LoxEe+00sVzi/v4F4rEQeM4XT7PjvLBmBU6gKxiy250L3OiKL
iC99MyicM5dMN9ADkMjvv2RsV4yupGe8U/GwFnNJiVHfRk2/RiMo6nPgJa2NqYBJbHfSqjL4pR5I
X8XFn+gXRfQ12Xg9XLqygCkU9V1eOdsqXsNpp6UtObEm7bJaTUTOHD1J6WTym56meWBsLHitx5/t
T7zthpurhEqyvVw0LqNpwXw4SWcevWotFMz0/MZUXWna3iOBGWjy0PjVAL5xATlNfNBLG4PcO46e
8Aaaho5JPKD5N3a9dGWV61ty4AkRMjjs5RIFEK+TMUtiOJLdDOr3gWgXIqdygVhMK9XL5aJe8fK0
9ttAm1kmch6RY8VSGpYUNsWRU9Wx+2ugZL31Ibb2K2aGr9Whm03yRpaLQyDz7GFqkgOqrEu1MXU6
BZu8RejCIFp8BucvWUPKgKz1doH/Zse8dkC/PwjNNG9XuCtCDyLkAmV5kGl2RUQpu49lHhL+EedF
ZkRdiABlBQwDIljEoH8giXs7FjDtfpAGBZLMJ4R7kZQyWbbTVxZJ++Ov1u3EkK3tYMvZoTyJMrPv
QaTpyq1k3FVJkyfcfXRY8zk0xw70IQiN5FrhHR6S4UHljOwRQgqtT2PRnvlNLhT1huBRjmo2KqDq
jcQ+c4LlfvU4RZi9Sl4iv8tQOHqn92S8/GevYcknuU8sS0/VcS3UCKzzaGsfjn/CzcNKiWEmqn8d
wFbddNYJGFIEEwDOYNtbvDTZ2irxzMRGRa6pU0bSKHuHA5thyMWMi8M8zTTfaJKYXzRpFlTmbNxn
1EIOikSMSdcvgslpZrP1hIDwI1exGxd211xYlTp2n/2yt93nqcyTkLhpAkYp80xDK8u3B7Iu30SY
5Ra/1F34J66HKHEns+hAhOyRj0nHydsYdhIQbMi0pUAK/JXW/nzu9mF20zeBxyNiiKPs+ZXFuNBz
Vt79mM4rkglbMM0xV0cqte+P3m+B0jK8A15qEcz8pqUF7O6uCfiWcu1Dh1sxtEjy0CW2yl2C/Ytz
2MB6vbQDdZQI5eyFZ5FKJEHD0LM6JHipzGaWt+S/y+Z1Req9Au028QyL9TCvpJ5Ff8tEj+yw7eUe
6RPte7Elf6X046ByEHD8eEToI9USQm2IwlUMIIuOeY73nW/+jMDUgCuv8DZ8J69gfoHVI1j7/OBc
FPVaAQvkVue8yRO+Q/w7T/ln9KBysTavaWwfDFKo1mlwM83e4+MVHnm6xhraCUopogk0bn+TExCN
0c7Ksll3WoqBeGbDr+J6DJC9fEYH1QRCIuvHhoTog0zGZErWt3sf1/zVgEVeWZ0APF0A1FEy/5w9
kqnrPdBbhCXVg34eqZ2+Xfljz9AbDicrfFBgxclemdsvE3E5Pm6bFM2CFyZK5NR86K8suvD9nCPX
PCGUFDMw3uiWgerl81nUSdmIQC4P7EZnEqDlMaKzbujBQtCFBIEL/fWRRc1mEifTYR4EWAPDSJqi
8S6Di/+ho+2x1B+vl+lL9PBYrtm+xRvMC55uSDgviKRxFUVPg/VXioNmNJmOOlrwa9SJyW6G3nti
gRYCj7WMQiklhKpCJlCb2w3iX9yqrzA98d/QePo9n4u7U7dWOYUct8Uc2HwfY7FQssRjcigBBmFI
+2R2y2BjNyiRdmHwmrmPuAdHTDd4gng3hGk2OW3uZWeUcFXxk/PoK50nFJ/B8mDTCaI2LGzojYG9
lK19nXUutkwd01izRS5HCrO8rnIFWYdd3XtrklECSJYcSmsDxwP0QnptFodbYrZexZyzMXTexdVS
jsLeaVU7UU4BN4eAMSF98RPGHu5n7tI0icG9fQLzeBNmGzVkCN8Nt2l2+MXOG6g3s+fuaS1vTsFW
ZOsqSocYzmCMcIBiqlr2iYM20KmuH77jQV5UbVJmsPtZpV65vei+gN15IXOqRmCpf2VJbtO82soW
vlip+DeDvSvrPDKFVye1cYbl0r1qPc3qRVDraFnfzdQhVRmjaNGhN6o5VTMPDCAQkc6i7esreLoE
9X0oX1Sd1POeiWygLVPKVq4OuWVuhWbh6K7Q6KDa+eT+3tJK17xdVMBXCRFYaHxOfwJhdU516wx5
vjxMcNuI2mFtVxBxdgApzOC5VUvCA1n5SP3cOScctAD1SJHPoaqhtPMr0TFsqtytySHoF6WYDmVI
BJb9oenCiRels5g4f7t9dsU4QMoScbueRewMUwaWOMf/Z1tbBE156sU7KVKvPM6B73hz8OjAmpDE
DGcOqQWx2rt4X6P5TvPNH/MTvqMiGdBDWbW+IkmzxzUyARASRWVw6SyatU+e7xviOzIEN45ufzkI
1JdSlYrWQk9np+yGTgkwHkQaykGh7SNOL74e3UQQVoJdfnRYw3tvIMmow3McH7aZZpocPZUjLkAI
DNViilTux+vuOB7hURZoJRVbS5C9F8wdAN4k1fi0AQ/RVPF/3EJfvMgae3H3DrQyTvt6wnTYsdU0
BXKA2YWkMLo7OL8HtXK8SxeB11wn9qgH/z09FDS0830CvaNWCfZaGfvy1CGXQ8tSJVZZOJ2KXzY1
ibIKOjBzatXOY1GqFu5z7Z6GLMuzPSgQzAE1EGGs4N2Okk8s9/npq26rqkELE5ELpa6UdnD1D6FN
YbienR9NI0++JaOKneGsvV8oKNs8jckiVrfQzlOoVdol3BGg/GW9ZZCxUr3Esv/1zpffw45MHzfJ
6GJHjbKtX8UNYz21raJEYv/gZ5x9OEOj33ahFjTdTAN8QXx+SAwOfAtL4d4q6XMDxTH73NqaihdG
1uRFD4PLx8OdYj2Z+HUmGDzUU/OXrn7A6f8Ov+/jk0KG+fATVN3Z77BVmuwh4lKLzTfhE76yPCcI
Uc/lfadk6ercOtVAag3H4eLCSCTWx7manhuvyObg/H2awLBVZNTMCUQwJGmpS2ET0SASmJqGv5Td
oFo6nWJUz7sgMFle+xCbQQM4wEpEXCfmLO5bKqitlhFLmLiD25+LOT3HrKUrdXckY5sRUFchjjxV
lV/dk71mW/yRpDel+cpZCG2meKyYgPmHigX2A1GLlgRo/JxocYsOPcGqTBpQm7+U0+2F4umyh3LS
eatWBc/vodVn0kpVsNJsRJIACOlmt9uqgKlzl1KZ1f8wWflaDvAWq5rZA0gjCIeUUEbZuZAaN1fD
ezuUqbSrug4mqk/7kXecEIYmpDRjm+gyTbCZ9Lku3k3H8oD2q8ii01hhq5rzBv49JjzTC153XLme
MKjMoCR9MivpDr5WQIX0S7dg6RbamB8nfPR8B8K0autQ+yJKxMCm2S1ixQVZqXATrAzRcHPyGVxv
OQDdm3njdDseVF7fbenEKCfoU4Q+AD+YxFjL3WU7Pt44CWi4A57brpgl0jP2OJ3ePt21x8VAA26V
sI6wHof1nBO2WwYncq2ykBNfMvLLSkFoxGWCPyk7Y2JMrXScIUBW7Fw1ovHcx/XhdS1aOVVfBXvo
gAmS8TCVkRK5ql1BQIIIbvBUe8QXdXIs95L6tLCytGkuMwaPJNqIZm6vsUpKuw8c6MJi12n9vxdR
h29z1uoSucF+qPRvOwgsav3rTHn12A05zNVuPWyZIXOV1XQcUPJy6O/4QZNFQE7mpWX3Bu8AxSZw
MQ15ZXUN1ad0kUVzEztrlK1zYrcuzGKVGVyoRTK/eCFlwjIw9EVLdnnbBXrXHXxcj1ME4myK26Me
Fqt1EOYIOWHolmhwEckPxj95/MS69kvRWlFlub0d2YjbUQ34UNoO7y6s/lUSLoE0aEJ1j2e9sPw/
iBcTts96lScJ29wEbT7ZTSmoWwd6nfPMAFMU1mLjSNS47KFbmsenylIVu1+dSQ7GvmNg9WZEHA7V
tI4ubzW9btFHWcb4524MkCd9UzfaYYcywcS3kryehbSYjkyBWesSfUUKDmmrqsppSdspcbsYxetE
YYvANsjCjqj+argNsYgwtF2Gf4AiWtoETRcs+u7cjGMBm+/ThJom9jbV02p/lApychr1pLxppamC
Nh/H6QvPuAhB1Nx+zbNU1M6y7fns1m5zvgx4mEZvLPsYY1pzwZbXoQ+6MRYP/NZbU6UoHz08PPwg
KI1fSSMzowlS9X7LK9UKWTfSNo7ZQlMyI5Kn1/Z/5Tkp1LOr1TLnGsHFieDcqm3132/kZt/aH5Kk
bNQPiaLjXgWlf3bHcnA+upaIFUQZqZO+4gDpb+f0fPCgebya9/bqANNnnMq1ismY7SiCkbqChMy0
QW3UWrwCtFEmO4KnC/AtFAUxis26hn0FjgKZKHKwG5UW7mehmKQmizvdRyWGRW+VYOCUXBWy/MvV
DqN/gD/fd5U8MG1K6LSbpRtaLyH+59WbTZI02pZ67CX3tjCUJrmlIv2uORa60+tAwFKzr70qz6S4
mzcEitpdf24qvez3/wg58xtfdQ+sE5YOplVgKJHn8rkdQSWAaayUwxJw9CWIivTt62p/hBy+FCVd
6wu+fHZIV30eao1d+MKKwKSRifapWsfWfdm1havbW1Bhc6ovn/ILP8uYYlmp7/0rlKs+3ZSi0X+C
+7ob8SgeqxpF9BCPPhC5OvRAaNwy9gM/GzfIhxQvH5Gvyfu7J+2kj+fkO4w4Cem8X9m0fBWDF9qq
0H/wDf8eFfbZ1ofA6fL8UOf+8PSq+BgJB51mbOpZfGuU48fTpjRlHPyHP2WNp+Xt4A4PaR6WfoQb
/5eBgm31L1Fb77ai7DG9tUVE1WR+SiKq7gVLtS4OCPjOiyI6QrR83jBdIHITFM4IMMei9nIMaM9p
uynBfiHEQzE0Mjra9YImf2pckzGMA0I6UvlP4aEMyRj2Gw7IpQfvshVwKi11ruF3cE+zhZodorrB
Ti9WyZ2y2HbySNJCEKYbHykBn/HXGrI/SUcwjlEyf8Mod4/7hNZtaheA4MyblAzmFmNP7VMUoxqc
fBOaCAOfoKwRJ+fv9/ipt8eyEjXnfIRx55+3JYgEQbMZMaqkZasP4M3AwmY4t4cTptQvqBdqQNiY
QRkeRTSJXbnOjLWOeJIQi8nT0UAhm5eRaazB7Z/QrQOSaMt2TM/heIgq5KWlj7nptCKb9MWtQZLq
cfpE6009qQTS9O+zYTWYRfG8Yg+oLodU3dfuZAwXIAQtEU5wfo27gc7UAxksvD2axHxbgyvEJPIY
dbNAjU1IuD9M22qK8Ow326KQ5JgaOltenfzuILOPBa8x1UhxftJRPrW2A2SmMXeEfReehAKuyRir
gvbAhxVDkfmZgzR1VZ3ntcxO5viJBbGM1A1Js2UlwBVMKcyk+Hrtpg146eokTYiEQCk4ISvLDouj
5k2EQHDqqr7W2+IuPv9+QyptrUgjb/cb16zb21e//rLeeufdeko72o0P5tvl3++sU4HDxjAFim5s
CMIC/e5ewCoonK0teYHI7HGDKYFTdKRj7VEovuFXsk7kqRst+RczvH3rNP9nxK0E181XaUZgbdLN
7eSOsEExwij7KOfT29EqJF7a0R5VOCICPQMCLiqZK1YB+xk1dUjMk0mVqoO0F2XKMmhZN8GPgvSF
5sRk2NtUYhuBNX7vwl8oP6PF9KYuQf0fezb8lq0o7o3L0IsaCvEu1spyiXOuCOP2BaZvxFbgXeiH
oxaNWS8QilHBdIYnCaeVSYl6wneQeunvO9hd0wKx8ZqKgF6T6bRUSQkkmPx4hPvfUPsID49UTyHZ
ZHEFBKHSd1EbBJ9PA5r/EYwNPfBwc1cYkJ0RgK+nmymZh5khms1ApzhQKUdPzKOKfzvS45UjTTsA
gESOs7XMJ/aWRQm1ahKylESBJQOgld45R6aqDLs58nybXUFIcy1K0avXI67SFVF27E53dSf3kq+1
DaDIC1hnIFjBPlVQNJxGmpFy61Ebr1xiGBLP1iZi03wPf3zxJ7cXvyiXiE4CqmMx7yjYfKniyXR0
uKxQTAz6RAboxcm30tYSNdo+MXIenTkPdwMPvWV4zPXKH7vBONm+mpAo/hblT5RCg14dF7hJo8ZZ
TWeIIh3SCX/Ms6E2NXBkZr4Mylm8B/feCFQS74FNNwGR0cdemYvJ7MbraCChxmTeUoHdFXBCDu01
JzxurNlf7Ybh7QR+BOSFReBLCc9o6vWHSQ1/ezKhFKei5GjIQtLtlc86MgXesauxTzgem3RDlRiZ
B6wCjRZV9TYnXE+mbrKpHG0BZbBWqlXf31C4pnxCc0V/6HXxCeKv5FxKZz/xXaA0v+nFFjqt4CLO
3DN0cpkSZANfPG9f1zjfbqgYxEtpAqvNnS2oPvmLcGbwfjxWTimjRd8m9icMYyOZKmqcHHR6x59d
jL7eGflfoCMaj8YdwC8FYoy5dcuCd6+Qw8pALVZra9ObE4MChkpVnBA7O9RnAnH3m0+Yeou/QkS+
o1uc+8qaqkvTUC2ovCdR8Kh9iGxHv6ZqiSL3LHY3v1hqVSTfeznuJ0L71GXqxs6IqZIs8RDnzpsV
DHyiqThNDekTRU/SmsiR2NNLFZpFXKnFWezfxr3MkmLSPsZC3M/3ET5JysLTlM1EYFCiO6A+OsrH
2kc5VuN12tunWxgoHOeGev00bjglq4gjGuKhrKH9EdYWnX8ZGtpfM6PHuIHY07CflRxsOZFGFZT2
Pvo2KEYFOiMEhWOqNAqcnjeP9LjInYejH8veecyGAw5GPJlZpuzT4uYV3oqs3v2zTdLEYOtkswGG
8lT71m8ZmvcjQPguQOBuqO4c258iAO3rSyxO4wiDbjOnbeCVHM43nN5S1mLf3GkiHDaIW6UZvDKp
QscyzvTnEIi2p7cH4S2tIe/dhcoGRROhZiqHPpMfcEeVD1UE0mtheRpEua/OerMFi7d21dk14cjl
kpPgLc1rNZzMUM8bHMqMkpwg2xnLSBxn1wMaGIu6B+thxuBDIPZ+YLJnmJD6/Llv6qfCGKz0C7fr
vr4CGexqFFmi4chCDWXT3cDPg6oMbIsig1Jeg2Mikn5N8TB6eDX2w/3EPxpXC98oDUQwDu1x2EG1
Rz4k8b4sFTi2gA741+JSnh8B/qwmLQFpfsY9qfRjdTCLhszm4H+x5MUDPdtxzHBOKJhvprIlBgjr
TeaWNLDDLEghDm0kwIQA0O0CnQXR6SNPPY54O37L0NRgMwXev0izTe3UfyZUFaX1uDY/br2cqDH9
vzHEsHH/lwAyOp2O+dJtQFRx1G/es5foOWGIY/KH+iRCAUlxvpLo7Zf25+J0AAgFtMVGHec1tQW/
sXTM3DYwWxTqSiKncanz/9V6OL/E+PpipPBfzSVBwMrCNLsQmJEx+w27fNJFekSVH9e1FE1Q6ZEI
ADh4dJMqBJlqQBj5mItzhdZ/AMREFzscHJ3V/FeDtbp0DgMa7Tr8COyVxsKpF5+LdOvCNFMlCngH
mzDJ+Op2yrptoAC/FWWnefLQdqdPl/GaxrquIKuGNREmucz1185mQ5TFDomQjPKc+CIWbMQMzpnV
Nnus7DNon/0lXqj60e/3BlHSt63NxiOKI1dNtECztISOwxT32fHwTC5gxcMUINKqf3TWLCEuxFu+
zaproQuujF4ddnzyGBs2iFCcjTMW7gYg78ZJZB0BsKpP+GGVb8HdHLJBTr+G3+lWBUppvl/KtNVM
mIcobgtrm5IvJJQ0ZPYNWK+jnfDd7VS5X5dAmZDzjYl6HiuK/FtvO3MgQXheg2uHT/rco4GqsNu3
rG6gDeey9FNE0IF9DJtYLu/G4UCoPcxhKTuG+/vQX8E6zEQ+DMoAtYVYghw5LuVh+O5+1yStA7vy
ycTpuo4110mP/kLEpi86rTv7HwSkBLHteUCmP41zezvplOVynjGZy0tMTGaPE9gNhnP3hYT6Gkc4
O3Avb+F/jIW657G8kQ1JMfCwSJA6SmEgP+w+X7qm/DH1NfC4v17AkYvPd3Pa+/EDkaT+OKYIKS9r
zcY1KKb3RP0XpWKZ58AP8Yb2vHasuU6Kws3eWaipxgZ6DRiaOewTQkERgbbKnPztaYIB4EaEguMP
vhm3jlJ/QmgAZQVN2GzWgNHIyukkOD6f88cXjU4Ql5BKKuZIGX/lL9oQyHFyrsnL9fRQgaiqRjGm
EvorDcf7D8xkBEXVFCDTn8ezZfsacpGu503n4lkeh0cRG5Y5HhAIiS5ynjMSe//MUklRNFYphRns
73/q6hJuntseepx8/DM/CBfU1v9Gdg7pi0uf+u9g2behx31S5JM3JFIX+epI8426XpfVdK4TqKnI
0ttcHQGz+6NfdJNTr6MHiEl/NrxO6yFjftTOJ/qH4w0rGYPnst97L/4It/S1kabwFOrdJLdhGIct
Vy4vfXK3eIkhMSrNfBmUoXp8LWC/XsWfKAFXn78tPpRCOHcT9p4wQgB1YcO4KJ4Sbt4I0i4mR95m
BygbHIP9rqecsDL1AQEqtqM9bDOB20aQ5o8IE6Y18d3mh75JGAMLY1Fch276AedX04+jExIM1Z5Q
CUWplA7+bUxTAneSRs4AAhisMcU7wWbK+zfqnNXYz+GMULBFUkQ3Jl63a1R+oMIzqO3UsgcpmLfQ
tK1BoVLH1WBhUiH06abu2HYXZOV7+ehhVn2pcCfgnbdlCyuVR7mN1TFFwRw0cXcSozzAdyT79aD0
osfsP9g9BRguDPW0SwBwgObZkTmlOYQdV2PdAnpQyu1UKSxMJHrnLcYBJyYz9Wi5Ay84gnwK1in1
ETnYRJXstk68vISDs3h9KTnQQW/01+Fz8BmTWwwT++DzVEU5leoJ+di/5OQq9ysiR4tMmVfoDk9k
KJaxbeZaOkp37efQMpSecHgtGtkBg3vTbK3b6cE1pE12q0aPjJkhvQdQgfsuxDsic3+INhsKofhi
fuzgiEkP+Es5L3gkHblzsWhFOkegpNDwj8J7Ke+3LIWsbQQTlaONKjo3WuDFukIipFXzkDJuS3WD
90vOrG6XIaOQMA9z4Yr+zRpzJ5KYo4DCi0BqQ4em7q/56b6wH0Zkk7LGd5IUnsly0sEXWYZDqShk
EKhHKdMnc2cDEA+oqmupTBET+TGHTWuno0StrRBwMhif9RI5nI6WiZTqGTZ86J1luvrYhiagdnAl
i758kgbToJapeuJkK8FQRxIgH7pb8JKTiw4z+DWtMoolm4I5RWrp3vY215RNnmoaC/0N0si5rQpC
IWfb+OE2oSoHgmh26QDXDdo3hExql1GSvHt6YmsUmvV0J+DUSri91W1Qaz7n1nmAtjU8/kD1RNE+
I5eptYUbDN6HhcX+i0JudGNBRLutxHKQgOc7LBw4g1l0IcUctV48acTUVL2Y53Rsh6U+Fu8Ls/H5
2SAb51xvhnxlh1xQ3U+W6gM2zG65cE0Btg5vH02aWcBj4IB243k1Wagh5t7kapwFiwr2Mwk2Xorf
6LGPA3QdN+L5kSG08u/ZIC+5fyV0BytZJm5mvr/STmCj77cQen2aaLt3NyhRdKTNHCr/uLt5CVn0
xNXiYgpCYG4cgunFWIrHmE5Ed3CedNINkegIJ3GOM4yiN4DhUUxfDiuQGKHD25bawAryRvMlsy+9
dV33emrDXdRSepQaib3CDfR3C2OswlcykZDLea67gzZifYnIp67cVw3U8aShDakuGI0OzL6AuAnC
gb4XurZJonoEoHysHhjYlNzNd+J9JWlXVK1n2iNDplPxDlvdovOwE47FrotBp6SLgD5DpMvxIJnX
COfSkUVOKW0+j2BkPoKAJ3B2WoO2D5y9AfdslwhWXzSPsQomaigPU/ii2gJqmfDcPWMa8p6gISnA
PZWdFrDyh18p9mJbViucei5svVOHqGk5UxT4E6UhizEvzenDSXEN+mLjz4LP7JZxHnjTXiz7afZV
YzREgprTlHqcful9E+tfh2ymWX6kjMi/2v6zqHlpSO8mHStFdifdyeR0kQ+/DMTEavTM7Fnw0XAn
3TDmuoLh3vX4cU/CrKs+qotCzSSaotTH3o+4bPzk4q+xffsIG/gg7gSlm2XNH88flDAix8aqVeyv
vtiFM/zmcRxTshuf2luQH33yZXFSRlKQPCf3ToSCzeY/gC9LBhRRiFkgS7rXULsjUmeo/LRX+36e
ZOLHyqQ2gzk3OUVzwAeAQ6EQyIYkcRkFNt/RViD+sRINwDPiV7U1zV68NtJgjkSIMN567KLF60dg
S5jORyPY8o4EZ3tYNCClj9CU+Ym/hm4MscUGdBZTMIL3aQjUFvPnM7x5hePBcI7XsbjI6u/IMUWD
7gzdxePZkOaxJodBQpHsw7YSvzilEIMMUNFtaSdX2QSrU2TjAekGQQzhLf//kB0JNl2NoEqM47nb
Kjv4+WjtO5l7S4CTP1MY8gBf/TRsKo1ode/w+of7XiwJ+nE8KoBFTuhuExDqj7Q3KWmZBU8mTCnL
CAMBvI8IAaPW5lSYVhjJTOTlV4U+UE1YrVtzegVXsKdSOtvDwEwYzaRmRLZDnAGCx3nXAstew4t6
YsSAL72yAgFniQUiKVn80TitJXwc08mtWVuyK2LTsSsMSazqkfGKpUIBmSWudrbZP+KNcFMIX75K
aJSyKBXDWowAbXf4CybWTf+uOgHFwPWZPiPvcsLP9eW7lA1oVZ/JZzFk/QhYdRH5n3Egzd1JdfRa
8kgpRmMes+Nw/jBSU3g3i5RWcxTpl+mhRv3XYkRYvLR9dmbC6OFHzvppt5v0tqnpDUTw/7NrhQfx
MbZcrhqtttbRL+iW4TMG1dqQ2r+WZcgdnUsV1WbBd73P264ANllpD6vWYbi07AuPQkuI25wDIiqX
2yRoUzyAs74/Hj+DTRs9PbJIHUzHHq+BcgO1HKkVMKHICeZbjk10r0auRdL/2EzUxuTlElPrsxCv
a2GjaYAKixxRI3mHRoR5Rz3V8XWaZ5qyMXYveAi8c0oSjqcr6zHyVqcS5yKa0o5Y+TeG1nwk1tYN
Hn93HPH4bS4Ms68DeD7oMyhCeApPE2ZhITGPG4AktevmAye2IuzeHyk+N4VCgJzJcV6B5gi/WpvB
ne4J0L/gWD9mY5XyYVHx9I9cKG2K60R70K9PCESEyD4UBcb2bea1J8Lr4gLnjsvBoVkVJre3KOK/
foQwXU5Z4jHwDb9XB3EXI1+F2B7PRxRRL6wvVmlI8k8R6yfmVuMWyB41N5YAYkKj/X2752OVo7mG
KszCCWUUrvJkrlyxnFOKiyfMBsxINJopdQkqHyIfHTmq2jKbCuWhF+m8/5IKprU1WMEvsqkrRGUC
lwSkbGzrD+xrVhSyfUBEgE+bf10fkqAMlCub4b+Tid4Jr33Me/ZKihBNxd7y3kR+wbyQz0mKXMvy
emtZmtqT9wyn/tGgN3/md9fGTnVwVsKQ9Yv1amTUJCFqZ0C2WoETlIL3EUrXQC7zgxxcrHYTuSRY
6veqAB9SThwYzIW7wDN17kmKU//wdZ6HSp06+T/n4I6UNELa3sxmTmTsjRo+oFMJq/YOq9fPhDT3
dFXRrW0pcQO0vNuRxpIHSVdSQygzYhkPBFZ98k6bV04+4BzKkEAPQESqR2AJ0SO+btJ28Mlw8AUG
9FQsI1SgruEKPPBfLG8oxvMC7PyGyQn+gWg471SXQqtGjl2Gx6mSu3nYpQy92eBL/GQOaP/Cl6U2
CGxFQIUVHOPKCRqTWEZx2IyMrZGLZlSyC/yLtzRe7PzOIId2ekwJHLRZajMGeqf2tjGz+m9aDYol
wFhFWxBbOvsWxN8cwZkgAxiCLx5B5Ri4AM3hQOz081GCje1EngBu53KiS0RXHINJmTpa55O/zWY0
IYGvu651U46ANrcacxxYwldZ1+wnUiSK/SeQ6PoD4W/40Vyl0vJAesoUjjgk2h/0RlIqOH2ivmIV
5W3eGhrNsEtBRLcKg1ejmlk1yATDL0ji8w7RzhiH1FFR4hnWeExaRWbRwU4Xd323G81OLBWxoAKs
JiW1X4d6cg6DRz5GqvC4/5SC3HyACKAha48tZivKpGZLs+RMhhyHUoPvO1U44sA+RbHUz3xy8ZQH
QmBZeRabDoMriXathx2yPUW4C4L/JVU9YYEodOAX+k5WvUPcd0Wl9ws4sGHGEsDdBRT3u0rQtFX9
bvzWF850PG9AXeS6SE7N/vOLj/pYcjsENoVgpppsmFz/ru8q/7SpmeEK/nTI3tmE02BazMitKLDD
eKHyOvxJMIWanlW1Klc5+U/BNmMxaMf6uRUDTpFfIUyytJnNWRcyo4ywFos2y5gK3mO1MsR4Y+HY
tIVjBafapXBNxs6d+VWg344hX2yLPmzMyzoRtDpDCeHMvKOsbwzjxeKwAv+ICVBW2cHpgFxX/ux/
anQ5uxS9o7Ir72m3T0MsyBB8EiEWLOkQu4uews+NfIwWzybBIaVDDT+x+RgWWXyXSoibvS6MJHsk
rIDGbYaFyY4Utp4i4t3OtQrSVFP47UAlCiwi5cUWyL1VebR8ifLMOcAGNSrFyMBBIxDe3jirkJvZ
64ynTCa4U03Ov+/maDlg9Szws44x5oOH/6oyP7zoeS/2kYu1Jo0OxvIFl9m0JSN1yJu8hm+/uz2a
ZBHTkkpD2mTPtzYHabctdiKYzjYALRJBbV8R1CBRf9VxS4kLDVoXTEuWcaDRfPrTlt19R/eLYGZT
CZuuh56vf8b6J/5aCfKyOoXp14wMxpVCo8OO5ouXMLtMczu5kFj8GsNuI9kw2RIozZClq/3IZ4Ta
W/saiWWiXItdzDNiD00hR34G+Vx2pL/P6gQ+5Jlb4jKDhqSaBil/WCUfFyrtOoFVtRtnymucWKQX
wMqc1F9RLpQZDv/UfLAPNVnuQi1W3tUzlayR9obK9jpAbpxUzhfuzhD6T8dyOvV0qLoidnu+4hCF
kvS4tdcm8O99W+rf5RR1v9GGwWZ9VmnbFWh2l0+xzquwMUz/ADYq27N9TzMGYcTi8dfRRUTlCT+w
/kLYTVumTJG1PV7KJoV+iUHPrjLW6+LM8JvJfS2Fzo6aA9R0xyk7HoClaE21n1gMr+h/6a1enVoD
aTfZGakYz38ro8uuL7iThDOQt4dADbbR/8vYTeD6svV5wtLBm4nI/Oni9O65BPf0cUghZ6bsJlrZ
LSe05bpJu7dzMMM3lc9G+7qUheGxyACxIIdeBeHNEEdT23tP7N1vdMAllYoKESNu92pWbe+m4Gvk
sl93ljwdoE67zGYWbg0F3TC+MkPBzpgZfNCCo4qWxn3zP9UmvjMjvdat9tK1f6u7w9CViQ2Ywl5X
MFxRuwG22x1LW54ukBYV5qs2r+Le2dSjxbOLXA9hneirxeAZek42vFxlaCirtJatwcj5C6J63Th/
1DTNnS4XyVRu+iHux4QFfuzfDNcHTWresMfiDr187RPU5sZpI/S4KmInSiDRsR8hGZGpuG+ZxWt/
Ya8sO0DBXPvc0XrAqUSsook1BP9Zxp3tqhO4pYWyASmbBdRUVXnTOHq4c1X/Pl0du+HeVh3M/Rtd
4EzNlumizNkJWr481/eJ6Mde3N3bo332ogPVb8YFg6J8uC5N3k50/czvLpErIluzdPgXOYfl5MDB
t0mImV1770c68gVkArnHcKq8359ghJQ0YuzPdM8HABGKXHpakw2HwR7ajxXnAnEbBo2ObpXzRuPC
o1Q7ou8RsfAB6ozzNWWgGT5mfM9600HT8q6i/kJe+xjLOQMhH6y/pPc16cCqVaOy9mLDozeN74qp
12GwKL7hXlVB0FG5LgKITQlwPPirJOtcHsOT4Rk+KSScsmqMgoFLQreNcZ73JzQBr1hphiLRWvgo
zHjxhg7eFLpA73zRLx52p6Hrr7N2II/yt00rvp6qxg6NeBISqBh0c2NpqPGwSfQ0RqcUn4vY/yEI
FInuHiFVd91vVLSYWuhYe/4scQv9kE8dGs781xO+GcXyJmgxH45qYlKRIJjTPM7OrRpkmpRGYAco
ClrO4hXuMZnCubjmB8aljfpqYtvGY6TPoFHSNDjciEiihVFEy96HQz4ilEp0OzWcIYZ8Z7eFSkLG
EdQUQPgVhcCJMN90Rb0SPHbpE8sR8X1B5tZcHtPj4hfPuhqwhwf56QxpHZTUZ/yBB4WfmVatrB8m
xaiOAQMSgM4LgrV+CNZPy1XsFZO+GrJ38ZsIk0SrKT0pAwwAYaNhJ75ZeqdVgyeQjxYFWUpG1SfI
ldMhiqJOGi0VmbEytpAwr60Oq45mU7CENdKWHLAJeI2Tf8gbBO3Juwgbu3no0Kyz3g8c0sUWeKtJ
2e+JeVzAey7owajVvc5wG+XivmA5i6kd3c/FgMhBlD1eNfL8pdYhvg6+UjMiFXjODL8URrMQALqq
nlTsGvmSTLFgeIgKqwNboJOXP5VVS9wyuhiCsyT6i1S92EnKduwAWdz7NaEeaxJ5mMgR0khiA0/M
TXssEQSYVuPt8tdvns0G8OLBmgbDyCO3adrGdqeJUgM7EUW6J7jUGTx+vWsksE0CVk5Vyk5ojBMX
R/lcGY5uQyMt8kKH7k566Hxa/hcrSYMQm2h5TxXz7h4H+11KNzGanezE4ZSmlslonv0xqkRGyOUH
gvI6yPQIHwh/ec/7r48iPW7sUzCzygJ2u8pCt1oIa9eQXKzbUwutjE9M6dvKDigsYIvnlKYEOjb9
SpD0Psfna45Ffaw0UQRt0/4alBbqCkI7SEabUxgp/WXQuOvP1FHVPJoTAaF+XjUwxioOGgTfm55J
XkBvbvJ/TXk3ca5UdPnrNdTTIE6YN1oLt4iYhGpM4fmmb5wHqpDlU5zAKFL0dDfBNJxyUnnMXLYM
5YD4TepPNm2EcQPZimVT1CkTzcDUIgWopgouGz3zIJSzzHA+IPpqjiIx/c64sJFcy8D1kko+ODAN
xRt0Ix9LPgQqqBi0T7Yr62e1OM5+EERIaKSPvuTULcbpLRwt/oOA5Am3hMhgKTyHHWoRaVsn59DT
ThlvBpiQt/FAnamSNmPaAmSGWq9JqzN7drDfbxRroQOS2a2829/8UYT0xv2BeEu3rjlnGy/bDETA
Cna0KRJAKZnTP2kut+WlIyC5X/GONFxszM4T/Gfq2tWYqs62wY+UaTeMcYEnPZMCRnvyyRpBjMGq
P7kXRXj+IigK9BQHRzIczDQ0FB5Z65B8EwWMdSVhPq6Wew9Mh+1xAQP+KNZW96Tg0yDinEmI8iNR
zXWvm2y14bvmwbypBd6gAg0PiOCjc92pph/P0oppBnZ7+uxbvDIcwoLw8OG22G57fbLZsja5PXmF
Cw6byfBAeTDgaIL+wlKEoicahhGGDMw+3OK4BgwvhKaO1vwLFpvsij8Nx7k5XO3NJLRyIRG4YHMV
b2SJtVZZ3DKB9/RmFDNE6KnWVR2eu0GFb4R/TfCy8z/F8BbJxRVX0D8yUCKE8kzrqsLDbImJSOJC
3uShkzMS/wgpcHI90/CWIlH5Ux+COulY2J2mbvsai//Qj6QTRZxYuflUKdZgq5S82t73jMTmvIop
iDHAdeJ43IcU06e09tuT17tmZGduxWTa0qo6Wej0pOPf8srXu5Uasi4Q0dlbDy3VXwN/6gWoDzZd
ih8E429VdqkI4Aut2y10bRQ9u7PQGdvX+OiVrpZQZiWM3Reev8jr8wsffcrE90rlyKFtYOuyGyb2
3CdJ58evU29oWV3H6K3btXxxBz04WjE+xDfIDPEUWHbQViPwICF32JmHwY+PNEQeJo2kYU3PHbLl
la/fr8jrepGM+FB4yMkPU1ldWClKzuxTf5SUks1eOx8cYxksPByUeKd+QgWljyVWY6wX8vBd5611
7EwKSgA/oEQ5STNX4OHIqyvv4EEoZM3SPZtSJkhPPy5mIQx7MYPrF2ieYiOzr74/poi2PBgtn4bY
5IwknK5BtAp2foVpc1D40y+bnr9Zf3MrhfyErauw/tToBGU45OSJl/yGzIAwFndaWEjn2y+LlSRk
28FeMFqbVjO/MIIhvbuc0XC4T+QlGXPE6nEVNytcy4qjBqhrH0GOnpylEqjN2Lxi7hP5MgA8bWOd
T4y3T8pyRws5VSEQLRqGVm2qj4Ex3+RwjnCGNGfj8euFuF56NWk26fvmXI5inDHaueWRTa2BCaZc
GmNqvC/kHVhevviO8DpgOgfUAgeMSA2b3hRd3CuX+DxFaGm42V5iV0tfx8jHs5/EtY7eXpAqcPki
i/0ksMX+D7MKa7H7iaHp2/+lxiFp08cdSqboaw1JaJYjN2n/7nEoJQyNuJgoQk6uTymBVcVCNK4y
nN1jb3EjROe3I+1rE1P0NSIk72mK8NTVKqLgd5AYzig180w4syGA0qavnnmPwYYjtzFne3npeVg/
XZXKcfJ+wzWvkornLjvDBAQhDmT46cl4ujPumntv7Q8uFZYUGZLZRJw53WQZeM4n3Zap3/WJc73A
oJ8yUhA5fOLrzNabc8shhz6RytddvYbgz0OOaO6Ms3Mujbt0n/+evBjoHkPshnlJzOkViO4w3xFV
t06IrtG97eOtK9fN/AqN51EsuZG4wlub/nWSVoXLbPMl1aKHD7cS7GHdhZbMKYxgURrm1rwLeNRT
IXH9Zmmyl57WuROcjNp3Exq5oRfDUl98wOONzrdOMvujSsrL6fHlen0NBXnaOerAH+sFOExvTQ6A
9/3KK+MqgMfHL3gmYiWEGbR060/Ac9jrMxEp7ABp2CF5+RzPkn7Kn4AjZABxbUYjyINaHROuBiGW
Zsh+bWjX1D/QblcNziGoEpKfOJorQGUoN+/7CbAoYW6+P4sGbhRXX6EXOXKyODEipxcd8ppq13AQ
oooPYgwmmeZd4KAqPy+FTDY4IMVWJlbC0gzSxJWSZi+ksJNPmDLLXnYO+vCACYAMTPQ8wAYqt9U9
DoGsdFtBiSGTxBhBjlyEhUNnCjJ53ZWCz7rl/NmoxSb8yvFGbkC156H9NEIqXgD4Y2yYSgQagBZX
IErf/tBLNyiNzCmFM7sn71gXiBtAv6bDAo2CQ2ebT2bT30TjXpeyPM2sxIW/zSiXCKCxDA5wEz5X
zJoa5YSpDxniQ2hjxC8zAyLRd7yaEmZUHZ0qm6Jb30SRt/RhveyrSGNGUNNd9ggVm8H58jTYprPq
llihSi21JYXu4cXR27HR6Nako21XTfoFidoxmVS3lpOqbwTz+yqxD2D341nxMDFK6HGk3dmc3Mnp
6KC2bIJLAmhsvoorabw60cgDqQeVnL1KDAOnG+EBnSr/SfT/QEs5VBreLyj48zlMyvbF1Xpj2x9i
lFxnJ6xl/ejXAzDaaJmFfrOL08LZuYOFg55VPtfiC7C673UmIREiHvAZqqUs2oK/SeijDHPw4tpY
/t+5QWak3UP+An0Zwzw9WB8STAx9Uh12LFTpv3MOlGZXZ3CosVgZPsM+fGF/+kiwUS1dFuoT3FmK
dGks9HIhImTGBBRYQn0o3/rDEWbphcMET9Iic1yGEflVVPn7COlPOU9lSmXK4Kxk8g2PRJBzRzNM
pGXcyBuGUB/LYTMdjRM+nchBs8yNyrX8Pz36WKfcvSEx7/tz1no6wAuHHUKA4gm8sVzz+C6gkol0
GTE26xgqFHgUc8jUzn1gVczxnh2+rlilzuDG+r4lvBqBP/EzSiRzI30xdAoaf4FyxyaIet7q3HwB
95U0e/y/B7C45UWR/QZvijX89ckR17yPBxVYAc2cch38S7ia4UarC5X3kGdLjhFIHAA88FzXFrtM
FRrQNA84x3lj3AA4h8nHobc3qWpF3fVeXbeclTpNF1SzetUBAAKS/z1GoXJ0k+Ou7fO0VBQENfNz
j9hi4VxFxIgGUlFPvwmU1IjZKSQSP5mQODVzpiO3Q7dpV37BnypIDcyRX5GPno+DvO1yMuH50dgt
xDkm+q9kXLusY1J0pVYtD6YpF88+QA08HP43rJgXBUoOyQDd6ptkvJqoLZkQ2/WVG07fIgkmw6wH
0FxFf4bevFzc7jGbN2bBjS2Lg0goDRHVI56ARNpZ2gIbELBalxAa4HwbKIeX/T1lUWUtZzw9D0+u
4Pa1kOYhNZnbZqYI0fCXflDwXQbvexC3zhL07e4ZzdqGcSU3kTZ2Ep5Rlf/CLCzby7QyzpC/8eir
zjTRSMHfGWuwXJdmZzRHF+FRKOALkKRQhNCXTcOuYHfkBL24PmTTBe6aSbvCV54SiPXZUC6mbka8
iwJkGD+4hpt/bijBLjvD49wK1eWuAncFwS+YGVxLvFiDQxeJSqEeYr80m8sUgE4TPRj4Coj2YEjP
DwLRB28i3AaGJkiqEeXnd7H3hPYyK+gzs289FLx9uYVqm0bfP+OGJm6Q9uXdtEzzz+9VqUywy+dO
K1vCaLldVShwhKBuzoUDdrU2JIxqlqXrzPqSR6/9IS2xMNQpW/2PE3v9TEo26INCsJyp0w38WY1U
NobBIKx0vtvBLja/11zPZEUXmf8Xu5NVYmVEqUQMOhQbjMNZQ1zb8hhy411DVpf+h3w9aL9cNf6R
GYzvjoHnEliIah1DKyOeN9OIg/yuEsE+7FEbNOPvUE0saWiksTaDRQRZLzvgXZ7oKtqQkKSwx6B3
3C87fSWcKGCeM9xUcIUzftuFAUOMioBwuZTG/HKmcTiE191pFJQMoYPuO+b7QV7LvHCfmrCQjYmj
uzSb532UIP5ETd6LE9z0MWilnbnviAw5npc5FBQsj0wzpL23+4UPFdblhFuI+Q4B7HYAkJ8/G8Dr
DTN0laHp6OMN7kU+5vm28hZYwxMcrNbbYq+qkbzEq08Zjf0t6VHWQAJMPTZqubcL8f0gyuFI1mXQ
sBe9M0TsfJuCAWp0j10E7sbcJwnk/BfT5VIRqy0XHSOtNOPZ/F8BRcvTvZkQYq2DgUYdy8jBZrHr
tagG931yTzIwwaTs4hIkvenPGrR1VcBc+I017YUIOgf226R6OhgYmlmTsua3jhGqH1/XUvbRUUIx
YGPyvGm3VcYhDjQzuWCR2IJcU1oC6b0xl7t8sWSzcWO8RSFAboWTARkqMTci23cyJrMg9IG33Pu7
gews+dX41wr50HkoJlypYYaGjCqcAdSrJHZfDGJpmZEFnaI5G8ArSGC3VNY429cOdaMbEgPsC03B
TAxLk4Asmnj0aytTvan52q3Rc5Kg4JoTwZtr7lCXPrLps9HYyQ3KIBth7GfyzfyL4upvOsJ7UZAl
p+G/QSPbW+wA2LnBbXZ0rOye0Fq9ITZqcakuQRh0d+UJg1A4lP055WUzWoFUs1LKYRTgKIOX8zyj
HAY8LG8sNT8ohpy8D+3YGBIhP+Mr9JnoTM1PnG5Kbt/WlJIkBEGpFBD4neunrwvVBSlo7/2JFdFJ
ux3rdPFW1mafeJjZuq5aHsxmuQwXbaJyoXOeCoUgZZvgrut/X55RA48+JVnL4g8ijyTNyK41/NAC
W78v7r/XiAL7Rb7RmW8Z8wTEEnDImClEQVllhH+pSAap2A1FAU8mJLeLo4H70msgQ8mJT387cDt9
BTEGOHe/2/AChMzzsSL6qHtirc99qRJo0Gf16tEpcwxwsNgmHSkxdyeRxzb2eJqeuCsyC5T2yaPO
GdgKXoDygUimXdCC+CHerhvH6N4Ct5TmFqeOTKRAaeI1e8Fc+dTX8AuFe4t+T2wQyIbMjZU7UvpO
Jw1pTlkvziOEFe/qWsbdKR/Iu5jqr8cMomsvWcbZkeSZxdLbZjAcPK6+aydVp/bGtHXXdkdRW2We
OH/JoTr1EAcyRsAXWabNL2ZsHUXSUvcQKPhT/e81d4M27VnrbARg3+PkVgHuTjf3+1J07Sj+rLqs
9XjnSl40z2ZukCuHJCFPy+eouxAsXfsVCDY/5cxBNR98+wTmuHQ9nYdhUyZHctnkTafTwMGYN7Yv
Xe564BAHr0F/g78LftzeKPUnfkcgS6QxbGLwOAv+ChZ0rV7HlqiVo20gWNccAh3FHeBk3y0Z9ZNq
+bdvpi6S+RR6QtaH6KvQu2FDV3pqvDrX/lyx7OKh4YB3c/KeQTgUzPfTsrgwFMBj9MlP2f2viKIb
sZjdclnJotKmx5I0GjR3sXykria6Rjh1IhqPpy1/jNihUTDuPYnTpFlR492/fNtTDHtxeKd/GWpb
pPPt1dEFy2aI946nJouleY32NREEjVV8EAa0MrD4KVy7TQIGEPU+45TFg8FGLU7GYmprbRVKsMyh
9azopdbGZVmvT+sC1EdRcwgYsivz1UEC8/8u/STQlwY6avUe4/yCC66tVQC+Er1VN4Ra9b4WT42e
zTkluLl6FeTb1tZH+mK2NBRLezG+wArF67T5tbs+tfQbLEIc6RoAcoG6O3GqHT1C3B7WWaxbIpT9
9lXc8yqvA5bRyyJWsPkut83KQRhfnadhx2mnTWeVnGqI/hS1CX4r1Vu/wxteIQ5+J2dEIsewQIpI
FQ+G34mmMWH/HpXBZX5j9E2d4rMBp56gVOzkRVSyeyH9MfWPD1PpP7rog9cZfdKLne/XzX09QOEG
SdopNo6pAyt4fFaJ5sY/vMbG4hDZuRk246xDutu0q7D7i/VNKJbcgzrQh1OHiGAu5NzUQWWPG75E
6e5t1aAv3Pj/zKzwrCXqGbbNxV/HHpKAXOTrwJ9ydcxlIySgyAR6Sz6yoOT5F8ei/feMjLC0uYS+
zFgCW2CCyng0r7pMVKwGxwD1eUJau3vIbLfOnDYVsGMrCwjNi32V/zBz9X1Q0bpgs3aZiJeRETk8
qDVCfQ2ZDgz1Pi04BXGkYUON6xFxp4RcE2l+ueLxKdzdcLSdwDOcLEg7Ib5foCONCefFI6OW38ae
hHYqNSIxfpdYRcF/ktlJERrPHjpX0U2jrW4vu6rM0ixM7RUCiawUdPz/yuatajqnODO0QPbsP0LW
IBK5nsat6KMPfIplf0vuW4iFkEK/tyxo3j2uhLLCiXD7r4thaqfWC2MYf2xg0fYC4NEZKsHZlEhJ
oLMZ7raCz5PpANnA4/IihkqPzvH8AceuCuy7mHE08ISh0L+1HrH//srVZMkAabYlTf7abtEoLe4a
vGJ54MsrZ1kbmdtn6vQB6JFf2xqNpuzO8IDuOZ76t7JuFQhg4DF2pE7CTk8bG5ou/nMs2przFWdl
b+GcmoEdY0QttzP4zHF4lbbjPJWouOeF7fDNDv9m26xkAq2ny9PfwG6yE0UlFAdKdyWOnO9IYFLF
Fbop3wSig/Phq4prjVK2aITmfguqt0CkZUvDxllPTnk6+G8JlZcxwLIdxU+s7Al3i1cjEr+Txa2N
86opARpkmz0xgZe5+3XJaApNSXSPpvAli+7d0N9YbafhAGXHICMFcVHm6ez48BZrpLz7dyST6+Rg
2Knuq+Ewp1znaVixXmehW8CN60JdbBhhINyl6SZ5Z1d/gxJNHAWssSNxDjBJCaeDt8L1nUdb5M2K
Avwy7NNxaLRlEykBVBTGNiScOYs0qNd/WEsz6UJQaY3eqeuGamX0TQaSN+TZ9OJl3oY/GUY9dgTt
+tG3kAOQUhBUMez71xoAcUxKHyvo2T0P+jnTH4tex8Xgbd/AV5mf/OfcPDXmA5ldNk4NHXJ1yq4F
WRORn8FvgUgSVOLHx09KioVcbSApIih4jbXmz27f0PxBj8VA1wgF6kzy8aOTtYtP0wNUQJfqNAUz
SlpPu6LkNRGasI120IgnI8ZHgvwZVSnQF87f1rzsHkdjoTrYNWWw3FOXeVNCqZF5D1n/qTHDoLcH
4PNP3p8OrU5wO3/wpZzmDL3EgnSJZ+ztaPz5Jyaky18XEEzz/0BUQKC+JQ79jDWr2FD2o72s/T4l
DI4pzCoGG/8ZTGtw3ZdMTqwyRevsbHiY0lQeO/q1VyPRCIcUJkF5kMiXiibq2V1hAnIlEJUZYF7y
vQgHVaR6NaEIM+1oAG7wsXYco2AZpCYyjZAZJogm7ijogWGNgGdauX0SQ1tTter/HfzeFklYcLF7
oZifH7b7WKV5ISFVHlEOo9erYMOOGZ9E4XCrxHB05RYlemzQSDNtN2EiYhLlFq/9ee8/FejI7cE+
o5MPs/CpZJ244R4Oou8dNF/CFyLLcBUhNEyDzG8Rll5JJ2ONFwfgpik3vB48DaeEv9hITSM0m9Lh
+4thC7w=
`protect end_protected
