-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
y8B+y0pwbYXDAGiDt+WLZoy7juqfOT5OIJ5iyt7Y5gfsjQRBwElInnTbwd7iBy+n3gZvNH781iPy
aDn36jpPVlOesS+uinUeZfQ+5msHfWPziH6thq2rC/RswIwYGvLFu+8jlyY9DqLQtWK7HkEsocSZ
odfvpT6GKdr8ILqVftAke3QXH42NqF9tI/G31cIMvYc+hz52jjyFIdfg63JxIKU/6kYCUVl/vUDZ
PR8EYkvwgCcmHqysvDcOSgUP1byuuPmsOrPh2HVniVMml9PN87+Q8+K/qNjXB4LCyZBUihmko7NS
+dk/Z1/e0/ck070RiIRQ0FVhfVm6TFIyWCYJEg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
AlqNUhyrKcC7mi3xjkjWOi6K6sPOHrbj6erP9A1K+Do/wQVQwdtqe0wpwk+jDtPaMCuNFCy7O7cT
4kfOSnKHEsHJdHdnJUyrtcyicaaiMqviyxo22cQrPElX/2sP9ETWazeO0fronb/XxAzxCwydi2Th
yY5Z11JHPrGATrgqiQRl1PRsiXRzZP++RGFM7CFNPfqjhoxJUQiXKk8z+nP1FPJImkND+znyDwkT
XsoPoWmuPSU3TAEE/7Tw/UOpNAnU4pWDb1uXgXi5FZ9tT7d78F25yTnJyt6FId3iWF8dNiI9oWzW
66fr2YHeYf7fvHIDRcD3ZILMvVvJuD7g0r13brh8jkkFcG3H62RmzDGJi6RHqziYzL2KM/O114Js
ds2lzejyontNv51lPb/Bz/E/gm2Zf5ceELg+SmAXo7aYUgRK2xebJHZUi+tqmQ+bvdkjcOkXjSc6
uvN/35Tf2ibPflo/+MzCFC1j+t9mLs8Etqps1TB4wap4/kOk7pd7uej2VWXjthqxu27Hq8mVP9zA
kMN+e9imLENjZT0HZaWG0qHu76lk9sMv8zVsP69GU3lSZEUta2ufVmH8Uiwr6nopFZepbaqyQ4/1
3U5S66pWDLXr9cP+Lct2DKAooPwkjTSnsZgDDkNK+SOXaOJ7Zs1OD1ZmDFwJ6hbx9Y9rPABmF6ex
xvL7aakVTb23V11ikqq8AVO//a6GE/Yi3va56cFqyGsvB+if0UDLSquWiSCgkQjDDS2r82ATsguW
0S2Vz9DVuTR9o7WjYci/aCd1NbnFYfoBz3vweQR7CyihR1bv/kmByRMfVIHIHxniQRugmVmZTpz4
48AZyzKXcIA0NyKXvw9mtcwWn2xjuKDXohrQiwr1/88smSu8DpGUJXB+JCfmCzfP1j9QxbyuNC+z
S6Rnrchlz/QqtiTJhK+/C5AdRQt4liElyANMWEzkErWOlXPypvMd5AgltjFPDGtU9c44j4cqRoZI
mbSBoT49DjFWIsvbQ/XmnDl3M1D21VPH2SsnQIxPJp6hOa59Ht0L73Jv4IIMvubziI26+wtv4/SV
Mk6VXeny5Zn36iErHEJLT9ev1v/wXvsKh9aIDycR6FYRoiUagxJrWNuO0y235aKhKkH8RpAa3yHn
ttx8wlWjm9Ex3ZO6htGd7oKxmzknpefyyQrIOHqSUmOjB/2qMLIviYbasQ697HjmpDAsHwNMePMV
AEHraiizbr6sQXdA7SSg7YY/REelgC/5ixMxxpCn4LViLHPdHa826BMAP1pYpG9TqjxKTMfbC/Yr
efMoNT4+fnWFQ1VTA/2MroMI4yHiRnvWN8fdeTaNmQUQTN1kYZO6xIszsl4xL4D0Hk1BSfZ/zsYX
tF2+K58h3SYhwZvp02amUHZcUDukVulH6aO1rqW42QRVbDUPAeF6G+6676h8Z+t8qRegTS0cTirY
Q0h8y7O+pHTwLjOvNexFBilT7xBXXuxGVH6yLI+af/QruEFil29tlkQCczYKgrOBcjsC5W2w0mdF
jnICeqDZ8CkuJUoN0jLRbkG1fAjRpEZ3poAQ/TOKpu0eP2RILYY19Y/NEtCG+0ZJgWEF0cy32O/H
iN6S/7kWqCVuCTKJChFN+Cu9Jr6uQfQ2xgNZAIBLqdne4bh2pF1+tU4ZHxKYG3QdTor+NLuO5dIs
5vzsISMjmpvhwTOZpjd8gViSTpW2sP355oUyPviCfDgA0bxMi1MxWu9e9RzdIJ4hzPaDwatGzO8v
N4nvo3R817rs5xSCanqMCEW45W8fc3J8w9da/oQ2Kc0sBfUE+GZayf2ZqAZ+MNFRF/jfviywnHVB
Aq35KFVf4IAnle+WQkQdd3yUmsmLITMtUrT/m2qlQuQeYv2uGEkuzRWONyrEY54bSlCCXWmNNYyo
ksmodZG7R5UuKTe2ADc72vUAvDKZEdUGhNiMp9bH8dPDvInpRuRegl9/XZfHTbuOXUEmIvMxsphf
aYAc/lVVFUE34MrPSpQebirrOV5wU4MFy+Eplzin10GrU7M+x3P40lACIMNAi561OwhPzDgHIgtI
sj9H6ziszeI76ft5eYTFaUbbORGsUD9s8gkNLNdTFqu0j/YC02Gjpqn1/Wal7sxg6l4l90XPE1bj
TJsi8eiiaUSoYVydG99XFnvlPcFtPbY/CdvPfNOzWmjmPlbL9B3YDj3PPxcwgr5UBjxsFPBzDp9w
2Tkm+L7fr8F8GVBG1wOQUiS7QNTdiutd/z1flAzlR+U8T9j6Hunj8F4Lwsxl7KweGT+l8EEEHrha
THVoA+T2iRwGshm3gYAWhb+NLEWuzqdXPzUzRsI1oGuNgqYd+EQ3EF4qS7ymvXy53WO2KT0jxQTk
zRM76I4ntaEdo2OIfqtdppCsOE4p6hlOu+eXtsebZVU/fhPF5IVVKoE3AivRpPku9XVGQXD+35gK
o56O+jkNCAF3zILD7ialCrKI2XsAVCqdm0rfOoubqR2Uo2KEcC0KD/09V+1w/Iok32ETiyMbAuki
f6Abl5Tws6ZS0BrFOPv4ZbsmUDs4v/e6+zDvQ/RISMMx2Abvn0YbKuSOM8KABbcTxjYCsbmUwZqM
HZfGhdxuDZixS+mlsUFiPXzAOIaQwyKZiJYnRGMY1ptmYQXh9O5T+eNZ725k0twdZ/A+CcH1O/rN
8tWVSOvcroMk797YGTxO0HmXi2yt4kC5B8PiRaiW53HEMbWIGT5kdgF/uEgbhDqfMWcEvQXSIu4w
Itn6+y8cJ7aByuHfvivXmyYc1HIoAjMkZiJiNEjdBPYZVxHM5pZCK97C2573Uhv1Qosgdkf1ntiZ
DJfYLV7h6q5ZGt34rAgLc2GIYR7qXjVdaBeEZos05I/NIx1td4ADiJK6N3FKBhpbk6H80TFOV1GT
uHGS/whRSUEZQogIO8sdxcqa3+N/PRcg9ImnLX+6QIWQ+WjLcKSNS4URMbsuVuWcoxLuGZ5ivRwI
fMmTkQ4M20Ek8xBMrLX9vucdun40sJ6wp6ZypV6MXPUcTs27kc45VkmBC4fXBa331qTnY51hnmrH
iHKwypHdNKkni2rmhJkiswRTGIW3kMA4CibQgcD9oZ9Z+n1tq8aacwSI18i9vwyAch8Lg07aDUtm
evHkXWV5fkqZqiE2sZilxa6vhMfOEYA56AwigDpUUAzEmUlUlthTlWHVIyfo6V9iESDi+Cac/boP
wt/++KeIILKgpDGuq5yorPdp1LpluQCGA3nGfR5JDX89a3YNWgSrYTEBjUQax0+qDO4mfDcmxbz7
zy7ZkKoPcshVDee+K+OO+VRLJSuLIilHZc72VZmlMzWFqz4xBN74zMt4ecCV7GC6iRKTjpnaaGKw
T2tpR0EU1d9IPlSBjug9XkkjGNHt/1nttFMe3Of86U11nDH3LTqyYpoGxH9G3BGVNzBwbYrQt3Ui
3Sh9WF3YKWssCTV6tXBBwCUdI5KhWg5zwLpnhT4FKKvTxL3Hk4Tk8AvyhB0uV8y3j2KaB1R0VZUI
NhwI3A+/vT+OT1Jb+TXPODighA41jEOTXoFLPqX3zYLt890QypumC99vKiUaROU7wOqGiScqpREf
2gHQr9/jGIYuYwQ3ew60kJ8zrVJmmN5cPL24JwHsdSscik4MpsNaMsfHdNW6d5MzS9pUHZcOnX23
x2EDJq9H/W7DAgUVjTPCibOfHWsXRkO0q7N4rRLwQo+grq1mCg8snVpl28CsdyO6ZERnUBkRZMan
eIDEyDK5SxjMlmYkxX56+lj1oDHnXPnPc5bHxji8Z3YNuM//2E56EJpJi28GsB+xDIjWUOTfOMci
ouf73qaLc2CI3ooM8Q/uM5Rs47AsPIcUO3ExLubMV/X1dmmwKknyegV25HCUUEtX2sWpJyYKDR/a
lwVPGuzweDFDkY5HBELhx2DC8Ugxd5DOzkkHJJRE+yJxFCMylwOKJ7FZ2Ca8xmd15y2jhawtmFaR
Xb/2AErRu6AUO7HDlhICHM0fqfQ+BBlQ3cwCZG8k5LsblJSwp6SoAiQz79lTYgUf2Ym2bPkOEYRa
0xAeqSFh2/1A7XAv/knUWgrbh8Ez6MHjKSUfIunQn4ujuu1tEWmb+R1q2KnSFasL6pf0b0W7qoHH
GiW0hFfjInQCzEXAiJPqq6gIiK9FkFbXBDkjjAlxZpB9gHwpHny2i0s7+fTvqXrdH02eHPdwgBzO
EXna8FAj8BPLkAMsjzOqL8fBTIy8PQjC6/Ql0957zQEqZnhGN+TYf32GOL9/fuB71lb7ygizrBIF
MsYfaD0zZha6fbdIfpnewWyEOXmHF4T3zJ0Oa6022vIAfVz4TTrqB9SnFSN2Jg6F8AT6ZY+2Lt0Z
5xMNN+A8ehT+D5f0BGilnlDEdY+1VTeh5pZZ5MQpNn8Fyz5DcZL7Bn9A4hmuxaxJr/Nn8NSpX2it
HdFXtmcbanqU7GTsWLjQwAoegD5Hcs2UcCTn+9cEakK8JuDlRARilxhvPMSx0tldrLkJqtAp/I3z
ro2h97MIX3O0aLgwP7iI+sdzXw1gUkvZ+CP5of5MWEp2cZLOqaHdC9QaWwNs32fmYvsoyFPSEmFM
Sc2zkXXrqoIgECPhZjq4Sfel8LxZ2yI1+YSdFLvs5HQoH7fckEbezFQtfOFHMq+jWfnL5EpZH+XD
WH/sEhKZRLwdb/BEMaVmKiaIHqPhhg8RY9crww6hZCtW6/r6mEeb+HyvBjxxwTLxAio8iMm4m7lh
pGtXZouNqxRyS+hohgfDPGmKj4+MTovHBcYDWqeTAmGDl4YAsz6KFK8zRO1WOBK0fzM1Ciy9CofZ
aWnza5Wkhvsd6cHE8aFLmHcxB0O+U9JQxxO4Wb4jq4UQIxUfYjgKKXuCWK+WBCGP+IEhs/X7jRwi
1O9/cIi7If3/GElhgelsTtMxjRWIjw8F0ZDpIKoVsD2SXO/mSHYhPtTRN1VLB9Uz2cb7u52hgK4H
ExpcSncLKBMTPzhlYMQEO9+3q5Dm1zCWiihVWLp7jPcJhG9gPZ3EYJ10p8e5FUiqrlL7vhLzEi9e
YKOlaIqBJpez34BVX/lklcSjQy2JmYHQKD7oyTx3qwHJsIud2wfin5cBgzP7JubKRj0DTfGYUtNR
geePTFdnWjLMwlFiWz93rlEyM3Wr1UkUN+buKmqsewcKyapxFfdAH/SCefa/Qq6NJzG3+pGAioy5
pARMYQ29+8W498l9XIu/uWe6vBlgIL9aXyZTcqzcWO4NJJhIbvf2XkPMia9U9YYdDoH/pe68H5bz
36BhB4keAJrneWq8Xf8gebrJXX/Hb0F18MclAdVfsIbp/bqk7CWqyN8rUhvGLGol/2U/+IDN5Omh
X4ZA/KOBggcII0PQY498nX0ayQgFx8Ybugq3QmbpuIS/6wODZCLBive18bnkco/nbV5t9neqdgZJ
INh3XnEoLxvTrGShn/gQ/loa9nuwxmkqDvHs9RZENWsscSNJoaBtB7tb9X+ocWmxJ/7TLgbHIu3j
vH4Z3l2O13A7d7Zd//2p/9X4D79WdmyRK4bN2OEbQ30oSdlyiiKi15ouoARSOnBwpZpr7i0dk4vq
YZk4Q5BTiMVowI5uHwYHy0S0E28bY6TZMWbAh9xuaPaV65VGQ5vN5MURbiivhOIqtlP/ckSWs4Ja
2B7TZRnk3zgO8KYgsWr8w9XuHw34zgXVMWiD1WJDFXQyEY6M43rNma0eS4qgjlbpcEB9UeOrKUae
LKaiWsgxCIGyy9eP5W3ENYk9C0nh/t2ppjvICpd/b+lze2GFHU1M4XZlyC094XzTkr3Oxwf+01Oj
h7aOl26bm7+aT5PKYGisZ7HwUt83JPyZTWW9PFmYIc0mCmM38RW6PQYYNC+uM8JzdnFcktaMkNvU
MdSW6PlhKLxUtLKc9K7zo/GfF6itm8fMKbDCina7K4QTmmKI7lKB5XXc/2urtDedoywPbx0gwwIq
125Y3D0z8UQS0Sv1UwiPuud/f72SyXtR+/L0qgYZoIkAHz7vjvcQNM4dopSbmfCV8c9ozNaZ9r5J
6D4OK9DV5SXJC/ZVOweyGu9YD4PdJgPFRSpjE3DKg8PmcCEsKm9bVgsQFQhlLM8hlM67N55xU/FM
/TLG+jhMKSgZQKrwMrBcxpaqbm4POrcYbOnNOPiaR2tn6dnvm6GkNJO80MOz6zFTBdQZu4L54jHz
f5Xl1Je0sEM/vaBgFwIU7i1C1yzsdLJr3VbuG0OPZrA0XyFGmOEjFJkK7kanmdx71zTfl49bHVdT
kYIrjmBI6vm/nuSJoxyMUjKyUMWV5OxluEADUCJgxIETN/NRjnVKPSOEhXvqX5qgE0hBVet7q1rr
0h9DcHhynpNhD7X4u72irj0uXg+Gc662PI18KPXUK9t3Tyilh5KySGPRHQS0n16CrsKNFbXAgkiB
e5RGKviqqtxRFPg3gA7GC2lzvI5o1o2zjN/k0xYWHAebA7mV8/1O9lMh702ci+NfP8Um9N4ewjA6
1iizdxM89Mks+Zc+95pCOmVeD7qu0Ky5i90WcbolbR0GkyILkhtf/wFHLMpEVukafcASRCAPPl6O
yHZax0XoUh4M6PNgmEOFS/0jBhdd/X+iez2/28dKoz1JpzwlXXhI8ZbBFyBXRnPhA5itLtWKMdyM
XRY8TFL0vIb4lNso+qr2aXXyozDkViACy2hSG+R0415lQAcKnAREZGw/XnZd/JcIzbhwupxw0JjI
TR0y1yVUqskXPO3WGkQHx2gUBvSW72HMcHTV7P816MATGRs6kccgDhr/jmldUHAD/hNGoP/xcl22
AP5gHwZHgwr0YBIAgjgpmmxTbR0IZCPMBURBS7RnfEhvlsn2jJFjnJh62+pO+sdBAtHEl/f+HwmP
9i1xuNfrPPvnzecHw8uZW/gfZRg1uWMUxqPxQKCIg8pzoYEew4nzjfnVeWntvM5vX2sG+mUKbkS4
SYB+zvN8lhAkNpNqrZxQduI5KAocpx0eZC/7aSZjeRIEwxTpIfhrkXPPIktqjRy+GUxrwUodHFhd
bBR0f0hDZFI+QBxn9HisiKJnRjKg5gQNUVwP/5nkjV1pBLLrHpXwuz13eij67EgVFsFPIv85fwpo
hneN6Fe1ssQylUkDK8EMf0hmveDJm7X/5mVVvkPwGpE1cCgWiXcpQP0J1/soap2Hx45QxvoFkgNL
31gh0jqlPzuA7aDoVYzPyhYPbckPJMB6DMy4rMrOKBzNOOKGtUsSmhEVd/N3QDA5HJbU6j7/c8VW
GTmXZowvyoCX2fimIa76SdG2rUdaxvwW8K5vtZWkjYUzHFtPy+ZUbsomX2bTSIAn8ypa13z1/1wx
Gz36BvG2MuVXdMz6LQ/GpPtr0t6HG+Os0J2Xwqu3xYzF1ENZS4mEcMHIDK9+JV4kZcJTUuPW7bL2
CXTKPUSJtrvlCz5dp689/SLyGbl06ACcdOnEhmL5sWegzdygUoD9XYSTqQsxM5iDx8ak++0bCqat
uAEO+AlJUUdt7VOL9SVMS7CBBO9BbFCt+H8aeTcM2PYch3sbdmJA8BtXTCvQRQ71FEV3LpW+lJj4
UwZe68V+pFfUv2y+n8JrU8jQdFk5yWAHwbc7kLcUCcXTcxSTl65JZPr8nUX17V8jkwZy6PrrCe9k
vR+u50a3fVJ7if/8v8ILUc9fEMaxjxDPrZugNrnF4o5Q2ECGeZXwP3phBHUS2hqu0LWYb/tfMIfW
WrzSIHGcBYUYkT6AP46f8R8y5JmH5D4CrsczgZdbwonrm0ogThT6JpJW0/b6U+DlOVjvAxh/kGmr
pqtdzR0WoDs+yrpML+gERZ3qeuu4KbJa7jEjCbmL8nVGFYCkqPMqVhP9LZXbe9ox5P5vEvJcO7bo
8WTt6sEU5nXpUNcXdcsFOUngAGZfiL4UfmbUu69SNoQpYEA8IhQzTkkoKKdL+ctCDAiQiSRTsEZM
6Os5EYCfGpKSaBugeb72utX3LL9eVephYxZDFNggscabSSqNKPkjZK9YhfkbvYqXPU8KjkFJ/9Yx
5bfp0Ryuw0eijgw3wT36TIcKGoEr0A87Iym0P5YowY1dpykuZT9onDQzHq9BcmbdnRaZoU2LpFn5
cSjxiVGOffvuDhQTQMsQ3op1FekTq1RXdExhnIVXd6vzMMQZRuw0WKyweqNp3hx3YQW8AoTuqs+U
ZF7QJdFOs0+RHbR5o6ZYjEwbqZPApkUlh8fRi+1EaBgKfo41gszyh3uZ7Qb/MJ5a/nZi7MqJ0+cn
p724xo4gc3xVjfp6IwWyRbLQgHErL4EcmtEVSg8CdcYS4o4iT46VBJvMgwKgSIr5GSlIwjBAGn+8
yQJAexkgEmiJ18EdQzp5Mdw9HenKyVPP9OBpejXC3clRHRpJi+gRrEmwQOWfnMrdEgOeYyBGtjE4
QlasLWGFCIhEjg3zQ30uj9IYj7b7sR2DPN6FNy4HN604u+2u+LXjSd8/RwBkTzj3Y7NT9FWKsdKh
uZ5IL21ioAQAQFvkhYbj9cM1l+h40IuWxv9gRwJKlbD0w5DFp07fPl3K/toe6G727/Paa4yBbCpk
JtokeBnorCIAJXWTQxw8p0Z/CtKzO6h5yvaL0AfCj3caomLO/m89z3MhexTrqMVFwZaDjIgeigbl
7TdPows9YiJPHGm7jDfa7ICWLpwOxn6OuVLk4HgVM9dwoK4koIcYcNb9WZeNbDCFuq7Cqw6nmJqN
roKFqOyoxd1Bb/fytDxRD8bgqVotiCM4UXyc2uVEtlsuXn7a1yMcaoN+j1dXOe0AuqHEwwB1ReXI
PxTREMcWkDFsWeMLgtOnTrP8ur4bUg4UR375ORZmMXAFkYVtwroW3Zw8bEm+eiR0jR6qnP9bbXWS
aCx1lqUMBMhhmM18Ji4kLKVjscCEgXRGeX9oWidMgMQK6BJETvyjhQnMiuKQE3f/Bz88kD0Ggjf1
jW21vX7GCIu1FU3jyk+dFirdOeCrFmdinovT1PsBL15PFaJSDFys4BTpg3YNusEWiQ3NlUj8cNft
80wxBv1sFX0LoBJDRa/M6xqMz10hVdYdWm2/xsjPYkkCiyU30yxftwaQR+Sz0O3i4LiEdI8lHBoq
EqkHqNyvkLK7yVv7TEYmE1avKxZ5f2rcKwVM/SVrM2iLWxJiPahz7pd0D1jtXPuN7LI03C0xPeo6
nrXqUZVEF8XvCDvKyOgbcF5HP2K88xK42gRJUDIUaz83rtvauAD49nFA175sS3vWg4cjTyO4USuD
A80G3f1ytaKYmtSQEihbaRY7hm/m6tltFEBrqIXSgM1V69iDpKnkvXkXePUqsogPm9cU0St45tCN
F/EyGkne5Is5GWi0zJqLN6GLcngt7m0AOG4a3qTVvSMeRfzRW1ac82U19vz4ahjeiQyVugpSKBRW
xiQZjrVD73YXQcHHQX1bZ0rgtureUVVwPycfwQy39aZ12XA68WqOJ6N0OrNCc2sfQ+uE6NKaAi/n
F9SIzEn0Jxh6nb1sDCAuYm2ggSr07TcP8N2DujBXHmbfxSCUKN1h0l9IsMTRI2k/aaF6e6rNy+PW
eWvh1zzQRo55Ca5O9bYwJFJtb4zRelH29vYamUFytDG1Mbw3ddsn9ZSkr8w+RXskAo2W6YNKjxJw
/XiwbTHhHmbmHy39hocoXRGBJTobh+GZPGRT0oybyqfR9gv1qb3AzVtq4tM2irHUHqGl2ljdFLxI
gtBtVULBJxwCwjSeqf6jpq8ak/IgyoeRWsXG9t9D58MjhAfC68ppsvUq+RrIjg//d5hy+yNpe5NL
PNE3DX+ES15YZak3wFQ2W29aeLv/O575QJLw/rdy7bsqNawD2EmrgiZhEk04PbE0uYCHroEi8ZPZ
Zsj82G1uh+A19bAFGYR9X88MKoHykiaLrYONH//UkZYZ4GLIIC1BjUbpyyV21Dj3BHRdh7SHPN84
mAD8wnioGnK83ne6ovHxwLBIzKMiD23OqmEyGZ15gtVMWUJwszDC0RPpzvJRAQJJsJL/TEJjAXPH
wSai/KZVyts3xPsBqbk5EPxrHuxg4BFP3rb1lYJJdoVWc1LTFmEG9UpwMcii+5cM0eLD8AA5nZ+J
ujhWl+USFpB0JMx0JJSIiGOngmzkieBpqfmdyvc39Ugzj+3v1B7oIhanf3KoTdqR1wgCrySxqZ/+
Gw101REtlDqw22Nht3QrUY5EQuuBwOiPzlAW/KQjJOvb5rvEPhprLyZaVjtt1gUiHwmxNQmYUKsh
faZqw/aI4uLaJ/SCJAzXiE/Bp29ZT8IU0nbc1lbV/7Cuv7cowYodZF8pHp+cvDtDkEVvxgucJSmW
I5hnLJfq0qIwjAPWnftMsqoR0y50Ftoq/oMAfUERU1beZfcuCajUs9Y6gc0VCUnZVzNSBnxyuL4s
vKR+RekMxLlK0K5keCRykf4x7/jDt3WOMheQPrl+op9WQGLb1IvXduykQgnpLL4WbO8rqe56QcFn
IyG5FquaN/igrMd0TXw9030CHiph/1/J+J3V/NqDxGR41MIS+tjs6xC2yr0tIFzFTIg/7J3RzGnn
2ZxMYG+GDlzZhU/rQE5KlB5jpt2eKhaD4fOi41ZA87Uz6ygcDwGAvHxq9YfgEMJiAJH8tNAAIa6j
X18m5uCUuNg64eeiTeqNqAUZGltAOYS96eYtMXv109MYY3wyPBIKj6sTO4gA0suzjcPmVIcBX8Oq
PpeoS0BOyiMIXYMHFz1xnxa3l56FHfE5i9q2Ox7CVgLyz76t2ElJaQS8ImZL0rNYVOK+NCENYKwk
BR4h/tT7vVt7/Uc4Idwl6z6FpmPheBoku5aCh+UlXu7lQ4aFyf3SXofBoKrGc6BGQBknVc7hh0Oa
zRW12Kxf9gm9B2m9npN3o55fLDT5ex8Y70VkXNYQuKM9ZhRumnpkDZvuxiAvPqNPuBtZroHeGch1
HwjBtMzgDWlEll9P3ERqlBVLeqxzVan7J8lQfKu2U0YwjXh0aSmS1NCvEEA8iAySGIHnNGx3fYig
VBbMtukpjtT3ygBhCTfT4GcHWTfBHHJVVRG90TrLZeSdQcQCc4bxnnrIGcO6cCq6U9HEQQiNGzsT
Qc5yr0bm3X1W6S3f4CcGbLzRYCaw97s7/RxRolrZTOpOpuQ3P6wDvK7VxvfKGgaeuklZsOffjZWZ
W9D9Vls6QN/ABoTePRv1UkCd5pj+PnfKODwkiiNoqdvS6c1xeVTuCQB4UJO2rEKuyhnNSxVPAD6D
I0TltTkHJoJjZB9yTaNYv2fjpEqJIeBEz5tPBpD9Z9WobZyLGjPdYPQuwFBncANjHfpISbrsR23L
V2uYIRPl1BuCM/miXMSI4tUfAPNbcO+y2nCXjI2LNmb381l/tYqSDt3zS4yAMho1iirW7WiftzWj
mGKYn1vtV0m/ByT9i/YjfaR/koVMBAv9mQGAl4y2sriszhfT5vDuT628/Cn1gTgOjOFGDeUmHJSw
bA+XlGlL7cnophK6rn5XBc59eY2PjkMoxiIdm3TJW7y2jUYpWdwEMOfeJ+tXoBC8GloVdIxVad8o
M4TI1Fbh7SCuGw1QuUZeSf9SrOFObEuM0cOlu4vgTBL1+ZIJtMGGbvLS/vKvB7yQPKDVzU8FxoLs
2lxglSlfcCh3L9AeQUmIzz/DfoNy9zwY8+7XDwoyVPJfe7CWdsFDepStp1uLi3QTfVd+HfTGlWAD
ZL0KMxyPM3B/nSEQagk8Ha4nXPkkIGmmcwAf76d7SihT6ktghTtrKBuOFZvyJn7Tv/lJmWEuYuLX
iUOcFJqKiWCul6Cbr69LtS6b2UcVp+BvKiy8/D7/fxP/4uj16uq0AvybnL2iglMpT1wTrm17U8mR
8tV2o1gBYDs7pJIY1vPO1+wmCpU6PvAnnPuKoBWt61wLGhVBTXdIBj1ibuTHB1ZTz35ON8I0x2Vj
uVqp6QDd8CqdDe29j9QZ/ovyvG5kxdEcMGeZPMKZRtJDcd9wCE1lOCzNkyZD4FLKz7H22V3x19kX
W+2yhfImzAeBHyiPxaBKdErqVxoHROZZ18xcM9aOvRSEDChpZC0/kCKfhjpHfqr1NXd8TBZtubjz
0hLfcLIjKfLwUEj0e3amAyPnVclHGLPIB9HG1YhW2MpG7T/HTJNvTbxs+2YVlN0jHTsvthmcnAl5
UmGhpVwEzxI5A7gewE/QlCwbkt+lJoEDBfch+LJwx1pXhR4igFsY4SHsC/4vcmVNyQrjAM0lTKml
LiFEUwX0WZdLYGNEEAiVCO625SGMx87UlHBeCQuLtlCo1bVIGwiuP7mtdN2D/P1N7RKT+jguOVJV
gL3zb/CujnUn+j0HPefJszSG2ZoJXrTH7dSYWE5icKDlyLMONxI4PNoFpdxqR534ogGQGENefi+j
hjk+mRpxItl7c1Gdf8ZRIi3h8FbiC7lkC0vYuSDkBaBJ5Iu5z5M/N0AdyrKFrzJNHRu2h5ZgKtu8
/ActarPgaLWFsLupKFE5TM3bWjKyFGifj2neS0z2JP6/I5196qbn3wkfF4bKWR9A3eWwOc++RTg2
DEwMoWmhbrgx2shNszPvyUfjgWNlZmbjSYx/35kkt1llAUEVF/xhKx0NjEvmiPr9ddJT9N5UllAY
U6BCBBs2dF69e8g6zQ2H3615UGQwHsrwWI4pldqzXi++b0gzUiUoAmiG/rgwEjwWi0tBtjO3ORrR
oVjckHnMdUqusIaxAmTY2xDsuFwgWZ6T/gPQc9dbgA6r5ouR1kv3Z3geZU/bmlfgGoiu4nxrWXwF
xmyyIB1ILy4izeODPd3hQrCOtfy3DnplNZFsQLzj2jfIFzTYELFRfmjIEIxCDWj3FpGDmQ+Ipjax
hmbVeAsDrcngoIcqT4vzruc4pYGXyepnOqv7zzFTdemOej7NuTbrynpzdkTKeCw4XoFdFNNW2Svp
6ygz3LWAmP75DQMnzpl2wQizfHHFnEmJO63/S9e2nY0UxgKs1u6kVy5fUcTjFMYHQhu0//xHZoC4
Tb77wCs/YZJvxEB0ZKJxiTnnLzS1JTq78seRBt4iIl1JC/rbVE6t2yoW5zw0p4jFnoXusg4MFgNo
6dXNdTS4w8KqG3FoZY2s0yQHZgVmhd4cOU/84ALXtMx0F7sOUBrs/u0LaP9B6cV1qR3c3m5B9+DD
XrPYVLMQzKuuKZ9irV1op9j8HMfFZ+BLYTT/rmHgTARpsEeqGH6Z3/LKzWWDKkume8iJViG2CqnF
NRHMolxcK+jTXoilhtoK2qLLlsG7EngcpkrOHotb4xzHiYp+6cUB2Jo23Ff/m+/V67E3qIcMKxCc
plqxgM7r3yXymdEsunUCjVs7ZtQd+H4f9TG+0AYyUrlMhgSY/X0SezkwBC5pVtPVXCFx2gxvP+WI
GLTBfdoWNwWCGzJjf4syNDpGDmA2JU0qE0TXMACs0BJ7a+h/n/OA36Dk7jvte0XkBsQNMeth6eBs
UQk2Sg9AmOBVe67Chx/ial2fybGQadQGVNj508hsYH9XCgn9eUnBo8HMWQ2EMpN7EVvaOTQBGLp5
BkD64KafFW05GI5E27Zv0c4Yo7h04+vshjeKZpDiPpOGeAjpKSQj04Zf6P4V2a45RKgpgNZqLDur
O2SHk5X9Tr1+frCtOvR2gWhHRLGJeuTD0hYvK6cuYmrBpE6NirtM1kq6ZFmAqe3XGrbPxcxFMcgk
MXEgMs2onZjGF8SdHypF8NgKpbqCLQFxVwrHlHLmvAacxBYV/zVzxESDgUYVWE4remV7P2s=
`protect end_protected
