��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=A�w�����ޡ����$n���՜%����~@�қ�IO���ɪ�H#X Vyʢ}�<��P�G'?��,���ɎĖ�H���6cT�.=� ��x$Q�L���S�!,���B����ڜ>�7Y�'T5�Og�I�P��=�S�'� j�G�g�m��[�F.��^�kF��$�9���[�ݓY���8�!�?�6�~��;�4�F
�hxt�K�0�����+h~�rV�o��M��jå;)��]"X52��Uk��O;�����aNt�VŠ'q��Cd�����*D���U0X��KU�7��G��I��÷iT��l1,����s8g��ȓΖ�4l-��S�W3��f��׸�.�sI]�t)�`�+���ؾ�di�	����"�dZD�&�˹�5�H��U�8�S�X��AE�8����E�����y�D�Ed��V�΢|/�#���!�O����h�)%�)��T0a�^V`J��&ى�Z�R���z �C�tp(���������3������X=�=�ex������ůO�k|H�ͼt4&�3�ߪܟ�Jw@�K÷2j;ɀ]j���$�`�s5�B�(-G~5��-~��8��0��������q�j��Wg)�Oގ
�QTF������a�)�o�6
b��&�)�҆��{`j�-V�#�i ��W��7����G~l��^��UVLgx�H��3֢󫟩q�&�t�tb����a�z����?�K���eڵU�h���B��u[��8D$�WH7ײ��0f�u{�y)�!�����(��;Ĭ$4α#�<�)0�㠡��1�^ÿ�s)c���Q����u�ЂN+�����'%xW�1z�ļ�x
�����D����@4Jy�]c�d~��^��)��G��^I��?�6q���S@����yag���� �*���ʨ��CD{!p���[_�\r��D�\Cy��_�<���%d�}W�~��e7���
��e��J��z:(��rT�F�)�<\�䛡z�6�!���z������t�_���=�<ĖʠV'�	�e�S�?-ˈ�x�N�!Uaɴ<�����׫���a�1��fA�CP"��*yҐ.���4��a�t�Pˁ��TA6�x
�F{����>v�F��=l�[�6�)9�ް?x�;]�"���%
ڵ$�𵹵�X<sZ0�`ˬ�z�s��q�HH�S�"�A���X��jN
�T �:�����Q��L`�n�u��9���L`3�o^�+
^� ���;̡` r��<�)�peN��\f�R�P���7E�-~��;E��̮��Z%��,�ov����^�S�&�d�%���W~��t__B��s�~�q}F;�1�>���̧B�uڈ�G�.���Ch,�<����1	"����K����\R�!��zziy�H he�U�������2��7�7h��p��Ӆ1�EtUI��V
��t�7��8\d�HY)�?�N�[i c�x��neDe"g�i�U`�C[���Hј%�:,�"������sf�S��Ɏ��&�8Z7'�����fЏ[��,)E~���V���?\@��)�7{���16���%�D^�]�R 's۬G�8�І���n=�@�2�d�jKl�{Df֘-���ُ���}QN���-��V�v����
�P4p$�9��#�<�����Y�R�����險;��kgvQPE����a{��L��`}�r-�������t��P��ۦ�ue����HU�H�1R���H��������>�
��c+�"Ob���P�&�N=5S�Xt���W	F�sSa�t�
AT4W��D�,=s1�1��9��^2���YU\E8���̄��)�&f�k�06dU'�^���@�����@�Zl �[|ɨa��#φ|y�X�FE��?K��tЈA7U��Ec��
A�ڼ�ܺ�e��1����p?.؀������21�)ǟN(R�'2C��إ���:W���v�`������8E�Jk=�5V�/�ɛ�������r�E�(��� ��Q�p@�.]�������e/��y�u��'I:��O���iX�)���/)47H�<V���5���W��,���9]0�{eo4%�]�Iش�Y}F4�pk�..�jF!B!L�ʐג�=u�U�#g<����Pؖ=K�)(���l�>lW����(��?`y������_�^�-?pW#ݧm��&�DU���U��Xr@AGǑQWZ�n�5�&�IlՓ1��[��g�R[��ſu MW�1�ۨ��ouI)Srcy�����@�򾺳7��}4�g�3��9'��(m���(K~�)U6ԤS14ɦ����t=Q<�#Ĭn6�L�.�������������$��|]�L�x�a��;sPPm�J�{E��a�'�ͣ0�S��Dex���.c���Vgw�s��Y�!���i�\�U��O0ͨsd��r���FY�+]��s��<���>f�C�2!J�= ��A<��p`�.g��Q�S�Y��KE{��6��w|�z�L�X�wtU�&�eB�E�c#T��m���*����r�TG�Z3dfem1}b����y+y�Q���H�0*�(��1�J'@"2o�}<��q�ڔ��W�6�U�ݲ�į�6 z�GAN83��i��T���|1�����LC�(��\����Yp6�@�+�@��n��/������g��(}��gVR�v��
��$�Z��o�U E�6��5�uYrVs�h>c��)��Y*�e�u�@�9�ݮMi3�VX�D`j�m��N�:*3vΐ�$��H[�WiZ;���,�2�M�Aθ��]��6G��X���L��~M��<ً���֙^z�rګ�7%J����c�F�����<����Qa�����cֹ�Z䪳A�)������JW����irt�ڳڢO�y�ݖ;���!�h)����IF:��?yO��W�H�T�[�r5�K+Ns!s1*��X�pΨp��w��v���)��gF1��k��r� �����g��B�lGh��'j󕥐�0<��A�|����X�6K�J*��_�6�@TH[�}�d���8�W���	�uh��M6�M��?��ݦ��)�z��.S� ���B�t�f��^�e���F�N�?OTu���z}�乾�TBt��4�2P��_u-�a!�<��S�"<���Ѥɝ%-�4g�T�~9��JJ\�)OWiY��S�]!g��ZF�{"8;&���<�nⵤ�+v�8��ݎ��a;��@����#T���E��-
�ӛ�u���S<��,Z�f��
`��=;PF\V�����P+A��S�g��5^�*O�9x�4�3���-�����(0��I�"����f.�)���
lq���re�Ґ�7�6`i�ц5�4��`�~�b�u�lpڼ�_1��򕞡�?�t�>���%5>0��:�S/v�	޲	c\�Y	���-7�H���e��K5�7g��U1֤4������K���+�w)�爵��l'\IKh	�А#�&�`R�mZ��=[���RK&�"�6�O�P�r�H�e��߻�6����j�ABI߭�^�mc�>�w�B�	�(�q���y�.K��%�@H���!niZ.?�.(2�Am��T]]<K7�^�B�5�TYF�,h6o��tv�v���OUKI�b��w�����_�Ÿ�f@�C�����T�g�X�R�K6��+�;�Or��h7О��]3(�]�lH��y�H�K;>�PW`�6[�K�ք���Ys`������$3�-����2�@V����5A���v�B�S�c=;M����≦�T��&o�wzQx4$y������i�Z�։�M���ߝn�\�z���.���$e�
�t��G��&[������jA��jR��}(�l��s8=;�{|]#����cg�j�EYݴ�)��3[�.w�z�]�r��O��z�O��4��
��ݥJ��S���F����ֶ.?�?��)zD&�vH�aҩ}11���|���.K].F#��To ���W���s	�� ��̭�BD�FO��-�bI�L\�/���j1��¬KS����`A}�n�lDB0o���q
-�u���=u�zM����c W����gٍ�c�����?q�ÏNea�us�� <���av�kDEO��;ڰ�]Y-0bȧnӅ�y�ߛq�>j�@��W�$�"_�Я[y�dPvxHA�+��K�2�%*������ƣ�ꊙ)��S�����X�`�\ڳ�5�͡�{DԴCl� @B��H^xiS�L��X�:р�q�~K�[W�'_̆.2�ʩ޻�fW��'�?��Z��^�v���|�	��p��a���Q^-ii�\�]z��ò�9�*�
�_�/AHQ��|�J���y$oM6�
���Q���h	���>躹��z8T--QuÃ��9��vn ���o���� �``�Zg�T��w	�dM�Xt5����`�.�J0Q��8��|�2��*��NU�Q�S�dᬅKL�%`�F�>`���nn�W��E�cH�D���{���������I��gḌ�����+��=��F���X����5f���p�"M�>g/��=�����@l{ai~,1<iPO5�a4K?�Z'��xou�[}2o(��huU�'7�D��%pi+�����dp��k����X���ݧ����{���V�w"��=/�n#����[BHy�{��vh�2�M�qm��J63�����4j�{�끖�����vq�yAp�2qmG�&�B(>	쎜�U����r��j���fM����V�.���H�[�,WȡZϰ��s���~ϋ��H��p�݇�J	�k��T$U���ڮJ�'/�̖�h�ԹސU'j�뿉�yIWI��'=	�S�(&�;�(��}!���
���,;��5W�'1�/�o�����-�ғ��5<
O$�y�������|�L�3��Ü�����X�	��nL���q>Q�7}Z��W�$�C���Y�|��eB��]�0�D�_d^��Tv�}��[S1?=T�k)�CzǑe��d�9ԍ��P��鋼x��v��"�!��fR�)���D��cL̸>�c:|ŵQ�: �|�(U�1}��0��V�b�7q碒���S<6�l�z��/��8�J�^�}ڕ���2`+��4�����K�q���J���6?��nq�h^�j0tx74��zޥջ�����9F8I��I��
��8\�W��$�ym���i���h��̼�b�&(���D�}�����W���o�I��#B7+R�G��+�Xa����
V.�I߶�Ќ��F��W]�M՛�������A��?TP���7�\)�u��+䬔��9#�J	&[����i@%m͝m����>��00P�2
ݭ�JH�;�p����	�18�2`�U=��&��רڜR��.�#�M4��'���8������%�kD=ҟ�)�"�	t�D���A��.�F�~�k�������J�P]c�zcl,� ��]�I��T��zʁz�I�ĳ����$1��~~a��5MH���ǳ�Nl��o���N\:��7�-���~��?��+�-���p�\����ˊY��)��x+��<{U�T�%�|�5x�y]����3�i,����m��#Z!"�h"�]�dvb���s��	�o=,�n�:E����c���,�X@��bKt���X������_3�= �R	P��|2�*���xqP�(CJ+ou$�t�
���=ͼ#.Zj�-xy{;���eS���ձ��;´=
��=���%�N��]{m��6�cc3�hj qH�GN���9��ǿ�Ϊ�k�>��-B&[�L]c׫P���x?�qy"��pfA ��̚V�Q�25D����%���W�I R��� ���P@@}�X�S����Wr���hrF<�Ԡ�=ͶOO]MJF���ɵ&\����݄A͕�Ƀ���(3p=��A���	�����D?+z�ql�4?��lF#�b��R�G 7FH�����%��Z����Ę�����ם%����ț�m��*-�V�wwSE��\e.JyDH�J���㠟�w���0#��e&���(f���7@�Ҡ���~�f3õ}��lD���tQgzs���8h"�?H(q���S*"]]#Σ
�E������r�z���Pb��U�B��ϳ�!���Yė�<ld$,�o����9�0w�u5ğ��>�I"��D���:�y4�3~:B����n]&�~�F�^kЊ{��|د���A�w<�(���_۹J度���(�Γh6�g���&Sc��e������ � ɠr [8o@�� B�b���r��^�1��G��3�(��ø;&Xi�&Z�D� ���� Yh��lykKwy����6��N"�(찅;y�u�;~��b(�!�7�@��=�"ĳ1Y�-)i�|[j� 3]��V�M��&0��EvA�rq���_��	���sc�D�t��*˴�`���U8��v��qg�pK���5AM�\L*vW�Q��P�z��ɊBv )����[!��L6� _��F���$Oֽ�o�|s��Hr8a��쨐ػ_L����x��Z���5gK��H�����!�J���I&~��|}�5��x}�4a�Y3�,#���v�:�N"��,_��(t�i