-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yL4O1nPK4X62urVT5EuXBZVABm/V5plo359FSQBuUKaK3XjOZb2YVc7ThJcDDzolyff9IPdRXs7T
0QlTKpbKbnPWauDfF+OGlidgXJZLfkf9l7c8qh1tNDUkrOJOS8zeXGXvAk66WMzkPkMCBD2W1aq+
buHhYfKWCq7vnhOsrL8B1Af7ltnSWo/Ni0gx7oodnzvTbkNNAG2UOhSlHBV9J92RhYgAHFh7GSoP
pWXGOrOlsM+90DY0ARox0+qCrXdX9l5mi6W8ihQQukwYLbfAtilQ6ZW8YlOKsbGCW9PX0ONQBb5x
J2f/Rzudei0CRzSw14HUgt3L8TWbsPYVXUPbng==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
B3iWuO6+aMX3xhph8M4tq5uc+Nnszp2Py7byFzMsrRd8owyBgzweI7UtflIXcXOn8ADpjmdJkE0c
UsKaMK33Ils1rUvVfugs3mfC3JOKp93q3b7lrCL098qLX+H5bfJziwq7XFEHgDRaXAKEj42n9RCP
lolUHWXcP7kuVeFhF94VQWYIWq7dQmhqQ80L4SJ/UJEWY8sVcNa63OmXyk+9CJZmCJR/Z+ltQOoX
7Tjb2WooxFv95sTJcJj7ljxkrQV2w0FTjUcXZK5IoYsOExp1LlDgXJAiJfVXpQHTKXpzdScvZt7s
vI/49B9kNlMEetX1OLqV8qGydwVbJSfaalUglWqFYse/NYL/BVWju+OzB50mVqZ50c0V64CQv2o/
/5CGxexc6wBLzEkRvUmBvsURRAXZKBDh4y3sci+f+YHt92gzuxt8lxo2mDkVYrW7wv/GvvDbY2sP
UT5Y3g6+5g+CjEDjzlqQwX73BgLKkrNKijyOzZjIbbx/S+F6F2hWu4MOowJyUPT9i7t4kGGDa/Gt
F8pscTdwEyL2dEycxgoj4v58EvsSnoUm6YEXOnLQdJ6vBygYRP8f6g9UzqNek4otRqle8SIZ7rIy
oNXf2CzPQuR2JuHEy4nen2XD4Nx2eJCkCsS6soJe2AK6Kk6HwWjbokbz8l6wIPruVjtZ71EkYqom
uutKjxITE8mnjRbrSw/rxVxpvOyRx8qP3/BjOpNJMqlhve9lyDRecZDlgOL6WiYrAP0Tz5YVUpGb
4AU0+qtJB+DR1dVAOVmcm9WbV//llrZEUjYlo7INz5Esu+s+++2hXebFQ4wx3A0DzjacR5aOBL/8
TRvS7oLIdUiLjRs36OJ6dk/5/KYECyp1frOj78NF9rQfamWJc5hh74yQP1Fv9pSylQEgq0Ohra6G
v97CDV6XDVkRn7gLdsbnMZlz+DJrW9fkKcn8SoqZz3IFXTI2NnO+liiqZ8pCs7lpFtoabRbjNTfI
LngBkLCNOak04GEtzhH3tgJMldjKNykoAIOssQoKA6O6tIZz2bFGqIwaIldMLqhyG31vHahhvvtJ
uegExoSw4vbGwa7TZehN9jkjCefEY2jCWG/T5iWl/iuGej0LTYShTRetjmPtqqAMgORfQd0YbCVT
ijus90odHv7T0UoqzWl226YRkcrfYkzAzXshs8KEDL0PUiWaj8XnVXgvkcDz4RWwEL5oO2oz6+fI
+adNYD0EWLFE8uG5rTf7/wp4bzvBuJiTTOe2Nir6fi+8X/aNqsMNvFWGWIiLI8zwjHahMBmGU5MB
bYdaBaiR8dutFf0CHZ+QPZMmeF1CmQwVlQfqgd7yEnzUMSfdWr0Rx+rvyUHmgIFabowtwftEmD9Q
UUCuStnfqK4gUEKFBVVBrCXCx7a4rWXf8q1BVHlLLINVgq6Vgqkcz7T1TaX/d7EOre1w2l3H09UA
hdYLm7ry3eefQcQt90hgUnCPZdBYHqVf44qdBACNzdaXZ9AuRy7BcLpFAS+eyOhyhhA2DrVtmOqk
5IklNOI/VJBhGrF4iXRfnA5vAvdhvGHX33UoYNkzQsGzk1QJDE0u0ZYuhZkElvvN1axoskFs8eHx
3wzb4OawizaTjA6H6zzYW48IP0mhm8uAFUGFz5hd2XwvwwtQn3eP1My10Gm42DRYlf94Rl+HBjAe
wdnCfmsSU7TTpRbNss9vCc43Gho4ZAGF5nOccZaXYPE3FBuKnPc+sWI0cwDmFYR0I1n4aN9erwjh
UpdG7dpEUyBYUg35EILrpk3OiAvLkxVz7fzz0oVqG+Pjs/VOWiMBKKyyX4ZkSpCi+2d2RLw2xf+c
AIBqvtFYQGOmNTdYxNT0VroL4kHlcyF4rFYZTLFIE+yWT5RideZUYhDz4kEjJEgSMzaBVursM8l8
xRgvLtU7DQ8HviB7hHuuSNL0ftMF7J1atoer/hwVZgqB2MT+yp4k3/SPxrk9Kxwaf13BVZtmXzU3
Ji4PdJfzou/TvH5OoOpVMO+cF9Tjr+TeGZdw8eaWoF23Gy3aaneobT6Rbnc0Kw02MO4HFXy/H7uA
z6kQFveLjwrMoc+XANptkkw68cyERnp1+ABWj9KBAA7ZDWewj2WqixnBUp5p1o3kGEv5SFTx6XvX
tUiTMY6bf7SwMANhEAcVQxulW5K71H3Eak82MWnMerfv8hYmJo876nJl55z7qQvhjQ69tG+P6pi7
K1PFkvAyhPHWIFOhuiGuM2dLGqLR6fUAZKUteljGmgq3QCVexVhgNhuSsZN41EtyBaJkyzdudBlc
9No88WzFMQphQYGnItMpAG2a
`protect end_protected
