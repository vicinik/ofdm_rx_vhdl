��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l��}~�	Z�[S���5�H���uaay-�L��q����~�@Z>(�6`�Q���̒��Ȭ�SWC
�4����2�葹��M_A���ؾ���J�Ϙ�����;�f) �R����A d�9�X�4��QR�Ј��]Z�f"�Z�A����R~R=���\ �]��Z�J�C�+�i_�֧��/q�b��Dv����K�\P�م�N��z��1���"�sO0�<���z�Rlپ�}��`��H��*�Ҽs8�̡D[3$'l�&���&D@�X/"pz!O1�����)p����^����5J�����)�6�#X�t��}���vAዴƽ��Y�h�쌊�a3�x��
���w!*��Ǆ�C��:�S�/f*"*����8�S��{��eKy�����.�<8���>���uK��1��6�m�;tq��S%� G����Cֺ�q?[����)0�S�2e�Se�+���hm�W��� �QH�SR�(���V�_������'��ٔv��ꎐ�p^���A$�ɒ���5z��{�/��2�#�)�=��i'�K>�Et0\/��yys΄~1x;N���H��G��q%����f]�|�+�ԁG��u�(���(̑��8��F�؇�p�uFi�1�=�N���_������5~B&&P�
B}�$J�osKpyÄmG���FUqs��.KP��wQ�I�,���PF��T/MYOu�#�qTzX:��w*�9<4�ǿ�Dȫ+Z0�?2&�E˽�KR�'��F 2$�oWU.a�|_ŉ`�0��g	8���\�7�G��f�>K���m x�h��=P�m���H�G���^���k9FB+��`��&�`��@Q�(��ϯ}��,�����2yC��CO�.��C-%�����D��A\�gR���U��*�5�ջ7̳��_���򉐒�z��b�a �)[L���-HUC�PU����.��O��bPH�Wd���Ѧ��_(��o�X+A��-*~�VlwѴ��S� �N{
^5�?�f�y�ˤ�����3o6�^�����<aP�'����Y��9o�!����.uF͊i�#�h�%&}R�퐮�+H��ܳ�(mɁ�c����(�(&<����Sz��W�:���ʨv����a�
܆��cC.��p,&0{.�v2O�!�����,y]e�=��E�V�c��ܒg�f�!�_��\��v��v8���ď��6��`�tK��㥵r��ac)C���޿���\���"��C֧���7r����,-��*��%�׺U��z/t
r\�~u��l�_e���3PS>��I�GBI�9��J���<
<0�
��"�sX�oΊ��؈w7w;��VY�$����9;�_�0d�#@�Қ��t�"k-�c���>�aрP
�O��9~�/��]ۄ8G����*�(E+'Q-1r�Dl�@�L�M�*�e~�@���������L���J��~t,�R�G�|�ʝ}�!�{[�.Ì�i3'�a�vT�;!��=���(�5���;<3��;����nB{�.V$8��ه��`��&�v5��Y���I^b�Z@���_�>��g�=�,L��i�Mqy�{��� F&�Q�@�*��ܑ�Hv�ןT���sY���m��gd��9܎��.WI���.7�㶜��K�L§����h�ڧ����i��}ZP�҅�����	z�ԒG'��d~ϛ�~| �.�<C�J���w<�g��ʜ���l����Z��Di HtSB̗�V���nrE|������A) 0z@P�v��j�)�h����p@F���1q	Jg�89�Zv�NW=��XX�MyWn�:{�l$�f���*(�_8�T-��b��6X��^���p�ȗET
cZb`ן�z͗B������reϫ �9��l�K�=�˱�&���^R� Z�i�27�f���~V���#|�ݠ��6��x���	�̽h7'����b$��"��Zz�}�~����y��\W��xp���ΰf��r�Ho��݀g��+_��%�1m��$��u�"��^�/��.�9�=�	YВ���&�}?c�RW)�?�t���'�S����\���i<���M��)�'P�w���X7cuby��Ϩ�ܺ#K��A;¹.����$u��\�I��@۵�{�#f��b���u]���*�:�C��O����=��'цx_�̆���z��z��#A��Ē7f)N��B�� P�i.r���l2�KkQ������Q���4����In��{X@��P%|��~:�<�1���n5��`'R���M!��<�J��U�����M�^�%ᏠH������c�9<��-�>3�Qw0 �yg�Ķ���n��9bY;�����[�����Ssþ��b=���g۫��&f�Ar��ר*8�m�ݴ_<⛾u��<fU����������]�!��=�l�6��v0���E��'�C�D�}�r;W�~��B^���p�,�9���'*�Q�q�|͡0]c'~&�����	���%�H�+;�T<��v?Q,�Rs�f�6��=8^&{�3ޝ���ы�V]�N@��>�Rd�d�\��p9��ܡ�|�UL&�Y6G	�E�U�-[o��|2��k��Gɻe�r����u+��/7���&7�Ab��i�$��y{Ejn�X�����^k��mu� #��s��:���&o���j]2ąy����1i��,{?�A1��}��y�~�a���G؝E����ۧ	�8_�F��$j�D�0v�W�B�M�ܑ ���V����7��䄥ʝ�.W��#�_��k�7ۄ8ԓ9N[Qi���6�պ�q.q} }XΤtO:���L�-(�91c"�~�FдMWs��U�\��w���0�ӑ�?�i+���{�zq#��|n ���Q��Fw�j`�/X�������u���@��'y<�΍܄�0 ��NR�����h�-ﺉ�P(6hF8�?�p	���8�	�� J��x-V��!-���-:L���J�4�ShKK�,�/�H�����]���UzcE:�ī�=��we�z@0��b�"ۻ�7dx������~�~�?�<����;e��X�%/L�"#j�LT�a�1z]�6C�d�E\1m8$�&�����^�T	�H=b�}�R ��?����(I��mK����?�B��R��`�����%��mX/�0$-��dw+��$�?�<�Ƽ�2Z����L��94Q�]Q�3[7�m�$x��^6�c��{6�&�ꞟ���R����;�;4�uv�T N�g�1Ncp���>�c����i��$Zh�`1مv�dMR�?<� s,;&�a��?�n�B��.9;���^_�x�_�(�f\�X�����mo��Qw&����>rI���A-o��"������ǈ����	\�I�ڲ�q���[�+Z;1�jB�����\����#b��{��h��-%�-W��l�8U��P @�����ZN��@4�p9=��ǈ�:����X��Cf�n�6v{��$?�l��L�!S4�qK��5��Qj�2��,\_�Z!d��������w�6s�kr@%%O{�[�c	Э,�Dyy(����3We��Ĳ;]0���sq�7��/��:<>�&������~�a| \b���:��]RI�J��,�PZ/��?|��A�Qt�ã��)tA��ㅒ��5�X�0Yj����SLC�+��	��yK��X2c�>ǬQpv��3��ʻӻ��գa6����a�^�Ӕ�J��%���21-�]��p�D��Ҩ��<Z��[$�W���M���2u`�(��?e����T1�G;jL��mfܦI���	?���L{Qpb�sb$�v?lv�����.[�Y��O��zb%����8�rv)E�����^@����0gZ�L*¥�y�qX�)��wc��F�.�!�8�(E@��J��K��h7�������<�O*U�f[Sb<:HX�!���P���l�8Ni�F�W���{.�?|>T&�cU��!����1�ס
�0�|����t�8Ů�0��<���*u0�S��_����1���=Uq��t�.z�E�ca\�=�W�4�x���A�x�|ff��Z������h2��W�Z���U�e�� ߬-�~�.lל(�|=�so�Ȣ��~8�.0��H�\��-Lo�+�?�����A�󆧿���e�9گ���������뱷�jx�p"E��^�X�=L�"�9���˂Y|%p��:�xn�'�J�w=E{�*����×W��Ã�2[ 	N��.���H���K��*{	_����VW�tJ�/�a�6��k�$�h�?D�I�c	��YLP�{E���^�<g�����6���\n��'���r��-�am��g��`jS���`ɿ�u�
�����Q-�:Z�����K�{צ��u�o.�y�/��[= 9��p���<a��
9�Zcg+̺���o�'Z�Ij���/"�)���%	:��<> �����ţ}h�]Đ���V�Y�Cd�F4_?{��7 1 h�9! ]�oN��hX;�j�3���	O�ц����s٣��C�][����Ʒf�w�F g=�{+�zi����%�G�D,~|�e�- D�(uLh�>�V�%��ǀׯ�~>�I��}��5P�Z1��8f%F�zq��[��PxgK:Lԍ��<�:��H!_����I��N&kl��n��T�����>2�,�l���Z��j핫7V,���~l*?Kɫ��\�2ɚLiAA�V]�4�R�Q�¨��v8n�9�a^6;�1-R��?����Kٺ�md(�2�.�Ij=��,�x,��)��� y�m4�乌�>��jz2���Р��e4Һߏ���|y�����܈�O�Uj�?��[��.��
�kL
�yL��T{��8בZst�B�������Ӵ.��K��vT�!u���	���)�LSo�
a1�ҩ�.�ŕ�ͼ�^��W&OUq�er���d���%��R��ۖ>�G��_9�X�-�Ш��}�D|�Ьޫ�B��y�>숡:���4%=*እ.I�|['�&~�h ?��3���-ݲ����.�ͭ��A��сud�1���u'"	���Np�5~��]|aYd�a��O��TA���a�R��Ωg�=��i��~�����'�RD�3�������}���}YC)f;U�9��, �N.T�f�΋�S��������:�~���-����������	��^P�R�&)��:L�7��/OZEc7�[a���
!�~g
�n��X0��x~'��^��4$/�7�٧9ԃE�5 ��?c|�&��ѢQ��A��W�t&���k�L����㞷$i3Q;Q4�ݔ�`�ӟV����?�!r�|���je֨���O��\e�����HB�Y-Kɏv	�R�V$�=�Fi�i�-�A�(|����\.��Q�@�7�-���	@ɾ��&����+=�Xk�:�йC�Ǯ'h=t�'[6?�w1��SX����vg�FMT����M?�R��$�.��栃!j�0�w����UӅM�F�ӌW������ ���c�h�����qbCxKfK�6�!a��a^#�i;y#'������u엌�G��~�$���K��YX��R9�P�*��,�c�m2UFf�/�U'f�a=i�f���,��:O6�.u�E����i���uF��;��0�`�(GA�t��*�`�3��R�بL��-�_˪�����FzE1�$]�P��0����T5癵�\���y��J7%�bp%=�`�ذ��"{�iI$����:Y��
J�e�rVʲ�����x��x��_}��<�W�C�
��I��	!��}<('�$,�J��ղ�"IP�;_�	�(0�(z�4�
��C��r?0��	ء�~���'(tJR��|P��V/�L'7�z�Ϭ�py��H��y��YTz	�������^�钂'�]�)qx����h��	�� �b���	o��+�%P�t��bR����!���y�q���[{9��|�H1��s���P�����)�4�̼��̙���2���^ x`��.ؼ���Ǽ:z.�����V,��U�������ɇ�
�98�}�M��34�]	�� W��w*'�23Aq<2���RM�� �����82�A������7 ziH�Q���Oc�)e�d���N�@���=y�u5���Z���XB�t�R0���s��B��_R#)n���t�/�jx��#ـ���_R3�T�ށ����K�x����ςXb�v�=(y}�ևao܍U�9�mh�G=�:@BV�(�9�/�o�Χ"?�0��.�֌� 7θ�$�Ԛ�1��7gv]���x���1�;��k��h��^����ٞF�~1i	?������F�9O�2[3��صH���D�����~��TCY1�����^;ڀ�N��a��Bn"cU1q/���=�eF�+j�*�ıW�1��5vx�S&��S�gVh;�����Ϡ�`A����m��jv�L�U�6g�Igf�^u��&�]]/��_�h�ˇ�D�"7m���b��;3ވ�����:W�������E s��F{�5ڭ� YӁ�L��ἵ��4"i��=M窗�Z���>������v���^f�7e,�y���Ӭ�7�c˵�|;'T�QOc/M��=��cwG#�҅���眽x�^�>ҋF�@ՌS�ѫU�y�!k�tqM���CHz�ł~���>����G�������B��R�n��w�rZ��Իm����0�rX@ѱ&���A?��\«G��Y~���|�G3;��j;&%����y��bS�����Z�ӹ^a���-��+xg
�lN
/��1�xz�Z�?9�{[����2UgY��=� �� 2d��ci�е���%��d"�bX����zOZ1>e��:���\��@؏��)w@�H/5⌍p��t���n`�Šڿ�H��~�V[�(*�<^ K�H���1j�pY�N���p��;t�`�Ýe2���ȴ���m2���b�41�=T��l�Y���� ��/�D�q>���Ǉ}�gN6V�(���E��
W�����Z��kr�H�\3��>6�q�>�ɋZ4t���DM����RE����6ϔw�o�M�O�)y���o> ����o  �K1 2q���؞��c�	����6���v���	Г�7")R/-C{�ٽ�9������_