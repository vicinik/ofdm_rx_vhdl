-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
A8c/9vZes5x2ulYhxpn55bdqDdND6bT3g8/RJMb/kPUDWuyTxAKvYdagEp14rKXVcQ2K9Z3mgs7Q
areMRVmjhSqxia7+J6T/Vo0th0Y7pTNspZba99691KGC4EJVyxIFf+zpkHs6+sqXnjolcJclkA9J
yhEwvtnCpbKd9n6pphwYZ+Lm0e6bR9mpluIKTGJvpZOQVw8fx6M+PPa/PERN+VYYCai//rwmgoCP
RRAVfIDn9G2Y0zPo0sa0p9af8tNOmK2ARtnY1rocz0NOxMw8pysZ6kEjiMg1bi2vCYj4RBq6BKss
MtEjGtgYcWKvTCoaOspFYW04nn/bvDxpqo/lpQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30096)
`protect data_block
3I4cb1Yi2oZHlGPkp+cr5azo86ts0rv3sgHb4+MczDAVyD738+KynS0b2FM6e4jF0o62XS9IEdpo
Rq82UcbQ3sNJsqA4IGIcV5oV0lXIXo3pwiR1Ehp1C5oZGCxfZLsb8XqjtKpVBMBqApVXqb0qfPVa
sETled5cg25QJCEQO0Jg5IyC+jf4vOT1wHiqP5I2cjoTqe8QK1SzBq2yIbykK64xA/FxnzYbZosu
HopcXje0BkfU5dQVzWhgA3Xcqquc6+C/3u9+7LugPB6NJxTxYx3itTi8ojEp4Nv3yPeJ0srlCEUq
A29IRq0S4RvqM+fFegIGUj5lVo5SsYEqeNGLahfV+mqCElEkR1Is6F9Mb755BAP19yOQW9H7doU2
i2Eqer3t+GX7ka7YraYKZVg5mymtT2PlwpJOuGBiEFvtM9TsoKdlGNaqAOE27QWKyfSvZVTDuXkM
wegcYyKJCbKAR0wwW4JBdGE4D7fSmsd2ymebQl3oRn+07fOgdvG7FmvIYl5GBCuoue4JI3nuyO5p
1tTqURYkWpjMoz+SWEpirxCoN8TxiGLJA6IS4BhWuQmyos7or2j5YPgFphLgOIT2XJ7G+30RXKJy
7tryRWH4aPj+jTqJeJhk4qynIB0sqIZ0J6JIXWvpX+Q9EpPxyRyCk1t/oe0m2o5ohsMRggTeWhIY
YCaMweGWnrDkL2XkpHibqamo4W7d21RoV6lJwaIq8OikX4YZdRCWrFoh5sjN40koNYKmlhD4di+d
H0ADTGdzl7mOHPYmLSIj0GxtHs07x5kP+wlR9VoRwjQUmBfbdig1q29XWfGC1546RUXiinfP6KdD
EIBe5gzW1SBjZlVq07E7lMFPEL/VYYPXCFWQ/4oCgDbi4fMh5CtMAPM1arpPzip9lPvzVVUkaAPR
dbzIX8a+cFtMWlQVKQ8JIUP5Ht0Q2ZNBB6xNSsGLJqzxOLrkHUV7M0Tr7Bda7DOTeS3VpVxc8qHk
CpL1SbPMIRPAdswcuJpR/XvYPVd9oCLj4rbJtBPubqVBWgtoDFSd/F88q5FHyXcNJea4bfbDtPsV
J/GO2nLCdI4nHC5hbZwlJySLPenGeFNx7vg28jHpya/bVoCZ5uEngmjJMIWfcS6tGtkXbipkGNz9
SkBkxmWhMBPnNNd2dQ7WRfSYGiS9sVjcAmlkZpLnWB2nupQL5Dq9VByISdtg1qHDiIbVnpl1/zxr
jcCIzkwXBlxfJxfWN6seGSyxH8GrUFmbpkZ7qQM1NeMFAkAAuR89ZotSD6c9yKcEJOzxctWhcPbQ
fFCt3R4E/nsCGUM8RAaQXIsRKT46fQ+IMMZKWUftrtoMMUvSt/kRh2h/SSgaGuj0tMgw2IMbGxFH
PhGzYE70zIp2/XGbTSkFVfgwJR1oN44Hp3FbovNQ613FYdVWinG919coEUWjkHGdSSgZSEs5XjtP
XmxTScpfliMjWnn5taDqZ7ugl/K/ncfRhmqLnKS4/rh8uob91tFvJfkKLfBGZDPywb8V+LZJBL7J
/y/i75y3mfIXwl4x8DvasTdSrG0OBuP1wK7yq496X6L7Z2mk8QUdx1z8E1l+4BOBuI7LVLPHLPlW
AbOz2kYXNoPfoc6cZxpdvl0PYevecBISvtVbc9psBHpJwR960PmY3M0y8EjH6CmOc1CkEfcNxKrM
9kD+twNQFrZb2Lej/gCqlffRYx+bJ/klZ+QsGIH94n+KrKmJ6A0Hwy8+cFCGtE4yZCGLEk4hgR50
Y1pTrVWUc4nYuPTuZOl6h+rF7ypULozL4lPIC/BibUX8ZpCj6xTd5TQ7Zz1lAuRbsNn4LXbPZnBx
GpqMLlXuaKOKASZK9zecbrSX4ZV0ZqM+30yPPthTi64Ks1mrByLKj3mv+gBhvg7a5YtTBscSe+Yo
GZDOeyOB5IICSvekM0z1EI5XIHmzWu631H9agGAKAod3sFX5v5IgYMzfqc9IwXphsWBctXTuJ5YK
tFnWtxgjqMou5aVSgJCg/i5Byl0bcPV4f8jPX+fbdoBQ8R2FYA7VG5zE5FBRlhjjoBNBViDksTMk
iN6Cjm8vpwXKr27MOTg9XkqJ6jIKfyvtfpz6Xf548eQQFyYDEXpZm5HOU0/gmwByXiX3vguSjGt7
eacAG/6LSBcg49kTwQMyQcsyTaQUJehjJ3/tBKsYcC/2zS/ebyO0Q4wNYBIKj3TnsUInIGhd1i9V
ijeCl341vCEZPIRIvTmd9RZmEapSxxaJN+NAFlf3IrIrCY2IUtsWLz9BHv7vzUIJ4tqIqH8oRCNx
rNFFkaOUwJGpRP1OOFabXIsS8PQQpt2acCj4Cvq365wJT9YXtoU1m0l+ZCOmhLQAIVghDn+idMGw
Blvj3KDysQ5KP4YaZdQbLxTPQmL5074uEf0a0tGItW5z85/wyhiw5WR00gDzsa+rrViPOvI+NCvW
xRiLZ+ayKmyZR4iJU1DQWl9Lknmi2Eh9Ia45psnjPiNKgmWUDMnITgFMt1YP8rTc+b30UGcr8c9O
KhTdoGip4Ifq+LADQ3unY3L07Ei87gcQrC1Zy2BlQCREMbjJVtBv2Y6F0N9Xx6ORMVClzlZAuceS
Jn7MrkNIMS288+5az95hg+jWvpz+uSKRYu7tRgoq81FUEBXOzOnhOIBTLdpYIuJE3nkMQoF312Hg
2ss9K3yjsiBnwRfYROTJ9pUceuABN40s2bCTiOD9Ll7VCYhGP2acqIZ5E8rmj9CbVk6AjA+SO3EI
Yq1OwwcHfQnmUMzJ19TyTVMlxEuQ1Qw9iN+JITLMPtuzosQS1fy4GYPo3b9ZJHA7M2n2WkJf7LZn
PpT7RxOS12RSR4CKVN6x/fV76PL1tnmWaKyWU2afM0Xy+HDc7UKslQvMgIG0vK61fQFze33yDrKK
v0RITsJsNH3BIj8CL2QV7yG7flTCBh90syQXPXC1L+AqemVbOg/Du92dqw+ph44nv/nojqIyDfI4
+sniI6ftzvq09nSslU6QhCGNfJL4WJPriltU1SDQ2snkDoxWCRTvks/KovjhMudU9hqUAUB+1f1U
GZlU+wgRULtA8L2iiKrw9iQzddsPviwrj2it3+LWFTXsZ/4ZekdMW4BYlvTblxkmiFXfFGYp29Yo
sreVvTJDcwUW99u2K4cyBGKGog0mlOTUXhakE+/p6hdn0RHfSI3+s37RtETmqSqpnqJPzFWPX0ce
y2OuJ4Cuj2AZ4TF13hk0oQ3RSgZtATmDmFBWMOu3YN0S9PZZRlKkVNAmlPxY3hrzPtwWj0/7kvuL
YYiGi7h/Qy+ym9sOrCOdXBEeygettoy0SwdbHT/SukK7F4BNJkMcMehfiA9E2J9vCnd1bNeH6w+g
WwSDXS1YiA8sRKI+TBWDic+uFvSnGFu5jBFG4jb1X3atvJ+A0rMRKdZNiC3dcfWdyOXHosKtEsQT
qHJQmsyHARqXphQiPby6glguiqUwbXBbVTVziJZG5V4/SxN/QQu9cUomYKIWQHuLgy5l51zMtrJB
kjZuuKHogLmOVhHnnQGqOUJt/3efw65TszLRg49yOzRq2MQ8aeXzYwL86/IgyPP/v0KylnbYQKS2
MIgHHFCj5bsjSoNS5uBsjeJwfOOI/xBJCGsrB9ZW+qTLdcxjkoZ6I0RZmpukaFu5GvRp+KehSrg1
B22S8eMP2hKMWroUAdHl2ID0THKsjpx3pjxEgZDg4QJuegch1gNowRxF+jZgtqR4T65uWGR6VryV
u6pm12z1pZNByx7T3CCjQxXxp5nyvI/jQAssDr0ay14nmiR7SB2fRSyUJBGs6oFO8EfMOrTaBLZX
fe5bbBHf5SFN0yGmHa/25vOICdYMCguH1bAvseUIlUNZoFCCRPzudQwYTX4tA7xKsoE3sPTVf1fq
1R6ZvgDtaC/fT0d4LB/W/E4PG+gUZtEN3L3FhxLsxUGlKLJi9jZYSW177oWSEit7AH8X5tBxrcA4
p7amf0lwgNt8gJMa4mz1ATkUravqNx5g6F56o5cowvwy0S7MD6xtxcLB8yBpe0YrgiZ/pjiIyZYh
xBJZ2T9A3sGTNrK1olh5JAfgmkV1ey6lL4Iw2J9wt+Ms6GzEW/BALh+6n8irKw0OfFJkyAZgUTcF
qkOhJOmQaNu6268oZMER7WXh99Ufsp6h8IWSOMd9iqa/TOocA5pDYBO/ag1Pss40GYPsxwvGQuYS
wSBeyJvg5VIlSBIhIZMA56K1a3FQgInWKH3sYMQ2HPcJ0yeIAniPdycOIYrCHez9EUYb5poxMCcM
IeJdlKIEt3qSrGcI0UNHwvaPhfWO638u25HmEdhjeDoZgFRzdFtHA/fkL7wbdsXnb9ETCpaiNpjn
yMMaE7kwzdxTb6hbKZz8QMjzTq1dohbpZk5Xng91C1l8ILxuSTEcb44YSc44jJedGaOSAcOYDjTC
mBh7Bg2/Vnt4XhfXQh39LAoEVohRtKmdd6cENgtUhL5QXwDaicAETNqwDPuXJonaDHVx7tk97Cpc
QgMRyTRWpt+H3T4cLoeqhw8HGs+abKlq6MVK8C6EqH0x3EwqLCE0kqDGSyiLb5cVvuMt0EF1tnc+
5jEKkcArecx7PZ0nSRw1w+dvO+UJ3EQZTHZvSo+EMLB5hkkNVTXrEIWzVqKjYGfgJtLwdeKThPcV
wZVv5jmsKrEPzAz+1/t/SAmskkc3s+LbgHPnsx8wj9ADIHB5/0SPQwrmM1a7I38djY9FvMIGo3/P
AUneom4Dd4905sTbCnvCXbllt4eRRS10oq0iHZO3Hr0Vf0KDLzK/o8g1VthzcbjiDSp126UG9wZH
en9AEl3tdeqElvQAcgJfLkipog4ihrDMtt9IKKY0zLaQl8hsBCjAfVwSM4nCGKYlFkXKPnVhhWYE
8DNaFIGBrZiBlkxNDMB3x2SIzpSG6wqoDHeCj5f4y2TC83lDXMn0dS6cHIBIg+6T6DtpMAPd5BTm
A4fd/6j0HYnCjxvkY2cBJfUK28GWKlIwq61eAUibGLkgsh49Zo4fn+sXAmkqdzMQpxfylbgDAkiE
EfQYAihLjRKy0eNGNBVdkDojdd8K98OJhescCd0YnRaRLjtx86y7j3xYStaUWev2BDmYZ6Tqoval
xlqur0CIj6CjVjpZz6VxXmHdaZf/aEVylbB7l3Uddvid+uhSMVLKUN7JPUZltUN7peA7jv71UBnh
eEf9SZPC1dJrbat5QTaWqce+x4k6GQj1n7gkgg9iOIseeMSwlFS27hA5E+9YVgvMdfeYIKgTXdg4
vCBNBOi4gamvnM9G6SFbiSJnQ4gDt3Ozc7wrY1H/BYfSL0SXwJKsuevL19S1122vAguLIyYYPhS1
qxq2oZg7gj0wger7PWqVN1+Uh0JJj3l4wUcoCI3BAxULQHch9DI8m2jzK/zfS4G7WMXeKfV60EyX
Wx3eYj6cfbX3wuSOPaI8KGR9ossKchqOp09rFX6L800dxT+HAPMzocPKK63P6uEx9EOF+9iMv/V3
qAJ53CSXywocKEksUd1x0+Kvre70yx2CqojjMg1KcqihItvNX4TEl9hM//4+Mh6TOQxGXS3tK9CN
3dDQrrQI2tSnYzlkIFKcPwVGeZOda56vE1qrEMt8cy9upnxGfUUgtyhO/MmMfJyzelVZMioFCqOT
gGobDRYYIKT64nycBH2/z2GAEJCLgUyNwFBfADhZ2KkKPH9Pyv1NSHcaejsMYyh9Mm4wJnuZwdTJ
FIlOM0laxwD2gyrjmIrvwPWkIMtJ92k6fQavl5bQOotFLHyWVWD37qTAQlybi/20Gr4xo3N1OBBn
mTjNQnZE90T6IxTRh9RGC2aIcb3mtdGVgZ63wkOFIQNj6YJRhfdI6aTvlor1KPfwdg/903k5y/66
Qt/q6OXL6f7HeQU2p8hINEoi0eKmKwr/xS8Srr4zkdmYO7GyZpnJgIyrVHQsdwpqkE4xDABrlxUX
hQsvTIL989zMzbLaLTXxdEO1T+RBzPXo4maV2I9MHdv3PNVR61by3PtlVCjsasMfQ4DhCSFpVuo5
GltKDU+B+3HnnAWnsVJh0TEAWUQKILTwJiQeaOCV4e2ANJzARi1HfQIQvvnI0KRZhh9zVlBVdF3A
CAkzwykk+YEazdTKuPwBg3ey5aV10hBjU7OFiKOTit7U79nem0h5leaRdNRqv8WKY8NRKrfCeoJX
IWM5ZS+jSC4oZ4d0+XpC1ohxW8ne3s7Iqbjqv17sYhoxOw1B6Dhm5mDwqyPaOh7zL81sKR4RQa3m
fBrBtWvZaJCzIk4d8XbOFFYbEYz9L7AlrW4hGgPNA2XeiW+SyGl7TkomhseA0ye3VYoOi/ehSh3M
ZNyW+e0ediwQ3pFL1EY1dQiJ22Z27sbHKXBsBZsUlkHbZijvD5OA1YkGo5hhbu/HyM1fpbe8cihR
rJ7slP7P3vzdXUY7zHaY3cVRHvOKvYHbGHUySu4+HduTAlXtO/pdORtMzGXhtW+1Afgytm1cE6bQ
Cp/RnC2UFbCuMiYSE6o6iMc+nZrIV+Bc/w9wTOXXZ48/mT8gXlfzclSTudA7iAI2elkoh2cPxsrJ
qNUxz2pWiO4qVBqZ+g4HikcCCOl2vBHq7L3qADOPmM+13SAgwNEZ/GyKjCu6A+8GGN9JBHIeZZHG
S9P1ER14bLZ/pQSzEWfV7P4PlRljmVHN7zlXRC5WTRb+wE7dZdkv82hObp36/h82dOfNa+xFQ4cX
BvKxH4PGcNDkx7d+d0722zLB6qrrHlOkgIF6Ug8Av0R7xnq7/4J3F8FppYtuxDj1JFGSRCZKC5TJ
mfZoK8Cx1P9AMaCcuq1TeDGQEQX3tn5u7UYd8ToJ7OBmzbCJr+JnY4xeeQQ9SMX4vHBVBf2mHR9r
dYuBXXd+gMGaXbg9/6sBDv3VOmtV6rP3ZpVKVIY+KgUDGFuRe9rcB+Evp2YhcHHLDEQPpJs8VEMV
ODdcpWPR9vEtmGVMmaNBt3b8S4m7SDS0VwTmL7zq1oit5G1DefPwK8AcSUhQXwcEHuL4rLl3W3P8
epk9UnKJxxsZnxnox1y+6mubG8Q+a/3XsK/FODCKRXtWrwgoRnRyUD27pi5pwcuRNY50emdT+5O5
pHByiL1XwuZd1atuOHZiqR1hQI9gj9g40967a4MEqdA0Y7/Xuk8JXVjXghmjxhjC+VVcEdT7zRSb
3+UURL01eTVVLYSReOLBOIE1HBdvh2kdzwxRRgRIN4Jz4BoOIsj/f6zK/LFWNl1r6KOWi3ME51UC
kEuTb1c2c6YAVEsv0d4k2DKBmLl+ElP6RadMlVH8dCA4l/W6+lZD9w6emqV+wdFt3w+7edFCMhX+
/H6nZ0qlJ99lZ+QWKX3Aazvjpnu6iajY+t8EdJFm7Kz6Zs6Mp+5Yujw/qcIjXkyryOeVtXWZs627
FH1TgzSHkHfWDq+nzw754vreHKZcIpZmHB/+anybLxGULqiVTAzZiA6HSn22A9BoPXy6cAGvpUdZ
3euoEfNnV82rsLOBKfTO6kcxg9YH5n9bKoe71D+uD5F8QZGbTog2GLfHVvhWWvzyUhZfR7GX1c48
8MGGKg0GlD2QpqzYfTJiak02RcOecicPZ5/TuFEdPcaV29IZMcYDDaDrb3d0Iqx+kbHmF5cTfMy+
WxdYa9RIZajccVOi/kcl2Y+QA5ILFmoFjwXQU94ioL/D8cik8DqJoaXvW2gBtwAymJxvnDgp8+45
77gIr4d5QNtb5g13CRxd4cT4u9JnjItK3lw5g4EasUSS+qKzhnPaR9enrh5yZ0XYHH/RIpHtC+hn
tzEE2i9FnoJLDTCIIT0lqJxvIJ0CNQ2idlKv+BflO1Uenqx4WBnA3Fbtt7UXDNVutU8WdPzJvhaT
tfC0v9GOj7lMxjEtU2NODR9Efrxk8PxYubNAlnf+r9rurjVZtc25tPaMGhHjVJYagBj5/mN5zViJ
ZKqLfDgSPjTatu451NNJZMJYxb2nGmrmQv9mqs97stkWu9jxGcMORDHqUsqL4YVEqcVi2VPuY0X9
Q859VKS+z2MtMEiJrJ/upvQDZh9Qcg/6c5t+QP2vt3wGWmNgH7WT0pAbSiCHqx4cTuLtqvP5nyR+
DtSwf6UJT89lLDr3GI9liSyBepakyPhuOQkZm1QWJd0XHWRakwyK+zTd/BF2oUfufAiKDz/O+5Ci
b8lOSUAtrFaM8wDLIsE82SWz2+6dQF67ZyySvx/OadBBmmpsZej6SucKwZvRU0C5zi0/itRlpBQP
q/ROKOOja+9gxwXb1hxb3YRsjtSlJH+azqtqFwxPdbMQpo2CPEeqKIfakQMuYD8vVpUiEQMT9n0a
b+YLCMVSekOwNX7siJgP109032UU9+yMMgOsfDFp8vjjZjdtXXc/XrFi8dkkOsk32ppJ2xwMc15k
OecaXfGEu+vw5tG/iF4EELJ28Fhsh+ZGIwsyxmOssB2tqdh5/J1Dcm/PP7fqRBbSgzGSJ+0PyboR
7oYFNdzKA13O4cucgH1ehpGPVjyo5njSF8DLd92SzNLSn4ZPYTv8Fdiol4p4sA1S+66EP4ZjEy2k
RDvra31ts3CY7TZnQxc4ywNQtVu58BHgLnMfcRLS7+8lAlFKr3vSVRr6XrcQXuj7o74x4aPHOqMH
wPtvuEcx8IWsJuL5Ia1UFqDXvEu2FFZzgYCLZyKoLeo8/bMU+qtcI+Jx7nMGJd7InZBbTZcPShpz
s8+V5TPJjMfCrSfjYnMIIzV1O4hkspHfyU56AJlJNVagCwfH+drGkspeXaehbJHjSz1fRhs//9X2
w2v6vOT9/3tQqXN/1szJY85sxR0LxEd7lzOFrYwpA0ZnFC4f+hnAUxs6OigdAkn3Qja1pRi15Tk0
o3YHUXkxrlOLgxa3DK1VEAMoHeYcWBIzw5OePkstID+Ops54MiU6bn4r/xz0RvUdn1CuTTYz6wmX
4uCJxRrX7zLTI3tzeqcjNJKlalDd5U6NczyzM0ly0phiOIq96GGjrGo20Ww3Ws6rfjs8ME57mt+K
Ec0UKfYqPMAipxmzCjeLwUVLxsvfrg2ozjfyPv1z8gHYmgHct3c29KIogrCOeFk4+rPByjgUBTPo
zkkqLTAWu/xWudmN7J+EjYa2EvjkqwVvSVOlCoEfyME04ryg4QGDtfi9NMBXMyBVGQtROxyXQnvd
uRRxU/VEZ9O0cRWmvKGHecBv9XiyCLnYe+hBSGL1Jf+HCJZCl/oszV9UJ9ZRDJJOuaCUds3O5nG2
oOal8w9Yxx4Fon/BMdghhj0jb4HMdamAutT3WbXHc0BRXlOQfUCo40FLgtGS82+2FS7BqsLVTXrR
fKsGLzfdpcq+3vsYCIaBrklJzgbrJI8el7VlmGb4RGZcvHm+6GCYWHPip6ak4Sa6MLirO0/yqzE8
Vz5F+8knk+Bd0u39kdy+uv1A7xYTkTFuZNbE3SFV852/kaHJDiR7VVvYciYz0WyxZ0O+7vNv12Rw
4LQ3/exbf/hqpZJEQSbUiCrNVyG+y+KDsMFuqSmvd5RsqjR494ZYHWn0rQ5KGp3TPK6e1ylvYDc/
EOCKzafsQ4bmdsTiaIxTDWS4tQP9j7Hd3A7XV6iWLdZL3n1lWWwP8pZplgRZQj/7CJHpBd2U+5MU
JwDcvKjCxyGls/RXjZMUpVG9+7jP0bbci4dL1cZ5Z0OpN7NYtWoZLAwWVt0j13Vak70jGbQaiTOs
gW4o/Fl3+N7rdcXhxJxZFikV4Ahk2sOLvQAovIOczyvPAxMhhrsjlAbxGkaXpKKXLvso/fenfBFr
0xHSOdw9RSh46RSVAdTRmgrbe+0eZSSARWfqk2PYHBhiQNVf+yGQCq7qxArW2wgND4hllPlI0Nn/
hfqFINhI+U/Fcfat4DXqydoX0dMEBFKC16sJf1MrcTYevtqJsxxEAhGnT2JXGutMU979jkTC3AKF
vIR49vwq8sUaScWqBdv40ddVmLD/x9JM3SwzDpTMxh9K7EvQjVvquJzqhejie6SpNWr+0joKW8bv
O2HAeepmlDKira/OrZ0YrudKXb1rtc4dXctYvL1FAQvnqUo3LnmtkVE0H/tQ2poXgCbvVf4inuAY
VAZ91TsgvTfAG5dO2dbSpZE3Q3M03KOlKJ7OP54YcZkps4oXnw7mBRCPit46+W1zacdIbJb6dfNC
2qKxAnbVw9dEMHLWvU7lUFZA712EaEReApCo/22sv00q8IrAWt8P0/SJEc6VU96sL6M8ROtYpiGJ
4YnOhuzQH5h+btYNTYGDhCV+TXyTRdPKgt1c8nprBQQ7n7GCsdrqJ1j1TDNgvzmsCXmPTO1MwgZ5
U90o74dok9xffFdbUmcaulaIzEjUg9jrblnRi1orx9gYAkRqiYKh1v/K9L3upQuAuxy/POdm5L5r
0pXVnOIuve46pV73Yl8pRfguwoC9mezaA5Ig9XS+x7ZXPURoZ0dNJz4xMHMfG//gQUEHBwHADcPl
y5uhwNY31G0BuvMelD4oJyeMjbXDow9LXMW63aUSciGBOTDAcnhC6EEHfO+wpyK8+9maDFPd2fdh
Hfi2hRJbVPNSCkvt3/MR9oFV5FFBUwFWy7IZefDnKqZ0grJ7MfDsxwEpG1V/fi5kMvYGxSBKPbog
F8S7CGBhLGiMOhV6CruWO1J83a47Yoq1z4O+H8L61beDdSY1hLAKDkIg9ySEO6OAGk9A67MpPQTv
gFUNvq89Ui2c058bBCNcJl/9UJsb9UW5AWHbEcHHebzz2yQfl8RpXC0DgiMd1EYkcKyhYjfTkxce
/mTrw2BnSuCZh028RF94D8zA+mq2HjYrCEPcZyKZvC6m7Nuov1wYmyHaJhXD/WX9Ay6pD0G6Y3VU
ZN8dfPC6HgX3bNg+60V5UwsHlcH+t5zKwuDmI0lGAb/lpNOJH40jTh1l3s2/QmwLre1oXBtr7Mo8
ixv5csNYQ8xNKkMEEkOgmeF9gCazi6k3XZ5Yhgd/6ycdbVwwEFrisOtgDgc579udVHgo15G2qg+K
LC7UhLGMLf8dKH/XtW9r7SMfakDqmmBRtG5E7dQ/jfI3FBLBzQFfScbNEdfvMtk8Yc9mDaDv4oCT
lpXqYw8w3Wv8UPe+deIJk1mQ195Ygh7l1Q2d5lrIUrPWjBmsq++8rX4FTp2Sm88I6U7X1O+XBf74
sKCJsirdSDFjtv5y2JXBWroZ4WxpWeFL3JNA+6Uev8Ud0XMtITQtx+v82XjH2nlGfrNQQ4ELCQeN
3WyTfSzxx4CXTzfA6vfhTzRZ8W+LuaiK9Y1Su2gKgNMPGWFY4nUQQgwTc+4phj292nBdEGsBAJKG
FYLTJIttr+gIEXhBS8EtIAn80EKhDdirSrj2oldE3cCSu0Sko3Z3EJ4prbQBRlc82soSTAZHJfIo
Livzro7yTRhhvSJfK9wLRk0WGgrQ9/Zz4hAr4UMOf5IulEcd3Atvk8HFW9KrPjQcYJYxhP2XzZQH
pg5tdzICUXJ2M7evjYU7/MMmh/Q4RnNpF41uuI5QhY5wUHYoxlQrNlxkBv48lw4ZsOM+9ROXb24b
g45WEueHRWPSh6qWAMd5EfYFrubMhYQZwK6A9r4GuOjrT36T2hXLx0rRADzBhLZkI8qJqa5knk3Q
N5uapusaTmAQtRDcty7tLM5oQMEPu076nKvPBjV95ggVQdTmLmanKY1y2/K1HrfozpleessiZLdP
FMkX0P8/NCgQPdi9A0hhwa2QEW4EWMa0DqJegrns26/ORtLw9AtAzDKP1Rwit6e6dQedNdN4Bjdn
jD7NINUNOcgcqlXDbWTD8G4dilctJ64e6f1+NG4CvPglfAQMYmrPEGegZExHOQJSxTYeGZO/pHXB
JKWutSRhFexElKwhT397+E1nWr7RkXjDArLZ60EdEB3BB6XOkM+nUP90LpVM8f+ATGQ8sSba8Q7b
XlXEYH336bGEeg1BMPxh049sHL+UDC0Ft2OOrl+Echu74VSWfs6ZbbmW5QIZt5ekXLA5vfouq3YT
Fx++dX+ZcLbvnnLPsgpgtm+o8YNuCj6S6j9+u5eHmfT81Awa6RyR1o3uM4zvVt7x/HjfgFYeBFrE
xHC7PSxx1fqyFEEHdMV9XbuyEKUPROgAivMlrumK6OetJ/zjdoDhwl46ZxaCcQy1xLDgLuHnLyal
6MYCx9DW6oucDBnY6BNuilNWZXxbF4MrYbay6AdDDICeByg5UDvkFXpjUTrQk08p6iNmLxiOl/tQ
jx9u5Fi0bhNAFTm4ev81KN2Pa0GWp53YKioQAkfOx5nWYBgUMxCgxhjqbSbKmglDu3gOjcKNmXy+
T/JxsFT7VBMC3qdYNl5uk41zAAXwbjaLZmVDXQT/RyU9dXJ8D27JfHiEhKB0OWEFwopbYvzuZagl
7ZudD8K4GeAwHLH3nMm4qtgdtJfAIaZe+j1FquDANHniLDf7NlT2Tmz3CfIar+32nX/TOvmIkbCG
9XUD2je74ARmsKU2m0aoomVlYUhJaG+ErjtSlqJB11Hf7Kvi5yCSmubHDxW/TvLdi8YHMUReoCw6
vtOaYQ4ycpMbuRv5EMvmCT+41Ob2SeB9nx3q+1E9o49UqjAlFPUVFbHTBaIZBF936E4DsX9QCqS4
lLnTwpjOLtCMrg4XCGqbcVr/pm7Jlb4lIV97QNqsDegPt/cOdtBE9K85UZJA7YIKPkyK3+nxxzjt
SmOqp5YuBQx2N0SI+dfmS9rImPvJm1fa2zCckcjxYabgdl7eotEMXbjPjSimTj6TBYyKKAV0dEiN
IQRqkACo2cYEg8hf3i29Nd9UKYb0i8y2Od8+HxlxUfrzdLzu/fM/Mnc4OZQZNob2revo6xY9aYSf
G3hK3iA4Qj+YR0KDGEhf/6NDbnntFwukguKz5Oxo/ogefYd6ipAL8DxLn+nBvE2RD9le6WlOYQub
OKQW+MoAPATZ1Mv77vNbelystbpHYfa+lOEo5mPK2MFZEophONeGkQd6VHGebcYKlhgyQxMK+ZV6
LHeCgIZeLR0EyljzDCt5IA+/Zws/lO7DroqBBay2TawQJBKcE+3r9oTPuzYdnwC7dsQPcA3X6pzJ
411onm7I78WkM9SJ4jnJkCNCxulARL5p/3E/X6jepa/pIjAONQrhuYAwvPOhoZGQjItYSWrV70WJ
j3o6s020TEjw0PcKdGRmmr7H3Ui0PVMUMbBTedMiMzzXqIs0sD2iN6vBlJIOH629TYlGMF1kOiLQ
CVsR8i2B3ruD2B3bIYgRgLNI++nBpMCk9xniIUZ859N0bAj7NYF7eSgztk2KuDkLOnbZAbEEPhqa
IlwXfh9lgg+0ZHiIxz+GBUbj4TtjubQMJmyisa/4fwHwHAE7GzfkGE9olM2CVTkzdL3G1czyJhK7
20v9v6XdOxkoemXiL3H4oWqJKjtAwgXCzS8Dv7t1FFqF5YcLYRR0kATWIoaDJzguuFG99S9HZKy/
nxRTCWtPRCK5sw6vDB+ksWi5wrFmk6r8E8cQoopmgq4MdYQVBlEr2XHF9jNcDsRsi9aXVOOR/amg
RdFlxo0bla6oj7hlLhW7MteO4u4v3fH2Q0rht6q/GD68wvBZQmv/+JS/ULue6lWqumM8aS67v4CP
nCOSsYtuxNEt7d7yGQx+vKdnvCcOAn+QJv16tNi/ZI5no8zOP1KpX+aMoXFmQlxSOaFDJkmHr192
SENY6hINmZlsyDf5XNxw5gBglYZRsu4opJNeZTxFFZaTXIfolPU/mNwV8ukqOnWSwiVoMi8LwOU4
GJA7zAdb8YE3PaMp5waaqXruXppo/xMiJOm3WgOXdZthmdJdl9E5LIVjWJoAlF43372dn2fFUxo3
vGFaxhCDoU/GO1FuC8nMVUvP4VOVP+PG/i2fC8fpijtECZMahlz09CaL1jAdRkmts91FExEw/s6M
+wMFGUrfyxAEgVK6nWwUwrvislDhpJV0JlLm2iPWpeZh5sy3v/8g4R52FFQjIMF9MST6sWQWEC13
CTxnfuVPOetUilqpprAakBNfgYM86tXFxESTwINKyZ/9L+IBwDBGGQbYVgnAXxKe+cJ6vsS4K0l/
5VvAy9AxoRLHwQEd5J+hTQONeEl18yP5F3oE698SY0+AsLsmPc29eny45NhafFxH5EtGh5gOf9VR
s/mRkqzi0N7MEgQu7amRfd1e8+IVKpSk+Le6fSytLkliR07EvJ6z0w80+btxr6fkuqrW+xVUoDpN
bsSyyRTkzgR+bipCHik4Bp+ZVa4V8WCZ4zYrIZw804tWSKnx+e/SHvO+m6LGj41t/LhfieHCBQte
H161J2LYhK7ptw2nJom4HgCSo9+Qo2pgIYUk+HCfvMkDWIsfHeQQVjLTtG1lDnGPjTjQz9B5XCXx
y6741twfXGhevdnvokriX6wSX5DNkfR0609BidF96JqXdPpzOgh1JqoocoOzlrfKibUHcl39ZyUc
YkfjmJJN39bNdqiTq8W+V6os54WbehPwy7GTTdWpInARochvYOJLLEVHuN/bzdTwCauUjNaS8tbM
D9jsUJ44YbgNuW8t3BGwamh439t8HbzxClfDcuiG911wYeyGKa0hcbfMyVmO6C1d+6wGpKnCt5qL
4GuNMZ67gntFb4yCkvPBgQBuzd21LZCJdcD+v52uxNEz3aZYBjmgfkl9NMio1PnBTVonOq84EAVK
VdDTJ9TjZQAlNmGb4yXr8la0Aq14Sf9QQQaHsQJnzI5C6wgpiWfHr6C5igLLzG0a4xr0sIXRE/Y/
JCY28Re7uOMrDd6XskcZsqINU8DiByih33yqqiZh2KxKVzpgTe67MP4+npV8kB0SrIM8u9qcTwsi
BumVMoi0XqfVoYrFoDk8MxeO8xngGIjPF8SLCOSw7PTJwbuZHZ5HRqRJEekKieW4bv3FJKxmvY3J
IDC+hbATMdxleReWZJVa5z0fesUTnPPgx9w1zIRtEMcYW89zLJz44zyZdwhXWxk9PTOr392R4Jgm
CaC0913qX9qvJzzUXO7bhpTNEb+0RK7Av36M8mmJPmt7X+ZGevXynJGH5TaHWI/SEuDf6TQYAs/z
2bGOPeo6CdavElNQbzFOOeHW0IQyJUcOb0OnMx4ZwNSIHrl4+vH3dQ7zaT1jloYKB8RY6CJpeXY2
Ohtm53RYf+M/vNuZvsOIfaQVivaMySnnq+6YeXJuajHCnVCAN79GH9nG9DrnZU2ShS6EL/GBxDnH
xlINVlmpx6mqPh3vZECFILgsRsdGG27zkxE/duNA3Vfp+SVaJWQiUkEQ087i6FCPjOD06arcxT0V
rKYcTPMu9HSfB0WLchisuHOIDiHoInjsxQt1mRAKxcfAj8jjert879ReYoSBMwQ9BHhJq8UCXvdY
5d+hnXeYZiSybbZ81wgqlcU/L7HpHazvz7cppliehx/320PAxAuzc3SpRHvL8fN5bGXUDQ92i6AZ
bdXW/HPvmpgW5YH9tMCxH0sULbrgjsYUwElYvTujFJe9Eh6Kunr9270HF6ZsDyKG32eN2pnEK2rm
h4f+jDcnnHsgJk0cPrBdirPBsYCUGtAiOqcM3XtwwakclFgj6GulIWo5vxnsu12ttSwFhzssu91b
BX2S+MD8x30ewH8/QVYGXFKTnbKrfEcFSjfwxzc+1iCyZipq1fS2LcMiVHkqtAgrNWM63EMeylHj
hna3xrpuHXCoHJFYA9CGR4KFc2kE89Lp3d3tbgwvu/oeGR1T/IQ/nzbU6rMryjkYgO4gHXVHEVwk
piY/c0S2HivT6aoKxei84EK0Y+AvWu+0+50Aamy2KT1rOt89ftYdMeclqSrMC6TWxqllnWt42J87
kdfhG6wq1wYP7nVXppZWRqTFq9tYb3o45L7Be/MWLKD+mAIrvARipr+qCYLGQkGJ0k1Vy1ENMO41
YMGO638QOBOu/K6T27KIYfT9UPvmDneFTlxGqJVvKZTW87IAGoRMLGWAhk9HNjZaxEY6VCq6f5ez
WX1x+Ga+QmN33qJkLS+rF8Z7CANux6ZdtDA4eN3WHQnxasnfO4SDLMjb4rMfBtXb24Mz/s/P6WVc
hy6hzoLKGcyGGCGooRPi3VTRZJXboq4QBorgTcB1DzVj/EsdG1EYbEC+0drYDQnsRXMU3rSUao/m
lopUnmMYf9UMfDvkUzOGjLCIIR7N6VOFQCyLdiHbm8S1QWxPj5mbwGP1Ym8uux4RfLnrXQPMbD4B
rA/XeY8VgEb3lsLrsW8zuX0dW/MorRlpYeQNNoDVRUldkaQcp/VSrTZ5vulzEmUAeMcQ+FxsrKXE
aHcqlNdP1dxkwqt6XwQ5H3XlPhaFDRvdAWnSOaTO3fiidCpA3vnZSrpjtrD1kauZNaFQLmTeyQmo
dKmyzedRKf2Hdaj4qI8kFSJCdiTlxmpuSzwDgzXq7pJqha0VNMW8IgAjm/OSLKLIGlxPUtOGv1Ij
g2mprF25YizINwYVB/E/8Kc49I9d7xzAZhBcnCC9T96P7tpanmPaB96L0LJ92cpDd4HJEmteC5JP
efE3k1GTb2yEZhpPz66L148wElwlc3m5e8sX6nSfYqe2LGvo9JpKSqvM+9fO7rNHi9jX8SvwSf1L
KrzlI/GE9YQqI9faJqOmj2GNA28l4Yp2RWm2pLonIIcnXT5wL5vxkX5CL3e1pGqEWdI+lQJBdszK
ZYTKIPyHfx00MYGU2ipqxXv7wq6vKTogeP2KfP5FdYjCVTiL9iCJMEc9eecNJapomxKXadeY91r5
a9hohZw2eWYz8wQJtXexs3M4Q5Dvql633MmE6dw37Q2ruhNxZrJw8yW7W8RBcTWQyqOj/zCuYA71
gWP4v2605mHWH/RdZG50qZWLJK9Kff8lFnlQqB3FncprvPhLLH5rML5d2gTGATwaBVkbXuDw1sRn
GlbrOabbdIbwgnwv4baz0ZXbsUjG/qewu34NyjVzL10HTX0Gp3Zh49pqwO6Dg9U2+31EgxVla9m/
HzbeZhuv1qjA8/O6yKKW7rt69FoogoKEgxNq9tiMFtGnD5IkqdkJJejMoohKS4cqpAN1pULzOfZy
FaNbrc3uRHh907eiR30XU6lmxrVd+INhuqTtg2pzppJZ7T0w/mWvYhn2oLu59NMzXiFWJdQ/31LX
GvHKwHFQqlIFOS3zT4XU6dQWST//LvXXEa0D7djOIRdIAzjlMv9XQw9SMOeCGWQOl5o/yLwbfRrZ
2ZXuj4Rsgn7+fWdzvGw25wGiZwCROpwaGIdu98LWIPpsNdibNGMa9jDqR0pyeTTvdHqtxT4nlS3m
1s1LIhRIxd8ecEyMTTiHXY8KR2huPzWbI/IDAkVOUlvMJBGB1QYf6ZyYAUl46qYnpv3XFLiZBIyp
GzsIiLteTdkYw198n7bFM6v2Z0Dv6UxcRDeBh0eCR65ck26IHIxG8I7u+U01Wdu6P6e1TRev0Y63
woJoajqJhEZC5BJWojyElK7ZmBCb5n8PKxC4K8EI50CsyJVvgRJWzlEIbZ87ZiIa2ol2StQil0uy
4FWZNzblP2S4cZKRuDRLPEP4DeVrndu+jVaE2ibYUaQKwVpYUuPtOpLALdNZjck8t1AUMr2lF1Lp
7PjJ9Cdgl+1aOJCPuUDXlstEkSnalbti+gXAA81pOGUz0pST0f25PADxCr2OWhI6pUBEP0iLp5NE
kc/qApz0VbUaAtvOx8qr1fb5c53OLLOwLaSQih/Ys8mWxQ5DCHsoJLJVNsZjR2pS61e39GEkCN9b
k5KL5vQJehtw95eweX6LDU8nmVKe/smAFHg5yvsaIcDG56BobygxDJBy1HyjDRGqfkyqO8wEtNmm
+e2+dY4AZa8gqVxnwedaIxIv4ZM3erODVK0MIBVkY0nOAYeG8jDi3aKeO5DLR8mUDolx7EKmRIIX
WRiZJ6jXqnF0YgI2GRg8L9XSCJyZ9JeoqmX8whD7c2dVIVhVhxtHaoBy4jOj88WMw0I4F1SRABqN
pFQjePyYkDur63ulKIzMBJBTEX6Sw+TRdxquq9U/Tyip4/hRLKdrVRpYD3qijjfy702ocYpNaQSj
71eCHFXoWLFknuok+vvE084BjvHe26JPK3zUpFcVZAdc598URYBN/KJJRqbw9eHwmJ5oxe7WBpjU
p33AKiVqsGICGgdC5OQQMfj9i90Ryu4Zdyt6Ot5kttabNle1YYunkPdyic5ZqO0u5s0/lqyJIAur
6n7o7fZrXzLjH6XHpjlz253RZwZAATA5QJvZEMLnTIU/EyGHGw+6cvgHmcwiEJ/7ZjxBdYx7IUDv
utzOvIldTsBv5WwKxZyNihy6/NpgmCN5u/h/mlym6ePQj7WZwHK16Ao696hI+UvVF3HiMmvlWzRG
56XIVWn2Mm+kQfBSa4Ma1Q5J12aFKVfYiwDD+JPH4aXO0jLUQWhkmoBjU/BuY5/vrMRDWEH8YzLD
KMrrRTdd8BLhxFHuO71W7i8uHiwbA5f7pd3YHxzf8TpqoU2kFs+iSjpr1egmRe6pjnRfBNBycyrQ
U3mrbnpvy4HPtGCuSsklD3ASgE/AYsIHfBDtBcNerstzZ4ZfAgLwbXnPSB/ZaTyqk2iiZBEUeUtS
KgFSPkTTK+CfRhR6Y5doguPR3x1Mmd++z+zwCNXWieiYE1zt41yYj4sIqoxCa5Hmm0jGvRtCFUL3
7DX6R/u+sZj+utgRpHj6ADsJrSdehQDbnH8Naoc16ODJFp1Yzw3QCHy7197H+5EXAjfcvYaeZh76
FIr6tobVQoTPi8lpgYTqML7+FRiOpsLkwADj8G7Rx6z3D82RY4gE7iVsULCvjxdr6JMsoSMdO2wE
AqDjuxVnlJj7OIALJCdaV31qRbIsEvCcgTiFhR6ry4RB4MgpsQ31Vlt/OA1Gehv5fEPoD1jk+m8H
SJKYnEIfWGE3lfIxzZObzSmMLjmc9TzbX3crwRx/A1bnfcfX1EnT4gTurv2vTwBO6xsiiWdAPdBh
BAy04J3nfdWdLbvrOJWFt5tYMwgs+3h/ozmEr+iXduu4wlyOMjAaegB1KqowUPOLfLBZJt6GO+M1
rs6BY2yuuD3HqYFVsNznoFVqNK2reb7/6pIMFszgbsGjJd9Z0kwLCMUUkyjGhuq7d/cS3vo2jZeK
DR9OYIGdqAHi/p14eReTv9MRYbPQcrlWb/v0nxdljftj6uhyoOeV5BOXt/Nc560w/g4bTZkgl2JA
3u/HKQRGUjs0J725DRoeqJ11Nd0ioDYACJfQx/6pSq4/ZADcUz18CgaM9ljr4yrtUajnM4lQ90tx
cCv1qru8gsZzp2BVl7dlmHlJuqGKk5cZh/MrYYUgdSSD7MUznGa4YcCV7xdgqt8DffcNC8wTPGUw
9NeoKjKxSvnMxg9UHXFILT5s4KYSn5CkwC3wFVcluQJz7NuVXpDBe+gd4fDguaKbpBkv2kOAQ/Ju
TAie0PhEIt7cNB4bO5jsEdCEjzGA+XV7dEwuglo2zmiCtx3nV21us+KiqzkJsK21hvo4vP2QD0L/
Qv7ONkn1I2soNvTwmzfnA/2wdi+f/tDOAfTZmHZHBHUx3bGgkiFJLmRMRhR+hYbjkr6ruulBRzZ7
hkXwdUbSmrZnz97H9tRdznFnsPVMu2Tj+37odeHitmur8itts+77k3m5U4+Qo8NdwM01sfBkZnMB
wju1DnfB5+j08NKwDE7rlqytxRAOMIyWIq9L6mTfmUJN3TSUCJT0UTHQZJKvUXwN9u8SqEJatEYz
VW54zYjNxJBQ4EcVr8W+NA5aCfUQz71DDfTr5gB7qFgs2VRGnOyQaS8jmtKde1cnkbJ8ns06TvEn
IJ/i5q/+t9P9DLlJxTG5OwjcfKLbUtWps+eZLKXCpYGG0SjRsgKxElv40wIf+C2WBb1XmqWV8qo6
Vn9sk5wmrv0U396WUjveyqefAehDBg2xyQ1GHiw0Z1mOOCPzhIAa75aMcJFIk9a7vgRusupZ25Dw
WDILq76oKiKfm2OYs5ihi1ZgnHVljjWlNcFpsjkbafU5XK9Q4SC94oRS4eeUwsUzTl9B2ronozzA
yiV5GCJZZODLXyXfU87eMibq7Gk0zH/JezCzKrYIC4nTLGOWfWTkHzQUbuqIP/B/MNWAYcijDhuN
8a1I+jTkLfcGuAWoSKjDVwv7rQG1zFu9qbahfxeqn9IMf4Lpe0TENFtUAGv0C3xiCYoztqzZe6sg
2p5mpLdJkrVWhotXzVsnnddo7mCRFcEqKxm8U1amy0ChaaO0x5K82CWI2h/txy24TVwohKZnA0fF
xx8RHMEV39MNRT75c4Nx6VRrnREPqiXFtV6AuvHg4tyNLwhk3zvRMI2/1of8dw4mwUk18Df8WJmz
Aspqs66/2+9rIjypSilWwZ3Iq31+3B2qgLz3MPvCtdpIQwTJorRFqcKH+TWnPi9mh83Wk+jxCm/e
uEvsZtWsqNHmlqXk5jcs8oGBGYavnHUEApc4FBz9MghO/T0QUyjz6rMd157P3vDsudw6yZ9keqVB
AbyoaqjtcLdWeM5V4PQ/JqS5jTTnHi9xP96/Z7NBFLqJsCynMQsaY4fbT/65Cr8i8eH0FOUcnyx9
2ny8ZMwO+rTkU91KuFrI/UCBEg0sQ5yGqC+acQ9H8nwiDH5b0tjWTXN1eVpca+4V1jFL8z23xbCe
U4wUwU+NpyJovUQxhYb9F1YWC7EsNz1RUB8I4oHOZCPfJEQE2UJoqTwOVZ0iDPxwM55p28seGBxe
48v2aNhormhQ4AGVebtK+EaM5YgaEowcaKg6SZxH5eydJmenH4bb28dFjfPBjY9k1TIU0Q285uSe
5yLwq2dj2ANt/oYF5WKJw2+ZNG8fZXwjnvpcI2LhIFhAY9AFVdvl1bh2qd7agGNyutlwxUVQa+2D
r60MCwFTXmqfxe4iKghO91UDMptCeIUH0EtpO/pOsX7kPXufPlX1uH53Qnxhw1wK76qZIEywZ4IE
hyl6xgw5twhJwBItkCvuJiXG7Bx1mZa5tYkE/qmdal2anYiNm1hgh2e79+gSHRjUl+GpDtfecucP
iyaH2mLmZixgX4s1UVRQGXbZRgR7WGNzPRGtN1Puev51kgctMtLeMwgGdMB3tQL/EnQu3+6oonYx
o+k+Bbdk2UctrWgyjk934hpgbVQJmW9nY8hIMM9fA6DBVJUVzTwBD/dPhxCJRGD26vjbt+j4ZkSG
gMvGEJNg4Yo7RckpOF9FogfdQLG75OZ/XMvAJ/cmZlAjOXe9xdRJLoeWHpPWW6AWkolx9GAfh3qS
jqfFtgFCG+siXs385aDAJR5K1FbUujK9emQu6w847GRjpHVVEQOPHFZ+GBTqw3KgxMUIZGHFb5BP
fhwl5qAo96EbbQo/251TtkfvyszVZk+u9CbTCWdk7SJ4EWSNCVLVtsc/HJwB0GVZRKnEa2aZSya4
JF3fE6dyOfOMJlUxob20ApjJnnuJs2PprBvg5j4f4TSIhrh9ZOXpXFEfBX4YjFGN8n+r8Qx2cGoy
odMtKze90F0ayH3e6HEDtB3PJ1bN8vsBz0KFu+XSCBUHmsnRcsvtotmlBbiFDauTBXbEsjVHkfUo
riNdqD8RH0KKBi2mkoW43sTDMJH84inEJXGSpg6NVuN79zEFJFMNS/3Uvq1nvqLdYSwAl6GhL/ee
/ussPM+Bj8ow0iKWwcbkxEIsq4FHDB/HoDFT+t4Fjcu8jvw5tWqNgmObMgaMERmqrlYzw3iPhbOV
TxQTipOtGKcPWIwSJlAmN+vCPINJqluPjsRDkOjDD1oMsS+JZZt3k8yvfRq+vF/E3POwjKC4zslU
xPjy9A8vUshNAHb3yuCMeKL++wQjVY3x7GGX8+7rkNg6ilYoeJ0SN8K7RR4QWDUZR5JkrNHNpy5c
hdASHwe9ctzw5ZcjQzKVnlLAEZ5ScZxqrcbeg2t1BOIIt3whOrIsDjtGnwBaPLnteGFAeUhUhNoZ
cPspgpKjEeTwQgW7pgUneSJsiBzWvlD2Rc2XEJNx8YgsD9yRdlJYLeC9cevMXH+bsmq9GXutmgvC
Om4SF2CihYuEFvv9f9ZgTFsfSlbMhid9iERyxB/fg9SZ5QBrNFhn33MYHGsX134JMq8AgEAxwSsY
Hhw4f1gMu1NQSyVzR8mTM31hTJh/OI2BCm2hpuX+aZwRAw3JHHdwzniMl9jOFg4heKRpE3AQHh3t
dmPdgGTm9+MuMtXOrIsY9TTPfq5UCB/3lk4JgLfS35jRFqL6O54dpcj6tpiJQP8Vxxnjp/zO3t8q
AlxZ18vUQhVwzEnQqazsFi7cXNoUf698fTCactp8VzaJr3o3+j7yHpqlN4cwsDwV80AmQATXZSRe
+3WVVEl+wVqYiLxWfZ1m8BfpiAUa/kDS4DIuGsr2NgdQE6YSreOxhRYLvYrxlTCijwof77WJKFlZ
8PSHUHnZVvdscu4eRmqHPQ0rvg+s/RmlypnoP/7yO7X/JReAeslgHbjtE+vzcCPwc6+EvsshSLDH
F6OiN7P7tG1EfgWH06FuqHJcz6cVOjG1w67SZt2oXFS5ZNBRXjkNE+ESx6ewq0E+lpWoW5L4/Rf7
3GfmbJIbMyrbSousFi1fmPPOBN0KB2V4aGQZebO0oOLMJTCc0nqV8ZN3zOQgsqul5RoGE6ljiRmb
ahZANM3U9YDrXfzLMlVCdGfZD8WG2Gfqq6m1nwk9YfV8CChrHbAFgpy1pOgKDd5pDsfWIQFei9Yt
Wnlfkuqkxq/o0C/74fEg6CzMWS5aklEsh2oRVxI461JQiFvb1iaXnSwBv9sQ/Bhh1tTx104yn3e9
UTSkIsWLeAOAD67X9iuZsTsyfTCl+/uCfU+bm785d4EVQvWnA+uIKpZa3c1u1xyC4gsoEIZa2ROg
Xq1BTXec067OSbtPwrRlVtzNk6Tcv/inZXiDBIJ44jvvpWbUKY3nSCBAXxvBO2RRdOEya/GhNNf0
AiQlDiQ5Cz07y8ckn3OPF7HYIaIOAKSnrDmNvCkZpEGd88R3/IegA0BLPasMBwbuBtm9IwhSAPSt
vZpf7q+gL7OtMOqn3hXTv65/mNGptLgsJN6rb+7zyAzmxUttXDCa9EGCUlJ+iyurYHbO0y+CM6Mj
Q3xJj3N30MpP3UiU+KFdAwcoXOxYiOgGHfpxd1l1tEK1Fjj/6P+3yea69xj0e61Pte7p/OkXZEQo
Nz84PyTcxl29QKa3yOfSfSdny/tPRI6r3YCPrTzdRcvT0Lw+nJ+N5DYdr1xJELCO87cC6+eVwHG8
YvWh9T4Omi3XXaF2g2JDvgdRWV6sFoh37Vq21KiVvurp6HN0I29PJb7LW5+E5VB0uh8pSHuFWBKw
vgc9JuSnaw2kMbWA3uKN9C6xKsrLR2sjDralRNUAn5GYrE6fOeJGpxnSduaPqSVRIFqFQSTVYCcp
pKzz7CXcvR0z8VCLp4zt36Fh7OPecmNWT6ZLH4AgZVEjur9ug6ROTV6DKA7cBjZV7mtt/IfDF2D5
BVqOyBaU1dUqFV82UXqdCwavewGPjWpwP6SAajxKKocg9lz0UFQpDbygBFHNLJv2b+Oi/1oe9blr
m+S3dS6WgKOtCBGIArXJ9qLEo3pDNcdPRqW0wXXD2VepEQRwxGYSSEhchlNAnJFZcQb2GcusFYz2
wb8xUi/RSmFZl7F8h0tR+sjBq4ol8m0N1dJLtKJP1yRBF5jYNwL8oe04xWW08nvCJTqOW0Ihou+R
K8PnWLcMQWLYD2ENUog8QveYlBseNPsJsmfPKQXmxxBh3XgXQv61OU+4Xx4HAzFWkNSjp+6AnX/+
CIu8AOVCLkDlwEHYriTIxw8QqTXGcestmyjdcaJNovmFBvKI7Wq6w4dCEgJ3/lS03bbiMDwQz/zU
5CqrTDwt7/rCwf5uxvGpDbJKEutJdp8Sps/mM6wdpGlfrPfTjgIG456iT3VpmbQB1aYCLZNmPTw3
BaNXWXDoUFnEvjRGFmHADWB9JxkTB7d2480/WRGMQMgkOqSHBGqXbpMGOPijnsCo8NdX8JBgndhi
PraL2VcyedyauvkiYj6EMGhGILu6vQ062HDFv/JbBFokT7GfcwCjxrXYdMLj3BDaF3oMOgqr3xKb
+4Lq/ax4h3wD6gHlFIoZ4Sskartddl2hK22Dk/03CB2bgEA+fEqGNmOx0YV6gMPktPdZ1dg/pb+1
kLfdegZWumucX0SQhIimqcr/Oc7KzVQLbmNfJIwCHzbbjyfLSihGyoU4zbLuxDwO39umgbNezazt
+64ZdhTYGzZj0JMYhgrsbvssK+Axto4rocI5t/gRiqVTcrnO3WOz6lZgM9b01CgU7Fhlbk5YgQgq
pG8g3RdIFGgGMl6DwVsa1DibUdaB0jghKKt/RP258W07k1FJ++Issc2aQ/nc4yTRdsTR53KTDl+m
nVTN9kZHA8vfX2kqIdclECNmk1VcRmd2SvvX2kaz2/9gr21Q6sfNmkeLvxd+7d2DxsPXl4h54CZb
bPEUVShdeyJmOrBlx7CwXl/4EbW4A6qqIzv7kdzvWTd80kN6KTmZ2kQScxa6I6tFL9UGm3nDct4d
+46i3Po1XkSDjaYCOiGF+l41gMXX0GSoChhAnfnftwpYT8Ra4SyJ/NvUoylbahT5tUEeNbgUw3YR
IFMb7vFiHfI//WizyfRSrxaLOEbG4uSQHrrmzn0XVln/BUCKyEWny7MwzR094U8M1YNlJz2JVcCV
iU9tCwyIpUykvnQEuG0YRRsygI00KmglZSKF0RWrqWNaCwOAOnYuIzBPlFxYdMzFoFEozXbMceh8
4AUWSONkoz72gBZwkAJG0P8jMqDBFAyuhzuAez74kseSCnsu301ficv1LQb9YY2UTJiPBNfQqgeW
clLgcuANVBETjpTRokGiS2BZAq425WBYP3bXxwYkd7jkmh8q9otG5/Lk2x3RTb92MJuad2NFjnmO
TKT/j6OVnQVVawTooZHXBVI823yFvq/NwvSOzuw8p5hx0BGHy1M9eyXvOKDTk9duBE00bwRXNGXy
Z5Qo2vzaDnc0IEwahpEADp+n6f3dRz5zfE9F4vo3Lpy6VokSy8CG1iF+FZFXRkMTJEYFC6j4HWyk
ghrRAuMwZ3PQgjZSImm0U/wTTQaNf9l9BmHTAOg8Rrz3D7RnYSbVNQCtm7qOd1LWAmVgSCv+ZGf7
tUlYQpkjuvxw47x1ZMV5oX0wQKK2xb62kMXkNrNvUvA0C8nbCtuKKk1o1I68aDizrgdXRdqQ66yw
Z/rRoozKQHTjmG8Fe76bez/mnHH3MciiDyozxECv/yJfPLOTfu0jGkWpoaC1sB/NswvzrNESE/Yg
yhXkUEE0tg0EluIaKfvf0AzOuzqZC4kksYInIPcR9XDSdm2tRv6S/suyenf1IXSplPMjEZ+uftIo
7Sb+D7mtV52Eq9D5HC0KRhP3/mB8wN4/hmQKvbpMo2KlshMlrPTAJjAD//XbxTeNViC86df49IHT
LZ64NeKp432qGVgQdA7yKrugd2QulkPMjlT1/V0rtXZx1ICCxL2Kh9XhlluolhGhXPXEc5BkD7Vi
U/x54vEbUB/xz4VyxdG7Gax6M8oT3CZ+ZQ84tXlU7AUP2pRlbMcr2FuWnm+bNyUr/A4M2e71cmCL
Orq2JwVRZkRrwVMKTbBvRFcxO8OgE3oxVolyn9XZQZoBvPIoBct350HBs8aPOt+BkMHuOhQVvSXf
gpOEe1Vy2KoecxCTcvmpjSS4P9Ad1fDQGvHsjLfJmN0OrCZoTcWqAi8dnVpMsn/KWPWOAaRkYgzl
WdHs4/dQcE/xLDX4GZ3g1rwklplFH5P+7stN9qY6NksOnW5w7Ue/qon1cPI3nBpDDwiNoSPT4FMr
3d/9X9i1ICFm+51Sp/uydB0IqwB0oEJ74ySKhP9uiX9+ygEb2B5eJyy19mU7+kbtQtfWxQmhZRot
/BpLwlKisRVqmEnJOOI5cCoykYjt1ZZ+SmoFDfx+PRDypU4REgzSA1NELrsZrAD6twGkTV3hjeKW
n2WasW2Nch4i+3fofHDWH1GS30ns5Omj1DfKjD1MPcJMn2mN7MxoEvYI5fnJwgjBMfAmY5EoTfyH
nhj4XIVQ8SQPLZpYy9sIt0OAYMzymsctGD+A7PdgubsibGHr7Ual0oPg7hxEtrAaUAlbtcsCHKpT
aeq1ArV6eTBDWKiYbvgvGrabH3nojy5KalQgJ0SErnOQ5Tg4hRjP3O/khSeb6z80wViIW6j4DIo6
qeB6sqa5XonUT1mTcFWoR2kQlztPYVwXmu0qo1jE25QlmPWLuHfQECoQj6ATKFu8rmFefeO3PStb
zjfW+dgkm7rhqkKNxGoMUnV5QFW8VpuW4p8djso0rmCJOwMlpwrhr6cZuMaQLLlhsEXlN2JV+8To
oS5ZRxNWT+BMDUTsmRrZgIam4GUf0ursGpAq1X4C4VLwyWYhjpRHMZo+CP5R3XSDy/xYOe2I39ad
12Yf6qtZpC1hYRubeVMi+pKdg9yWAIOwVS/hS/ZMGrpBnGYd1UUtmChfQrqILy2fntGkiB3H6Fw7
zHMZdyj11Kdm7PXd4ZPkYCAoXBvY3dBSCObRuKop805U/TS+LjULm4qseog4eTsLt9aFGlURKk/2
adlqj+wB2h53ROKfcl5a/+8FqnACxL1/VLWzNxt1FtkEQg1LI/ifY0l7Bd8P7+uvwvNqW7oamkgt
RDQU3GvSS3hAds2rUKDUo/gIigzjgBtVTK3s5uTtv3moHDS5RohoCXEC577Ubqi1EX3df9ag8X62
DFt5hNQ+y17FqmD77ac4PsRTy/EK9GSruZUrqvQLp7GXD2L5VyniWsBtZcCkO0Eg80AiCRFwGOwv
b/evYB4LiVRMIsFiUvMldb9MnjFZxTagGMOw6+cHeU0pevqMDsFHeqEOIeBfQMd2pZe15HmHFGoM
gwar+3PivBNEbj/SmfPHh/ox40bxHI74lnZ/W9HsgU56qWRid92Wuuc1xTwu2kPDPtrfapg1+6x6
pnftQiH/gfzVEVkPgzJtKj/s8FGEJWFgqbSruACWjtRVadECMW+t/nDH4OZ0Xphs7bsRwt3rS4zS
o4dCP1U3jxvFBsSnJsmOboOoV5Z2psoO7Cw8OFO1ds2PPukL3WPWc22PvmwBblOrXdjeeKI2Zymt
g+9cJw+MPg2O1rfJJVyoYB2n1FyvmXa8DvYvEmsjkFZG6wo9NjdS5gh7pTQzIoM8Zl0N4OTIi/A7
9NkyoSlhSUVoTxqU45Kw1R4EdGjmC9Mu5OL/S0dmm1U5U4MnmxI2LXbOiCA0/BKTJ87l/1SpMoL3
FTQssKpXek6AN88La2P65BqF1cPmSAGQPYRhe8jt01opPQenLh59/ja889Zi2gE8r1V15I+mm8Kt
DVAkMntXn16F1RoZpmCLKTocTDzipUd5IOqhYvJRWyNgTFonGGdDH5IgdFIf1cRJ2fNJpzhXYOt2
5ulO5w+6S21oMeyd5aKhB42VnCDWlrUFWjV/m3njl3TKvlSKQvGgEzU7NOHxJWwVGKy0eS7wcNxt
jqweu0BuV1PKFdwnX0zUZ5k+Iij0FaOeB4r3bW9O/XvbrZTNHVGwjCFMzXM5vxBKG2a/1heXQBsX
BYx42vfBJg6Y8vHjDOdQKQSD6G2MtW7lYWyvDqVA9YsN5fgrbD1EeA2Cbyk5G6e7zqCIu34yuQWK
oHrCvVSerWp5uc6beZtybYQz7woHRccOhmqtHn3RY8khzOD/yT3DrsfgANOtajppa731FhcyDvb/
GtnBVhSrMm3U0usE5iCwR5I4kwWn1vlUNMeICF28de19ZfqSFx0Ug7WDhckPRlSwE4ex5/5zdaBz
5fg1w+yl6sArl13nZsYnxFmHEMEMDs+Tt/wDZz5BLFTCltgbE+WUNRtMUeYG0pcAhZkABYWwV9wL
IB4beG6LPHYgjrfGdEV1rnO1uhjoA12ZoocNVsn7QwNgzwhZj9/0nmsOe9T4a4S8KZhl3xc4cCeJ
vDF/EirtmpwaulCQO7WKliAE/EfpDyZkSDmNrwa6NBqiQEHIf3oPojJ4pfAiVF0/5LVnJmO050rt
2onQbikAvNCwpok/CRxKDBZ4oPhIUOyVN5mPSmiwO3W1cbu6Iw35f0X8fbJDwXSHKDWCUQVRTy9P
CLOy9bCmmfamlYTU13r3jM2FTGcF9W7RPsqhNRIjrC0XLZSL8UjkTnOuGjRGIXpifgxbaHcbhY9r
TYcC4IwQuptzVmanTPJ0NgENGXekblkYWxbPn4HA+KVx8134Np3L/BL2CBkWGiRgwolYO5QrqKsZ
XvmUfI8oTLaOaBPUJH3zuIvPMCRlPBM1/b06s6SD47HovlLm3PN65XDdemJ0nwTc1il4nyPP39cC
UYIS3mREU6iillex/M06WOsa2PA22nrfUhnfv9vS2VgyEqAgbsW4cwd9g+e2zcskQgMA9RMwfxaY
kvL1EoeVzeF10SO1eI/Lwi/B1bvoxRuyzfNZHgfirhvVf0BsHftplE28uj5bO9xhsSG6lT2Nqdqq
tbWdd8Ft131AIQbYo9uvnjP8HnTu2ByQqo2Yp3aB7azbei3vu49pgZ9IWhYXiwRFaAU36ktj2g8S
6iXvLoh6XYxVESvoop8SQMvVM1PTy3hkuzJhO98UeJmfVFtaXs/128nBCm5K/BjOh7skhMHpYrcX
USMjmeGE0T1thnMjg5kykJAYNQbYNL9mD+LM7gF/CByX6jGg5MZS9ZxFkTfvIJw4oGfBjqZY7ts6
n+7gTdlMDx+KV76g/agRndy3K/OGS5WQMaprpnvYNI9+zbZzSqbj3XZV7xCr6wz18HJTxdcy83Wx
YVVD5W+taCFvEt9kzhyxeEZ9B5Z8+ziKCPzo8gnXUp5xbV80lxfSVFNUNxNV/eHmTUZunNeK0Tbx
1t95Wd8XJsXtDxnEgnuh8CDI/LLnT26+qZLoiG968xV1kpDiA0fWSKmyadP/p6BaYbrORFIsjyG9
vYyAolTwAkg8zUUEUWPDr2GMPiKtc6G0M+o7EjxFBJPoOzpVMsAOdLJC+Y30xFN1tcapI/fWdxI6
sMMYn0nWbcQIy8cZZRIFniG22sFhfXX3KvYfN6qdAk4JTy76EuZneiOxP0FZWbcwXdAh191JPj+j
jdxrZFO6GPCT2IvK/HwoRYb61e9BxyX+FUSgMTrMdqPw9k59ODD1TzylPG4PA3ONoI2YXPKVcNoi
G1dCxfU1otvByf9RqSXUkQvwMXSuVfBOGcXWj75ArDNfqqlkWfmMAPDBijOMi+TZkpVKLTbkrN3+
3KUus6hh4kg3S8+MbEjYYLVewuX9HKfUzXUpp1vqc0ajIV4UE3L6exQ98vWWmO3/tPw0TAngnHpy
RPWF20yFI+KIFibKba0VuBoPaqfdZlNAYeiV0gV9JBqpSWMAPFz0iRBdn+a2+y03tUQZ/zFyzop5
a/AjF1vGwQOUaao48EOhv8xqXicRBNBk58A6DQi6NqO1nWBoYa8K5A5EbkovBKdOWBwcPB9NQiMZ
6qLaNhjf9UVK+7bNTS5ckCjDcvG06FsTyqMTOaCq/ibqOuihAv91yGuaDOfXrZFyvy6XLXrgTS3/
OOqQxlMeTLIFD8LTGVhaBw2/3XrCbNr9Aqww/VqTI6Cumj0NrklcQEk5Lz0/YQQv5dv0kW9ePU+2
figWTGmZWrrEtfZHFs3Do1wmIpK472LuD4GAFhQq4Bq3cPyfMiv9qraMdvZk6Nq0uKURh3dV1vnO
nRbdAdCFlZ0qyUFIZFQs7QGy1GbjXCq/0ODpdnj38+HBoL9rUYkyHDqleCtyKamAX/LPuTd7zPNf
B6+UlW84dchyS3NBH+uNBeZOcC+AwZezJTbfL/KAyKcCyNGFgenyXjQ7U70yyEdrykKAjtSFOUtd
qh5QdtJko8kE0jhPJ0BueMqAEVVdCnmuEW+ouO0fIZh5xCM945wjL2tQ1Zox/lb4c2lV4cQNgQS9
1erLebpAXHBra/4s1AoRlxiXhqlqc0Ye55Lg8NI7DyFTv/c7y7y/PDhbiTfOmozOQ91Y24LY4pAp
JzPPTbX29+Az10ps2oksmFDiO4fWDM+6WjQYjXL0vWdct9HbYfDB6MfL2faN74O4DfZHCAqxorPZ
HuiuNt9NdoIlJQZSb/igIHZAnbZxNqfaLpBbPNWbVwfT3HBqKMadIWIKw/asUAbeoWHBRIsiHzVd
unYJbfbNdJ+0cnzFigZQXOzrUt9bH7Hn/o4bgM85xxOzLDuWLZIusEXFCFL4S2X6Aeg7MQr8R09n
FDNTXVgIC1pqsS08BBCvUKYHRW8Xle+bDqwAN3NFgeu3wxN0WmuaJgdRdJtCzbREk/0grZBfAa9J
c0WWsAYGDsapQ318EjHLAcx85qEX/KvAtYXP9sL+9e/er92c6m5qWHlqHkxYQoQUQ3k+GmyJtrmG
hhO09UTR4AxRi3iByGX9OEECDoVHnrKAeWn3CzcFgQ5tDY5D3zpwFNSZBfNhUA8tzP4RxKVqrC+w
OTOUNCKm6f1apzOg08FSJifS8Fyofx25ExHE2CIkCAoK0ygJBuW8wXQuWunfRFj7Pg7n45y2ok4U
25ndCwwHhRkcxJ2LS3+EmxzKYD4y0N6n1Q6KibQe7wQvmkPSstFmuenRTbWUhNrePz4fu0ublbz+
6fxzyQn9B46hUxuTxi9/gID21vUSb7fdCaIXWJdN7Ks45p5N2PmOj2Z2L3iMORtzwid6DCfB0oAi
vVgaJjTObBWdm7T5yQ+o2AKPk/y6g5d3yvcpKRJga2360huUq9JEu0PLy4jvysghYfxZi94t7JrE
lY5KwcLlSE9LsjuBbH+5fX7QZWgMcCp8FL1h9h75mC/uAYo0sfaK2BA/uUM+9vdcS6a34beP5W4/
a5Neg2HboFH0yEzlrzXaqX8FfTJeNS3zD6P637detDhdZHiM09obxAv+WZDOuWrVVBHvlvYiyWIM
k+WKMnYTndApvqmFh543K7JguOiuawZwQ32bIvaBiV8nCycGUkR8MjZPFd6FfpE3/viuXeBfBwSV
m+kRbN+/sPFBf/WJh49Knh5R41YtEZKXOzAaKOwNAFVmrIQhQMPQhM1+FyjjqyZmgwXOSTfdWW/E
qu/r137PGqkPb106ukwiTBtUhueWJAOTd3Ei67g+TEbmyj4hkrmfim7NV9eEocYDp5HqShCkA6us
oYH9wAKgXmPykpnl+ihiPWwsVirw3MbvOkhhgMxOgXyY3dQDHi/G7zKV5/+v3oZA+xOSRI6HyF9k
fzGz3huApWAb3PACsvH4eJ8qgPICyioHMl5qx08XAD5ruZpn3TjFbVqh9cKMzUlK39tQDwDKe26r
wd07alCQkzAjbQBnfmxv9Ix1LlfI5WPJ11nMe94ArUmgf9Wf5Q7ntGkTqJiCX3xRLyevAzfN1oMr
/CcGQUcLbsr/XlFwT2ykuUwOT65L/zOcwQG8gAop1RzV3mEICJZ9q17d+IavuAvo5mlip+1zxs8C
7n4ow+KNx1QDY48LUgQZeNaNDrkC75J4bIKwhmD+iQXk+IZmrXwtH596iSNu7JumdWlSGMQVWNGL
aF07rj0FgElE9jADaDhC1jWNNEqxCv+21tdvgpHa9YD3VDT+ja8NRjNzI9a8g38wFnBSA0d+h8jN
Ber2LC0MNJGg6Yso+V0/hy2i7HqUqvjJUL1oOh76XRwB3uafRwljbv4zX6UyhTunuioDzURhjcjF
orfP0QNz2rUsx+X/LHN5LyB9bz+8zmwOUun8xXbD7zORoNwPSLKAXn+mdG8RIdvzN+YWaJ8OYtqx
5XNyOJ8YuPYUWuCZtmXTDK/wtj0wW8heB4j5stW/pY+ECMiQ4q6dFKui4XZzkpPxQz6trr9WFmfy
ujHDyVISj1CGAL106AytfSYn1XbrJ+ORnxxNynkaACn2UyQfErNSlBOfXZ909swsnhULC6RKFhsa
BShLCea9dqStyUADSXtHSfqkYZ8OLt+f8/dfaosgmSB9Cr96D4S64/kI2qE7l+ZNFCQB1tZXABqt
HMq5EYZGCgBaF9qkZKMhV93aqhbyFr6be55lF4hY1Qt/szHoeMGqnlvjU4mi9HkOEDjZDVtOQqgh
eX45h8OJ9UeHfvoXvu+ehsNWsvqhuk1zDCm3a1UGX9FdxXCvvi9bWiXDCs6GYphuqXeG8HZdAfj/
BUA3CETGP9bRizSdU/Eq+rvLXuyV7bSexxkfcxiPvd4wZdx9gGA+7qSW2WDswmgY2mDp8cjttpQA
b8i0YM4B5eelBfKGrPESDINWZUC+QwH8ht7kNLa8JAD8/QoiVTWrW/qpdJA8CiMF8BR9H6OpE79t
7Lllh/P6Hw2mT38IUD4Oepg0r5qjO5XSWKJT5282BcMJ2kqQ6A3XRUSWQiJ5oq0vS8GCgQfMVKIk
coCD4pUh4fa+SjkY6viE8rEm8TaOiws0KYR5xJZOywmz9uq/xDNmXoeWT4SikNEjAR9DAPH6/MKq
KHd73hZVwWl0iGFSIMMMLYJFooTDlQSFaRs5Bssvyr5EPUjIXzsjcOBHPDQIUq9Pkl+G+tja4xvb
yrraDpSDQblqpWAdVF6drA3+VsENf5gblYnPuc+5NYntEXkEOXI4g4zf5dHTeBw03LG6+TdDDO17
2fKcppeoONNqIrbZaBGPXyfEOocpzJKHF+8tZvYN5/DKTwBfoRhoAr038CEa4NcZSFiSqHe26R5t
64Lb98xFVRBUD02a6AeWZJA67HltWEdJmU+ceLPO+yxZZ5uxfgAKZI7u2mZRXvf7opaDyQVjhVqZ
G6ffWdIVOa68EqUCTYh0ay71U8vtzC2ehS1kOcWTRvEQmlklFNtrGWqzgFkfp/A/S6YFuZucEdUv
AJ3DyX1cBk9mF2UMWskLEKz3f54R0q22pFK2fTFlOOFhtRLVn+jVOQsSQAl0Dil9GzZZF2l1Hb9e
uTupkFV1AzosP4BcxgqUfVGQlwMtfSEnM0bXz78W6c1gIx0iTt6AAyxHFZk5OlQVPyRQ9oEbC2XL
KLpo2YZinCBMfGbwKdSlE2o3cwMvJFS0SRbOKO1G+zorcYyMz66dLoQ4RZfY/xzH1YYG3L7H/QMU
sR4DXZXV/Fuhd6ukmh2NrkVrvh92O0gH+rLKDPKrAYIhPoPQHUMqAhBDlJ6lXN/ReTPReiTrJWpj
vlERs1vBQVJs8Znzy+561GZpa0sJBKiaMIyMHyN1ErZ9R5Dd9K2n+NUwSC8YHmdYnu9BNV2qsFv2
xsZy4q5QwvPn+9RcfvAQEtOloyVUvP674nAAQPfiVkkEU0VspJffKCkiMN1qwv8psybZXFslgetN
r16phzVwBX+yF/NNiHs2dtzgFEcAEeBy/aE4klEX276uyS2zrUTI109/cWMZ51tdTjscXVsVfG5b
BsTryA+Don/piZYEsR7AAbq+OHzqISrOz3YGf9P3xIbsSzvozLiIN/69cCaww/NTxRtg+fo4XHlX
DeVoMP38+alXb+8ni0j9wobIwTnqNGztiGVGxAC9a5oZH22YBjGSQB/m5G21f4cvW4ljnpMTXk7J
o29Y4W4rmYr5iaTA4tJ6GW11awmtcqYqK+JT9aejmNKc1sljA1PD/BeGaIRCjhljAY8YIqUFdZXS
msN6LOuelIytQz/oVL87aUzOJbO5/nKoRTTix24MAinlb76HXRHI2+fYpfGCER5rk1dMe+298M3f
1EpP+QOVT4/3udR6rW8gel32fzKQ3J9LfJlxd+wTQoXwFeh4ukA+ezZXhCtlASLxK9iTcK8dbmda
yjSHMqiV8dbjvncptOmFtBssKFzFvrYA5LPcHpgogziy67SKp9nXdMODXTJiLCto24N0MbI3wSNQ
HkcDkw5hEhEnyC+rYUlOklf9D0PrHkfX4iN0843vxp+EEuXgGf6DgQYT8GaAAn2l4Qpqzld8kXO+
6kxIhavXK7/WtmgLnsp7gDHC/z0AxLO7jxS7XWHL+Ezkj93wcqM6ZJaehgxqB+0PNPItt/kRqtyd
4iP8wxqdLOT7GIJz5isl5PdJBoJmhNmbcSvoPhf8cEDxlZ86FlsCIoVFsTaeyYUJJShTvpj6fTtF
E4AvkQtKVW80ALcjT/t545Jo4lFOrmNPs3DHHBc0Y787S7HMvN48HR5AUWrU/suXltlOvWwitJog
istUDf2ta4nLqLhfRirNxNB3mWXecg2otek11dS7r1IKX+OPwD7EQLYrqU8cwWKbddttNR5e0pL5
rUa5DAitWfYUksVjPd23D20AAYysmLNgtAVdc4qrdR9qfAyJVkszYxTvwRppDU+xAQn02aKQeMeF
GHmHCXW+vyOk8pHUUA0c3dV37dpmdOfkJFZYdItPiUIisCiAS4MRYRM84rNObgIrL6R+zxIju/Y+
iLlNk6SgVLQiNShWHoc2Qcgor3WLrhS9KEDGCmyvatSiMUUeCkG93TMlhIiaylIZr+bb/JCYZtdq
KKx+3DphaEw9RKbPnRL98lci3qljm5u4MMPBLO9exlHyVVrZIsWAC3TERq1IH0cdBM2/YNfDLevW
QUvQ8W6Y6S71YHoSNhwQYUxCkUsBhpvRI4bf6lYDgPrGM79kwYRoXU9QP6dMpjsR5ZeFfap1zZ4A
WVnXfyH5WIjNg0KaBpOfFkNH5kEugkGq+UytCxMlnorUUHiVa5HHAyJKMXVmRF6MeXXbgJDRG9h1
6JJ6fBZ9RWx7KLhYCjOLjWxFfWv+aVpX/e8vfO5CX2P7tK82gwklkOXFztyMES4C87h5L7aS7+Fd
PUaT9kLJ3lD1VnvqQUm6Sbf1h2CjiwegnntTvRO1dxO0iTY7uSJkHA2ZRryPIMp4NITRSr5wY30t
3f0an5Lp1iY8RCc5OvkBza3bvXh1VUjuPskPkEYXoywLbfSuFswPbkx1f4gI81MBQP7za7oMJwis
IIYkh9PwS1LhJ638UyllotOKK9fX04a62U373UpeE55aUt/Hj2YzZAcTnsUqieMkeTdFnW0UeoB3
262c8FC2wj+1xFBe3OxnLECkNXXtjCs30TrUfTYDHTr6UohvIXR0YRfg/mviwG5+pZ+9WZbQwltx
m33APqUTI5FZoUJhoLGlNLbMHaZcKTsqQPVG3TLQKwXZcw3SgyYQxZQSbTbjbyhLB/rMLiWBh9ch
vZa3LEgBKACsdSKxtP4fOVvMxJ/U9mbd7aiaEOy4nT73xsDnaI6Wvktslbs5dQ8GwFGsyHShQaNQ
KmM3orRf2kML+DfR53AtA8muU6F2WzF2GO1OXoPv3dCmXgR8OoWIti8QunQAm+LZ8PRWCnxH0ZHD
ZaqniHKK2MkH+0SK5uoSIYTib+uIoYy9lyo/bgtX+CT45oTu0BT9m6u/cg23WBE1uM6YUv8Hx1lx
4EbhY3m6a2dof9Ck4U8F0GQIUmjUbxAZuouVz9TvqsEUF79HTa14VIW8CUiApzskEKmXvexCGMYw
ZvJHiA41V800CJawr5Bqpt1vUImd67/UYAzmGHx/58GZ6i9ienHHq3AJ3MQWjCXZVL2Uyx3E8IYR
+nX2Rkr2GO90yJP8XHtdNgAKQmvINJFlN7mq+CDApY3xrsXpI9wOTe2pXeT3mXYt96z1oh3nRazw
ZGGNJHTHduNEvaaqkOJlVWN4A/jSRhw4QMi3qC6P8sKuWIuzAO0sH+xVV6mvbbBKtzgYjFt6S84y
zi0KFxXe99wy2YosI4raoS2FryswlEa7PJtdcEqyYsjQcpuOS0CXCttnvgbeoRLWC8h0eOc70ADp
rOr7Rl1O4Lt+xPw6eS8AqmIUGefR78G3BC2zr0o5ey1fN3ZQAj3q4aja41/V5FTwMNHy6PS8WYC+
N7/3vhxoOP+68/oh0lIxZIHOY+E1hEeO+teai8jk0aboxgiNW6pl6lIoP7hM8sD4+15/ijKtEy2z
8Fu8pCmqRIHz9+LxObzVTO0CiTeleXRButVFecPo3vHArrblX/w9FoJLl1nOqR34wvxLYN5OYpr/
LWbZV1bdIIHDoHN2muD9bU63I0UyAPeNIUKY7w7durCqFWwEhj8zHkbvTKMKUrPMTCUS7fyCMJ+o
1j0iNfcqrhklK99bN0CtuqyL0L+PgvDLgEiW39LHQfVK37VHyx3i76Hp+vXm+/qlPiVxFR9s39pK
2wvqRdNV8oxmhWhYKKpn41zh71ol9sLHoF91TYqQYtrgsdxVGMR42JrDch9K6GNudt1oh3A2+d5l
q2zI40MdQakUgJrr9Mz6iw8N+zrBXUKDtiEyihYvZFNFpxOTJW9gzhedW5/ijGy38aiWzQMsVyxj
Tmlcl9Vt/9AYtgkTT/w+PqSvKuixj7fHS0IONzYlp/ouJLE4/l+JmAutiOwOQpPFNzWwmO4T2Ii/
yHEGDMAklyRCv9L+mkHzp6UzfVoTfSt62fGpNn97ukCxdgLBW3DpEeCfLRlgF0NLNFYefXst+MIu
LvqlUC8qpLqNM5HE++WjBAI8XiaYpzhwtWPk5SUZK5dTepvgN2MflCm7RxS6GJH5fqtNlCwWZbsN
BTfQ3TOmQcXw9ws/n8C66Wp0uQFxTR4wrTPEsVbV+qFHUO6BYlWwhxM85IQVv3yqECTWkiJuioZ0
3ttuIuIuoL1MhAFiN2RFH3xAf0YRNVZixftDtyyXrKB2PvCCXBQaKPPHgYMCZh5QY6ydAfl9tC8o
oBBV3tpvUMMS5FHjliqpju3U0cyAe8zxPrWf0WiOKsEe3aWjpBU0Wv1mVNxob+RpvLrJEImXceN7
mL9L2fMAofl5v6Qw5H/kSTij4BBFG4m3X/KAZjthCXP9R1klcVk+cdyR4vTwlVD/BO2zmORCJmOR
IoixavRQBktAwLjP8xnSRJ9rwEJZH1j8NAyeCaqa4MoK+IVyhBag9LMmlmNJBg6BXR3UEdwyo7kB
Hbz9OnV/E+FVpTwSXzUrzn8k0UyfcxU/4JyBlQQbDxgWDBIY7/Lc9vp8+eG9uW4UQ/9YlQBGmWse
KwlgYYcBwnLAYfYH1qBBugFSacIGps7QBwxss8J/h2gZ2CkZdzo9OmSPEmJsCKMUOccMrU3Sezpv
vnmKf01bE1Izw4Ni4Agh3TsgbT7hR0OXuZJHL+K/rhRSSvIY2oSHQpRtbrvgYkrIdAwKE0LjR0KB
O3oOpzu2mc/ztX3UtbQ4r0datz/R67xWrWTZoBrzS9fxBzACnjGRC6+njmiQ8Yng48AKA5H6mYlf
2WcIJjeMAT79ZSi26j72Jj6ZyFljWodviB7PhaWhsVhapBUdjY1/g3I9OJ2QaTWYblRxhFkDHx+S
BhYO9yryVpzk4l069YEurrSOZCI8GpwfCDGsur/LixWj8jvTRvRTdBsRekhRM6/EkU2q9n6EV3z/
XF71gUDFBcwMYwAhqf+sxBt+2yIr5j3p3xYpRHH2uYutmyFbzjQ6co3XBat1b1Obwjd6IDlzJB5A
XFMgP0e3FzY2fKn7IPYO5Jkh4tcxp7I/ZR0hZavhl+I2PCCNZItRDVRyXF+dv2JLAUCo17jRj45S
nYwiLTSSNnNmT6uZpYUuGbc3GAflSNZFRAhke+9qMe6saBV9O1ZkvYM4x245nNkYM/Cm0E6xPz+g
O/xzQsTY9XlLjrjMa3vUVB5jxFfzuEnAw4Laez3l/e/+zE0EOFAHjZF2SdTmKwVomkK7ZUrHn8KP
rS9zzEJiKoZUtHJ1jCo+sEeotaMcwslRjuWHYa1pZ0pbEO4GsDgrzlVOfEwUYQAGfgrry93VLAMb
TSheV+mROA7nzEytL71aNwbHdIdU8L2FfIt5VjIf+1JLXhxH30hBjZESE6qOhizwHO703XxCxYsf
fQcF9thbuPLUUKb1cb3HXKU65YT0YWNRQNye7xvekbTL94UHexR1rHnnBiTdq/xAxWWKPXBe+j1b
5ZjD0MsZexpKbt4WOWRTTcvtvn+iBLX/j1AuZ94ID/y2m+JM4TeXxu5JGLpr6QLyfy6Vdp/Ia1tk
xVW7B2c7yuQX5Z7Eenu99GcLiHAjEaSBKAMVJEfL1tpEyv+cJhuwnBDtvlae4aIcNhgjRBqrovh0
OleiqmP2izShsONUgbgdo0aNz7gfCQTmE0u2mttJFqGxUPFsurg5XsdSHW0uUvrt+mNxELkfjWzQ
r1HecTtGkkR+zGBfuqH/j4XVIRW4z0TWg98BCjtUwiHNwFG080c6fXMrT5X+XQ5ND+k+p8JfaR0K
oNAD31Fvkt5qcm0Hx7/7ccnIOIyVQEiKUBIGgIwEZGi8ZFn8ubHA8/nVdYOeA7jCa8ggK8SwJJMp
U/1RCtjaIWEyYIRbYxaw9mnNdPbTXUMK8fnmN0o3pwLMKj3p9haB5wj6FEl4iWCbd4QKNB2hukS7
sUptlYB/Vjo0VCeGW5r1Tr6nno7t/vD5OgD26rWFmdrWCZzpFPfnuUtJY8ecwrB3g59kWYlnZOU7
0fy5yTMfrWez4fpokeHaQyWqqvFwWEIXyW6J7Slp6Yb9A4gdrb5kzQ7AVkY/m3ITjAA//VF+KZbv
QlscO+bMo9hgOgV8ZJi3KSXNlFjH/+TDGmJFof6a7Lg5ZFYgbDrYPC7Ihwd8/iozyrBk/Ssn1Zq8
LJzbAxuh8EmRIQOkQv5bpvwo/i7zeWjsVSflFjvXSA/OII6YbgdCqwkfwsu8AGDcjGXfY4Qn2BXZ
+7wiwQ/2CocAibuh3MtNmaee9GOTHpjJQkDc5VJtLtAPRTD3XZBY3J//POPRHNuEc9T9ps3Mq1zv
+MWOBkCIev66pQiMYuvMVySzbFZciwDpFAOFWVm41NJU+lRhjQ7i0zFZL1F5sZEinmHswd5IadD9
gqi072RkgVNISbXR5fYYKpdpNrmRPZvDYBD046BwsWwOcDuSSSbWpqQh3gGK8wDnOA5ANZy4j2kN
yrAVykXUtDgMFoGULvGJyBbIMY3Wphjk+Ksg7G7zMLLmaE1A5E/HISlKh5zlN4sw6J9bdFocNFRy
5NMdWOhFXKa5Orr8EI9C2wuJ5q59vMWye3il3pNoY3OxUD1yKlwfPTEpkkjvXFl4lJK7D1VM0bH1
La9PfOBpF18+iBQo8Ct6SPQchtz+NUj3txX5ZFb/jLYMgvBptluDoF7zF3xayYHUr2WLYXznDWvh
FLRSjvDc2pjrmeLypv1xYIlQF6o+HQleIewWK0A9yKDpAzlpQbDoR93Z4gBeP3DZPmQm51hVmA6h
Q+NZszNoWUTqAQjdRBQVTMOn7ada2Cn5/oSB8gdRLu3zsuXZSGvJqYqHUfLD6hg0vep9eo79dEdy
avlpyN/PjSzbUzQeld/1sgoclYw5OsO3dbRs40OYRPiMGMCsYi0pq7qOF1r0Bphyi709Psle6Fcq
WeZ4HZVPzWfoQZRTEr8VthlFnpu2br+d4Xbyhttk51csJBuzM6ihOnmIi3zoqBy7umPdseNYrQjL
iis6rzz+dzfTobogiRVxjlzMwIho+Thb3zMgGqWGeqx/Ad52HR0dd0slmbIHAWdkLm263Yra92vO
V9Ks5vHZwF9SdCA0unYeOj2gkbKXEm7jAU7u8fuygjiP7tfBm7E8Rqff6pfQrqvw/rIYwdmcLW2X
50PQIzsdHxan+h0lTDBsB5OJ7jjbWpP8A9HtM9ojvSs4fQs2BtjWfaNSUr4BRmHtCWGCVa2WYDPA
oHSHu+iuZrWT4qDCo/Y2pDJX+fxQhkC9te+z6d01v9wQ0hxy50PtltxYeAnBLcj9SLOSwthyhEuI
d8qbBml62NuCVxCQNlXprk5XjqMLjRnsuXVJrh3hwrAM01jcm1LJssweuLEAmvi8ZpGfGaQVCz5k
Whhn3kTSs+4ygvXRlLOO+3bx95aYCfpnGQLHshNOAtEG3bYzzVw3gA1wwpS4MjoBgQm1xoeYnd0w
+1TB3VXtZTSbauTQzfnjwAvEX5l4EDW5aKdz9s+40bh+2Odgst1SX04hnyGSLgoKXqM5jBW5wRzW
XSUrIjuIG3Kc3AnS8GWUORYxu3q4GDLEJpp7d4C0i45yQDGUjlmtRsKVKR9cFlL8lb/NbaYZRNvl
vlB/Rd1GT+O+mB7vac39FG3NNfyNwmoha+M/tUs70KlvShzXBVQY/+/zLh9mL+ZQzVNQwBGvAp/t
vOFKAE2yJ2Rk/X71eF2s4CJ6jVtGKhm/plMu6kbvygAEgAQUIaf/LbYnsaE2xcfe6hhqnFVLGFq2
il5d+5lrHRLN/Bm/We5cqtC8gKLwlZ7q5yK3fLYWgUI/l4DGd0lKeg17BlLyFI1rNMwOOKxqUH9b
+2zELkv5ms/uguvTHTarOK1xDLIHYU5ZqX51ZOVJysFm6zEcjmZxiofROZJjM1LxLBPxbtHH659p
`protect end_protected
