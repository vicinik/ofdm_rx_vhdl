��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_do�q��+�����T3M���ZC����	!�*]'_��0L��A�vT9����<Hov����Xj>[�=���u�s���!�Y�}>�i�	7�&��jْz!-����}f��*<-$F����I|�hQq&A��&��D��1u�wUM6:'��g��ڊ��fC��D��K6��� fvv.����7w�nE*�b����l��]�gI���)�nԌL�
ʚ�Gː�.�!)��#Ͽ$#�2�8��$e?%���g�i������o�#�����z�Bl}46Z Ad)I̺]�_�\�W��_��{;"��B�`��g}jߜH<��kJ��*�.�O�
<_��Ět����8��{B�6A�����gPP�� 5�v'�2Wek̅ak������d9%��`w,n�)W��D�2'G�uǂ�h���%���\������7AH�"��XͿk�f U�ss�٬��{\�g�����/�xI�7�W�'�����rC�BZ+�"�랟O�RW�vhNJ�#�A�j�ݨ��_m4JU٢��F]#A��8g��4�������Et�
 A�|�tC���W�s *����)���CS�
p!��c�p_z�x���r� �nc7ϬTf�@%N�������,���q^B�p���Ih�]S?�.ʁ��q�1�K���� 2�M^��_ǵ��%ƯE�m_�GrhX�Z�ƍ�6�V��yC4nk���ʜ��>Jً��9e+�����C�/x-�sUm=j�ʔ��q�~�B��&�&�G�S�(7Rl�ZTĦo�%ij;�*�1  �F

����%�Gw�!9N2󳫷_��<�rv��VBS��&�s��}��
�c�9�����=���B>�@=(!��K����]�� \��`{��Y�Ys�k���\G
��3w����-'����F�4��CS��$�;*]��x-�J�8��W�y�.��>ک9��o�;$�g�����}�� V���t/�����K���X�����Ѽ?��� ���Sl^Z��-AnbT���]4	*t �JjP>�<��"I<2_>�G��f��$I����C0vsg��B;�PH&�J#\Vj�t�(�A#miX�m8j��>���kh�)@Ք,�3'�Ut!I���+�UZȢ���c��??^mX�':Y�V��4�; �X,iu"Ώ^� ��2�ڷc;���Վ�}^@P]��0����F�8��N�\��Y>c�M�T�ۜJۯR���{Yx=��R�C�D�*�i&�/[[�E[g$�:)'�@@ʫ�m��eĳ�d�ҡA�ЊVQ$��
-6��e��0i('�]Fd@��O�f��sP��1h�Y� TF�ǭ1�' �T��R�Y��W/1����M��R�{���O�s��&Q�MIm4��F�	kt�
�}�F�\�H�����n��ő�3�U ���6��n�l�X���-��	��N]�����c��+h��	�~�+��%�<�&��K�n;#_][�,�����2�b�6{����4�*�^����n��̖+�I�R�����W�KO�Z2�+��i��>y���r���[��(�	Y����!��ڡw{�$_�S`��%)+`yEx.���Ѻ�&^N-ZGƯ�&��?&��O���!�ᢷ�u�ρ��f�Ĭ�v����Ed�i
�k���R��C�OB��T���õ-���)xz��(���ĥ�|	Y��|v����b���A>Z�zu�QJ��2�w<�X\�����v&�h	L��F�^��H�>��/�^K��ÑA8�C*����t�%�τ>�R�,0aޙ�X3*��%�U��g�h/k�'ӬD��\���>{���2gG8�7����),�'?+w29!l���-F����o���l0kݢy�jX�lѵ���#����|�$ɘsH���q�c �e3�����Կ�����)`d�+��>]��ku�~'+�o$�[t���D��J:���x��L��;�҄T�(t���[�&p���Ծ#oD,j?6(^��Oy��i=��J�}��O�؊.�?����V]^���2��x�Q���q�~H�I�$�2К;p ��DM��O$ړ*.z�o&F�O��~!�'Sa�\��t��0f�=��k��cR����4���%ݵX���4�|g������!E�?WI���[�%�ib��
?�z��`��^/��Y�Rf����$j4�AF��Dj���M���	V�hvRK6Ԃ㾛���y;_�N�/N
�bh�����|#�	�����o"f�Wf���B�	d������6�D1��Y��J<���o	`n\B��#F��s9�P'a�}�#�9��'p��X�6��iJp�5�� V��oZ񕱄��d=����շ`�t��,�������'��������!E���+��I��O+�6�C��'",��ҊB-�����U��� e�w�%]�6�����e"�r6 Ȱ�����4\A���ÜX�߻u����+i{��w����C%8��A�.�U�<���R��J��<��U��vfnZ�g��8��[�ދa��J��( ��Y���dT�OC~`k���W�D�3������%���hc��=������Ң�`0�X������
!LU�P�����,�1R��_ԮBhAᏄ�}V��m��.��]q1�u�'F���쩔��t
XUD���'*�.i�̍�7旍~5�r��1�J�xvj�⋴)2v�ܵ�8�G	���������Ah���=�uo	��9MKkQ��p���L%��.E�JS*��ɞ[7?��_T^�Î��*b�� v�>N�Ph�a�%M�m�(,�߁	ߘ�Z���m&1UDo��X����N��H��럛AhGR
�/��@�hb�0�����kg!�L^�0j�S0���'�ԍ�Ӧ����5~���ݱ�a�(+�z6��=V�4��M�g��5g�9�N�EE%Ьe��!b��Mg1�4����V�,����2��!i�$�����@t�D4TV�&�A<��5�l.�ryJ�N�=����M�&����"/�>���>3rw-"�񱃌hJP�yV][aE��E2�x���&���.��<���k�Ǳ��4�s��|���7��t&T>���u�.)H[�����q���e�Bu~��� �RLs��o���5Z�a~L�h`����<n��GlV�����^�u�BR-�<�uT����Te*��T������"	fi�,3m��K���D
�G4�V��e���
��O1�B?9�|)�;Ǽh ������-�@�ů"�1}:�/<�x{��n� A��	��������Z,,
�1��<���ii�P�L�����慍��g��;@T��U���b�l~xNO�r��2P�`�]�ʦ[v!��E:q�0���ɥ�*�֪Ʈ^
�	ܺ&??]�4nN�].���6�vI稁��v�y�5xT	.�l<���"��부:"�f�Γ���0jC����2�'���<��1 ���O�j�}c�D\�����c�S��.5�S�e)���,�1��m�M���Z�W���r˹l�@g�`黰#��Z4�%	n���o����&yv�^�LD����=�o�л!���?FE����1�#6�KL�ۘt��O�Ws�#�����&�������+�V(y4����*���#�hj�UȽ{���/T�p�����p��_�O��P�i�&�-��y�Kе�'P���SJy��g��o�-�.Y./?~����W�N�!�&�-�8��JHn�Eu��qIw�o�� u���␫jŦ5���*t�ҳ��B������}��ohQf$��lL��g��.z>��qS��Ksr�q��V�	"f�����R#��/��:������mr�L'�R)����e�����l�b
K��ɴ��\�OE��p���g���U�����E��4dUP�H���𑢷��_!q4K�~�	�n>�Y\
-Ӌ"��@�L;��8��R��KSX'��y�氢��!>��� 9�l��}���tKel�F�����t��|c,Q[��/�W����nՒ�m������s*r�G�~�ɌX��:z؁�fG+FB.��曘=�S7Ja�+�����ppT|���2�6G����lbD/�