-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sbCKXIeHV1yZWsDTuvUQ/F7KJyG5p3gjNVlbOhdVpgONWU6UphAggnKHm5WfE9e5MKwdSaK4fkSE
n+OYhqNXCqiE6xsoyL5xnWA19atG+yGaUBQmp9DQ0Frl7uUBCAFo5jbtafhxs/2Bh9FJ/TsJydPK
FMWJzqyloETTgXdW10WHNlIOrRvmH+gaxxSoEa71mSYt+6xlc6rtjCDouEMSV2JwAkYLFiVfejS+
101ibVHyYhGj9ESs+2+6w2sQLQalmQw5Iujj7wj7B57MQAZ57hD2oTG6WEF/+MYmrUB5drgaEnI7
BdbAk/jcwgLJe2taM9XarFHozs51TdTc6gqzoQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 50592)
`protect data_block
EHgU1XVK0hzIE5UfJbGZP/D+M0zLDlVwxRVsYLgIZg3Ca1Av668HlewWpVG2EBGnCDuE2+jxu+cU
LGds/SbibmVnxvWq34zjoR6HRoQk9b5L9KGmIU3Vj1hFfF8QaVT5kaWtyP0FkatfEDY4hTIYB0mU
NUuSuZnQHTCUTNEVVhVYUndDhRNLnknFubN7NCgb0tX2ZoG4cn2QxEwmIVe715CD9zMLzLO3vfXU
8f3wurSUVsKQYp8AK6pSXHxfNC0wC1onGzQKIz4/mOl8OfOAKBuMEvTr1efSyx2gWdgk1YE7FolK
Z7t6GiyIbNtbtSFivs6ADSwT7CX5WR2Xf/gOrfLGxlTYpnQBNFs57FRvIT/PXb1dYl8ME8vgz0ko
/QS4B515/opWigSoKd49A5TpbP9n+7B3mYinrjGSqpkeBwyz7HDSVUxOhz+5kX+3SQMdi7WIbNTE
sNkO2cpxFTYFaEXLcgZu+U2aLzo0aHOiWARRyxzyIXBO8JzR7iafDNoq3BDZAOVnsYSW5dKJFbk2
DbdSzGtWPcNlGMAiqzwgbbAcsLY88W01ursmnS5+wdtVswqvH9oZPOtrb8duL6m2leiAg+A3yVuS
V58WN1USIL5Ss7ZdqzmRmgr+WtUEkRpuKVjcGWEAIkS/IgX6/ZfkKKSqTVbUIEzT9meE8z7eT0uR
mIJJUv5B/h26uZyc9oxf9gXha76xZJbzIHy/Hg9RcqoC6zUEXU955j0KWw3+4mCKdPvDCgNVW/Hk
p5IbD24aZAGFrB9ltfeNPwlufpOe2+v04hhXuKzK2cLZe/BebPTOD/AgDGb1TQXjzqptQbhCEkcx
e5RANXEvY0Ij1HRDVZYMKjOOBLMnTPJlm7+GfwfUx6W9r7qlAGCJK3ZINxEHnWl2bHY7K1XK+J9k
t5Ts0oX84xrTwbc/6FSxJKIp75GVAI9i0ps+jw4m+A6HPi42pyxYlYb8+otMIqvn8iiKwAO+jlkT
1cjUme47wxwMAtVa28TVwI/1W7+xrvB3CczaEpiBf5jFbypRDRGCCRNj0OG6tjzDa+M2qPIi63Zs
97uehMi0MVOwRp2WILIDnvSFM4MZAANE9/iEjRIzTq6Gc/+TZUSkonAG76Pip/p7yAMcL+EyCg/F
WbCJQDJk9gYPM8qzel9kUkeXnT8Rtlq6V3K3PUXhgzelNb2Lpp6cDJH5U5z8gf98EIdM2T2DoImY
6w/Prh/8Q6AjyBT0hqBtvAa0x6Xu6InIf0i9Gy3ycdAXrJHSscmSazf2sa6cISZA8osyS7mT0KSt
nCyGFpwGTj8y1+hwSxndSFi+ydhokvqOrCIucMUL9E4qbzKyqFNTgUrd1oo45S/cZKTAuyyZjDlZ
Ss2FIEx9Sv2tAxQQjDpn4CYH0VDzhD59aGrycAdz0nciSi7EuEjWVXhbFBMmtefWYy96VizYccS4
GIjGD3N5EiNtANH2xhUsxk4y+V4isFYCIip81OaAIll5Z9Pjhj4QShn7p5FmmtS76SXnfL8lg0xk
6clpcmz7nFDhMNZJ0M/UqskjmChjbT3iVJ36G/MpZUoYzI9disruk9OIY5TQO0qaHCSuO2CIOYeH
5E/iH0C85GFYUHVjB9OG+/0uVKIThEN5Cz7BMehh0PCe/2NzhzaZtRPVdCFLxY+DxrOWlCNj31h4
mBE+WWmpsRRXTDkOjhvMOQev3c7gIZiTAyXh+Wr5Fs3VqYOu8uP+gQDm4oRS1hm2mUoukD6JxRbn
CUtyb6KB9b3kGxYsvfZLun2eNa6oby6TJucozb+xka7wJqU27jZsyMggIv7V0y2GPJzfvAP512IK
Ko5zMGdyxcp6YJpoGg0Akn2wQkffYd1sRrxi4yJHPQ4AR38mnvr/VkvLGsipWhL3sTy3GXqv9Ggx
uBPjSTVcMfa4zMl3AUENJOa1ddTdjIGdVrFc3NEfT88kpWqViwzeZfWOHJ4XR0X0UZOKU5JQoHa8
D5GKFw7vsgj+scgMCWWsmCzPniiquN4ei0EA/tCjJqlkweFjB+cEF7DY6vjvNPBeW3anmBLxSjzR
QCqV8UVxxWCcct2OjO8rKA7wwNkvoB7ZAqcMUOKVfOX1xpt3tPAqowNxAHSd3Qov9ihT2ujRO3hV
d+Hfp1BLPuf6Pxww6RXYto0OZEYo4E1rXZYly9RhxDFvDPOhcjzEI6mR60FbOwsQVlL+ElJLpWvb
XF4a97ZzonS4bS9bS74NXObwUsNH25XZYpctwuFBVk9UgnYb+6arnHy/MQYy06RTPbtjsHZGu9I0
NIBEuxqjjLyTd2/WqzV5IUv4XkyRPJ3It8q7PDRGsfKLzk5SLWAfShktJ1hcuyO38nC+CmLB6TqC
23Nqs56izBIxoNfZt1RIiDP/UaF6ZEUU/UKDXUCubbkXKg8nYInRP6XTpWWFw0lg2+fV+TLGPkyi
Q3beSRCWJou6OeMPI5Ly8meCeYxtaQayffFYpE9fHjAKIWJC+BO1gfLYSeJw6nhLKJZUx9TuoOuq
OHwUEx0H1ALvUrWf9obsUAX9fcB/1dmWBd/qLLGS+QaXEkzOgHKeHkmUb5KZsBBRXBsH4Jyp7nmg
3SpXb/FbvhpK6J/wyZSICnd/YZf0ZoOzLpjY4ODfsEUAfERsb6zg6/f42YPwQWzKkCL/qAC9mzh1
0S99Un8DTji/TKX0IoGAhMNERIe4N4lDajfs9hxqntl7NejYfMI1Y5YGBnJcWHbKvGv850Jd/SlV
edyAqfFNS+bdx3abZXhgecQ8z9TDqql53U100+2TTIJTnILeqZh0lVO351OeVn69zbUquS4Mcji3
ppZ+t0y94DjZ9W/IuA0tuvSD5Hekk++mTX1FY5vbJ8gATxjBfjRviRP8diIiW6XCxZWAFnnpvH0a
c36sfw3LwC/XjLbrY0k01f4eToinFyLv4a6jzh6sUZQ8DwBG8ZZgJLfH/MtrSsMVZWtePo9xDmex
fDgiMXd7vP/1TJTS5rnhxIAhx/UM/AzwqzFcuPNyDdCDq8x1o208Y8cQUIv5xnsD7+pNTX/G8hjc
CwJlhSLmDgW4FPo2fEgt2saWJBpc1dmM4ZuesxoYIfncYYaIxWU/ivpG1DPIhvuHlwlXMstJA6Ju
c5djtfXq9hKrXlBEXgkVNtIN1VI89m048PZwxzxNWTUrnEX/xW9K7HsuJH0yPl8Q3RkVpfRzsvw5
IXTfWcJ2NYpaUEfN8/I9kDc/S4TiboeMKkgOu1V8BU4MI+yKvlJ+cmmn/HHKgTO9j6liqySnhASx
Xv0IYWKlHGTvBLjyrp8ABzAE8bXnkTNIxyNqwzIsaT+CU1U2IA14OiqbC9KeRQITVMsThNUeKAhO
0G4tAYgZow6kaJ70ryn9DoEQuoLm0Sw07PVTH6HHQyFQzMiMM3ouY25rRnTN8z2fCeXu+rYNpOtF
k/H4x7k6IsGEcVsF2B7pTInuD0iNbwOnTBKa6IWn+dsBGUmAPVUxjuKEJaToZLU/7yBDymKsT4zi
8BaucrQaaWMvYcy0SilNxAiAWp/hJbuUOkCu+Mfkfd9qXn5pbgjJ1C51+G7OZr52jONrtbgIiHec
EjJcS5MoOCOzSx1XTHjd9SGFGliFoSsY5x4kEBHAvoJ4fJUVbKcPtncV9B2vjMnRIJCrcRLY8ZZd
8T/DT5+qIBp2Csyh4PZ1JTROEcA7w7nfdA4W+75R6hdjO8ZqsLcdH1cuUog2H/Sqzut88q9+r2jy
lfdzCammDD9b6ReBEsj60bD0zerFAFM9snC4jCUBShr2omzK36rlTd/BhNAMxTdOiGKIDze2PP1o
1XFwDvB7jpVqIWkyV9DtfzqBLwAXvjcqTGdeKFuhXMxYAt+UsUgFjKLdgQCFwPILy1VzxH9TE809
cqzivSdexyt0mOgEUtxjf0v0m9EierPzuDUH4j2yHS0f8WOONTk0qNWUsvMOiT4WD5ClfKvpzLGu
b0NJpZ8EGUIj/vQiTB591dgrbGQn0tK0CTTUkaWkYcymkWm/a2zEiuYdA5W6RxukTpRfjnRircqF
hGQKEMvGLfEMmd2TZoCyRDS1Sb0xOmhyoSATR4D2mNiORUooYqDyRj7aHUH6Any6YDgu+8vMxIBt
p/R37o4g8YBysJ5mTLPso3nTXM5S4Hp+5r30ViDcCYBHt8pg+OxW/KjGbBFRBxEGukW2a0IK7hOz
e2mBfPbi3Q62lUATZbudD+z+MS0eO+G8Cpn0mDugHJMHOEjMU6V6Of83IFepw3xYd/cluuxoAnM0
9Kh7tE+QzrmCoIKsuFhw/yKqRrn8G+JMH/aySQShLyS8b2P2RQqy4MgeX85+1IgCzZoDHkNSRVSh
CPR+6yXqMXjYGGje4lzkmXWybBXfW1nciRZ2yzcABpNNFo/ievQ/jkpjokgtOu0mTasIC+W6/vUd
IJZhXuyZJOChuk7TNfllLjxsCd/2aoHUoQnjNXI+F2uAy7d5pzAia3jbrKQYLDeeo5VbSLS9nNXa
0HEwXPyVqTiQgy+DPbbZtYdDK9x5wm6/ZSuRb12zvD4whoGKuXyOhWd/1wcr3PlK1F9zubESGXwX
YZnmcCBSLxKoYpiByf+zrZN3V7spJs/bjXIu9xDbJLzXD7KdbSwOaheuclkrTqvO4fqho5Inb/ik
QUdC+ihhIBvqpe3GPyxUnmo3vI9y/Y++BNqkv6GFY+v98n4nqCkWCJ8aoSoSZnntOcdVvMkEb7po
S0VISu2B7b5LZRmHOHMmWkSRGHZ+CqCpoV0x6Q7+oMTbXfMT26EhJKxcvAEliVlNf8wDnWMNaPKp
+Z5YFRZ0dWcigib2VTfOJXK9akNsMzQKLxM5yCPAoqjr2NCXkpxUdI5LwdPY+4VNG/oyXe9HWMcy
laQkleESiROXxYMZ6iifWD44/owQQO9X4qFsAItgDm3KX//5ZPDCClU2q6aI7mIkRfMBDB6pKx2t
C100/U/L6iDW4CeeOT/Df0bxJCD33Ntz+Puj6L7tGss7y+MgkDpW4oBgWLgXE8IJnwrRtnnkqY9M
YgzBeDvfr2xNskHdZ0jZErL+Zoj8KAnYjfi9YvhKyQSMZP2XmHFzK1kaaWwgK30lZYAXkyeatqXL
Y9FO8LSHOWAA0p/6OZiHz27XPkC1XmFVhEXiywokZM7gBDs+4nxGMb/QTj/VtALxnupPBXhU6Uez
46hgRQb5A6cyMEHDzRym+UAmiqXUKHyqIKJR7UwSZ3V77ML5BRPY/dOIphYbI2gpyOo1T40QtmQ2
6xqS9DvIKaytqjjjrsvHLTkVRw639Oe0rIbeIJBV6DOPBDn+19m0txH0dosiEs5EzQP684ETV0Px
VXml2PXrGOEsPu0kU1Hjnjs8fDv/wjIH5CZc9sqQMvFxoRPMPNGmMiiKX+Z3+yahj4GMXKo58g81
lOrlL/sdWzb5vUsh7ruZfGTYAOheIQfblVC8lT6tqSmvrQ93iMJ9CRnUetUlbYRdlR1lKVtVipeC
hwspocePLmowafimaQjWXgW1KgOlQZQx9wVbgTS4e2W0idVRhgsJHrm67WYLMNPIpI7l/Wwf0bpN
Th01N5UkA5IO+geo+LmPvGAa4uz/wbvPInFjmGXiO5DpH76MBGGF3AzuwS5XzVS0D8bWMKx7CcXd
xIhPmvfGqArMa94bEjDVR/yqdQp9rvfP/Da9CSA01txZw8M7lTA+u1DRsj8HxfR6zqpABvTgovRG
8UrpyeCNVkpk4/pfmJWUSaMVSv8fyIZhy/EuERvY1ptzZHJIvhDRjMkoZRwCjCzUFyrIxdGz+vMq
zl4YZo38c5uvAQu1A10TWXMffmwUf8qZtXGp8DJ5u4VklOMVZhBMPnjrzxf1sk3QJ5ytX0y2jMKD
FtmkAOeLdC+oEhsssbZ5xEew7uFT5YnaUwuGNgeXyBDmiAQnqlHXcz+T3LJxN2/jKt37kWCrw92o
CuUY4b/OIzIasBCQ6lrXPVsmemem9dYm+mb1uGZsCWUc/set9zdN2QcK3FaxUr69TDRUi8ZNLUvD
YeBVN/WVuDA75Q7pQ10WuUydwC0e4RZRt1U+w7sevcaNku64Qxk+tCvbmN8oOz7NSdnM8Z3vbVzL
V8nhseNqPzLvBh3jDNciU20ImtbS22eZuO8EGph+zQi3txm0jE+PRQYAs+uOpvF+OFP8JwwzHZ9B
egrSTx24FyigOkCFGbox7nZz+USGacgeQKBH7qun0hbubo0jcrbnDBbsDTZaQYdDpN10DUXhlsZE
IBzw7zPU1aUGF51hMdnN6C9FZeqiUi3oEEaa064L4cKAOqz5Ba4OpPQMRjbuxoQ9wLTpyuBDO3Bv
tRMhn6f6xf1uD4pgs3ikQZKarKRV0xEg3l9472MRpBZEyR4CS7zCK0CSIVGOIMJEbSo8Arx5TKDv
Oq1aA0diUqvHgljmwwiteIEZ649WrDjyYPFb0thsKyFZBbZ+2goRZfikibz6N2eYE/yFhcUxEjPB
Qo/P+0H5J/RVUFtoNkEK2jJ5pXgSv5xutHv3nd4gG3w8TtvMfbdAs+0S+gdpkrNSej19QLpCRlfZ
DqJZwdkaA4lPqmIoYwFAWBwQGEf2P5jZQOgFBd/uVTuOFvDGJivJ1ANpoTQuo8LziJtROapYhFtD
msbnir4Rx26GbiRYnqyLD+JG/NlXGnSNSyvN02m7EyU2FA4OOHzebTCLDvvCMMiBt4P1q5uiangD
J7T4EqgmhPR4xE0eaup62rgsr4EmJtJEy19TKKJEsgwzd6kkV0mBip8UwMgoFmCYyHvHRTSeAtx5
sTabLOwdCa2tqSAd3r3QPBfRB8zknP6ouUYua2ZsQvuzGOMXbMmv8nN4biLUl5DH/udU7rQ7nJPp
Llm9bRz6WRT2WnMW55glr5/gycQA/q7A7aMzxv/zuIUsnj/0iuWL2D+jSEIp1yMFMAZXqEgvWBpz
zz/hBV5LcwTw3I568Vi6potXFNNQidFopYOEFU3n2HUQ3Ig6JjFaqqkDTpTV/YyVwI/utuwqAwaY
MQMKiFHyoAGxg7QQYRBa2hbuOUTcVxg+52sFC4pl1RrM3MIycvNw8zsFhRYS1FezlylBaSOnwCFA
mQEwm7VIv+CaTK/RLGm6kWUgm32y7kqhn3E0BWDRb4HjRBs8HaJGX2yHiwEi4Tub1d7DuzU3IhBI
HnUERTuOKjRk4iHP9OglWB5QZbcGMv03VgwzzUI6m+Fc/zT8mSdeaV+9CPLKA6NpW1xK5MX7WFSz
ggl5eYvczO0S1+awZvM4kWh+spyzyhUsD23qy0r8MoH3vifh0D2O9QqkQE/cVEshkdZ++UocA35v
rraShED0yHICg19vDFYKd7/M6x+3/Q3Oe+uNrgmx482cRAL5j1bs4WjYI80avGHCgm1oSfb+bxyQ
ZXlI1UAV4wAilAXFPNHeL42JjFdf/dvCNhjVDm6VbbQHwiHDOa4rw0nWzgfzpjNsndWK3vs50QjB
ZCf+gV3zK5pB+e6SqXrfjJlmU0/xroYQzxdQqdoCf7UgrUSk2cmzMMh3tgQWd9aKzYidXTHarpGQ
uT95EEXkVFkVP1jPfeR/QgCj9Aqz58oaOqyVGkfnRj/skJxSVSEBMmdf7Hr0n5O5W1hsTm8OmAwV
4MjzIFQyEwxi1yG+wTK+PNZxs5AA1ox66FTRKdEf7MUE4HY7VEVpEx8QUmy5L9ZT35DFSbQDA2wC
z00tdqLxIHcSvQI4ERy2wTx8bEFLkHEE5FY0Uolm+zpvwJvgR6HTyWmYpKdelqLMnLi5ML/Jf/nt
YtIxbgTbKBQqxyVwUknn7iGvCLXenfTZxnHuS8OetdarXyYpMFXT9SuB+jhfhj8pEdTnRH7VY6Ld
f59MImN0pw6l193cD4qNQ2IGIoFt+7BXdgO6pQypMy0T5mSYukMp5udJkpVi5+KpC91BEikVPDBL
7A5W26qXmp6ktG4K898yLrvmvFmluQRcvAXfEOjNDfl2uyFtaacNBspzVQVuos7ZWIMLSzuq8qdd
mFUKuz8sSCbwss4I6KK6EIm4VEw9E6G7LVoZ/q/WCucEi6mvIjEfuE200rrE0eAUKDzrDxaK1Sfe
ckMj7uRd2v46HSqcaEjV15yW3snXTNzIqAXv4mNGhMDcwEUp9JYkpdUTsq08smrLHUUBxL26jILj
aFf/aRMnCQRZBAzSBDF+cpQCSRbCKOqJqLwWNW8n0Z0HhEBx2r1+Ax2Fkpsjm9pmLMoZabbev5Ls
lX6zLAAgNwEeTrVtCjC0vuFRnW+uJ1/J6dPvmMzp+AUAMSCak6PxRGnYHsy7G/Bcz9ThnNyyzV+v
d61cXZO+YEQ5oOvpSg2C+bR9ipvXlEa13nSRE8z0bw0maurvS3lrntk5K3ZiAaknEwMjGCw7EDzN
E/k/IoLF5ZI0+ujzhaYvnDjZJEacErCWCkrpUUcy2z0aIsWOWJI5Wk8OLiaVuT7auhCZexRiAnmI
p8oliw/aF2BYePkCqbWzZfAR2OU/p0eUVImukEzUiA9jHYdzoRj8tD5Hby3ac9tSUtvhbjLepfBH
qEgtfdeNX1KCct1aDRopejumHC34FChP1fiAmRmPzH8oQj20Sipj/x3Ox3CWMuH4Z7J5+hvWwLb3
PeQUOrE/v/eTSf2I+AXplpCyPqVQVVKePwfCKUWi9wOjYQz6AknWC3lOiAUl+3OWtZAsFW9P3JsW
t69pFnMS5hlCi0HmC8UuJII2pGj4ocYvCMjogAKJSAfI+uHwcxNAjwMGbWYFYaFrHQ7PDSSfzhnC
C9ZXt8sIx1fYGotSXqKLgMKbrgR18Ey3WUgl8ADR2YXiWz1oPkxr6gCX/FI7bDbyLEv5DS1sXUxX
25i2o2LDhm0wA3tH/voOaj0J1We9tVJ8hT/7POMknR8Yutgw5P8C0S8KLWVI0eqgBwRSoDANed3n
0KDPWGsgdI5nrmWEiFTv5nNYrJvco80H6ku897lwAruCbMmyx+Y9BmS2U/dsffOij88jWG5wx2ds
4J0qSVRkg2HVEcSwXAnz3kvm3P8nMVjA0JqfIS0UvdwfjTXbysrx0IPESg/QfT50zhHdWGoLoJ2n
ShXhsZyQUo8MaJPpa4GZAI9rUxUGRKb/FAsOpPqcDMRlVw3QNRgfSXNJ12Ev59hGqbecxIgjdeSJ
ySjsxkQcyUSbx6g6OB5oVq+5I9N2h5tGqrNyAhTkdDdYzNnz2uOfMBe0yPPMi6yykZd2vhBWIf1T
oVC2TtrqiC9FZ9oFgsnMC59Ez2/FJfNz8iXzZE0TNz8nLpt/LZnrll/1Cjav4mUtBQq43FcIAZIV
0pOCQnrRQIo7TwxwJmBssTma5umRycyp8J83Pgts+yzpho1lF5YwXivpYgGP0HG4aqy/CVK+oPrL
pWdxp1LElPdV/nAzjFJXUjs6lR/zYPvLMTbATw71lLtB7YSRi1xIkWVtbjFyJWRxvlnB7xnzsiJi
t7MXtNmeo04TgOOhu+fADFE5/SARV82V5F1PYAKkY3iFl8lgLPiKsCAwyu40WJqraIapSUnyE6Zm
gL2QszGkX7adOwKWjcm934SbphMWr1q0f0FvqIkb8L9SANyBKfc7UBKX2GOWdVKuYRdOLbpmVh+O
NQ8lA6xLwnhzY5VDFkdRYSB/NRppAuUoFgSZ8ggI8sv24ZcJySvbC8uFrhIoOph9f9FV3FcxfddF
2j2z6CWk10XJgD2bDkF7hkOGSEDaiQe9JizUWV+6R1CCWbKTHTfCAq1+1ua6PF9F0j/wmDcU3cPC
/j/tSU1kxUsT5PDLJZ7oerPdcK2nT6fmmfLhJlWhpC+KWEGZrYt4v/tVDV71RLbDh3jcyXXx/e8N
c5CLYWU1324EDTnaufYmOndxS0xf6spK+nhBhlnpTi7mbuvdAZoKPAy2UgZpRL258+rSkGY/ka5d
YV+buHA8ntlIFU33kzO/Q2nmJwP94h/Ip53LTvUFYcY4Akk097kn3pF39qj/9MLANHpOFDryBQ+2
GhJjXIz1WBZsjCpaVx9BqZDHhnALOqv2nukeKdWLqRTRBJlKVcq/iSPCU9WCcgJvnIODEsY1QJWX
dLxqmDQNFeo14LdXJHx2KgTkJGYLH8bnCYhh6qB8t8W8Y2RMr7TOb2gU+Ttq9UNWaeogBPrd8QWg
Ym4FsyBCG8u1FLJI0ucwP+IFZVT0ZXBU0vOIQEkyqS0bHp0rK05KfZHKhoh9Gun5MgueP73uGYir
cfzE6HLjAarhzGC3Fxy3NLzQR93zP0Aai1zyAlTJs0NnwLoF+4UUO5GxJ0V5kr2f0zH01XdZblh6
SWY3WKkTDdD2Kvbv0mRQt/zCZlNmn01lohbvEsvNQnKhCQoyL5fh3sub/kO8N9I3+UbpGfjKGPs9
Ut/rLOxvYJ78ZcHsP8J0JE5WuDeQxRgnNJbjJ0UpTJvHSQRjRvqxWXK8K8myQE48a4Cp1b55SD6k
2jbRjvqReFfkzq7TjlRivAlB/KWGsFmenPwLlCmxe+loWugv2p76Vq/Ilbgm4r0BTLbF1Z/PesJU
XwOarlVAswErWBa5ObDkFBFLkBwP8QcoAYXoDfg1LEtraA4whyb+2co6FFYNv2CtMb2X8uj81yit
2z5lnGwmf3aOgMXGgAlF0VVcYLhOPlDjOiP8exuyG0DRzCi8PrBN/Cfx4U3wuCt+9dUb5e/s5W4C
sg2lhhXJsLmp+BT2vFrory6Su0Nm2+S5e3zN3kO5HAH8xcTsAFr6Xp6FvL2nXhCCimP+CD2MRsQR
aeNcfXQNm12c5knUj62DknqKhq3EhBxmtAV4qku+ETAEQk+0zz1/BEyjRYfwZZLWVGiCS6yqG+jN
OC8tkwk+Tb+PydofMftCR1P5v89MWs4kjm24Afak3e10zo0hyg5wM7p7KJ4KpYhaPke4LLqIPgn8
HNrHRTak0Vd5yRRZ41AL6gfQctJ/HnHt86B90j5SyuJtPeU11yflSsGfRsyiRfCcPHL9oySKyyZA
CBCXKH/guTkeh0UzjBIoNYKtSxPbd2mfoIA9iu/ZIgUE9xMmOvq+PNXKjWOJExsxsn1GVD+0Y8oU
0EUmvd5k6vlIR4SwiARRU6zv73vi157P1UKdum+Gn+d/nzOLYQ9e241GQbAP4sxD724/eoJOv/LQ
zwR15dbvlKtb1YD5ZKGNZTdopjpEbiWTB1sPm75IsOOiWP5GaUR+Ibt/lsOiGBV1m4o8xySroxih
r22mQq1Y1Bx1rHP1r+3902bJhS4+ksN1k6m9Z6N2obZSwKzmA8heYXHjS68g+AmMaXkRZdAMruOd
U7gDEVyTxXD3D81lRH15OH51iui9RCqRbEq+PxHqTxqnvz+UrrRye7AjXVJNR+lT7yV/ZzIw+n/p
XZNkIABgKKNe0uamxDoB4g5o6rFfj+bPA2WAKOSt7Aa3Qzor39S3q6Qt76byw0pTiM4YGKTUycmI
UbLD2Vx5+fBjePQYIHWXo1WS2DUehSgmwFxljcWOOrET31A4p5w8TGxsSr2TUWHvFpyf50t1+tAP
16Me5I/jFXhUKb4bmG/Q2aQ/J73vdOIwX3lyE3MDXBEtkwxfkMCZAEicoKXl4DeNEiAKAF+Xir6g
bOfZOaWbcnaYDxcNpYCH4sAnx37sm/n2bjJ8ZtB89L/CEwQOcBDcxaTZxNMTYJ32CM/k889dSpZN
Qvz9I7Gdq/9It7YuiJOSzzNkR8qSkLkqTYLYCvwAeYVrZOHyzH6vJdT7uciDXZO3sOV5FfM7BzT7
iFd9iAhwyeONXPhBNzNfCbRjPJpiVmBQzV5U5yU+S6TLgRZBsJmBkWAxbwP21WV01pY9gcpTW0fF
o8LwJO4tf9AqpOoG8Ip0ctAD25+kP3vbMmX5mZM87cDXiA6tt5JglusUcKSLAO580FTSQ8Z7oioT
WNrtVXG+AfV+at7J9B5g1XCCsLpDcXFFsREpVLwUnPMBKb51DjAxgUVIAR54jYW7lIrZY4OT0NMs
YghU+rRcI/Fz6KKR2opo33I1Bk4AWmqLe7EIvqN3Uap0tloyughY9lhNuxAQpus65DtRPNYxoSez
+so7gN0g6/S6HQSlqx/VxWByzpOv2OmH+/YTj6LU4GZtirzI0pWAxvynPdIy17XyJiT24qx77BWO
kEj+cvTZ5NMhZE0jZcRh8Lpf1UqS6GfK98XBs/5Lc/nzekL7WUfNanhQUt6txvYVQf0HiAm393c2
KqgBYUa4MrBjGwm84Q4hwkHeFBBJAU6KBRJOXZuZwPY9t5wiZ0EO/IPF970whhu9c1kwFDqcoY2b
TyJhICjF0FqgS0rvkei6bnJ7avsGfvNJtqr3zet2TTpFugKlm2fDVG0i3TpffJiSzjWpzpaDhOsM
8we0XHb5Pzozz5CrHAwWHJUGvFkeblii9tg4ogHssqa62MISPx69g6O6l9M52lB6upONM70Kcx+2
/RDvsvw9kmhgBsc2FU6VSV9jiLaJ2TJ2RwNNznHQ1LYx+FSC0j0Lj5h2QYzb2Nx635wxURrzJ4Zl
4dnUlRFoUrHuy8d03ZiwhI4ZIAtRWXvYOgrQUeHCa0HDLUus2wi0xvTxWZrwIgrZcbk2dMto30CX
IYJFxisGXJb2YUqz90g4No3RTz2fYY35uCscWSd0ORhLykBnBMLq+sqgoBaKz2E52Q/s8T1T918K
nkiT8gziWypGEKwR/7n2kif7rHmHFbT9AnkozWy1iz4rRGV0xTrvqYORjyJEdCrmXLWpVM2uVXcn
oZzSvu3Xv031NTULB47/2QfKhHVqQPONcxf19fMid4QMLINLz3aRMg1vcCImfuexYhTTZmozF64Y
tKMtB5oJBdTGcKPe44bLqZRXkmH9MX/QXLCZesSAWaWvjXedUqmQ+aq0JPpOLs/L4esj0EjJOS+5
6sAlyDwgbIgxVKBo0Ad8VNU/XTLpERjTIDEWFj+OY7onLL1XrWVzGxr8VYXIkTCkiyhOWdRrouuM
C5VQdlzQUCOy9RGT/tFht4ji9YNXDyV/1Yq/ke2CKIDbM/rF5jOxgjoK38yyT2d8gTBHBQu/cHED
DxARPLkBwln0DMGeEWn5MFknwIWSGxoNU1EmuBnH3yw79B+tBdBJvbuPbFxjtvOJ1klCii8P8tYB
YIcvHz+gdbkaiutfKcpXEZtmdnZGLoYaTkbgZ4nN9sPt+Bx7WWId77LEuHtgg/NZ5DXK6SABKHfY
+T9tpEFZGXjeh0DoG4UB2TLnXeg+6QLgV0yvuRqumXauB5q40vQ3TeSnwcf8HuJTTAditx5f86Y/
F8LsLYdOPUPVCDf//hpgy8lqD0DQz1SnoAmdvvQLU19Px3jCYx85GZP/Df8f3SecTqd6f/pNyG/l
4p3hW5woPLVItUb1BNLAtxnNwmw+PBAO8C/k2tNfIvBbKX9WOcDn/W/NJ7b9XBZYLsIGP2hwR/pl
EafCkzrzSMFf58DAe1WQAF6SZ8oaC6AIRHU0ukMK1jhel0zo2NHI/OKvvs1k04cAN16lYJrTSoii
2RiiOUWB2/PmMJvDhUCz8339Aa5TQmQNzfim2Ovtl2SxaNnGzxh2BuN5vcJ7dNbSP9d0pAJasyVB
XDUb+xzzy3rp1/+uUWt6ywExhdxO8gV4n7MhjfnMMtk8SInROsV+RbkvxmTllDWr5mPYCWfP20gi
R80cDqCfDDcRuMTX0MmrfsIjMon7Lut/DUwQJpr1V7K2xOfVkurDks3nAZRo4f37e2HIcW+QarPG
VHyaQM2aAqCaGKrP6uf22gKPoUynKJjk4pMZjUfeLATlLhXV60JepKEvEETumzu/z2/G90wPSq9I
LNc7suWvmDsdvIvEBLFXcwnOVR7bsn2RzwWcjXXzEAMe3s2RxVjz5ku0BOOyS2AT1S0EC9Cxm9AS
No8iinOLqrSfa/X2r0Rz6p7vo8kl4OnFB8mAOSXL5hSl7uWYRz5XMO/hQa7YeWXIO4mRaMNk7ckX
3XF941Fw+OIQJ/DMV55sPXROAH11W3ZfLahx8FNmpXAYVF1RumYzE+ZMpoLskrNR7y/hJFYqQ2be
4ZUYf6hO0v43VWoC8wYwWS24L3puGf3RwgL1j0uzWkKNZbA5oK3y939eeuzn0XT+hHVURJtn6lmC
s2yPoltdOZHkKvRtYq/JMtbOAaSobRwbf7XdA5thcuY1Mnc9RRLXCiOQqKy2k9FaLEtH29lKvVKq
/BeboIT7sF/XR8ahWXXubMGlhJFonCfypMXfTLMBHgnL6WG6PEv9wJ0sX7aMunrJZHCAxWMFtyEp
1R5gRtLIc/tvRZme7MIrFLoEpiUpcqbV8KMcdWyVFecc69rM/CdRwDPP3+bTKtUmt8W8sCZOLZbC
pmGhVWvdw16Obx18cgapxzXdfnvk2SMvp0rXlClm8xvY1s38Lhm2SFa35IQPu6I+wV6y7GqcqmaI
IcyqntDhlhd/yIQC9JQCNd6WL7ZUprSuR5pdxgiKdo6cS6PwcC0nNRrFuFVFUIZCKisqVTD5grzm
9XqeTXi+lrA2uTh2DTlVmrwSUcfzIvxL3R28KpNH44M6FTPt9VvTT97btFyJS0s+4c9XfR9KU5B+
On/k0MlXlLGC2e4e9xdp4YkUL6+Q3folk80KFrAN4HjNUCgvA/SoLCnU6L1zNHkUwHmP2zLEdhwz
z9ualU0pK7bWwl4+INzscnaP/pzPK58xeTD4xIDbh3xH27csUkPGSzTtJzWw65V4dIRmXw9VBbRF
yXmI1HfOrQomhEV21Zds8Bgu7ruAX+4n+AJHwVrv9Pmms+mWd6hOpkjr2zHBKd2Pgyz7wH+1PilL
QxZQNEM6bnK28Q2W1ATPR8k+47ZAWNpUPfrg42PJMPSJ/Jup21XivP+c5FwdPAcJgZpBc8AzPQKj
zYBIlfIt2lIbk/jXX9mD2dCbbt2Iu8QKTHntnLL47LZQ/HGBzfKxIwijZ1rl1qMmDb00ulVYYc9e
BalCYUiljpyu0FEXMUrEbNd/KdmaznMwmJ7GiRnjSGy4FfzAw+yi0MhoQnPI+3sEnIGN6OxKlBHe
luVxZOokydjYS/+sowS4NPZXshpi4hjgh7F6CbbWWAsLivigy+8q43RDG8kErQbfe6Oay+o528g5
V29BwQcYUeLTcmRuxf1oMej8E75K1FCTcIqoMVqHmHNnnKst0tGJ/Sn7F6MPsaIrUigm11BDzc6z
slal7SLo/CD3d12erm8E/u6bO0J2h2oSDmDC+9pIskNHKTSJH+AvuygcslE4RCYoN+iesKbHPV9K
4G4WMlz5Ba81AHlLSmrkbIoylm+gn+aSj1MYHpfguGolj9Vb5qXWkv3zfhPiNSQiD6cpXQQ9b99e
Zl0P0VlCVeoZs12NDh7BrgLI5dY6GUC0QNnPx8pXpbzsHlo6nxnGM/wEhuCTXqvXf3SWawAPoR7U
bxiLWruT41IYJZLIvezPc2g/S4gLl2tqouxUuaWr2NTcs+rPmMJw2T1bkUwHcoU/JZ+4XyRAkxSj
aBhfnZfwU/B54V2h90RNwVAVYuSqR6DcnI+8+ei6gkXx+XsiuQDA+kL7XT78RtDpIHY5UTpvv4er
26UiiGlEkJjrVDMP0qu17tiPGG0bb8NiLyXYJkXjGb6cllYmFUi1uPctBPX6/OWIWN/ozBnA0ii/
AL1mJVPOtPhW+u5qV3h5BkmOfcFavLdQRhVUUECc3mRxfjVe9VAXaXLYFPcjlS3BLlkeWyA3MEaf
mkUmnuhWSn9sXXTEMz+gvr9/BNWDtc5YTF7y9l0O2DWz+7UuRwJW+DwpNH9UOsAzj/LOv5XM6bJF
5brDr1Jbn9vjLOstU1qEW+BPrEariGDH0Axsz0h7YT+pENFeJR35lmlgVp/XbhknwSP2VHv9Y+bs
QKvwXmyV8P6u6Im5A1NaELxcd+97WYIFSfM5tUSSvmIobHQra1sRIUimEU/Xa8uBtFjsKVRLIG4V
ytcw1XQK0pbrQA9S1i/pA8pfOTbMCqsiJJyv6fEU3bdSA35yt84GucqEyfNc/BLG+nkYpVC44em4
Ch2nAmtqtt45OocMQEFZ0DkftML5VpYUcb0tMcAebV6+0prLOg9u38mHn2HVAiuFbTGZm0g2aztj
7/0YgxJkaQa9topwngfNfnzb/uDQtOChqSFE3ffoj3uck30264YcvkaGE+irHGEy+O96XyxjnbWk
BlkXjE8IrKkCEzYKoIRvZ1qtLTHUIQf6PyFCNBBdOXwVDgIOtmacJ4tNNJJYuMVvH5kjJJkNvRek
5j6TfIj3rW1oDav+wiBIVMILb1+RXFG6lqgJt0Vxph9x2H0lMlPjV3ibg5e7BaNzko4AUVsNoyxN
/wQMltvcQwMXBeFPue3l4CmWkW5nQzz72A6R2gMKJTs+Y/q0IW+crCwQoTpNRAE6jNGvVWGqza6f
D72G1/v2v03GMswlJF/sMLcO9YItTjCSZast3w7siSWLH9ErA93Tss85oLuhZ/0ypxprzvuwFZ6T
10dfC3Le1OFsHeLT8CFZHkbt3q7xotDKJwVMcnEJyKYcg+mvcc39n+cMQUJHMiqryNQMtUxyUrCb
TsuUdVONil6m6sudMlE27b8p2V7OaYzrhhxF4ByC5PVyjD0hGpUQkHXDDjZJpLjHMaX4yu/Bg0SM
hOTuS7Cv+HvqQ6BFZi0gAZHdWcI9JmCwU3ibuuBzxkjFMfOKQohhRf0okNKnJys/XT91l5qwc6gp
duFgw03wffb7XiFGFgcJGPiA9pEs5nqiH1HCufa2Mml1ZmpVm9UjW9MRhuzc32GBv+awugj1PsGn
bEKbDc2mHNa/S/PYTCWjA/ttJ1RIJ/PxrYvzlqSL+Er4muyjx43626ihnV42+O23iFo80XMV8ae+
D929fXgSNLhVYDlvOoow0Q+aHX0gUuIl6i2wLXVEy4qxWKbbTP4ugVom26fRBpWyWtAde3xozSmq
BRr5ORNcYETmRLh2o7QIIQwTK6W7rFUC0tkdxDnjSVHKShBX//g0MQYMMVy2EZVvFEz+IezA9B3W
XERhhf+SFnWR/Hy12yXt05Hffzkpn/wiSfHYYKmo/8O6m7/P+iJ2nFktPLFZlfT7lYWLD3BiKOe3
g9OLAJ2oJhOV4bI6VUZUcE9QRBDp7BNtGJFM7e0i090y6Id+208EMJK+VYuxnITcD/Mq6T7SLx4p
aLWDnqTXzhxc8ouOV89fPi9PjtIE4qY7gIg5QQjAr+gLoacUQNRRY72nu4x6eM6ezEQ7K8Fp/KVy
j5qXKcwjm0re8jmHibETM+4QT07XZDoJxjGiCzUmmcKpg+AYCRxzftqBkCav0nSkFPvtIAGDSbcu
I7ojQDX/gyqsX/8kbw5yESg7JqZQxxgmfc9nWS4vDCM6y8omyCgdF874W4QLgi/5iJc2X4es4ZQ3
GHl+dBfjkrgrBsb2JVwgm2o0C5nh4bTVQzjxTV+E3funaf3/r76TprB0HMQ3wg6j3GJpQYBTBd1E
aEFRNSySQ5VwpmeWUAwCQp+uDUBekxGhwv5cLIzE1a/lo8p88RJ/AUu+eusve36bBpY0HjgTxXYC
tEEYM4pjqK3BTsCpQ6lH+4IYAVmxO8YB8DxWcFk8mLjAavPdvFCf6fJsAx0Ty6LuEHo9F8w6eF4j
mM/+/BayyOmlMvMDKWqGkPoAWqRkRcET52WgT/nQoPuAUk2mAE7XfodS1S2Xxj4vRmRZge946ycU
Ohzd2mBfcvKVuWVGqF/eGqZT2iPmA8EBDE0fTmBGq904rJ0NYDVl1dGELS/81GOiQglCzlNbwlx5
t5Rpj3cr52V6DoPtshgm6fkD2BRNChEZgbuD6T3YPbnZ8QmJyH6cHPM1kprXeGNYaJf00pkD6f67
FgBzgPMjaDN2W4H8zQoP8zL5T139kyK4kje6TKjezpStya5HGBkxih2y/6Anos+mgxGRGGXOmhyV
UOR/Q6VfkR+1rlBO1mC30CNJHverIwVohYxpg0bxM7yXKOmcTfDGKKNFqfBjx3/YI1bvikL9QhJ4
anWShNfueqMUJknL3f7zKvdwxYxBdzQb8/aZeulK1OdjNChEi7NMc+tTs43fpIXZH2eYFsi1wmth
6m/4iwXtEi7apB28pzbAgb8Zfo3UpQAMy0bVYrOWvzh8UX+TLIEg4EQ/iP1iEvAsOBfStCY+HJtb
/iv2kd99wsAqu294KJ3UvSuz5R59fhKQ4BLRPmLX7f5sWimv2OENTO+8B5BIFHNMLLn49i/470fZ
99THPHYErxjA97jAkQV/5VBPiCdDAEAKFvs2XR7V99lbwEk4Mu9ZZLKe7nQKY32h4YdVA7SgVyYm
3imxQJjXYvv9wi4p9rjfkRLOKcBqb3Vbu/0GhN21zk7uW80O15bvmFUA7/qQudwSI7VbSBnAP6o3
qRqkLHF6WeGj4U+/XqiFQCKL8zznQl4qaTupJSCkVaq/mIgT07s+4C44wWDavueDKDW6z90SejhF
OEwsDAfipfrkboD+oYooLsnQ1ZWAz8XiWOrtyq49e7OgwSxCilMauWSTldd4FgHHLOQa39tcl57w
tPuJHCPjcghKYSaiviWoI1i5qGaPPIOI4g9ZtCQsP/PSRKu6Wxpu3PhPDsADCof8qsTcY6xqDAm5
lFSvVRdQCM0kAJFzSGfDsOKJ1YwxJ5hUKf++oPbRzBwX26jLjkANzXPX+DmeSsFrbKBlPjIHylPh
+F1DTZ4i1vHonEC+CxW7ikG4h82kWVLjsu0auK1sfVyl1bwQHksZaipZVD3iR8Up3p2tAqk5r/1M
NZE/Av7FJvVE4ruH7dxCLMqdmDC8XmkfRyoO2f66saTinQRyEOUlsRYik+oMzJ5Fy0Puy2W1d2CN
DHCWtlZ1SdiItD5wWfBj8CHvTFIl+Fq3CSL21f1uhCybTGiUYFZBE9wrtzopAiYB+Up8V637GirY
7qn2Bt3af79zflaBJCtH/amhXH/lwBx+fIk91V29t3ZVIJlo8LcQRJfmscKZYH04/HB4NhN4i0h5
gg9lFAJinr4RI3AMjxVM89bjjeoskBM5RpOMNe7d9uctsLlHptQs+b6f9U5mMr0Z96j0G1a2qThI
HOqYe0OGEvlRYG3nwskL8KINUoDP+Ch1ErrYSwyIMhsrcvZAyzzrLWUO9K57LmdVQtriPIMKc4LC
1O3M1hMUeFu9ayTVZNA8IHPvHH6t0feLpktpJfgCnz5jNlbRHqZMmt0gyV76tBW/pgBYJoTk7YqB
USWt+iPo0agPNgAUX0qGPMsJ/J4wbNy+LmhSw5Eu7Z6sr3CgwUHMTpzBlj+9sc1PaZw1TSz5rJXL
f1O+Xwapp1BGH7/CzIZuOHLcjzTQOfyxcry6hfb4cND32IkrmRaXH7S3ZRhTsijqrhZ0jz+v7WI1
AjjBsqxKVAXkOOE29Wa0n88PQ69tbkG5I96sOq2JpwnX+IGKjMyg62YyzP/POMxOjp+qcj5obN0e
MSSFgbrA8JrnW6Pi9qz7I1uRGFVZBoz4Lj1451UoG6sZJUa0NjJ4KsRueTnhDE/bXvQdLk5kY3gw
StTvOZ4PyyEl+3Um4ttikb2uNo3QkTwi2VHRJnezdEhHfqPDHpZ9SxPoncCyeA5NR8+ndnaNBsk6
AJ+SlovVF+98IhQup1Lgr4QEZqWB5yW0neW+g+bLYH2VSS3NcKt+QidD0QTsEkoGoXLwrnNM55NQ
kOMhR3w/w8uhqmYyeVPQEyP01HRugGGI7iBF2wiAOfN6wuHd0dPla543lH6uDqAM8+ByLpLz/Hhr
3Sngzke18QOhvK7tvnNABQtDLSI0rdWqgFqm5rdSFoy7SfEECQjSDI8QkHLFUnqBeCjVcnE4hQJe
oNiKCzjuRipxnymLU8YZXV90ENPPsC0ulEBQ3HuMkIUdM8Jxqqd4Tslqo+cqFyoFTF3BUxg/H8GO
5uOJv7OscLZNoXIL6nLL5k33pHNL3+AL09uXpbWRdoIl01K7w1NSr2mUI/EoPSZnId1k6v2jDGpi
oMCvmt3GgLLGPuOgs9szqwI4axnkWjC/1Oohygjjqklld/YqRKV/TPpog++jU7y5Z0Osq6Y9ph4J
67KBOSGQ7XX62y5O+0Fxj+LWoWiRalaBaTOyG17BXwjjJTk5PZaS3FvyQg3QwSJXiZHoChu6RPTv
g133uXgvUuYf89P4Xoc5iLHfKwuqSU+eoihCcw6PDrHJkm6LKDxD4BXq9MoiKCAJOdN6GYjwzwpb
Xbon7NwATrqXFwbLkjmSo220+KzOLVU1/SQ15qnnr5YijwP7ZqbDFEXJleeaJHkkmolgL9yzHoAa
YQVavw2HUnyk+TuOXDgjYRrDU4NAxJeXvoQ7ifj6ueOlUT1Yz/zN80FLeanr9JjgGop1QyfJUVtN
/SVzYv2UHOmArVmsLFWzVBREnMC/XVdUzKLBcO2spJai3gFCJPz8yIwGxEe8kjBEIFxb/tMS3Obc
XGBOmBr3L9GNmOLiBKuc/ffNi8JNx5PYlun5tOsh00XDe88GDMOgwVK6Htmrvv+6fC5NZyD5UHzZ
yZPlTt/pB+9cL81pXnWcfj3/sV4enrxkBcaR7PzY94/UmlDuD+CiwFqu0Kykl6RuMiom/MNwSIUH
2fkHqXmoPK3sRhI5t9NP0+NzgYZnuSZZLK//6vMg2d0KsZ2pqmgTMrGX5l7QMiJPQzt1N4EHZJOA
AwsFhffiuKVnUnyAWGypnB+01amTbWcgXaolxK1oFPfVM0Z7vJv0yp0T47RVeP/PXpppvrzmW7fn
woZ6iJIJVyTel5Y07L4NHl9JqhWoZ/Zyx3MZUWAymy9VvAO1VQ8GDZA1A6w6b4PyptqSKVTIV7TE
9PYPFsos0VOxc8vkaVJUvcHNlbroQ17h7k1TqK8WcjXccTCeZA2UZ1cXy1lJXyprqBwdMb/eHNLo
PtbYcy4HX4Sh3TeTOPv/bzM5WO6J/zjNWYeyUq5QJRb0hSnZsI8n6UUEAm8edxHhr7XbVXT1I84h
xcW5gWcYvTBXFCjFRxpyq2oG0X1Kw/FySmsYtEL8Ez5CQ0xftGuWpPtQss+O25MWmsOtSyY6Lkwn
Ovo4PpH9Dm+CQOSGWRpoaj6f99j3Qijg57ssnA2TLZzqVGNkWRdAa1odGwQcXNpogHzNxLcJ+TG8
2nWUnM9fZ7T3mH2QB6sncdBYRVEs2XjmT6LZBYre0QVRJVyhwQouhomkzNLLOP96ZrwHUNphd+Kc
zJpyZufkqRexn/5bEwIjMEv2s/qQcjNHAgWMcVwcJNxpeYxzd4Vz/RLq2jZY5mB0zLSDm9FwGiqg
wPwfcBav1r0rQlJlvvMwbcKAgYdVBXyEsSouu/NtteRwIoc3BhTQEnrV5CL2hcVFBARreNTvPxTC
180dvrg9UyZFgs8QWceL6HHwGxgZH5N9qsp5c2blI9LsogahOp8SXetGVtrxpSlQ79lVyPs36BsJ
laWRyBVuwuVGlE72xEFi9UGPF/JzEBEQCT74psHZzEdzOssiDBmokjANgXtKM7EjWglIv+kHFJSK
MuDJt6eztwSB0XPstLD1dRReDMfUgbfEb84c4o6DxSvubEcmQgozihhhtKdhlhHbx9FJsy+ksxdM
yh1cFd19ePTi1tVZ5HRa1J6y6E/fT7zKurM2H982lQzrSk+gE0kLi1oEK1X3ZQMB2HLGlydhnq7R
1OuFbhC1x4ajikIp0TqItlHP+rjK4ZhAPa8m1YxAO5a+hfoeLVFQr6oZ3zu+XGDU5wvnSKiOe96H
0bJeMwucS23ZQlMVlxg3NiwwSBoAwKVr4+edTrIRU3sSXo4haIFmj8fa/oI/LdFZPUKqupwWSWAL
pnrjNH4gXrb92jFAW1zK1vgTL5G0oMYZVaQ9ABGg/JUeiqIWiCS0CI8egPBnAt0oxtNmqzDK8rf3
7R3uVDjZNH8tLU73GH1cYx3W7TM6LVz8p5oA4QCdz1N2dvRDA4EkB+XYmn2MJJgBQQUoSyCyZ63M
D518oFoqgsrZf8WMRMU0qoRGg9g7PSh9TA3rkzut0xTdnQzi/Ujj0qdJUilR4ntdvQn1SswY22t9
QDS50Wd5+kcp2twBz2nXbGeita9EArEzFEEd3rBY39tr/8+B0gezknUjchz9Zd1aviqe3fo1pEs1
LULHD+jzaB4TtxeBa76j16WyVKJOoNL8ldkWBGyQu2tOZnj5aCXa0Gn7cEdY68q8LJ+pBHTwFFQX
gMmPFHm9XjP7wpdWQrCQmnaURX1o9BiCNQ3E+35V7wvjt3wMUUM6Sz8RolGSbO39YkFMnOUOHvQg
rVGcWRln20pRBhHARX1GIWk9CofS/FneguWDbokuv45HPOKkwvxh/DDpPxxr0G/RDLr/+TJZ8+cd
IsdvZa1VixazDVpMC16WV+iPEuQwylAK6zFAaBPcm/d9CoaMzS4vC8KbYlH5QbLTQA4A1sNZuVL4
1GtnXPs9XeVeOfgiZ5JCWqOR2ChADzr1dcMMl0M5qyBAqjjGXHtdLLciygLlIMDtK6elcx4j3HTs
Zo3yDBxuamCFxeZLarfF14xCN+PVAMNBCPCiVE1qfw/UYqmQh8ghKBJSMi/DkZfrBHjCJQy85T5X
hFUggfActVHwL0GycBoLbJvrOoV7M9XJmY+z9nRgOIlIXG8gDoO1DXJJUNfcy/VmuuheX/a16TTU
73gDjllncJtVxHXzjx9/hnuD84VH64Y9OfXWJ1YMW3ZFyhNRLQRadKSQpslblusQPwNGUbIRF6AB
9V0yq9Tspn64RVpdA9DoE+rSeRxXZHcLQLSC9mImgWsoKC3StST3vLYtFZ/z+wmzkz8MQpRDbXsc
FM4ENl9PKqTD7K9ZQfP3J3MLUl84JMbwXcJd0AjPma7ZBT2Oax7E9SvdLe/cUQXWfv4Iq5KN6K8x
jKqhIFALfWfbTKYkcqQ0x8wwewe2yE78ZhCdNc0t52DVGIqzQRhImoz6UMArzSghGCw8KHo0vk4J
iNx+wy6Uvtr5Dg+eZziTyY0RHRfLdozv3HBcaIa1wPO8SNC8Xt/30KOIJcegqPuH4azzVfGbVY4D
cze8zE5v/plagN3hk5sqORvQ/Sp8knO1xFioIv9NmV/CsgA2nLzfg9lrlai7wnXeHOEYaZLUnJpt
SPFUi10TB1WL135ZtsxILJH16nNfmVhiWPosOo+REP0vIdugEaqOUQsnPgh0CBXTIAnaN1UMX1ny
7yjRg8/1hg47ewzrfG+9LUfV5EQ5B5NTXGjSPXayv6AOAcZe1zSWeS7Jw417miyt+DN69y+CcZbW
ZkdBoRLiEi0J7o4R9I+1p/gqTRdSaETWd6gqtW0XMGUt8cXRbg2nDSXiQkTf/A+OIgtODw4y0rZc
Ycns14fbUFUesejIcxZPgVVEgDArP8ze7F99eKuss3xhzYtoBK4CUwMRwA0gHSLYDrAmYmr+oaM6
E/A95HqlamVeqXRPolHdMbm2KIfeCh9vzaC8z80z7o08+dhJC2oSCyp4T5nPw4p5/+ZSb+2TeYVs
ChB+lMHbTMY+GcP7o/jcsmsUnTzsvOc7Q19synEZhpFmlQ+cLkR776p96UJF2omvZJo5OltpvmH8
oEOxDZUwPCEoVc053ZP8IED/n/G7pnKAZD5Rq9ZR45E76uppc7VHDLE1/WyDbgMWQNgQCgKbvhEJ
2LnP2YH50JomzjTZFeFOJ88htoxpqZgbDT/l7s/JmGNue95VCM0Bf3HxZpCfqsDSRydWHXeljO31
kerSsYgjhWvLFVZWreAYu96ZyS3wln/DlhlEqTzP5VMV1h0V5mN5s+mHfSCjfxDNu/cWEWlh9iiz
v826NvDcRT/WhUt3wFNjjN5zv/uFCljxnqoERiIeUoD6vJZzUnH8P5hOu0ZgVr+PqOdCK6ri8Akx
DuehiFSjbcEJQt4xdt2wfc3B7HMDCOxi0kf9BU+71aB0aEtwq6sLvXAOLBr95gkBxuDbSyJ1qf7m
2luElNGRxl7Hyeubv2E+dRPks6LK/L02Ct/46CwpdlP3H2iXyDaAXunWa/hWIdBEpL+5OQVdhmtB
cv4EVKcI+87XSxayPQRCkniSh4jFGXQCuJW+ETU6lQpp4hgI5uHUE7pBKruwy00rrjA21NneRMBP
/sh/ybilXnj9OxqTXiIgOzXjOxgKqmNpl+frNypmZm3D7Vf5c2nYVUxMGpDphEIt3RmhoJFOrsKW
e3s33Hrh7EV3GWP8qeZH8lmpKRYfGq+qM4POrpfjcZQcuf+qXVFQStdS7SeHR0rpd4FT0TO+18k2
m4e9lIxVXufdtXH+4SkHJMh2YXXgBD++uhB5BfYfaQCre8raFutIOekRZvYStlmI/BkXYDBHpi/G
x8hQVVIYc5jaRllpcdiXZR5OTjutotTYcjZcSfOomgeXI2NpTXu4fTysk/+fqIAD3n1jpgjGxl5g
apfAR8wNbN49pPCuZCdPzBmxQpgk+S1z9Vc3p5qLuCyo1uAhaS6dFBJiblRg+9d/uG9xvg4VT2Dz
KQ9tgfldpqtNsnuTE120U7sGvDM6rOHaGoSxy/2XGk1jW5xjXvRiO/rzeYMj8/Hj2Cp3PNkOQJDe
VVvaQOcdrQIMkSHX9nzw2pNllceWEhu4rgEt8ZhLXwacO/tVeroa4YcC6mlFhfFqGx2KUAGSVV1D
7+rI1VV5yqJevJCEeyoozYK+pjmwpBGRXKMvnx54xILIFeGTkZKABIcdFDUuZ13r61dk9hSONfdW
KgfdmyY1MRi167E8HEcWJJwwEoSl0BBQWFmeb4EI7N0PbsLG0E76lxraysrxRlEGkqfQZaBBliAF
Q6HiYcq0D8QdppaqRY9MfxJL/lTD4mN222wQ1YkaZncHZufKxJ/LXXhACK+ZehQb1FUHA1z+nXKA
wNeyx1QYWHPYTXlMoaUS+Bq+gQ9bOzHLUOGYwcMHuPGmqEjZP6OTDKliNbtTbvO/VhWpAtvyrE86
H2ACT8d5fD3152eaQ8teRILS4tBErhTqMo2nqJQ8viMwJlxFLtYQe/3kp/CpfnzoqAtLA+m5PyLE
w7ARgRq4LVePUKb2GCRmHaMVFHENkl1B6oeGTFD5JTN645Gy7QX/rd9U3ffPQ73zoFj0nJrGH/Ys
psOhbCPSyaYDsyDh7+NVCEO9PIFyadxXPpL9THG3v6C4LQ0sYz9PHGz7rD9Q8zcIgieFWW0RbnEJ
rwMbg+2MMkkRdR1n+a5ClK6DLEob30bfESf9p+0lcJmyQUFF3jhg4aURxgJoc/3EQfNvevmegEjY
dxV21fJddrWo8VLY7HH3m7ME7cGCx95sUhD3/jNL52/TXQJypeWrbC1ybFa2QzJm3CX7YOPn1AJA
k3WSp2Ta4mgbavpkcWKDinwQQAd9sQbX3jSCcSZPj0/gMyT6sJdnZnEOBQgBhHZ/qB4YRo2SHLcm
84HkFcueJL2fD9kIQR1kTET5Jy3OTg/zJpTxWp+T33YjMh4bqlIuYD+JV0RgFmmbPq9XV68VPZ67
P9RkFR3p0j2fvGC487h8pH/gExCgOjfYyrEA6XErn9khpf3gcjQc9cJRZnxgP3XaXiugQuiSUTap
xG6qClIrNiyt+Mj5BahNjS2X1Yl904vz0t8WHFYcLCmTpVrFSp3SxoFKrGnm+7DURZPEM+pgbQhN
FIqMssz5zuk+tCw4/E+zMulF8F5ocuUlecA+pVC+ZTk7C5DyGgSLmFFIiX6Vn+7fJdcE/lYRkmMV
lysrfKfvwKcjnmuwjDXR441CKBZuKO+zLlyUexUNhtcRzVj+aslu2gVbPn9Fq8aD64ddqydR5qef
Og86Ruf7mR+uhFbfKbuBkD8PyWdu9v0Z59C0OZsNaBJXW9ZaAXXIad8v7DhRxK4g8oqVSkehf+w/
sGkTJVmlcEVO7IQcVO+SVWX2SmKXgX5SKzksOIRmQzf/FWqP5ztqgQyRfuB2D2tl9rrL6DWcpS55
vs8S3i9rna/4JhWhgKcfDf83k2QEd7VJz8lYjbdbalOnvfFozqcsnJ5CHekacysbDpuZu2drV5Ha
VIKn2yP5VtQwZoKsgM4YPJp8uZNwhFoHshe0KJ51FMKOKhUkBqu5+VBZa2+71oVqE7PRy+wio6+f
Lzxlx4iz6TuPadevExuKNKx7rfW2Nu1L/4bLnJv/8ShkNPhYE7MPPXUo6O2LOfH/vbvz9WLrIi+S
/GKzgQkERhMso9yNDPht831kh09DJtFAxbtEvqgo1JPDPANZdtYZRCvgkXiXCVDCytt2quEJhbFq
O9easThBkQbqyO3VI1aulwhSG+RzQn5BMPWnv+aGZt29qRxHdTxcPWLp4Jz2dvjUCMhALV35Ftqo
p50I2AeLkFwy2KecI7GSoNYvdf+3JtuZKvWGVI3kiddlmN/3pjBXs8VOMx2IymmtyR8E7hPr13/j
IboWKk8ljXFDoNAsKNBmM2HiYLm1ZWPZ/eED5tk5WD1QEMGx0tH2qAg6odaAvN9dRa7Hq8rfxAOG
yr8bWcw80LWxb70zf9R5f+UmQTYL6TPqGJ2nuzDFooB1bNHTvV79xXzI5oqnr33IDRDoKposL1hS
6619GFwHFZOZla3jleTong+ogNTfV7rpkP5PAcKE5HUgIba6KnDrA3L8I4xWHG968hfBdFNxCEGD
2u/fRxeMts6M3ia+VvKO3wFD7g9yuA6OsBTHsPHFKrUJSiTyOrVbIvDVru2G1m+DqhdBPg3T618C
dl8+ksXe1U8yitfvnO5mYrUBEf0bLKAHfM/uQ1up5k1C5NHENCPb1S8Y8AXMozJW0m+Pn27ZdoNL
YuCYY5xuVilXia/jTUp1npsPIswHCxV1vG1c/RhUb767HO+PpN1UgTxIu+8OxfJJsjPr+yxFhnfa
Td2SOTdCxrVrs6n1Pvlvgf70ns2mhj9TvGFOg7r/ff4TE1HGbfTrgVyLONjpUgg5XxfssptFrpYF
Bhj33U4BHvdexArMo8i++7nzn7k0CENjNNmMe3NVz0s853Fu8oiht1ZZdDnLk3FSHwI4g8HkantD
Hy3gJH1DytEHd2peYqTw2BYerzBLev19CtKEnismLEYtsUpqaoI9RxSSNJWWI5o1JQ4OSKU/+m+O
+MmhfrRAmpUPLS11VL7b57qhCZ27lluFywuiVfZ5QcPA0C4j2qCISQtU91v0w0EiKk+hKvB4xAni
YRSedxkhCEGXon5yEzP0IVl6W4go98ajAoaZ1t0Nq1SNQzl+QTMTRttqcA4Z+dGzTJ4s4oKngrZu
QyCdyGH5p2rd4Oi/MWEesgiPLTHzwYnEYD2oUsaV8XTgnSEbgcUpvx7un9SQYYVF4hz+LTMdfkaL
jVc+cAjz1xmLi6ca0nu93VhL97YQglIL+pWgthbYCGr+qdN4sh/RvJW5F3fW5RBj3D+rTFToFHCN
xTiMzXqDwiuk4/heTJhrJLtwzYw+HbR//wmaAA230lle0qRzbNL2YNla5Dt44Y08DZfDnAAzYlOS
Gh0TgVlPNm05ccRgqkPtyWV06HcUf8n6IbjbgkjMQ5xtLGXHHxv6wTLkxShqxKrV2uVjllfyMHMY
lP7TdrvFqRnxaBVtjRyS1/4aA1ky6/uJ54KpJXytzru2U/UiWQaElOUnA1AYtTXMzwZ83Edx2w7M
CHHJTmdDgTk0ZCpuIMRajLmzvPjjrMvV3ZMxBp4S1ShtLQMFdeHdooNPMB35M3aGMuCDgAcc0+ax
WUAGeJXw2MrDJlAEpsyqxy1yHQZJsiQUYxf7AykUJxpkAXo45IfxsPTIqlu45aHVzPidBLKQCQgh
lZ690O54tQtZLf1LP6ja5MGzs0VDo5v+Go35FL4NHpkowJvMIZrGY0vun7RRUPQ+cyM1SQ3PEZm9
+fxESSViBEjIV8Wimfpd41s9dn06HFySAbRosQywDFVYvBvVPBi5j0SPmpVG5WogWL1N3MqPRZY2
VuRBQ2KuZZS4x7IFWGTbic/cYN811fgVDDt3uLJ+X4UFh4lBdRNkssSYNB/PAsUiBVjxTa8BVNa/
PwiUtXek18PiT0Uq6e5Q/tO/ZNkEoLY7lSrgNiH35MSnR67WZWm3U6dtIU8hW8AnZIl0ta62kkRB
2Wubsz5QUr8BgmVmLlbBz20KbWVwX7Bf1nPAEK0oP0CMvOoVDxrx3DI+f4HSnTjHJUgl85PDWh+l
qaiZ5m7Prw46FIwbNpWVYUqzhQUAjVoAjkP9g06hPqmlMe/vFgQIFNsqk8GKQBDq2aUZdRmLAwAR
HEckzl5GSuikV+YAUL9ap2ep3Io9aNyiBdKQ61ACc3vD9sfRQE82v5CUaeu3YBdwlJCHs7ly3eHJ
fb2SdyvVSqK85x7VdkchoeNUuplLFwswF/0f0l4jjHQRWSIZb5fCP9CP9WmaSImF+exdrwpaFYFA
RVJUKFtEdUt24jm2idhSqXfBVtbrVPc9qm7GjwVF+iLUJ+/CbLh7fyVEWW0OanBGHKSX53nONtYh
uG5eQYDbd5UTqI/ZPnZYz1A/BF4RY4CzRMF23gVBB1yhJd37HZyKZHSgSoYAbuxrXNSCvCVSTRFl
v2MruMgQ/NOVpbi1XL9865BZwgdVp7boXZrf3Mif4zHhQzfUhhn810t1J6sEfzt41V5hE36/RClc
vNJsJDExvjGLR/xsE6RUdkX5j8/4xzAKtCdwuLMA4G4QwPkcC6c9P9zrwZPHuExEc1zzRnIXFyfc
9qHJb1DbtX+/C9QPkS0pH3WZSG/T2c1tnYy5HAn53BVzc44dP33LvrRdIte1S0XhWruwaQTPDq8g
M8lhqj1HcJK+7bTUaAXDdKWgIeya6QKesYi43wTbHQiUddKzDe0MHCYtPAuUXduC0VofWGl5NuVE
7Gm+5CgZsD896duNZzeOWOgwV6cMhkKy4PVIDOA1epyF4CNtO4zai+GNfNBaGs6+d1n19ng3K3xc
jZpjgc4M9y3JdqVPchXSpF3hkPR+o7N8WXkOMWfDOkRzYMs8Ux7qJV7sh80OPZEQbPHMVlT2h7pT
VAARtGoogEHpmdReudWVwh1Q7W0rdk59devmzX+3epbNpfmBOoJgMKvcxb/TBMaNFaKGiG1SefNd
B2FZL2O7r2VrttPjwExmk2rb+4Nt1CWU4uELp9aS2gKEr7M5mTfB6xTAVWOrFLF8Yr8rDDX0PJ8u
up40m+pDhSznbrtkpqgOlZJrnykOniUEPTM29joXH99JBgVr1wVwdB10IJwkX50UjbNNvU0gDXQu
FedHLGG9vsz7KMJYrsOJHK7u+myLPNZQEmyfbjZVGOoFzkLyI7fWy6yMAVpdZ4KOP1b0/DP54EDJ
Tx1wqqIuhXWy6T/WUCxkMp3T3QqZUGi8StYAwC2QRZkfbWO3MRHYSXAgXoyxN/siJlLVMsZBhxNc
OxQhT8W500QiJgVQEtMddBCHq7d8YnxJuYadVrStZoVm9IuuFtiGvYpDAU5p5c4rRqoVxEi0JBEY
tKS3IkAcyArCg1roC3Wkgi8rAYt+V+yHqtdhoOFigNry8u6GW6mgDPkcSpgNeiQEuSWEd+Pp+9/o
DW32x3dC94gEzOHKCEZ/6PpME+A7a+EAbHVi5/nt6TozHJsSBLn8thp3ZBbyHZkTy6mqfM7dv8ch
TPXsOa7Ouf+o1FHg3XTOkAQ26cwbgyJMk5q6o/sTMOvqZUKxKa7JD+zZoFAUp3GISQnEG5zbkRO5
La4RvHNTUx+j4KAxlwfGa2os54Dr7vc4IcIBMOvJEMVerydc5sveTl6eXgigENWlfF5xCqTiAam3
ZinoQuW74gHjL4gAz6y/YEHT3fQcR0u2YSr2+MaDrqKahYYbZuq50cWWAi3OwPT1Z/D2Kld5/MTP
bajh2lwVIDMoRYZ9WtRYksoKs+x8p9hfs5Hspe4pR/Z9s8cUIUX19+IOpjE6GclgjED9YZp+gs17
3WHAfU0uk8Nog+mmLxCYoUvtLPisJO0FmrPxtojgGuyqQH6OF++Jvfnfi8WFSIi4oU6mXuE6Fvai
27lLv9ulIvUwZrnHckTQIJlg7eYKzYVVlQ+OowlB2qvTaYDHQZJNf9IG9meDhqc+y/NHY8xMj3lk
FoUbKLlwPsZAqkh6TSuRhcVN+KvmaYcJD2kT6Gj8ReoWhBbUG6zCJrr2GFXxSQeAEBOBHt2r6jMy
OHeWQBUEFGq/xhE63UhbCdPLJtXROLI3XMOVcA0J78G7KF9WfDcsDqvb338wVkEF3vRLytwk0TSX
iMbnkDlIMLOaj97BZ+4x8vCL8S7PXM/FmeEa8WWprY+Rj88D/GBUhdMECT+Z8DZddWSjpVT9j3DW
EjULhGU1MhfL2TwKhCLXtnwIIBPuhDRW18w9QYHiLPtkkapyBdwFjI+oKoqjiXeRCghpDEZHQb5d
S4hCqzkr7p/3mAyj6F2eIzuUDleorAs6VQGoTaBkSLDr5Sy2cDOMJJxgtiH0DzoKFtR/ndvpSYSy
SbJSf6xs0qdeZgvZ5HXEg4AioxibeimgtSwIVCagRZvNNSkN6zJavmgtdy1Na73C0GMXAMmtghVo
gZDl/9I5/8dBgCobD1GVJwx7DzTNm1mUyr5UQliDeW73+m0pKGFvq0clTP948JWfFiVZPH8GeBNj
B/Kl5AnUVWfnlWU3mm+48RkyfRFlRtOyNlmX0Swz27oyE3T+1B8sVN1Vs2v/djpCAJchNLZw1dH4
Dvfzuc9H/er+wF14wnCua1pKhMOCcopBepOFnz4muuyHuYJ3ZIl7H1GsaUbwzD/TRJ7BaX0jd1Ns
NwSW9sga3NlKV0si72oBvAe7J+E8sD/BEdf3hwqp4I8Ghq4pHq2wvSPbG/xsf2aVo3sPJa+9yISM
CKs3b0mlllN8UZfhlhmule2Xy/NrLHXoZrvBERvA25VZmby6cknXIhrRQxy9MH4P/jRJben2FhzZ
Ls9fzleo4hNcEif+VbSoCoArlLt7LWps8w+tzvdagLCqRnGjRBRKCk/oj+8RIaY6/LI2Jke+cxfT
LIei6vHameQUIpuDpmqiEOtMY7e1HkAxXnnZ/YD46wU8tqJJ6jNMzv//A4j0G4jHUvuQrPhQAJNC
hBsBikqzuaVxOYoo8WL9f7yU/kC6JoBHHlP/JAXH3nxfXNkLxjOo4Q97vflRqArmlx5zxW3ap2I9
/wUb1e50XsmCLkrHCXqFajP/vMPEp+gAFBP9rSKN25lRBrIBCHYlJuVLgSgjHcTF9NtnpR5c2giw
/UDDijfd1buUdCoBIcj67FEzQtDxlRnriz5cGYOIWPv60XbDT0eTP+dblJThiJzIQrggcM/fomOs
B3OQMJNqHD8zElG0aXmQJIOwvprqprxWO0O4o2hUWiFLqIL3aGkRAGGKZTqXg7uONqameEpZz8H5
zWr3F0slSmrXf5D6+9jZl3RMEL+Nc58tHiwp5uIPtNGmV80GBSwFUKmrEjPsKjidVau2vUeZ7zTV
J1fvrWHucRZyUKc/NzwHDxhVNez9TOlpytNGEo5gYusWPe9gjkgHHeR1EtPell3d5tWNx/dWeBy4
C1PF2iTsv3yST3bn6R4BMHrh2JigLOREPzhxsixV7A2ftAe7afTeZD/4JcYgoEHCUYKx3MwWOH/3
nS3bi6/Hg4VBPhrOe2XORnPw2TOqHJz0Dvn2E+DFptp/Qu5zdwcYuW5nQOOfNHd2CXEXNmhQmXpv
fthtpLVeMK92CLb/rKjTUJR8Ve37ciy/ZlaOXBpC93wd4r0AWUXPMwszHRJXiVHhT2nKuv1YjQS+
gwvXFoZVckhrCs5+dVxCN/C0yKPHKJ8Kcl1BdNGpTgU0smab8EHF6XH61+a/z7HxJsLWq3V6MTIi
M3B12BNGJJ8b8yZY6rxe+fcKn0H57LRIabP2Wk5X1TMsqcwXK4bcM8itmrq0fWr9KresTbr+pOB/
P5LfjSx6to+XCS3SWOqiN5d0WPZTL8haOuPb+ymjCR+8CXo/CUmIHXyRVE88ypmxjyUd2KBHAhwM
w7IVo6D+EN3rLoccGkMeqlsklx33dmjAumkAtHenwpiSnYNgL2FEt7/3DK+jjEi4UGOMODKBrCNf
rxpZTKhING1lHsUS/N5yGlde1N8KQ0x104AOdq9hFGnMgOVVGXcb3nuEdBOoTiVn0lkVGkW5nksq
TsW+oF6yp7ULKFH2JzI8Lv1605REOjS0rWL79e58xYPtziy8BCX7KI639bZmqbtFEvubEAqK72po
g2Jq8L0WCSnu1b28+tl9I5HHNKLHf5TU56+tCPetEu7Ps7LzMYWqkyKNkzUGNjIDvxxXHWF3rFPf
1SXum0m5iegBsB5Mo13zIH/zKLJ4po7q8mvkjXmrfPQF9J/D5cwtXmBm6kPUk5i0aePeHumu05wo
ltr2FfAgnWXE5KxrRDKsObVMmSHrfv4ErZx2gFkTDRdXcXkkfU/YMBTZflKTQy2c6LQI2lcgZhFv
UpXg68hUuvPxcrVcEeiquBACFzG3tt6DCy/PG7A67z9o58e38OIoV35MbWeYcrfvDPeKwXexypDC
j8BVq4TY8nENs+h2sDSpDeqPHlA2ks5NrgG1MHM3kTsAlAkmGNm0k76dGLh/IgPpVxMjs9vwXyib
n1O3m/a+X3eRt/G9v+ST8Y2/C//O4YcDdns+65b66/V9LSQTND90MKauviS7dj2+IQcYbtyYz89s
lbAw1p3MkXGU2MOItbaynMHblQSoFy9FumzOx70FQfvaYqpQmQHpdwny/rgp6mBk9g9qc/DFvLx3
zZDHs37OEI1NskqerfMpm1pKCsE4UbTAdtFNzj7NYIO6+VA2G/3V0Ulf7XM4w+WM1Ro+At1qmA9u
Z/5eo0nB01Zipcbt6qHBx52KqP3t0OfrewBK6FJGYP5NXVOuRMelkGjjBvyPK1LFKBXzKXPcHOxF
g5+CpScB17i1KX0FbPFtN+dkowy1aEua+vHe8LdzLn0/fATnDtEQaUAfd6wgZE7qs+fB9BKsmPCD
Lec4c7mkGCIiBcbhKI0F7XnX/3NEpMyCT12qzaZxjTeYS+yrBD4418y/o2/jyo+VtSzfkXd+9bsN
6zlWDbreS2GWReeW02JhRyBsoZypU4UR3IOqgGw0HSecPvZLQk+hQb+csh+W8g+kvnTA+ZLvv1md
jEq7aK+j3ztgITvB7io4QC9pjuLW0lc1/gh2wfkutylWskzZ0YZq04Buxn++RmIBKhzv+WPYkInM
KGpFJ2+CBrRfI6hqmBf8XLZUcXLmUr1IRdpvTSFJzLn5zfuyPjxAfwMkUOFdApN9Gw/w8ePJlUH+
DKo8vRU7Xwd1AHv0Rl4b0oNPJJktaKk53FmhiNlYOO1NTkh+sPGY4Iwb8Ny11lj/rcqyUyMxWlII
LjVDR9NDreagKSFbmoFyo2KjJ475zs05fZg/IxbWlPGET+FQS8yDZD76nev0nlFnbQfaTivXk8dE
aYDJZidR8cuvhoG+FvRzCvi9nCsYluxNMD1KRw8AAMIUJnD/oOhVTQMbTNLJlcaWAJG2EyVr1B4l
5nHFv8nqBhozLoqBqGi5vGIGVivFILPnmO01sR8tcH7n0x0WWtR9TA++SL27EjJij4vEAe/rMM60
4R7MeMV87ZN8k5wSOLFx/I9Bj1q+W4CzjVjgCjLQ8bqQ8vF/p5YThY2KCN9o1CXgfc/h5mn79vlm
wZrCAdSkeo2EvWIuKCyC4ycD2urtLzJNpx6pq5mwgTRMkT7/brFLnmUNPDyxGEPQ6EjbuSwWq4vb
y1jmZdlEuUUJJ5GzC9AknXFhalV8mEx++xYEsWUA0/vBUysmqRlQdU6+1LlA8dNI9QFWeCdy07Sf
MIruKX0IJOYOm9Hgo6jLMYETWafef72+e18kz50CK+r5H/sRUV34zt+dDqFtT6ThaHnqCQXL3Pwg
jxyYTxHBIYYyqmHoJjkOBA3jk25ZDq/x6V/Bilut/s42ylcnH26hB3DpnRy65Bnu4oYeyfeBsZnS
6+8OVgqVqyWB+B9dkQPQh0CukpMktLl1eoGOUyUVu+mAtSE0LuBXM0dviYQ07QHLHn/4kSt6efIe
0gTZ+bni8K44wRvGcL6k9PN9RddbPBp8DKo3saXFbgYchvW/oEPVkprQN15UjoFaWd9NFxZm+GO3
QlVqZhbUhb0Bfh2g+1gK3boHKG4hMRrUs10CSNXWyBZl6wan970NTXxRiyhFS/J/0Ogjfz1JwZfd
VbENeOx0hzxizgDDZdlIZroPFw7zS3+Gb1ERcklKhXdsqcwssbiwgCT3a4jjWtzAUo5c4siGg35T
PehNE141nupG12MGp1GA7O163D+e32P1H9PR8btwKdljk1UaXgUbhPWLuwciMfbRk84DfZXEs/fL
dU8J5VxdhGnyxvWsz8OGoMwykbjO1VYym/87vTvrhdE1qJ1GV8GbioXiXJd9RW/fDpwxRqk+BCzN
u8d+YoDspY7s1kS8I1GqJ++AZzwLoqiEYo3GcBWSNtzDoVMnYbtv3Ur2I2JmYM7SsATQnfv/bPcf
X6QH4ClmkX6ZiXWe4TgSH8COspBnjx4x043qgilwbBZJoZZ3F4xXN6ujF+83PitpKb7NrXwPMBth
RLeXbrVdG/ZTji5htu3MShSKTUL/kiee8kez1O7jBBbrOn0EsVQsFSASuHhAtbAlWY9IzvYsJM53
eFzPDhzzBlvYkGrZsWOHuxPDHAj8RFoiCRcFizeysUyvkhPFNoHGBpaHKRnfZgFN3LLfxPFDjCb2
hD+Rjbnkd2638OjcSVUZII/w3W/qWm5bn35ylXrMjTZAinDNDsvA0dD63BxHPVodadCOIzPkfi7d
6kxQJbV1MKo3o/rlcAahuZjLM0PYAd8KnVvMs09MHKAwzxJs04jyGwAS8OxHVMHIsVQ1XIDy1z83
XZradmd85dOTxUM2beX2DKqP+V5MjWrpgV+H6cOvHoFZQYrR4XACuUYR+ZeWLl3R4+S9PdmNgleW
rshpKVwwgjgPO5hUFWQ/rGLCZQQsLjUycphp/TnoTXAt71zxj8oQ9qA0crqmKXVFhgsPnJ77dLFU
Bvjw5+o5w/GWnj9Mq02HnvSu8gDhpxHHxAiANEimvCK3WGG78VsT28mo0els/+3pWNmtXjIEJ3uj
+s5Yw9MSUTVZkMrGChyaS3EOtAtZ4ip3djrnhVDHK0vXh0KkEyE2Vxe8HasREB+bCTL6gccVUBFQ
RgDnUR1iSS/TOjMsXhc95R1o6CwEjAd1L39u5BN8Xy02b9j7pm+3dyDeX9pz0gKUebBU6rUh5ATx
vXBYDvZE/gD2mah7f5wkkrcaY3vwj9ruLUGYd1l1G6EZCZT0o84JK44ydh9sWaOOCmX2dbLJpd2s
DxfqAh1p6Orvr1medthyxQHnfvRNAkWFMtwUURTgJWonVIi1wzJ8rhWUH1IcBF2vQ+uFc0keX+lD
dbxJdrTjJKi6ezelI5tEC6nKCc8+fXO1/KUwo4dvU0hmit0Dbzc/qnGzy1YyIT3D5inTKbNof5pt
+sIuJbN4aW9OiZ1GUc+Mi5j/HLodMbp6HzZxHC5MwLCSltpYVHkM7AKfhJ5+anv8gZP6ryBTqhkq
f0ulrRbPY2+ofoXLJL1YRAZP7pWCWeX+mm1UCbI86ZezFFz87OcpEbwO/TjU42G4gUriKpi7I4ue
dTkRIfyOqKVNyYSq2G1QEfJOQ77DrfMAQORQSLpjjb+Q38mj6tV+i5yFEKAP0kvTQ6pSUDUGUsCp
sjBpJcxvoq6jf2HnP6Ib0fcU0jxk3chD5BmcdcIEzD54hVOlCnM8IzbAra0ZqG4UiZw6u9ncrF/M
Lvyp8LJ7peZ62cEMWvbpwcc4+KDuUi8V4bEfhKeEpA8TDwF9okQSIZckYNefekj+zGAZ/NXQIfJy
XipvUFQTbz3L+ElF+Ebj5OUmbhdYrEUgsXOa4oKj1WJJjL6KfWuMZ/n2qNvRBgRsdYlxGmB0+3Jl
qwgyiTXnN0rouAcHQ/mE3IROXFByTTQH5EUowJXaF/Qe2YfRordXHeamFlgTiRiFQIh+gp3mDBZq
mNoO0AoUWCvdChmNkGJ84ov6+ibZBIMSKAhRVBBDn13sLKWwaLaoc1Hxkop2eIber3BDnwJaGXaO
W3QMnK7oaioomKzYgzznGhjs2uhaeq24dfpRIiBoVtnl7dRY1TdcYBAHbLceaZDw6Igb01TpBcjg
fHl0KuSxaXb+qspV49uHfLQ9tNFe6LGysTgtiWLeOdxnGBQutRnIPzQDjcZ5///HnTrEME/4gho6
ll+TUqwRWia+12I39iRCxyOaeHr726GUcLE2V8dgKgenxXk80R0GlOhvyWi/JXlbQLRQ80/UZA8P
QsNo7HuBDQCQpIZ4qHvsj2/N6mNTOem1ZwmtdBmSm9bLi3iQnzGVf186HciqwC5gnhLUZGOmAyAd
waYKeEWOKRtfGXqvJ/gIZ+mu+O4tfXjGoRFAiVTUGOmoo4ydldSdOk0/VVwUeUjsZ9P+Yd6TuUuE
n+g9cT3s8NmUEAYQhvPA2a2ZXdoFeRh5aZn2EZLKV8JwMBvBr5U/IMyy8npUidGnAE44M65MOe6U
ngSw8+HatDliQDhYV7PR8KcE7eFSSTtDyB5WcldLCJrbBgc6SVuJjsfzA0qYmQKTTlrb1oeW0Z4X
P4MlFIVn5kIYO9NLOxPnuMcO/H2RBYu6Y/l0NJsgwbOpWmjdMUpLfNo/dxvfqy6pZBVR2NDmnwuo
MHQGlefcUTyHAEPDgkatiL1fYWye1N/AVLbIeYRk93IrIfnQhllAJzTlhPl4q7z3ocb7gdpLiBa3
M3HdZQkfpuoS8p33kZyRDVw7Yg0Y77O0iAlSTlM6lnB8axOzsI0IHh86kSRkNSnMy/SdS0nIWICG
AUcSsSU8tQJqmOFD0fL8I9q+9YQAUCHeS+O5gdV5rvqbSx2dncdVj3luU+qF9eVazoR7fln01uCl
ahGQo/GZuUyJ43F7PBUHQI1QMK1sOK9NUyZ2VRYXNJhNf/0by7w+p6jpXyf6QTFBeUD2z7cTLc/s
1rDzcsZu8o1z9MBSYZp6RVpRdFDBHK3YxNkCZhUJzT30bW383lU3B4CZL3ijVrEwdB7wzMU3r9Lc
xSoEnADbjF3QGt60zP8nVZoCZaVpudLqVQQjpCYfc/FPULIFL02q6tbtiBgdOSQoc3Y0UpBQsWlE
cEE55E7rJs5MzJY0LRRwK+igIIen6baClb6aVLaIuUtW3OIMepvPTK1vxFTMJiehBrrldVr0+Pml
qg4t9iUMHIvf3gf0P/PeeNHlKOEKAOpbQxxQbbysXQACHY/X7XIjB7DCDRadoQDPgJWSkzO+AVCM
nCikz1/47gxHbPCzoyva7L8rAAr8CJ7TPId3nSP+mQqjr7xTMfzccMU0Gb7dbRQqeC18qIrpy6Qn
I/Z2UUnHxy3HXT+bqQdnABGpwySKYp2CrYf9zsKg+SQR5k+PT4O9IDxQrEP/IWQP3zObZT0hjkew
2wfd1mvHucdXpriEYL/K+YdTO2hfKPovjXx5WygqQzcX+oL1vvqRJq8nm7oZQlClL3b+EPOBOv4x
39zaySZy8LAaZ0BtRNxfcyXSh6wRIF0ipXqsxUUBrbFNIfMIdq9hQxrmdivsvB5esXzhs1QI5ot4
3JC6hdeDZqdpc4qiRfC1Nathrc9YVWZCt8E5DlKajjX9d+szaunLoQVYR3YDMu9QTlflIUvv5Kwo
0z7tURQv9NLIUJb4yNrmp9Y1cAzSVPwmKc4jTnaKsfNvC/VSbm+uIYoZKstpAuKthuFjBaSHp/l2
sB1jUOcV02JJblsXWRsQ4mgrRro5Jz6rZXdAE+ZBkqW5yIh4hHMlcXesgzQ5UjXwlRRM2emZSxSr
kXSv1h8X1ChjDMfQfGGrQZCVUe5KXe0Xv5d/bQg49yfAqAldMp/5qXcoa9ERiN9a8euXO6LajTWh
nVd6+z93qrMIhoHlPyt3LaHLOex1HWamiBgoSOoCA+N5W2eZ5hOqCvXDnvKJPVdKL+zeHKUSncmI
qUbY6Pv/WZpNp1P44QkHwV15UesRM2rC+hy2I29L4CdUzpASUNYfwsl/YuajFC799pCchhW7y443
fKoW+gb2d3YZYzJemVJT3PYjrlGyjFMVDo0q3wSIQnWib1MjSf7kMwljI88Ggbt4GUVphO7YkJkm
4nIhZnM2c1knD1vQA+kCua2xSgmRygEK4BeoCwKWA+f5DYQwOVS0qIjwC+T9C5xhF2CeJya8nMEk
kPAbvj615aJK7CXUda/WnelUHV3gbQF2yBxNFc7I3sfrNDHuKT3Nr2D85gG310oLnN+1aa3ZxPEx
YDymLcjV0Guan53pprHv8ziTP+qaSeSpXwnJAuppbWleYXynOoQbdcBS1Y5Vw0vd3q9SUvVWzE2Q
sVj9KI2YQdhdJjCpYxp3HQ4mrc7GoRyI82j/cIdWz0kVCIcC7J4FwS8O0nYk301MwCyEgafjjvfD
9CyvO2y3q5km4lxJ3lYa6JLcYT5F6Klpm9Bhvn6t0H1D/PGkMYyexuUM/LBa62z1qDQm54TNJ+VE
bW4VOGzBQIoyyxksazCxdWi5aEcf+fThonCKMkhRrgYjCBYI6qCYRPuqCBu5apXDSChSiJ5MnMZZ
0ZQNSLNyf2Brmt7rBEz1936ZCHSHB2QmspHPnJDFGjieEYQmN8iQpXx68J9rHd4xH1/KqTviE6+I
wfKh2T2Gm7ysfyCBPm3HaFw7eQdK8gWPbSlp6k6fON9agntIFPLMlABDvgcu0ZjC3lObbMHppLn8
wKHB+YeymvYpUZM5v9VjiF7F83NKQkAhzwCdI84/dk4JPgFbG2/IWM6tZHtVO7QYrSfRmSqLAt8Q
hjq0VICklx9wYJJzU50xQeG3eZ5JLwtPrTQmj9hN0qfhBh5joCt/kWhH1Z1O4ld6aggg0diHDXnG
//pww4Wm9Diw0JatXSzyIl7YrXx+6O0pqvUai+qt+S67EHR1Z0vnzkOsY6vvMLfIi3w3mw9p+de6
iRJYoHWcFNnC1iIlu88CcmSrhGOl0L6x+5s1a4TyU8Fg7r3bvmKjkE8NKt1eofaAOfzqABFa3pb7
st5JYwfZXScelWHHVyV2EG6g99oN+wEBCRMmGhD5mXN1u0xF3h/ixdLijUxLDALSETyFTQYC4vPG
WE+bqaMU3vNEVwed1QimJWy/fM5BT1uJjra9LbMNBDZVht2rc5rEk+7nOLcVCbNTWNyi/TzpW1dx
Zex6WbT5l2/9jbiA+ILJ2L7somILVgF3qmY444h/k1Ov7q1r8JkIwKCKmKr+WPmxkRWZqE79LnJW
PzI9SjB3ktcF8PRe1fzO2IAEgFuTzHUhUoRqlVvZlT7SED+hAGHmmqExx1Wjh56WER08eDqD2TaR
vcEKC7aqBklCRRjppFL62dh8Wyf0HnWgQuagngTrv45uQWTAmnRDYXTQHtFg4oPiMBs9lgtBAivt
9qBa4sIK6jaG7eudrL7oxyOyg2x2mIrzCKX4h2SFRaR6r5vPOUBVMjtYIWC3gviUgmSLV3B9jIB6
4+aoiP745JTLg2RtEn+pAjvUPsxweK0zL2K3oCvwbIN+HiumTxyvraBbZKzZcXjUDK2eNkiewKPv
Vx9VJ/CbuhLGtoB1jagJqRVYi2Fd3QDaZ0XZmzP0NXb1zTOxhrlSkJkSZpGO0lK0J3NTF63oPYdb
bWjfIXHMiSvpg7mj7qudqg031iy+qtLB8AY1AQ+tlDd4I4elOXVXwDy5vqIdR5u0E2/9N8WZBtuv
rpfKGFudkH0+xzUENRFG5rgzh5opIAIKUobg4zrxDozhW6Tv9RvUi+bRgwiYsRl7Ill61ShuxBYR
8rugDFRDeWvsB36LVqE7AfkINUkxv+MENCI+n7N5nIPsfcYSXD0Mn4KsJOyLKH/OtL5lQcvn7FA1
M8U90ZkFspxFGmwoZHS0uQLgJsyvvyx5Ff2l0N7JK6Iqeb9ekRZB3cBYo+y00xhKVPdz7VzSeEko
HerppdqYfMVxTtab9BzsVWGFNMtsBq+PiDjxngfpO2+J76pTQkDz1ggnYk0b9eGJNPRCaz9ZlIKw
lxPUD2Ob0qk0DYsTb9Icag4AgWz+Hu3waasspdtZgFOTckHGSO9688RuR4Gd9tTqCV4DX8DMvh2T
2eCR7j3kPwYRjGl7viIyoWKgPpd9inrGCc+fWxtv4Upgpj0YMDSf2xS9IUpFNqPimsZIwBq9XqhT
Q8iurulHiPkRwY16OHs/JzRZznoxtTgdvLlS8vmLGs+tWOi8ENTFgfX8s5MPoFcAMBowoSeZdsjH
TMq+jhoY5C1ERafPau27oiP0HokJA+xxgy99Dp8Uo6QLyUZ7ZwsuqOA+nijgspmFrbPek9X2tIva
B2e6wfQ08YeBCMD9+5YwXmcj0mU5NKwg75MTn9+pgKIYP+K5PzlHKFUDERaMyiAcWZM1YMMdSpxS
wxIukYMHvxg4azbBo9tgOn5R6FXXj6JooxI9cpCo/g/oOzCCGVv0iG+asThrrjPaM3ghrry3O9V7
qH0UTXPoS1ewWxMAi2c2WMUzwYu7jX7soFK8F7BPqiS7dQz28SsftoIBIdO2AGCuxSBk9eLWPPp8
0kBBXlGQmS0ijFL0sGewf7e3zFutBbLDFpN1zO+e7wz2DXvKpV+vcz8HSGMIsjFmcLFpzAr7ZefH
WydxfB3VAnIF1UgeOIN0OuxCCSVvdcRSyDFfD7HnG/5A8f0aeQVl33ULULPjP28hn43xD+UcIrCL
QpMFUgxFBPvu9BxYC5bVIs2iZnxsRuiNukfX20Xduyi6is1VbaI+TqTZMPmLtlNE7mVBkASA7cz6
MTN6jawuJ0FvA4UvmxY2aqgnps+w6aECCtAHX7aYlzmyO1vLRCoE0LsP2CGFwIecDU4KplH1hVdw
y4o90pXBIij7fw7yXAcjSgsJ6j8FpUQfY0Oe0rXC+2AgIWekbmA7UTJAZzxB660s1iZ38uhNe1fF
q0eaYXcqha4k67+EA9wgSeRPRWcktD4E/6VGDU5z56JyR4zaFEFA4bXXJEDlJH7SUPldbBv7wUx/
246ASH+/Sy4r3xx1B2QnYLhOilomaRnWK09IYmi1AOTLcG+qNO9hWJS803glR41xSZTy2Sa1PhUb
zycwsJlGX68cxUO5iqOUe2ZoaQHTjZL095T/X50icRH2ILG3kikjXtvGaM2Ab0SUI39xT4aXEF56
imdox8s7nd0un/iriMR54OwgUGQ+ybV96V6RKOOP0Q0m7nIlT8iZwKZv/y2j2ybdIv3g8DYzlXxk
ze3WX12eazFkSAHa7e9TutBeHE/NcQGO4TI2PUu4vbL0dIgZCDIg69wk2aOx6zlK8NvrxPj2wiv9
L1Ms8/PncpafOYDfQ7dViiy3lWaYTK1js9X38/O2MlCrtXVHV6YOYzibGVcOxr4G5cgqibfB+UNn
03bm2bgXWuJ9QIHZUtlm4QVSMzB4G5yVeB+nB+IiVlQi69H1sgcO8lCMFPLypjf14jZgZlmsDopC
7wzue5/Rcxgb5iHmbTJ0Sf+UH2ht0V6BDC9us5GXcilsxxFxghy+pidQhRzwuuTzr/05XQOBMr2o
VWu9yBRfN8KIzghEdk9s/hTcVwcqlkZCdSu0rIbcD9EISsCajIQ6JVlDN3btrgtjnp3P+6mwWiHX
e2Z7nXCOVDKSCGz3WmMvovYxTPu7Hpn4PA3Ku6vImhPrHxXT6xawQY4mDhRBo8AYVsVimul3BdKt
+sAjtZQRqAweFFH1gInRVmOkad3q9KVTyhpdo4LF4Y9HpZYSbDoiUffpkh/D4y/B9w5CcBUKb0S7
8/EnfOaA+b660KZx9twUX2Xc9++3SeoZdcWfG7cntsmJBWD31mZkVt0HX4ZDPaneYXkWyRTF814z
tFnEy6SnyNa3AkK/97v8/GkmDgdSOaE+RwZgl5lOELm9QZG/zL4TzuRlXNMoM3dIMrXgYI4Gub3M
nEsqEGf1/0JJbbRwBVxJIw41YQCIihfiwID6LjesgYyudtcnrbJtbxT8p9j39lU83ftNl1OrKCrq
3HwQIJCCuWgyNjkjkw1XOM+mYWEZpfHsnGF5ZtEGL5uZsd+AiR9uYsbme/RwYeJbTm0ujUpZdMlU
pOR34r8ZAYnXZdvhODYP5/T+GmPjA9YGGQ2d4kzxuv48FBDBN7vp584ZWsIgeAeXuMbRfQakWIW7
QCMs3RwqEj6ZBpyi05I3TS0eeBtXw78ra9lhE+6IaL/qbncwExlDfOPMB6ehLHocYdtUibvJghnQ
PzNS3Z4xA6HpZMZV28yb5CHjySl38p5oKJVeRzGpLtc2ywUsynAOXppcMU0JooyRGTluAQlNP+ms
M80VSna2BbpfboLwhtqdbCAuTzN+SjLla28GIclxbBRPZ0A2T+8fPksQkvOjJmS4C7wUfeOfT0m/
sUotRF7IW11vylO+HQUT9KxBQHyumo466vym/q8cjREHDJk1vpiM2jJanmA7OjqMX2UJMLExzwpw
/aE7g9e/NYfmH9NKc275ilxn/c+asB+i+/JMZIM3F+hqOwzw4KQq94TWVZsPj69QoCcW35AO3gHi
i03kA0L5h0Me2kGd/Ed/1IzBxwVa34jTkAx/XS8G+qTiw/pnrp1JFiybp1mmhBeo2VHefS4ujo2j
yGDSjf0+roEl3d1zhZqlrPqmHZakzdvOaGki8bvvEMFiA324Z38h0QmT7lR2pO1vWY+pUFEO2u+O
iFVLHq3Uqhfw0tX28w9hKgxpjX2Q/yffn3p0nLS/vckZcmWnpxPyaBfx2YQbGW2l1H341rczx916
Mc5QiSCdc9BbtDkIg9rynZ0HvQzw5WpiBCd4uDvUUZmJZvV6apEZZ1EgjaIrIqPFa6UVdXUWOJ34
jXV042AQbcPujIV9PJvH+EJZNPEc1pZLVa8RLhX9lFbh5dX8AjQAJOzSUlXnqrFGGLFI0RiCvZTz
LFNSC0d7I4M+hFYMhRl0rHlP5NjbT7vRfL0y13WdqUbAhE3NhG3vTVM+K10Ue6wnB6Cx9VNzUVp+
0PHi3npSv3z1d0X14T4O4H2OLos+4i1IqfJbmYzbfKbB2WFqj4GW5zCDV3Ot6j2oIWxVXhb8jfxv
4FjbGcn4iDG1lJ4H+YOoHaEN2AJuFk2KFIcEd1A3S0N4Tqc0GPfprZ+ln9SICYN7ysbn71/tC29h
rT/XjQGQqAxOzTUPt5zB+dvu3vClMCMP4uDZB56e10Km2pe22dnntA6EBUShkJd4aBH5N/PdlYle
BSjOABBamFtPWJW+UovViPjavDhENujZw7n4wWGqilhmiDIdSbHT/DZvvqOHM5mry85/fplQ+eGT
0/Axput0UnXQlzKzHUXbqQiUGLpbL6WZTyMJH2PIIOXmecBqgCdM/zUwl2loatd8aXgOJMnOtEuM
ousFnHqNEHQngeEzoiXevXRSr8O2yELmyPn5wxb9UVi9rZ8vQle1HU3HMGKADKq5plvMjZgXlOpZ
r6crS241uYXLIZbTHWJw4MCyr8krU3n+lFz+pshY4XOMCFlLpBjHhcRXT6UtdrOv96Y/FFJUeKoP
0KxuzjOmj+egZhCA8BZUV6GiEef3W7IW6DO/OJHzJ9qBSmR9XRqiR9CrGOTLBEygZLAEpJ07mR4h
/oEANGRORHZMnro4kh9p5CqtCBGHitVn+576zqDV5erL5u1G1W5kusZ1bRcMwTf53ebB9Wjlo6mz
KhTh98eAs4b8vWPoFY5VuCp/wjqWGq5uzR40mcN+f76zKB0N/svKDqyDXEEztoww9QuUANY4ytI1
hcnQLE1nSk15LgqEimQmlomxUF9WsCVyUHYep5qcAQ/6lUkdXK4GyQS7x7iW0iiLBOya7cl+iwig
u/y9BprDsIehdqEP194/GtWkYMkYpWhFlYHl6O7kn1elKGuVzLIHHtHu/pAXL9TfnW+nSh8S9tGm
A2YtLwIlzJeD6mWLpsq3f02aZAQPMqiz7T41u4w8O0vB2OtR6HW3CWllf3xSrfTKnbLRimhPTx4u
uciGHdH5fE5Lr4dNzIsXZM03lLSVmvqXLcTVAPQRQlIcMOs9VaLaxLd0+qsmimGZ4Z9PCIKfkeSc
ZJKR/NNNlGpVDxdw2ycMkSeKl4XeccTFXL5LRZcaGDrshNi/TjwM0xYcJkjLuZ1cPxww2jrN5lCY
qUp6PSqvRCACEfGNCAkkWMn+/QuFs/6nF4MbzjNoCV9fBB2CbK0er2oUssnH5cpVSukf7sX7N+bv
Bw1PLRumwJwrSp5aL/T6vPUVcXy57sW0zLitET2dAMPgGmXGMLF/GkFzg9fwNbW0ZKhbueO1kWjB
tpymHqWO4L1gs/ecRa7GkoAIYBYIAl4kQC9Zf5uLAohhztKQtajINnYLSOQGiIj3z2ZiA1RVndIC
EWocQl0AHIvjQubDv/zt1X0cp3pMgMxB944M47hswW0KKwPfYsJkl/ghGFKlwXfD7Mcy2Gih+B1H
oGnnXvkNvbyW7qsr/wuPdlz37X0X0AXC5jYCmhAU0xMLpZfuf1QUNUoDDmpBm/KQtguh+BMpm/m/
LD7IaNmlZJRaMnK0qglQDcs34/i7J7yfhD0CMwdYSTjUfOY6Pub8GngIxMTZuNR+UL24jWVGNF3o
Sb6QXmBqoNw/3uJRPrGwtUDpayE5ICJO+BJKhHvupBuRg5s0jtpqGSBDgjWyXKeoufLR8Mlq/Uio
5IvhXaYjxkTdtJqXGkZvpS0xR8KWkvWZ46JsnpJrwp69z9WKtIakx6vZI6CA91fmdv+L1eu++4Z7
6jE41re54FydL8LnTT1GtcdtTYFI+StWi+W4tGZQaux2uSXNj8b11sSIZuzuq6IEhbIquK2ai/Ob
YeFHHIs/ouIdqV1VOi4Wr0l1HKzKACg/Nf6ffSMVIhxx1hb7Qfnp3X9a1lOXek0VEr/s8gW0h7yd
ZvauoZot6LYF1l6gg+tBHeHLjZh2sdTX1TOV/+TCUfiFm1Y/0E9SMNgpLwY3ewcgJxx4daKnsqXS
5R06VYvqskbqjsNVGZtF1TnIJlML0HVt/Cy1LUpbEjVDQ1MR5k7QGBzbKmTMutB2oA1LDQYqnGyt
gt76ba+BcNDNN8wphdgrKgyhbsGzdwqOEzEwwoufTTzsbA86IqMF+uXanvQwBo2SQ5YpO0o6MuXp
JPzDx2en9MP8kHVhKadCe5dtPJBDvk8BmOF23nv8QYQ195PSYQ77jwiI0IaKqIK2hE6NU347Uxww
rTOBNp8ocYa4DGKot4x/TZoFn2SOSjozVIIenMFGK0eZbSCJ1PJg/0HrwrOoBLaO2+uaKkkvwxDD
uV70QPKWGxwjIhwlPQilgU3DX+Aori2SvPI5eOyWB5aOVxQh3ecv4AAEKUIWtR2lsTw0hqLpfhPu
rjN8rsMlh1VD8pVeLv4iReXbklKy69PvGSOwQdA+ZNASsu5tbM6QEn9ZXH5pcxiAW/3VszU1P/8l
JAK+nplei1EP8JuARabmOtxnHsCiyQkzKEmhBKhidSugYDP9Wwh/YJVxXWaCbUJCvjUxT036cBc2
TxJ2iOGaaT/CO7hq+KSxxUVxzolT+S5+z8Ar8wLbSspv5lyrjF0aJ0qykBS3D+BMVF9O1bUpUMqc
h1wnyK0TcJzkz+qgH02k/Ymm/qXRHP9RGs679XUs4huEKUr1z8TiVnOjVsDK7rli84IsccHMXo8n
gyaii/WrJCD7ezjiFRvI5eG+QFrgVyuya5G1dbvl/KxVhh5zaTTpld55tb0hpzT/uX35/0KyMxoA
4DuvRlPUSif3T3a3VQHd8W0Nj7U81AlQrD9ts7aChATQcXrssRg2+z0eR6BqlCoiPL9EUT/tZ3E+
Vbp0FCw14nX+BY/nHmG63mzp/xckSUkHOu43cedtPR9xX2ww1UKGl0MKnRGjjO5Z6/2DOhqovT1W
EXOXYNCW0FeyobjU3R2G3Nm8zySuWSDpLq+YooyKqvZdzKMkZVIxhrj68ROrmxROff7cEA+Nacfk
3MjwGoDZqPnoFgylxvzmv9wl3W3uhHKTC+UqYCjnjhnmRpwu9RgCRvtmwCMa4xOZgInVzsBVKu38
9iC2sSGK+X5jB/Vxpc+h0Hgi2jq4U8Wj+X2soIPKPfZYJjzCMDmMGSaAolMXqIo0qMPubCSZmMUm
x4Avq/fc9h5A0tLBWBFhOk7gbC+7SJfoyjcwcIUX4MwF5ptbnHzY3by1gpMTZirjqvzDZGlckYRD
KDdwq2oj/FTV0TyALjc/d+/Dr+1oDxJ88ZuwpwnF5cGY67rAGsA6T0AhKemHAD/xt3BDYL8VnFbZ
oJzFvv+ZjhqKDmktuef0NZui6Eqkvg+/krlCwQ87goaPgWgA9mzG1N4cL9+c0iSDC5ZOq/0lyP6H
DiyBf+swDkwDNKrfZ7Lc0U2vI/VlNeBRDvKgwfB0ERepnJXhJY66YRh5g2coqrhpqRMPu8XBao8X
Hjm8ocpoN7OmOU+0hGhhdueD2USSfD4iRKj+8sepw63mxw3h5k5uMKX9gqbSkYeFPQguyMoelPo8
AdRDWpcjgYDJp7Uy9BSwqIWOEM/FXMa2TQsYc7yo3EKaDV2TUc8Uu4+TqcfFvi7tZBuGdkOzhCLh
4cdgG/j274GZHxwwCeIExgZ9wstie6yKKkEAyW/+f02DyTL4S0nkSgtyU2fOYFW7OsBowQqFhxnJ
PMr11vy26nAF9mvIWr5egw/8xnjmb0Hl3EJ96QNGYJypDaHYMAQ9PwQwmVvFMSTdeCKPkMIJJLQ7
3hEv3pCwnJ0KRV5MPfWbio81msvx2ao1IRMY9L7HQv4rNUk6rmroKNs522zHkBlkl+SgGfgKWJcz
F72c8wt9Dyc+u210EycvP5k47U5SD/7veyvZQG7zbmezO0eyen1+7OUE0/CA7yPOAQi+KRXgdiEC
ml0wdqApMyPS8wyQ+gt41XKLy3zZtgMqkmziMUuPspJmu3e4cAf1N1RoZ9LXJMqU7G4N8wtmF61d
pL8G+a+bczb8mc/vUf+8CCuuVPzXzh9Pr66QHB6qKVRwStfFElTwHI1FlGnWpER9Uh9rMz6lmWr7
YrHVwqv6Ij/63QZl8esd6QI/8Fk9otrAjM283QLAGp6BK0QyYIN4bBWJMnbH4V8MBD8HKVU4U4E/
LVDP8+P2lDSJW1Gl+WX3+DhZiJfgx5GyKZxRhsyFPdakbNr3Cgt9z42y0QuwQ2lTA8PXkISNb6KJ
EJfEiFhRnsMPNcf3UssGz32bc/GsR9MuI2AGanRz9m6FuSm/QOMm/Oo6c/HBj/leGnzzblrZx6r1
RK8KAh46W1J6GswcADHy+wpI9Xc3a7D1KUUlWp7F/PxSYYXrIzdJLujcgl1S+eenn66T/taXKLQF
3a7xahCy08/56SiISsANJF7BeS/FC7nW6AoJ8coaLVS4/9ME7wB5R/FFDB2+BwU382t02f0MpsQ5
Z3c5GSQJOpoejnD2c46Yal0Iml7FUxG64l5VFuw7Tw9p4LPTKQpGoxvsz8jM/KGYuimtTBHnCc6X
ly+vGNxAHBISr8Bs3CVndejnXjuSN6991znzLCvVuwunxB9TvO+CZOYD1FS6vXORoaZxwpVNfyww
9DLZnvr97uZFc2GvHKps7LNxAIb3tm7T0436yaXsdLJ1wYLZn7YbMHP//SjxVGKiqRzgGPG4bmqd
bZ9s/l6+Lo4HwdeoFpdWYM/8JR6+VBPXqBd2RNf5CE0DdlFwsED9Rhh/uPyv7GAThvJuC0M5UFOJ
oOh04UMIPlSgFGH0vc8YJrqeDrect2OOf908bFwm4+OYu3kd03GtxBpLZ2tsCaElDSGBA4pJ/43I
ZxfG8Z3WBn8u5ZZmcIZ8c4MQ/ycagQurvwLSlfsZEGd5yhYRa8Gps9hhSvVHXXHzfpfwJqZSbNNB
LITo11It4CWB89MhurZ2afyk9cswY/R8Kp7KSPQNawHLKK1O4aMHefva8Ufta883nGjrASRcLTbc
IkOL83DUMzpA7BDxSkp6gmaI5rOwfq+nFZQ2crCRgvX1VoNFxuTn2zDCdBYL5VhD7UYD+z2T93Z4
hVnu+MuwNh7AS5+SvQgFilStON/stvQlfPnkgUH++6FBaHCrveULpxL46DydhAYqZkR9cmsxYJ1T
x7T/J1NYT53EBj5cnlJL7VHmdWtPcmnhYT+TLZy+L6mnDTsVTDMpe9mu8CcL8hWxg6GIAkiFFbtY
0sC2vWfeU9kVm2R/j2QNNxU1hrGf41krh9mzFUD6GrpS4+3noEhYSBTtLYS0CwiSAX2N+saHziOw
et1Yxg7yBTlxpEpMHRimY/sXYtCg3qRf+nh18z1NFLPg29XgUDn+IJaF/Gxv0yRRewikNLJ0rhnu
UBJznpxuWMmljXTPXYMWmnaJ0kMsQDNC0495zZM95JRPRbA/Rj1mv6EqRZQkMcMEMMaam7E4Xm2S
QxzOLN541K3lua/t3yyuYcGjrTYEHxEqgwO17aPigrkB1ng5T7bDvqvb59BbQea9eAd37fw825X8
MEaWYp+VQVxDJB1rcfp1YRkVUiOZ4dG3gHGUj88suRePcx98XPmnn8qwfzqGXbJw8rBKkfoUe3M/
UV92UBgRHfCE4ZkFm89AZCzUHqg3TzexbwyNxKvDhRnAHWEw9Yqsf9Quv4SH3RRPZkAIxGFzFr3j
ymQqWvO1pHGHENIzIKV3DwBkvCynKi/99YoJAd4zOBNB6/4Gck3QmH2rvdkwo6/4cy7uXQ74A8QY
LtxEBysa03gXgb0zWY0cameNfQFcmEqEfBsQJoIkkb/19nYqDReLjjlShgEyeDpwuwOA4TVtHPzq
9qepQP1z3ASgC30H4aQgx5EadKS3170GqjX6269aplivKse9kXhMiI2HNKJ7kNOO2Xh/IIxpyXYf
dIlm1zMMGJ7JJ9fh+2DPeq7280jXFf4rG4My5rtTiEBXM3rioGkEWbc/CV5Jt/xMc+oeFWfrxdWq
7p/pjw1UaUrLzcuLpiypYIWFaZMfEcLvNUzmeAtcMoaYNEyF3nM7vPycWRUqEdSlHD0oiTN8XbKI
RuwoSBYMG/93pbS4adfNJPf5aXkguZXogep0nqjxMcnX0aNmy9k5aEac2Ewb0v6jgWDj+Vd1Lgy+
vt7NKc6tx/a52UKv9rBFkd+7z03Y7o0IJsLjcyFAZr1DFtdtGLiGzrAr7W3y7pI9ubvnEW6VKks2
+owHy+yFGUS7uhSXsKWZb3CDXUKnpdrNTyAuzJ5mDPbeC20XmaCJLPdQ7Oy8YrmfmqHHS3nkwWo1
sQ4qjkzOeXdk9LpMn2+i+dFTmPJiyk8c69cY1VPeRCM9dibig6J6M/Fy7Vgf136Min2vCBdwmhbc
V4E3VJ4QGVwpZgCcDaZ+CUOckJ/6Y2az1bkp4sPVWyu53ZV4ITwdqkfG71uW6bgSmQa002ww8jOX
c+H+bD/iGrJcS8KTZS6u7XqHdUSBrmZyVJaOLkyQ12OVj0H9hN7MszLIbZY5AGXv2Kb17/f5hV1G
znPd7kcHgQnJCc7FPbEEzPgLaMWyzLMuRFCa8vKs5VnzabzQEWLvNXaKvB1x4CjNJKYlRZjYxY2o
t6pnn6ScpsNuMkTR5+f4nMbMvpZel95HR4KgfChRDNOuuzKkKn5Q6c9qIQbTmWpEtIFiA5EK8bCi
MJyGpBs45bSAM7kDPwj8a9yKuNVPhrVFEclXzcz8Mjj+zEv+QkC6NHAWGK4a9z5YbCQunE+4eI4c
2Fux9W/FHOLRRwdoXkVL7KZ/FmT9cH1ePlsmHbUmLsjJvHAIu4f+dxndu3X5QSr4xYnneQppkhil
YM6VgC8qj6/J3Vt0KD+I+B3xRoewGQvkUo+rPtH3KR7oJzM7P41+e4pshx9gYTAknDz47G4HXZoG
BF7yHLomqWnWGaD3kMaox0glh/UJzAPnqXMWCo63GpbLOOzbCh3tWMb72xdGpbDqPsY3rAQYewVM
Ua7WjisuQ/SGNvrW+zvEtUOqtpWMaK3ZAxVll8WVadUc43RSAs7jpMkNNhfOXtfWskIG3/KfwhV8
j8s25Q/SY8cMIw8F1kJXa4XpizQYuhrKF0qo9AdNOqbxlBQx7GReS2lCp9s765VRG12G0fSHsCQo
/nkM8BFBlmmHUT8ODxC3GMo/IT23qX7bMT6GRhHLjCDkfAmtZAm9JpxyI4bQ4CY4bm8NxwW6Qfd8
VqH1QT/msYl0a3h8wl+OXC8GlCA8cZlqpY5HN7ak5oz0xvKP2yedJvywmvt2AbI+JU9BQj6ym0cH
EAV+Y7CJ0nIt3MrKSQuD4OTWuojNihRbB3zj+bpv1m33KdJTg9Km8aYCvLAnkCe0cBD8EavhcvVe
kCqV/acTgC9tGjBEkBw84J6PkQpI4axmffqVWFecSY6TAGjVZMt3twT/zGTPMsJjwN3HwFqH6F5c
wqDM05tJ72oHpgKcmYlVZ0hHtPUsIHgzlYGKCPqmeSQ3JZpjmBamJ+8vfr4h04DnfRO5R7Ixv2xy
IFNq0/PQLx1b/5GXY+qjN4EnKGUeLIwyknTvjTeXpnDvwplYvrgctbE7PZmSKeNz/h4tkC0tplgd
NyEHP+9fNKXSDxOI8zrYH3f7x6EBXJGrGtpOzMVX9DXt+eZL4EwqUUfx0SzWW9MVjt3ij2+SwZMS
57itE+AROmhtnbXtuAbOshkBT5Asi6gL9yABAkNOu9yoiF595BdcJnXEM8H+791QLbxGOhPnqzx5
WRcz9WDl1IlnDNGg39Vkl5Dg5+thK9ilzWwqvwYwBY0S5raMtm0Q+TU6nx7iPDkTFwxgPt8jPe0S
BVrilBFrcLGVDqoXGku5bF3SsMlDFSUdXg33c2R94FdyE/Xk0j25ye2X0w2DtobUzliXvNChM2KM
9r1FH9Fr+phkeFWeUPGvckXsHy01OmWrWKGXZYafqSAfIeOt4iDuNyXb7oZoN6lhxbA6C2P9F8k9
ynBdavjoyF1MBEF/c9yoRfJSrZUTYsGyomNgbeI6P4Qm+MOLV+1TYZ34vkxTtAQ6xjWoTGHXrO+E
KBTFlVGmMiRMYLFVTf3NHFexYFDMiRIOTJzlniO+52vZgWOrV7Z6ZuCNxpcZr9VMThALLM1s3cL3
5ZT49yj/WcrSaMVx6bDufpZmcVNq3sIVmi4iyvby6HbFkzU4cMQ+9vz/A9s/XzP715cT/Yah3hd7
RbApFXeUhkhCuhwuRWk9gKc7Oel/IjGDhoYwBrPCfWJEtF2wnSiXp+/6U+HZ3WA2WE4hHPBJ7ucN
FSVFj7eM0KbWwEldaLcJW4bPRfa79fqURnQcEdRLdIi/mzPBq6OEgHM3aDF9NNgp9ov8SnpIMGtc
a+NjRjEQnMj5w0Cx/FbJSzXh+1dGBkACfK+lDkR556evNG1mv46TU1iflQh/IoGj6M25eLRoQPnk
GXdOK4gaHFpVv6BTt/TqHkB/Y5/hxPh0OIMOcbMdMmGue0SHW5aM+D61z+EuR6W1hzL2E4I//6JK
sZYUTXW0SUXYMT46XKwsiu3/pFrXQvaH1xDLBECV9FGfYDcjb6ZGRU3o4v8fmH/7ioLJmukCEDit
OW7W0ZUPHmbeP94sNpUfb0Xi5ANrnjGKvx1cL3XFwPWdAEhNiPKYtsfn89twaTLi8vVN9//bm+DD
xs26Q0ljP7s0j4Cg57N8Xgzox0MtKAJtzcTPMr2OPZWPTWKdRNpJGZtYRorybZKYFOI4g2Dw4mRg
41DopzzVKtLhTS95jahAuQBgsqZDuV4hERvuEIIXCapbLOjWG57y1ZvD36OuX7Nk56eF7pUjjY0T
lNFKqbux5Dny6x2lHN3gouKiSIFBMa7yUyFUaQq/xhmFv0lgMPSZanucktDnv5eWCRxRIHZ24ptG
Z4PTn4LNukd5Jb3duwUDUrVmDEFb2x2TuPQNTy3fRx++BxG9spXCpK3D6Jnefi6J9nHahvJyTSJ8
6UOHdyfQrWUETZgOIg6V0k1A5d1NjQfbWkFwJpnNxnMOTXe1b+sh95Ya4uzr2R+LAoVeRcqNzVz1
fOqtJqs8YVcQPE84GDPsSAoHR/cr8An3X9JUnqXoKJz7fkuaEaDr4YPxPJmKxZJn7PS3/BJB+z1f
AyEZLCP1oqg8QfZhO5lTVB5UbCJg28Eg94tUyvhdVYNsx/HEgSWO6n4wqKD+Eb3I59L5SWFLh3do
1KCEtjRxYNH1NVxpuPo8GjRBhJQFTz8PFgUyV1OjSkKKGKqdJhh3eWbvkqujsFgLGGU1jXOnH4Jt
MakbhOvNwbZPurOiGFIPC7BcH45LpX0EFeFxHbJYBSLSyVa+/EDed6aUbVrWLfm1lTA+oQ1qbxgG
Kt9DL/32PyKMFNau+MdAbG5NXH9LpFsiovsLBmYFe2RQilVGiBX+bxMq2FNMg8Bu4eczjXBlhSF0
mz+2D/8HOHX+x+GSXQnOb+BJLiHBNV8PGVeFXYS9IqIP8vzN2+eERV2FW8t/wtLefB6yekOigYtc
n7/osf++ALwdOkW1HbSQai73MgR0ZCiIXwZQC7JdIHs3QMCgnM5C5iuVVs+XqD1tjrU1vWgbtnrJ
1NmRR6PXe3+NCUCrrTzF1winxisncJ5FVjHtJf4Ghg4+lMu/UA9589KzQjXfpFNd9HbcPpW8oH+A
yMDyaou/MgGC+yV55KyNjzbd64CI+RzdaADGjtZQrLuj+SK05XP6dwTCv8mIxeFzQZpz4kQ1yvwn
TTJYXqJSS+0EOIHbyoGnmvc0a2ik9kIJzawaEPUZ9DmrBuryFNplCp4M2CKgbUlPC7gaoB+ycB27
BUusKhRoa9FHwBgLylwjc7nBy390xkcUDCVCmIJll4H1PfvjLwrxAU4gky3OHj7bqv1LJcEBDdfq
O7Q0JxScIC6WKLorWoasCywfATJ9edQR8PbR5CBwWxryXyquVlMEsGQANC2+SD3b0TvVpOlZF/ZI
Iu/vzWO7MAEbxQUCVkV97+Nt1cCUwcw0DKuzTBBhVOdDfy20iZ+/+H6HNJXG/RVkqRBHynfhDdBi
T2GCnE5B7Z8/2O0Cjhvt/5KYa4egX9dcRyLcZIOrGOQrvJ5leE7bKJr96xG7dLx9W15cffeiEczM
UHa2tIrwLXWLbrhky1eb+fUqqvsKRdcsZZNcJ8VUzklNPl88yNZJb6LHGU2nowuxnO3PlW8gbQLH
oBg1RV1+VEmFhJnJSDWvHqPJ6fyeuNdYQNPx9IRNQBHGAtMBd/6l6Bz5G3Z51gw/0WOprYoWBsLk
HMSDx12ZU5MCBQFdvtCh3ZPAjdF8rqMPPgCXIVSd7MO8CzpVMXIW/3+RoW678AaQjrBbBPac2G2B
LgUXn49vpru57DaKZR8tWTP9a+fjutzzA9Ac1LhwHUhztO8dz9cP6uMFmg+OKiRRBPKOh6CG8bSk
zRBjyVWq1aa8E4XY4FlavRubabOxeM1OEUsQQCsZuNMf5++WSYKN1ppxmqtUQpIn0+cke9XH6idQ
jjRyARjNUbY8AbhmbbDYANvWPS2ZVw5zxCOepMrjdL/pYA3mYFmCKK4n5XkfGf3l0lrfU1PqUfHD
c7NRLi2I7CWLd5hJyg0U5pAi/Pj1mFXrtPmFVteE49u/gEiyPFaf7ZhfpbmNxix0IXnKaK2ll+5Q
Ay7mQR4ohoeZi+fs8DYQ/w/VFZ42OhIXFPR+9GZD+m+pTjccYF8j2pkEtU1kOyu6I6D4ZSX9qQM1
e/33Czl8XB7C6KnWjrfrWxhR+c8kCItbiImCDgcVyEsMq+gH7fZ6eIWCpKT5oSBlnpQpRyqupTBB
RLXLPUiub8z/m4bk+xKrZ/c7g+4nMYGKh626ruaO/O919zRsS1Tmj7ZmC30XlH6YyQc0cSeJRHrC
tKHURBKAjk0SzFPRdIWm7l5o6p8IxcsH3xW4yL8lKipoujW+P6cBUYPFjvRGCoWwl1eWKx7mqL1U
UrSgdW5R/1GSFDBOcGPF8HVBGPkXuIagCSiSc2UEYRKfjyy+Y15oMAN+WxRqgaZGZPOhAZdOlWfp
b9sW2U3MLdYk9u78ro/5kiT+05kSFDoXl+kIncwE0KjL9gHLMdV5OpbnJEl8ytU2AroWoJ6V9NNl
b/4u7cuBQdZGf++d3tRT19YAbMSw/bgY9JWu6Gv/21127gPuLWMT5rkM+i3X0wsUCqPH3RdQx4Hq
hHiiX4WB6EzdO/2m5hE9ayqGdzL4R22S5sLQVTP6xupSQKVn6po9OdFWsQ9XTJvvRvrqk8tK2bvR
FM3qQwN7MIRrP2P4/L6Kx2KfYwsHo+WeIiNDYtPV6RE9+titLizAVsLulj4IbrbFW+how8S9KD6+
OnqP++P6ue5M/RfaddNd8Wo0Bi8VmKmxsIk9F0Kx9Mo8zyRoaTvCoN4TIE/FcW/MdKMPwZhErdOp
EBS42EfTtVTUimWBvDxI6xtT6DWv8tMnYi6o3TRqUCG0zzDc7KJlZNKSDrWzVfOYcgoJthO6Gea0
3jHYV3bBhlpTJ6HhqeaWopY8uEkJ0CR9lwjup0bVH0DlRjlUJG1fRKp6DuvVAqtWxWNAXI9JBHJ8
QNN0EOIAw99TpUYrCP7vPjUe6Oy3JXl0aVl1by1amyNzs8Z7uoSXhnaph8KzSuiMyv0KJmwZpE8m
S5irsDS2OMawJi5H0y3jLuziR6VaFqKe8BaLvu3XFi9OPMHmn402NLZ1k00fjY3Fkf3+YgYdBtkp
rTxXxuIV3Da3ujH6qHybhGUhK3kvKkN37KUOaGszUer2Z7ISxM8mEUQZCbpTQIoZVl2cA7NGFS4v
HWWMHwTRG15NwvbGPcLYT+yGXxsSiBApGl9l8T1oQOU2pmtDVVSarO4n0EBuuw5hYDMw/XID9tbU
ak7XWO2BfbYXn9BcsWm4KnyTN/hFA1oPnPN1Ya2ADII49O04Fumlj19YSmYrlzgLr63Btg6uVdZq
Xzi8+Cf8K3MfLWcwmFQLqxn57aQcMIjt7mPCcuq7cNmI+RnfmqtEbFMGNsZ6QwUOofqe5RfpW6Pd
gWsk/GtrB27zcf2ifO8LcUzPSOlvVOCojIs1GzNYEo4OFaf+KAC1m92HfrR2cLrS3LKkrptnj4Ym
fB5beOb3rM2Q0BndTRyEPtWsf7REIbIrlXh4ft3tmPCEeGIUJqYTDLG6X8+kMza5vl2F6vYdHh8v
D7AHyUwT7B7S97OEDxbw8SHX2CQrWxdlHv5ItnPbdJqK0XpiYnJMejF4oWtewyBUN3mMq3pyiR7k
/zWqPqNT87ia+wu5fjUdKPD4rzROcpR1ao1/dAl6JfPuHJlYcPJprqlj0vSGKFTPK+N7fCnI1bWq
9mvBiw4+p+ysS1k4Ls1ad9afBGmHYaFLxBX75VVEa1afLeY6NPbv+469CQMX9mg7kY3tr9D3i8/B
z5IGJB+F+GunGppBWAOql4PMxjoQfVJBZo9CrUoiVL9/nhUsRjJclHtdr7WxAQ/icYvKUzW8tpdn
dk+YQRTdnSkqt7wSVgmH+zso42FXir1OB08U1uMxO9Nd5GChrdlPMVHD12eiSxia9wF9v7toIfUK
ugzmgcfh6CmOC/UaUQYuUGfNkLaori9JntESM1uYGGGu+aPz6soEEot7n33RFYhxWbMskTWoTbXk
Z8u9oEyxe4KuQGsI0q4F7er9CZqs6aAcW7A1Sssm7T0fr6xwXNi0BP3PYvG22BAj/WW4SzvQLyvw
1HFWQQPaO5/yDgtxJFXWaAJSXLCT+G3LohqLn7itAMezGjYTalnT6RTF5bxpzOFFghlxqzKk8hOU
ziO2rzRHdOGVHYiiScp5E55DwjYpjEqdbBBBZJMPCLKFZB8IOEkMW6UO8EHbLnXKBxdxQVOr2r0+
nAJdeLTaOXAzlENr3FIAxozvYZwW5yufzlt2WzWYzuxKmkjSVzCyxxwCkbvXwDqDPHxB5LxZFGNm
bpXdxChVCWXsSESyGKRwsHz45IYzRZigVpFiG04VX+s6O6Vmsn42IkhtajwUo2y/YPJLswRH35Ld
fC7MHBBPosg+wCShkSV6g4Q8/F5TgdUr4yo1ndybWEl7ctNuAXhtIZ9zYQ1rjDy1xYGgTdObSEFc
tZv+/qdvDaAyxEjcY40wMGXVzCOK9P0Kgckhmfc7IBgI+MSXFPDQbBRYlA8Ox2FQtbJf/Fm/1GFT
c/3mNGh5IwIG8TusAO8XTFNW7izMvAi36YO1kbK5A0recPvd0TEFFLdk7Yzib+HmnEdDgPUd9MF8
VUYmdz+x3UwPAHlzvSVYXPG9pQwpspW1Gnoc1QJnB4p6qqc3sgMQ+O8lQJtUy2tpVRusj7tOPNQQ
lYAi/xEfIvHPz7kgMZu4WeO0ULw/853S4LfjAxekVT1HBv2t4uXljGciwHGySPo8G4+vU3SQ4W5T
XCUvxjB7NDQXF7lCIXuLD/34MCSAkzEBitI+IkG+CQaOd7+curAr8XAUSgm2eiEkJ8FX2fE9z6v3
ToE7OBM+qNtc4vYAUxE+qJ32lNKoi2/tzgwE0Tu3TbL6PskcvPZJYYMtqIuhrlqddIPNpIGDBVjZ
E8X+xAN9dEzhQ1/ns4xINiH1hRcaoiLpwqT1DBouT4YJG9lHNscwH89811GVdcsfyhR8hRIyghW8
NQnAVjkxTMfYlrFhTpDMOi1p8TevCE8nCAStdZoJd+PI7YqoftaDOKmQY7fQGPgwfg855zltXpYy
P5ogrjFH3s9NXraKiw4T6H+DT6CK29cLL1/xI3sjKVdMgwIgsvQfjK4Yg+ewDbWHNBOL9MhnVsGa
Et9Rq8BdeYBcxTqxT91HA4DBMk4pTJPY53kNhvQNwSu33Oop3CgkObtsxdn0U5p+47ZF37jfiIM5
gBMMgMZdAw0N5sNOxZKqIj4ep7GJtcU71PAI9YMqmS5V6oqhmntSy9ATImOHIHlRDBqe4GegljFn
UN5ztHBEbCYoXUcs/aKgaysWK1qwahOt/xdOMPq10EE7eYIPu8Tp6zob/shlMJAI3DGGKcgSKlxb
kR3KnoDaFB6Ac0ZDFuLgjtg30FbjfOMS2nBdZ15LBiaAKDpx3GyIWfdo3NKAikTUAIbPkOAfI83G
ZVhwA8N8mnjG5nn1YyQbSLXWptp5RTs0TJFFRKQoZ4L0JgRTFl7n8XYX+TR26bvq+NECJ+7wHrn9
J/G12qmk95LBye9O/cxbXUE8idyYELUWil3VSZLse5kt4fBOwVr3Rrf2OQnhr5ZrTJTZND0cU6U2
v3SrSOYkPY0Uy7hghGbbyCa0B2l//cJ3nrTklcEcL2PzSbmq5o0f2LYj0RBa9rG261uu3KANZxJH
DSnYZCV8t/ziqLozb7O+r8cy9y3TppW34pImmDXziNoyWmDxXjrUC9VGNQtokzqYWvfZ8CpvENuG
UQpU2+L2HPJGkTOjb2xtYsV+1664wrx9qh9gm52wSEbbCgv5r1tdmG8IKGUNPcORtbYYMtMnttx3
outb6Zr7E3ceaoKYWk8IVLLq+MM3zdnu1TsKQPMU8d3m/jlgubvIlzMBbq6AdrZTeDFcwjGFBlng
yjd+/lUtL7e5vo6Je9D6bH/uMeoQFQgSLMvKMSE7Sk3e2t8Zi7r/dRO9F8E6oEzEesw1CD7LCMg2
jQUriuxSwy7cdZRXVQnUFynHmlh0IOhSbYrhgcgS/4EGCqlJCZOqDWVV137FX0P5TTxFLarIZYFF
wgecpKP4gLKWMC+1umKfhBESZ53TcsFNwIctQYhDEgDxN2fdnuz9n+ErNgizg2YkViRnei9vfQBz
eTbokNcEnxA4eJ5JsPCVIWQ/jnYh2hAFCC+ZI7LAHuaNo2JCTkQL4hiAQlPC9i+nzAmLvWmfwt/p
/E1qL8E1zkmWKNPGbPsanB3HigTodaG5jaa0GZIeOzyPaJIRTElL7+8GLthwCeGgIq+aUzAFkalN
QyFLHOxzExz4AZJRjIQ/MjZ2di7j24VO+fTMMnvc8goYorGF4kyWqqKigpah3gnBPjuLzKoMysTG
TPHkgZWF+x7nPk1KhqgVjnHLBeSLFC3kIDCjGORDUCWLtGyecYD104kBju0sOj0vFmqRa+Pk+N1c
Bj9Hu5NcRr/kb4vzKcMQCM8uFd8OMLVnQMieJqSv3+rrOKygWxMtCeOqexH1WLkJfqHVXGD3fcCH
090TyofFS+Ge2EhfAcxg6QVIVJkzQ3uL/n4Tc4cWpIXU3ldBMbHXnYxtFQ0iPU+zKuOh/Zb+yTSJ
1durOwvWjBIAZ4baTOQhKFouZEhpdnCw1H3w/zsBnxU1taDRCzVkvyv51n1AP8U0Vmd6BsOJQ7to
08eDoVXjCdu+Lnuquk2iIjvB36BJupQxqD6GmcIlhCWLZX8g0DZKikBoXvgt+gqliBNrXMZYnDWP
qIn4KlgYUC/p1KoezOWe5vciwLDBBNL1OEnkLn0IdBzbQ4C9F8SpiKwN3TgX0odLTp4PCg/XICiu
LnfnYaVLDLXSwE1q9s7/oRcCwCkeuQCA+jIwsj8mEw8KlC0+ecSBqG0JkQhcJ0fgJ5+oVzUCe5MH
gd147uozAZkYugBmM+3+bAx6r33bm2EwBhpa0SxvavJLq/Gkrr1ljfZnXG2xeOGZVjhdbEfqEoA3
14KKjHfyXHmzgxhB/uKD7Qb5ilPZfFtNT7a7y+tXrSZvdczZlaefXPbXu4/7mRIXi6AfcuqDst2/
fASOMeaxZYs9DliFf/eY+gVpI6/P6WJeaNoKDKJPNIyhkb7+344nKA3tN+K6UjSZoujLHQPN/Kzs
jgE1EazKK6+pxEHLxWg3pJa1jDLmDxnY9VIjx3BotVRdoDfF1VM/CroXzGGTaFqgH0C92QAKlBN1
K3tGeLtf89rjoFVZYTgRvC+pIDjiIzYclBtu03Kc4OrPLP9eP8leLzw6NBSpi66EWqfe7C5KA7c/
SxhOwMjdadVljgQnmVtgWpG5esme1kRxh9vJYVu4ocbBuCie5g8raUQ77cxUDDQG7vJjEz5hGc3m
bvH9ed/V8cjMOQQk0DiSzcVeRB4aKopnauwalcaLX9H93pVGfQaNnkGO7SB5btVtHLtM48NtxNv0
MY7tnVRMZAFjB+CdseIhAvG20TKr8VrJlofOhnrQqjW4iFiblDnvdIbeei4MWNgedyFg/HwL4PK4
Pf6gl5gmT2Ts7vU5ntlJ4zymJn5lTg/GMeV+GB5zlESA3SiOPc+a0sDsY6cMFbth85MUU7xouPUB
k821qzk4gTeJdIsufRWpsXesg3Fk36bGkbEBj69vW+MS+qRWLMyj54B/AZJ7tqPHZ+3bHaq1Qypp
xDNEkt1eVQInDKZr4YDE2SeaLDdbiVt6dydC/xvCznBiHb7hp9XtSdSavdTIMzDwH571sE34W6Cc
R59jgfnukz9eZNWhwC9HRlpXjZKJ95XbcxPXIYr9GzwoUYLha+FmH0wmuO4pNxak5005JzAtNH9y
KeyR6TLKItkhAx6Y30/DJ3tY4xsAudC6BVkcIJOzrBnQRev2UtpM+d/8rHu6pjwlG+TkHzhXQKR3
R+488N5ex6Xhtr0//skAQiMx/B94GhsF83WrEaIGwfzbmtpwXP1LrUYcUqqXyL6SpGign6d7gVBr
rW2RUstobELaIuv7ZtKJZz1l9Zizq2OWK21NBfaOd2c8znFp1oLxvEPAqdh0TJTfQ0JwLOJ+yID4
d6fGNm8QQes69paZvOYArKvwsKh+iJLdtTyhTfo6t6Reuyc5KriPcod2d+VNeYzTlryVTpr36ICa
KCI/rXXOIC6fshqCQfv/LZXRzJPRgNcABs9L0FOm71lvMn+8ExCr2ij1qWBjFi+o7I/gAAJSzC+R
6lWXfhgJfJ/qo8odutZacI7KkVYFYZqucs9T2J5XmpUUwgiM94qir8/X0EWe7dwDJrqwiJp3lj/e
xAzNzTiaP/jjfuQltFZhLihPa6MIfm2PAkTLW+VQViVJYKhx0gaC3hdXybQ41lZsX6UiBHWRs4rR
qh1ZjwresqFsH4fC7jizc9HXMId+qrj88wGtAK1oyc8cKPHVENNhdLHDDYkZMzyLfWQd/7lwZyHR
PABrFP0WLnEV3WY1FM/aqkfJJ2gwLX4HnJOPB+ix7noc/fQ8yjqdbp8d7aKKVxXtxWkDZsI4uEGP
eNZUDUsF8TLwgeZfAJLpu6rO03lZc10Z+L8x2XTHpOHX1tAS1ytgQHx12g2F/3xRzk/t9KMzmwZn
//bUPDPX2O1O7sDQfApbllHjxaHraI7zwsKDH+yERe0RwXzNGa4pzow2jgb6HveTJcUs1P4Dcncb
WRTFVLZMw3cnbYEIE/pdHZCeM5ALOgDxQEpc+EzEf9mV1SxqIaT91Lsv8GucDj2v67DMoNghFW1y
y6cOcVh5L90x/NSTVASniXqj+kqjTVf8ZMU1GcFPd7sWk5ZqcqpOmD5U7PTY6b1R6owNsXxkzGiy
tLTucYfTLQDfon4RArk65YMp9GEkHuVq+ZImM//gmVZ/ig+rm+44qzfo8+0fXebXpUBk8FTxaWrE
2zTaLEenyclABw4oqLgsCmw4hcIVNM5CDarY9TH01V/q5Y+L8SU/8e1YwRmSnIFFCAuoU51RMtnO
s7DjJKkShqIom0FsreT//ra/foPmV7UMgtSmEDXtmv6b7zgKW67biHbtuD7GIVLfjQ1LzngZC1pG
B5nF6aMBhWJipxixou9yTrLIZKuo6f3qe7f+/X8kzeAJv8Vuu45HF093ancS8X5vfeIVICYsHW0s
5GCkJhnPgJVSzbsX6cSSQGR+gTYjD9FsMocdsrEehx1MJzogRbTPO8qQGJsoWvZiHzeM2l/xTsI1
VgnnUgZIxkd9O2b1j8GV5sOT8bL7V/GrJ1NZ6WlF7f2xAgl6AeHYpE87UTWY/1TPW05LM7hkRok9
xrIHKDymXBx2O+Yr2q/a3tr1wTz/elIPRQV+5UpACv75txsqagPFcwG/CuoBXXGeOGvl1TyGsqhQ
22Aapwy+LDIiq5DmAbO87Y3aAl5KHdQwSaNTu9dVoLO6ekxzwCyUG3glCzeiOPymSXtchXbD+11v
0JwND3AXZPEtPgVaSf9JkIEqrCa9wNaJZB0BLbP4kHhYGgbjvamgQxSo0jvGh8jZ6xEwIAVXfGFw
NhkUUEPNUkMeT/Zp6L/x2f8KdNrJzFYaXnDC/R5J1P7DnDw0OMKZXrjSm/yciVWgxjVNFgSLW0hO
bRcTKNxbSJb5yWV/6fOAFnx7+KxOBS0MhRxWcwNTpvHqj6L6MQbMaxlvXzuq1eE/Bhydk6AHhi9u
55dZRddQfGeIHY7Ydr8T66UziSl78y2Ync02HM41oPZEz8ltF/5kVB8zVA8+DqVPPNjkxvTrVYc7
buks64acjIIAiM9dlB52fgcE81FlxENFIGZddoDpiqhvT2+PNBPMSznX8lI9TxvBQunalWq+v4UR
cpUWrnkBVct3tCAW7v7QhAKQ0rE8DMKODiS5nJjfNZ3L8BDdjqRZ52lalN0858fFe1xLGJ3PGXt3
o2+gqsvZXJBa4dsDvPpyF5f5sfCokANxhkS7N+8hYfwqLlkPAuExXj6zfmzlBHhEvjx3b5Ned6ro
L3sNYubJ3AaKNg9SMxehPmmnV1vq53yX8n54jLYRBp7zFWD/xgfMZuJs+TeElgZmjmnDUEG5AP8a
A8wC9W1AAqdaeUK4jccWO9Rf9QU9288IuGFimZQk0bdUM6UiUG3fLAm7e1Ie1E8w6egOtLf1LTC8
Ykobfykd8w+79WEBZsrM5L7e75U8bBnbddgPEvhQmwIJ/QpoHRYdH3iJJtLmquKYdFP+ctBcgeO8
iHzu9NwCmcBC3Vf7M6H2mvJ9N/Z3rtiqENzZpiEcd+YZ457/gIH7UO51pFH2jxKxc8oT5YutkXLB
XeSY4ZV3kx3pRLghRmXQ2Zo+U94JPmKXwlQ8avXCzxz7ThNsiY27ZV8DeFa+Zk/kE1KGZ5hfprU0
uCt/D34VewIvzhY9e1RR9eZ4imV3IRuh5P7oZFNynLc/AWgsbzWGXVAdM22WnMCpKJKYw9PhcDCg
t7yjeI81UvXPbW28JqYNYQmYgwoBtYhgJDI46sRKLPlWwk3NFEg+709aXNIco8HK54LSt8cTK7CS
w/NjxJSC/laswlNAenoSPXGuUxDZnhA8b/lDiaHgcX/qqSamU8udgiYR+6bk4eW6wUANkVSj5Ffl
PXO1ijWnfBgmk0u1GEv4wLsH0ExpsJdAPwSms3WgrX6Swu7uAa/AXGS4lgs8/lfxufmFct41V4ir
Ow/xx/XdE8CCU1IsIfd2hsn8b2g6bJS4usHJdTsw+rgPK69GbFJbNtTarGlS1Px8F4MB3iHvxLjp
vC0FzBaW/H48kAmjxRHCPeglAAHeuFPkgYXkTtl4ZZVFte9K/FRobe3gsJ0b2xxPfdTZeYtSKSny
Qv9XkruGCIT94NjHyHbMFDrhgsjjtD0x7zt0mWRfpf/uKIXrJBa8zHmhsZX8Jc8cp0LPHmHenoHg
UDupEdgl/4mOACaKK99HVzz7gmbV6cBk8iTFE4HmE6c++MOboqqrpQs0Fop84RomrwBKXfKzMAX/
cuGForFHs5GYCTkf3RxCBJ/9qLQrZnI768HCVGE8rWt6QiynBGZ/Wndj3jMtSQmJCa+XSpNXHU5x
zJJkF+f1hznLyYp35oUytGBAlL8AEt2Bh72NuEpFowFX/jg8XeDWRPqPRUnBlAjGL+E6dhQVrCPH
N04LX/w2uMVzCEEFpII5/lOeOcow4+Tjz1Gy9ZdFJ7bSdOBf063DwkRNfeFTzKWNwpcM/TSTafQk
5HwfdYFzpRnXuaaGyApQOZN6thfHuPufDqjkv5Ek3TxbzcnVQM+mTNa+wODEC7NH2LTNdJ/6lTVj
Nj6ykA/TAspK54hLtp8OlJ3+EEYqLupDQxGrM6BZT6FasdSPGzCcq9N1fb++8HRKTxeV4Hc4rAdq
MFmf1dU5G4Cs+t1vbMrJhgNdbqZSzk5g14k4G5SGcjTfT4tIb/LAxuRYNStZyzAX9hL8nWn2PC/i
7Dq2wVwm8Ze9BdX5/9dpGeC6PZ9OtU6liklN3MtAswapS/ednd/97HA+Vo++DmtNN23QdfShe8Wr
y2eIEi7vbSW1ostvWuk0i7NXNojItgyA5RaPTlCHSzYzjnoW4KhIU33oh1LYzPw11XPDQMVUHTUI
L1u3tyJ1SC2BvmzeN6wYl3o+NckBZ4a5ORdg5vZ4QtV4pwi9BWvniFrrinHc3fM37KEc0AGXDYb6
s7A1ZJVEjIkkZ3NjwGqiz6pgN7wX1WXMAWm8pPB+fGrHU+aYCffm3xyIu86m+0vHTG29VvPGhYUZ
udE/3HP8lROYmL6Ry/jlEuHWMMabS8YjNlY9Rd5u5hcL4IJNWqM8DaRTcax5GKHpTQTlrDuIoq4f
QBhNXwmsClvyC7qQCwcjZEBL/5mfNnG9OreT3RMt7H9ii/wwietzORY4TJbsNcJtW+PRSQ+XlSYu
JkKO7VFNrYgByWEBjciWeUwrH19bnb8nypuASZb7K/B6ifJSY9bsl12T8WnAOe2AWA3IcNz1FW21
79SYDl1Xa9v9i/bF42nOTlGJz3qga4lN99z/YWSoTuUDvGczoKlMCNL94fhiIRH1IAIZ15g+ctwj
d2UUm+sVHI0rDoGllYBFvK0IvR7rqldhDYbrGYX4nHM8xuqy2n3AuGOku3XXbYf+X40AYI2y7C26
CY9YlygOGfGRCYiBp+yRm4WWg6wai7ZGcHKSVEeuRHRfD/yOKgEC1y78UAeTHNF0297Roq5a83DA
6UX8DTp8B/OsML9A81eEoTdLF1z2rzUrqrnLMrE9EYcsFT9gNNhUCLA2P9cqPX55FOxFagAwsur/
Uwu8ou8Mep/AIC3rxSfYnZ2ELyzMlicRRn3GoY2oRcNj1+uHVUzrrilkFtRmfE5zryRcn3QFYPSk
WE3TXa2qAkUfoFwUsxBB+ypzdijhOj1NcDudhegV9vTObehYrGcc25ms1Q7egiYGOS565Mii0BkY
3+WZ6d6UQjS9IxZCHy0IoczKPvWMdXSZQpxUo6EWeeUx0aVnI1boA01LVAlFlT3jKlbJn67k1y3S
CPgVQcOiQHNpN1dn8funCgu9c0Kk4vIfK9lfVl6nLDC7H30hBJYRs7rY0VbF2wbXkBMkbbOAeDCZ
MuMXbvLO1rffISURq3EThkqITYvcEhlwvy3VGCVpEYUxLqcohnfQKcV3CXfj2Qktam+QMqP0Q99u
0i5JQFtxdTj5FMvSau/38XjPopCRriIlSq8anq/pnDtT/Bbt7tDqMvI2MuAoLA81WntaIfY0t3IY
CeuokBEVcWjmlmt7JGGfVJUDPABzZet8qX0qaNKF5aoqEqJIA9IGsiARPpCspGOlvnakow2whyLl
J35vdpkZ2MbZLFnlfPuwCzQ0eWypG2pW2wJD9o2/YIEPaJOvHY/WMFajVSLIQ0+fOuFkdFFzRQPo
pvIyBbFrd9J3Rna/QzgVUaghxpIFccyQHahFN6M0oHh6uNgz9h5VZ8Hr7zKc9ejKI3qtQrmU/ez4
mOLp7pv4cP0002huX/AdEyT1FtyxnwGdr3cnZdBSBHh5sV0TMvMmd2pLVXjUbQXw5/d4SopLA16n
QIG2kd5IfC6LqVzVFoIj8cUrP91rVEKkfcsc1+HL4iX2IR4ieyQHGPUHPvfv5vBQDznvD4zyKy+x
Typ6xgyGj1KCCP2D3HXsKJ8l6JaCFvp2hb/K4oPjE27cVdOTAsoIH+Y3f5hDfZnpghq4wQ0wbxWf
XHU9pM9LTqC4KVSsEf5+CD5t3nNJ1z6bV0aJLnTJGJvIUyuCUOu4lbojPSMy4DL2Mw5jsGkK8rNV
gzxdqXlTcJWo8omUQv4OgiJYAyCWDQ/Kl7/5dG4/Cjr21ROkCYH7Yg0Ee1z94nHr+22VG4csZFpF
Jpo7avThXvvLyWfASiZts3YyansMRHxnhno8yDq9M58tsoCPB5iSuMqxKhtIUxioHRlY6T6kRpbW
3SApD7yJeUEbPUXqiFDa+wzS10dynz8VUcMlF76OIsSSG/yzxZOomUMAbkukrIahOXU66Wdm7yAa
YoupnpUQSNuAz1dOXMy4oRQYFaMSBsviEPodoK1aPFBtkILSxsG6lEghWb3QvfsMOce9Rh+0KljJ
7mYsTjnDFCe6i/lyi8zwqieNQCoxh4DL0CvYIRzyphdebbLBuGot0k56Mca4bcifvFHyioNfP7rK
VxFZPdQnQeFOe1BTrjmihIfb7g6BTi2sNTrDZ05eGEavFD3dwSI4CzULQu6qEOnCqp5Z+cOBIfCK
AteoTBMi+phecjLE4KV0vORccLyIenwb78iBhYrMryNIpcPQ9SCEk5i55WgmmRtb5z5jYBLbWGMs
XdhvT74OfcIcjHWdb3O8zuyJnt69fMOSPlQD6dgmg4ebqAnaHfaFR9lB+RTpHMMQmwKK7Gx9/Qfu
I0tn9mEx9sYRDIUIge3+pM55jEjU5hQKjFYgFKIxOhMAPpYpPWAgKAOwC6TXarEjoc+q5QwKROL+
7tSBTKfw4NRq0RyAUYJaUl8RLKs6pSxGnCuGfHRdxdtmRu7VhywH3wI++o49u4Z0LHv9sAGkpxUq
560GQp+bWD8KNtJKNyN7BpKbzPryopIUju6YOs7wktLgF4WdhsvfCmYr3ZifbgrEmjlKjCbKSCfC
nOUjhVdT/U3TNGfdnqzaC7dS4BGpCw07QCtJIbGnQ7KgqmpaRq9mB+OlPJwwAocxs7c9zk8+blY8
cFWYGxbiEfvcRP+VPdb28vXxmkx/sYnKxZq9XiQghZ5O9JMvlV1a1LJQ1Bdrwxgm/E9SjHmZR3t4
4VqMKgP8JUMIcaPG73CTQ3nuU1D50xeAdPCxjrdJ9nNBCfOwL4AXhnSTkNoFDL+0jkl/MMeZWA3T
XqRd15NiciwfslWjIvsTJIwZy8hLCgKCpMEetEu/IGVs7fQJvDvgEicPnpO7gllqLgnaoVev5Cvv
XV+IM83TcnkDH7NO6NM+doa3+n9ZcJLTlrE2xD+P5UzhOt/o1Vf8374ue+Z8pNCJ+iT9cRIF4J/2
KMXbf7PTW6kuQl5E0Pz40lPakBDgiUFegJVdtaOutOFlP6aG+OJNgfBTISnZZ05My++qzXcdavAA
6J4j7E/x4gbx0O7P+Lx8rlInLvXdXqGGoyeKIwu/v8Cd1Vlh3GP9hJ/w4J1/rUfbfBDhhi5xCSMV
hwWyIRSuAQtO0N7vi339amcdhPtKCZkqHGY+yP9FlhPwETVqFOwZBE+0Q8xB0HKb7pARcHV11uFu
YLWICIbeeDhNMoEZhRb3vkLdid6a7SZ5txHWs1NXCY8j1y9awEgEhhtHYRkJg11fhDTHkH2YWd6W
2aRJBixsYkKZFFecKTFJTAD4vEgpPJBtclWKdH2wvq93ewB5z5y0nEWYnyIqm6XzfUvguM14b40l
i3iQdzJkHKvy1dTq/S0ry0zwXcRDjEiq1dtdcNOdsFeYcDbiIj3fi89GCyb6P61wL+qJQANHxDVR
PAKBAT11Im5lcdWpQsHc5ranTpJ5TZK9xbu20RG019Ru/whmt18pKBihED6khCAtaBgE2PufnPiE
DqWeW625H+iIO2uG3qMz8s+WHW4SBxsIz7nabVxpdhqesSE0SbcmcQnpsOBsba6gRYv1Lbzum1/g
twaUgVyczMIslkuwQCWGTP6igzLzQg+k8SWW9f89MIDkC9RJ5KSJplSPlgLEiyRgFuPwpc2aqC5f
N5Qv6zuYiRqNngAc0l8p3ajBQvvg6uWXnLbgYQ2+SUUoin+ZpS5pSobGTZ3i8Hx8C89RHVHOLY37
fvz5gXlXOGiUp+7yT/5dvdIRGrZvH4JkLU3BWh+Bd3hSQvI995hcuRSmDbmClsTtwhEBHgLB/Xin
63ZLA880shp/cAg5JOHomlftfUpWbKJFOfju5OOD2cIr28WP2xiYro38Wfdh3fuzPm7PYIxBxDIm
ZMfBEQXBiKiFOqadGroHR9Vn9nIoafv9HIYgEkVQNaK/UhpnKnzAphuWGHec9G0mQ1t32MDMQB3F
VtO3MF3m9Of4wBdji+nhszOI89EuylCs4L1qOeiD6b23PEMmodtwGNMb0K8ilPPBtOlykqVn9bA5
iOO0iYuJReqC9gNj7syTcBSZUn38GAJ4jPu6yaJncv1Ac/RKNmOrMRGaZG+tpkoCkPKxq+CHkHoY
j35nPcGSLIumMk4P5dkLujv5UJV3dRgOAubIUHrDNf7Y54T9rQbN8c5Byf9G2FIVg+dJN4CL1WkC
8aQ8thMI6aNeQbFpOX1/aApQP/5v1B3MrS3egFQpVRwF4zk2RAWvr/8qVy1t5IrWLsgK32jbSCDs
BZ4GUxlRUcl+d9y2T33bsbnVfOXlkhxP9xBa6x0UzL1NneOPo6Dug//EGoVfblU76DJz1EmG19bj
P+f4Qv0rsfJDYIIVN7GhshJHbzpqGlW59F1PZtzOTNuzFYeGf6m3FYePaxjYM/plVFdjZjryrQal
oCE5pkaysuLm169rhZ95x99NeOzuOK2Vq1gWmj7rQlHr9n+lVxmNNWiBZzAPzkt8hELwAbPOaf5H
nQE9rxAEIyMtTodneRp8f5CJFEE3vpnLxEPjD7exERgDT6ytAYe77DqnaMpYcQH5m14jf570z/Xn
XmTqFA0I61qaAwoDqydz2tLzTCWJm9L+wWcxJcpcAKNY
`protect end_protected
